module basic_5000_50000_5000_200_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_1202,In_399);
and U1 (N_1,In_9,In_141);
nand U2 (N_2,In_743,In_2228);
or U3 (N_3,In_145,In_2757);
nor U4 (N_4,In_608,In_3288);
and U5 (N_5,In_3645,In_81);
nand U6 (N_6,In_3714,In_4282);
nand U7 (N_7,In_2733,In_477);
or U8 (N_8,In_2261,In_325);
nor U9 (N_9,In_4559,In_719);
xnor U10 (N_10,In_494,In_1639);
nor U11 (N_11,In_4741,In_3024);
nor U12 (N_12,In_1729,In_4830);
nand U13 (N_13,In_2529,In_3831);
nand U14 (N_14,In_4272,In_4325);
and U15 (N_15,In_1295,In_3346);
nor U16 (N_16,In_3196,In_2346);
and U17 (N_17,In_2575,In_4350);
and U18 (N_18,In_869,In_2643);
xnor U19 (N_19,In_3194,In_1293);
nand U20 (N_20,In_2353,In_3495);
or U21 (N_21,In_3965,In_2125);
xor U22 (N_22,In_3870,In_3300);
or U23 (N_23,In_2775,In_4307);
nor U24 (N_24,In_4194,In_152);
nand U25 (N_25,In_1890,In_1327);
nor U26 (N_26,In_2738,In_1269);
xor U27 (N_27,In_2622,In_4806);
or U28 (N_28,In_4757,In_2595);
nor U29 (N_29,In_3486,In_863);
nor U30 (N_30,In_2914,In_2662);
and U31 (N_31,In_4062,In_4509);
and U32 (N_32,In_3999,In_1065);
xnor U33 (N_33,In_1466,In_740);
nand U34 (N_34,In_4820,In_3268);
or U35 (N_35,In_617,In_1152);
nand U36 (N_36,In_4858,In_3096);
xnor U37 (N_37,In_435,In_3215);
and U38 (N_38,In_4175,In_4635);
or U39 (N_39,In_8,In_2634);
or U40 (N_40,In_2967,In_1740);
and U41 (N_41,In_561,In_378);
or U42 (N_42,In_653,In_4122);
nor U43 (N_43,In_106,In_4640);
or U44 (N_44,In_1346,In_718);
and U45 (N_45,In_1881,In_4156);
or U46 (N_46,In_4823,In_3287);
nand U47 (N_47,In_3200,In_1785);
xnor U48 (N_48,In_1161,In_4026);
and U49 (N_49,In_4021,In_3542);
nand U50 (N_50,In_1811,In_4440);
or U51 (N_51,In_2908,In_3158);
nand U52 (N_52,In_1587,In_4412);
or U53 (N_53,In_2688,In_2838);
xnor U54 (N_54,In_1220,In_2416);
or U55 (N_55,In_842,In_3626);
nand U56 (N_56,In_3572,In_4643);
and U57 (N_57,In_409,In_3849);
nand U58 (N_58,In_1406,In_2601);
and U59 (N_59,In_4956,In_1929);
nand U60 (N_60,In_4117,In_303);
or U61 (N_61,In_4489,In_1681);
nand U62 (N_62,In_926,In_3858);
or U63 (N_63,In_1362,In_4653);
or U64 (N_64,In_3104,In_151);
and U65 (N_65,In_1433,In_3208);
xor U66 (N_66,In_4336,In_3140);
xor U67 (N_67,In_2611,In_4925);
nand U68 (N_68,In_4873,In_1781);
or U69 (N_69,In_2322,In_60);
nand U70 (N_70,In_788,In_1252);
and U71 (N_71,In_3253,In_1786);
nor U72 (N_72,In_3769,In_4472);
nor U73 (N_73,In_3796,In_2997);
or U74 (N_74,In_1492,In_4096);
nand U75 (N_75,In_1809,In_1463);
nand U76 (N_76,In_3226,In_3129);
or U77 (N_77,In_958,In_252);
and U78 (N_78,In_4700,In_997);
and U79 (N_79,In_4153,In_1550);
xnor U80 (N_80,In_1725,In_1808);
nand U81 (N_81,In_263,In_520);
nand U82 (N_82,In_2909,In_4362);
or U83 (N_83,In_3808,In_868);
and U84 (N_84,In_573,In_3247);
or U85 (N_85,In_1084,In_1619);
xnor U86 (N_86,In_4373,In_921);
xor U87 (N_87,In_401,In_4543);
and U88 (N_88,In_4248,In_620);
and U89 (N_89,In_3321,In_4326);
nand U90 (N_90,In_3939,In_742);
or U91 (N_91,In_4620,In_3243);
nor U92 (N_92,In_2404,In_3970);
and U93 (N_93,In_2603,In_4345);
and U94 (N_94,In_496,In_1966);
and U95 (N_95,In_3940,In_4014);
xnor U96 (N_96,In_2717,In_3005);
xor U97 (N_97,In_4384,In_1902);
nand U98 (N_98,In_4475,In_4482);
nor U99 (N_99,In_4526,In_1170);
and U100 (N_100,In_4538,In_3976);
nand U101 (N_101,In_2397,In_4797);
nand U102 (N_102,In_2396,In_2823);
xor U103 (N_103,In_2459,In_3314);
nand U104 (N_104,In_173,In_922);
or U105 (N_105,In_4042,In_3925);
xnor U106 (N_106,In_4708,In_3441);
xnor U107 (N_107,In_2441,In_1634);
and U108 (N_108,In_1381,In_4285);
and U109 (N_109,In_691,In_1903);
xor U110 (N_110,In_567,In_952);
and U111 (N_111,In_3905,In_4805);
or U112 (N_112,In_3582,In_887);
nor U113 (N_113,In_1916,In_3618);
nor U114 (N_114,In_119,In_4340);
xor U115 (N_115,In_2911,In_1410);
nor U116 (N_116,In_1880,In_2624);
nand U117 (N_117,In_2319,In_4651);
nor U118 (N_118,In_3012,In_877);
nand U119 (N_119,In_351,In_3595);
nor U120 (N_120,In_1561,In_3340);
nand U121 (N_121,In_3139,In_625);
xor U122 (N_122,In_2537,In_3260);
or U123 (N_123,In_4680,In_4353);
nand U124 (N_124,In_2916,In_983);
and U125 (N_125,In_3900,In_1037);
or U126 (N_126,In_787,In_3952);
nand U127 (N_127,In_965,In_513);
nand U128 (N_128,In_4693,In_506);
nand U129 (N_129,In_4106,In_3931);
xnor U130 (N_130,In_916,In_1008);
or U131 (N_131,In_2067,In_3025);
and U132 (N_132,In_3074,In_4841);
and U133 (N_133,In_32,In_1913);
nor U134 (N_134,In_2850,In_2379);
nand U135 (N_135,In_3275,In_4317);
xnor U136 (N_136,In_4990,In_4075);
or U137 (N_137,In_3732,In_4138);
nand U138 (N_138,In_431,In_4267);
xnor U139 (N_139,In_4675,In_1366);
nand U140 (N_140,In_1219,In_1520);
nand U141 (N_141,In_4608,In_4623);
and U142 (N_142,In_2704,In_1479);
and U143 (N_143,In_4807,In_2273);
and U144 (N_144,In_4828,In_977);
nor U145 (N_145,In_3010,In_153);
nand U146 (N_146,In_4533,In_3592);
or U147 (N_147,In_3701,In_4560);
or U148 (N_148,In_2267,In_3118);
and U149 (N_149,In_1883,In_4006);
and U150 (N_150,In_370,In_97);
and U151 (N_151,In_2479,In_2072);
and U152 (N_152,In_3446,In_1280);
or U153 (N_153,In_2150,In_4595);
and U154 (N_154,In_489,In_4392);
and U155 (N_155,In_3812,In_3865);
xor U156 (N_156,In_1595,In_1566);
xor U157 (N_157,In_1950,In_2526);
nor U158 (N_158,In_2071,In_3765);
nor U159 (N_159,In_2034,In_269);
nor U160 (N_160,In_1073,In_71);
nand U161 (N_161,In_1245,In_3202);
and U162 (N_162,In_4212,In_2138);
nor U163 (N_163,In_2922,In_2571);
xnor U164 (N_164,In_4637,In_1979);
nor U165 (N_165,In_1649,In_643);
nor U166 (N_166,In_1558,In_4647);
nor U167 (N_167,In_586,In_2556);
and U168 (N_168,In_2776,In_3424);
and U169 (N_169,In_1545,In_936);
nand U170 (N_170,In_3710,In_4327);
and U171 (N_171,In_637,In_4419);
or U172 (N_172,In_3407,In_3033);
or U173 (N_173,In_3046,In_2184);
nor U174 (N_174,In_2936,In_1849);
or U175 (N_175,In_4203,In_3088);
xor U176 (N_176,In_2395,In_1792);
nor U177 (N_177,In_192,In_2790);
or U178 (N_178,In_2844,In_1666);
or U179 (N_179,In_4984,In_309);
or U180 (N_180,In_1713,In_3415);
and U181 (N_181,In_2992,In_451);
xnor U182 (N_182,In_1272,In_1872);
and U183 (N_183,In_2263,In_4468);
nor U184 (N_184,In_2149,In_3459);
and U185 (N_185,In_377,In_3772);
nor U186 (N_186,In_2166,In_3357);
or U187 (N_187,In_2094,In_4044);
and U188 (N_188,In_254,In_4594);
xnor U189 (N_189,In_2123,In_834);
xnor U190 (N_190,In_4793,In_3944);
nor U191 (N_191,In_2028,In_3277);
and U192 (N_192,In_2308,In_4306);
xor U193 (N_193,In_480,In_246);
or U194 (N_194,In_100,In_2075);
nand U195 (N_195,In_3949,In_4737);
xor U196 (N_196,In_2950,In_2927);
or U197 (N_197,In_4907,In_1186);
nand U198 (N_198,In_883,In_4020);
nor U199 (N_199,In_3623,In_4657);
or U200 (N_200,In_3453,In_701);
nand U201 (N_201,In_4865,In_1006);
nand U202 (N_202,In_739,In_1428);
xnor U203 (N_203,In_4439,In_1045);
nor U204 (N_204,In_471,In_4047);
or U205 (N_205,In_4545,In_1648);
nor U206 (N_206,In_4527,In_4866);
xnor U207 (N_207,In_281,In_410);
or U208 (N_208,In_1657,In_4069);
nand U209 (N_209,In_3210,In_402);
nor U210 (N_210,In_2439,In_1047);
nor U211 (N_211,In_2700,In_2709);
xor U212 (N_212,In_2248,In_1958);
xor U213 (N_213,In_3670,In_367);
or U214 (N_214,In_3768,In_3479);
and U215 (N_215,In_1175,In_4137);
nand U216 (N_216,In_2943,In_1565);
nand U217 (N_217,In_3455,In_4920);
nor U218 (N_218,In_3803,In_2367);
or U219 (N_219,In_4132,In_1503);
nor U220 (N_220,In_4239,In_1231);
nor U221 (N_221,In_2793,In_4981);
xor U222 (N_222,In_735,In_4279);
xor U223 (N_223,In_1771,In_3122);
xor U224 (N_224,In_3295,In_1691);
nor U225 (N_225,In_2581,In_1167);
nor U226 (N_226,In_2951,In_2120);
or U227 (N_227,In_3169,In_2314);
nor U228 (N_228,In_4556,In_3876);
nor U229 (N_229,In_486,In_4729);
nor U230 (N_230,In_3004,In_1744);
and U231 (N_231,In_999,In_4324);
nand U232 (N_232,In_4958,In_4931);
xnor U233 (N_233,In_2989,In_4293);
nor U234 (N_234,In_3085,In_3334);
or U235 (N_235,In_3270,In_4750);
nand U236 (N_236,In_2630,In_3536);
and U237 (N_237,In_2767,In_2270);
and U238 (N_238,In_3912,In_923);
and U239 (N_239,In_4150,In_1640);
and U240 (N_240,In_955,In_644);
xnor U241 (N_241,In_4682,In_1533);
and U242 (N_242,In_1931,In_4867);
and U243 (N_243,In_3037,In_1304);
nand U244 (N_244,In_1456,In_2186);
xor U245 (N_245,In_3190,In_3390);
xor U246 (N_246,In_1350,In_1723);
or U247 (N_247,In_1995,In_3339);
or U248 (N_248,In_1342,In_4663);
xor U249 (N_249,In_2904,In_4844);
nand U250 (N_250,In_3629,In_3365);
nand U251 (N_251,In_4689,In_4374);
or U252 (N_252,In_1993,N_81);
or U253 (N_253,In_3678,In_4963);
or U254 (N_254,In_2074,In_178);
nand U255 (N_255,In_660,In_1412);
xnor U256 (N_256,N_245,In_2430);
xor U257 (N_257,In_4056,In_2369);
nand U258 (N_258,In_1394,In_3475);
nand U259 (N_259,In_1090,In_4518);
or U260 (N_260,In_213,In_2583);
or U261 (N_261,In_2198,In_3452);
or U262 (N_262,In_1961,In_884);
nand U263 (N_263,In_4234,N_68);
nor U264 (N_264,In_2415,In_3754);
nand U265 (N_265,In_4762,In_3615);
xnor U266 (N_266,N_220,In_3972);
nand U267 (N_267,In_3432,In_110);
or U268 (N_268,In_476,In_4731);
or U269 (N_269,In_1338,In_2057);
nor U270 (N_270,In_1130,In_2910);
or U271 (N_271,N_51,In_631);
nor U272 (N_272,In_1548,In_3638);
nor U273 (N_273,In_3738,In_1821);
and U274 (N_274,In_1353,In_2500);
xnor U275 (N_275,In_10,In_1340);
and U276 (N_276,In_659,In_1651);
or U277 (N_277,In_2582,N_99);
or U278 (N_278,In_2932,In_4230);
nand U279 (N_279,In_449,In_2532);
and U280 (N_280,In_1116,In_3955);
xor U281 (N_281,In_3862,In_712);
nor U282 (N_282,In_789,N_25);
nand U283 (N_283,In_873,N_142);
nor U284 (N_284,In_4095,In_230);
xnor U285 (N_285,In_3651,In_4494);
and U286 (N_286,In_1114,In_1605);
nor U287 (N_287,In_4783,In_4583);
or U288 (N_288,In_2168,In_3863);
and U289 (N_289,In_698,In_2533);
and U290 (N_290,In_4114,In_2117);
xnor U291 (N_291,In_3628,In_2035);
nor U292 (N_292,In_1398,In_3576);
and U293 (N_293,In_4849,In_3977);
or U294 (N_294,In_612,In_2938);
xor U295 (N_295,In_2751,In_389);
xnor U296 (N_296,In_3204,In_3050);
and U297 (N_297,In_3241,In_1076);
nand U298 (N_298,In_3434,In_432);
nor U299 (N_299,In_2955,In_380);
xor U300 (N_300,In_3119,In_1064);
or U301 (N_301,In_4514,In_4786);
and U302 (N_302,In_1516,In_1095);
nand U303 (N_303,In_2562,In_969);
nand U304 (N_304,In_3347,N_227);
nand U305 (N_305,In_198,In_4032);
nor U306 (N_306,In_3750,In_4207);
nor U307 (N_307,In_2987,In_1180);
or U308 (N_308,In_208,In_210);
nor U309 (N_309,In_4935,In_1042);
xnor U310 (N_310,N_66,In_615);
xor U311 (N_311,In_2313,In_3286);
nand U312 (N_312,In_1329,In_1486);
nor U313 (N_313,In_4109,In_1816);
xnor U314 (N_314,In_1782,In_2392);
and U315 (N_315,In_3837,In_2082);
nand U316 (N_316,In_1305,In_3668);
or U317 (N_317,In_316,In_1275);
or U318 (N_318,In_1759,In_2543);
nand U319 (N_319,In_2464,In_4537);
or U320 (N_320,In_1920,In_314);
nor U321 (N_321,In_2093,In_751);
nand U322 (N_322,In_4268,In_1633);
nor U323 (N_323,In_3507,In_3117);
xor U324 (N_324,In_2015,In_1221);
and U325 (N_325,In_4201,In_2716);
and U326 (N_326,In_3724,In_1154);
nor U327 (N_327,In_301,N_226);
or U328 (N_328,In_2818,In_2307);
nor U329 (N_329,In_4582,In_3396);
xor U330 (N_330,In_4423,In_4691);
xnor U331 (N_331,In_2458,In_3587);
nor U332 (N_332,In_1457,In_556);
and U333 (N_333,In_4342,In_4474);
xnor U334 (N_334,In_2788,In_1235);
xor U335 (N_335,In_3648,In_1915);
xor U336 (N_336,N_76,In_3378);
nor U337 (N_337,In_3580,In_3218);
nand U338 (N_338,In_3249,In_4435);
or U339 (N_339,In_2390,In_4536);
nor U340 (N_340,In_2323,In_3419);
xor U341 (N_341,In_663,In_63);
or U342 (N_342,In_1549,In_396);
or U343 (N_343,In_3687,In_2465);
and U344 (N_344,In_4186,In_3265);
or U345 (N_345,In_1779,In_12);
xor U346 (N_346,In_4800,In_484);
nor U347 (N_347,In_2453,In_1306);
or U348 (N_348,In_4804,In_639);
nor U349 (N_349,In_4829,In_3634);
xor U350 (N_350,In_2437,In_582);
nor U351 (N_351,In_3822,In_811);
xor U352 (N_352,N_133,In_2640);
or U353 (N_353,In_4798,In_4980);
and U354 (N_354,N_84,In_2229);
xnor U355 (N_355,In_716,In_2670);
or U356 (N_356,In_326,N_79);
xnor U357 (N_357,In_382,In_2447);
xnor U358 (N_358,In_387,In_4396);
xnor U359 (N_359,In_3502,In_4055);
or U360 (N_360,In_4181,In_2868);
and U361 (N_361,In_3211,In_959);
nor U362 (N_362,In_836,In_2427);
nand U363 (N_363,In_2940,In_2631);
nand U364 (N_364,In_1465,In_1504);
nor U365 (N_365,In_2328,In_2244);
nor U366 (N_366,In_4781,In_2320);
or U367 (N_367,In_4483,In_3351);
xnor U368 (N_368,In_1528,N_180);
xor U369 (N_369,In_4037,In_4975);
or U370 (N_370,In_2480,In_4826);
or U371 (N_371,In_754,In_894);
nor U372 (N_372,In_3319,In_4053);
nor U373 (N_373,In_914,In_3108);
nor U374 (N_374,In_2121,In_2118);
nand U375 (N_375,In_4270,In_4219);
xnor U376 (N_376,In_4398,In_488);
or U377 (N_377,In_3983,In_2252);
or U378 (N_378,In_4774,In_705);
or U379 (N_379,In_2217,In_1761);
or U380 (N_380,In_890,In_395);
and U381 (N_381,In_4889,In_553);
nand U382 (N_382,In_3379,In_1214);
xor U383 (N_383,In_893,In_3105);
nand U384 (N_384,In_3369,In_1320);
or U385 (N_385,In_2663,In_176);
nand U386 (N_386,N_108,In_3761);
nor U387 (N_387,In_1795,In_2745);
nor U388 (N_388,In_1276,In_2451);
nor U389 (N_389,In_2029,In_3568);
nor U390 (N_390,In_293,In_544);
and U391 (N_391,In_262,In_3951);
and U392 (N_392,In_4128,In_4111);
or U393 (N_393,In_3094,In_183);
or U394 (N_394,In_645,In_3857);
or U395 (N_395,In_1420,In_4579);
and U396 (N_396,In_1249,In_4308);
xor U397 (N_397,In_1029,In_2608);
nand U398 (N_398,In_1877,In_3708);
or U399 (N_399,In_1974,In_4961);
xor U400 (N_400,In_2064,In_23);
nand U401 (N_401,In_3233,In_741);
nand U402 (N_402,In_134,In_610);
nand U403 (N_403,In_624,In_2735);
nor U404 (N_404,In_522,In_1091);
xor U405 (N_405,In_2664,In_3234);
and U406 (N_406,In_2220,In_1604);
nor U407 (N_407,N_212,In_1527);
xnor U408 (N_408,In_1685,In_1793);
or U409 (N_409,In_2463,In_2902);
nand U410 (N_410,In_3707,In_1449);
nand U411 (N_411,In_1259,In_1341);
xor U412 (N_412,In_2905,In_3462);
and U413 (N_413,In_3942,In_3349);
and U414 (N_414,In_89,N_202);
or U415 (N_415,In_1375,In_2185);
xor U416 (N_416,In_4170,In_4086);
nand U417 (N_417,In_3526,In_1142);
or U418 (N_418,In_2301,In_4546);
or U419 (N_419,In_4957,In_2829);
nor U420 (N_420,In_448,In_264);
or U421 (N_421,In_2888,In_284);
nand U422 (N_422,In_1970,In_3516);
or U423 (N_423,In_3700,In_606);
xor U424 (N_424,In_1424,In_80);
or U425 (N_425,In_3132,In_130);
and U426 (N_426,In_4744,N_11);
nand U427 (N_427,In_722,In_2178);
xnor U428 (N_428,In_186,In_1203);
xor U429 (N_429,In_1311,In_3429);
nor U430 (N_430,In_492,In_831);
and U431 (N_431,In_4463,In_2059);
xor U432 (N_432,In_3842,In_3000);
nand U433 (N_433,In_2930,In_2632);
and U434 (N_434,In_1956,In_1952);
nand U435 (N_435,In_4955,In_4706);
nor U436 (N_436,In_193,In_4993);
nand U437 (N_437,In_696,N_214);
nand U438 (N_438,In_4742,In_1171);
or U439 (N_439,In_2633,In_752);
nor U440 (N_440,In_3603,In_2782);
xnor U441 (N_441,In_508,In_4681);
xor U442 (N_442,In_1331,In_1544);
nand U443 (N_443,In_2771,In_662);
and U444 (N_444,In_3272,In_534);
nor U445 (N_445,In_2363,In_2351);
xnor U446 (N_446,In_4195,In_4502);
or U447 (N_447,In_3709,In_3292);
nor U448 (N_448,In_1495,In_3672);
nand U449 (N_449,In_4211,In_4283);
xnor U450 (N_450,In_3305,In_986);
nor U451 (N_451,In_2187,In_1172);
xor U452 (N_452,In_2510,In_3399);
nor U453 (N_453,In_1546,In_2045);
xor U454 (N_454,In_771,In_2901);
nor U455 (N_455,In_988,In_4415);
and U456 (N_456,In_621,In_2903);
nor U457 (N_457,In_1325,In_3177);
and U458 (N_458,In_1236,In_930);
nand U459 (N_459,In_3671,In_3728);
xor U460 (N_460,In_3820,In_1317);
or U461 (N_461,In_4262,In_3515);
nand U462 (N_462,In_3066,N_63);
nor U463 (N_463,In_565,In_979);
and U464 (N_464,In_629,N_177);
and U465 (N_465,In_1144,In_3815);
or U466 (N_466,In_4102,In_2488);
nor U467 (N_467,In_3072,In_3593);
nand U468 (N_468,In_911,In_4238);
nand U469 (N_469,In_1517,In_2249);
xnor U470 (N_470,In_1498,In_3236);
or U471 (N_471,In_487,In_3408);
xnor U472 (N_472,In_390,In_1836);
nand U473 (N_473,In_3280,In_3763);
nor U474 (N_474,In_730,In_3376);
nand U475 (N_475,In_4408,In_3715);
or U476 (N_476,In_1025,In_4531);
nor U477 (N_477,In_4944,In_4411);
xnor U478 (N_478,In_4382,In_4924);
nand U479 (N_479,In_3731,In_3644);
or U480 (N_480,In_4512,In_1923);
or U481 (N_481,In_2552,In_1351);
nand U482 (N_482,In_1885,In_1616);
or U483 (N_483,In_2509,In_22);
nand U484 (N_484,In_2981,In_667);
nand U485 (N_485,In_2722,In_2063);
or U486 (N_486,In_218,In_1308);
or U487 (N_487,In_2344,In_1906);
xor U488 (N_488,In_3303,In_1513);
nand U489 (N_489,In_1896,In_3929);
nor U490 (N_490,In_690,In_4261);
xnor U491 (N_491,In_3464,In_3049);
nor U492 (N_492,In_4455,In_2389);
nor U493 (N_493,In_1113,In_3789);
nand U494 (N_494,In_545,In_3637);
or U495 (N_495,In_2553,In_2666);
and U496 (N_496,N_140,In_2499);
nor U497 (N_497,In_3945,In_4602);
nor U498 (N_498,In_2680,In_3581);
nand U499 (N_499,In_3690,In_2193);
and U500 (N_500,In_3248,N_432);
nand U501 (N_501,In_69,In_3913);
and U502 (N_502,In_2294,In_475);
nand U503 (N_503,In_2159,In_274);
nand U504 (N_504,In_4557,In_4550);
xnor U505 (N_505,In_3666,N_157);
and U506 (N_506,In_1011,In_4566);
nor U507 (N_507,N_497,N_60);
nor U508 (N_508,In_4257,In_1244);
or U509 (N_509,In_1717,In_4809);
xnor U510 (N_510,In_4292,In_1508);
or U511 (N_511,N_364,N_406);
xnor U512 (N_512,In_1763,In_289);
nand U513 (N_513,In_987,In_1963);
and U514 (N_514,N_457,In_951);
xnor U515 (N_515,In_4591,In_4456);
and U516 (N_516,In_2491,In_3722);
nand U517 (N_517,N_33,In_3720);
and U518 (N_518,In_2276,N_104);
nor U519 (N_519,In_535,N_424);
or U520 (N_520,In_3219,In_111);
xor U521 (N_521,In_3839,In_3834);
nand U522 (N_522,In_1611,N_138);
and U523 (N_523,In_973,In_250);
xnor U524 (N_524,In_1756,In_589);
xor U525 (N_525,In_1297,In_552);
and U526 (N_526,In_4876,In_2505);
nand U527 (N_527,In_2516,In_1436);
xnor U528 (N_528,In_4810,In_2519);
or U529 (N_529,In_3167,In_4490);
or U530 (N_530,In_4399,In_282);
nor U531 (N_531,In_4316,In_2160);
or U532 (N_532,In_2817,In_3392);
and U533 (N_533,In_2675,In_1388);
or U534 (N_534,In_379,In_4376);
xnor U535 (N_535,In_3427,In_3696);
nor U536 (N_536,In_2784,N_264);
nand U537 (N_537,In_4420,In_1898);
nand U538 (N_538,In_3206,In_2317);
nor U539 (N_539,In_2941,In_148);
and U540 (N_540,In_1129,In_2796);
xnor U541 (N_541,In_185,In_1910);
xnor U542 (N_542,In_2669,In_3142);
nand U543 (N_543,In_2254,In_1538);
nand U544 (N_544,In_2142,In_255);
xor U545 (N_545,In_3620,In_630);
nand U546 (N_546,In_2890,In_3316);
xnor U547 (N_547,N_454,N_383);
nor U548 (N_548,N_330,N_125);
or U549 (N_549,In_2147,In_2030);
xnor U550 (N_550,In_3450,In_90);
and U551 (N_551,In_1086,In_3783);
nor U552 (N_552,In_4365,In_776);
and U553 (N_553,In_30,N_178);
xnor U554 (N_554,In_773,In_1695);
nand U555 (N_555,In_4298,In_4157);
nand U556 (N_556,In_4617,In_1738);
or U557 (N_557,In_2754,N_95);
and U558 (N_558,In_3604,In_350);
or U559 (N_559,In_369,In_1873);
nand U560 (N_560,In_862,In_3162);
nand U561 (N_561,In_4254,In_4917);
nand U562 (N_562,In_3213,In_3126);
and U563 (N_563,In_1482,In_3133);
and U564 (N_564,In_53,In_165);
and U565 (N_565,N_283,In_2703);
xor U566 (N_566,In_1983,In_4159);
nor U567 (N_567,In_510,In_4904);
or U568 (N_568,In_3673,In_4346);
nor U569 (N_569,In_2656,In_374);
xor U570 (N_570,In_3967,In_3416);
xnor U571 (N_571,In_3688,In_2756);
xnor U572 (N_572,N_472,In_4329);
xor U573 (N_573,In_4210,N_421);
nand U574 (N_574,In_191,In_1053);
or U575 (N_575,In_3082,In_2058);
or U576 (N_576,In_1692,In_1718);
nor U577 (N_577,In_3461,In_2176);
nand U578 (N_578,In_1960,In_3310);
nor U579 (N_579,In_2194,N_389);
nor U580 (N_580,In_1572,In_227);
nand U581 (N_581,In_1474,In_2697);
and U582 (N_582,In_2226,In_1435);
nand U583 (N_583,In_2858,N_209);
nand U584 (N_584,In_577,In_40);
or U585 (N_585,In_4467,In_2163);
nor U586 (N_586,In_728,In_947);
nor U587 (N_587,In_1030,In_2098);
and U588 (N_588,In_2760,In_450);
nand U589 (N_589,In_4510,In_485);
xnor U590 (N_590,In_4728,In_4252);
or U591 (N_591,In_300,In_4906);
xor U592 (N_592,In_4480,In_745);
or U593 (N_593,N_388,In_3633);
nor U594 (N_594,In_2302,In_1984);
and U595 (N_595,In_3343,In_4795);
nand U596 (N_596,In_3570,In_3180);
xor U597 (N_597,In_3546,In_2894);
xor U598 (N_598,In_344,In_4125);
and U599 (N_599,In_2189,In_2420);
or U600 (N_600,In_2218,In_459);
xor U601 (N_601,In_2001,In_3797);
nand U602 (N_602,In_3589,In_3788);
nand U603 (N_603,In_3602,In_3959);
nand U604 (N_604,In_3988,In_6);
and U605 (N_605,In_4430,N_211);
nor U606 (N_606,In_1878,N_373);
xor U607 (N_607,In_2152,In_3745);
or U608 (N_608,In_4241,In_767);
and U609 (N_609,N_122,In_3641);
or U610 (N_610,In_4260,In_28);
xnor U611 (N_611,In_190,In_2802);
nor U612 (N_612,In_3775,In_658);
and U613 (N_613,In_4355,In_2915);
nand U614 (N_614,In_692,In_4683);
and U615 (N_615,In_593,In_1753);
xor U616 (N_616,In_4083,In_1467);
xnor U617 (N_617,In_2988,N_416);
nor U618 (N_618,In_4972,In_1447);
nor U619 (N_619,In_3987,In_4803);
or U620 (N_620,In_3622,N_273);
xor U621 (N_621,N_469,In_4041);
or U622 (N_622,In_2215,In_3908);
nor U623 (N_623,In_2321,In_744);
xor U624 (N_624,In_4438,In_1074);
or U625 (N_625,In_3361,In_1564);
nor U626 (N_626,In_3506,In_4734);
nor U627 (N_627,In_1328,N_24);
or U628 (N_628,In_3907,N_162);
or U629 (N_629,In_3727,In_253);
nand U630 (N_630,In_1636,In_1489);
xor U631 (N_631,In_1628,In_472);
xnor U632 (N_632,In_3543,In_4661);
and U633 (N_633,In_182,In_2102);
nor U634 (N_634,In_4577,In_4414);
nor U635 (N_635,In_3729,In_2612);
nand U636 (N_636,In_4050,In_2973);
nand U637 (N_637,In_2618,N_413);
nor U638 (N_638,In_4046,In_2655);
or U639 (N_639,In_3428,N_159);
nand U640 (N_640,In_2821,In_4878);
xor U641 (N_641,In_1364,In_2378);
nor U642 (N_642,In_2277,In_1669);
nand U643 (N_643,In_2460,In_880);
or U644 (N_644,N_186,In_1374);
nand U645 (N_645,N_310,In_2288);
xnor U646 (N_646,In_113,N_363);
or U647 (N_647,In_1442,In_3843);
and U648 (N_648,In_41,In_302);
nor U649 (N_649,In_3293,In_126);
and U650 (N_650,In_4982,In_1036);
and U651 (N_651,N_272,In_2180);
nand U652 (N_652,In_4937,In_4466);
xnor U653 (N_653,In_3156,In_327);
nand U654 (N_654,In_4187,In_4129);
nor U655 (N_655,In_4233,In_4530);
nand U656 (N_656,In_2763,In_415);
or U657 (N_657,In_2848,In_3792);
nor U658 (N_658,In_442,In_1677);
or U659 (N_659,In_461,In_4667);
xor U660 (N_660,In_678,In_1404);
nand U661 (N_661,In_4066,In_3125);
nor U662 (N_662,N_13,In_618);
nor U663 (N_663,In_3578,In_4013);
nor U664 (N_664,In_56,In_2171);
nor U665 (N_665,In_2213,In_88);
nand U666 (N_666,In_2535,In_4771);
nor U667 (N_667,In_440,N_324);
nand U668 (N_668,In_3498,In_2820);
xnor U669 (N_669,In_3494,In_3971);
nand U670 (N_670,In_1062,N_5);
and U671 (N_671,In_2100,In_991);
nor U672 (N_672,In_3847,In_3779);
and U673 (N_673,In_4223,In_4303);
or U674 (N_674,In_2157,In_906);
and U675 (N_675,In_3212,In_1376);
and U676 (N_676,In_2843,In_502);
or U677 (N_677,In_4847,In_2484);
xor U678 (N_678,In_4900,In_1299);
and U679 (N_679,In_4246,N_279);
nor U680 (N_680,In_2673,In_2474);
nor U681 (N_681,In_1163,In_3302);
and U682 (N_682,In_772,In_1143);
and U683 (N_683,In_128,In_4286);
or U684 (N_684,In_2900,In_3123);
xnor U685 (N_685,In_1948,In_93);
nand U686 (N_686,In_4085,In_2620);
xor U687 (N_687,In_116,In_4130);
nand U688 (N_688,In_3996,In_849);
or U689 (N_689,In_481,N_153);
nand U690 (N_690,In_3047,In_1614);
nor U691 (N_691,In_4843,In_1372);
xnor U692 (N_692,In_804,In_3652);
and U693 (N_693,In_47,In_3313);
and U694 (N_694,In_2544,In_4017);
nor U695 (N_695,In_666,In_1148);
and U696 (N_696,In_1714,In_4462);
or U697 (N_697,In_4120,In_592);
and U698 (N_698,In_3359,In_3782);
nand U699 (N_699,In_4406,In_1609);
nor U700 (N_700,In_2511,N_94);
nand U701 (N_701,In_3871,In_710);
xnor U702 (N_702,In_2456,In_1209);
nand U703 (N_703,In_3019,In_1742);
nand U704 (N_704,In_287,In_4167);
and U705 (N_705,In_516,In_4880);
or U706 (N_706,In_4945,In_525);
and U707 (N_707,In_2557,In_623);
xnor U708 (N_708,In_2274,In_4119);
or U709 (N_709,In_1554,In_202);
and U710 (N_710,In_530,In_1243);
and U711 (N_711,In_2134,In_3229);
xnor U712 (N_712,N_408,In_841);
xnor U713 (N_713,In_1274,In_927);
nand U714 (N_714,In_4662,In_889);
nor U715 (N_715,In_1379,In_3662);
or U716 (N_716,In_3205,In_2893);
nor U717 (N_717,N_228,In_1160);
xnor U718 (N_718,In_354,In_4850);
nor U719 (N_719,In_4504,In_3616);
and U720 (N_720,N_117,In_137);
xor U721 (N_721,In_2281,In_1360);
or U722 (N_722,In_2201,N_380);
xnor U723 (N_723,In_4091,In_640);
or U724 (N_724,N_451,In_604);
nor U725 (N_725,In_3228,In_3006);
xnor U726 (N_726,N_494,In_755);
or U727 (N_727,In_428,In_1298);
nor U728 (N_728,In_3163,In_2984);
and U729 (N_729,In_2897,N_274);
or U730 (N_730,In_1403,In_1827);
xor U731 (N_731,In_1141,In_4007);
nor U732 (N_732,In_163,In_1239);
nand U733 (N_733,In_4301,In_1396);
nand U734 (N_734,In_3034,In_2878);
nand U735 (N_735,In_566,In_1754);
xnor U736 (N_736,In_4631,In_4555);
or U737 (N_737,In_1371,In_1530);
nor U738 (N_738,In_4696,In_1573);
and U739 (N_739,In_311,In_4385);
nor U740 (N_740,In_982,In_2423);
nor U741 (N_741,In_2853,In_1598);
xnor U742 (N_742,In_4377,N_126);
nand U743 (N_743,N_32,N_268);
or U744 (N_744,In_1654,N_160);
or U745 (N_745,In_1085,In_2224);
nand U746 (N_746,In_4378,In_2815);
and U747 (N_747,In_4460,N_225);
nand U748 (N_748,In_3069,In_3383);
or U749 (N_749,In_4764,In_736);
nor U750 (N_750,In_2683,In_822);
or U751 (N_751,N_265,In_2692);
and U752 (N_752,In_1735,In_2119);
xnor U753 (N_753,In_2600,In_1701);
xnor U754 (N_754,In_2006,In_1107);
nor U755 (N_755,In_2424,In_1309);
nand U756 (N_756,In_15,In_1886);
nand U757 (N_757,In_1653,In_1001);
nor U758 (N_758,In_2860,N_550);
xnor U759 (N_759,In_2657,In_2579);
nor U760 (N_760,In_4860,In_3145);
and U761 (N_761,In_150,In_1627);
nand U762 (N_762,In_2691,In_384);
nand U763 (N_763,In_393,N_329);
xor U764 (N_764,In_3437,N_331);
and U765 (N_765,N_699,In_1737);
nor U766 (N_766,In_3992,In_677);
nor U767 (N_767,In_602,N_12);
nor U768 (N_768,In_364,N_479);
xor U769 (N_769,In_237,In_1383);
nand U770 (N_770,In_181,In_1300);
and U771 (N_771,In_2257,In_4927);
nand U772 (N_772,In_2449,In_2096);
xor U773 (N_773,In_809,In_4229);
and U774 (N_774,In_455,In_2925);
or U775 (N_775,In_2002,In_733);
or U776 (N_776,N_90,In_4400);
xor U777 (N_777,In_4413,N_570);
and U778 (N_778,In_568,In_3529);
nand U779 (N_779,In_1937,N_604);
xnor U780 (N_780,N_28,N_102);
xor U781 (N_781,In_2113,In_2490);
nor U782 (N_782,N_611,In_1687);
or U783 (N_783,In_238,In_279);
nand U784 (N_784,In_2124,In_1358);
nand U785 (N_785,In_1112,In_1021);
and U786 (N_786,In_2615,In_2685);
or U787 (N_787,N_586,In_1841);
and U788 (N_788,In_503,In_4024);
and U789 (N_789,In_497,In_3787);
nor U790 (N_790,In_3698,In_4214);
or U791 (N_791,In_3762,In_2759);
nand U792 (N_792,In_4524,N_593);
and U793 (N_793,In_372,In_3556);
nor U794 (N_794,In_1612,In_2660);
nor U795 (N_795,In_2610,In_2433);
or U796 (N_796,In_3182,In_4976);
or U797 (N_797,In_3468,In_843);
nand U798 (N_798,In_4505,In_357);
or U799 (N_799,In_3342,In_902);
nand U800 (N_800,In_2255,In_4521);
nor U801 (N_801,In_944,In_2644);
xor U802 (N_802,In_3358,In_3514);
nand U803 (N_803,In_4402,In_4178);
xor U804 (N_804,In_453,In_3176);
or U805 (N_805,N_233,In_1791);
xnor U806 (N_806,In_3764,In_2667);
nand U807 (N_807,In_595,N_613);
nand U808 (N_808,In_3370,In_1434);
or U809 (N_809,In_881,In_4940);
or U810 (N_810,In_4882,In_2070);
nand U811 (N_811,In_2803,In_4523);
and U812 (N_812,In_4424,N_256);
nand U813 (N_813,In_1334,In_4989);
nor U814 (N_814,In_3985,In_2247);
and U815 (N_815,In_4711,In_4789);
and U816 (N_816,In_127,In_3440);
xor U817 (N_817,In_2755,In_1922);
or U818 (N_818,N_246,In_897);
xor U819 (N_819,N_561,In_1775);
nor U820 (N_820,In_1212,In_292);
and U821 (N_821,In_775,In_541);
xnor U822 (N_822,In_4151,In_531);
or U823 (N_823,In_4253,In_3191);
nand U824 (N_824,In_4607,In_1166);
nor U825 (N_825,N_358,N_259);
or U826 (N_826,In_3583,In_4908);
nand U827 (N_827,In_896,In_3682);
xnor U828 (N_828,N_97,In_3975);
and U829 (N_829,In_3625,In_3291);
xor U830 (N_830,In_85,In_3448);
or U831 (N_831,In_3993,In_2876);
nor U832 (N_832,In_2869,In_1261);
nor U833 (N_833,In_391,In_283);
or U834 (N_834,In_4323,In_2230);
and U835 (N_835,In_1022,N_493);
nand U836 (N_836,In_3209,In_1989);
nand U837 (N_837,In_1150,In_3675);
and U838 (N_838,In_3481,In_1285);
or U839 (N_839,In_2192,In_2574);
nor U840 (N_840,In_4464,In_144);
xnor U841 (N_841,In_3246,In_2602);
nand U842 (N_842,N_167,In_275);
or U843 (N_843,In_189,In_905);
and U844 (N_844,In_2162,In_242);
xor U845 (N_845,In_3497,In_4274);
or U846 (N_846,In_3184,In_1033);
or U847 (N_847,In_1563,In_94);
xor U848 (N_848,In_4590,N_531);
and U849 (N_849,In_2482,In_3869);
nand U850 (N_850,In_3885,N_165);
xnor U851 (N_851,In_4846,In_626);
nor U852 (N_852,In_2054,In_1445);
xnor U853 (N_853,In_898,In_2661);
and U854 (N_854,In_4300,In_4702);
or U855 (N_855,N_412,In_76);
nand U856 (N_856,In_4008,In_1760);
nand U857 (N_857,N_610,N_456);
xor U858 (N_858,In_2594,In_233);
nor U859 (N_859,In_138,In_261);
or U860 (N_860,In_3864,In_3751);
or U861 (N_861,In_2538,In_4245);
xnor U862 (N_862,In_3878,N_114);
nand U863 (N_863,In_996,In_4108);
xnor U864 (N_864,In_3410,In_1562);
and U865 (N_865,In_4218,In_4712);
nor U866 (N_866,N_670,In_422);
xor U867 (N_867,In_2934,In_1944);
xor U868 (N_868,In_2982,In_4790);
nand U869 (N_869,In_2814,N_607);
nand U870 (N_870,In_3179,In_1665);
xnor U871 (N_871,In_4845,N_440);
nand U872 (N_872,In_1265,In_820);
nor U873 (N_873,In_3375,In_4941);
xor U874 (N_874,In_1483,In_2073);
and U875 (N_875,In_3982,In_3344);
or U876 (N_876,In_3854,In_1683);
nand U877 (N_877,In_4686,In_3154);
and U878 (N_878,In_1092,In_3353);
nand U879 (N_879,In_4428,In_2182);
nand U880 (N_880,In_960,In_4313);
nand U881 (N_881,In_199,In_1056);
nand U882 (N_882,In_953,In_1908);
nand U883 (N_883,In_1355,N_248);
or U884 (N_884,In_4951,In_801);
nand U885 (N_885,In_1242,In_2489);
and U886 (N_886,In_1542,N_229);
nor U887 (N_887,In_557,In_4996);
or U888 (N_888,In_4458,In_2560);
nor U889 (N_889,In_3068,N_216);
nand U890 (N_890,In_3947,In_4985);
nand U891 (N_891,In_1858,In_4616);
xnor U892 (N_892,In_925,In_2110);
xnor U893 (N_893,In_3517,In_4065);
nor U894 (N_894,N_338,In_676);
xnor U895 (N_895,In_1015,In_1850);
nand U896 (N_896,In_3106,In_2349);
nor U897 (N_897,In_2834,In_4149);
xor U898 (N_898,In_4319,In_975);
xor U899 (N_899,In_4877,In_1694);
xnor U900 (N_900,In_4902,In_2452);
and U901 (N_901,In_793,N_643);
nor U902 (N_902,In_4295,In_3774);
or U903 (N_903,In_3705,In_474);
and U904 (N_904,In_847,In_4516);
or U905 (N_905,In_1578,N_532);
or U906 (N_906,N_4,In_706);
nand U907 (N_907,In_4679,In_2825);
and U908 (N_908,In_3500,In_2400);
nand U909 (N_909,In_2554,In_1004);
nor U910 (N_910,In_3171,In_838);
and U911 (N_911,In_4539,In_3631);
and U912 (N_912,In_2534,In_3242);
nor U913 (N_913,In_1590,In_2455);
xnor U914 (N_914,N_210,N_501);
and U915 (N_915,N_37,N_552);
or U916 (N_916,In_4077,In_1250);
xnor U917 (N_917,In_3588,In_2798);
nand U918 (N_918,In_1832,In_174);
or U919 (N_919,In_4331,In_1128);
nor U920 (N_920,In_4231,In_3770);
nand U921 (N_921,In_4554,In_4390);
nor U922 (N_922,In_2678,N_146);
nor U923 (N_923,In_1199,In_3896);
xor U924 (N_924,In_4240,In_2010);
or U925 (N_925,In_2746,In_4370);
nor U926 (N_926,In_4838,In_3143);
or U927 (N_927,N_624,In_2165);
nand U928 (N_928,N_199,In_2065);
nand U929 (N_929,In_3492,In_4625);
nor U930 (N_930,In_4926,N_235);
and U931 (N_931,In_3639,In_1613);
and U932 (N_932,N_164,N_332);
nor U933 (N_933,In_968,N_124);
nor U934 (N_934,In_2358,In_825);
nor U935 (N_935,In_2155,In_3345);
nand U936 (N_936,In_220,N_26);
xor U937 (N_937,In_1864,N_569);
nor U938 (N_938,In_1405,In_4427);
xor U939 (N_939,N_500,N_444);
xor U940 (N_940,N_105,In_2472);
nand U941 (N_941,In_4756,In_211);
or U942 (N_942,N_615,N_711);
xnor U943 (N_943,In_4960,In_499);
nand U944 (N_944,In_796,In_1444);
and U945 (N_945,In_4885,In_3642);
xnor U946 (N_946,In_3496,In_1917);
and U947 (N_947,N_441,In_1027);
or U948 (N_948,In_308,In_3067);
xor U949 (N_949,In_2545,In_3386);
nor U950 (N_950,In_3726,In_360);
xor U951 (N_951,In_2405,N_445);
and U952 (N_952,In_4648,In_179);
nor U953 (N_953,In_121,In_2862);
nor U954 (N_954,In_1255,In_3197);
nand U955 (N_955,In_1178,In_2599);
and U956 (N_956,In_937,In_4361);
nand U957 (N_957,In_993,N_682);
xnor U958 (N_958,N_348,In_1188);
nor U959 (N_959,In_1601,In_2578);
nand U960 (N_960,In_4665,N_459);
nand U961 (N_961,N_649,N_400);
and U962 (N_962,In_2107,In_3317);
nor U963 (N_963,In_2645,In_3795);
nand U964 (N_964,N_744,In_4277);
or U965 (N_965,In_1596,N_1);
and U966 (N_966,N_710,N_559);
nand U967 (N_967,In_3630,N_276);
nor U968 (N_968,In_4227,In_4684);
xnor U969 (N_969,In_1699,In_1867);
nor U970 (N_970,In_408,N_43);
or U971 (N_971,In_2040,In_1149);
nor U972 (N_972,In_700,In_3362);
and U973 (N_973,In_162,In_4184);
nor U974 (N_974,In_3657,In_2139);
nor U975 (N_975,In_482,In_2337);
and U976 (N_976,In_3712,N_365);
or U977 (N_977,N_335,In_2577);
and U978 (N_978,In_3235,In_3245);
xor U979 (N_979,In_2996,In_3718);
nor U980 (N_980,In_600,In_3957);
or U981 (N_981,In_4950,N_632);
or U982 (N_982,In_1524,In_4033);
or U983 (N_983,In_2019,In_3980);
and U984 (N_984,In_3391,N_619);
and U985 (N_985,In_2293,In_1322);
nand U986 (N_986,In_4213,N_253);
and U987 (N_987,In_828,In_569);
nor U988 (N_988,N_16,In_4812);
nor U989 (N_989,In_406,In_4366);
nand U990 (N_990,In_3933,N_92);
or U991 (N_991,In_3259,N_275);
nand U992 (N_992,In_3859,In_3052);
nand U993 (N_993,In_3201,N_269);
or U994 (N_994,In_1888,N_511);
xor U995 (N_995,In_1696,N_302);
nor U996 (N_996,In_1427,In_386);
xnor U997 (N_997,In_2069,N_168);
and U998 (N_998,N_407,In_3819);
or U999 (N_999,N_204,N_328);
xor U1000 (N_1000,In_4519,In_1429);
and U1001 (N_1001,In_4881,N_814);
or U1002 (N_1002,N_807,N_708);
or U1003 (N_1003,In_3230,In_1770);
nand U1004 (N_1004,In_3053,In_2883);
nor U1005 (N_1005,N_931,In_1784);
nor U1006 (N_1006,In_3867,N_646);
xnor U1007 (N_1007,N_673,In_1866);
and U1008 (N_1008,N_73,In_3607);
and U1009 (N_1009,N_526,N_224);
xnor U1010 (N_1010,In_4584,N_815);
and U1011 (N_1011,In_2810,In_559);
or U1012 (N_1012,N_529,In_1749);
or U1013 (N_1013,N_366,In_803);
nand U1014 (N_1014,In_3322,N_911);
and U1015 (N_1015,N_702,In_2679);
and U1016 (N_1016,In_3746,In_3294);
or U1017 (N_1017,In_1177,In_3807);
or U1018 (N_1018,N_470,In_3183);
or U1019 (N_1019,In_2131,In_2282);
or U1020 (N_1020,In_1348,In_2312);
and U1021 (N_1021,In_2929,In_3439);
nand U1022 (N_1022,In_4716,In_1757);
nand U1023 (N_1023,In_1589,In_4508);
and U1024 (N_1024,In_1475,In_2354);
and U1025 (N_1025,N_830,N_293);
and U1026 (N_1026,In_2748,In_1655);
and U1027 (N_1027,In_3483,In_1125);
and U1028 (N_1028,In_1647,In_1986);
xor U1029 (N_1029,In_4088,In_4222);
xor U1030 (N_1030,In_1098,In_2913);
nand U1031 (N_1031,N_986,In_3262);
or U1032 (N_1032,In_2589,In_2926);
and U1033 (N_1033,N_997,N_872);
nor U1034 (N_1034,In_2744,In_1216);
xor U1035 (N_1035,In_2627,In_4698);
nor U1036 (N_1036,N_863,In_201);
and U1037 (N_1037,N_647,In_3151);
and U1038 (N_1038,In_2266,In_99);
nand U1039 (N_1039,N_286,N_630);
and U1040 (N_1040,In_3669,N_333);
nand U1041 (N_1041,In_2576,In_1103);
and U1042 (N_1042,In_761,In_3686);
nand U1043 (N_1043,In_1462,In_1798);
xnor U1044 (N_1044,In_3363,In_2361);
nand U1045 (N_1045,In_827,In_1680);
nand U1046 (N_1046,In_941,In_4070);
and U1047 (N_1047,N_696,In_1525);
nand U1048 (N_1048,N_956,In_1121);
and U1049 (N_1049,In_4193,In_1797);
and U1050 (N_1050,In_313,In_903);
nand U1051 (N_1051,In_3579,In_3093);
and U1052 (N_1052,In_3892,In_1982);
nand U1053 (N_1053,In_139,In_3350);
xor U1054 (N_1054,In_288,In_2231);
or U1055 (N_1055,N_299,In_2099);
nand U1056 (N_1056,In_4529,In_546);
nand U1057 (N_1057,In_4244,In_414);
nand U1058 (N_1058,In_3435,In_2839);
or U1059 (N_1059,In_4155,In_1823);
nor U1060 (N_1060,In_854,N_343);
nor U1061 (N_1061,In_2734,In_4794);
nor U1062 (N_1062,In_1292,In_512);
nand U1063 (N_1063,In_2481,N_518);
xor U1064 (N_1064,In_1289,In_3501);
and U1065 (N_1065,In_1124,N_385);
nand U1066 (N_1066,In_596,In_3284);
nor U1067 (N_1067,In_547,In_2285);
xor U1068 (N_1068,In_3575,In_3207);
and U1069 (N_1069,In_2536,In_985);
or U1070 (N_1070,In_3112,In_294);
or U1071 (N_1071,In_2518,In_3586);
and U1072 (N_1072,In_456,In_2350);
nand U1073 (N_1073,In_1246,In_4787);
nand U1074 (N_1074,In_1752,In_3433);
nand U1075 (N_1075,In_299,In_3882);
nand U1076 (N_1076,In_3318,In_4394);
nor U1077 (N_1077,In_3887,In_671);
nor U1078 (N_1078,In_1710,In_4547);
xnor U1079 (N_1079,In_4630,In_1140);
xor U1080 (N_1080,In_4052,In_3115);
xnor U1081 (N_1081,In_3544,In_2731);
or U1082 (N_1082,In_3805,In_3897);
nor U1083 (N_1083,In_3237,In_1933);
and U1084 (N_1084,In_4646,In_1553);
nor U1085 (N_1085,In_2794,In_4426);
and U1086 (N_1086,In_25,In_4311);
nand U1087 (N_1087,In_4470,In_426);
and U1088 (N_1088,In_2227,N_152);
or U1089 (N_1089,N_697,N_853);
and U1090 (N_1090,N_542,In_1192);
xnor U1091 (N_1091,In_68,In_1018);
nor U1092 (N_1092,In_3227,In_239);
or U1093 (N_1093,N_147,In_2555);
nand U1094 (N_1094,In_2769,In_1251);
xor U1095 (N_1095,In_359,N_662);
xnor U1096 (N_1096,N_772,In_490);
nand U1097 (N_1097,In_1635,In_77);
and U1098 (N_1098,N_889,In_2504);
xor U1099 (N_1099,In_1807,In_3269);
nand U1100 (N_1100,N_789,N_919);
xor U1101 (N_1101,In_347,In_1624);
nor U1102 (N_1102,In_2596,In_3716);
and U1103 (N_1103,In_1023,In_147);
nand U1104 (N_1104,N_672,In_3170);
nor U1105 (N_1105,In_1863,In_2609);
or U1106 (N_1106,N_414,In_1764);
nor U1107 (N_1107,In_3178,In_2714);
and U1108 (N_1108,In_1577,In_1602);
or U1109 (N_1109,In_1105,In_1815);
xor U1110 (N_1110,In_1772,In_1706);
or U1111 (N_1111,In_1724,In_1767);
xor U1112 (N_1112,In_1225,In_2939);
nor U1113 (N_1113,In_2558,In_441);
or U1114 (N_1114,In_3283,In_3561);
and U1115 (N_1115,In_83,In_4666);
nand U1116 (N_1116,N_173,N_966);
or U1117 (N_1117,In_2626,N_603);
nor U1118 (N_1118,In_388,N_429);
and U1119 (N_1119,In_291,In_4759);
nor U1120 (N_1120,In_1936,N_503);
xor U1121 (N_1121,In_214,N_627);
nor U1122 (N_1122,In_1446,In_558);
and U1123 (N_1123,In_3063,In_1234);
nor U1124 (N_1124,In_2990,In_4701);
or U1125 (N_1125,In_2985,In_3798);
xor U1126 (N_1126,N_287,N_307);
and U1127 (N_1127,N_731,In_159);
and U1128 (N_1128,In_1871,In_817);
or U1129 (N_1129,In_2032,In_837);
nor U1130 (N_1130,N_169,In_2638);
nor U1131 (N_1131,In_2315,In_3328);
xnor U1132 (N_1132,In_1946,N_884);
and U1133 (N_1133,In_2290,In_4534);
and U1134 (N_1134,N_763,In_332);
or U1135 (N_1135,In_2114,In_1515);
nor U1136 (N_1136,In_2362,N_812);
nor U1137 (N_1137,In_1783,In_216);
nor U1138 (N_1138,In_1854,In_2800);
or U1139 (N_1139,In_1453,In_4477);
nand U1140 (N_1140,In_3539,In_867);
xor U1141 (N_1141,In_2617,N_882);
nand U1142 (N_1142,N_20,In_1063);
or U1143 (N_1143,In_699,In_507);
nand U1144 (N_1144,In_2221,In_686);
xnor U1145 (N_1145,In_2077,N_112);
nand U1146 (N_1146,In_1506,N_83);
xnor U1147 (N_1147,In_3282,In_3161);
nand U1148 (N_1148,In_2684,In_4909);
nor U1149 (N_1149,In_3866,In_2101);
or U1150 (N_1150,In_4068,In_1413);
nor U1151 (N_1151,In_3460,In_4609);
or U1152 (N_1152,In_2112,In_3793);
and U1153 (N_1153,In_1997,In_3073);
or U1154 (N_1154,In_2086,In_2466);
xnor U1155 (N_1155,In_4182,In_427);
or U1156 (N_1156,In_4498,In_4854);
or U1157 (N_1157,N_640,In_2879);
or U1158 (N_1158,N_638,In_1555);
or U1159 (N_1159,In_4784,N_848);
or U1160 (N_1160,In_2765,N_107);
nor U1161 (N_1161,In_2126,In_4112);
nor U1162 (N_1162,In_2933,In_3454);
and U1163 (N_1163,In_3447,In_4761);
or U1164 (N_1164,In_4127,In_729);
xor U1165 (N_1165,In_2946,In_1810);
xor U1166 (N_1166,In_3374,In_4357);
or U1167 (N_1167,In_1081,N_565);
nand U1168 (N_1168,In_3298,In_3901);
or U1169 (N_1169,In_4473,In_277);
or U1170 (N_1170,In_790,In_3075);
nand U1171 (N_1171,N_933,In_1557);
and U1172 (N_1172,N_890,In_2450);
nand U1173 (N_1173,N_992,N_557);
nor U1174 (N_1174,In_2418,In_2569);
and U1175 (N_1175,In_3097,In_3472);
or U1176 (N_1176,In_727,N_826);
nand U1177 (N_1177,In_257,In_1894);
xor U1178 (N_1178,In_1650,In_562);
nand U1179 (N_1179,In_2024,In_4404);
nand U1180 (N_1180,In_2712,In_3395);
xnor U1181 (N_1181,In_2041,In_2461);
or U1182 (N_1182,In_2388,In_4136);
nand U1183 (N_1183,In_118,In_1799);
nor U1184 (N_1184,In_4966,In_3744);
and U1185 (N_1185,In_2917,N_738);
and U1186 (N_1186,In_3489,N_839);
or U1187 (N_1187,In_104,In_4335);
nor U1188 (N_1188,In_1734,In_4851);
and U1189 (N_1189,In_4154,In_1780);
nand U1190 (N_1190,In_2590,In_4567);
and U1191 (N_1191,In_3173,In_3371);
xor U1192 (N_1192,In_928,In_4417);
nor U1193 (N_1193,In_1176,In_2245);
xnor U1194 (N_1194,N_723,N_201);
and U1195 (N_1195,In_4256,In_3308);
nor U1196 (N_1196,In_226,In_1072);
or U1197 (N_1197,In_1288,In_1967);
nor U1198 (N_1198,In_1079,In_1100);
and U1199 (N_1199,In_1336,N_865);
or U1200 (N_1200,In_363,In_495);
nor U1201 (N_1201,In_3070,In_1472);
or U1202 (N_1202,In_2084,In_4165);
xnor U1203 (N_1203,In_3521,In_4492);
or U1204 (N_1204,N_309,In_4281);
nor U1205 (N_1205,In_738,In_3881);
nand U1206 (N_1206,In_4146,In_1169);
xor U1207 (N_1207,In_4278,N_989);
nor U1208 (N_1208,In_1828,In_3038);
xnor U1209 (N_1209,In_3121,N_888);
or U1210 (N_1210,In_2841,In_2762);
or U1211 (N_1211,In_1087,In_3806);
xnor U1212 (N_1212,In_2240,In_2017);
nand U1213 (N_1213,In_3092,In_3003);
or U1214 (N_1214,In_168,In_514);
and U1215 (N_1215,In_818,In_4421);
nor U1216 (N_1216,In_365,In_4258);
or U1217 (N_1217,N_625,In_4642);
or U1218 (N_1218,In_4796,In_1347);
nand U1219 (N_1219,N_56,In_3829);
nor U1220 (N_1220,In_3443,N_965);
and U1221 (N_1221,In_1223,In_1860);
xnor U1222 (N_1222,In_2025,In_1003);
xor U1223 (N_1223,In_2223,In_4884);
and U1224 (N_1224,N_949,In_807);
and U1225 (N_1225,In_4736,In_3699);
nand U1226 (N_1226,N_317,In_1777);
nor U1227 (N_1227,In_2980,In_1790);
nand U1228 (N_1228,In_2053,In_1556);
nor U1229 (N_1229,In_2145,In_976);
nor U1230 (N_1230,In_1174,In_231);
and U1231 (N_1231,In_3840,N_527);
and U1232 (N_1232,N_282,In_654);
nor U1233 (N_1233,In_446,In_509);
nor U1234 (N_1234,N_417,In_4409);
or U1235 (N_1235,N_376,In_1851);
nand U1236 (N_1236,In_2406,N_466);
nor U1237 (N_1237,In_3504,In_3192);
or U1238 (N_1238,N_655,In_1262);
nand U1239 (N_1239,In_2619,In_2135);
or U1240 (N_1240,In_4769,In_1344);
nand U1241 (N_1241,N_609,In_1870);
nor U1242 (N_1242,N_779,In_337);
nor U1243 (N_1243,In_413,In_1817);
nor U1244 (N_1244,In_1688,In_1567);
xor U1245 (N_1245,In_1812,In_1145);
nor U1246 (N_1246,N_616,In_2944);
and U1247 (N_1247,In_1408,In_3001);
xor U1248 (N_1248,In_4710,In_814);
xor U1249 (N_1249,In_3962,In_1855);
nand U1250 (N_1250,In_1385,In_1632);
and U1251 (N_1251,N_930,In_1591);
nor U1252 (N_1252,N_381,N_885);
nor U1253 (N_1253,In_4822,In_3323);
xor U1254 (N_1254,In_2693,In_4645);
or U1255 (N_1255,In_2646,In_2141);
nor U1256 (N_1256,In_3153,In_1719);
nor U1257 (N_1257,In_2384,In_1502);
or U1258 (N_1258,N_935,In_4160);
nor U1259 (N_1259,In_1625,N_410);
nor U1260 (N_1260,N_1090,N_832);
or U1261 (N_1261,In_1409,N_52);
nor U1262 (N_1262,N_845,In_4946);
and U1263 (N_1263,In_3844,In_1582);
and U1264 (N_1264,In_4471,In_2899);
nand U1265 (N_1265,In_1418,N_590);
xor U1266 (N_1266,In_3525,In_4087);
or U1267 (N_1267,N_473,N_659);
xnor U1268 (N_1268,N_247,In_49);
nor U1269 (N_1269,In_2412,In_3917);
nor U1270 (N_1270,N_1189,In_875);
xor U1271 (N_1271,In_4273,In_3079);
nand U1272 (N_1272,N_654,In_3608);
and U1273 (N_1273,In_164,In_3936);
and U1274 (N_1274,In_4949,In_1644);
xor U1275 (N_1275,In_4605,N_1092);
nand U1276 (N_1276,In_1774,In_2278);
or U1277 (N_1277,In_2127,In_460);
nand U1278 (N_1278,In_462,N_1053);
or U1279 (N_1279,In_2275,In_2470);
nor U1280 (N_1280,In_1017,In_336);
and U1281 (N_1281,In_2444,N_1024);
or U1282 (N_1282,In_2681,In_1934);
xnor U1283 (N_1283,In_1703,In_4185);
and U1284 (N_1284,N_575,In_166);
and U1285 (N_1285,N_379,N_533);
nor U1286 (N_1286,In_1519,In_4688);
nand U1287 (N_1287,In_848,In_436);
nor U1288 (N_1288,In_272,In_4078);
nor U1289 (N_1289,N_899,In_2199);
or U1290 (N_1290,N_391,In_1126);
xnor U1291 (N_1291,N_881,In_1930);
nor U1292 (N_1292,In_1845,In_2942);
nor U1293 (N_1293,In_918,In_3948);
nor U1294 (N_1294,In_3953,In_673);
nand U1295 (N_1295,In_2865,In_697);
and U1296 (N_1296,N_996,N_402);
nand U1297 (N_1297,N_206,In_3736);
or U1298 (N_1298,In_1575,N_1026);
nand U1299 (N_1299,In_2299,In_4025);
xor U1300 (N_1300,In_1016,In_3009);
nand U1301 (N_1301,In_3755,In_2036);
nor U1302 (N_1302,In_4179,N_368);
nand U1303 (N_1303,In_424,In_1168);
and U1304 (N_1304,In_3605,In_1238);
nor U1305 (N_1305,In_1954,In_683);
nand U1306 (N_1306,N_382,In_2658);
nor U1307 (N_1307,N_1022,In_3530);
xor U1308 (N_1308,In_1395,In_4191);
nor U1309 (N_1309,N_1108,In_4515);
xnor U1310 (N_1310,In_2089,N_634);
xnor U1311 (N_1311,In_3186,In_298);
nor U1312 (N_1312,N_687,In_3165);
or U1313 (N_1313,N_485,In_4751);
nor U1314 (N_1314,In_1991,In_4638);
nor U1315 (N_1315,In_655,N_175);
and U1316 (N_1316,In_209,N_1089);
nand U1317 (N_1317,In_4375,In_2253);
and U1318 (N_1318,In_1332,In_2629);
or U1319 (N_1319,In_4589,In_1469);
or U1320 (N_1320,In_4852,In_4391);
and U1321 (N_1321,In_4621,In_4655);
nand U1322 (N_1322,In_2330,In_3566);
xor U1323 (N_1323,In_3875,In_4674);
or U1324 (N_1324,In_1599,N_244);
or U1325 (N_1325,N_1183,In_2831);
nor U1326 (N_1326,N_1086,In_934);
nor U1327 (N_1327,N_879,In_821);
nor U1328 (N_1328,N_936,In_1307);
xnor U1329 (N_1329,In_1131,In_646);
and U1330 (N_1330,In_2892,N_877);
xnor U1331 (N_1331,In_458,In_2742);
nand U1332 (N_1332,N_128,In_949);
and U1333 (N_1333,In_465,In_2382);
and U1334 (N_1334,In_866,In_1115);
nor U1335 (N_1335,In_3327,In_1437);
and U1336 (N_1336,In_2365,In_4912);
nand U1337 (N_1337,N_156,In_4432);
or U1338 (N_1338,In_3827,In_3099);
nor U1339 (N_1339,In_464,In_2370);
xnor U1340 (N_1340,N_1203,In_2885);
nand U1341 (N_1341,N_353,In_2052);
nor U1342 (N_1342,In_4971,In_1069);
xnor U1343 (N_1343,N_176,In_3403);
nor U1344 (N_1344,N_346,In_656);
or U1345 (N_1345,In_1630,In_1067);
nand U1346 (N_1346,In_2023,In_2438);
nand U1347 (N_1347,N_115,N_1017);
nand U1348 (N_1348,In_3007,In_1583);
and U1349 (N_1349,In_3015,N_898);
and U1350 (N_1350,N_1101,In_2804);
xnor U1351 (N_1351,In_2050,In_3071);
nor U1352 (N_1352,In_4597,In_1837);
nand U1353 (N_1353,In_3051,In_1824);
nand U1354 (N_1354,In_177,N_480);
and U1355 (N_1355,In_2108,In_4791);
xor U1356 (N_1356,N_1003,In_1895);
xor U1357 (N_1357,In_468,In_1183);
or U1358 (N_1358,In_4259,N_1113);
nand U1359 (N_1359,In_587,In_1450);
and U1360 (N_1360,In_3258,In_860);
nor U1361 (N_1361,In_1766,In_4581);
and U1362 (N_1362,In_2642,In_3367);
or U1363 (N_1363,In_112,In_3650);
nand U1364 (N_1364,In_4202,N_817);
and U1365 (N_1365,N_10,In_2088);
nor U1366 (N_1366,N_734,N_313);
or U1367 (N_1367,In_2251,In_1354);
or U1368 (N_1368,In_224,In_3821);
xor U1369 (N_1369,In_1892,In_1678);
and U1370 (N_1370,N_502,In_856);
or U1371 (N_1371,In_4888,N_489);
nor U1372 (N_1372,N_1004,N_290);
nor U1373 (N_1373,In_725,In_3077);
nor U1374 (N_1374,In_2799,In_2727);
or U1375 (N_1375,N_1041,In_528);
xor U1376 (N_1376,N_521,In_4034);
xor U1377 (N_1377,In_529,N_515);
and U1378 (N_1378,In_2375,In_3655);
or U1379 (N_1379,N_846,N_8);
xnor U1380 (N_1380,In_140,In_2181);
nor U1381 (N_1381,In_2747,N_974);
or U1382 (N_1382,In_2078,In_1659);
nor U1383 (N_1383,In_3621,In_2508);
xnor U1384 (N_1384,In_1294,In_2051);
and U1385 (N_1385,In_4144,In_2859);
nand U1386 (N_1386,In_661,In_4587);
xor U1387 (N_1387,N_909,In_4901);
nor U1388 (N_1388,In_2003,In_614);
or U1389 (N_1389,In_3045,In_335);
and U1390 (N_1390,In_3584,In_4354);
nand U1391 (N_1391,In_3174,N_39);
xnor U1392 (N_1392,N_728,In_3540);
nand U1393 (N_1393,N_741,N_304);
and U1394 (N_1394,In_4064,N_1170);
nand U1395 (N_1395,In_4163,In_3767);
nand U1396 (N_1396,In_2137,In_2376);
nand U1397 (N_1397,In_1324,In_2605);
or U1398 (N_1398,In_3916,In_2454);
and U1399 (N_1399,In_3020,In_3981);
nor U1400 (N_1400,In_50,N_938);
nand U1401 (N_1401,In_3531,N_600);
nor U1402 (N_1402,In_4848,N_597);
nor U1403 (N_1403,In_2269,In_2148);
or U1404 (N_1404,In_3,In_157);
and U1405 (N_1405,In_222,In_1597);
nand U1406 (N_1406,N_34,In_1945);
xnor U1407 (N_1407,In_4564,In_3473);
nand U1408 (N_1408,In_1147,In_2999);
nor U1409 (N_1409,In_1522,In_4487);
xor U1410 (N_1410,In_1722,N_1216);
nor U1411 (N_1411,In_4895,In_3488);
nand U1412 (N_1412,In_4368,In_2625);
xor U1413 (N_1413,In_2027,N_261);
xor U1414 (N_1414,N_514,In_584);
and U1415 (N_1415,In_404,In_3387);
or U1416 (N_1416,In_1048,N_608);
or U1417 (N_1417,N_298,In_2191);
or U1418 (N_1418,N_512,In_3562);
nand U1419 (N_1419,In_1552,In_1909);
nand U1420 (N_1420,In_4315,N_1033);
and U1421 (N_1421,In_2882,In_2935);
and U1422 (N_1422,In_416,In_2280);
nand U1423 (N_1423,In_2022,N_1227);
xor U1424 (N_1424,In_4740,N_1045);
or U1425 (N_1425,In_3032,N_291);
nor U1426 (N_1426,In_1787,In_668);
xor U1427 (N_1427,N_722,In_1839);
nand U1428 (N_1428,In_3120,In_4198);
and U1429 (N_1429,N_831,In_215);
xor U1430 (N_1430,In_3742,N_926);
xor U1431 (N_1431,In_888,N_678);
and U1432 (N_1432,In_879,In_2565);
nor U1433 (N_1433,In_3855,N_426);
nor U1434 (N_1434,In_4388,In_2129);
nand U1435 (N_1435,In_2875,N_1103);
and U1436 (N_1436,N_1238,N_1208);
xnor U1437 (N_1437,N_492,In_21);
and U1438 (N_1438,In_778,In_913);
nand U1439 (N_1439,In_3095,In_339);
nand U1440 (N_1440,N_1185,In_2918);
or U1441 (N_1441,In_2047,In_1451);
or U1442 (N_1442,N_751,In_2033);
nand U1443 (N_1443,In_885,In_865);
or U1444 (N_1444,In_195,In_2167);
nor U1445 (N_1445,In_2122,In_1088);
nand U1446 (N_1446,In_92,In_1266);
nor U1447 (N_1447,N_109,In_950);
and U1448 (N_1448,In_1987,N_88);
or U1449 (N_1449,In_4090,N_21);
xnor U1450 (N_1450,In_2948,In_3203);
and U1451 (N_1451,N_306,In_114);
or U1452 (N_1452,In_4578,N_963);
xor U1453 (N_1453,In_4084,In_1514);
xnor U1454 (N_1454,In_1584,In_634);
xor U1455 (N_1455,N_297,In_3846);
xor U1456 (N_1456,In_2097,In_1264);
xor U1457 (N_1457,In_4775,In_4871);
xnor U1458 (N_1458,In_2316,In_791);
nand U1459 (N_1459,In_2393,In_826);
nor U1460 (N_1460,In_2046,In_1392);
or U1461 (N_1461,In_2653,In_882);
xor U1462 (N_1462,N_241,N_1119);
xnor U1463 (N_1463,In_2854,In_1576);
or U1464 (N_1464,N_1124,In_2235);
and U1465 (N_1465,N_262,In_2435);
nor U1466 (N_1466,N_100,N_797);
nor U1467 (N_1467,N_555,N_991);
nand U1468 (N_1468,In_4660,In_1380);
or U1469 (N_1469,In_3801,In_920);
nor U1470 (N_1470,In_3518,N_378);
xnor U1471 (N_1471,In_1226,N_449);
xnor U1472 (N_1472,In_526,N_143);
nand U1473 (N_1473,In_2133,In_1932);
or U1474 (N_1474,In_96,In_1707);
nor U1475 (N_1475,In_3315,In_3332);
xor U1476 (N_1476,N_405,N_1182);
and U1477 (N_1477,N_23,In_4235);
nor U1478 (N_1478,N_671,In_3299);
nor U1479 (N_1479,In_39,In_549);
and U1480 (N_1480,In_572,In_3600);
and U1481 (N_1481,In_2515,In_1228);
xnor U1482 (N_1482,N_93,In_3850);
nand U1483 (N_1483,N_1093,In_2710);
xor U1484 (N_1484,In_2960,N_436);
nor U1485 (N_1485,N_1145,In_3990);
and U1486 (N_1486,In_4478,In_4699);
nand U1487 (N_1487,In_3150,N_1180);
and U1488 (N_1488,N_520,N_296);
xnor U1489 (N_1489,N_184,N_462);
xnor U1490 (N_1490,In_1438,In_1942);
nand U1491 (N_1491,In_4571,In_3830);
and U1492 (N_1492,In_1638,In_1407);
nand U1493 (N_1493,In_207,In_1286);
nor U1494 (N_1494,In_3388,In_1283);
nand U1495 (N_1495,In_3022,In_3031);
nor U1496 (N_1496,N_1161,N_985);
nor U1497 (N_1497,N_87,N_468);
and U1498 (N_1498,In_2037,N_483);
or U1499 (N_1499,N_849,In_4360);
and U1500 (N_1500,In_2923,N_1381);
xnor U1501 (N_1501,In_397,In_3841);
nor U1502 (N_1502,In_3538,In_2446);
or U1503 (N_1503,N_1377,In_3924);
nand U1504 (N_1504,In_91,In_4995);
or U1505 (N_1505,In_4501,In_693);
nand U1506 (N_1506,N_1050,N_1269);
and U1507 (N_1507,N_395,In_1448);
nor U1508 (N_1508,In_647,In_764);
nand U1509 (N_1509,In_2889,N_1319);
xor U1510 (N_1510,In_2260,In_1661);
and U1511 (N_1511,In_1218,In_3166);
nor U1512 (N_1512,In_3809,In_172);
xnor U1513 (N_1513,In_2279,N_1470);
and U1514 (N_1514,In_4897,In_3743);
xor U1515 (N_1515,N_141,In_3697);
or U1516 (N_1516,N_48,In_4221);
xor U1517 (N_1517,In_2972,N_360);
nor U1518 (N_1518,In_4169,In_2864);
nor U1519 (N_1519,In_3181,N_1066);
and U1520 (N_1520,In_4905,In_2855);
or U1521 (N_1521,In_55,N_1347);
and U1522 (N_1522,In_1743,N_541);
and U1523 (N_1523,In_1623,In_3663);
nand U1524 (N_1524,In_4899,N_821);
xor U1525 (N_1525,In_2805,N_1097);
nor U1526 (N_1526,In_2991,N_85);
or U1527 (N_1527,In_4452,In_2584);
xor U1528 (N_1528,In_2976,In_3914);
nor U1529 (N_1529,N_1361,In_2200);
xor U1530 (N_1530,In_3659,In_4497);
nand U1531 (N_1531,In_1201,N_962);
and U1532 (N_1532,In_1194,In_3804);
or U1533 (N_1533,In_1884,In_466);
nand U1534 (N_1534,N_1249,In_1904);
and U1535 (N_1535,In_4016,In_1814);
xor U1536 (N_1536,In_3880,N_925);
xor U1537 (N_1537,N_1154,In_844);
xnor U1538 (N_1538,N_1312,In_1481);
xor U1539 (N_1539,In_240,In_4197);
nor U1540 (N_1540,In_1889,In_3758);
xnor U1541 (N_1541,In_2011,In_1732);
nand U1542 (N_1542,In_3998,In_2795);
or U1543 (N_1543,In_4833,N_1221);
or U1544 (N_1544,In_915,In_7);
and U1545 (N_1545,In_329,N_955);
xnor U1546 (N_1546,In_3835,N_791);
xor U1547 (N_1547,In_4023,In_2779);
and U1548 (N_1548,N_1369,In_3100);
xnor U1549 (N_1549,In_44,In_1139);
nor U1550 (N_1550,In_4939,N_767);
xor U1551 (N_1551,In_1089,In_1491);
xor U1552 (N_1552,In_493,In_780);
or U1553 (N_1553,N_864,In_4987);
xnor U1554 (N_1554,In_1838,In_3848);
or U1555 (N_1555,N_782,N_1272);
nor U1556 (N_1556,N_1146,N_1257);
nand U1557 (N_1557,N_495,In_4725);
nand U1558 (N_1558,In_4176,In_2377);
nor U1559 (N_1559,In_1693,In_3560);
xnor U1560 (N_1560,In_245,In_1094);
or U1561 (N_1561,N_482,N_957);
and U1562 (N_1562,N_319,In_1359);
xor U1563 (N_1563,In_4372,N_825);
nand U1564 (N_1564,In_4910,In_3157);
or U1565 (N_1565,In_931,In_726);
nand U1566 (N_1566,N_1348,In_4309);
or U1567 (N_1567,In_3466,In_342);
nand U1568 (N_1568,In_2492,In_2613);
nand U1569 (N_1569,In_4932,N_1062);
nor U1570 (N_1570,N_1168,N_422);
and U1571 (N_1571,In_3541,N_1229);
nand U1572 (N_1572,In_4002,In_2507);
and U1573 (N_1573,N_823,In_1480);
xnor U1574 (N_1574,N_857,In_3406);
and U1575 (N_1575,N_1177,In_59);
nand U1576 (N_1576,In_1257,In_1891);
xnor U1577 (N_1577,In_3904,N_403);
or U1578 (N_1578,N_1489,N_1068);
or U1579 (N_1579,N_1451,N_78);
and U1580 (N_1580,In_4959,In_929);
or U1581 (N_1581,N_701,In_2259);
or U1582 (N_1582,N_556,In_4141);
nand U1583 (N_1583,N_704,In_1992);
nand U1584 (N_1584,N_1149,In_1947);
nand U1585 (N_1585,N_35,In_3444);
or U1586 (N_1586,In_3954,In_330);
or U1587 (N_1587,In_4371,N_999);
or U1588 (N_1588,In_3325,N_111);
nor U1589 (N_1589,In_579,In_3421);
nand U1590 (N_1590,In_3756,N_1309);
nand U1591 (N_1591,In_2222,In_1674);
or U1592 (N_1592,In_2649,In_204);
nor U1593 (N_1593,In_2978,N_425);
nor U1594 (N_1594,N_171,In_981);
nor U1595 (N_1595,In_1281,N_471);
nand U1596 (N_1596,N_1118,In_2852);
nor U1597 (N_1597,In_3532,In_307);
nand U1598 (N_1598,In_3057,N_804);
and U1599 (N_1599,In_3267,N_399);
nand U1600 (N_1600,In_669,In_2295);
and U1601 (N_1601,In_4486,N_513);
xor U1602 (N_1602,In_4328,In_4347);
and U1603 (N_1603,In_2729,In_3014);
and U1604 (N_1604,N_1139,N_336);
and U1605 (N_1605,In_2286,In_1580);
or U1606 (N_1606,In_2421,In_1312);
or U1607 (N_1607,N_932,In_812);
nand U1608 (N_1608,In_4887,In_1061);
nor U1609 (N_1609,In_1426,N_467);
or U1610 (N_1610,In_2469,N_1080);
nor U1611 (N_1611,In_3373,In_4704);
or U1612 (N_1612,N_1438,N_594);
or U1613 (N_1613,In_1049,In_2049);
or U1614 (N_1614,In_107,In_3926);
xnor U1615 (N_1615,In_2846,N_1262);
or U1616 (N_1616,N_657,In_1002);
nand U1617 (N_1617,N_1079,In_1083);
nand U1618 (N_1618,In_3402,N_851);
nand U1619 (N_1619,In_78,N_1459);
nand U1620 (N_1620,In_3508,N_910);
nor U1621 (N_1621,In_4220,In_1949);
and U1622 (N_1622,In_3790,In_2339);
nor U1623 (N_1623,N_49,In_517);
nor U1624 (N_1624,In_3172,N_1426);
xor U1625 (N_1625,In_3694,In_241);
and U1626 (N_1626,In_473,In_3799);
xor U1627 (N_1627,In_194,In_1415);
or U1628 (N_1628,In_3791,N_762);
nor U1629 (N_1629,N_507,In_3423);
nor U1630 (N_1630,N_1351,N_1314);
and U1631 (N_1631,N_1473,In_734);
and U1632 (N_1632,In_632,In_2849);
or U1633 (N_1633,In_687,In_265);
or U1634 (N_1634,In_3377,In_1670);
xor U1635 (N_1635,N_367,In_1848);
nor U1636 (N_1636,In_2236,N_805);
and U1637 (N_1637,N_1005,In_4429);
nand U1638 (N_1638,N_981,N_1165);
and U1639 (N_1639,In_434,In_2210);
and U1640 (N_1640,In_2549,In_232);
nor U1641 (N_1641,In_2721,In_109);
and U1642 (N_1642,In_381,In_3078);
nand U1643 (N_1643,In_4447,N_809);
or U1644 (N_1644,In_1826,N_1477);
nor U1645 (N_1645,In_4305,In_2872);
nand U1646 (N_1646,In_1500,N_89);
or U1647 (N_1647,In_805,In_635);
or U1648 (N_1648,N_1284,N_46);
nor U1649 (N_1649,In_599,In_2813);
or U1650 (N_1650,In_1682,N_251);
and U1651 (N_1651,N_937,N_423);
nand U1652 (N_1652,In_3960,N_1099);
nand U1653 (N_1653,N_144,In_2272);
nand U1654 (N_1654,N_185,N_139);
and U1655 (N_1655,In_2004,In_3149);
xnor U1656 (N_1656,In_2886,N_1156);
nor U1657 (N_1657,N_148,N_990);
xor U1658 (N_1658,In_4628,In_961);
or U1659 (N_1659,N_567,In_4856);
and U1660 (N_1660,In_3941,N_1299);
xnor U1661 (N_1661,In_333,In_3336);
or U1662 (N_1662,N_342,In_622);
xnor U1663 (N_1663,In_574,In_3550);
or U1664 (N_1664,N_904,In_3382);
nor U1665 (N_1665,In_1778,In_2542);
xnor U1666 (N_1666,In_1532,In_4709);
nand U1667 (N_1667,N_1070,In_27);
or U1668 (N_1668,N_509,In_3594);
and U1669 (N_1669,In_2807,N_411);
or U1670 (N_1670,In_2146,In_2520);
nand U1671 (N_1671,In_2877,N_238);
and U1672 (N_1672,N_749,In_1526);
xor U1673 (N_1673,In_4813,In_3685);
xor U1674 (N_1674,In_4903,In_4735);
and U1675 (N_1675,In_3585,In_3035);
nor U1676 (N_1676,In_4113,In_4636);
or U1677 (N_1677,N_1367,In_2018);
nand U1678 (N_1678,In_1387,In_1430);
nand U1679 (N_1679,N_591,N_1242);
nor U1680 (N_1680,In_2887,In_4011);
xnor U1681 (N_1681,N_560,In_3135);
nand U1682 (N_1682,In_3199,In_54);
and U1683 (N_1683,In_305,In_591);
nand U1684 (N_1684,N_818,In_4312);
xor U1685 (N_1685,In_4045,In_4330);
and U1686 (N_1686,In_523,N_639);
nor U1687 (N_1687,In_1521,In_1803);
and U1688 (N_1688,N_539,In_581);
or U1689 (N_1689,In_1155,N_760);
or U1690 (N_1690,N_484,In_4291);
nand U1691 (N_1691,In_609,In_2095);
nor U1692 (N_1692,N_1131,In_188);
or U1693 (N_1693,In_4063,In_3677);
xnor U1694 (N_1694,In_3723,N_288);
or U1695 (N_1695,In_2172,N_478);
xnor U1696 (N_1696,N_1402,In_3920);
and U1697 (N_1697,In_2348,In_3414);
xnor U1698 (N_1698,In_2962,In_3547);
xnor U1699 (N_1699,In_1301,N_1025);
nand U1700 (N_1700,In_2411,In_4118);
xnor U1701 (N_1701,In_3961,In_2966);
nor U1702 (N_1702,In_3852,In_792);
nor U1703 (N_1703,N_1359,In_1646);
and U1704 (N_1704,N_667,In_2572);
xnor U1705 (N_1705,In_3356,In_4009);
nand U1706 (N_1706,In_4685,In_3653);
nand U1707 (N_1707,N_1179,N_573);
and U1708 (N_1708,In_4837,In_2380);
and U1709 (N_1709,In_4441,N_1027);
nor U1710 (N_1710,N_1460,N_1250);
and U1711 (N_1711,In_3886,In_1747);
xor U1712 (N_1712,In_4913,In_267);
and U1713 (N_1713,N_345,In_4287);
and U1714 (N_1714,In_636,N_642);
and U1715 (N_1715,In_3935,N_775);
and U1716 (N_1716,In_3252,In_1189);
nand U1717 (N_1717,N_592,In_3081);
or U1718 (N_1718,In_2965,In_102);
nor U1719 (N_1719,In_1939,In_4027);
or U1720 (N_1720,In_4344,In_4356);
xor U1721 (N_1721,N_61,In_295);
nor U1722 (N_1722,N_1293,N_688);
nor U1723 (N_1723,In_1897,In_3320);
xor U1724 (N_1724,In_2725,In_895);
or U1725 (N_1725,In_1468,In_2806);
nand U1726 (N_1726,N_1479,In_1727);
nand U1727 (N_1727,In_1258,In_273);
nor U1728 (N_1728,N_695,In_4772);
nor U1729 (N_1729,In_3921,In_2175);
nor U1730 (N_1730,In_675,N_98);
xor U1731 (N_1731,In_682,N_1420);
nor U1732 (N_1732,In_1345,N_747);
or U1733 (N_1733,In_4974,In_2986);
or U1734 (N_1734,In_2428,In_1973);
nand U1735 (N_1735,In_1833,In_3274);
nor U1736 (N_1736,In_2326,In_4670);
xor U1737 (N_1737,N_1445,In_4349);
and U1738 (N_1738,N_1078,In_3146);
xnor U1739 (N_1739,N_1253,In_945);
xnor U1740 (N_1740,In_3549,N_255);
nor U1741 (N_1741,In_2947,N_658);
nor U1742 (N_1742,In_3368,N_870);
xnor U1743 (N_1743,In_1641,N_1065);
nand U1744 (N_1744,In_3329,In_1319);
nor U1745 (N_1745,N_620,N_984);
and U1746 (N_1746,N_1423,N_861);
nor U1747 (N_1747,In_62,In_2005);
and U1748 (N_1748,In_750,In_1263);
nor U1749 (N_1749,In_318,N_170);
and U1750 (N_1750,N_1433,N_1497);
and U1751 (N_1751,In_3490,N_1123);
nand U1752 (N_1752,N_1516,In_2517);
or U1753 (N_1753,In_2031,N_1169);
xor U1754 (N_1754,In_571,In_1802);
nor U1755 (N_1755,N_357,N_614);
nor U1756 (N_1756,In_3355,N_783);
nand U1757 (N_1757,N_894,N_205);
nand U1758 (N_1758,N_579,In_576);
and U1759 (N_1759,In_4633,In_715);
xnor U1760 (N_1760,N_1021,In_1955);
nand U1761 (N_1761,N_198,In_1663);
nand U1762 (N_1762,In_3950,In_2761);
or U1763 (N_1763,N_792,In_479);
xnor U1764 (N_1764,N_1375,N_1683);
xnor U1765 (N_1765,In_2364,N_1214);
nand U1766 (N_1766,N_1596,In_948);
and U1767 (N_1767,In_2161,In_3614);
xnor U1768 (N_1768,N_928,In_4152);
nand U1769 (N_1769,N_636,N_1623);
nor U1770 (N_1770,In_1603,In_886);
nand U1771 (N_1771,In_3469,N_356);
and U1772 (N_1772,In_1868,In_3873);
nand U1773 (N_1773,N_880,N_1181);
xnor U1774 (N_1774,N_1582,In_2983);
xor U1775 (N_1775,N_1532,N_1107);
and U1776 (N_1776,In_1499,In_2014);
xnor U1777 (N_1777,N_742,N_1114);
nand U1778 (N_1778,In_4348,N_1023);
nor U1779 (N_1779,N_1109,N_716);
nand U1780 (N_1780,In_1926,In_1256);
nand U1781 (N_1781,N_1416,In_1907);
or U1782 (N_1782,N_972,In_3760);
nand U1783 (N_1783,In_4875,N_700);
or U1784 (N_1784,N_1663,In_1110);
xor U1785 (N_1785,In_3107,N_1577);
and U1786 (N_1786,N_1117,N_327);
nor U1787 (N_1787,N_840,N_866);
xnor U1788 (N_1788,N_1018,In_4641);
or U1789 (N_1789,N_301,In_2957);
or U1790 (N_1790,In_711,In_243);
nand U1791 (N_1791,In_2374,In_4652);
nor U1792 (N_1792,In_3064,N_1611);
nor U1793 (N_1793,In_2884,In_3888);
nand U1794 (N_1794,In_1007,In_1750);
and U1795 (N_1795,In_4705,N_1212);
and U1796 (N_1796,In_4333,In_4997);
and U1797 (N_1797,In_1421,In_2528);
and U1798 (N_1798,N_38,In_2173);
nor U1799 (N_1799,N_1624,N_606);
or U1800 (N_1800,In_781,In_3457);
nand U1801 (N_1801,In_1057,N_1741);
nand U1802 (N_1802,N_1435,In_555);
nor U1803 (N_1803,N_1469,N_1200);
and U1804 (N_1804,N_1239,In_1386);
nand U1805 (N_1805,In_786,N_1648);
nand U1806 (N_1806,In_853,In_3691);
and U1807 (N_1807,In_321,In_3599);
nand U1808 (N_1808,In_2636,In_1626);
nand U1809 (N_1809,In_681,In_4263);
or U1810 (N_1810,In_3264,In_3335);
or U1811 (N_1811,In_371,N_730);
nor U1812 (N_1812,In_398,In_2995);
nor U1813 (N_1813,In_1751,N_1604);
nor U1814 (N_1814,In_3890,In_1708);
nand U1815 (N_1815,N_464,N_1569);
or U1816 (N_1816,In_1643,In_3054);
or U1817 (N_1817,In_783,In_3609);
or U1818 (N_1818,N_1412,N_794);
or U1819 (N_1819,N_234,N_254);
or U1820 (N_1820,In_1373,In_2197);
and U1821 (N_1821,In_2300,N_1608);
or U1822 (N_1822,N_1366,In_2256);
nor U1823 (N_1823,In_1310,In_4520);
xor U1824 (N_1824,In_1205,In_1755);
or U1825 (N_1825,In_3326,In_2383);
nor U1826 (N_1826,In_4632,N_370);
nand U1827 (N_1827,In_3721,In_585);
nand U1828 (N_1828,In_4322,In_4173);
or U1829 (N_1829,In_1938,N_803);
nand U1830 (N_1830,In_1458,In_1494);
nor U1831 (N_1831,In_695,N_1235);
nand U1832 (N_1832,In_4099,In_3676);
xor U1833 (N_1833,In_3565,In_4717);
or U1834 (N_1834,In_4952,In_1151);
nor U1835 (N_1835,In_4969,In_3065);
nor U1836 (N_1836,N_813,In_4164);
xor U1837 (N_1837,N_623,N_1084);
nand U1838 (N_1838,In_2953,In_61);
nand U1839 (N_1839,In_1924,In_1401);
and U1840 (N_1840,N_189,In_1026);
or U1841 (N_1841,In_2614,N_1529);
nor U1842 (N_1842,In_4304,In_3891);
nor U1843 (N_1843,N_941,N_1467);
nand U1844 (N_1844,In_3027,N_1593);
nor U1845 (N_1845,In_1038,N_1283);
and U1846 (N_1846,In_3520,In_1840);
or U1847 (N_1847,In_258,In_2174);
and U1848 (N_1848,In_500,N_1195);
xor U1849 (N_1849,N_1194,N_732);
and U1850 (N_1850,In_4615,In_429);
and U1851 (N_1851,N_854,N_80);
nor U1852 (N_1852,In_4777,N_1658);
xor U1853 (N_1853,N_968,In_4265);
and U1854 (N_1854,N_544,In_4603);
and U1855 (N_1855,N_1105,In_2580);
nor U1856 (N_1856,In_103,In_763);
nand U1857 (N_1857,In_2736,In_4216);
and U1858 (N_1858,N_1141,In_3574);
nor U1859 (N_1859,In_4948,In_4190);
xor U1860 (N_1860,In_3239,In_2563);
or U1861 (N_1861,In_3551,N_1616);
xnor U1862 (N_1862,N_1152,In_4722);
xnor U1863 (N_1863,N_1138,N_921);
nand U1864 (N_1864,In_995,In_3647);
nor U1865 (N_1865,In_2494,N_1507);
and U1866 (N_1866,In_4562,In_2816);
nand U1867 (N_1867,N_197,N_1464);
and U1868 (N_1868,N_1060,In_38);
or U1869 (N_1869,N_602,In_651);
nand U1870 (N_1870,N_1526,In_4339);
and U1871 (N_1871,In_3776,N_1649);
nor U1872 (N_1872,In_1397,In_813);
nand U1873 (N_1873,In_4746,In_3110);
and U1874 (N_1874,In_457,N_190);
or U1875 (N_1875,N_824,N_1273);
nor U1876 (N_1876,N_1681,N_1281);
nor U1877 (N_1877,N_1379,In_129);
and U1878 (N_1878,In_4853,In_4228);
or U1879 (N_1879,In_4057,In_2956);
xnor U1880 (N_1880,N_1539,N_27);
nor U1881 (N_1881,In_2341,In_4289);
xor U1882 (N_1882,N_1219,N_1255);
or U1883 (N_1883,In_1071,N_1698);
xor U1884 (N_1884,In_3649,N_1258);
nor U1885 (N_1885,In_3899,In_2355);
nand U1886 (N_1886,N_362,N_759);
and U1887 (N_1887,In_1162,N_295);
or U1888 (N_1888,In_2483,In_4522);
and U1889 (N_1889,N_1210,N_57);
nand U1890 (N_1890,In_3397,In_4723);
nand U1891 (N_1891,In_3255,N_1357);
and U1892 (N_1892,N_906,In_1232);
nand U1893 (N_1893,N_1728,N_448);
xnor U1894 (N_1894,In_1043,In_1844);
or U1895 (N_1895,N_1230,In_310);
nor U1896 (N_1896,In_2468,In_2212);
nand U1897 (N_1897,In_3559,In_2949);
or U1898 (N_1898,In_132,N_1191);
xor U1899 (N_1899,In_491,N_1462);
and U1900 (N_1900,N_446,N_252);
xor U1901 (N_1901,N_1259,In_759);
and U1902 (N_1902,In_1096,In_1711);
and U1903 (N_1903,In_4481,In_3503);
or U1904 (N_1904,N_1160,N_1538);
xnor U1905 (N_1905,N_1543,N_977);
or U1906 (N_1906,N_960,In_334);
xor U1907 (N_1907,N_1384,N_1431);
nand U1908 (N_1908,N_1495,In_2413);
nor U1909 (N_1909,N_1365,In_2271);
xnor U1910 (N_1910,In_2408,N_1335);
xnor U1911 (N_1911,In_2104,In_75);
nor U1912 (N_1912,In_4553,In_932);
xnor U1913 (N_1913,N_1344,N_869);
nand U1914 (N_1914,N_1484,In_2493);
or U1915 (N_1915,In_286,In_323);
or U1916 (N_1916,N_1151,In_3144);
and U1917 (N_1917,In_3449,In_3042);
nand U1918 (N_1918,N_585,N_1602);
nor U1919 (N_1919,In_709,In_463);
nand U1920 (N_1920,In_3060,In_3348);
or U1921 (N_1921,N_1638,In_748);
nand U1922 (N_1922,In_4672,N_580);
and U1923 (N_1923,In_2792,In_4236);
nor U1924 (N_1924,In_3485,In_3619);
or U1925 (N_1925,N_442,In_2694);
and U1926 (N_1926,In_3130,In_4992);
and U1927 (N_1927,In_845,In_2521);
and U1928 (N_1928,N_398,In_3372);
and U1929 (N_1929,N_714,N_1627);
and U1930 (N_1930,In_4816,In_34);
and U1931 (N_1931,In_1422,In_1535);
nand U1932 (N_1932,In_2398,In_4576);
and U1933 (N_1933,N_1632,N_598);
nand U1934 (N_1934,In_1531,In_1976);
nand U1935 (N_1935,N_519,N_1397);
or U1936 (N_1936,In_2567,In_1852);
or U1937 (N_1937,In_1672,N_787);
nand U1938 (N_1938,N_1749,In_533);
and U1939 (N_1939,N_1354,N_166);
or U1940 (N_1940,N_1013,In_2391);
xor U1941 (N_1941,In_133,N_188);
or U1942 (N_1942,N_1387,In_1507);
or U1943 (N_1943,N_1447,N_1289);
and U1944 (N_1944,N_551,N_558);
and U1945 (N_1945,In_3919,In_2568);
nor U1946 (N_1946,In_650,In_4970);
nand U1947 (N_1947,In_3680,N_1556);
xor U1948 (N_1948,N_1677,In_87);
nand U1949 (N_1949,N_833,In_1551);
xor U1950 (N_1950,In_4476,N_1047);
nor U1951 (N_1951,N_1558,In_4454);
nand U1952 (N_1952,In_3734,N_915);
xor U1953 (N_1953,In_3223,In_3636);
nand U1954 (N_1954,In_543,In_444);
xnor U1955 (N_1955,N_929,In_2958);
xnor U1956 (N_1956,In_1270,In_197);
nor U1957 (N_1957,In_4131,In_2243);
nand U1958 (N_1958,N_18,In_3244);
xor U1959 (N_1959,N_1535,In_4140);
or U1960 (N_1960,In_1296,In_3098);
and U1961 (N_1961,In_1559,N_901);
nor U1962 (N_1962,In_2840,In_2331);
nor U1963 (N_1963,In_4383,In_720);
nand U1964 (N_1964,In_4242,In_1248);
xnor U1965 (N_1965,In_4469,N_1536);
and U1966 (N_1966,In_3400,N_668);
xor U1967 (N_1967,In_4134,N_318);
xor U1968 (N_1968,In_4658,In_2208);
nor U1969 (N_1969,In_4892,In_3979);
nor U1970 (N_1970,In_3113,In_3160);
nand U1971 (N_1971,In_1862,In_4000);
nand U1972 (N_1972,In_3601,In_3384);
or U1973 (N_1973,In_1788,In_2559);
xnor U1974 (N_1974,N_41,In_4570);
nand U1975 (N_1975,In_1044,In_3984);
xor U1976 (N_1976,In_3114,In_3198);
or U1977 (N_1977,In_1370,N_1465);
nor U1978 (N_1978,In_785,In_1490);
nand U1979 (N_1979,N_1076,N_1503);
nor U1980 (N_1980,In_2811,N_1006);
nor U1981 (N_1981,N_773,N_1591);
nand U1982 (N_1982,In_2103,In_704);
or U1983 (N_1983,In_3928,In_3405);
nand U1984 (N_1984,In_1726,In_315);
nand U1985 (N_1985,In_657,In_1097);
or U1986 (N_1986,In_3814,N_74);
nand U1987 (N_1987,N_914,In_3823);
nand U1988 (N_1988,In_4442,N_118);
and U1989 (N_1989,In_2352,N_836);
or U1990 (N_1990,In_3023,In_1055);
or U1991 (N_1991,In_2686,In_1135);
or U1992 (N_1992,In_1668,N_537);
and U1993 (N_1993,N_1285,In_670);
or U1994 (N_1994,N_1684,In_1842);
and U1995 (N_1995,In_3794,In_1510);
and U1996 (N_1996,N_1323,N_1701);
nor U1997 (N_1997,In_4215,In_501);
nand U1998 (N_1998,In_4923,In_2671);
xor U1999 (N_1999,N_6,N_1243);
nand U2000 (N_2000,In_16,N_1889);
and U2001 (N_2001,In_1728,In_3667);
nand U2002 (N_2002,N_1849,In_2969);
nor U2003 (N_2003,In_4003,In_2785);
or U2004 (N_2004,In_4928,In_297);
and U2005 (N_2005,N_693,In_4600);
and U2006 (N_2006,In_4760,N_1600);
nand U2007 (N_2007,In_1034,N_834);
and U2008 (N_2008,N_1197,In_2297);
and U2009 (N_2009,In_2414,In_4139);
xor U2010 (N_2010,In_1990,N_1476);
nor U2011 (N_2011,In_855,N_1153);
and U2012 (N_2012,In_2937,In_4593);
nor U2013 (N_2013,In_3777,N_1534);
or U2014 (N_2014,In_1035,In_2109);
and U2015 (N_2015,N_788,N_1571);
nand U2016 (N_2016,In_3041,In_564);
xnor U2017 (N_2017,In_3467,In_2541);
or U2018 (N_2018,In_714,N_477);
nand U2019 (N_2019,N_1353,N_746);
or U2020 (N_2020,N_635,N_450);
xnor U2021 (N_2021,In_4678,N_1828);
nand U2022 (N_2022,In_361,N_1994);
xnor U2023 (N_2023,In_3877,In_2242);
nand U2024 (N_2024,N_1818,N_774);
or U2025 (N_2025,N_1926,In_3385);
nor U2026 (N_2026,In_891,In_3337);
nor U2027 (N_2027,In_1208,In_1656);
xnor U2028 (N_2028,N_1860,N_250);
xor U2029 (N_2029,N_1756,In_1054);
and U2030 (N_2030,In_1523,N_1224);
or U2031 (N_2031,In_4491,N_563);
nor U2032 (N_2032,In_1675,N_1403);
and U2033 (N_2033,N_1932,In_3533);
xor U2034 (N_2034,N_116,N_1848);
nand U2035 (N_2035,In_2777,N_737);
nand U2036 (N_2036,N_1896,N_664);
or U2037 (N_2037,In_4097,In_4921);
nand U2038 (N_2038,In_4058,In_2443);
nor U2039 (N_2039,In_527,In_1363);
xnor U2040 (N_2040,In_1658,N_1821);
or U2041 (N_2041,In_4196,In_470);
nor U2042 (N_2042,In_430,In_4973);
xor U2043 (N_2043,In_4043,In_4588);
and U2044 (N_2044,In_3853,In_4592);
nor U2045 (N_2045,N_1899,N_1732);
nand U2046 (N_2046,In_3470,In_4484);
or U2047 (N_2047,In_306,N_1776);
nor U2048 (N_2048,N_1775,N_1167);
xnor U2049 (N_2049,N_736,In_2912);
nand U2050 (N_2050,In_2206,In_2797);
and U2051 (N_2051,In_1271,In_1059);
xor U2052 (N_2052,In_1820,In_1278);
and U2053 (N_2053,In_1768,N_1132);
and U2054 (N_2054,In_3895,N_1693);
and U2055 (N_2055,N_1842,In_3185);
nand U2056 (N_2056,N_648,N_828);
nor U2057 (N_2057,In_603,In_1326);
or U2058 (N_2058,In_2764,In_3306);
or U2059 (N_2059,In_205,N_1643);
xnor U2060 (N_2060,In_146,In_4669);
xnor U2061 (N_2061,N_1345,N_67);
nand U2062 (N_2062,N_1488,In_3127);
nor U2063 (N_2063,N_1949,In_994);
and U2064 (N_2064,In_3535,In_536);
nand U2065 (N_2065,N_1699,N_312);
nand U2066 (N_2066,N_916,In_1741);
nand U2067 (N_2067,In_1887,N_1597);
and U2068 (N_2068,In_4654,N_582);
and U2069 (N_2069,N_200,In_2547);
nand U2070 (N_2070,In_3266,In_850);
nor U2071 (N_2071,N_1868,N_1645);
or U2072 (N_2072,In_4418,In_964);
nand U2073 (N_2073,In_1432,N_1422);
xor U2074 (N_2074,N_36,In_2357);
nand U2075 (N_2075,N_1406,N_867);
and U2076 (N_2076,N_1277,In_3752);
and U2077 (N_2077,In_2652,In_4629);
nand U2078 (N_2078,In_4954,N_958);
nand U2079 (N_2079,In_707,In_3730);
xnor U2080 (N_2080,In_4459,In_2828);
xor U2081 (N_2081,N_819,N_77);
and U2082 (N_2082,In_4249,N_1618);
xor U2083 (N_2083,In_4124,N_618);
and U2084 (N_2084,In_1846,In_537);
nand U2085 (N_2085,In_2607,N_852);
nor U2086 (N_2086,In_394,In_1537);
and U2087 (N_2087,In_1352,In_1443);
or U2088 (N_2088,In_3915,In_4549);
or U2089 (N_2089,N_1839,In_2359);
and U2090 (N_2090,In_1969,In_1879);
nor U2091 (N_2091,N_196,N_1727);
nor U2092 (N_2092,N_1653,In_1323);
and U2093 (N_2093,N_1376,In_1822);
nor U2094 (N_2094,In_72,In_29);
and U2095 (N_2095,In_1041,N_1903);
xnor U2096 (N_2096,In_2587,In_4770);
or U2097 (N_2097,In_3810,In_206);
nand U2098 (N_2098,N_1440,In_4811);
nor U2099 (N_2099,N_1480,N_1444);
xor U2100 (N_2100,N_1218,In_1935);
nor U2101 (N_2101,In_2009,In_4947);
or U2102 (N_2102,N_1978,N_1724);
xnor U2103 (N_2103,In_2998,In_43);
nor U2104 (N_2104,In_1493,N_447);
or U2105 (N_2105,In_721,In_1416);
nor U2106 (N_2106,In_4158,In_2020);
nor U2107 (N_2107,In_3511,In_2043);
xor U2108 (N_2108,In_392,In_4612);
xor U2109 (N_2109,In_2091,In_870);
xor U2110 (N_2110,In_1343,In_907);
or U2111 (N_2111,In_1773,In_2592);
nor U2112 (N_2112,In_4713,In_1698);
xnor U2113 (N_2113,In_95,In_688);
nand U2114 (N_2114,N_1811,In_758);
or U2115 (N_2115,In_1615,In_2061);
xnor U2116 (N_2116,N_1574,N_745);
or U2117 (N_2117,In_2604,N_1914);
and U2118 (N_2118,In_4237,In_4318);
nand U2119 (N_2119,In_940,N_1215);
and U2120 (N_2120,N_1008,In_4687);
nor U2121 (N_2121,N_1955,In_4507);
xor U2122 (N_2122,In_4840,In_4999);
or U2123 (N_2123,In_3571,In_1204);
xor U2124 (N_2124,In_3553,N_1992);
xnor U2125 (N_2125,N_893,N_1551);
or U2126 (N_2126,In_2772,In_4694);
nor U2127 (N_2127,In_4162,In_4367);
or U2128 (N_2128,In_3238,N_488);
or U2129 (N_2129,N_1282,In_2513);
xor U2130 (N_2130,N_681,In_4724);
nand U2131 (N_2131,In_1187,In_3826);
or U2132 (N_2132,In_3661,N_1386);
or U2133 (N_2133,N_1720,N_847);
nor U2134 (N_2134,In_4801,In_2701);
and U2135 (N_2135,N_121,In_852);
and U2136 (N_2136,In_747,In_3002);
nor U2137 (N_2137,In_2687,In_3737);
or U2138 (N_2138,In_3224,N_1454);
or U2139 (N_2139,N_1990,N_1130);
nand U2140 (N_2140,N_776,In_223);
xnor U2141 (N_2141,In_4979,N_1342);
xor U2142 (N_2142,N_1343,In_5);
nand U2143 (N_2143,N_545,In_3279);
or U2144 (N_2144,N_571,In_521);
or U2145 (N_2145,N_802,N_1098);
nand U2146 (N_2146,In_3872,In_2690);
or U2147 (N_2147,N_1733,N_674);
and U2148 (N_2148,N_1544,In_4297);
xnor U2149 (N_2149,In_819,In_2179);
nor U2150 (N_2150,N_1807,In_551);
nand U2151 (N_2151,In_2801,In_3733);
and U2152 (N_2152,N_1722,In_1313);
nor U2153 (N_2153,N_1159,In_4276);
and U2154 (N_2154,N_1121,N_1316);
and U2155 (N_2155,In_2702,N_1875);
and U2156 (N_2156,N_1071,In_760);
nor U2157 (N_2157,In_2672,In_2385);
nor U2158 (N_2158,N_1816,In_835);
and U2159 (N_2159,In_2324,In_4834);
and U2160 (N_2160,N_1287,In_2895);
xnor U2161 (N_2161,N_1840,N_712);
or U2162 (N_2162,N_939,In_1106);
nor U2163 (N_2163,In_4839,In_3548);
xor U2164 (N_2164,In_919,In_1874);
xnor U2165 (N_2165,N_1918,In_1484);
or U2166 (N_2166,In_4825,N_1743);
nand U2167 (N_2167,N_415,N_1819);
nor U2168 (N_2168,In_0,N_1275);
and U2169 (N_2169,N_1125,In_14);
and U2170 (N_2170,In_4778,In_3195);
and U2171 (N_2171,In_3624,N_1579);
nor U2172 (N_2172,In_19,In_3711);
xnor U2173 (N_2173,N_1500,N_1104);
nand U2174 (N_2174,N_1773,In_782);
or U2175 (N_2175,In_3749,N_369);
nor U2176 (N_2176,In_2329,In_2169);
or U2177 (N_2177,In_1875,In_4998);
nand U2178 (N_2178,In_1928,In_312);
or U2179 (N_2179,In_3124,In_4135);
or U2180 (N_2180,In_1206,In_3893);
nor U2181 (N_2181,N_1784,N_1721);
nand U2182 (N_2182,N_1788,In_1570);
xnor U2183 (N_2183,N_1934,In_2866);
nand U2184 (N_2184,N_131,In_3964);
xnor U2185 (N_2185,N_1486,In_954);
and U2186 (N_2186,In_3740,In_3838);
xnor U2187 (N_2187,In_1227,N_1321);
and U2188 (N_2188,N_1318,In_1197);
nor U2189 (N_2189,N_1937,In_2597);
xor U2190 (N_2190,In_1367,In_4054);
or U2191 (N_2191,In_967,In_167);
and U2192 (N_2192,In_4619,N_1046);
and U2193 (N_2193,In_2402,In_1617);
xor U2194 (N_2194,In_1540,N_1171);
nor U2195 (N_2195,In_1273,N_1970);
nand U2196 (N_2196,N_1641,N_64);
and U2197 (N_2197,In_872,In_4359);
nor U2198 (N_2198,N_270,In_2283);
xnor U2199 (N_2199,In_4183,In_3040);
xnor U2200 (N_2200,In_1999,In_1962);
xor U2201 (N_2201,In_2287,In_816);
nor U2202 (N_2202,In_4015,In_746);
xnor U2203 (N_2203,In_2921,N_1950);
or U2204 (N_2204,N_523,N_1510);
nor U2205 (N_2205,N_316,N_1619);
and U2206 (N_2206,N_1810,In_1211);
nor U2207 (N_2207,In_4448,In_2749);
and U2208 (N_2208,N_543,N_750);
xnor U2209 (N_2209,In_3973,In_1600);
xor U2210 (N_2210,N_1324,In_4779);
nand U2211 (N_2211,In_515,In_4574);
or U2212 (N_2212,In_2000,N_1331);
nand U2213 (N_2213,In_4039,N_1952);
and U2214 (N_2214,In_4142,In_4859);
xor U2215 (N_2215,N_517,In_4493);
nor U2216 (N_2216,In_1000,In_784);
and U2217 (N_2217,In_3438,N_1010);
and U2218 (N_2218,N_1748,In_3056);
and U2219 (N_2219,In_2836,N_781);
or U2220 (N_2220,N_1237,In_2425);
or U2221 (N_2221,N_707,In_4436);
and U2222 (N_2222,N_1463,In_3555);
nand U2223 (N_2223,In_1927,In_2730);
xor U2224 (N_2224,N_729,In_4074);
xor U2225 (N_2225,In_3974,In_4542);
nor U2226 (N_2226,N_1432,In_3043);
or U2227 (N_2227,In_3703,N_953);
xnor U2228 (N_2228,In_3380,N_1923);
or U2229 (N_2229,In_857,In_3128);
xor U2230 (N_2230,In_972,N_1352);
nand U2231 (N_2231,In_1423,In_1512);
nand U2232 (N_2232,N_1204,In_3471);
xor U2233 (N_2233,In_3256,N_1570);
and U2234 (N_2234,In_1853,N_1682);
or U2235 (N_2235,N_1573,N_1659);
and U2236 (N_2236,In_345,In_3188);
nand U2237 (N_2237,N_1147,N_510);
nor U2238 (N_2238,In_3250,N_1584);
nand U2239 (N_2239,In_4121,In_1066);
nand U2240 (N_2240,N_1246,In_2665);
or U2241 (N_2241,N_522,N_1116);
xor U2242 (N_2242,In_3719,In_800);
nor U2243 (N_2243,N_1630,N_524);
nor U2244 (N_2244,In_4269,In_3341);
and U2245 (N_2245,In_4743,N_496);
or U2246 (N_2246,N_691,N_855);
and U2247 (N_2247,In_4726,N_1651);
or U2248 (N_2248,In_3956,N_3);
xor U2249 (N_2249,N_219,N_566);
and U2250 (N_2250,In_66,N_1981);
nor U2251 (N_2251,N_419,N_1135);
xor U2252 (N_2252,In_2963,In_4863);
nor U2253 (N_2253,In_684,N_1514);
or U2254 (N_2254,N_987,In_2974);
nor U2255 (N_2255,In_2289,In_4659);
and U2256 (N_2256,N_260,N_637);
xnor U2257 (N_2257,In_2431,In_4389);
xnor U2258 (N_2258,N_1398,N_644);
xnor U2259 (N_2259,In_511,In_2550);
or U2260 (N_2260,N_158,In_3493);
or U2261 (N_2261,N_340,N_1867);
xnor U2262 (N_2262,In_628,In_115);
xor U2263 (N_2263,N_1150,N_971);
nand U2264 (N_2264,In_3409,In_2539);
nand U2265 (N_2265,N_1276,In_2296);
and U2266 (N_2266,N_2231,In_2310);
or U2267 (N_2267,N_2144,In_1039);
nor U2268 (N_2268,N_1231,N_1921);
nor U2269 (N_2269,In_3087,N_1301);
nor U2270 (N_2270,In_1014,N_1813);
nor U2271 (N_2271,N_355,In_4862);
or U2272 (N_2272,In_2448,In_1715);
or U2273 (N_2273,N_1954,N_2198);
nand U2274 (N_2274,N_1256,In_765);
nand U2275 (N_2275,In_3598,N_1916);
nor U2276 (N_2276,N_1738,In_2781);
and U2277 (N_2277,In_1621,N_2233);
or U2278 (N_2278,N_2178,N_1155);
or U2279 (N_2279,N_715,In_679);
xor U2280 (N_2280,N_1095,In_616);
xor U2281 (N_2281,N_1408,N_1750);
nor U2282 (N_2282,In_2758,In_340);
or U2283 (N_2283,N_2173,In_3706);
xnor U2284 (N_2284,In_4585,N_96);
nor U2285 (N_2285,N_2069,In_1464);
nand U2286 (N_2286,In_4618,N_1162);
or U2287 (N_2287,N_724,N_1244);
or U2288 (N_2288,In_136,In_2371);
nor U2289 (N_2289,In_2409,N_1134);
and U2290 (N_2290,In_1391,N_137);
nand U2291 (N_2291,In_320,In_2641);
nand U2292 (N_2292,In_2919,In_1800);
xor U2293 (N_2293,In_438,N_434);
nand U2294 (N_2294,In_2506,N_280);
or U2295 (N_2295,N_584,In_4930);
xnor U2296 (N_2296,N_1671,In_2732);
and U2297 (N_2297,N_1016,N_733);
nand U2298 (N_2298,N_1675,In_2809);
nand U2299 (N_2299,N_65,In_419);
or U2300 (N_2300,N_1338,N_1341);
xnor U2301 (N_2301,In_280,In_1571);
xor U2302 (N_2302,In_2432,In_4580);
or U2303 (N_2303,N_1308,N_944);
and U2304 (N_2304,In_538,In_1739);
or U2305 (N_2305,N_917,In_385);
or U2306 (N_2306,In_3818,N_409);
nand U2307 (N_2307,In_366,N_820);
nand U2308 (N_2308,N_612,In_2971);
and U2309 (N_2309,N_145,N_1472);
and U2310 (N_2310,In_4551,In_3018);
or U2311 (N_2311,In_924,N_1085);
xor U2312 (N_2312,N_1707,N_969);
xnor U2313 (N_2313,N_2049,In_689);
xnor U2314 (N_2314,In_3331,N_1292);
xnor U2315 (N_2315,N_311,N_705);
nand U2316 (N_2316,N_645,In_4038);
and U2317 (N_2317,N_1758,N_2038);
and U2318 (N_2318,N_1953,In_3534);
xor U2319 (N_2319,In_86,In_3689);
nor U2320 (N_2320,In_1859,N_475);
nor U2321 (N_2321,In_4664,N_1757);
xnor U2322 (N_2322,In_823,In_2832);
xor U2323 (N_2323,In_4604,N_2183);
and U2324 (N_2324,In_4363,N_1332);
and U2325 (N_2325,In_3217,N_1052);
nand U2326 (N_2326,In_1215,N_1261);
nor U2327 (N_2327,In_4511,In_2306);
and U2328 (N_2328,In_3537,In_1222);
nor U2329 (N_2329,N_2103,N_1074);
xnor U2330 (N_2330,N_650,N_1407);
and U2331 (N_2331,N_2240,In_2305);
xor U2332 (N_2332,N_2107,N_1960);
and U2333 (N_2333,In_4496,In_1120);
nand U2334 (N_2334,In_3477,In_2791);
and U2335 (N_2335,In_824,N_1441);
and U2336 (N_2336,N_2191,In_2060);
nand U2337 (N_2337,N_1673,N_1900);
nand U2338 (N_2338,In_2561,In_2650);
or U2339 (N_2339,In_1284,N_765);
xnor U2340 (N_2340,In_4081,N_683);
and U2341 (N_2341,N_1729,In_974);
or U2342 (N_2342,N_964,In_1869);
or U2343 (N_2343,N_2072,In_1805);
or U2344 (N_2344,N_2155,In_229);
nor U2345 (N_2345,In_4894,N_1672);
or U2346 (N_2346,In_4898,N_271);
xor U2347 (N_2347,In_3832,N_1946);
and U2348 (N_2348,N_1966,N_790);
nand U2349 (N_2349,In_3505,N_564);
xor U2350 (N_2350,In_2115,In_58);
xnor U2351 (N_2351,N_1841,N_2176);
nand U2352 (N_2352,In_3816,In_3643);
nand U2353 (N_2353,N_766,In_3753);
xor U2354 (N_2354,N_1443,In_2728);
xnor U2355 (N_2355,N_1522,In_3845);
nand U2356 (N_2356,N_1461,In_2659);
nor U2357 (N_2357,N_2134,In_3946);
and U2358 (N_2358,In_4022,In_4004);
or U2359 (N_2359,N_1714,In_3590);
nor U2360 (N_2360,In_749,N_690);
nor U2361 (N_2361,In_4284,N_540);
or U2362 (N_2362,N_549,In_1919);
or U2363 (N_2363,In_3664,N_858);
nand U2364 (N_2364,In_2740,N_2168);
or U2365 (N_2365,N_1943,In_1547);
or U2366 (N_2366,N_1687,N_1196);
or U2367 (N_2367,N_384,In_4752);
xnor U2368 (N_2368,In_1361,N_1874);
xnor U2369 (N_2369,N_1315,N_1491);
nand U2370 (N_2370,N_1617,N_2249);
nor U2371 (N_2371,N_2097,N_2236);
nor U2372 (N_2372,N_1557,In_105);
and U2373 (N_2373,In_1077,In_1704);
xnor U2374 (N_2374,N_860,N_1612);
or U2375 (N_2375,In_2720,In_2436);
nand U2376 (N_2376,In_4835,N_433);
xor U2377 (N_2377,N_1999,In_1689);
xor U2378 (N_2378,In_4719,N_2230);
nor U2379 (N_2379,N_1524,N_240);
nand U2380 (N_2380,N_1747,In_3513);
xnor U2381 (N_2381,N_404,In_3187);
nand U2382 (N_2382,In_3683,N_923);
xnor U2383 (N_2383,In_4143,In_212);
and U2384 (N_2384,N_562,N_1260);
and U2385 (N_2385,N_2137,N_2221);
or U2386 (N_2386,In_2774,In_3527);
nand U2387 (N_2387,N_231,N_349);
and U2388 (N_2388,In_219,N_359);
and U2389 (N_2389,In_4506,N_427);
and U2390 (N_2390,N_387,N_430);
nor U2391 (N_2391,In_4914,In_3558);
nor U2392 (N_2392,In_830,In_2874);
nand U2393 (N_2393,N_2058,In_846);
xnor U2394 (N_2394,In_2719,N_2013);
or U2395 (N_2395,N_887,In_4561);
or U2396 (N_2396,In_2881,N_1976);
and U2397 (N_2397,N_1560,N_896);
or U2398 (N_2398,In_260,In_2531);
or U2399 (N_2399,In_2410,N_278);
and U2400 (N_2400,In_2338,N_1786);
and U2401 (N_2401,In_3934,In_2303);
and U2402 (N_2402,In_4031,In_627);
and U2403 (N_2403,In_2979,N_1734);
and U2404 (N_2404,N_795,N_392);
and U2405 (N_2405,N_1888,In_2209);
and U2406 (N_2406,In_4093,N_325);
xor U2407 (N_2407,N_1799,N_2139);
or U2408 (N_2408,N_179,N_2003);
xnor U2409 (N_2409,In_3695,In_1690);
or U2410 (N_2410,In_1620,In_4107);
or U2411 (N_2411,In_64,In_1569);
nor U2412 (N_2412,N_1575,In_4226);
xor U2413 (N_2413,In_4668,N_2123);
xor U2414 (N_2414,N_2006,In_642);
nand U2415 (N_2415,In_2833,N_661);
or U2416 (N_2416,In_1964,N_1793);
and U2417 (N_2417,N_1136,In_1629);
nand U2418 (N_2418,In_4721,N_1686);
or U2419 (N_2419,N_2001,N_1030);
and U2420 (N_2420,In_777,In_753);
nand U2421 (N_2421,In_832,In_3138);
and U2422 (N_2422,In_1606,In_1731);
nand U2423 (N_2423,N_487,In_4030);
nor U2424 (N_2424,N_735,N_263);
xnor U2425 (N_2425,N_19,N_2078);
or U2426 (N_2426,In_1529,N_1853);
nor U2427 (N_2427,N_873,N_499);
or U2428 (N_2428,In_3304,N_2200);
and U2429 (N_2429,In_423,In_605);
nor U2430 (N_2430,In_797,In_125);
xor U2431 (N_2431,N_1304,In_3011);
or U2432 (N_2432,N_1370,N_816);
nand U2433 (N_2433,N_1428,N_1977);
xor U2434 (N_2434,N_1808,In_2676);
nor U2435 (N_2435,N_1642,N_1622);
nand U2436 (N_2436,In_619,In_2495);
xor U2437 (N_2437,In_717,In_1207);
and U2438 (N_2438,N_1355,N_1851);
xnor U2439 (N_2439,N_1267,N_1297);
xor U2440 (N_2440,In_3833,N_2002);
xor U2441 (N_2441,In_45,N_1187);
or U2442 (N_2442,N_1690,In_2156);
and U2443 (N_2443,In_2718,In_101);
or U2444 (N_2444,In_1454,In_4479);
nand U2445 (N_2445,N_322,N_1452);
nand U2446 (N_2446,In_2440,N_1513);
or U2447 (N_2447,N_1905,In_4387);
or U2448 (N_2448,N_1940,In_2462);
nand U2449 (N_2449,N_605,In_1104);
nor U2450 (N_2450,N_1656,N_1552);
and U2451 (N_2451,In_1953,N_1655);
or U2452 (N_2452,N_827,In_1082);
nand U2453 (N_2453,N_2088,N_390);
and U2454 (N_2454,In_2566,N_453);
xnor U2455 (N_2455,In_403,In_4718);
nand U2456 (N_2456,In_3366,In_1471);
nand U2457 (N_2457,N_134,N_1586);
xnor U2458 (N_2458,In_135,N_1087);
nor U2459 (N_2459,In_433,In_1195);
nor U2460 (N_2460,In_1330,In_1009);
nand U2461 (N_2461,N_372,In_1972);
or U2462 (N_2462,In_3597,N_534);
or U2463 (N_2463,N_718,In_4290);
nand U2464 (N_2464,N_1837,N_2067);
nand U2465 (N_2465,N_516,N_1689);
xor U2466 (N_2466,N_1599,N_1588);
xnor U2467 (N_2467,N_709,In_4071);
nor U2468 (N_2468,N_1633,N_871);
and U2469 (N_2469,In_3569,N_31);
nand U2470 (N_2470,N_698,In_1834);
and U2471 (N_2471,In_304,In_203);
nand U2472 (N_2472,In_4942,In_1431);
xnor U2473 (N_2473,N_1996,N_2141);
nor U2474 (N_2474,In_2136,In_4855);
or U2475 (N_2475,In_570,N_1430);
nand U2476 (N_2476,N_799,In_373);
or U2477 (N_2477,In_4453,N_136);
xor U2478 (N_2478,N_1975,In_2475);
and U2479 (N_2479,In_2842,N_1787);
and U2480 (N_2480,N_303,N_1007);
nand U2481 (N_2481,N_1661,In_2403);
nor U2482 (N_2482,In_1478,In_1384);
xor U2483 (N_2483,In_2366,In_17);
nor U2484 (N_2484,In_3773,In_1138);
nand U2485 (N_2485,In_4768,In_2262);
nor U2486 (N_2486,N_2216,In_4443);
xnor U2487 (N_2487,N_1525,N_785);
nor U2488 (N_2488,N_2115,N_2076);
or U2489 (N_2489,N_267,In_3596);
xnor U2490 (N_2490,N_1997,In_904);
nor U2491 (N_2491,In_4622,In_1291);
and U2492 (N_2492,N_1938,In_2214);
and U2493 (N_2493,N_2044,In_4204);
or U2494 (N_2494,In_4528,N_2082);
xor U2495 (N_2495,N_595,In_1123);
nand U2496 (N_2496,N_1973,In_1136);
nor U2497 (N_2497,In_3739,In_4465);
nand U2498 (N_2498,N_1057,In_2087);
xor U2499 (N_2499,N_439,N_2192);
nand U2500 (N_2500,In_4407,In_2945);
nand U2501 (N_2501,N_1863,N_2214);
xnor U2502 (N_2502,In_2835,In_13);
xor U2503 (N_2503,N_1742,In_802);
and U2504 (N_2504,N_2397,N_2037);
nand U2505 (N_2505,N_1271,N_2439);
nor U2506 (N_2506,In_1337,N_1939);
nand U2507 (N_2507,N_1615,In_2205);
nor U2508 (N_2508,In_3296,In_3026);
nand U2509 (N_2509,In_1411,N_281);
nor U2510 (N_2510,In_2477,In_3412);
or U2511 (N_2511,In_1318,N_2167);
xnor U2512 (N_2512,N_1206,In_1335);
xor U2513 (N_2513,N_1631,N_752);
nor U2514 (N_2514,N_150,N_2022);
and U2515 (N_2515,N_2251,In_2106);
nand U2516 (N_2516,N_2000,N_970);
nand U2517 (N_2517,In_3606,In_420);
nor U2518 (N_2518,In_3577,N_755);
xnor U2519 (N_2519,In_664,N_2284);
xnor U2520 (N_2520,In_1700,N_1082);
nand U2521 (N_2521,In_2706,N_1247);
nand U2522 (N_2522,N_1102,In_4161);
xor U2523 (N_2523,In_4532,In_3364);
and U2524 (N_2524,In_268,N_2339);
xor U2525 (N_2525,N_2102,N_1236);
or U2526 (N_2526,In_74,N_1173);
or U2527 (N_2527,N_2043,In_1230);
nor U2528 (N_2528,N_2314,In_131);
and U2529 (N_2529,In_1477,N_1458);
nand U2530 (N_2530,In_1279,N_2160);
and U2531 (N_2531,N_194,N_2394);
xnor U2532 (N_2532,In_3324,N_951);
xnor U2533 (N_2533,N_1945,N_1562);
and U2534 (N_2534,In_2502,In_1287);
nand U2535 (N_2535,In_4177,In_1684);
nand U2536 (N_2536,N_1223,N_829);
and U2537 (N_2537,In_2486,N_2481);
or U2538 (N_2538,In_3036,In_425);
xnor U2539 (N_2539,N_1137,N_1126);
xnor U2540 (N_2540,In_1671,N_239);
xnor U2541 (N_2541,N_1240,N_2170);
or U2542 (N_2542,N_2332,In_2698);
nor U2543 (N_2543,In_4232,In_124);
nand U2544 (N_2544,In_4870,In_2188);
nand U2545 (N_2545,In_4296,N_1856);
or U2546 (N_2546,In_861,In_3646);
nand U2547 (N_2547,In_24,N_1172);
or U2548 (N_2548,In_1459,In_445);
or U2549 (N_2549,In_4624,N_2362);
nor U2550 (N_2550,In_483,N_2360);
nor U2551 (N_2551,N_314,N_2273);
nor U2552 (N_2552,In_542,In_2906);
and U2553 (N_2553,In_4690,N_689);
or U2554 (N_2554,N_2291,N_850);
nand U2555 (N_2555,In_2739,In_1819);
or U2556 (N_2556,N_2154,In_324);
xnor U2557 (N_2557,In_200,In_122);
nor U2558 (N_2558,In_2787,N_2016);
nand U2559 (N_2559,In_1758,In_1721);
and U2560 (N_2560,In_1267,In_3278);
nor U2561 (N_2561,N_1792,N_207);
or U2562 (N_2562,In_1857,N_633);
nor U2563 (N_2563,N_2025,N_976);
and U2564 (N_2564,In_3800,In_4986);
nor U2565 (N_2565,N_1142,In_1748);
or U2566 (N_2566,In_2773,N_2324);
xor U2567 (N_2567,N_1054,N_2212);
nor U2568 (N_2568,N_508,N_1515);
nand U2569 (N_2569,N_2477,In_2707);
nor U2570 (N_2570,N_1901,N_1264);
or U2571 (N_2571,N_62,In_2668);
and U2572 (N_2572,N_2417,In_3725);
or U2573 (N_2573,N_222,In_1985);
or U2574 (N_2574,In_4381,N_1767);
xor U2575 (N_2575,In_1357,N_2425);
xnor U2576 (N_2576,N_1274,N_952);
nor U2577 (N_2577,N_1995,N_924);
or U2578 (N_2578,In_1134,N_1568);
xnor U2579 (N_2579,In_594,In_1303);
nor U2580 (N_2580,N_1127,In_1019);
xor U2581 (N_2581,N_106,N_2101);
xor U2582 (N_2582,N_2205,In_2164);
nor U2583 (N_2583,N_1475,In_4988);
xnor U2584 (N_2584,N_50,N_2453);
and U2585 (N_2585,In_2250,N_2052);
and U2586 (N_2586,N_653,N_1228);
xor U2587 (N_2587,In_1541,In_1068);
nor U2588 (N_2588,N_1417,In_768);
nor U2589 (N_2589,N_1796,N_1198);
xnor U2590 (N_2590,N_1838,N_1968);
or U2591 (N_2591,N_1667,N_72);
nor U2592 (N_2592,N_1061,In_3164);
and U2593 (N_2593,In_1321,N_2014);
or U2594 (N_2594,In_3656,N_1211);
nor U2595 (N_2595,In_2598,In_703);
nand U2596 (N_2596,N_2005,N_1178);
and U2597 (N_2597,N_1382,N_753);
xor U2598 (N_2598,N_2290,N_1668);
or U2599 (N_2599,In_251,N_2261);
or U2600 (N_2600,N_1739,In_3868);
and U2601 (N_2601,N_1471,In_4445);
and U2602 (N_2602,In_3360,In_36);
nor U2603 (N_2603,In_4425,In_1762);
and U2604 (N_2604,N_438,N_1158);
nor U2605 (N_2605,In_4116,N_1528);
or U2606 (N_2606,In_4714,N_1075);
nor U2607 (N_2607,N_1831,N_1270);
nor U2608 (N_2608,N_2246,N_1390);
and U2609 (N_2609,N_1744,N_1908);
nor U2610 (N_2610,N_1302,N_934);
or U2611 (N_2611,In_3394,N_801);
xor U2612 (N_2612,N_2312,In_1806);
xor U2613 (N_2613,In_4513,N_2432);
or U2614 (N_2614,N_1561,In_4676);
and U2615 (N_2615,In_840,In_3487);
and U2616 (N_2616,N_2117,In_2334);
and U2617 (N_2617,N_344,In_2753);
and U2618 (N_2618,N_2021,In_4936);
or U2619 (N_2619,In_1876,In_1765);
nor U2620 (N_2620,N_2320,N_800);
xnor U2621 (N_2621,N_2471,N_1726);
and U2622 (N_2622,N_2456,In_2786);
or U2623 (N_2623,N_2187,N_1106);
nor U2624 (N_2624,N_1864,N_393);
or U2625 (N_2625,N_2070,In_4166);
or U2626 (N_2626,In_228,N_2441);
nand U2627 (N_2627,N_2460,In_3059);
or U2628 (N_2628,In_3704,In_4697);
xnor U2629 (N_2629,In_4280,In_33);
or U2630 (N_2630,N_2436,N_1329);
and U2631 (N_2631,N_2450,N_2248);
and U2632 (N_2632,N_1404,In_4076);
nor U2633 (N_2633,In_1032,In_3611);
and U2634 (N_2634,N_975,In_1393);
nor U2635 (N_2635,In_3044,N_727);
xnor U2636 (N_2636,In_3436,In_2026);
nand U2637 (N_2637,In_1789,N_2229);
nand U2638 (N_2638,In_1746,In_2239);
or U2639 (N_2639,N_686,In_3091);
nand U2640 (N_2640,In_4753,N_1009);
or U2641 (N_2641,N_1855,N_2343);
and U2642 (N_2642,In_4059,N_2392);
nand U2643 (N_2643,N_1326,N_1566);
xnor U2644 (N_2644,In_1975,In_3610);
xor U2645 (N_2645,In_4040,In_1165);
or U2646 (N_2646,N_2018,N_2275);
and U2647 (N_2647,N_326,In_1377);
and U2648 (N_2648,In_917,In_4288);
xnor U2649 (N_2649,N_2416,N_1794);
nand U2650 (N_2650,In_3168,N_1286);
or U2651 (N_2651,N_242,N_1567);
nor U2652 (N_2652,In_4535,N_1911);
xnor U2653 (N_2653,N_2132,In_1133);
and U2654 (N_2654,N_692,In_349);
or U2655 (N_2655,N_2385,In_4266);
nor U2656 (N_2656,In_2345,In_1536);
nand U2657 (N_2657,In_3103,In_1046);
xor U2658 (N_2658,N_1843,In_1099);
and U2659 (N_2659,In_4224,In_4857);
and U2660 (N_2660,In_2570,In_532);
and U2661 (N_2661,N_2061,N_22);
nor U2662 (N_2662,N_2415,N_2389);
or U2663 (N_2663,N_1481,N_1936);
and U2664 (N_2664,N_1778,In_2170);
nor U2665 (N_2665,N_2346,In_4890);
xnor U2666 (N_2666,In_1861,N_135);
xor U2667 (N_2667,N_2219,In_3474);
or U2668 (N_2668,N_2213,In_4732);
or U2669 (N_2669,N_2293,In_1745);
xor U2670 (N_2670,N_1034,N_174);
and U2671 (N_2671,N_2331,In_2076);
and U2672 (N_2672,In_3080,N_1759);
or U2673 (N_2673,In_2399,N_2257);
or U2674 (N_2674,N_1035,N_2452);
and U2675 (N_2675,In_3084,N_2064);
xor U2676 (N_2676,In_4302,In_2042);
xnor U2677 (N_2677,N_2152,N_292);
or U2678 (N_2678,In_2343,N_431);
nor U2679 (N_2679,N_2321,N_621);
xnor U2680 (N_2680,In_270,In_4572);
nand U2681 (N_2681,In_1543,N_2444);
nor U2682 (N_2682,In_4051,N_2099);
or U2683 (N_2683,In_4061,In_2092);
xor U2684 (N_2684,N_2024,N_739);
and U2685 (N_2685,N_2414,N_1000);
nand U2686 (N_2686,In_1378,N_2304);
and U2687 (N_2687,N_352,N_2279);
nor U2688 (N_2688,In_4379,N_2458);
nand U2689 (N_2689,In_4586,N_161);
xor U2690 (N_2690,In_649,N_418);
or U2691 (N_2691,In_3401,N_1325);
xor U2692 (N_2692,In_970,In_4883);
nand U2693 (N_2693,In_2496,In_2851);
nand U2694 (N_2694,N_2440,N_2189);
nor U2695 (N_2695,N_1011,N_868);
xnor U2696 (N_2696,N_1678,In_2044);
nor U2697 (N_2697,N_1494,N_2094);
nor U2698 (N_2698,N_1797,N_726);
or U2699 (N_2699,N_1094,N_2374);
nor U2700 (N_2700,N_1780,In_4060);
and U2701 (N_2701,In_4953,In_4369);
nor U2702 (N_2702,N_1222,In_1241);
and U2703 (N_2703,N_2238,In_4649);
or U2704 (N_2704,In_4824,N_1852);
and U2705 (N_2705,N_2263,N_1592);
nand U2706 (N_2706,N_2140,N_1806);
and U2707 (N_2707,In_1024,N_2398);
or U2708 (N_2708,N_2222,N_1421);
xor U2709 (N_2709,In_4755,In_3906);
and U2710 (N_2710,In_4916,N_2162);
and U2711 (N_2711,N_2433,N_758);
xnor U2712 (N_2712,In_376,In_4891);
nand U2713 (N_2713,In_3420,N_2029);
xor U2714 (N_2714,In_766,N_1662);
nand U2715 (N_2715,N_1188,In_2085);
nand U2716 (N_2716,N_1072,N_995);
nand U2717 (N_2717,In_2637,In_4968);
xnor U2718 (N_2718,In_1720,In_1012);
and U2719 (N_2719,N_2051,N_1280);
or U2720 (N_2720,N_1625,In_2356);
xor U2721 (N_2721,In_1102,N_1327);
nand U2722 (N_2722,N_912,In_1801);
or U2723 (N_2723,In_774,In_4395);
or U2724 (N_2724,N_435,In_4874);
and U2725 (N_2725,In_319,In_2485);
and U2726 (N_2726,In_674,In_2079);
and U2727 (N_2727,In_2723,In_400);
xor U2728 (N_2728,In_1080,N_53);
or U2729 (N_2729,N_1725,In_2588);
xor U2730 (N_2730,N_2473,N_504);
or U2731 (N_2731,N_339,N_1825);
or U2732 (N_2732,In_1153,N_2296);
nor U2733 (N_2733,In_3101,In_2190);
nand U2734 (N_2734,N_2245,N_769);
nand U2735 (N_2735,N_2463,N_1580);
and U2736 (N_2736,N_1626,In_2907);
nand U2737 (N_2737,In_4763,In_4147);
nand U2738 (N_2738,In_4627,In_3811);
and U2739 (N_2739,N_2335,In_1712);
or U2740 (N_2740,In_1971,N_1511);
or U2741 (N_2741,N_1450,In_3309);
or U2742 (N_2742,In_892,N_631);
or U2743 (N_2743,N_1791,N_2438);
nor U2744 (N_2744,N_1716,In_2394);
nand U2745 (N_2745,N_748,N_1254);
nand U2746 (N_2746,N_1578,N_1971);
and U2747 (N_2747,N_2497,N_1740);
xnor U2748 (N_2748,In_3627,In_992);
nor U2749 (N_2749,In_2863,N_856);
nand U2750 (N_2750,N_2175,In_524);
nor U2751 (N_2751,In_4393,In_4922);
nor U2752 (N_2752,In_4978,N_455);
xor U2753 (N_2753,In_117,N_2010);
nand U2754 (N_2754,In_3311,In_1282);
xor U2755 (N_2755,N_1063,In_1010);
nor U2756 (N_2756,N_1029,In_1179);
and U2757 (N_2757,N_1910,In_798);
nand U2758 (N_2758,N_1680,N_2448);
nor U2759 (N_2759,In_4271,N_2621);
nand U2760 (N_2760,In_864,N_1559);
nand U2761 (N_2761,In_82,In_1901);
nand U2762 (N_2762,N_1718,In_4831);
nand U2763 (N_2763,In_439,In_4431);
and U2764 (N_2764,In_437,N_706);
nand U2765 (N_2765,In_901,In_1439);
xnor U2766 (N_2766,N_2359,N_1548);
nand U2767 (N_2767,N_1115,N_1349);
xnor U2768 (N_2768,In_2713,N_859);
xor U2769 (N_2769,N_719,N_536);
xor U2770 (N_2770,N_323,In_3681);
nand U2771 (N_2771,In_4994,N_2352);
nor U2772 (N_2772,N_1268,In_2386);
or U2773 (N_2773,N_237,N_2413);
nor U2774 (N_2774,In_322,In_4915);
nor U2775 (N_2775,In_2012,In_1111);
or U2776 (N_2776,N_1906,In_839);
xor U2777 (N_2777,N_2618,In_2013);
xnor U2778 (N_2778,N_1340,N_2300);
or U2779 (N_2779,In_909,N_1456);
nand U2780 (N_2780,N_1782,In_4352);
xor U2781 (N_2781,N_2106,N_2470);
xor U2782 (N_2782,N_1985,N_2412);
nor U2783 (N_2783,N_553,N_629);
nor U2784 (N_2784,In_4049,In_221);
nand U2785 (N_2785,In_851,N_2104);
nor U2786 (N_2786,N_191,N_1418);
or U2787 (N_2787,N_1328,In_829);
nand U2788 (N_2788,In_362,N_113);
nor U2789 (N_2789,In_2130,N_1307);
nand U2790 (N_2790,N_2247,N_1055);
nand U2791 (N_2791,N_2363,In_3717);
and U2792 (N_2792,In_4180,In_1389);
xnor U2793 (N_2793,N_1766,N_2323);
and U2794 (N_2794,In_539,N_2695);
or U2795 (N_2795,N_2340,N_2329);
nor U2796 (N_2796,In_1157,In_1473);
nor U2797 (N_2797,N_2634,N_2745);
xnor U2798 (N_2798,N_1252,N_954);
nor U2799 (N_2799,In_18,In_4558);
nand U2800 (N_2800,In_4780,N_1745);
nand U2801 (N_2801,In_3028,In_4123);
or U2802 (N_2802,N_1961,In_3781);
and U2803 (N_2803,In_3301,N_42);
and U2804 (N_2804,N_2283,N_2319);
nor U2805 (N_2805,In_1440,In_1662);
or U2806 (N_2806,In_3573,N_2210);
xnor U2807 (N_2807,N_1380,N_2174);
or U2808 (N_2808,In_2258,N_1385);
nor U2809 (N_2809,N_583,N_998);
nor U2810 (N_2810,N_2418,In_341);
or U2811 (N_2811,In_876,N_2505);
nand U2812 (N_2812,N_243,In_2264);
nor U2813 (N_2813,N_1802,In_4446);
or U2814 (N_2814,In_4818,N_2307);
xnor U2815 (N_2815,In_2457,N_2009);
nor U2816 (N_2816,In_2442,In_1981);
and U2817 (N_2817,N_2274,N_1691);
nand U2818 (N_2818,N_2691,N_1564);
and U2819 (N_2819,N_2113,N_2120);
and U2820 (N_2820,In_3389,N_277);
and U2821 (N_2821,In_1093,N_2688);
or U2822 (N_2822,N_2053,In_2048);
and U2823 (N_2823,N_1930,N_2663);
nor U2824 (N_2824,N_2587,N_1695);
nor U2825 (N_2825,N_1541,In_2143);
nor U2826 (N_2826,In_652,N_2333);
nor U2827 (N_2827,N_2703,In_2234);
nand U2828 (N_2828,N_2042,In_2203);
xor U2829 (N_2829,In_2871,In_4189);
xor U2830 (N_2830,N_2179,In_143);
and U2831 (N_2831,In_1369,N_1755);
and U2832 (N_2832,N_2580,In_1476);
xor U2833 (N_2833,In_708,N_663);
xnor U2834 (N_2834,N_1770,N_215);
and U2835 (N_2835,N_2041,N_2721);
nand U2836 (N_2836,In_2016,N_2316);
nor U2837 (N_2837,N_1038,N_2655);
nor U2838 (N_2838,N_2036,N_2555);
nand U2839 (N_2839,N_2334,N_2490);
nand U2840 (N_2840,In_2770,In_1843);
or U2841 (N_2841,N_2435,N_1213);
nor U2842 (N_2842,N_2538,In_1705);
or U2843 (N_2843,N_546,In_1918);
or U2844 (N_2844,In_1830,N_1120);
or U2845 (N_2845,In_971,N_703);
and U2846 (N_2846,N_2357,In_98);
nor U2847 (N_2847,N_2467,N_1834);
and U2848 (N_2848,In_4397,In_4206);
xor U2849 (N_2849,In_37,In_1518);
or U2850 (N_2850,In_3404,N_2511);
and U2851 (N_2851,In_3554,N_129);
nand U2852 (N_2852,N_2309,N_2195);
xnor U2853 (N_2853,In_762,In_2639);
and U2854 (N_2854,N_2543,N_2472);
xnor U2855 (N_2855,In_2654,N_481);
or U2856 (N_2856,In_3591,N_1251);
xor U2857 (N_2857,N_2218,In_4072);
nand U2858 (N_2858,N_588,In_73);
nor U2859 (N_2859,N_1442,In_4814);
or U2860 (N_2860,In_1198,N_2465);
or U2861 (N_2861,In_4461,In_1539);
nor U2862 (N_2862,N_2289,N_2689);
or U2863 (N_2863,In_2928,N_2220);
xor U2864 (N_2864,N_1589,N_2684);
or U2865 (N_2865,In_3512,In_2241);
nand U2866 (N_2866,N_1822,In_3281);
xor U2867 (N_2867,N_2354,In_2724);
nand U2868 (N_2868,In_4868,N_232);
or U2869 (N_2869,N_2298,N_2040);
nor U2870 (N_2870,In_4192,N_2399);
and U2871 (N_2871,In_1441,N_1389);
and U2872 (N_2872,In_2207,N_628);
or U2873 (N_2873,N_2541,N_1696);
and U2874 (N_2874,N_2605,In_2822);
and U2875 (N_2875,In_2880,N_1644);
nand U2876 (N_2876,N_2017,In_1181);
and U2877 (N_2877,In_3674,In_3747);
and U2878 (N_2878,N_2600,N_1241);
xnor U2879 (N_2879,In_120,In_1118);
xor U2880 (N_2880,In_4896,N_2153);
or U2881 (N_2881,N_2674,N_1809);
or U2882 (N_2882,N_913,In_4626);
or U2883 (N_2883,In_4205,N_1988);
xnor U2884 (N_2884,N_1654,In_2008);
nand U2885 (N_2885,N_1883,In_155);
nor U2886 (N_2886,N_2503,In_328);
xor U2887 (N_2887,N_1001,In_723);
or U2888 (N_2888,N_1248,N_1964);
or U2889 (N_2889,In_1988,N_1928);
nor U2890 (N_2890,N_1760,N_2096);
nor U2891 (N_2891,N_835,In_1592);
and U2892 (N_2892,In_3943,N_1640);
xor U2893 (N_2893,In_563,N_2126);
nor U2894 (N_2894,In_1968,In_2128);
xor U2895 (N_2895,N_2258,N_2673);
nor U2896 (N_2896,N_1845,In_4171);
nor U2897 (N_2897,N_1233,N_334);
and U2898 (N_2898,In_4749,N_581);
and U2899 (N_2899,In_1119,N_2715);
or U2900 (N_2900,In_317,In_51);
or U2901 (N_2901,In_4799,In_1402);
nor U2902 (N_2902,In_2977,N_2733);
and U2903 (N_2903,N_2146,In_3692);
nor U2904 (N_2904,N_1958,N_1372);
xnor U2905 (N_2905,N_2656,N_1091);
xor U2906 (N_2906,N_1482,In_4217);
xor U2907 (N_2907,N_2027,N_1313);
or U2908 (N_2908,N_1414,N_2606);
nand U2909 (N_2909,N_883,N_2502);
nand U2910 (N_2910,N_2379,In_1509);
nand U2911 (N_2911,In_2525,In_1618);
xor U2912 (N_2912,N_1779,N_1902);
and U2913 (N_2913,N_1081,In_3910);
xor U2914 (N_2914,N_474,N_1850);
or U2915 (N_2915,In_1040,In_1769);
xor U2916 (N_2916,In_3828,In_1921);
and U2917 (N_2917,N_2227,N_2517);
xor U2918 (N_2918,N_2446,N_1300);
nor U2919 (N_2919,N_2442,N_2642);
nand U2920 (N_2920,N_756,In_235);
xnor U2921 (N_2921,N_2081,In_1631);
and U2922 (N_2922,N_2671,In_770);
xor U2923 (N_2923,N_1993,In_1058);
and U2924 (N_2924,In_1051,N_2482);
and U2925 (N_2925,In_1425,In_3426);
nand U2926 (N_2926,N_2237,N_163);
xor U2927 (N_2927,N_2235,In_2867);
xor U2928 (N_2928,In_2514,N_2008);
nor U2929 (N_2929,N_1873,N_2569);
and U2930 (N_2930,N_2143,N_1028);
xnor U2931 (N_2931,In_4596,N_822);
and U2932 (N_2932,In_331,N_1164);
or U2933 (N_2933,In_1588,N_2464);
or U2934 (N_2934,N_1371,N_2127);
xnor U2935 (N_2935,N_1904,In_2265);
or U2936 (N_2936,In_3354,In_980);
xnor U2937 (N_2937,In_278,In_3289);
xnor U2938 (N_2938,N_652,N_1692);
or U2939 (N_2939,N_2130,In_4450);
xor U2940 (N_2940,In_3381,N_743);
nand U2941 (N_2941,In_2780,N_1112);
or U2942 (N_2942,N_1731,N_2524);
or U2943 (N_2943,In_3509,In_4540);
nand U2944 (N_2944,In_2381,In_4730);
and U2945 (N_2945,N_1509,N_2287);
nor U2946 (N_2946,N_1362,N_2582);
and U2947 (N_2947,In_4575,N_1508);
nand U2948 (N_2948,In_4341,In_2931);
xor U2949 (N_2949,N_2461,In_4422);
or U2950 (N_2950,N_2519,In_1716);
or U2951 (N_2951,N_2635,N_2539);
nand U2952 (N_2952,N_2632,N_1650);
nand U2953 (N_2953,N_811,In_3290);
xor U2954 (N_2954,N_1542,In_1237);
xnor U2955 (N_2955,N_874,N_1193);
nor U2956 (N_2956,N_771,In_4650);
and U2957 (N_2957,N_2730,N_371);
nor U2958 (N_2958,N_1388,N_461);
xnor U2959 (N_2959,N_1572,N_1703);
and U2960 (N_2960,N_2528,In_3491);
nor U2961 (N_2961,In_156,N_1425);
xnor U2962 (N_2962,N_2035,In_518);
and U2963 (N_2963,N_1814,In_4707);
nand U2964 (N_2964,In_343,N_2598);
and U2965 (N_2965,In_3141,In_1574);
nor U2966 (N_2966,In_42,In_2132);
and U2967 (N_2967,N_2551,N_2285);
nand U2968 (N_2968,In_2154,N_1869);
nand U2969 (N_2969,N_1485,N_2411);
nand U2970 (N_2970,N_1320,In_4343);
nor U2971 (N_2971,In_1260,In_4251);
xor U2972 (N_2972,N_2372,In_3083);
and U2973 (N_2973,In_3089,In_3658);
nor U2974 (N_2974,In_1356,In_3263);
and U2975 (N_2975,In_2898,N_1774);
or U2976 (N_2976,In_1070,N_1527);
and U2977 (N_2977,In_2284,N_1880);
nand U2978 (N_2978,N_713,In_1996);
xor U2979 (N_2979,In_938,N_2513);
xor U2980 (N_2980,N_2050,In_4209);
and U2981 (N_2981,N_1336,N_2564);
xor U2982 (N_2982,N_2619,N_452);
nor U2983 (N_2983,N_2142,N_2612);
nand U2984 (N_2984,N_2109,N_2365);
nor U2985 (N_2985,In_3214,N_1768);
nand U2986 (N_2986,In_4962,N_599);
and U2987 (N_2987,In_2993,N_1483);
nor U2988 (N_2988,In_4766,In_4338);
or U2989 (N_2989,N_1424,N_1322);
nor U2990 (N_2990,N_2512,N_2361);
nand U2991 (N_2991,In_4001,N_907);
and U2992 (N_2992,N_2562,N_1358);
nand U2993 (N_2993,In_4208,N_208);
xnor U2994 (N_2994,N_808,In_3431);
xor U2995 (N_2995,N_2434,In_266);
and U2996 (N_2996,N_2400,N_1506);
or U2997 (N_2997,N_721,In_946);
and U2998 (N_2998,N_2370,In_607);
xnor U2999 (N_2999,In_2407,In_4788);
nand U3000 (N_3000,N_1761,N_2522);
xor U3001 (N_3001,In_4145,In_4337);
and U3002 (N_3002,In_4819,N_2457);
or U3003 (N_3003,N_2701,In_4005);
and U3004 (N_3004,N_1405,N_2402);
nand U3005 (N_3005,N_2610,N_2900);
nand U3006 (N_3006,In_3430,N_920);
nand U3007 (N_3007,In_2635,In_2387);
or U3008 (N_3008,N_458,N_2858);
or U3009 (N_3009,In_3563,In_3545);
and U3010 (N_3010,N_680,N_2675);
nand U3011 (N_3011,In_3883,In_2434);
xnor U3012 (N_3012,In_1339,In_2768);
xor U3013 (N_3013,N_2373,N_1220);
nand U3014 (N_3014,N_2387,N_2407);
and U3015 (N_3015,N_2911,N_2629);
and U3016 (N_3016,N_1111,In_2476);
nor U3017 (N_3017,N_947,N_1374);
nand U3018 (N_3018,In_3785,In_638);
or U3019 (N_3019,In_3741,N_1493);
or U3020 (N_3020,N_1554,In_1568);
nand U3021 (N_3021,In_2808,In_1912);
and U3022 (N_3022,N_1012,N_685);
and U3023 (N_3023,N_1803,N_666);
xor U3024 (N_3024,N_2789,N_538);
nand U3025 (N_3025,N_2685,In_4092);
and U3026 (N_3026,N_2970,In_3251);
nor U3027 (N_3027,N_1576,In_1146);
or U3028 (N_3028,In_1702,N_2938);
and U3029 (N_3029,N_1306,N_1972);
nand U3030 (N_3030,In_2524,N_2768);
nor U3031 (N_3031,N_1647,N_1409);
and U3032 (N_3032,N_2090,In_149);
nand U3033 (N_3033,N_2682,N_2079);
nor U3034 (N_3034,N_1546,In_2333);
nor U3035 (N_3035,N_2306,In_2593);
nand U3036 (N_3036,In_2695,N_1639);
or U3037 (N_3037,N_2065,N_1225);
xnor U3038 (N_3038,N_1517,N_2709);
xor U3039 (N_3039,In_3528,In_4019);
nor U3040 (N_3040,N_2084,In_4133);
and U3041 (N_3041,N_1772,N_2846);
xnor U3042 (N_3042,N_2318,N_2763);
xor U3043 (N_3043,N_2832,N_2743);
or U3044 (N_3044,In_4115,N_236);
xor U3045 (N_3045,In_3909,In_2522);
or U3046 (N_3046,N_1798,N_47);
or U3047 (N_3047,N_768,N_2250);
or U3048 (N_3048,N_2705,N_2839);
nand U3049 (N_3049,In_1679,In_2870);
or U3050 (N_3050,N_1723,In_1);
xor U3051 (N_3051,In_2335,In_1622);
and U3052 (N_3052,N_1795,In_2497);
xor U3053 (N_3053,In_4983,In_3398);
nor U3054 (N_3054,N_2196,In_3261);
nand U3055 (N_3055,In_2651,In_874);
nand U3056 (N_3056,N_2592,N_2637);
nand U3057 (N_3057,N_2046,N_2973);
nor U3058 (N_3058,N_2820,N_2825);
xnor U3059 (N_3059,N_2891,N_2683);
nor U3060 (N_3060,In_2083,N_2243);
nand U3061 (N_3061,N_1174,N_2136);
or U3062 (N_3062,In_4919,In_421);
nor U3063 (N_3063,N_886,N_2823);
or U3064 (N_3064,N_2186,N_2342);
xor U3065 (N_3065,N_2811,In_3445);
nor U3066 (N_3066,N_1657,N_2760);
xor U3067 (N_3067,N_2506,N_1753);
and U3068 (N_3068,N_1777,In_4886);
or U3069 (N_3069,N_959,N_2813);
or U3070 (N_3070,In_859,N_2998);
nand U3071 (N_3071,In_2530,N_2294);
or U3072 (N_3072,N_2579,N_862);
nor U3073 (N_3073,N_994,N_1594);
nor U3074 (N_3074,In_296,N_2916);
nor U3075 (N_3075,In_407,In_2677);
and U3076 (N_3076,In_1835,N_720);
nand U3077 (N_3077,N_1549,N_2647);
or U3078 (N_3078,N_2177,N_1935);
and U3079 (N_3079,N_2681,N_2772);
xnor U3080 (N_3080,N_1186,N_486);
xor U3081 (N_3081,In_1302,In_3333);
nand U3082 (N_3082,N_669,N_2914);
xnor U3083 (N_3083,N_2849,In_2551);
or U3084 (N_3084,N_1051,N_2338);
and U3085 (N_3085,N_341,N_2262);
and U3086 (N_3086,N_2739,N_2479);
nand U3087 (N_3087,N_1368,N_2633);
or U3088 (N_3088,N_2896,N_2574);
nand U3089 (N_3089,N_2376,N_1265);
and U3090 (N_3090,N_1715,N_1448);
nor U3091 (N_3091,In_3778,In_1050);
nand U3092 (N_3092,In_1813,N_2943);
and U3093 (N_3093,N_2728,In_2195);
or U3094 (N_3094,N_2716,In_2845);
nor U3095 (N_3095,N_2384,N_1088);
xnor U3096 (N_3096,N_1520,N_2299);
nor U3097 (N_3097,N_2487,N_1765);
xnor U3098 (N_3098,N_946,In_3232);
or U3099 (N_3099,N_1933,N_2019);
or U3100 (N_3100,In_4613,In_2090);
xnor U3101 (N_3101,N_1635,In_611);
and U3102 (N_3102,N_2485,In_4911);
or U3103 (N_3103,In_1028,N_2267);
or U3104 (N_3104,N_1205,N_1717);
and U3105 (N_3105,In_3442,N_2459);
or U3106 (N_3106,N_2894,N_1439);
nor U3107 (N_3107,In_447,In_1277);
nor U3108 (N_3108,N_2847,N_694);
nand U3109 (N_3109,In_3458,N_2946);
and U3110 (N_3110,In_1951,N_2180);
nand U3111 (N_3111,N_1769,In_2527);
nor U3112 (N_3112,In_1127,N_1833);
nand U3113 (N_3113,In_3231,In_588);
xnor U3114 (N_3114,In_3220,N_1735);
xnor U3115 (N_3115,In_633,N_1637);
or U3116 (N_3116,N_2744,N_2165);
or U3117 (N_3117,N_2940,N_2313);
or U3118 (N_3118,N_1609,N_1360);
nor U3119 (N_3119,N_2350,In_225);
or U3120 (N_3120,In_3147,In_2606);
nand U3121 (N_3121,In_2039,In_1893);
xnor U3122 (N_3122,In_1217,N_2962);
nor U3123 (N_3123,In_65,N_1746);
nor U3124 (N_3124,In_52,N_2790);
nand U3125 (N_3125,N_2699,In_756);
xnor U3126 (N_3126,N_1296,N_2884);
and U3127 (N_3127,N_1719,N_1143);
xor U3128 (N_3128,N_2770,In_3856);
and U3129 (N_3129,In_1159,N_1110);
nor U3130 (N_3130,In_3825,N_375);
or U3131 (N_3131,N_1790,In_943);
or U3132 (N_3132,N_2239,In_1941);
nand U3133 (N_3133,N_2758,N_2842);
nand U3134 (N_3134,N_1610,N_1700);
or U3135 (N_3135,N_15,N_1983);
xor U3136 (N_3136,N_2149,N_2020);
and U3137 (N_3137,In_236,In_3923);
and U3138 (N_3138,In_259,In_3061);
or U3139 (N_3139,N_2401,N_127);
xnor U3140 (N_3140,N_979,N_2206);
and U3141 (N_3141,In_234,In_779);
xnor U3142 (N_3142,N_1660,In_1831);
and U3143 (N_3143,N_2383,N_988);
nand U3144 (N_3144,N_2597,N_876);
nand U3145 (N_3145,N_1446,In_184);
and U3146 (N_3146,N_1666,In_2699);
nor U3147 (N_3147,In_1020,In_806);
nor U3148 (N_3148,N_1895,N_1892);
and U3149 (N_3149,N_940,N_2723);
xor U3150 (N_3150,N_2660,In_2144);
nor U3151 (N_3151,In_4103,In_1709);
nand U3152 (N_3152,N_2850,N_2623);
xor U3153 (N_3153,In_2715,N_2188);
nand U3154 (N_3154,In_1184,N_181);
and U3155 (N_3155,N_2992,N_1184);
xor U3156 (N_3156,N_2930,N_2523);
or U3157 (N_3157,In_3062,In_2952);
and U3158 (N_3158,N_2197,In_1882);
or U3159 (N_3159,N_2987,In_4601);
xor U3160 (N_3160,N_1140,In_963);
and U3161 (N_3161,N_2755,N_2520);
xnor U3162 (N_3162,N_2345,In_3702);
or U3163 (N_3163,N_1974,In_3297);
nor U3164 (N_3164,In_2752,N_321);
or U3165 (N_3165,N_1002,N_2777);
xnor U3166 (N_3166,N_2901,In_4634);
nor U3167 (N_3167,N_1278,N_1674);
and U3168 (N_3168,N_2371,N_2700);
and U3169 (N_3169,N_2566,In_2711);
or U3170 (N_3170,N_2159,In_989);
xor U3171 (N_3171,N_2668,In_4544);
xor U3172 (N_3172,In_3665,N_1636);
or U3173 (N_3173,N_91,In_3465);
or U3174 (N_3174,N_2161,In_900);
nand U3175 (N_3175,In_2523,N_386);
nor U3176 (N_3176,In_3813,In_1994);
nor U3177 (N_3177,In_984,N_1907);
xor U3178 (N_3178,N_2971,N_675);
and U3179 (N_3179,N_2874,In_31);
xor U3180 (N_3180,N_2757,In_161);
nor U3181 (N_3181,N_2927,N_1565);
nand U3182 (N_3182,In_368,N_2277);
or U3183 (N_3183,In_1400,In_1013);
nor U3184 (N_3184,N_2575,In_4386);
and U3185 (N_3185,In_2473,N_2870);
xor U3186 (N_3186,In_1253,In_478);
nor U3187 (N_3187,N_2640,N_2381);
nand U3188 (N_3188,In_3632,N_973);
nor U3189 (N_3189,In_4314,N_796);
nor U3190 (N_3190,N_1519,N_2317);
xor U3191 (N_3191,N_17,N_2818);
nand U3192 (N_3192,N_2311,N_2303);
xor U3193 (N_3193,N_119,N_1827);
nor U3194 (N_3194,N_2667,In_2994);
or U3195 (N_3195,In_2291,In_4938);
nand U3196 (N_3196,In_4080,In_4745);
nor U3197 (N_3197,N_943,In_2573);
nor U3198 (N_3198,N_2989,N_132);
nor U3199 (N_3199,In_2847,In_4503);
and U3200 (N_3200,N_2217,N_2604);
or U3201 (N_3201,In_505,In_3679);
nand U3202 (N_3202,N_2581,N_1621);
and U3203 (N_3203,In_1182,In_4610);
xnor U3204 (N_3204,In_1497,N_2419);
and U3205 (N_3205,N_1199,N_1898);
xnor U3206 (N_3206,In_271,N_257);
xnor U3207 (N_3207,N_1058,N_1835);
or U3208 (N_3208,N_2704,N_1897);
or U3209 (N_3209,N_2807,In_4991);
xor U3210 (N_3210,N_300,N_1944);
and U3211 (N_3211,N_2821,In_2737);
nand U3212 (N_3212,N_1547,In_4433);
nand U3213 (N_3213,N_2639,In_1825);
and U3214 (N_3214,N_547,N_2544);
xor U3215 (N_3215,N_2859,N_2302);
or U3216 (N_3216,N_2819,N_2627);
and U3217 (N_3217,In_4692,In_732);
xor U3218 (N_3218,N_2712,N_1857);
xor U3219 (N_3219,N_677,In_2373);
nor U3220 (N_3220,In_1349,In_1505);
or U3221 (N_3221,N_1043,In_1382);
xnor U3222 (N_3222,N_2364,N_2591);
nand U3223 (N_3223,N_656,In_4100);
or U3224 (N_3224,In_3090,N_2114);
xnor U3225 (N_3225,N_2322,In_4656);
or U3226 (N_3226,N_7,N_2208);
or U3227 (N_3227,N_895,N_2702);
nor U3228 (N_3228,In_1488,N_2860);
xnor U3229 (N_3229,In_2158,N_2677);
and U3230 (N_3230,In_2422,N_2845);
and U3231 (N_3231,N_1311,N_1394);
xnor U3232 (N_3232,N_1984,In_1368);
or U3233 (N_3233,In_2961,In_3759);
xnor U3234 (N_3234,N_2445,N_2599);
xnor U3235 (N_3235,N_2443,N_320);
xor U3236 (N_3236,In_580,In_519);
or U3237 (N_3237,N_2281,N_75);
xnor U3238 (N_3238,In_4832,N_993);
nor U3239 (N_3239,In_1804,N_2326);
or U3240 (N_3240,In_2304,N_2466);
xnor U3241 (N_3241,N_950,N_1192);
and U3242 (N_3242,In_601,N_2071);
or U3243 (N_3243,N_2202,In_1137);
nor U3244 (N_3244,N_1613,N_1049);
or U3245 (N_3245,In_858,N_2651);
nor U3246 (N_3246,N_679,In_338);
and U3247 (N_3247,N_2185,N_2341);
nand U3248 (N_3248,In_4104,In_3613);
or U3249 (N_3249,In_4548,In_469);
or U3250 (N_3250,N_2091,N_3008);
and U3251 (N_3251,N_554,In_1911);
xnor U3252 (N_3252,In_2826,In_1247);
and U3253 (N_3253,N_3109,In_79);
nand U3254 (N_3254,N_1909,N_2877);
or U3255 (N_3255,N_2047,In_4485);
xor U3256 (N_3256,In_1078,N_1042);
and U3257 (N_3257,N_2791,N_3106);
nand U3258 (N_3258,N_120,In_1667);
and U3259 (N_3259,N_2958,N_1688);
and U3260 (N_3260,In_1031,In_2705);
nand U3261 (N_3261,N_2135,N_2869);
nand U3262 (N_3262,N_1832,N_2925);
xor U3263 (N_3263,N_3094,N_2913);
xnor U3264 (N_3264,N_3239,N_2390);
nand U3265 (N_3265,N_3172,N_2672);
and U3266 (N_3266,N_2810,N_2780);
xnor U3267 (N_3267,N_2131,N_2880);
nand U3268 (N_3268,N_3169,N_2851);
xor U3269 (N_3269,N_927,N_1434);
or U3270 (N_3270,N_842,N_568);
or U3271 (N_3271,N_2166,In_4018);
or U3272 (N_3272,N_2358,In_4073);
nor U3273 (N_3273,In_1925,N_2451);
nor U3274 (N_3274,N_1712,In_2968);
and U3275 (N_3275,In_4785,In_998);
nand U3276 (N_3276,N_3199,In_2743);
xor U3277 (N_3277,In_247,N_2793);
nor U3278 (N_3278,N_3095,N_2975);
nor U3279 (N_3279,In_2741,N_2108);
nor U3280 (N_3280,N_1713,In_2105);
xnor U3281 (N_3281,In_4380,N_2826);
or U3282 (N_3282,In_2237,N_3156);
xor U3283 (N_3283,N_2552,In_4250);
xor U3284 (N_3284,N_2571,N_3249);
xnor U3285 (N_3285,N_945,N_1785);
nor U3286 (N_3286,N_2892,In_4321);
or U3287 (N_3287,In_4739,N_3145);
xnor U3288 (N_3288,N_2650,N_2034);
or U3289 (N_3289,N_2430,N_1429);
nand U3290 (N_3290,In_4105,In_560);
or U3291 (N_3291,N_2573,N_1634);
nand U3292 (N_3292,N_2835,N_1752);
nor U3293 (N_3293,N_2609,N_2956);
xnor U3294 (N_3294,In_375,N_1333);
nand U3295 (N_3295,In_1316,N_1401);
nor U3296 (N_3296,N_3019,N_3133);
xnor U3297 (N_3297,In_3086,N_2773);
or U3298 (N_3298,N_1226,In_383);
nand U3299 (N_3299,N_3244,N_1736);
nand U3300 (N_3300,N_980,In_1315);
or U3301 (N_3301,In_1240,In_672);
nand U3302 (N_3302,N_2954,N_717);
nor U3303 (N_3303,N_2182,N_1804);
and U3304 (N_3304,N_535,N_2549);
nand U3305 (N_3305,N_1175,In_2789);
and U3306 (N_3306,N_2255,N_3230);
nand U3307 (N_3307,N_2883,N_2797);
nor U3308 (N_3308,In_4457,N_2794);
nor U3309 (N_3309,N_2853,N_2990);
nor U3310 (N_3310,In_170,N_793);
or U3311 (N_3311,N_2421,In_554);
nor U3312 (N_3312,In_3654,N_3009);
nor U3313 (N_3313,N_2030,N_1991);
nand U3314 (N_3314,N_2150,In_2827);
nand U3315 (N_3315,N_2752,N_1669);
and U3316 (N_3316,In_3824,N_2889);
xnor U3317 (N_3317,N_30,In_1943);
or U3318 (N_3318,N_3122,In_2111);
and U3319 (N_3319,N_3167,N_786);
or U3320 (N_3320,N_2366,N_2045);
and U3321 (N_3321,N_3215,In_966);
and U3322 (N_3322,N_2906,N_3063);
nand U3323 (N_3323,N_2957,N_2455);
nand U3324 (N_3324,N_3226,N_3241);
and U3325 (N_3325,In_3989,N_2608);
xor U3326 (N_3326,N_463,N_2266);
nand U3327 (N_3327,In_1686,N_2719);
xor U3328 (N_3328,N_2948,N_155);
or U3329 (N_3329,N_1096,N_2567);
nand U3330 (N_3330,In_3285,N_1157);
or U3331 (N_3331,N_2966,In_3393);
nor U3332 (N_3332,N_2981,N_1595);
nor U3333 (N_3333,N_3005,N_2834);
nor U3334 (N_3334,N_2662,N_1392);
and U3335 (N_3335,N_2507,In_171);
or U3336 (N_3336,N_3096,N_2742);
nor U3337 (N_3337,In_1108,In_4565);
nand U3338 (N_3338,In_154,N_2630);
and U3339 (N_3339,N_2844,In_2332);
and U3340 (N_3340,N_2646,N_2548);
and U3341 (N_3341,N_2769,N_1614);
and U3342 (N_3342,N_2775,N_3065);
nand U3343 (N_3343,N_2292,N_1858);
and U3344 (N_3344,N_374,In_244);
xor U3345 (N_3345,In_1210,In_1645);
nor U3346 (N_3346,N_3023,In_4703);
and U3347 (N_3347,N_3101,N_2937);
or U3348 (N_3348,N_2572,In_3938);
or U3349 (N_3349,N_1877,N_2209);
or U3350 (N_3350,N_1378,N_2885);
and U3351 (N_3351,In_2975,N_2644);
xor U3352 (N_3352,N_2720,N_3090);
nand U3353 (N_3353,N_2977,N_221);
and U3354 (N_3354,In_694,N_2408);
xor U3355 (N_3355,N_2953,In_3997);
nand U3356 (N_3356,N_2643,N_103);
and U3357 (N_3357,N_2492,N_2086);
nand U3358 (N_3358,In_3523,N_3157);
nor U3359 (N_3359,N_2310,N_2766);
and U3360 (N_3360,In_4174,N_1540);
nor U3361 (N_3361,N_2917,In_799);
nor U3362 (N_3362,N_3010,In_1132);
nand U3363 (N_3363,N_2736,N_3245);
nor U3364 (N_3364,In_4733,N_3085);
and U3365 (N_3365,N_982,In_3137);
nand U3366 (N_3366,In_418,In_4836);
xnor U3367 (N_3367,N_3184,N_2056);
nor U3368 (N_3368,N_1553,In_1496);
nand U3369 (N_3369,N_294,In_3968);
or U3370 (N_3370,N_2803,In_2116);
or U3371 (N_3371,N_2947,N_2706);
and U3372 (N_3372,In_3786,N_2740);
nand U3373 (N_3373,In_1233,In_3894);
and U3374 (N_3374,N_2784,N_3170);
or U3375 (N_3375,N_3072,N_437);
or U3376 (N_3376,In_4048,N_70);
or U3377 (N_3377,N_3165,In_4082);
or U3378 (N_3378,N_844,N_2693);
and U3379 (N_3379,In_3273,In_2830);
or U3380 (N_3380,N_2129,N_2244);
xnor U3381 (N_3381,N_2804,In_3159);
nand U3382 (N_3382,N_3151,N_837);
and U3383 (N_3383,N_1064,In_1905);
nor U3384 (N_3384,In_3879,In_2081);
or U3385 (N_3385,In_4765,N_1201);
and U3386 (N_3386,N_3076,N_2454);
nor U3387 (N_3387,N_1581,In_685);
or U3388 (N_3388,N_3207,N_2336);
nand U3389 (N_3389,In_1581,N_3037);
and U3390 (N_3390,N_918,N_3062);
and U3391 (N_3391,N_3036,In_2360);
xor U3392 (N_3392,In_4035,N_3227);
nand U3393 (N_3393,N_14,N_1817);
or U3394 (N_3394,In_2216,N_2475);
or U3395 (N_3395,In_933,In_1399);
xor U3396 (N_3396,In_2812,In_757);
or U3397 (N_3397,In_2970,N_2124);
or U3398 (N_3398,N_3211,In_70);
nor U3399 (N_3399,N_2841,In_1560);
nor U3400 (N_3400,N_1847,N_2199);
and U3401 (N_3401,In_285,In_1460);
xnor U3402 (N_3402,N_2073,N_2908);
nor U3403 (N_3403,In_3021,In_498);
and U3404 (N_3404,In_2856,N_2904);
and U3405 (N_3405,N_2959,N_2396);
nand U3406 (N_3406,N_2994,N_2491);
and U3407 (N_3407,N_1383,N_2272);
nand U3408 (N_3408,In_2861,In_3884);
and U3409 (N_3409,N_2337,In_2478);
and U3410 (N_3410,In_2068,N_1449);
xnor U3411 (N_3411,In_2824,N_1989);
or U3412 (N_3412,N_2750,N_2286);
or U3413 (N_3413,In_4264,N_1419);
or U3414 (N_3414,N_3203,N_3079);
nand U3415 (N_3415,In_1268,N_1979);
nor U3416 (N_3416,N_1605,In_2007);
nor U3417 (N_3417,N_2039,N_626);
and U3418 (N_3418,N_2403,N_1915);
or U3419 (N_3419,In_3640,N_3190);
nor U3420 (N_3420,In_1254,N_2496);
nand U3421 (N_3421,N_1346,In_713);
or U3422 (N_3422,N_3137,N_2420);
nor U3423 (N_3423,N_1505,N_1820);
nor U3424 (N_3424,N_2999,N_2602);
or U3425 (N_3425,N_1956,N_3103);
or U3426 (N_3426,N_3219,N_2909);
nand U3427 (N_3427,N_3231,In_2819);
nor U3428 (N_3428,N_1512,N_203);
or U3429 (N_3429,In_1586,In_4294);
or U3430 (N_3430,N_2876,N_1967);
nand U3431 (N_3431,N_1455,In_4437);
nor U3432 (N_3432,N_2918,In_1676);
xor U3433 (N_3433,In_1730,N_2048);
or U3434 (N_3434,N_1685,N_2062);
xor U3435 (N_3435,In_454,In_2591);
nand U3436 (N_3436,N_2031,N_3150);
xnor U3437 (N_3437,In_4817,N_2899);
xnor U3438 (N_3438,N_2827,N_1871);
nand U3439 (N_3439,In_2056,In_3966);
nor U3440 (N_3440,N_2864,N_2714);
nand U3441 (N_3441,In_1333,N_2694);
xor U3442 (N_3442,In_2503,N_2661);
or U3443 (N_3443,N_1395,In_169);
xor U3444 (N_3444,In_4720,In_2682);
or U3445 (N_3445,N_1705,In_2621);
nor U3446 (N_3446,N_2997,In_4748);
xnor U3447 (N_3447,N_897,In_3312);
nand U3448 (N_3448,In_2616,N_2652);
xnor U3449 (N_3449,N_2351,In_2674);
and U3450 (N_3450,In_597,N_2761);
or U3451 (N_3451,N_2978,In_1959);
xor U3452 (N_3452,N_1339,N_1015);
nand U3453 (N_3453,N_284,N_2223);
xnor U3454 (N_3454,N_2867,N_361);
nand U3455 (N_3455,N_2731,In_2211);
and U3456 (N_3456,N_2268,In_4754);
nand U3457 (N_3457,N_3222,N_1676);
nand U3458 (N_3458,N_1330,N_1702);
xnor U3459 (N_3459,N_110,N_922);
nand U3460 (N_3460,N_1763,N_1393);
or U3461 (N_3461,N_589,In_1652);
xnor U3462 (N_3462,N_1620,N_2253);
xor U3463 (N_3463,In_583,N_1391);
xnor U3464 (N_3464,N_1665,N_3129);
nand U3465 (N_3465,N_3098,N_2607);
nand U3466 (N_3466,In_1417,N_3108);
and U3467 (N_3467,N_1530,N_2405);
nor U3468 (N_3468,N_3049,N_2083);
nor U3469 (N_3469,In_4568,In_2891);
nand U3470 (N_3470,N_577,N_601);
xnor U3471 (N_3471,In_3991,In_2548);
nor U3472 (N_3472,N_195,In_3757);
and U3473 (N_3473,N_641,In_3413);
nand U3474 (N_3474,N_2546,In_2471);
or U3475 (N_3475,N_1879,In_1452);
nor U3476 (N_3476,In_4738,N_3185);
xnor U3477 (N_3477,N_2890,N_1882);
or U3478 (N_3478,N_1711,N_3007);
or U3479 (N_3479,In_4351,N_2732);
xor U3480 (N_3480,N_1629,N_2995);
nand U3481 (N_3481,In_2726,N_3030);
xor U3482 (N_3482,N_1710,N_2976);
or U3483 (N_3483,N_587,N_1865);
nor U3484 (N_3484,In_908,N_2508);
nand U3485 (N_3485,N_3246,In_575);
nor U3486 (N_3486,In_1697,N_978);
nor U3487 (N_3487,N_1823,N_2690);
xnor U3488 (N_3488,In_2445,N_1913);
or U3489 (N_3489,In_4563,N_3039);
nand U3490 (N_3490,In_180,In_4495);
xor U3491 (N_3491,N_2631,In_4247);
xor U3492 (N_3492,N_525,N_1646);
xor U3493 (N_3493,N_1207,N_3139);
nand U3494 (N_3494,N_315,N_2878);
and U3495 (N_3495,N_3208,N_3191);
nand U3496 (N_3496,N_2696,N_2194);
or U3497 (N_3497,N_3034,N_1129);
nand U3498 (N_3498,N_1801,N_2764);
nand U3499 (N_3499,N_2422,In_3771);
nand U3500 (N_3500,In_815,N_2147);
xnor U3501 (N_3501,N_2138,In_1461);
and U3502 (N_3502,N_3088,N_2792);
and U3503 (N_3503,N_3465,N_3112);
xnor U3504 (N_3504,N_2537,N_2785);
nor U3505 (N_3505,N_2809,N_2941);
nand U3506 (N_3506,N_2983,N_3447);
and U3507 (N_3507,N_3323,In_1664);
and U3508 (N_3508,N_2936,In_2298);
and U3509 (N_3509,N_2871,In_3193);
nand U3510 (N_3510,N_875,In_1290);
nand U3511 (N_3511,In_1455,N_2974);
nor U3512 (N_3512,N_1232,N_3406);
nor U3513 (N_3513,In_731,In_2225);
or U3514 (N_3514,N_1959,In_356);
or U3515 (N_3515,N_3297,N_3484);
and U3516 (N_3516,N_2746,N_491);
and U3517 (N_3517,N_3038,N_3093);
and U3518 (N_3518,N_2625,In_680);
xnor U3519 (N_3519,N_2395,N_3011);
nand U3520 (N_3520,N_3240,N_347);
and U3521 (N_3521,N_806,N_3148);
or U3522 (N_3522,N_3432,N_3302);
nor U3523 (N_3523,N_2377,N_2133);
nor U3524 (N_3524,N_1020,N_3453);
nand U3525 (N_3525,In_3222,N_3216);
nand U3526 (N_3526,N_2164,N_2806);
nor U3527 (N_3527,In_4089,N_3257);
xor U3528 (N_3528,In_4606,N_2824);
nor U3529 (N_3529,N_2484,N_3311);
xor U3530 (N_3530,N_2059,N_891);
and U3531 (N_3531,N_2469,In_3748);
xor U3532 (N_3532,In_3552,N_3330);
and U3533 (N_3533,N_2529,N_3368);
nor U3534 (N_3534,In_978,In_2055);
nand U3535 (N_3535,N_2128,N_3056);
or U3536 (N_3536,In_3918,N_2204);
and U3537 (N_3537,N_337,N_2462);
xor U3538 (N_3538,In_4334,N_2380);
nor U3539 (N_3539,In_1736,In_1229);
nand U3540 (N_3540,N_3232,N_1291);
or U3541 (N_3541,N_2596,N_3074);
nor U3542 (N_3542,N_1217,N_3031);
nor U3543 (N_3543,N_3182,N_3025);
xor U3544 (N_3544,N_3242,N_2967);
or U3545 (N_3545,N_45,In_3817);
nor U3546 (N_3546,N_2558,In_4541);
xor U3547 (N_3547,N_1555,N_1603);
and U3548 (N_3548,N_2815,N_1737);
and U3549 (N_3549,N_2532,N_2888);
nor U3550 (N_3550,In_962,In_3836);
nor U3551 (N_3551,In_1419,N_3044);
nor U3552 (N_3552,N_1518,N_2725);
nand U3553 (N_3553,N_1881,N_2531);
or U3554 (N_3554,N_1128,N_2817);
or U3555 (N_3555,In_3995,In_3932);
or U3556 (N_3556,N_1133,N_2015);
xor U3557 (N_3557,N_55,N_2861);
nand U3558 (N_3558,N_3186,N_2965);
nand U3559 (N_3559,N_2748,N_3442);
xnor U3560 (N_3560,N_2692,N_1373);
nand U3561 (N_3561,In_939,N_2423);
xor U3562 (N_3562,N_3418,N_3341);
xnor U3563 (N_3563,In_2623,N_3033);
or U3564 (N_3564,N_1457,N_3365);
xor U3565 (N_3565,N_983,N_192);
or U3566 (N_3566,N_942,N_2252);
nor U3567 (N_3567,In_3076,N_2570);
or U3568 (N_3568,In_3155,N_2501);
nor U3569 (N_3569,N_3201,In_4967);
and U3570 (N_3570,N_2388,N_2879);
or U3571 (N_3571,N_2711,N_3456);
and U3572 (N_3572,In_1776,N_2066);
xnor U3573 (N_3573,N_3401,In_1914);
nor U3574 (N_3574,N_2710,N_2653);
nor U3575 (N_3575,N_2282,In_1796);
and U3576 (N_3576,In_3994,N_1427);
nand U3577 (N_3577,N_3205,N_3162);
nor U3578 (N_3578,In_3417,N_1521);
nor U3579 (N_3579,N_3195,N_3324);
or U3580 (N_3580,In_3889,N_1917);
xor U3581 (N_3581,N_2593,N_2698);
and U3582 (N_3582,N_1762,N_2985);
nor U3583 (N_3583,N_3123,N_1781);
xor U3584 (N_3584,N_3413,N_2969);
and U3585 (N_3585,In_57,N_2125);
xnor U3586 (N_3586,N_2375,N_3408);
and U3587 (N_3587,In_4869,N_3197);
nand U3588 (N_3588,In_3425,In_355);
or U3589 (N_3589,N_2427,N_3352);
xor U3590 (N_3590,N_3428,N_2767);
or U3591 (N_3591,N_948,N_2814);
nor U3592 (N_3592,N_2584,N_59);
nor U3593 (N_3593,N_3086,N_3420);
nor U3594 (N_3594,N_2068,In_35);
nor U3595 (N_3595,N_3472,N_3357);
and U3596 (N_3596,N_3064,N_2533);
xor U3597 (N_3597,N_3303,N_3210);
and U3598 (N_3598,In_4320,In_3557);
nor U3599 (N_3599,N_2181,N_3391);
nand U3600 (N_3600,In_3116,N_3171);
or U3601 (N_3601,N_2353,N_1545);
nand U3602 (N_3602,N_101,N_2032);
nand U3603 (N_3603,N_3419,N_3067);
xor U3604 (N_3604,N_3289,N_2510);
nand U3605 (N_3605,N_2615,N_172);
nand U3606 (N_3606,N_1771,N_3223);
nand U3607 (N_3607,In_3902,N_3355);
nand U3608 (N_3608,N_2437,N_1490);
or U3609 (N_3609,In_2696,N_1148);
nor U3610 (N_3610,N_3127,N_3021);
nand U3611 (N_3611,N_2722,N_770);
xor U3612 (N_3612,In_2964,N_3492);
nand U3613 (N_3613,N_2118,N_154);
and U3614 (N_3614,N_2798,In_1314);
nor U3615 (N_3615,N_2080,N_2665);
and U3616 (N_3616,N_3069,N_3212);
and U3617 (N_3617,In_4188,N_2516);
xnor U3618 (N_3618,N_1400,N_617);
nand U3619 (N_3619,N_3066,N_2480);
xor U3620 (N_3620,In_1585,N_878);
or U3621 (N_3621,N_1815,N_2234);
or U3622 (N_3622,N_3471,In_2204);
nand U3623 (N_3623,N_2301,N_1083);
nor U3624 (N_3624,In_4199,N_3433);
nand U3625 (N_3625,N_3295,N_2356);
nand U3626 (N_3626,N_249,N_230);
and U3627 (N_3627,N_2986,In_3861);
or U3628 (N_3628,N_3385,N_2504);
and U3629 (N_3629,N_1894,In_3660);
nand U3630 (N_3630,N_2923,N_3015);
nor U3631 (N_3631,In_2628,N_3073);
nor U3632 (N_3632,N_476,N_2931);
nor U3633 (N_3633,N_2563,In_1005);
and U3634 (N_3634,N_1886,N_2898);
nor U3635 (N_3635,N_3002,In_4449);
nand U3636 (N_3636,N_1039,In_2778);
or U3637 (N_3637,N_3425,N_3327);
nor U3638 (N_3638,N_2509,N_2961);
and U3639 (N_3639,N_3378,In_3519);
xor U3640 (N_3640,In_3422,N_2852);
and U3641 (N_3641,N_1878,N_2624);
or U3642 (N_3642,N_3270,N_3298);
and U3643 (N_3643,N_3177,N_2344);
or U3644 (N_3644,N_2697,N_3141);
nand U3645 (N_3645,N_3449,N_1891);
and U3646 (N_3646,N_1590,N_3269);
and U3647 (N_3647,N_2308,N_1598);
or U3648 (N_3648,N_1830,In_2196);
xnor U3649 (N_3649,In_3131,In_2233);
nand U3650 (N_3650,N_2535,In_4644);
nand U3651 (N_3651,N_1800,N_3029);
nand U3652 (N_3652,In_4808,In_3567);
or U3653 (N_3653,N_3138,In_4776);
or U3654 (N_3654,In_1173,N_1492);
xor U3655 (N_3655,N_2550,In_1794);
nand U3656 (N_3656,N_2163,In_4727);
and U3657 (N_3657,N_2754,N_1585);
or U3658 (N_3658,N_3124,In_2153);
nor U3659 (N_3659,N_780,N_2093);
nor U3660 (N_3660,N_3273,N_2816);
or U3661 (N_3661,In_1998,In_3451);
xnor U3662 (N_3662,In_2512,In_2);
nand U3663 (N_3663,N_2921,In_3484);
or U3664 (N_3664,N_460,N_2426);
nor U3665 (N_3665,N_1957,N_3434);
xnor U3666 (N_3666,N_1037,N_3181);
or U3667 (N_3667,N_465,N_2887);
nand U3668 (N_3668,N_2119,N_3265);
or U3669 (N_3669,N_1708,N_213);
nor U3670 (N_3670,N_3444,N_1583);
nor U3671 (N_3671,N_2787,In_1978);
nand U3672 (N_3672,N_905,In_3257);
or U3673 (N_3673,N_2211,N_1266);
nor U3674 (N_3674,N_3022,In_11);
nor U3675 (N_3675,N_3192,N_3309);
nand U3676 (N_3676,N_1399,In_3008);
and U3677 (N_3677,In_1865,N_961);
xnor U3678 (N_3678,N_2636,In_1593);
or U3679 (N_3679,N_223,N_3328);
or U3680 (N_3680,N_3452,In_4275);
nand U3681 (N_3681,In_4029,N_506);
nor U3682 (N_3682,N_3443,In_4879);
xor U3683 (N_3683,N_660,N_1884);
or U3684 (N_3684,N_3358,N_1044);
xnor U3685 (N_3685,N_3480,N_2781);
xnor U3686 (N_3686,In_1733,N_2242);
and U3687 (N_3687,N_1859,In_217);
nand U3688 (N_3688,N_3496,In_2151);
or U3689 (N_3689,N_3334,In_2501);
nand U3690 (N_3690,In_2219,N_2649);
nand U3691 (N_3691,N_3200,In_3713);
or U3692 (N_3692,N_3314,N_3179);
xnor U3693 (N_3693,N_3164,N_3499);
and U3694 (N_3694,N_3168,N_3250);
or U3695 (N_3695,N_3481,N_676);
xor U3696 (N_3696,In_4358,N_3189);
or U3697 (N_3697,N_1550,N_2518);
and U3698 (N_3698,N_2075,N_1498);
xnor U3699 (N_3699,N_3390,In_3874);
nor U3700 (N_3700,N_3140,N_3259);
xor U3701 (N_3701,In_417,In_871);
and U3702 (N_3702,N_1998,N_2305);
and U3703 (N_3703,N_2559,N_2278);
xnor U3704 (N_3704,N_1413,N_3131);
or U3705 (N_3705,N_305,N_2259);
and U3706 (N_3706,N_740,N_3326);
and U3707 (N_3707,N_1824,N_1872);
nor U3708 (N_3708,N_2734,N_3473);
nor U3709 (N_3709,N_3440,In_1900);
or U3710 (N_3710,N_3349,In_548);
nor U3711 (N_3711,In_4434,In_2920);
or U3712 (N_3712,N_2489,N_1706);
or U3713 (N_3713,In_2857,N_3448);
nand U3714 (N_3714,N_2172,In_4255);
or U3715 (N_3715,In_4225,N_1607);
xor U3716 (N_3716,N_3217,N_3238);
or U3717 (N_3717,N_3213,N_2808);
nor U3718 (N_3718,N_3052,In_2238);
or U3719 (N_3719,N_3376,N_3366);
or U3720 (N_3720,N_2157,N_1704);
nand U3721 (N_3721,In_3111,N_3409);
xor U3722 (N_3722,N_2225,N_2838);
nor U3723 (N_3723,N_2406,N_3284);
and U3724 (N_3724,N_3415,N_2949);
and U3725 (N_3725,N_3441,N_3359);
and U3726 (N_3726,In_2487,In_4517);
nor U3727 (N_3727,N_2077,In_4573);
and U3728 (N_3728,N_2942,N_2922);
nand U3729 (N_3729,N_1846,N_266);
and U3730 (N_3730,N_2996,N_778);
or U3731 (N_3731,N_3110,N_3454);
nand U3732 (N_3732,N_3092,N_1965);
nand U3733 (N_3733,N_1279,In_1610);
nor U3734 (N_3734,N_2759,N_3234);
xor U3735 (N_3735,N_2530,In_3510);
or U3736 (N_3736,N_3339,In_3922);
nand U3737 (N_3737,In_1109,N_9);
or U3738 (N_3738,N_308,In_4782);
nand U3739 (N_3739,N_397,N_3178);
and U3740 (N_3740,In_1957,N_2862);
nor U3741 (N_3741,N_2679,In_3802);
or U3742 (N_3742,N_443,N_3294);
or U3743 (N_3743,N_2848,N_3374);
nor U3744 (N_3744,N_1290,N_3204);
nand U3745 (N_3745,N_2856,N_3460);
nand U3746 (N_3746,N_3435,In_4110);
nor U3747 (N_3747,N_58,In_1122);
and U3748 (N_3748,N_3255,N_3486);
and U3749 (N_3749,N_1844,N_1504);
xor U3750 (N_3750,N_3679,In_808);
and U3751 (N_3751,N_2945,In_160);
or U3752 (N_3752,N_3618,N_3388);
xor U3753 (N_3753,N_1764,N_2920);
and U3754 (N_3754,N_3235,N_2494);
and U3755 (N_3755,N_1606,N_2756);
nand U3756 (N_3756,N_218,In_4028);
nor U3757 (N_3757,N_2431,N_3635);
xor U3758 (N_3758,N_2726,N_2325);
xnor U3759 (N_3759,N_3194,N_3081);
xnor U3760 (N_3760,N_3237,In_4827);
xnor U3761 (N_3761,N_2595,N_3500);
or U3762 (N_3762,N_2855,In_276);
nor U3763 (N_3763,N_622,In_3136);
nor U3764 (N_3764,N_2576,N_1854);
nand U3765 (N_3765,N_3669,N_1166);
and U3766 (N_3766,N_2737,In_3048);
nor U3767 (N_3767,N_2527,N_2280);
nor U3768 (N_3768,N_3641,N_3602);
nand U3769 (N_3769,N_3593,N_572);
or U3770 (N_3770,In_1224,N_2735);
and U3771 (N_3771,N_1876,In_352);
nand U3772 (N_3772,N_1628,In_4671);
nand U3773 (N_3773,N_1893,N_3583);
or U3774 (N_3774,N_3279,N_3301);
or U3775 (N_3775,In_2873,In_67);
or U3776 (N_3776,In_4611,N_2628);
nor U3777 (N_3777,N_3649,N_3305);
nor U3778 (N_3778,N_3146,N_3028);
nor U3779 (N_3779,In_2232,In_1213);
and U3780 (N_3780,N_1190,N_3483);
nand U3781 (N_3781,N_3107,N_2926);
and U3782 (N_3782,N_3567,In_912);
nand U3783 (N_3783,N_3654,N_3535);
xnor U3784 (N_3784,In_2062,N_3596);
nor U3785 (N_3785,N_3476,N_2666);
xnor U3786 (N_3786,N_2007,In_3254);
or U3787 (N_3787,N_3431,N_3503);
and U3788 (N_3788,N_3676,N_2776);
nor U3789 (N_3789,In_2954,In_4639);
nor U3790 (N_3790,N_2583,N_3264);
or U3791 (N_3791,N_1912,N_3696);
nand U3792 (N_3792,N_420,In_3225);
or U3793 (N_3793,N_354,N_3153);
or U3794 (N_3794,In_2648,N_3014);
and U3795 (N_3795,N_1533,In_1579);
or U3796 (N_3796,N_1410,N_428);
nor U3797 (N_3797,In_2372,In_4410);
nor U3798 (N_3798,In_1193,N_3531);
nor U3799 (N_3799,N_2121,N_3707);
nand U3800 (N_3800,In_2292,N_3262);
nor U3801 (N_3801,In_1101,N_2622);
or U3802 (N_3802,N_3651,N_2950);
nand U3803 (N_3803,In_550,N_2895);
or U3804 (N_3804,N_3024,N_3152);
xnor U3805 (N_3805,In_2546,N_3533);
xor U3806 (N_3806,In_2368,N_2347);
nand U3807 (N_3807,N_3570,N_3429);
or U3808 (N_3808,N_3657,N_2707);
nor U3809 (N_3809,N_2893,N_1531);
nand U3810 (N_3810,N_3603,N_3513);
and U3811 (N_3811,N_3490,In_2924);
xor U3812 (N_3812,N_3693,N_3622);
nor U3813 (N_3813,N_3315,In_1899);
and U3814 (N_3814,N_3482,N_1890);
xnor U3815 (N_3815,N_3479,N_3625);
xor U3816 (N_3816,N_3532,N_2802);
xor U3817 (N_3817,In_1642,N_1363);
xnor U3818 (N_3818,N_3310,N_3395);
nand U3819 (N_3819,In_3338,N_2515);
nand U3820 (N_3820,N_3658,N_1922);
and U3821 (N_3821,In_3780,N_3688);
or U3822 (N_3822,N_3523,N_3026);
nor U3823 (N_3823,N_2486,N_2369);
or U3824 (N_3824,N_754,N_3749);
nor U3825 (N_3825,In_3522,N_3489);
nor U3826 (N_3826,N_377,N_3516);
nor U3827 (N_3827,N_2428,In_648);
nor U3828 (N_3828,N_3597,N_3439);
xnor U3829 (N_3829,N_71,N_3554);
or U3830 (N_3830,N_3573,N_1920);
and U3831 (N_3831,In_1485,N_3048);
and U3832 (N_3832,N_2378,N_3020);
nand U3833 (N_3833,N_2193,N_2498);
xnor U3834 (N_3834,N_2536,N_2348);
nand U3835 (N_3835,N_490,N_665);
nor U3836 (N_3836,N_3542,In_2586);
nor U3837 (N_3837,N_2708,N_3467);
or U3838 (N_3838,N_2929,N_892);
or U3839 (N_3839,N_3053,N_3398);
xnor U3840 (N_3840,N_2295,N_3099);
and U3841 (N_3841,N_3508,N_3740);
and U3842 (N_3842,N_1962,N_1812);
nor U3843 (N_3843,N_2404,N_1870);
and U3844 (N_3844,N_3470,N_3650);
xor U3845 (N_3845,N_3714,N_2542);
xnor U3846 (N_3846,N_1942,N_2779);
and U3847 (N_3847,N_2724,In_2318);
xnor U3848 (N_3848,N_2158,In_1673);
or U3849 (N_3849,In_899,N_217);
or U3850 (N_3850,N_3662,In_2401);
nand U3851 (N_3851,In_3524,In_1190);
and U3852 (N_3852,N_3159,In_2268);
nor U3853 (N_3853,In_4200,In_3911);
xor U3854 (N_3854,N_3493,In_196);
or U3855 (N_3855,In_4929,N_3682);
nand U3856 (N_3856,N_3691,N_2367);
or U3857 (N_3857,N_530,In_1660);
xnor U3858 (N_3858,N_1862,In_4416);
nor U3859 (N_3859,N_3417,N_3719);
nor U3860 (N_3860,N_2782,N_3361);
nor U3861 (N_3861,N_2786,N_1694);
nor U3862 (N_3862,In_833,N_3125);
nor U3863 (N_3863,N_908,N_3130);
or U3864 (N_3864,N_2023,N_2116);
nand U3865 (N_3865,N_1951,N_3741);
nand U3866 (N_3866,N_2270,N_3715);
or U3867 (N_3867,N_3610,N_1697);
or U3868 (N_3868,N_3027,N_3474);
nor U3869 (N_3869,N_3609,In_2647);
nand U3870 (N_3870,In_4243,N_3253);
nand U3871 (N_3871,N_3166,N_3529);
or U3872 (N_3872,N_2687,N_2190);
or U3873 (N_3873,N_2151,N_2774);
xnor U3874 (N_3874,N_3605,N_3576);
and U3875 (N_3875,N_1436,N_3477);
xor U3876 (N_3876,In_1117,N_2749);
or U3877 (N_3877,In_2340,N_2429);
or U3878 (N_3878,N_3461,N_3236);
nand U3879 (N_3879,N_651,N_2594);
xor U3880 (N_3880,N_2393,N_3717);
and U3881 (N_3881,In_4079,N_3091);
and U3882 (N_3882,N_3317,In_2564);
nand U3883 (N_3883,N_3667,In_4364);
nor U3884 (N_3884,N_967,N_3188);
and U3885 (N_3885,In_3927,N_3515);
or U3886 (N_3886,N_3723,N_3040);
nor U3887 (N_3887,In_3029,N_1294);
xor U3888 (N_3888,N_3626,N_82);
xnor U3889 (N_3889,N_3394,N_3060);
or U3890 (N_3890,N_3506,N_3530);
xnor U3891 (N_3891,In_4488,N_2905);
nand U3892 (N_3892,N_2224,N_3332);
nand U3893 (N_3893,N_2678,N_2654);
and U3894 (N_3894,In_3456,N_3620);
xor U3895 (N_3895,N_3252,N_3745);
or U3896 (N_3896,N_2963,N_2934);
xnor U3897 (N_3897,In_3221,N_2840);
xor U3898 (N_3898,N_2988,N_1887);
xor U3899 (N_3899,N_1468,In_4598);
nor U3900 (N_3900,In_4792,N_3643);
and U3901 (N_3901,In_2540,N_3504);
and U3902 (N_3902,In_1856,In_3240);
and U3903 (N_3903,N_3697,N_3307);
nor U3904 (N_3904,In_4552,N_3337);
xnor U3905 (N_3905,N_2902,N_3321);
nand U3906 (N_3906,N_3360,N_3117);
and U3907 (N_3907,N_2565,N_3661);
nor U3908 (N_3908,In_4126,N_3116);
and U3909 (N_3909,N_1751,In_4943);
xnor U3910 (N_3910,N_3671,N_2882);
and U3911 (N_3911,In_3102,N_3747);
or U3912 (N_3912,In_248,N_3640);
or U3913 (N_3913,N_3505,N_3621);
nor U3914 (N_3914,N_3612,N_1987);
nand U3915 (N_3915,In_4401,N_2717);
xnor U3916 (N_3916,In_2347,N_3436);
nand U3917 (N_3917,N_2648,N_1927);
or U3918 (N_3918,N_3607,N_3142);
xnor U3919 (N_3919,N_3363,N_2499);
nand U3920 (N_3920,N_1829,N_3600);
xor U3921 (N_3921,N_3585,N_2514);
xor U3922 (N_3922,N_2145,N_2980);
nor U3923 (N_3923,N_2778,N_3519);
or U3924 (N_3924,N_3070,N_2795);
nor U3925 (N_3925,In_935,N_2241);
nor U3926 (N_3926,N_3043,In_187);
xnor U3927 (N_3927,N_3639,N_3512);
nor U3928 (N_3928,N_0,N_3224);
or U3929 (N_3929,In_540,N_3336);
or U3930 (N_3930,N_3744,In_1534);
nand U3931 (N_3931,N_3271,N_1067);
xnor U3932 (N_3932,N_3459,N_1234);
nand U3933 (N_3933,N_3149,N_3501);
nand U3934 (N_3934,N_2122,In_4977);
xnor U3935 (N_3935,N_3457,N_3498);
nor U3936 (N_3936,N_1202,N_1295);
nor U3937 (N_3937,In_1060,N_2686);
nand U3938 (N_3938,N_2972,N_3082);
nand U3939 (N_3939,In_3851,N_3126);
and U3940 (N_3940,In_3058,In_810);
xor U3941 (N_3941,In_3564,N_3574);
or U3942 (N_3942,N_2545,N_3382);
xor U3943 (N_3943,N_2718,In_3784);
xnor U3944 (N_3944,N_3630,N_3491);
or U3945 (N_3945,N_2391,In_3307);
nand U3946 (N_3946,N_2012,In_4934);
xnor U3947 (N_3947,N_3059,N_3353);
xnor U3948 (N_3948,In_358,N_3710);
nor U3949 (N_3949,N_2055,N_2638);
xor U3950 (N_3950,N_123,In_1977);
nor U3951 (N_3951,N_2626,N_684);
xnor U3952 (N_3952,In_1637,In_249);
xor U3953 (N_3953,In_4148,N_3389);
nor U3954 (N_3954,N_2328,N_2751);
nor U3955 (N_3955,N_3280,N_3312);
or U3956 (N_3956,In_2309,In_2419);
xor U3957 (N_3957,N_3742,In_956);
xnor U3958 (N_3958,N_3128,N_2865);
and U3959 (N_3959,N_2657,N_2011);
and U3960 (N_3960,N_1537,N_1730);
or U3961 (N_3961,N_3701,N_2547);
or U3962 (N_3962,N_3681,N_3437);
or U3963 (N_3963,In_3766,N_3160);
or U3964 (N_3964,N_2590,N_2521);
xnor U3965 (N_3965,N_3320,In_4893);
nor U3966 (N_3966,In_4861,N_3592);
nor U3967 (N_3967,N_2837,N_3281);
and U3968 (N_3968,N_2805,N_3656);
xnor U3969 (N_3969,N_3143,N_3041);
or U3970 (N_3970,N_3595,In_3016);
xor U3971 (N_3971,N_3083,In_769);
nor U3972 (N_3972,In_4168,N_3261);
xnor U3973 (N_3973,N_1969,N_3243);
nand U3974 (N_3974,N_2843,In_256);
or U3975 (N_3975,N_764,N_3673);
xnor U3976 (N_3976,N_3193,N_3229);
nor U3977 (N_3977,N_3343,N_2828);
xor U3978 (N_3978,N_3410,N_3426);
nor U3979 (N_3979,In_2708,In_4310);
and U3980 (N_3980,N_1303,N_2830);
or U3981 (N_3981,In_346,In_724);
and U3982 (N_3982,N_3202,N_3608);
nor U3983 (N_3983,N_3724,N_1032);
xnor U3984 (N_3984,N_3663,N_3047);
nand U3985 (N_3985,N_3345,In_4569);
or U3986 (N_3986,In_2585,N_1866);
nand U3987 (N_3987,N_3527,In_3969);
and U3988 (N_3988,N_2585,In_2038);
nand U3989 (N_3989,N_2903,N_1601);
xor U3990 (N_3990,N_3522,N_1305);
nand U3991 (N_3991,In_1847,N_3689);
nor U3992 (N_3992,N_1948,N_3003);
nor U3993 (N_3993,N_3502,N_2327);
or U3994 (N_3994,N_2568,N_2783);
and U3995 (N_3995,N_3313,In_990);
and U3996 (N_3996,N_3455,N_3734);
or U3997 (N_3997,In_123,N_3300);
and U3998 (N_3998,In_3175,N_1122);
nor U3999 (N_3999,N_3478,N_2993);
nand U4000 (N_4000,In_3478,N_3422);
or U4001 (N_4001,In_2467,In_2327);
nor U4002 (N_4002,N_3699,N_3214);
and U4003 (N_4003,N_3400,N_3892);
nand U4004 (N_4004,N_3526,In_4067);
or U4005 (N_4005,N_3584,N_3648);
and U4006 (N_4006,N_3922,N_3611);
nand U4007 (N_4007,N_3989,N_3628);
nand U4008 (N_4008,N_3286,N_3863);
or U4009 (N_4009,N_3844,N_3861);
nand U4010 (N_4010,N_3826,In_4767);
xor U4011 (N_4011,N_3571,N_40);
nand U4012 (N_4012,N_3316,N_2315);
nor U4013 (N_4013,N_3925,In_3276);
or U4014 (N_4014,N_3970,N_3852);
nor U4015 (N_4015,N_3928,N_1056);
and U4016 (N_4016,N_3154,N_3812);
or U4017 (N_4017,N_1836,N_528);
nand U4018 (N_4018,In_3684,N_3726);
nor U4019 (N_4019,In_737,N_3354);
or U4020 (N_4020,N_2919,N_3268);
or U4021 (N_4021,N_2801,N_3118);
and U4022 (N_4022,N_1310,In_4036);
nor U4023 (N_4023,In_504,N_3713);
nand U4024 (N_4024,N_3674,N_1919);
xor U4025 (N_4025,N_3939,N_3735);
or U4026 (N_4026,N_3111,In_2750);
nor U4027 (N_4027,N_2028,N_3176);
or U4028 (N_4028,N_2256,N_3911);
and U4029 (N_4029,N_3858,In_4010);
or U4030 (N_4030,N_3104,N_3704);
nand U4031 (N_4031,N_3274,N_1163);
xnor U4032 (N_4032,N_3134,N_3487);
nor U4033 (N_4033,N_3854,N_1783);
nor U4034 (N_4034,N_3100,N_3845);
or U4035 (N_4035,N_3933,N_3732);
xnor U4036 (N_4036,N_3809,N_29);
or U4037 (N_4037,N_3818,N_3132);
or U4038 (N_4038,N_3736,N_3319);
or U4039 (N_4039,N_3581,In_1414);
and U4040 (N_4040,N_3746,N_810);
and U4041 (N_4041,In_1965,N_2897);
nor U4042 (N_4042,N_2620,N_3947);
and U4043 (N_4043,N_3057,N_3807);
or U4044 (N_4044,N_3796,N_3275);
xnor U4045 (N_4045,N_3771,N_149);
or U4046 (N_4046,N_1652,N_2641);
and U4047 (N_4047,N_2613,N_3777);
xnor U4048 (N_4048,N_2476,N_3900);
or U4049 (N_4049,N_3885,N_838);
xor U4050 (N_4050,In_175,N_3538);
or U4051 (N_4051,N_3350,N_3733);
nand U4052 (N_4052,N_3624,N_2169);
xnor U4053 (N_4053,N_3793,N_3712);
xor U4054 (N_4054,N_3891,N_3551);
nand U4055 (N_4055,N_3711,N_3874);
and U4056 (N_4056,N_3801,N_3367);
and U4057 (N_4057,In_665,N_3497);
and U4058 (N_4058,N_498,N_2866);
or U4059 (N_4059,N_258,N_3427);
xnor U4060 (N_4060,N_2098,N_2493);
or U4061 (N_4061,N_3882,N_3445);
or U4062 (N_4062,N_2554,N_3464);
nor U4063 (N_4063,N_2729,N_3372);
or U4064 (N_4064,N_2112,N_3990);
and U4065 (N_4065,N_3559,N_3552);
nand U4066 (N_4066,In_3017,N_289);
or U4067 (N_4067,N_3931,N_3783);
nand U4068 (N_4068,In_158,N_3463);
nor U4069 (N_4069,In_3134,N_3781);
nand U4070 (N_4070,N_2184,In_795);
nor U4071 (N_4071,In_2426,N_1048);
nand U4072 (N_4072,N_2553,N_3767);
nand U4073 (N_4073,N_2540,N_3451);
or U4074 (N_4074,N_1415,N_2087);
nor U4075 (N_4075,N_903,N_3335);
xnor U4076 (N_4076,N_3964,N_578);
xor U4077 (N_4077,N_3545,In_3735);
nand U4078 (N_4078,N_151,In_3418);
xnor U4079 (N_4079,N_3017,N_2033);
nand U4080 (N_4080,N_3666,N_3078);
or U4081 (N_4081,N_3706,In_4614);
or U4082 (N_4082,N_1502,N_3823);
nand U4083 (N_4083,N_3485,N_2886);
nand U4084 (N_4084,N_2526,N_3975);
xor U4085 (N_4085,N_3283,N_3743);
or U4086 (N_4086,N_3541,N_1474);
nand U4087 (N_4087,In_2246,N_3897);
or U4088 (N_4088,N_3299,N_3198);
or U4089 (N_4089,N_3698,In_3152);
nor U4090 (N_4090,N_2614,N_3940);
nor U4091 (N_4091,N_3550,N_1356);
nand U4092 (N_4092,N_3105,N_3631);
or U4093 (N_4093,N_3589,N_3924);
xor U4094 (N_4094,N_3645,In_1829);
nand U4095 (N_4095,In_2311,N_2915);
nor U4096 (N_4096,N_3864,N_2944);
nand U4097 (N_4097,N_2873,N_3517);
xor U4098 (N_4098,N_3848,N_3700);
nand U4099 (N_4099,N_3815,N_3553);
nand U4100 (N_4100,N_3450,N_3860);
and U4101 (N_4101,N_1487,N_2057);
nor U4102 (N_4102,N_2875,N_3616);
or U4103 (N_4103,N_3945,N_3905);
nor U4104 (N_4104,N_3511,N_3521);
nand U4105 (N_4105,N_3386,N_2);
and U4106 (N_4106,N_3556,In_4965);
and U4107 (N_4107,N_1826,In_2080);
nand U4108 (N_4108,N_3950,N_3322);
nor U4109 (N_4109,N_3862,N_3870);
and U4110 (N_4110,N_2924,N_3617);
xor U4111 (N_4111,N_3683,In_957);
or U4112 (N_4112,N_757,N_3944);
or U4113 (N_4113,N_3619,N_3407);
nor U4114 (N_4114,N_1925,N_3816);
or U4115 (N_4115,N_3825,N_3782);
or U4116 (N_4116,N_3889,N_3759);
and U4117 (N_4117,N_2964,N_3561);
and U4118 (N_4118,N_3855,N_3342);
xor U4119 (N_4119,N_3068,N_3880);
nor U4120 (N_4120,N_3371,N_3548);
nor U4121 (N_4121,N_3920,N_3887);
nand U4122 (N_4122,N_2271,In_3013);
nor U4123 (N_4123,In_4098,N_2074);
or U4124 (N_4124,N_3267,N_3308);
and U4125 (N_4125,N_3488,N_3004);
and U4126 (N_4126,N_3936,N_2907);
xnor U4127 (N_4127,N_3225,N_3325);
nor U4128 (N_4128,N_3976,N_3565);
xnor U4129 (N_4129,In_1940,N_2060);
nor U4130 (N_4130,N_1073,N_3903);
xor U4131 (N_4131,In_4677,N_3546);
and U4132 (N_4132,N_2800,N_3750);
nor U4133 (N_4133,N_2616,N_3820);
or U4134 (N_4134,N_1176,N_3594);
nand U4135 (N_4135,N_54,N_285);
or U4136 (N_4136,In_84,N_2796);
nand U4137 (N_4137,N_761,N_1036);
xnor U4138 (N_4138,N_2409,In_3463);
xnor U4139 (N_4139,N_3969,N_3046);
or U4140 (N_4140,N_3183,N_3895);
or U4141 (N_4141,N_3738,N_3907);
nor U4142 (N_4142,N_2765,In_443);
xnor U4143 (N_4143,N_3114,N_3254);
nor U4144 (N_4144,N_3525,N_3006);
or U4145 (N_4145,N_3655,N_3982);
nor U4146 (N_4146,N_3446,N_3292);
nand U4147 (N_4147,In_4405,N_2753);
nor U4148 (N_4148,N_2588,N_3822);
xor U4149 (N_4149,N_3909,N_3543);
nand U4150 (N_4150,N_3840,N_3932);
xor U4151 (N_4151,N_2424,In_348);
xor U4152 (N_4152,N_3462,N_3346);
nand U4153 (N_4153,N_3784,N_3647);
nor U4154 (N_4154,N_3851,N_69);
xnor U4155 (N_4155,N_3035,In_4);
nor U4156 (N_4156,N_3402,N_396);
xnor U4157 (N_4157,N_3364,N_3722);
xor U4158 (N_4158,In_1470,N_3859);
nor U4159 (N_4159,N_1941,N_3251);
xor U4160 (N_4160,N_2488,N_3514);
or U4161 (N_4161,N_2822,N_3495);
xnor U4162 (N_4162,N_3967,In_4747);
nor U4163 (N_4163,N_2500,N_1587);
xor U4164 (N_4164,In_1156,N_1986);
nand U4165 (N_4165,N_3971,N_3998);
xor U4166 (N_4166,N_3381,N_3955);
nand U4167 (N_4167,In_3271,N_3416);
nand U4168 (N_4168,N_3709,N_193);
and U4169 (N_4169,N_3403,N_798);
and U4170 (N_4170,N_3917,N_3953);
and U4171 (N_4171,N_574,In_2689);
nand U4172 (N_4172,N_2297,N_2762);
xor U4173 (N_4173,In_4815,N_1317);
or U4174 (N_4174,N_1411,N_2788);
xnor U4175 (N_4175,N_3604,N_3896);
or U4176 (N_4176,N_3824,N_3915);
and U4177 (N_4177,N_3753,N_3850);
nor U4178 (N_4178,N_3158,N_3758);
xor U4179 (N_4179,N_3404,In_4012);
and U4180 (N_4180,N_3209,N_2601);
nand U4181 (N_4181,In_1200,In_3039);
xnor U4182 (N_4182,N_3690,N_3708);
and U4183 (N_4183,In_2783,N_3865);
nand U4184 (N_4184,N_3831,In_2066);
xnor U4185 (N_4185,N_3811,N_2525);
nor U4186 (N_4186,N_3856,N_3578);
nand U4187 (N_4187,N_3121,N_2928);
nor U4188 (N_4188,In_1158,N_3913);
nor U4189 (N_4189,N_3660,N_3668);
nand U4190 (N_4190,N_3876,N_2932);
xnor U4191 (N_4191,N_1499,N_3977);
xor U4192 (N_4192,N_3055,In_1191);
or U4193 (N_4193,N_3318,N_3575);
and U4194 (N_4194,N_3113,N_2713);
nand U4195 (N_4195,N_3282,N_2863);
xor U4196 (N_4196,N_3972,N_3992);
and U4197 (N_4197,N_3703,N_3077);
or U4198 (N_4198,N_1298,N_3918);
xor U4199 (N_4199,N_3331,N_1496);
and U4200 (N_4200,In_3617,N_2156);
nor U4201 (N_4201,N_3636,N_3761);
nand U4202 (N_4202,N_725,N_3054);
xor U4203 (N_4203,N_3805,N_3803);
nor U4204 (N_4204,N_3814,N_3119);
nor U4205 (N_4205,N_3598,N_2617);
xnor U4206 (N_4206,N_3797,N_3665);
nor U4207 (N_4207,In_405,N_2577);
and U4208 (N_4208,N_2004,N_2560);
and U4209 (N_4209,In_1075,N_3032);
nor U4210 (N_4210,N_2276,N_3569);
nor U4211 (N_4211,N_1664,N_3912);
nand U4212 (N_4212,N_3615,In_4758);
xor U4213 (N_4213,N_3839,N_2089);
nand U4214 (N_4214,N_2410,N_1350);
xor U4215 (N_4215,In_26,N_2449);
and U4216 (N_4216,N_3642,N_3544);
nor U4217 (N_4217,N_3770,N_3728);
nor U4218 (N_4218,N_2265,N_3537);
xor U4219 (N_4219,In_4802,In_4444);
xor U4220 (N_4220,N_3588,N_2207);
xor U4221 (N_4221,N_401,In_1501);
nor U4222 (N_4222,In_46,In_4101);
or U4223 (N_4223,N_1040,N_3344);
and U4224 (N_4224,N_3788,In_3330);
nor U4225 (N_4225,N_3632,N_3810);
or U4226 (N_4226,N_1947,N_3664);
nor U4227 (N_4227,N_1437,N_3080);
nand U4228 (N_4228,N_3988,N_3702);
or U4229 (N_4229,In_702,N_3727);
and U4230 (N_4230,N_3799,In_1980);
nor U4231 (N_4231,In_3958,N_3147);
and U4232 (N_4232,N_3684,N_3547);
and U4233 (N_4233,N_3562,N_2771);
or U4234 (N_4234,N_777,N_3580);
nand U4235 (N_4235,N_1963,N_1245);
nand U4236 (N_4236,In_4500,N_2676);
xnor U4237 (N_4237,N_3756,N_2968);
and U4238 (N_4238,N_3951,N_3883);
xnor U4239 (N_4239,N_3637,N_3599);
xor U4240 (N_4240,N_2960,N_3288);
nand U4241 (N_4241,N_3961,N_3790);
and U4242 (N_4242,N_2148,N_3430);
nor U4243 (N_4243,N_2105,N_3370);
xnor U4244 (N_4244,N_2799,N_3291);
xor U4245 (N_4245,In_4872,N_1263);
nand U4246 (N_4246,N_3921,N_3926);
xnor U4247 (N_4247,N_3987,N_2203);
or U4248 (N_4248,N_841,In_2336);
nor U4249 (N_4249,N_3634,In_878);
xnor U4250 (N_4250,N_3539,N_3769);
or U4251 (N_4251,N_3411,N_3087);
xnor U4252 (N_4252,N_3973,N_3827);
or U4253 (N_4253,N_2611,In_4403);
nor U4254 (N_4254,N_4180,N_3960);
or U4255 (N_4255,In_2021,N_3614);
and U4256 (N_4256,N_1982,N_3369);
and U4257 (N_4257,N_4140,N_3591);
nand U4258 (N_4258,In_3693,N_3875);
or U4259 (N_4259,N_3563,N_2386);
nand U4260 (N_4260,N_4078,N_4142);
and U4261 (N_4261,N_3144,N_3414);
xor U4262 (N_4262,N_3716,N_4175);
or U4263 (N_4263,N_3938,N_3115);
or U4264 (N_4264,N_3837,N_3821);
and U4265 (N_4265,N_3786,N_4046);
xor U4266 (N_4266,N_3564,N_3572);
or U4267 (N_4267,N_3705,N_3916);
nand U4268 (N_4268,In_1365,N_3833);
xnor U4269 (N_4269,N_4146,N_3536);
or U4270 (N_4270,N_3720,N_4126);
or U4271 (N_4271,In_2325,N_3772);
nand U4272 (N_4272,N_2092,N_4194);
and U4273 (N_4273,N_4232,In_3898);
xor U4274 (N_4274,N_4242,N_4116);
xor U4275 (N_4275,N_1364,N_4056);
nand U4276 (N_4276,N_3524,N_2201);
and U4277 (N_4277,N_2330,N_4064);
xor U4278 (N_4278,N_4236,N_3577);
nor U4279 (N_4279,N_4134,In_411);
nor U4280 (N_4280,N_3405,N_2603);
nor U4281 (N_4281,N_2738,N_4205);
nand U4282 (N_4282,N_4062,In_598);
nor U4283 (N_4283,N_3795,N_3013);
or U4284 (N_4284,N_3333,In_942);
nand U4285 (N_4285,N_2829,In_290);
and U4286 (N_4286,N_1288,N_2495);
xnor U4287 (N_4287,N_4168,N_3751);
or U4288 (N_4288,N_4108,N_3686);
or U4289 (N_4289,N_3045,N_3886);
xor U4290 (N_4290,N_4107,N_3965);
xnor U4291 (N_4291,N_4186,N_1396);
nand U4292 (N_4292,N_2833,N_4244);
or U4293 (N_4293,N_3934,In_3903);
xnor U4294 (N_4294,N_3762,N_4189);
xor U4295 (N_4295,N_4083,N_2478);
nor U4296 (N_4296,N_4123,N_3731);
nand U4297 (N_4297,N_3768,N_3842);
xor U4298 (N_4298,N_4022,In_353);
nor U4299 (N_4299,N_4048,N_4105);
nand U4300 (N_4300,N_3835,N_2984);
nand U4301 (N_4301,N_4208,N_4203);
nor U4302 (N_4302,N_1789,N_3136);
nand U4303 (N_4303,N_4145,In_412);
nand U4304 (N_4304,N_4217,N_4176);
or U4305 (N_4305,N_3687,N_3748);
xor U4306 (N_4306,N_1337,N_4060);
nor U4307 (N_4307,In_2177,N_3836);
nor U4308 (N_4308,In_3499,N_4006);
and U4309 (N_4309,In_4864,N_4219);
nor U4310 (N_4310,N_3421,N_3383);
nand U4311 (N_4311,In_2202,N_3968);
nor U4312 (N_4312,In_3860,N_4003);
nand U4313 (N_4313,N_3830,N_4047);
or U4314 (N_4314,In_4933,N_2664);
xor U4315 (N_4315,N_4138,N_3163);
nor U4316 (N_4316,N_4132,N_4014);
nor U4317 (N_4317,N_4097,N_4121);
xnor U4318 (N_4318,N_4165,N_4193);
nor U4319 (N_4319,N_3586,N_4100);
nor U4320 (N_4320,N_4181,N_2872);
or U4321 (N_4321,N_3263,N_4081);
or U4322 (N_4322,N_4133,N_4069);
nor U4323 (N_4323,N_4034,N_3566);
xnor U4324 (N_4324,N_1980,N_4124);
xor U4325 (N_4325,N_3509,N_1523);
or U4326 (N_4326,N_4122,N_3957);
nor U4327 (N_4327,N_3774,N_2026);
or U4328 (N_4328,N_3285,N_4169);
and U4329 (N_4329,N_3943,N_4136);
nor U4330 (N_4330,N_4188,N_576);
nor U4331 (N_4331,N_4197,N_784);
or U4332 (N_4332,In_4695,N_1805);
nor U4333 (N_4333,N_2288,N_3018);
and U4334 (N_4334,In_2140,N_1563);
nor U4335 (N_4335,N_3775,N_3780);
nor U4336 (N_4336,N_3221,N_1478);
and U4337 (N_4337,N_3304,N_3277);
or U4338 (N_4338,N_3089,N_3677);
xor U4339 (N_4339,N_3675,N_3997);
nand U4340 (N_4340,N_3633,N_4177);
nand U4341 (N_4341,N_4087,In_2429);
xnor U4342 (N_4342,N_3287,N_3380);
and U4343 (N_4343,N_2468,In_142);
nand U4344 (N_4344,N_3694,N_3568);
xnor U4345 (N_4345,N_3730,N_3692);
nor U4346 (N_4346,N_3879,N_4141);
or U4347 (N_4347,N_3173,N_2741);
nand U4348 (N_4348,In_3978,N_4089);
or U4349 (N_4349,N_2260,N_3958);
nor U4350 (N_4350,N_3832,N_4247);
or U4351 (N_4351,N_3638,N_3872);
xnor U4352 (N_4352,N_4218,N_3755);
nand U4353 (N_4353,N_4118,N_505);
nor U4354 (N_4354,N_3075,N_4007);
nand U4355 (N_4355,N_4237,N_3986);
nor U4356 (N_4356,N_3084,N_3399);
xor U4357 (N_4357,N_3919,N_3623);
xnor U4358 (N_4358,N_2382,N_3763);
xnor U4359 (N_4359,N_3555,N_4111);
and U4360 (N_4360,N_3904,In_108);
nand U4361 (N_4361,In_2183,N_3659);
xor U4362 (N_4362,N_3558,N_1754);
or U4363 (N_4363,N_3266,In_1608);
and U4364 (N_4364,In_3189,In_3411);
nor U4365 (N_4365,N_3206,In_1487);
and U4366 (N_4366,N_3800,N_4054);
or U4367 (N_4367,N_4249,N_4211);
nor U4368 (N_4368,N_4095,N_4163);
nand U4369 (N_4369,N_4091,In_4673);
xor U4370 (N_4370,N_3293,N_4227);
nor U4371 (N_4371,N_3935,N_3351);
and U4372 (N_4372,In_2766,N_2952);
nand U4373 (N_4373,N_3579,N_3362);
nand U4374 (N_4374,N_3721,N_2232);
nand U4375 (N_4375,N_3906,N_4055);
and U4376 (N_4376,N_4156,N_3000);
nor U4377 (N_4377,N_3995,N_4153);
nand U4378 (N_4378,N_4222,N_3468);
or U4379 (N_4379,N_4192,In_4842);
nor U4380 (N_4380,In_3480,N_4027);
and U4381 (N_4381,N_3392,N_3387);
xnor U4382 (N_4382,N_3974,N_3278);
and U4383 (N_4383,N_4042,N_4226);
nand U4384 (N_4384,N_4112,N_4171);
xor U4385 (N_4385,N_2912,N_3813);
nand U4386 (N_4386,N_3942,N_4040);
xnor U4387 (N_4387,N_4028,N_4238);
nand U4388 (N_4388,N_2669,N_3582);
and U4389 (N_4389,N_843,In_2342);
nor U4390 (N_4390,N_3120,In_4599);
and U4391 (N_4391,N_1209,N_4065);
and U4392 (N_4392,N_3672,N_2561);
nor U4393 (N_4393,N_3923,In_3612);
xnor U4394 (N_4394,N_4020,N_4031);
nand U4395 (N_4395,N_4052,N_2264);
xor U4396 (N_4396,N_3601,N_3475);
nand U4397 (N_4397,N_4102,N_1059);
and U4398 (N_4398,N_4129,N_4213);
xnor U4399 (N_4399,N_4101,N_2951);
nor U4400 (N_4400,N_4012,N_3787);
or U4401 (N_4401,N_3838,N_4094);
nor U4402 (N_4402,In_4499,N_4029);
or U4403 (N_4403,N_3927,N_4079);
nand U4404 (N_4404,N_4173,N_3258);
and U4405 (N_4405,N_3102,N_3785);
and U4406 (N_4406,N_3520,N_3754);
and U4407 (N_4407,In_613,N_4172);
and U4408 (N_4408,N_3910,N_2228);
or U4409 (N_4409,N_3397,N_4098);
and U4410 (N_4410,N_3884,N_3979);
and U4411 (N_4411,N_2368,N_3765);
and U4412 (N_4412,N_3937,N_4013);
and U4413 (N_4413,N_3438,In_1390);
or U4414 (N_4414,N_4113,N_3959);
or U4415 (N_4415,N_4160,N_3187);
nor U4416 (N_4416,N_4204,N_2534);
nor U4417 (N_4417,N_3952,N_3737);
xor U4418 (N_4418,N_3276,N_4131);
or U4419 (N_4419,N_3161,N_4009);
or U4420 (N_4420,N_3412,N_4229);
or U4421 (N_4421,N_4190,N_3290);
xnor U4422 (N_4422,N_4117,N_3175);
nor U4423 (N_4423,In_3352,N_4166);
xor U4424 (N_4424,N_3776,N_2854);
xnor U4425 (N_4425,N_3135,N_4053);
nor U4426 (N_4426,N_2215,N_2836);
xor U4427 (N_4427,N_3868,N_3841);
or U4428 (N_4428,N_4127,N_4202);
nor U4429 (N_4429,N_4191,N_4240);
nand U4430 (N_4430,N_3985,N_3248);
or U4431 (N_4431,N_4088,N_2727);
nand U4432 (N_4432,N_3653,N_3757);
or U4433 (N_4433,N_3873,N_3466);
nand U4434 (N_4434,N_3272,N_4224);
xor U4435 (N_4435,N_3507,N_394);
nor U4436 (N_4436,N_3348,N_3946);
nand U4437 (N_4437,N_3962,N_3898);
nor U4438 (N_4438,N_4025,N_4164);
nand U4439 (N_4439,N_3384,N_3789);
xnor U4440 (N_4440,N_3718,N_4207);
or U4441 (N_4441,N_4155,In_4172);
or U4442 (N_4442,N_3012,N_3954);
xor U4443 (N_4443,N_2171,N_4159);
nand U4444 (N_4444,N_4152,N_3652);
nor U4445 (N_4445,N_1069,N_3469);
or U4446 (N_4446,N_3627,In_467);
and U4447 (N_4447,N_1670,N_2935);
and U4448 (N_4448,N_4216,N_4035);
nand U4449 (N_4449,N_2939,In_578);
or U4450 (N_4450,N_4023,N_3980);
xnor U4451 (N_4451,N_3778,N_4019);
or U4452 (N_4452,N_3991,N_4024);
xor U4453 (N_4453,N_4241,N_3908);
or U4454 (N_4454,N_4147,N_2979);
xnor U4455 (N_4455,N_4004,N_3798);
or U4456 (N_4456,N_4114,N_3396);
or U4457 (N_4457,N_4075,N_3725);
nand U4458 (N_4458,In_1185,N_3001);
nand U4459 (N_4459,In_2959,N_3329);
xor U4460 (N_4460,N_3494,N_3670);
or U4461 (N_4461,N_2226,N_3050);
or U4462 (N_4462,N_3779,N_3247);
nor U4463 (N_4463,N_548,N_3379);
and U4464 (N_4464,N_3510,N_3914);
nor U4465 (N_4465,In_3055,N_3228);
nand U4466 (N_4466,In_3030,N_2645);
xor U4467 (N_4467,N_182,N_4209);
nand U4468 (N_4468,N_3773,N_4051);
nor U4469 (N_4469,N_1709,N_3256);
and U4470 (N_4470,N_3042,N_4090);
or U4471 (N_4471,N_3999,N_4073);
nand U4472 (N_4472,N_2910,N_2254);
or U4473 (N_4473,N_1931,N_4005);
xnor U4474 (N_4474,N_4032,N_2589);
nand U4475 (N_4475,N_1014,N_3458);
nand U4476 (N_4476,N_1861,N_4243);
xor U4477 (N_4477,N_4074,N_4115);
xnor U4478 (N_4478,N_3893,In_4094);
and U4479 (N_4479,N_4231,N_4154);
xor U4480 (N_4480,N_4120,N_4130);
and U4481 (N_4481,In_4715,N_3941);
or U4482 (N_4482,N_130,N_3808);
or U4483 (N_4483,N_3528,N_3424);
or U4484 (N_4484,In_4918,N_3994);
nand U4485 (N_4485,In_1607,N_4151);
and U4486 (N_4486,N_3857,N_3338);
or U4487 (N_4487,N_2680,N_3549);
or U4488 (N_4488,N_2111,In_3635);
nand U4489 (N_4489,N_4125,N_3878);
nand U4490 (N_4490,N_4162,In_641);
and U4491 (N_4491,N_3849,N_3629);
nand U4492 (N_4492,N_4210,In_3216);
nor U4493 (N_4493,N_3817,N_3560);
nor U4494 (N_4494,N_44,In_3986);
xor U4495 (N_4495,N_1501,N_1929);
nand U4496 (N_4496,N_4038,N_3218);
nand U4497 (N_4497,N_2670,N_3590);
nor U4498 (N_4498,N_3766,N_4071);
and U4499 (N_4499,N_3097,N_1453);
or U4500 (N_4500,N_3794,N_4439);
or U4501 (N_4501,N_3948,N_4393);
nand U4502 (N_4502,N_4279,N_4033);
and U4503 (N_4503,N_4449,N_4421);
and U4504 (N_4504,N_4375,N_4149);
nor U4505 (N_4505,In_3930,N_3680);
and U4506 (N_4506,N_4371,N_3174);
xnor U4507 (N_4507,N_3375,N_4016);
nand U4508 (N_4508,N_4398,N_3613);
xnor U4509 (N_4509,N_4256,N_4352);
and U4510 (N_4510,N_4150,N_4477);
nor U4511 (N_4511,N_4036,N_4092);
and U4512 (N_4512,N_4263,N_4293);
xor U4513 (N_4513,N_4220,In_910);
nor U4514 (N_4514,N_4057,N_4257);
or U4515 (N_4515,N_2095,N_4178);
nor U4516 (N_4516,N_4382,N_4471);
xnor U4517 (N_4517,N_3829,N_4255);
or U4518 (N_4518,N_4323,N_4473);
and U4519 (N_4519,N_4137,N_3557);
nor U4520 (N_4520,In_2498,N_4315);
or U4521 (N_4521,N_4428,N_3340);
or U4522 (N_4522,N_3196,N_4063);
xnor U4523 (N_4523,N_4326,N_4061);
xor U4524 (N_4524,N_4450,N_3877);
and U4525 (N_4525,N_3984,N_2586);
nand U4526 (N_4526,N_3869,In_1164);
nor U4527 (N_4527,N_4310,N_4372);
nor U4528 (N_4528,N_2110,N_4200);
nor U4529 (N_4529,N_3233,N_4438);
nand U4530 (N_4530,N_4252,In_4299);
nor U4531 (N_4531,In_48,N_4445);
or U4532 (N_4532,N_4309,N_4329);
and U4533 (N_4533,N_4459,N_3373);
or U4534 (N_4534,N_4157,N_4044);
or U4535 (N_4535,N_4360,N_3760);
and U4536 (N_4536,N_4328,In_590);
nand U4537 (N_4537,N_1077,N_4225);
and U4538 (N_4538,N_4491,N_4342);
nor U4539 (N_4539,N_3071,N_4308);
nor U4540 (N_4540,N_4453,N_4403);
and U4541 (N_4541,N_2658,N_4085);
and U4542 (N_4542,N_3180,N_4321);
nand U4543 (N_4543,N_4008,N_4206);
or U4544 (N_4544,N_4433,N_4402);
xnor U4545 (N_4545,N_1031,N_4377);
nand U4546 (N_4546,N_3930,N_4422);
xnor U4547 (N_4547,In_3963,N_2483);
nor U4548 (N_4548,N_4364,N_4376);
xnor U4549 (N_4549,N_4365,N_4233);
xor U4550 (N_4550,N_4317,N_4346);
or U4551 (N_4551,N_4454,N_4158);
nor U4552 (N_4552,N_4110,N_4119);
nand U4553 (N_4553,N_2991,N_4262);
nand U4554 (N_4554,N_3894,N_1144);
or U4555 (N_4555,N_4397,N_2831);
and U4556 (N_4556,N_4215,N_3678);
nor U4557 (N_4557,N_4254,N_4290);
xnor U4558 (N_4558,N_4099,N_4432);
nand U4559 (N_4559,N_4261,N_4399);
and U4560 (N_4560,N_4353,N_4246);
nand U4561 (N_4561,N_4482,N_4492);
or U4562 (N_4562,N_4331,N_4344);
nor U4563 (N_4563,N_1679,N_4182);
nand U4564 (N_4564,In_20,N_4026);
and U4565 (N_4565,N_4404,N_3949);
or U4566 (N_4566,N_4411,N_2868);
or U4567 (N_4567,N_4304,N_4301);
nand U4568 (N_4568,N_4458,N_4086);
nand U4569 (N_4569,N_4388,N_4351);
nand U4570 (N_4570,N_3843,N_4363);
and U4571 (N_4571,N_4370,N_3377);
xor U4572 (N_4572,N_4367,N_4278);
or U4573 (N_4573,N_4385,N_4495);
and U4574 (N_4574,N_4401,N_4059);
xor U4575 (N_4575,N_4461,N_4339);
nand U4576 (N_4576,N_4408,N_4348);
nand U4577 (N_4577,N_4460,N_4297);
xnor U4578 (N_4578,N_4068,N_4228);
xnor U4579 (N_4579,N_4302,N_3901);
nor U4580 (N_4580,N_4457,N_900);
nor U4581 (N_4581,N_4199,N_4299);
nand U4582 (N_4582,N_4467,N_4474);
nand U4583 (N_4583,N_3963,N_4369);
nand U4584 (N_4584,N_3016,N_4084);
nand U4585 (N_4585,N_4407,N_4378);
nand U4586 (N_4586,N_4425,N_4283);
and U4587 (N_4587,N_4488,N_4287);
or U4588 (N_4588,N_4041,N_4082);
nor U4589 (N_4589,N_4135,N_4010);
nor U4590 (N_4590,N_4077,N_3819);
or U4591 (N_4591,N_4324,N_4295);
xnor U4592 (N_4592,N_4322,N_4271);
or U4593 (N_4593,N_4313,N_4248);
and U4594 (N_4594,N_3729,N_3752);
or U4595 (N_4595,N_4462,N_4368);
nor U4596 (N_4596,N_3888,N_4285);
or U4597 (N_4597,N_4284,N_4330);
nor U4598 (N_4598,N_3981,N_4480);
nand U4599 (N_4599,N_3881,N_2933);
or U4600 (N_4600,N_1885,In_4451);
nand U4601 (N_4601,N_4409,N_4465);
and U4602 (N_4602,N_4230,N_4030);
nand U4603 (N_4603,N_4395,N_2857);
xor U4604 (N_4604,N_4187,N_3356);
and U4605 (N_4605,N_183,N_2557);
and U4606 (N_4606,N_4274,N_4049);
and U4607 (N_4607,N_4496,N_4250);
or U4608 (N_4608,N_4357,N_4017);
nand U4609 (N_4609,N_4350,N_4039);
nor U4610 (N_4610,In_3109,N_4174);
and U4611 (N_4611,N_4000,N_4201);
and U4612 (N_4612,N_4338,N_4405);
xnor U4613 (N_4613,N_4015,N_4291);
nor U4614 (N_4614,N_4335,N_4483);
and U4615 (N_4615,N_4334,N_4266);
xnor U4616 (N_4616,N_3155,N_4389);
and U4617 (N_4617,N_4312,N_4286);
and U4618 (N_4618,N_3695,N_3983);
nand U4619 (N_4619,N_3996,N_4002);
nor U4620 (N_4620,N_4307,N_4185);
nor U4621 (N_4621,N_3871,N_4358);
or U4622 (N_4622,N_3792,N_4469);
nand U4623 (N_4623,N_4264,N_4484);
and U4624 (N_4624,N_4198,In_4332);
xnor U4625 (N_4625,N_4143,N_4214);
or U4626 (N_4626,N_3220,N_4333);
or U4627 (N_4627,N_4493,N_3606);
nor U4628 (N_4628,N_4251,N_3058);
nand U4629 (N_4629,N_4391,N_4355);
xnor U4630 (N_4630,N_4394,N_4272);
or U4631 (N_4631,N_4167,N_3061);
or U4632 (N_4632,N_4431,N_3993);
xnor U4633 (N_4633,N_4485,In_3482);
nand U4634 (N_4634,N_4300,N_4464);
or U4635 (N_4635,N_4341,N_4337);
nand U4636 (N_4636,N_3978,N_4332);
nor U4637 (N_4637,In_2896,N_187);
and U4638 (N_4638,N_4109,N_4490);
and U4639 (N_4639,In_1818,N_4441);
and U4640 (N_4640,N_4294,N_4179);
nor U4641 (N_4641,N_4325,In_4964);
and U4642 (N_4642,N_2063,N_4340);
and U4643 (N_4643,N_4345,In_1196);
or U4644 (N_4644,N_3802,N_1466);
nand U4645 (N_4645,N_4234,N_3306);
and U4646 (N_4646,N_3587,N_4381);
xor U4647 (N_4647,N_3956,N_2881);
nor U4648 (N_4648,N_4103,N_4298);
nand U4649 (N_4649,N_4183,N_4466);
and U4650 (N_4650,N_4018,N_2355);
or U4651 (N_4651,N_4316,N_4066);
xor U4652 (N_4652,N_4489,N_4415);
xor U4653 (N_4653,N_2812,In_1594);
nor U4654 (N_4654,N_4273,N_4011);
nor U4655 (N_4655,N_4379,N_2100);
nor U4656 (N_4656,In_2417,N_4410);
nor U4657 (N_4657,N_4387,N_4067);
and U4658 (N_4658,N_4374,N_4303);
and U4659 (N_4659,N_4259,N_1100);
and U4660 (N_4660,N_4412,N_3646);
xor U4661 (N_4661,N_4481,N_4076);
or U4662 (N_4662,N_4414,N_4045);
nor U4663 (N_4663,N_3867,N_3804);
and U4664 (N_4664,N_4390,N_4311);
and U4665 (N_4665,N_4442,N_3966);
nand U4666 (N_4666,N_4281,N_4096);
nor U4667 (N_4667,N_4277,N_4343);
or U4668 (N_4668,N_4448,N_3051);
or U4669 (N_4669,N_4396,N_4080);
nor U4670 (N_4670,N_4354,N_4050);
or U4671 (N_4671,N_2447,N_3899);
nor U4672 (N_4672,N_3260,N_902);
and U4673 (N_4673,N_4161,N_4362);
or U4674 (N_4674,N_4196,N_4288);
xor U4675 (N_4675,N_4470,N_4478);
xor U4676 (N_4676,N_4318,N_4058);
nor U4677 (N_4677,N_3806,N_3828);
nor U4678 (N_4678,N_2982,N_4336);
and U4679 (N_4679,N_3902,N_4386);
xor U4680 (N_4680,N_3929,N_4072);
and U4681 (N_4681,N_4327,N_4319);
or U4682 (N_4682,N_4384,In_1052);
or U4683 (N_4683,N_4392,N_2659);
and U4684 (N_4684,N_4447,N_4400);
or U4685 (N_4685,N_4292,N_3347);
or U4686 (N_4686,N_4093,N_3853);
nor U4687 (N_4687,N_4144,N_4452);
xor U4688 (N_4688,N_2349,N_4417);
nand U4689 (N_4689,N_4184,N_4276);
or U4690 (N_4690,N_4444,N_2955);
xor U4691 (N_4691,N_4486,N_2578);
nor U4692 (N_4692,N_1924,N_4413);
or U4693 (N_4693,N_4424,N_4245);
and U4694 (N_4694,N_4423,N_4347);
nor U4695 (N_4695,N_4487,N_4427);
or U4696 (N_4696,N_4406,N_4258);
nand U4697 (N_4697,N_2269,N_4436);
nor U4698 (N_4698,N_2474,N_4359);
or U4699 (N_4699,N_2747,N_4440);
nor U4700 (N_4700,N_4416,N_3791);
and U4701 (N_4701,N_4435,In_2837);
and U4702 (N_4702,In_4525,N_4221);
xnor U4703 (N_4703,N_4475,N_4260);
and U4704 (N_4704,In_3476,N_4148);
nor U4705 (N_4705,N_4499,N_3540);
and U4706 (N_4706,N_4468,N_4306);
xor U4707 (N_4707,N_4429,In_3148);
and U4708 (N_4708,N_350,N_4268);
and U4709 (N_4709,N_4195,N_3846);
nand U4710 (N_4710,N_3423,N_4305);
nor U4711 (N_4711,N_4282,N_3518);
and U4712 (N_4712,N_4269,N_4443);
xor U4713 (N_4713,N_4380,N_4070);
nand U4714 (N_4714,N_4043,N_4128);
and U4715 (N_4715,N_4001,N_4455);
nor U4716 (N_4716,N_4275,N_596);
nand U4717 (N_4717,N_4498,N_1334);
nor U4718 (N_4718,N_4037,N_4280);
nor U4719 (N_4719,N_4021,N_2085);
or U4720 (N_4720,In_4821,N_4320);
and U4721 (N_4721,N_3866,N_4426);
nand U4722 (N_4722,N_351,N_4212);
nand U4723 (N_4723,In_3937,In_452);
xnor U4724 (N_4724,N_4451,N_1019);
xnor U4725 (N_4725,N_4419,N_3764);
and U4726 (N_4726,N_4267,N_4497);
xnor U4727 (N_4727,N_4356,N_4446);
or U4728 (N_4728,N_4418,N_3890);
or U4729 (N_4729,N_4296,N_86);
nand U4730 (N_4730,N_3834,N_4361);
xor U4731 (N_4731,N_4239,N_4476);
nor U4732 (N_4732,N_4265,N_4472);
and U4733 (N_4733,N_3534,In_4773);
xnor U4734 (N_4734,N_4479,N_4270);
and U4735 (N_4735,N_3393,N_4456);
nor U4736 (N_4736,N_4104,N_2054);
nor U4737 (N_4737,N_3739,N_4437);
xnor U4738 (N_4738,N_4373,In_794);
xor U4739 (N_4739,N_4139,N_3685);
and U4740 (N_4740,N_4383,N_4106);
nor U4741 (N_4741,N_4494,N_3847);
and U4742 (N_4742,N_4430,N_4434);
nor U4743 (N_4743,In_1511,N_2556);
and U4744 (N_4744,N_4289,N_3644);
xnor U4745 (N_4745,N_4349,N_4235);
xor U4746 (N_4746,N_3296,N_4463);
or U4747 (N_4747,N_4223,N_4170);
or U4748 (N_4748,N_4420,N_4253);
and U4749 (N_4749,N_4366,N_4314);
xnor U4750 (N_4750,N_4549,N_4623);
and U4751 (N_4751,N_4720,N_4696);
and U4752 (N_4752,N_4532,N_4569);
xor U4753 (N_4753,N_4505,N_4728);
and U4754 (N_4754,N_4706,N_4625);
xnor U4755 (N_4755,N_4530,N_4718);
xor U4756 (N_4756,N_4660,N_4556);
or U4757 (N_4757,N_4554,N_4630);
xor U4758 (N_4758,N_4681,N_4680);
nor U4759 (N_4759,N_4580,N_4540);
and U4760 (N_4760,N_4703,N_4624);
xnor U4761 (N_4761,N_4677,N_4541);
nor U4762 (N_4762,N_4509,N_4545);
xnor U4763 (N_4763,N_4678,N_4654);
and U4764 (N_4764,N_4508,N_4652);
nor U4765 (N_4765,N_4745,N_4515);
and U4766 (N_4766,N_4558,N_4514);
nand U4767 (N_4767,N_4691,N_4721);
nor U4768 (N_4768,N_4638,N_4744);
nor U4769 (N_4769,N_4562,N_4560);
and U4770 (N_4770,N_4565,N_4719);
or U4771 (N_4771,N_4741,N_4581);
nor U4772 (N_4772,N_4666,N_4570);
nand U4773 (N_4773,N_4566,N_4689);
nor U4774 (N_4774,N_4688,N_4636);
or U4775 (N_4775,N_4544,N_4674);
and U4776 (N_4776,N_4538,N_4606);
and U4777 (N_4777,N_4628,N_4687);
or U4778 (N_4778,N_4704,N_4643);
xnor U4779 (N_4779,N_4551,N_4573);
nand U4780 (N_4780,N_4631,N_4608);
xnor U4781 (N_4781,N_4507,N_4726);
xor U4782 (N_4782,N_4559,N_4679);
nand U4783 (N_4783,N_4520,N_4603);
nand U4784 (N_4784,N_4592,N_4697);
xnor U4785 (N_4785,N_4513,N_4649);
nor U4786 (N_4786,N_4723,N_4621);
or U4787 (N_4787,N_4646,N_4604);
and U4788 (N_4788,N_4732,N_4567);
xor U4789 (N_4789,N_4640,N_4734);
nand U4790 (N_4790,N_4733,N_4589);
or U4791 (N_4791,N_4516,N_4637);
or U4792 (N_4792,N_4684,N_4525);
and U4793 (N_4793,N_4627,N_4710);
xnor U4794 (N_4794,N_4598,N_4673);
nor U4795 (N_4795,N_4634,N_4594);
and U4796 (N_4796,N_4612,N_4664);
nand U4797 (N_4797,N_4534,N_4500);
and U4798 (N_4798,N_4511,N_4523);
nand U4799 (N_4799,N_4522,N_4561);
nor U4800 (N_4800,N_4690,N_4685);
nand U4801 (N_4801,N_4577,N_4583);
xnor U4802 (N_4802,N_4671,N_4709);
nor U4803 (N_4803,N_4686,N_4512);
nor U4804 (N_4804,N_4542,N_4553);
and U4805 (N_4805,N_4714,N_4731);
and U4806 (N_4806,N_4742,N_4582);
nand U4807 (N_4807,N_4632,N_4571);
or U4808 (N_4808,N_4555,N_4518);
nand U4809 (N_4809,N_4669,N_4614);
and U4810 (N_4810,N_4699,N_4656);
nand U4811 (N_4811,N_4503,N_4730);
nor U4812 (N_4812,N_4552,N_4617);
or U4813 (N_4813,N_4543,N_4692);
and U4814 (N_4814,N_4700,N_4529);
or U4815 (N_4815,N_4644,N_4504);
and U4816 (N_4816,N_4675,N_4657);
nand U4817 (N_4817,N_4536,N_4575);
or U4818 (N_4818,N_4531,N_4572);
or U4819 (N_4819,N_4672,N_4695);
nor U4820 (N_4820,N_4626,N_4749);
nand U4821 (N_4821,N_4563,N_4712);
and U4822 (N_4822,N_4601,N_4587);
nor U4823 (N_4823,N_4639,N_4622);
and U4824 (N_4824,N_4715,N_4641);
or U4825 (N_4825,N_4659,N_4633);
xnor U4826 (N_4826,N_4737,N_4588);
nor U4827 (N_4827,N_4683,N_4629);
and U4828 (N_4828,N_4611,N_4597);
nor U4829 (N_4829,N_4574,N_4738);
nor U4830 (N_4830,N_4506,N_4519);
nand U4831 (N_4831,N_4528,N_4548);
xnor U4832 (N_4832,N_4698,N_4510);
nand U4833 (N_4833,N_4605,N_4722);
or U4834 (N_4834,N_4568,N_4618);
or U4835 (N_4835,N_4591,N_4593);
or U4836 (N_4836,N_4526,N_4662);
xnor U4837 (N_4837,N_4501,N_4610);
nand U4838 (N_4838,N_4645,N_4655);
nor U4839 (N_4839,N_4584,N_4596);
nand U4840 (N_4840,N_4602,N_4642);
and U4841 (N_4841,N_4727,N_4539);
xor U4842 (N_4842,N_4502,N_4707);
nor U4843 (N_4843,N_4708,N_4701);
nor U4844 (N_4844,N_4740,N_4550);
or U4845 (N_4845,N_4746,N_4537);
xnor U4846 (N_4846,N_4702,N_4579);
nor U4847 (N_4847,N_4600,N_4739);
xnor U4848 (N_4848,N_4711,N_4653);
nor U4849 (N_4849,N_4748,N_4670);
xor U4850 (N_4850,N_4533,N_4724);
and U4851 (N_4851,N_4713,N_4517);
nand U4852 (N_4852,N_4524,N_4599);
and U4853 (N_4853,N_4667,N_4651);
xnor U4854 (N_4854,N_4736,N_4694);
nor U4855 (N_4855,N_4682,N_4527);
xor U4856 (N_4856,N_4620,N_4743);
and U4857 (N_4857,N_4546,N_4578);
nand U4858 (N_4858,N_4747,N_4564);
xor U4859 (N_4859,N_4693,N_4650);
nor U4860 (N_4860,N_4619,N_4735);
and U4861 (N_4861,N_4729,N_4586);
and U4862 (N_4862,N_4717,N_4705);
nor U4863 (N_4863,N_4663,N_4716);
or U4864 (N_4864,N_4607,N_4665);
nor U4865 (N_4865,N_4521,N_4613);
xnor U4866 (N_4866,N_4635,N_4647);
and U4867 (N_4867,N_4725,N_4615);
or U4868 (N_4868,N_4576,N_4535);
nor U4869 (N_4869,N_4585,N_4668);
nor U4870 (N_4870,N_4557,N_4616);
nor U4871 (N_4871,N_4609,N_4547);
and U4872 (N_4872,N_4648,N_4658);
nand U4873 (N_4873,N_4676,N_4590);
or U4874 (N_4874,N_4661,N_4595);
or U4875 (N_4875,N_4564,N_4578);
and U4876 (N_4876,N_4556,N_4589);
nor U4877 (N_4877,N_4681,N_4590);
xor U4878 (N_4878,N_4513,N_4528);
and U4879 (N_4879,N_4682,N_4586);
nor U4880 (N_4880,N_4705,N_4546);
nand U4881 (N_4881,N_4726,N_4738);
and U4882 (N_4882,N_4685,N_4637);
nand U4883 (N_4883,N_4749,N_4734);
nor U4884 (N_4884,N_4735,N_4647);
or U4885 (N_4885,N_4723,N_4630);
nand U4886 (N_4886,N_4648,N_4668);
nor U4887 (N_4887,N_4675,N_4525);
nor U4888 (N_4888,N_4584,N_4739);
nand U4889 (N_4889,N_4737,N_4695);
or U4890 (N_4890,N_4620,N_4510);
and U4891 (N_4891,N_4540,N_4553);
nor U4892 (N_4892,N_4616,N_4642);
or U4893 (N_4893,N_4716,N_4705);
or U4894 (N_4894,N_4649,N_4536);
nand U4895 (N_4895,N_4655,N_4505);
xnor U4896 (N_4896,N_4583,N_4697);
and U4897 (N_4897,N_4715,N_4541);
nor U4898 (N_4898,N_4505,N_4711);
and U4899 (N_4899,N_4578,N_4722);
nand U4900 (N_4900,N_4595,N_4722);
and U4901 (N_4901,N_4553,N_4603);
nor U4902 (N_4902,N_4614,N_4742);
nand U4903 (N_4903,N_4565,N_4639);
nand U4904 (N_4904,N_4729,N_4662);
nor U4905 (N_4905,N_4632,N_4588);
and U4906 (N_4906,N_4672,N_4668);
nand U4907 (N_4907,N_4539,N_4506);
nor U4908 (N_4908,N_4743,N_4520);
nand U4909 (N_4909,N_4738,N_4677);
or U4910 (N_4910,N_4737,N_4698);
xnor U4911 (N_4911,N_4634,N_4656);
or U4912 (N_4912,N_4589,N_4668);
xnor U4913 (N_4913,N_4738,N_4687);
nand U4914 (N_4914,N_4626,N_4660);
xor U4915 (N_4915,N_4516,N_4721);
nand U4916 (N_4916,N_4680,N_4628);
or U4917 (N_4917,N_4582,N_4661);
nor U4918 (N_4918,N_4516,N_4661);
nor U4919 (N_4919,N_4745,N_4720);
or U4920 (N_4920,N_4667,N_4650);
or U4921 (N_4921,N_4661,N_4736);
xor U4922 (N_4922,N_4532,N_4739);
xor U4923 (N_4923,N_4574,N_4700);
xor U4924 (N_4924,N_4603,N_4544);
or U4925 (N_4925,N_4646,N_4513);
and U4926 (N_4926,N_4559,N_4608);
nor U4927 (N_4927,N_4593,N_4746);
nand U4928 (N_4928,N_4639,N_4641);
nand U4929 (N_4929,N_4743,N_4713);
or U4930 (N_4930,N_4578,N_4695);
xor U4931 (N_4931,N_4524,N_4613);
xnor U4932 (N_4932,N_4540,N_4562);
nand U4933 (N_4933,N_4711,N_4557);
nor U4934 (N_4934,N_4594,N_4604);
or U4935 (N_4935,N_4549,N_4725);
nor U4936 (N_4936,N_4651,N_4731);
and U4937 (N_4937,N_4575,N_4504);
and U4938 (N_4938,N_4641,N_4642);
nand U4939 (N_4939,N_4557,N_4713);
xnor U4940 (N_4940,N_4534,N_4507);
nor U4941 (N_4941,N_4595,N_4558);
nand U4942 (N_4942,N_4693,N_4709);
or U4943 (N_4943,N_4653,N_4612);
xor U4944 (N_4944,N_4564,N_4733);
nor U4945 (N_4945,N_4660,N_4643);
nand U4946 (N_4946,N_4565,N_4541);
nand U4947 (N_4947,N_4695,N_4736);
xnor U4948 (N_4948,N_4517,N_4643);
xnor U4949 (N_4949,N_4602,N_4545);
xnor U4950 (N_4950,N_4618,N_4626);
and U4951 (N_4951,N_4645,N_4642);
xor U4952 (N_4952,N_4679,N_4702);
nor U4953 (N_4953,N_4502,N_4511);
and U4954 (N_4954,N_4535,N_4630);
xnor U4955 (N_4955,N_4657,N_4649);
nor U4956 (N_4956,N_4584,N_4741);
nor U4957 (N_4957,N_4637,N_4668);
nor U4958 (N_4958,N_4606,N_4741);
nand U4959 (N_4959,N_4536,N_4721);
and U4960 (N_4960,N_4711,N_4673);
or U4961 (N_4961,N_4684,N_4601);
xnor U4962 (N_4962,N_4531,N_4718);
nand U4963 (N_4963,N_4514,N_4629);
or U4964 (N_4964,N_4553,N_4616);
and U4965 (N_4965,N_4564,N_4611);
or U4966 (N_4966,N_4631,N_4656);
and U4967 (N_4967,N_4679,N_4570);
nor U4968 (N_4968,N_4532,N_4626);
nand U4969 (N_4969,N_4715,N_4612);
nand U4970 (N_4970,N_4504,N_4551);
xor U4971 (N_4971,N_4742,N_4546);
nand U4972 (N_4972,N_4661,N_4502);
nor U4973 (N_4973,N_4703,N_4699);
or U4974 (N_4974,N_4602,N_4567);
or U4975 (N_4975,N_4636,N_4657);
xnor U4976 (N_4976,N_4542,N_4574);
xnor U4977 (N_4977,N_4700,N_4565);
or U4978 (N_4978,N_4654,N_4516);
or U4979 (N_4979,N_4731,N_4544);
nand U4980 (N_4980,N_4500,N_4552);
or U4981 (N_4981,N_4652,N_4557);
and U4982 (N_4982,N_4576,N_4649);
nand U4983 (N_4983,N_4524,N_4614);
xor U4984 (N_4984,N_4521,N_4731);
and U4985 (N_4985,N_4642,N_4620);
xor U4986 (N_4986,N_4644,N_4683);
nor U4987 (N_4987,N_4716,N_4725);
nor U4988 (N_4988,N_4529,N_4561);
nand U4989 (N_4989,N_4748,N_4713);
and U4990 (N_4990,N_4582,N_4668);
or U4991 (N_4991,N_4667,N_4689);
nor U4992 (N_4992,N_4721,N_4529);
nand U4993 (N_4993,N_4538,N_4580);
nor U4994 (N_4994,N_4738,N_4504);
or U4995 (N_4995,N_4519,N_4679);
nand U4996 (N_4996,N_4748,N_4693);
xor U4997 (N_4997,N_4544,N_4626);
nor U4998 (N_4998,N_4623,N_4727);
and U4999 (N_4999,N_4698,N_4597);
and U5000 (N_5000,N_4831,N_4979);
nor U5001 (N_5001,N_4996,N_4991);
xnor U5002 (N_5002,N_4786,N_4788);
nor U5003 (N_5003,N_4775,N_4935);
nor U5004 (N_5004,N_4817,N_4792);
xor U5005 (N_5005,N_4924,N_4778);
and U5006 (N_5006,N_4829,N_4989);
nor U5007 (N_5007,N_4978,N_4830);
nand U5008 (N_5008,N_4772,N_4847);
or U5009 (N_5009,N_4961,N_4988);
xor U5010 (N_5010,N_4942,N_4796);
nor U5011 (N_5011,N_4931,N_4807);
or U5012 (N_5012,N_4771,N_4939);
nand U5013 (N_5013,N_4761,N_4815);
nand U5014 (N_5014,N_4809,N_4816);
nor U5015 (N_5015,N_4838,N_4958);
nand U5016 (N_5016,N_4921,N_4836);
or U5017 (N_5017,N_4770,N_4928);
nor U5018 (N_5018,N_4883,N_4755);
xnor U5019 (N_5019,N_4977,N_4751);
nor U5020 (N_5020,N_4832,N_4812);
or U5021 (N_5021,N_4981,N_4957);
nand U5022 (N_5022,N_4824,N_4923);
nand U5023 (N_5023,N_4850,N_4990);
nor U5024 (N_5024,N_4776,N_4825);
or U5025 (N_5025,N_4798,N_4851);
nand U5026 (N_5026,N_4801,N_4911);
nor U5027 (N_5027,N_4888,N_4965);
xor U5028 (N_5028,N_4803,N_4878);
nand U5029 (N_5029,N_4834,N_4853);
and U5030 (N_5030,N_4891,N_4861);
nor U5031 (N_5031,N_4932,N_4948);
nor U5032 (N_5032,N_4835,N_4925);
or U5033 (N_5033,N_4997,N_4890);
nor U5034 (N_5034,N_4802,N_4955);
nand U5035 (N_5035,N_4768,N_4926);
or U5036 (N_5036,N_4910,N_4777);
and U5037 (N_5037,N_4762,N_4944);
nor U5038 (N_5038,N_4940,N_4870);
nor U5039 (N_5039,N_4758,N_4767);
or U5040 (N_5040,N_4892,N_4887);
or U5041 (N_5041,N_4992,N_4863);
nand U5042 (N_5042,N_4860,N_4856);
xor U5043 (N_5043,N_4793,N_4773);
or U5044 (N_5044,N_4949,N_4908);
xnor U5045 (N_5045,N_4962,N_4821);
or U5046 (N_5046,N_4766,N_4753);
or U5047 (N_5047,N_4894,N_4947);
and U5048 (N_5048,N_4909,N_4881);
nor U5049 (N_5049,N_4983,N_4993);
or U5050 (N_5050,N_4904,N_4898);
nand U5051 (N_5051,N_4889,N_4967);
nor U5052 (N_5052,N_4849,N_4859);
xor U5053 (N_5053,N_4897,N_4896);
xnor U5054 (N_5054,N_4846,N_4929);
and U5055 (N_5055,N_4938,N_4885);
nor U5056 (N_5056,N_4884,N_4917);
nor U5057 (N_5057,N_4839,N_4765);
nand U5058 (N_5058,N_4998,N_4906);
xor U5059 (N_5059,N_4805,N_4854);
and U5060 (N_5060,N_4913,N_4886);
nor U5061 (N_5061,N_4903,N_4780);
nor U5062 (N_5062,N_4862,N_4987);
xor U5063 (N_5063,N_4877,N_4995);
or U5064 (N_5064,N_4876,N_4901);
and U5065 (N_5065,N_4789,N_4785);
or U5066 (N_5066,N_4964,N_4914);
xnor U5067 (N_5067,N_4818,N_4782);
nand U5068 (N_5068,N_4959,N_4794);
nand U5069 (N_5069,N_4869,N_4804);
or U5070 (N_5070,N_4943,N_4764);
and U5071 (N_5071,N_4919,N_4760);
nor U5072 (N_5072,N_4757,N_4956);
or U5073 (N_5073,N_4968,N_4855);
xnor U5074 (N_5074,N_4810,N_4972);
and U5075 (N_5075,N_4826,N_4774);
nor U5076 (N_5076,N_4907,N_4865);
xnor U5077 (N_5077,N_4837,N_4980);
or U5078 (N_5078,N_4873,N_4867);
nor U5079 (N_5079,N_4999,N_4945);
xor U5080 (N_5080,N_4848,N_4966);
xnor U5081 (N_5081,N_4974,N_4827);
nand U5082 (N_5082,N_4916,N_4946);
nand U5083 (N_5083,N_4769,N_4822);
and U5084 (N_5084,N_4905,N_4795);
xor U5085 (N_5085,N_4941,N_4797);
nor U5086 (N_5086,N_4790,N_4902);
xnor U5087 (N_5087,N_4882,N_4915);
or U5088 (N_5088,N_4893,N_4927);
and U5089 (N_5089,N_4973,N_4871);
nor U5090 (N_5090,N_4880,N_4844);
or U5091 (N_5091,N_4784,N_4920);
xor U5092 (N_5092,N_4813,N_4823);
and U5093 (N_5093,N_4976,N_4763);
or U5094 (N_5094,N_4982,N_4950);
nand U5095 (N_5095,N_4828,N_4934);
and U5096 (N_5096,N_4971,N_4937);
or U5097 (N_5097,N_4899,N_4833);
nor U5098 (N_5098,N_4918,N_4841);
and U5099 (N_5099,N_4874,N_4872);
and U5100 (N_5100,N_4864,N_4933);
nor U5101 (N_5101,N_4857,N_4781);
nand U5102 (N_5102,N_4756,N_4994);
and U5103 (N_5103,N_4858,N_4754);
nor U5104 (N_5104,N_4752,N_4960);
nor U5105 (N_5105,N_4868,N_4820);
xor U5106 (N_5106,N_4952,N_4875);
or U5107 (N_5107,N_4936,N_4759);
nor U5108 (N_5108,N_4791,N_4879);
nand U5109 (N_5109,N_4814,N_4750);
nor U5110 (N_5110,N_4895,N_4845);
nor U5111 (N_5111,N_4951,N_4799);
nand U5112 (N_5112,N_4985,N_4954);
nor U5113 (N_5113,N_4806,N_4840);
and U5114 (N_5114,N_4808,N_4866);
or U5115 (N_5115,N_4843,N_4842);
and U5116 (N_5116,N_4970,N_4975);
and U5117 (N_5117,N_4930,N_4912);
nor U5118 (N_5118,N_4900,N_4783);
xnor U5119 (N_5119,N_4779,N_4969);
nor U5120 (N_5120,N_4963,N_4800);
and U5121 (N_5121,N_4787,N_4953);
xor U5122 (N_5122,N_4811,N_4986);
nand U5123 (N_5123,N_4922,N_4819);
or U5124 (N_5124,N_4852,N_4984);
or U5125 (N_5125,N_4764,N_4839);
or U5126 (N_5126,N_4990,N_4943);
and U5127 (N_5127,N_4925,N_4840);
and U5128 (N_5128,N_4890,N_4986);
nor U5129 (N_5129,N_4893,N_4766);
or U5130 (N_5130,N_4858,N_4977);
or U5131 (N_5131,N_4840,N_4919);
and U5132 (N_5132,N_4777,N_4947);
nor U5133 (N_5133,N_4963,N_4937);
nand U5134 (N_5134,N_4764,N_4903);
xnor U5135 (N_5135,N_4755,N_4864);
and U5136 (N_5136,N_4851,N_4761);
nand U5137 (N_5137,N_4895,N_4989);
nand U5138 (N_5138,N_4804,N_4917);
or U5139 (N_5139,N_4915,N_4902);
nand U5140 (N_5140,N_4776,N_4866);
nor U5141 (N_5141,N_4987,N_4947);
nor U5142 (N_5142,N_4818,N_4792);
nand U5143 (N_5143,N_4788,N_4877);
nand U5144 (N_5144,N_4973,N_4759);
and U5145 (N_5145,N_4874,N_4756);
and U5146 (N_5146,N_4871,N_4854);
or U5147 (N_5147,N_4883,N_4997);
or U5148 (N_5148,N_4912,N_4826);
nand U5149 (N_5149,N_4970,N_4899);
xnor U5150 (N_5150,N_4906,N_4923);
nor U5151 (N_5151,N_4829,N_4789);
or U5152 (N_5152,N_4974,N_4985);
and U5153 (N_5153,N_4934,N_4855);
nor U5154 (N_5154,N_4798,N_4915);
nand U5155 (N_5155,N_4912,N_4963);
nor U5156 (N_5156,N_4806,N_4934);
and U5157 (N_5157,N_4901,N_4853);
nor U5158 (N_5158,N_4936,N_4924);
or U5159 (N_5159,N_4997,N_4993);
nand U5160 (N_5160,N_4983,N_4950);
nand U5161 (N_5161,N_4754,N_4911);
and U5162 (N_5162,N_4799,N_4830);
or U5163 (N_5163,N_4892,N_4891);
and U5164 (N_5164,N_4842,N_4981);
xnor U5165 (N_5165,N_4780,N_4881);
nand U5166 (N_5166,N_4924,N_4761);
xnor U5167 (N_5167,N_4862,N_4878);
nand U5168 (N_5168,N_4995,N_4931);
nand U5169 (N_5169,N_4853,N_4933);
or U5170 (N_5170,N_4967,N_4752);
and U5171 (N_5171,N_4784,N_4930);
xor U5172 (N_5172,N_4968,N_4932);
nor U5173 (N_5173,N_4776,N_4976);
nor U5174 (N_5174,N_4945,N_4789);
nand U5175 (N_5175,N_4934,N_4873);
or U5176 (N_5176,N_4971,N_4895);
and U5177 (N_5177,N_4966,N_4951);
or U5178 (N_5178,N_4927,N_4988);
or U5179 (N_5179,N_4841,N_4830);
nand U5180 (N_5180,N_4910,N_4839);
and U5181 (N_5181,N_4766,N_4967);
xnor U5182 (N_5182,N_4923,N_4892);
xnor U5183 (N_5183,N_4913,N_4940);
or U5184 (N_5184,N_4939,N_4828);
nand U5185 (N_5185,N_4796,N_4861);
nand U5186 (N_5186,N_4841,N_4796);
and U5187 (N_5187,N_4911,N_4812);
nand U5188 (N_5188,N_4881,N_4926);
nand U5189 (N_5189,N_4828,N_4998);
nor U5190 (N_5190,N_4876,N_4902);
xnor U5191 (N_5191,N_4864,N_4850);
and U5192 (N_5192,N_4880,N_4996);
nand U5193 (N_5193,N_4774,N_4816);
xnor U5194 (N_5194,N_4801,N_4948);
nor U5195 (N_5195,N_4848,N_4958);
nor U5196 (N_5196,N_4826,N_4840);
nor U5197 (N_5197,N_4999,N_4986);
xnor U5198 (N_5198,N_4940,N_4780);
xor U5199 (N_5199,N_4789,N_4962);
nand U5200 (N_5200,N_4949,N_4954);
xor U5201 (N_5201,N_4993,N_4928);
nor U5202 (N_5202,N_4807,N_4904);
and U5203 (N_5203,N_4985,N_4972);
nand U5204 (N_5204,N_4957,N_4838);
and U5205 (N_5205,N_4936,N_4990);
nand U5206 (N_5206,N_4785,N_4922);
nor U5207 (N_5207,N_4781,N_4822);
and U5208 (N_5208,N_4772,N_4799);
nand U5209 (N_5209,N_4768,N_4816);
xor U5210 (N_5210,N_4967,N_4937);
xor U5211 (N_5211,N_4878,N_4952);
and U5212 (N_5212,N_4884,N_4876);
and U5213 (N_5213,N_4888,N_4775);
nor U5214 (N_5214,N_4782,N_4947);
nor U5215 (N_5215,N_4916,N_4985);
nor U5216 (N_5216,N_4812,N_4990);
xor U5217 (N_5217,N_4828,N_4900);
or U5218 (N_5218,N_4844,N_4751);
nor U5219 (N_5219,N_4784,N_4949);
and U5220 (N_5220,N_4843,N_4932);
nor U5221 (N_5221,N_4990,N_4926);
or U5222 (N_5222,N_4918,N_4868);
nand U5223 (N_5223,N_4828,N_4792);
nand U5224 (N_5224,N_4826,N_4833);
nor U5225 (N_5225,N_4863,N_4832);
nor U5226 (N_5226,N_4958,N_4772);
nand U5227 (N_5227,N_4781,N_4940);
xnor U5228 (N_5228,N_4929,N_4971);
nor U5229 (N_5229,N_4798,N_4938);
and U5230 (N_5230,N_4968,N_4945);
or U5231 (N_5231,N_4987,N_4954);
and U5232 (N_5232,N_4766,N_4768);
nor U5233 (N_5233,N_4912,N_4925);
nand U5234 (N_5234,N_4955,N_4782);
and U5235 (N_5235,N_4793,N_4771);
and U5236 (N_5236,N_4970,N_4952);
nor U5237 (N_5237,N_4900,N_4909);
or U5238 (N_5238,N_4881,N_4992);
or U5239 (N_5239,N_4885,N_4956);
nand U5240 (N_5240,N_4795,N_4944);
xnor U5241 (N_5241,N_4860,N_4855);
and U5242 (N_5242,N_4755,N_4769);
or U5243 (N_5243,N_4951,N_4924);
and U5244 (N_5244,N_4864,N_4862);
nor U5245 (N_5245,N_4924,N_4781);
nor U5246 (N_5246,N_4974,N_4960);
nand U5247 (N_5247,N_4874,N_4837);
nand U5248 (N_5248,N_4858,N_4890);
nor U5249 (N_5249,N_4831,N_4860);
and U5250 (N_5250,N_5004,N_5074);
and U5251 (N_5251,N_5153,N_5042);
nor U5252 (N_5252,N_5244,N_5103);
or U5253 (N_5253,N_5065,N_5242);
nand U5254 (N_5254,N_5137,N_5161);
or U5255 (N_5255,N_5040,N_5022);
or U5256 (N_5256,N_5176,N_5214);
nor U5257 (N_5257,N_5182,N_5235);
nand U5258 (N_5258,N_5018,N_5194);
nand U5259 (N_5259,N_5102,N_5046);
or U5260 (N_5260,N_5197,N_5248);
nor U5261 (N_5261,N_5078,N_5032);
or U5262 (N_5262,N_5070,N_5014);
nor U5263 (N_5263,N_5213,N_5067);
or U5264 (N_5264,N_5057,N_5198);
and U5265 (N_5265,N_5174,N_5105);
nor U5266 (N_5266,N_5047,N_5052);
nand U5267 (N_5267,N_5024,N_5238);
nor U5268 (N_5268,N_5169,N_5144);
and U5269 (N_5269,N_5060,N_5071);
or U5270 (N_5270,N_5084,N_5013);
xor U5271 (N_5271,N_5231,N_5215);
nor U5272 (N_5272,N_5216,N_5100);
and U5273 (N_5273,N_5224,N_5126);
nand U5274 (N_5274,N_5033,N_5055);
nand U5275 (N_5275,N_5056,N_5012);
xnor U5276 (N_5276,N_5173,N_5116);
xnor U5277 (N_5277,N_5187,N_5066);
and U5278 (N_5278,N_5209,N_5124);
nand U5279 (N_5279,N_5145,N_5002);
nand U5280 (N_5280,N_5006,N_5119);
xnor U5281 (N_5281,N_5148,N_5072);
xor U5282 (N_5282,N_5247,N_5142);
nor U5283 (N_5283,N_5149,N_5234);
or U5284 (N_5284,N_5122,N_5051);
nor U5285 (N_5285,N_5164,N_5027);
or U5286 (N_5286,N_5021,N_5133);
nor U5287 (N_5287,N_5045,N_5156);
or U5288 (N_5288,N_5019,N_5107);
nor U5289 (N_5289,N_5097,N_5108);
xnor U5290 (N_5290,N_5157,N_5143);
xnor U5291 (N_5291,N_5186,N_5243);
xor U5292 (N_5292,N_5225,N_5087);
nor U5293 (N_5293,N_5167,N_5029);
nor U5294 (N_5294,N_5016,N_5058);
nand U5295 (N_5295,N_5123,N_5043);
or U5296 (N_5296,N_5104,N_5053);
nand U5297 (N_5297,N_5112,N_5220);
xnor U5298 (N_5298,N_5199,N_5177);
nor U5299 (N_5299,N_5218,N_5050);
or U5300 (N_5300,N_5237,N_5099);
and U5301 (N_5301,N_5236,N_5110);
or U5302 (N_5302,N_5191,N_5219);
nor U5303 (N_5303,N_5189,N_5203);
nor U5304 (N_5304,N_5227,N_5159);
or U5305 (N_5305,N_5121,N_5120);
nor U5306 (N_5306,N_5184,N_5230);
or U5307 (N_5307,N_5000,N_5217);
or U5308 (N_5308,N_5001,N_5008);
nand U5309 (N_5309,N_5246,N_5151);
nor U5310 (N_5310,N_5163,N_5106);
nand U5311 (N_5311,N_5059,N_5140);
nand U5312 (N_5312,N_5165,N_5201);
or U5313 (N_5313,N_5210,N_5168);
nor U5314 (N_5314,N_5079,N_5111);
or U5315 (N_5315,N_5023,N_5171);
nor U5316 (N_5316,N_5113,N_5205);
nand U5317 (N_5317,N_5075,N_5170);
or U5318 (N_5318,N_5146,N_5212);
or U5319 (N_5319,N_5017,N_5134);
nor U5320 (N_5320,N_5077,N_5125);
and U5321 (N_5321,N_5192,N_5025);
xor U5322 (N_5322,N_5090,N_5098);
nand U5323 (N_5323,N_5010,N_5132);
or U5324 (N_5324,N_5034,N_5085);
and U5325 (N_5325,N_5228,N_5094);
nand U5326 (N_5326,N_5041,N_5083);
nor U5327 (N_5327,N_5101,N_5005);
or U5328 (N_5328,N_5204,N_5152);
and U5329 (N_5329,N_5036,N_5135);
and U5330 (N_5330,N_5211,N_5208);
xor U5331 (N_5331,N_5179,N_5076);
or U5332 (N_5332,N_5185,N_5136);
nor U5333 (N_5333,N_5037,N_5068);
or U5334 (N_5334,N_5035,N_5180);
or U5335 (N_5335,N_5096,N_5223);
or U5336 (N_5336,N_5249,N_5115);
or U5337 (N_5337,N_5048,N_5088);
or U5338 (N_5338,N_5221,N_5232);
nor U5339 (N_5339,N_5039,N_5147);
or U5340 (N_5340,N_5114,N_5026);
nor U5341 (N_5341,N_5093,N_5160);
nor U5342 (N_5342,N_5206,N_5086);
xor U5343 (N_5343,N_5131,N_5241);
xor U5344 (N_5344,N_5109,N_5020);
nor U5345 (N_5345,N_5061,N_5073);
nand U5346 (N_5346,N_5089,N_5011);
xor U5347 (N_5347,N_5081,N_5183);
nand U5348 (N_5348,N_5155,N_5158);
or U5349 (N_5349,N_5229,N_5190);
and U5350 (N_5350,N_5196,N_5080);
nor U5351 (N_5351,N_5128,N_5172);
and U5352 (N_5352,N_5240,N_5031);
nor U5353 (N_5353,N_5139,N_5129);
or U5354 (N_5354,N_5162,N_5175);
and U5355 (N_5355,N_5188,N_5038);
nor U5356 (N_5356,N_5044,N_5233);
nand U5357 (N_5357,N_5028,N_5007);
nand U5358 (N_5358,N_5003,N_5069);
or U5359 (N_5359,N_5181,N_5063);
nand U5360 (N_5360,N_5062,N_5193);
nor U5361 (N_5361,N_5130,N_5166);
xnor U5362 (N_5362,N_5082,N_5226);
nand U5363 (N_5363,N_5239,N_5064);
and U5364 (N_5364,N_5141,N_5030);
xnor U5365 (N_5365,N_5154,N_5222);
xnor U5366 (N_5366,N_5138,N_5150);
and U5367 (N_5367,N_5009,N_5200);
nand U5368 (N_5368,N_5015,N_5092);
and U5369 (N_5369,N_5245,N_5091);
or U5370 (N_5370,N_5178,N_5054);
and U5371 (N_5371,N_5049,N_5207);
nand U5372 (N_5372,N_5195,N_5127);
nor U5373 (N_5373,N_5202,N_5117);
xor U5374 (N_5374,N_5118,N_5095);
xnor U5375 (N_5375,N_5036,N_5195);
nand U5376 (N_5376,N_5033,N_5141);
xnor U5377 (N_5377,N_5218,N_5225);
nand U5378 (N_5378,N_5085,N_5189);
xor U5379 (N_5379,N_5093,N_5241);
nor U5380 (N_5380,N_5242,N_5182);
nand U5381 (N_5381,N_5002,N_5110);
xnor U5382 (N_5382,N_5095,N_5087);
xor U5383 (N_5383,N_5118,N_5142);
nor U5384 (N_5384,N_5210,N_5180);
and U5385 (N_5385,N_5183,N_5078);
nor U5386 (N_5386,N_5100,N_5145);
or U5387 (N_5387,N_5154,N_5197);
nand U5388 (N_5388,N_5247,N_5172);
nor U5389 (N_5389,N_5018,N_5168);
or U5390 (N_5390,N_5082,N_5184);
nand U5391 (N_5391,N_5133,N_5232);
xnor U5392 (N_5392,N_5176,N_5164);
nor U5393 (N_5393,N_5059,N_5157);
nor U5394 (N_5394,N_5181,N_5108);
or U5395 (N_5395,N_5138,N_5182);
nand U5396 (N_5396,N_5194,N_5124);
or U5397 (N_5397,N_5242,N_5196);
nand U5398 (N_5398,N_5238,N_5122);
and U5399 (N_5399,N_5039,N_5223);
and U5400 (N_5400,N_5037,N_5106);
xnor U5401 (N_5401,N_5058,N_5212);
and U5402 (N_5402,N_5040,N_5158);
xor U5403 (N_5403,N_5102,N_5245);
or U5404 (N_5404,N_5153,N_5003);
and U5405 (N_5405,N_5173,N_5085);
nand U5406 (N_5406,N_5223,N_5107);
and U5407 (N_5407,N_5146,N_5111);
or U5408 (N_5408,N_5200,N_5044);
or U5409 (N_5409,N_5220,N_5053);
nand U5410 (N_5410,N_5134,N_5069);
nor U5411 (N_5411,N_5230,N_5143);
xnor U5412 (N_5412,N_5219,N_5117);
or U5413 (N_5413,N_5170,N_5018);
xnor U5414 (N_5414,N_5007,N_5095);
or U5415 (N_5415,N_5133,N_5002);
xor U5416 (N_5416,N_5227,N_5117);
and U5417 (N_5417,N_5204,N_5086);
or U5418 (N_5418,N_5011,N_5246);
nand U5419 (N_5419,N_5181,N_5137);
or U5420 (N_5420,N_5043,N_5059);
xnor U5421 (N_5421,N_5196,N_5171);
xor U5422 (N_5422,N_5040,N_5068);
xor U5423 (N_5423,N_5155,N_5193);
xnor U5424 (N_5424,N_5151,N_5063);
or U5425 (N_5425,N_5032,N_5084);
xnor U5426 (N_5426,N_5028,N_5074);
or U5427 (N_5427,N_5039,N_5216);
xor U5428 (N_5428,N_5033,N_5109);
nand U5429 (N_5429,N_5069,N_5188);
nor U5430 (N_5430,N_5228,N_5214);
xor U5431 (N_5431,N_5108,N_5026);
and U5432 (N_5432,N_5202,N_5084);
nor U5433 (N_5433,N_5191,N_5160);
and U5434 (N_5434,N_5145,N_5128);
xor U5435 (N_5435,N_5234,N_5109);
and U5436 (N_5436,N_5229,N_5223);
nor U5437 (N_5437,N_5045,N_5091);
or U5438 (N_5438,N_5000,N_5190);
nor U5439 (N_5439,N_5200,N_5101);
xnor U5440 (N_5440,N_5132,N_5194);
or U5441 (N_5441,N_5138,N_5013);
xnor U5442 (N_5442,N_5223,N_5038);
nand U5443 (N_5443,N_5198,N_5223);
xor U5444 (N_5444,N_5113,N_5201);
nand U5445 (N_5445,N_5160,N_5170);
or U5446 (N_5446,N_5110,N_5006);
and U5447 (N_5447,N_5107,N_5102);
and U5448 (N_5448,N_5093,N_5010);
or U5449 (N_5449,N_5041,N_5165);
and U5450 (N_5450,N_5219,N_5130);
nor U5451 (N_5451,N_5126,N_5199);
or U5452 (N_5452,N_5168,N_5223);
and U5453 (N_5453,N_5165,N_5100);
xnor U5454 (N_5454,N_5106,N_5183);
xor U5455 (N_5455,N_5040,N_5144);
nor U5456 (N_5456,N_5204,N_5080);
nand U5457 (N_5457,N_5147,N_5034);
xnor U5458 (N_5458,N_5089,N_5233);
nor U5459 (N_5459,N_5161,N_5209);
xor U5460 (N_5460,N_5172,N_5077);
nand U5461 (N_5461,N_5189,N_5105);
nor U5462 (N_5462,N_5193,N_5004);
nand U5463 (N_5463,N_5073,N_5087);
nand U5464 (N_5464,N_5083,N_5073);
and U5465 (N_5465,N_5000,N_5096);
nor U5466 (N_5466,N_5073,N_5023);
nor U5467 (N_5467,N_5105,N_5232);
or U5468 (N_5468,N_5233,N_5203);
nand U5469 (N_5469,N_5246,N_5134);
xnor U5470 (N_5470,N_5026,N_5191);
nor U5471 (N_5471,N_5004,N_5050);
and U5472 (N_5472,N_5005,N_5146);
or U5473 (N_5473,N_5159,N_5186);
xnor U5474 (N_5474,N_5010,N_5034);
nand U5475 (N_5475,N_5131,N_5098);
nor U5476 (N_5476,N_5105,N_5061);
or U5477 (N_5477,N_5052,N_5182);
xor U5478 (N_5478,N_5083,N_5015);
xnor U5479 (N_5479,N_5188,N_5070);
and U5480 (N_5480,N_5196,N_5217);
nor U5481 (N_5481,N_5128,N_5015);
and U5482 (N_5482,N_5028,N_5016);
nor U5483 (N_5483,N_5040,N_5199);
or U5484 (N_5484,N_5107,N_5070);
nand U5485 (N_5485,N_5068,N_5239);
nor U5486 (N_5486,N_5070,N_5074);
xnor U5487 (N_5487,N_5151,N_5136);
nor U5488 (N_5488,N_5187,N_5059);
and U5489 (N_5489,N_5208,N_5201);
nor U5490 (N_5490,N_5147,N_5005);
xnor U5491 (N_5491,N_5117,N_5037);
nand U5492 (N_5492,N_5085,N_5026);
and U5493 (N_5493,N_5006,N_5203);
or U5494 (N_5494,N_5154,N_5088);
and U5495 (N_5495,N_5148,N_5161);
or U5496 (N_5496,N_5219,N_5085);
or U5497 (N_5497,N_5208,N_5042);
nor U5498 (N_5498,N_5018,N_5103);
or U5499 (N_5499,N_5070,N_5199);
or U5500 (N_5500,N_5366,N_5266);
nor U5501 (N_5501,N_5417,N_5381);
and U5502 (N_5502,N_5470,N_5358);
and U5503 (N_5503,N_5308,N_5480);
nand U5504 (N_5504,N_5254,N_5345);
and U5505 (N_5505,N_5402,N_5310);
and U5506 (N_5506,N_5304,N_5473);
xor U5507 (N_5507,N_5374,N_5465);
nand U5508 (N_5508,N_5256,N_5413);
or U5509 (N_5509,N_5359,N_5336);
nand U5510 (N_5510,N_5388,N_5276);
xnor U5511 (N_5511,N_5466,N_5471);
nand U5512 (N_5512,N_5279,N_5347);
and U5513 (N_5513,N_5267,N_5327);
and U5514 (N_5514,N_5289,N_5269);
or U5515 (N_5515,N_5434,N_5485);
nor U5516 (N_5516,N_5460,N_5328);
xor U5517 (N_5517,N_5364,N_5394);
and U5518 (N_5518,N_5406,N_5319);
or U5519 (N_5519,N_5429,N_5362);
or U5520 (N_5520,N_5383,N_5463);
nor U5521 (N_5521,N_5421,N_5341);
xnor U5522 (N_5522,N_5457,N_5389);
or U5523 (N_5523,N_5492,N_5493);
or U5524 (N_5524,N_5378,N_5451);
and U5525 (N_5525,N_5399,N_5387);
or U5526 (N_5526,N_5324,N_5286);
nand U5527 (N_5527,N_5273,N_5301);
and U5528 (N_5528,N_5283,N_5281);
or U5529 (N_5529,N_5445,N_5295);
nand U5530 (N_5530,N_5302,N_5444);
and U5531 (N_5531,N_5390,N_5258);
and U5532 (N_5532,N_5271,N_5352);
and U5533 (N_5533,N_5326,N_5474);
or U5534 (N_5534,N_5317,N_5334);
or U5535 (N_5535,N_5385,N_5263);
xnor U5536 (N_5536,N_5433,N_5405);
or U5537 (N_5537,N_5348,N_5342);
xnor U5538 (N_5538,N_5330,N_5380);
nand U5539 (N_5539,N_5333,N_5370);
nor U5540 (N_5540,N_5409,N_5291);
and U5541 (N_5541,N_5490,N_5278);
or U5542 (N_5542,N_5322,N_5251);
and U5543 (N_5543,N_5284,N_5436);
or U5544 (N_5544,N_5277,N_5272);
or U5545 (N_5545,N_5343,N_5397);
or U5546 (N_5546,N_5264,N_5391);
xor U5547 (N_5547,N_5384,N_5270);
or U5548 (N_5548,N_5369,N_5478);
nor U5549 (N_5549,N_5250,N_5489);
and U5550 (N_5550,N_5346,N_5368);
xnor U5551 (N_5551,N_5339,N_5300);
xor U5552 (N_5552,N_5398,N_5375);
xnor U5553 (N_5553,N_5462,N_5325);
and U5554 (N_5554,N_5446,N_5303);
nor U5555 (N_5555,N_5453,N_5491);
and U5556 (N_5556,N_5497,N_5365);
nand U5557 (N_5557,N_5288,N_5297);
nand U5558 (N_5558,N_5257,N_5481);
and U5559 (N_5559,N_5332,N_5309);
nand U5560 (N_5560,N_5484,N_5475);
and U5561 (N_5561,N_5472,N_5262);
and U5562 (N_5562,N_5275,N_5344);
and U5563 (N_5563,N_5494,N_5442);
or U5564 (N_5564,N_5487,N_5454);
xor U5565 (N_5565,N_5408,N_5379);
xor U5566 (N_5566,N_5321,N_5392);
xnor U5567 (N_5567,N_5439,N_5313);
nand U5568 (N_5568,N_5448,N_5431);
and U5569 (N_5569,N_5456,N_5461);
nor U5570 (N_5570,N_5299,N_5427);
xnor U5571 (N_5571,N_5476,N_5354);
xnor U5572 (N_5572,N_5496,N_5298);
nor U5573 (N_5573,N_5292,N_5259);
nor U5574 (N_5574,N_5468,N_5360);
xnor U5575 (N_5575,N_5335,N_5495);
xor U5576 (N_5576,N_5411,N_5437);
and U5577 (N_5577,N_5320,N_5282);
and U5578 (N_5578,N_5420,N_5349);
xnor U5579 (N_5579,N_5418,N_5412);
nor U5580 (N_5580,N_5376,N_5287);
or U5581 (N_5581,N_5340,N_5268);
nor U5582 (N_5582,N_5416,N_5261);
nor U5583 (N_5583,N_5372,N_5395);
nand U5584 (N_5584,N_5438,N_5419);
nor U5585 (N_5585,N_5294,N_5305);
and U5586 (N_5586,N_5410,N_5355);
xor U5587 (N_5587,N_5440,N_5415);
and U5588 (N_5588,N_5255,N_5274);
nand U5589 (N_5589,N_5422,N_5373);
xnor U5590 (N_5590,N_5424,N_5425);
nand U5591 (N_5591,N_5403,N_5396);
nand U5592 (N_5592,N_5435,N_5323);
nand U5593 (N_5593,N_5331,N_5316);
or U5594 (N_5594,N_5338,N_5361);
nor U5595 (N_5595,N_5400,N_5293);
nand U5596 (N_5596,N_5459,N_5377);
and U5597 (N_5597,N_5467,N_5428);
nor U5598 (N_5598,N_5499,N_5486);
or U5599 (N_5599,N_5479,N_5318);
xor U5600 (N_5600,N_5469,N_5356);
and U5601 (N_5601,N_5458,N_5498);
or U5602 (N_5602,N_5280,N_5265);
nor U5603 (N_5603,N_5404,N_5426);
nor U5604 (N_5604,N_5464,N_5353);
xnor U5605 (N_5605,N_5329,N_5296);
or U5606 (N_5606,N_5357,N_5367);
nor U5607 (N_5607,N_5423,N_5393);
xnor U5608 (N_5608,N_5382,N_5371);
and U5609 (N_5609,N_5285,N_5350);
nand U5610 (N_5610,N_5351,N_5307);
or U5611 (N_5611,N_5482,N_5443);
nand U5612 (N_5612,N_5252,N_5447);
and U5613 (N_5613,N_5314,N_5477);
and U5614 (N_5614,N_5414,N_5450);
nand U5615 (N_5615,N_5449,N_5260);
nand U5616 (N_5616,N_5407,N_5363);
and U5617 (N_5617,N_5290,N_5306);
and U5618 (N_5618,N_5386,N_5432);
or U5619 (N_5619,N_5483,N_5430);
xnor U5620 (N_5620,N_5488,N_5455);
nor U5621 (N_5621,N_5452,N_5315);
nand U5622 (N_5622,N_5337,N_5312);
and U5623 (N_5623,N_5253,N_5401);
nand U5624 (N_5624,N_5311,N_5441);
nand U5625 (N_5625,N_5370,N_5455);
and U5626 (N_5626,N_5467,N_5495);
nand U5627 (N_5627,N_5400,N_5469);
nand U5628 (N_5628,N_5447,N_5478);
xnor U5629 (N_5629,N_5362,N_5405);
nor U5630 (N_5630,N_5409,N_5495);
or U5631 (N_5631,N_5434,N_5314);
and U5632 (N_5632,N_5254,N_5310);
or U5633 (N_5633,N_5459,N_5277);
nor U5634 (N_5634,N_5421,N_5311);
nor U5635 (N_5635,N_5388,N_5396);
xor U5636 (N_5636,N_5394,N_5301);
nand U5637 (N_5637,N_5302,N_5432);
nand U5638 (N_5638,N_5456,N_5341);
and U5639 (N_5639,N_5494,N_5291);
nand U5640 (N_5640,N_5297,N_5318);
and U5641 (N_5641,N_5336,N_5314);
xnor U5642 (N_5642,N_5417,N_5317);
and U5643 (N_5643,N_5353,N_5338);
and U5644 (N_5644,N_5259,N_5385);
nor U5645 (N_5645,N_5473,N_5426);
nand U5646 (N_5646,N_5254,N_5332);
nand U5647 (N_5647,N_5280,N_5471);
xor U5648 (N_5648,N_5375,N_5319);
nor U5649 (N_5649,N_5262,N_5277);
or U5650 (N_5650,N_5299,N_5364);
nor U5651 (N_5651,N_5377,N_5402);
and U5652 (N_5652,N_5412,N_5382);
or U5653 (N_5653,N_5253,N_5344);
xor U5654 (N_5654,N_5290,N_5291);
or U5655 (N_5655,N_5331,N_5355);
or U5656 (N_5656,N_5423,N_5487);
and U5657 (N_5657,N_5345,N_5253);
nor U5658 (N_5658,N_5426,N_5413);
nand U5659 (N_5659,N_5449,N_5486);
xnor U5660 (N_5660,N_5457,N_5382);
or U5661 (N_5661,N_5391,N_5314);
xor U5662 (N_5662,N_5400,N_5382);
or U5663 (N_5663,N_5274,N_5356);
and U5664 (N_5664,N_5353,N_5383);
nor U5665 (N_5665,N_5438,N_5291);
nand U5666 (N_5666,N_5456,N_5440);
nor U5667 (N_5667,N_5469,N_5287);
xnor U5668 (N_5668,N_5414,N_5333);
nor U5669 (N_5669,N_5462,N_5281);
xor U5670 (N_5670,N_5472,N_5334);
nand U5671 (N_5671,N_5352,N_5394);
nand U5672 (N_5672,N_5301,N_5390);
xor U5673 (N_5673,N_5291,N_5458);
nand U5674 (N_5674,N_5326,N_5365);
or U5675 (N_5675,N_5382,N_5438);
nor U5676 (N_5676,N_5336,N_5394);
and U5677 (N_5677,N_5374,N_5358);
or U5678 (N_5678,N_5286,N_5271);
or U5679 (N_5679,N_5344,N_5331);
xor U5680 (N_5680,N_5393,N_5326);
nor U5681 (N_5681,N_5447,N_5301);
xnor U5682 (N_5682,N_5460,N_5475);
and U5683 (N_5683,N_5393,N_5312);
or U5684 (N_5684,N_5414,N_5424);
and U5685 (N_5685,N_5293,N_5483);
or U5686 (N_5686,N_5386,N_5401);
nand U5687 (N_5687,N_5411,N_5431);
xor U5688 (N_5688,N_5339,N_5290);
nand U5689 (N_5689,N_5408,N_5295);
or U5690 (N_5690,N_5341,N_5323);
or U5691 (N_5691,N_5300,N_5496);
nor U5692 (N_5692,N_5441,N_5437);
and U5693 (N_5693,N_5273,N_5499);
nor U5694 (N_5694,N_5470,N_5301);
nand U5695 (N_5695,N_5308,N_5322);
and U5696 (N_5696,N_5435,N_5281);
nor U5697 (N_5697,N_5354,N_5356);
or U5698 (N_5698,N_5269,N_5358);
or U5699 (N_5699,N_5342,N_5290);
and U5700 (N_5700,N_5489,N_5308);
or U5701 (N_5701,N_5401,N_5480);
or U5702 (N_5702,N_5308,N_5397);
and U5703 (N_5703,N_5391,N_5495);
nor U5704 (N_5704,N_5394,N_5413);
nand U5705 (N_5705,N_5497,N_5451);
nand U5706 (N_5706,N_5365,N_5438);
nor U5707 (N_5707,N_5322,N_5378);
or U5708 (N_5708,N_5386,N_5340);
and U5709 (N_5709,N_5272,N_5472);
nor U5710 (N_5710,N_5335,N_5294);
nor U5711 (N_5711,N_5495,N_5497);
or U5712 (N_5712,N_5406,N_5250);
xnor U5713 (N_5713,N_5274,N_5282);
or U5714 (N_5714,N_5407,N_5345);
xor U5715 (N_5715,N_5392,N_5352);
xor U5716 (N_5716,N_5383,N_5278);
or U5717 (N_5717,N_5360,N_5412);
xnor U5718 (N_5718,N_5308,N_5499);
or U5719 (N_5719,N_5433,N_5422);
and U5720 (N_5720,N_5478,N_5311);
nor U5721 (N_5721,N_5403,N_5303);
nand U5722 (N_5722,N_5389,N_5251);
and U5723 (N_5723,N_5306,N_5272);
or U5724 (N_5724,N_5298,N_5475);
nand U5725 (N_5725,N_5365,N_5289);
xor U5726 (N_5726,N_5488,N_5476);
xnor U5727 (N_5727,N_5266,N_5491);
or U5728 (N_5728,N_5329,N_5449);
and U5729 (N_5729,N_5482,N_5377);
and U5730 (N_5730,N_5257,N_5488);
nand U5731 (N_5731,N_5265,N_5391);
and U5732 (N_5732,N_5373,N_5402);
nand U5733 (N_5733,N_5499,N_5350);
or U5734 (N_5734,N_5324,N_5403);
or U5735 (N_5735,N_5314,N_5320);
and U5736 (N_5736,N_5445,N_5279);
xor U5737 (N_5737,N_5291,N_5322);
nor U5738 (N_5738,N_5338,N_5306);
and U5739 (N_5739,N_5366,N_5454);
nand U5740 (N_5740,N_5301,N_5302);
nor U5741 (N_5741,N_5443,N_5459);
xor U5742 (N_5742,N_5445,N_5336);
and U5743 (N_5743,N_5373,N_5409);
and U5744 (N_5744,N_5342,N_5405);
nand U5745 (N_5745,N_5297,N_5368);
and U5746 (N_5746,N_5385,N_5374);
xnor U5747 (N_5747,N_5309,N_5333);
or U5748 (N_5748,N_5322,N_5361);
nand U5749 (N_5749,N_5348,N_5391);
xnor U5750 (N_5750,N_5538,N_5644);
nor U5751 (N_5751,N_5527,N_5632);
nand U5752 (N_5752,N_5590,N_5683);
xor U5753 (N_5753,N_5657,N_5748);
nor U5754 (N_5754,N_5731,N_5699);
xnor U5755 (N_5755,N_5548,N_5585);
and U5756 (N_5756,N_5529,N_5616);
xnor U5757 (N_5757,N_5743,N_5660);
nand U5758 (N_5758,N_5698,N_5719);
and U5759 (N_5759,N_5726,N_5613);
nand U5760 (N_5760,N_5667,N_5707);
or U5761 (N_5761,N_5673,N_5596);
nor U5762 (N_5762,N_5638,N_5706);
nor U5763 (N_5763,N_5532,N_5615);
or U5764 (N_5764,N_5542,N_5508);
or U5765 (N_5765,N_5691,N_5623);
nor U5766 (N_5766,N_5630,N_5588);
nor U5767 (N_5767,N_5601,N_5606);
xnor U5768 (N_5768,N_5663,N_5507);
nand U5769 (N_5769,N_5600,N_5633);
xnor U5770 (N_5770,N_5693,N_5723);
nand U5771 (N_5771,N_5736,N_5517);
or U5772 (N_5772,N_5564,N_5676);
xor U5773 (N_5773,N_5520,N_5629);
nand U5774 (N_5774,N_5689,N_5686);
xnor U5775 (N_5775,N_5655,N_5642);
xor U5776 (N_5776,N_5697,N_5591);
nand U5777 (N_5777,N_5652,N_5557);
nand U5778 (N_5778,N_5619,N_5576);
nor U5779 (N_5779,N_5682,N_5654);
and U5780 (N_5780,N_5622,N_5717);
nor U5781 (N_5781,N_5746,N_5627);
nand U5782 (N_5782,N_5561,N_5625);
xor U5783 (N_5783,N_5578,N_5549);
nor U5784 (N_5784,N_5537,N_5595);
xnor U5785 (N_5785,N_5546,N_5536);
or U5786 (N_5786,N_5742,N_5687);
xnor U5787 (N_5787,N_5666,N_5650);
nand U5788 (N_5788,N_5540,N_5565);
nor U5789 (N_5789,N_5580,N_5571);
nor U5790 (N_5790,N_5656,N_5711);
nor U5791 (N_5791,N_5525,N_5521);
and U5792 (N_5792,N_5643,N_5727);
and U5793 (N_5793,N_5603,N_5651);
nand U5794 (N_5794,N_5513,N_5505);
nand U5795 (N_5795,N_5688,N_5636);
xnor U5796 (N_5796,N_5749,N_5543);
and U5797 (N_5797,N_5647,N_5547);
nor U5798 (N_5798,N_5579,N_5514);
nor U5799 (N_5799,N_5744,N_5637);
xor U5800 (N_5800,N_5648,N_5570);
xnor U5801 (N_5801,N_5718,N_5678);
and U5802 (N_5802,N_5587,N_5518);
and U5803 (N_5803,N_5695,N_5554);
nand U5804 (N_5804,N_5530,N_5680);
and U5805 (N_5805,N_5611,N_5553);
or U5806 (N_5806,N_5541,N_5617);
and U5807 (N_5807,N_5690,N_5574);
xnor U5808 (N_5808,N_5685,N_5552);
or U5809 (N_5809,N_5669,N_5702);
and U5810 (N_5810,N_5604,N_5724);
nor U5811 (N_5811,N_5662,N_5694);
nand U5812 (N_5812,N_5701,N_5737);
nand U5813 (N_5813,N_5696,N_5664);
xnor U5814 (N_5814,N_5713,N_5586);
or U5815 (N_5815,N_5589,N_5524);
xor U5816 (N_5816,N_5634,N_5740);
or U5817 (N_5817,N_5516,N_5598);
nor U5818 (N_5818,N_5612,N_5593);
or U5819 (N_5819,N_5640,N_5741);
nand U5820 (N_5820,N_5668,N_5738);
and U5821 (N_5821,N_5631,N_5610);
or U5822 (N_5822,N_5583,N_5523);
nand U5823 (N_5823,N_5703,N_5665);
nand U5824 (N_5824,N_5670,N_5710);
or U5825 (N_5825,N_5658,N_5715);
nand U5826 (N_5826,N_5544,N_5645);
nand U5827 (N_5827,N_5735,N_5563);
nor U5828 (N_5828,N_5608,N_5684);
xor U5829 (N_5829,N_5692,N_5510);
and U5830 (N_5830,N_5620,N_5551);
nor U5831 (N_5831,N_5729,N_5705);
nand U5832 (N_5832,N_5621,N_5733);
xnor U5833 (N_5833,N_5599,N_5677);
xor U5834 (N_5834,N_5716,N_5671);
xnor U5835 (N_5835,N_5605,N_5528);
xor U5836 (N_5836,N_5567,N_5728);
and U5837 (N_5837,N_5511,N_5515);
nor U5838 (N_5838,N_5573,N_5641);
xnor U5839 (N_5839,N_5725,N_5635);
nand U5840 (N_5840,N_5675,N_5609);
nor U5841 (N_5841,N_5584,N_5721);
nor U5842 (N_5842,N_5720,N_5597);
nor U5843 (N_5843,N_5581,N_5562);
or U5844 (N_5844,N_5674,N_5639);
nand U5845 (N_5845,N_5592,N_5672);
nand U5846 (N_5846,N_5504,N_5512);
nand U5847 (N_5847,N_5569,N_5577);
or U5848 (N_5848,N_5502,N_5526);
nor U5849 (N_5849,N_5730,N_5556);
and U5850 (N_5850,N_5659,N_5626);
nor U5851 (N_5851,N_5534,N_5722);
nand U5852 (N_5852,N_5535,N_5594);
nor U5853 (N_5853,N_5602,N_5539);
nand U5854 (N_5854,N_5501,N_5566);
and U5855 (N_5855,N_5503,N_5681);
or U5856 (N_5856,N_5555,N_5661);
and U5857 (N_5857,N_5614,N_5531);
nor U5858 (N_5858,N_5500,N_5653);
xor U5859 (N_5859,N_5704,N_5646);
or U5860 (N_5860,N_5732,N_5739);
nor U5861 (N_5861,N_5506,N_5560);
nor U5862 (N_5862,N_5700,N_5628);
nand U5863 (N_5863,N_5708,N_5568);
xor U5864 (N_5864,N_5575,N_5519);
and U5865 (N_5865,N_5712,N_5509);
nor U5866 (N_5866,N_5607,N_5559);
nor U5867 (N_5867,N_5533,N_5582);
nor U5868 (N_5868,N_5709,N_5572);
nor U5869 (N_5869,N_5522,N_5649);
and U5870 (N_5870,N_5734,N_5550);
xnor U5871 (N_5871,N_5624,N_5545);
and U5872 (N_5872,N_5618,N_5679);
and U5873 (N_5873,N_5745,N_5747);
nand U5874 (N_5874,N_5558,N_5714);
or U5875 (N_5875,N_5744,N_5536);
or U5876 (N_5876,N_5602,N_5598);
and U5877 (N_5877,N_5695,N_5659);
nand U5878 (N_5878,N_5609,N_5581);
and U5879 (N_5879,N_5709,N_5538);
nand U5880 (N_5880,N_5615,N_5623);
nand U5881 (N_5881,N_5644,N_5577);
or U5882 (N_5882,N_5661,N_5551);
or U5883 (N_5883,N_5749,N_5680);
xor U5884 (N_5884,N_5546,N_5582);
or U5885 (N_5885,N_5507,N_5702);
nand U5886 (N_5886,N_5659,N_5578);
or U5887 (N_5887,N_5726,N_5740);
nand U5888 (N_5888,N_5749,N_5649);
or U5889 (N_5889,N_5502,N_5651);
xor U5890 (N_5890,N_5591,N_5554);
nand U5891 (N_5891,N_5531,N_5735);
or U5892 (N_5892,N_5670,N_5714);
and U5893 (N_5893,N_5550,N_5542);
xnor U5894 (N_5894,N_5585,N_5682);
xnor U5895 (N_5895,N_5506,N_5527);
xnor U5896 (N_5896,N_5651,N_5719);
and U5897 (N_5897,N_5714,N_5567);
xor U5898 (N_5898,N_5554,N_5650);
xor U5899 (N_5899,N_5575,N_5585);
and U5900 (N_5900,N_5611,N_5618);
nor U5901 (N_5901,N_5561,N_5679);
nand U5902 (N_5902,N_5557,N_5632);
and U5903 (N_5903,N_5631,N_5675);
or U5904 (N_5904,N_5529,N_5507);
xnor U5905 (N_5905,N_5636,N_5522);
and U5906 (N_5906,N_5586,N_5532);
nand U5907 (N_5907,N_5539,N_5500);
nand U5908 (N_5908,N_5525,N_5655);
xnor U5909 (N_5909,N_5598,N_5636);
or U5910 (N_5910,N_5506,N_5692);
or U5911 (N_5911,N_5587,N_5647);
and U5912 (N_5912,N_5636,N_5502);
nand U5913 (N_5913,N_5739,N_5678);
or U5914 (N_5914,N_5687,N_5635);
and U5915 (N_5915,N_5620,N_5623);
and U5916 (N_5916,N_5727,N_5649);
or U5917 (N_5917,N_5562,N_5557);
or U5918 (N_5918,N_5554,N_5692);
nor U5919 (N_5919,N_5665,N_5612);
and U5920 (N_5920,N_5639,N_5582);
and U5921 (N_5921,N_5511,N_5586);
xnor U5922 (N_5922,N_5711,N_5613);
nand U5923 (N_5923,N_5625,N_5650);
xnor U5924 (N_5924,N_5661,N_5594);
or U5925 (N_5925,N_5644,N_5678);
and U5926 (N_5926,N_5746,N_5609);
and U5927 (N_5927,N_5650,N_5563);
nor U5928 (N_5928,N_5742,N_5521);
and U5929 (N_5929,N_5592,N_5731);
or U5930 (N_5930,N_5713,N_5732);
or U5931 (N_5931,N_5562,N_5541);
nor U5932 (N_5932,N_5525,N_5528);
or U5933 (N_5933,N_5512,N_5740);
or U5934 (N_5934,N_5724,N_5581);
nor U5935 (N_5935,N_5553,N_5523);
nor U5936 (N_5936,N_5543,N_5527);
and U5937 (N_5937,N_5561,N_5583);
or U5938 (N_5938,N_5645,N_5654);
or U5939 (N_5939,N_5536,N_5703);
and U5940 (N_5940,N_5578,N_5586);
nor U5941 (N_5941,N_5632,N_5520);
or U5942 (N_5942,N_5553,N_5642);
xor U5943 (N_5943,N_5634,N_5584);
or U5944 (N_5944,N_5616,N_5610);
nand U5945 (N_5945,N_5558,N_5582);
xor U5946 (N_5946,N_5513,N_5638);
xor U5947 (N_5947,N_5553,N_5594);
and U5948 (N_5948,N_5694,N_5563);
or U5949 (N_5949,N_5509,N_5628);
xor U5950 (N_5950,N_5715,N_5652);
or U5951 (N_5951,N_5662,N_5663);
nor U5952 (N_5952,N_5528,N_5539);
xnor U5953 (N_5953,N_5583,N_5575);
nor U5954 (N_5954,N_5519,N_5610);
xor U5955 (N_5955,N_5661,N_5743);
nand U5956 (N_5956,N_5637,N_5570);
or U5957 (N_5957,N_5730,N_5513);
nor U5958 (N_5958,N_5596,N_5573);
nor U5959 (N_5959,N_5555,N_5594);
nor U5960 (N_5960,N_5656,N_5539);
and U5961 (N_5961,N_5634,N_5597);
nor U5962 (N_5962,N_5650,N_5700);
xor U5963 (N_5963,N_5738,N_5670);
nand U5964 (N_5964,N_5741,N_5641);
nor U5965 (N_5965,N_5708,N_5727);
nor U5966 (N_5966,N_5739,N_5567);
or U5967 (N_5967,N_5675,N_5655);
nor U5968 (N_5968,N_5559,N_5710);
nand U5969 (N_5969,N_5543,N_5672);
xor U5970 (N_5970,N_5529,N_5666);
xor U5971 (N_5971,N_5509,N_5749);
or U5972 (N_5972,N_5738,N_5747);
nor U5973 (N_5973,N_5566,N_5529);
or U5974 (N_5974,N_5502,N_5642);
xor U5975 (N_5975,N_5636,N_5716);
or U5976 (N_5976,N_5708,N_5683);
nand U5977 (N_5977,N_5594,N_5653);
or U5978 (N_5978,N_5505,N_5504);
or U5979 (N_5979,N_5650,N_5529);
nand U5980 (N_5980,N_5551,N_5652);
nand U5981 (N_5981,N_5729,N_5562);
and U5982 (N_5982,N_5620,N_5726);
nand U5983 (N_5983,N_5654,N_5504);
or U5984 (N_5984,N_5627,N_5504);
and U5985 (N_5985,N_5603,N_5648);
nand U5986 (N_5986,N_5502,N_5739);
xor U5987 (N_5987,N_5547,N_5614);
nor U5988 (N_5988,N_5653,N_5544);
nor U5989 (N_5989,N_5535,N_5561);
nand U5990 (N_5990,N_5625,N_5698);
xnor U5991 (N_5991,N_5698,N_5637);
nor U5992 (N_5992,N_5679,N_5698);
and U5993 (N_5993,N_5505,N_5732);
nand U5994 (N_5994,N_5645,N_5725);
nand U5995 (N_5995,N_5694,N_5610);
or U5996 (N_5996,N_5717,N_5590);
nor U5997 (N_5997,N_5706,N_5586);
or U5998 (N_5998,N_5678,N_5542);
and U5999 (N_5999,N_5635,N_5512);
xor U6000 (N_6000,N_5891,N_5769);
and U6001 (N_6001,N_5852,N_5850);
nor U6002 (N_6002,N_5954,N_5776);
or U6003 (N_6003,N_5851,N_5909);
nand U6004 (N_6004,N_5911,N_5790);
nor U6005 (N_6005,N_5932,N_5955);
or U6006 (N_6006,N_5773,N_5849);
or U6007 (N_6007,N_5882,N_5996);
nor U6008 (N_6008,N_5788,N_5857);
nor U6009 (N_6009,N_5887,N_5951);
or U6010 (N_6010,N_5876,N_5984);
nand U6011 (N_6011,N_5783,N_5949);
xor U6012 (N_6012,N_5836,N_5920);
or U6013 (N_6013,N_5860,N_5793);
nand U6014 (N_6014,N_5976,N_5943);
nor U6015 (N_6015,N_5966,N_5774);
nand U6016 (N_6016,N_5960,N_5754);
xnor U6017 (N_6017,N_5829,N_5761);
or U6018 (N_6018,N_5824,N_5884);
nor U6019 (N_6019,N_5843,N_5902);
nor U6020 (N_6020,N_5822,N_5979);
xnor U6021 (N_6021,N_5794,N_5883);
nor U6022 (N_6022,N_5903,N_5972);
and U6023 (N_6023,N_5771,N_5778);
xnor U6024 (N_6024,N_5861,N_5845);
nand U6025 (N_6025,N_5812,N_5995);
xor U6026 (N_6026,N_5848,N_5875);
nor U6027 (N_6027,N_5913,N_5872);
and U6028 (N_6028,N_5914,N_5839);
nand U6029 (N_6029,N_5844,N_5760);
or U6030 (N_6030,N_5838,N_5923);
nand U6031 (N_6031,N_5963,N_5803);
or U6032 (N_6032,N_5928,N_5929);
and U6033 (N_6033,N_5987,N_5953);
nand U6034 (N_6034,N_5892,N_5762);
nor U6035 (N_6035,N_5968,N_5781);
nor U6036 (N_6036,N_5975,N_5772);
and U6037 (N_6037,N_5965,N_5919);
or U6038 (N_6038,N_5944,N_5897);
or U6039 (N_6039,N_5795,N_5858);
xnor U6040 (N_6040,N_5874,N_5950);
xor U6041 (N_6041,N_5898,N_5853);
nor U6042 (N_6042,N_5910,N_5786);
nor U6043 (N_6043,N_5904,N_5927);
and U6044 (N_6044,N_5999,N_5820);
xor U6045 (N_6045,N_5888,N_5937);
xor U6046 (N_6046,N_5988,N_5957);
xnor U6047 (N_6047,N_5905,N_5863);
nor U6048 (N_6048,N_5986,N_5756);
xor U6049 (N_6049,N_5907,N_5877);
xnor U6050 (N_6050,N_5813,N_5916);
and U6051 (N_6051,N_5895,N_5994);
or U6052 (N_6052,N_5862,N_5952);
nor U6053 (N_6053,N_5819,N_5826);
xor U6054 (N_6054,N_5871,N_5989);
and U6055 (N_6055,N_5997,N_5973);
xnor U6056 (N_6056,N_5921,N_5945);
nor U6057 (N_6057,N_5789,N_5880);
or U6058 (N_6058,N_5969,N_5924);
xnor U6059 (N_6059,N_5942,N_5805);
xor U6060 (N_6060,N_5935,N_5936);
and U6061 (N_6061,N_5757,N_5828);
or U6062 (N_6062,N_5970,N_5869);
xnor U6063 (N_6063,N_5814,N_5753);
nand U6064 (N_6064,N_5792,N_5796);
xnor U6065 (N_6065,N_5859,N_5815);
and U6066 (N_6066,N_5870,N_5981);
and U6067 (N_6067,N_5775,N_5879);
or U6068 (N_6068,N_5835,N_5817);
xor U6069 (N_6069,N_5833,N_5971);
and U6070 (N_6070,N_5930,N_5938);
nor U6071 (N_6071,N_5977,N_5800);
and U6072 (N_6072,N_5847,N_5777);
or U6073 (N_6073,N_5992,N_5961);
nand U6074 (N_6074,N_5865,N_5983);
or U6075 (N_6075,N_5758,N_5808);
and U6076 (N_6076,N_5752,N_5856);
nor U6077 (N_6077,N_5889,N_5809);
xor U6078 (N_6078,N_5922,N_5802);
nand U6079 (N_6079,N_5918,N_5751);
xor U6080 (N_6080,N_5827,N_5867);
and U6081 (N_6081,N_5958,N_5925);
nor U6082 (N_6082,N_5791,N_5787);
nand U6083 (N_6083,N_5908,N_5896);
nor U6084 (N_6084,N_5830,N_5941);
nor U6085 (N_6085,N_5807,N_5837);
xnor U6086 (N_6086,N_5782,N_5939);
nand U6087 (N_6087,N_5926,N_5811);
nand U6088 (N_6088,N_5825,N_5946);
xnor U6089 (N_6089,N_5810,N_5799);
and U6090 (N_6090,N_5940,N_5956);
or U6091 (N_6091,N_5900,N_5846);
and U6092 (N_6092,N_5947,N_5873);
nand U6093 (N_6093,N_5821,N_5784);
nor U6094 (N_6094,N_5933,N_5964);
xnor U6095 (N_6095,N_5831,N_5818);
nand U6096 (N_6096,N_5764,N_5834);
xor U6097 (N_6097,N_5982,N_5823);
or U6098 (N_6098,N_5779,N_5750);
or U6099 (N_6099,N_5980,N_5755);
nor U6100 (N_6100,N_5780,N_5917);
nor U6101 (N_6101,N_5993,N_5785);
or U6102 (N_6102,N_5934,N_5890);
nand U6103 (N_6103,N_5866,N_5974);
nor U6104 (N_6104,N_5854,N_5763);
or U6105 (N_6105,N_5978,N_5894);
or U6106 (N_6106,N_5948,N_5840);
and U6107 (N_6107,N_5770,N_5832);
xor U6108 (N_6108,N_5998,N_5985);
xnor U6109 (N_6109,N_5806,N_5766);
or U6110 (N_6110,N_5855,N_5798);
nor U6111 (N_6111,N_5959,N_5768);
or U6112 (N_6112,N_5886,N_5893);
xor U6113 (N_6113,N_5816,N_5962);
and U6114 (N_6114,N_5915,N_5991);
nand U6115 (N_6115,N_5797,N_5804);
nor U6116 (N_6116,N_5801,N_5912);
or U6117 (N_6117,N_5885,N_5868);
or U6118 (N_6118,N_5841,N_5990);
or U6119 (N_6119,N_5967,N_5767);
nor U6120 (N_6120,N_5765,N_5842);
nand U6121 (N_6121,N_5881,N_5906);
nand U6122 (N_6122,N_5931,N_5878);
xnor U6123 (N_6123,N_5759,N_5899);
xor U6124 (N_6124,N_5901,N_5864);
and U6125 (N_6125,N_5763,N_5937);
nor U6126 (N_6126,N_5816,N_5770);
and U6127 (N_6127,N_5952,N_5971);
and U6128 (N_6128,N_5974,N_5969);
nor U6129 (N_6129,N_5958,N_5833);
xor U6130 (N_6130,N_5949,N_5904);
or U6131 (N_6131,N_5864,N_5862);
xor U6132 (N_6132,N_5849,N_5986);
nor U6133 (N_6133,N_5850,N_5760);
or U6134 (N_6134,N_5805,N_5913);
nand U6135 (N_6135,N_5819,N_5815);
nor U6136 (N_6136,N_5815,N_5998);
nand U6137 (N_6137,N_5973,N_5953);
xnor U6138 (N_6138,N_5879,N_5766);
and U6139 (N_6139,N_5955,N_5925);
and U6140 (N_6140,N_5961,N_5829);
or U6141 (N_6141,N_5961,N_5982);
and U6142 (N_6142,N_5916,N_5751);
nand U6143 (N_6143,N_5775,N_5830);
or U6144 (N_6144,N_5950,N_5949);
or U6145 (N_6145,N_5902,N_5926);
or U6146 (N_6146,N_5923,N_5994);
nand U6147 (N_6147,N_5766,N_5977);
or U6148 (N_6148,N_5989,N_5760);
nor U6149 (N_6149,N_5833,N_5889);
nand U6150 (N_6150,N_5973,N_5894);
nand U6151 (N_6151,N_5859,N_5981);
nor U6152 (N_6152,N_5982,N_5918);
nor U6153 (N_6153,N_5943,N_5909);
or U6154 (N_6154,N_5925,N_5836);
nand U6155 (N_6155,N_5874,N_5843);
nor U6156 (N_6156,N_5787,N_5835);
or U6157 (N_6157,N_5920,N_5752);
or U6158 (N_6158,N_5884,N_5885);
and U6159 (N_6159,N_5751,N_5777);
nor U6160 (N_6160,N_5774,N_5819);
nand U6161 (N_6161,N_5869,N_5824);
or U6162 (N_6162,N_5882,N_5798);
nor U6163 (N_6163,N_5837,N_5993);
nand U6164 (N_6164,N_5978,N_5820);
nor U6165 (N_6165,N_5852,N_5760);
nor U6166 (N_6166,N_5758,N_5967);
or U6167 (N_6167,N_5919,N_5780);
nand U6168 (N_6168,N_5750,N_5758);
xnor U6169 (N_6169,N_5762,N_5898);
nand U6170 (N_6170,N_5919,N_5879);
nor U6171 (N_6171,N_5981,N_5932);
or U6172 (N_6172,N_5938,N_5936);
xnor U6173 (N_6173,N_5819,N_5910);
or U6174 (N_6174,N_5806,N_5850);
xor U6175 (N_6175,N_5785,N_5860);
and U6176 (N_6176,N_5928,N_5761);
nor U6177 (N_6177,N_5947,N_5879);
nor U6178 (N_6178,N_5855,N_5859);
or U6179 (N_6179,N_5953,N_5845);
nor U6180 (N_6180,N_5816,N_5872);
nor U6181 (N_6181,N_5971,N_5844);
or U6182 (N_6182,N_5969,N_5871);
xnor U6183 (N_6183,N_5964,N_5865);
and U6184 (N_6184,N_5822,N_5837);
nor U6185 (N_6185,N_5907,N_5844);
nand U6186 (N_6186,N_5967,N_5762);
or U6187 (N_6187,N_5753,N_5784);
and U6188 (N_6188,N_5811,N_5896);
xor U6189 (N_6189,N_5956,N_5828);
xnor U6190 (N_6190,N_5950,N_5797);
nand U6191 (N_6191,N_5828,N_5897);
xor U6192 (N_6192,N_5997,N_5856);
and U6193 (N_6193,N_5837,N_5862);
and U6194 (N_6194,N_5801,N_5830);
and U6195 (N_6195,N_5882,N_5820);
nand U6196 (N_6196,N_5847,N_5857);
and U6197 (N_6197,N_5989,N_5962);
and U6198 (N_6198,N_5831,N_5825);
or U6199 (N_6199,N_5863,N_5939);
nor U6200 (N_6200,N_5930,N_5856);
xor U6201 (N_6201,N_5857,N_5770);
nor U6202 (N_6202,N_5767,N_5962);
or U6203 (N_6203,N_5848,N_5968);
nor U6204 (N_6204,N_5851,N_5813);
or U6205 (N_6205,N_5885,N_5785);
or U6206 (N_6206,N_5757,N_5816);
and U6207 (N_6207,N_5901,N_5983);
xnor U6208 (N_6208,N_5915,N_5863);
nand U6209 (N_6209,N_5949,N_5828);
xnor U6210 (N_6210,N_5751,N_5817);
nand U6211 (N_6211,N_5851,N_5889);
and U6212 (N_6212,N_5876,N_5846);
or U6213 (N_6213,N_5880,N_5832);
nand U6214 (N_6214,N_5929,N_5947);
or U6215 (N_6215,N_5916,N_5761);
xnor U6216 (N_6216,N_5794,N_5770);
xor U6217 (N_6217,N_5980,N_5832);
and U6218 (N_6218,N_5874,N_5894);
nand U6219 (N_6219,N_5759,N_5910);
and U6220 (N_6220,N_5864,N_5836);
nand U6221 (N_6221,N_5802,N_5793);
and U6222 (N_6222,N_5948,N_5991);
nand U6223 (N_6223,N_5887,N_5766);
and U6224 (N_6224,N_5772,N_5787);
nor U6225 (N_6225,N_5977,N_5909);
or U6226 (N_6226,N_5788,N_5862);
xnor U6227 (N_6227,N_5853,N_5940);
nand U6228 (N_6228,N_5765,N_5773);
xnor U6229 (N_6229,N_5995,N_5904);
xnor U6230 (N_6230,N_5768,N_5831);
and U6231 (N_6231,N_5846,N_5883);
nand U6232 (N_6232,N_5930,N_5886);
nand U6233 (N_6233,N_5959,N_5908);
xnor U6234 (N_6234,N_5920,N_5866);
or U6235 (N_6235,N_5858,N_5960);
or U6236 (N_6236,N_5862,N_5866);
nand U6237 (N_6237,N_5921,N_5916);
and U6238 (N_6238,N_5976,N_5754);
and U6239 (N_6239,N_5945,N_5930);
nand U6240 (N_6240,N_5877,N_5853);
and U6241 (N_6241,N_5925,N_5807);
or U6242 (N_6242,N_5801,N_5834);
nor U6243 (N_6243,N_5783,N_5782);
nor U6244 (N_6244,N_5753,N_5931);
and U6245 (N_6245,N_5765,N_5783);
nor U6246 (N_6246,N_5981,N_5778);
xnor U6247 (N_6247,N_5919,N_5812);
or U6248 (N_6248,N_5936,N_5799);
or U6249 (N_6249,N_5893,N_5890);
nand U6250 (N_6250,N_6010,N_6191);
or U6251 (N_6251,N_6069,N_6122);
or U6252 (N_6252,N_6098,N_6225);
nor U6253 (N_6253,N_6068,N_6008);
nor U6254 (N_6254,N_6058,N_6137);
nand U6255 (N_6255,N_6129,N_6094);
or U6256 (N_6256,N_6207,N_6194);
nor U6257 (N_6257,N_6140,N_6082);
or U6258 (N_6258,N_6245,N_6062);
and U6259 (N_6259,N_6190,N_6220);
nand U6260 (N_6260,N_6127,N_6072);
nand U6261 (N_6261,N_6096,N_6126);
nand U6262 (N_6262,N_6232,N_6104);
xor U6263 (N_6263,N_6040,N_6027);
xor U6264 (N_6264,N_6236,N_6043);
or U6265 (N_6265,N_6026,N_6198);
or U6266 (N_6266,N_6235,N_6193);
and U6267 (N_6267,N_6186,N_6172);
xor U6268 (N_6268,N_6167,N_6200);
nand U6269 (N_6269,N_6124,N_6176);
nand U6270 (N_6270,N_6076,N_6163);
nor U6271 (N_6271,N_6011,N_6174);
or U6272 (N_6272,N_6215,N_6083);
or U6273 (N_6273,N_6239,N_6202);
nor U6274 (N_6274,N_6044,N_6196);
or U6275 (N_6275,N_6237,N_6079);
nor U6276 (N_6276,N_6020,N_6209);
and U6277 (N_6277,N_6070,N_6180);
nor U6278 (N_6278,N_6107,N_6133);
or U6279 (N_6279,N_6241,N_6014);
nor U6280 (N_6280,N_6115,N_6086);
and U6281 (N_6281,N_6222,N_6030);
or U6282 (N_6282,N_6165,N_6065);
and U6283 (N_6283,N_6005,N_6000);
nor U6284 (N_6284,N_6218,N_6130);
and U6285 (N_6285,N_6092,N_6113);
nor U6286 (N_6286,N_6166,N_6002);
or U6287 (N_6287,N_6145,N_6021);
xor U6288 (N_6288,N_6118,N_6114);
xor U6289 (N_6289,N_6057,N_6231);
nor U6290 (N_6290,N_6217,N_6168);
and U6291 (N_6291,N_6012,N_6153);
xnor U6292 (N_6292,N_6154,N_6138);
nor U6293 (N_6293,N_6141,N_6059);
nor U6294 (N_6294,N_6242,N_6224);
nand U6295 (N_6295,N_6152,N_6089);
or U6296 (N_6296,N_6018,N_6112);
xor U6297 (N_6297,N_6189,N_6050);
or U6298 (N_6298,N_6071,N_6054);
nor U6299 (N_6299,N_6042,N_6185);
nor U6300 (N_6300,N_6017,N_6009);
nand U6301 (N_6301,N_6240,N_6169);
and U6302 (N_6302,N_6234,N_6134);
nand U6303 (N_6303,N_6210,N_6181);
or U6304 (N_6304,N_6045,N_6187);
xor U6305 (N_6305,N_6188,N_6146);
or U6306 (N_6306,N_6171,N_6119);
or U6307 (N_6307,N_6073,N_6004);
and U6308 (N_6308,N_6136,N_6074);
nand U6309 (N_6309,N_6025,N_6162);
nand U6310 (N_6310,N_6048,N_6080);
or U6311 (N_6311,N_6227,N_6214);
nor U6312 (N_6312,N_6006,N_6206);
nor U6313 (N_6313,N_6230,N_6109);
and U6314 (N_6314,N_6033,N_6244);
nor U6315 (N_6315,N_6249,N_6221);
nand U6316 (N_6316,N_6106,N_6216);
nand U6317 (N_6317,N_6055,N_6173);
xor U6318 (N_6318,N_6147,N_6170);
nor U6319 (N_6319,N_6229,N_6144);
nor U6320 (N_6320,N_6031,N_6039);
or U6321 (N_6321,N_6157,N_6197);
and U6322 (N_6322,N_6024,N_6238);
or U6323 (N_6323,N_6121,N_6120);
and U6324 (N_6324,N_6051,N_6116);
nor U6325 (N_6325,N_6226,N_6077);
and U6326 (N_6326,N_6093,N_6060);
nand U6327 (N_6327,N_6164,N_6123);
or U6328 (N_6328,N_6228,N_6067);
nor U6329 (N_6329,N_6087,N_6016);
xnor U6330 (N_6330,N_6132,N_6243);
nor U6331 (N_6331,N_6184,N_6117);
xor U6332 (N_6332,N_6212,N_6182);
xor U6333 (N_6333,N_6110,N_6046);
or U6334 (N_6334,N_6028,N_6178);
and U6335 (N_6335,N_6001,N_6159);
xor U6336 (N_6336,N_6063,N_6203);
xnor U6337 (N_6337,N_6177,N_6108);
or U6338 (N_6338,N_6248,N_6183);
or U6339 (N_6339,N_6007,N_6155);
nor U6340 (N_6340,N_6125,N_6084);
and U6341 (N_6341,N_6208,N_6037);
and U6342 (N_6342,N_6175,N_6075);
xnor U6343 (N_6343,N_6158,N_6029);
nor U6344 (N_6344,N_6233,N_6085);
nor U6345 (N_6345,N_6078,N_6205);
and U6346 (N_6346,N_6036,N_6064);
nor U6347 (N_6347,N_6199,N_6213);
or U6348 (N_6348,N_6102,N_6211);
xnor U6349 (N_6349,N_6111,N_6105);
nor U6350 (N_6350,N_6139,N_6179);
and U6351 (N_6351,N_6148,N_6081);
nand U6352 (N_6352,N_6150,N_6023);
nand U6353 (N_6353,N_6246,N_6056);
or U6354 (N_6354,N_6161,N_6049);
and U6355 (N_6355,N_6149,N_6131);
xnor U6356 (N_6356,N_6160,N_6223);
or U6357 (N_6357,N_6022,N_6143);
or U6358 (N_6358,N_6192,N_6103);
or U6359 (N_6359,N_6066,N_6099);
nand U6360 (N_6360,N_6041,N_6156);
nor U6361 (N_6361,N_6061,N_6100);
xor U6362 (N_6362,N_6135,N_6090);
nor U6363 (N_6363,N_6052,N_6088);
or U6364 (N_6364,N_6247,N_6219);
nand U6365 (N_6365,N_6013,N_6097);
nor U6366 (N_6366,N_6015,N_6095);
nand U6367 (N_6367,N_6047,N_6091);
xor U6368 (N_6368,N_6019,N_6142);
nand U6369 (N_6369,N_6035,N_6128);
or U6370 (N_6370,N_6151,N_6201);
and U6371 (N_6371,N_6038,N_6053);
and U6372 (N_6372,N_6195,N_6034);
xnor U6373 (N_6373,N_6032,N_6003);
xor U6374 (N_6374,N_6101,N_6204);
and U6375 (N_6375,N_6066,N_6063);
nor U6376 (N_6376,N_6077,N_6031);
and U6377 (N_6377,N_6134,N_6143);
and U6378 (N_6378,N_6215,N_6237);
nor U6379 (N_6379,N_6048,N_6017);
or U6380 (N_6380,N_6049,N_6204);
nor U6381 (N_6381,N_6010,N_6196);
xnor U6382 (N_6382,N_6033,N_6162);
and U6383 (N_6383,N_6247,N_6190);
or U6384 (N_6384,N_6042,N_6089);
nand U6385 (N_6385,N_6049,N_6006);
nand U6386 (N_6386,N_6036,N_6126);
xnor U6387 (N_6387,N_6132,N_6089);
nor U6388 (N_6388,N_6082,N_6180);
xnor U6389 (N_6389,N_6138,N_6173);
xnor U6390 (N_6390,N_6222,N_6166);
nor U6391 (N_6391,N_6083,N_6124);
nor U6392 (N_6392,N_6113,N_6136);
nand U6393 (N_6393,N_6209,N_6198);
and U6394 (N_6394,N_6010,N_6039);
or U6395 (N_6395,N_6152,N_6025);
nor U6396 (N_6396,N_6135,N_6074);
or U6397 (N_6397,N_6108,N_6190);
and U6398 (N_6398,N_6161,N_6007);
nor U6399 (N_6399,N_6103,N_6008);
nor U6400 (N_6400,N_6061,N_6017);
and U6401 (N_6401,N_6231,N_6051);
xnor U6402 (N_6402,N_6194,N_6146);
or U6403 (N_6403,N_6237,N_6149);
xnor U6404 (N_6404,N_6182,N_6028);
nand U6405 (N_6405,N_6109,N_6153);
xor U6406 (N_6406,N_6141,N_6249);
nor U6407 (N_6407,N_6175,N_6055);
or U6408 (N_6408,N_6217,N_6202);
or U6409 (N_6409,N_6087,N_6129);
nand U6410 (N_6410,N_6112,N_6158);
nor U6411 (N_6411,N_6064,N_6081);
xor U6412 (N_6412,N_6178,N_6245);
and U6413 (N_6413,N_6015,N_6173);
and U6414 (N_6414,N_6198,N_6228);
or U6415 (N_6415,N_6100,N_6249);
nor U6416 (N_6416,N_6056,N_6086);
nor U6417 (N_6417,N_6198,N_6204);
and U6418 (N_6418,N_6079,N_6096);
xnor U6419 (N_6419,N_6176,N_6024);
and U6420 (N_6420,N_6198,N_6238);
or U6421 (N_6421,N_6134,N_6231);
nor U6422 (N_6422,N_6015,N_6213);
nor U6423 (N_6423,N_6027,N_6121);
nor U6424 (N_6424,N_6088,N_6217);
nand U6425 (N_6425,N_6004,N_6028);
nor U6426 (N_6426,N_6069,N_6013);
or U6427 (N_6427,N_6097,N_6244);
nor U6428 (N_6428,N_6232,N_6249);
nor U6429 (N_6429,N_6229,N_6061);
nor U6430 (N_6430,N_6059,N_6145);
xnor U6431 (N_6431,N_6030,N_6138);
xor U6432 (N_6432,N_6102,N_6203);
xor U6433 (N_6433,N_6100,N_6219);
nor U6434 (N_6434,N_6219,N_6093);
nand U6435 (N_6435,N_6059,N_6165);
xor U6436 (N_6436,N_6134,N_6139);
and U6437 (N_6437,N_6238,N_6041);
or U6438 (N_6438,N_6219,N_6240);
and U6439 (N_6439,N_6115,N_6137);
or U6440 (N_6440,N_6100,N_6174);
or U6441 (N_6441,N_6235,N_6012);
nor U6442 (N_6442,N_6054,N_6154);
nor U6443 (N_6443,N_6038,N_6234);
and U6444 (N_6444,N_6011,N_6212);
nand U6445 (N_6445,N_6059,N_6125);
or U6446 (N_6446,N_6221,N_6132);
and U6447 (N_6447,N_6085,N_6222);
and U6448 (N_6448,N_6129,N_6019);
xnor U6449 (N_6449,N_6099,N_6162);
and U6450 (N_6450,N_6218,N_6090);
nand U6451 (N_6451,N_6046,N_6001);
nand U6452 (N_6452,N_6083,N_6145);
and U6453 (N_6453,N_6067,N_6216);
and U6454 (N_6454,N_6158,N_6224);
or U6455 (N_6455,N_6111,N_6180);
nor U6456 (N_6456,N_6076,N_6008);
nand U6457 (N_6457,N_6060,N_6130);
nand U6458 (N_6458,N_6089,N_6162);
or U6459 (N_6459,N_6070,N_6131);
and U6460 (N_6460,N_6133,N_6179);
nand U6461 (N_6461,N_6102,N_6230);
nand U6462 (N_6462,N_6072,N_6103);
nand U6463 (N_6463,N_6050,N_6125);
or U6464 (N_6464,N_6108,N_6034);
nor U6465 (N_6465,N_6124,N_6133);
or U6466 (N_6466,N_6052,N_6071);
and U6467 (N_6467,N_6034,N_6085);
nand U6468 (N_6468,N_6050,N_6143);
nand U6469 (N_6469,N_6010,N_6247);
or U6470 (N_6470,N_6167,N_6022);
and U6471 (N_6471,N_6034,N_6107);
xnor U6472 (N_6472,N_6077,N_6240);
nand U6473 (N_6473,N_6041,N_6216);
xnor U6474 (N_6474,N_6218,N_6140);
or U6475 (N_6475,N_6128,N_6082);
and U6476 (N_6476,N_6231,N_6011);
or U6477 (N_6477,N_6230,N_6031);
or U6478 (N_6478,N_6116,N_6008);
or U6479 (N_6479,N_6068,N_6029);
or U6480 (N_6480,N_6124,N_6137);
nand U6481 (N_6481,N_6049,N_6158);
xnor U6482 (N_6482,N_6154,N_6211);
and U6483 (N_6483,N_6017,N_6195);
xor U6484 (N_6484,N_6104,N_6133);
nand U6485 (N_6485,N_6065,N_6192);
xor U6486 (N_6486,N_6010,N_6055);
nand U6487 (N_6487,N_6035,N_6185);
xor U6488 (N_6488,N_6014,N_6221);
nand U6489 (N_6489,N_6159,N_6117);
nand U6490 (N_6490,N_6013,N_6057);
nor U6491 (N_6491,N_6239,N_6221);
and U6492 (N_6492,N_6032,N_6234);
nand U6493 (N_6493,N_6126,N_6110);
and U6494 (N_6494,N_6187,N_6245);
nor U6495 (N_6495,N_6029,N_6173);
nand U6496 (N_6496,N_6112,N_6228);
and U6497 (N_6497,N_6211,N_6182);
nand U6498 (N_6498,N_6160,N_6241);
xor U6499 (N_6499,N_6230,N_6211);
nor U6500 (N_6500,N_6474,N_6359);
xnor U6501 (N_6501,N_6269,N_6268);
nor U6502 (N_6502,N_6299,N_6366);
xor U6503 (N_6503,N_6451,N_6470);
or U6504 (N_6504,N_6483,N_6342);
nor U6505 (N_6505,N_6309,N_6305);
and U6506 (N_6506,N_6306,N_6307);
and U6507 (N_6507,N_6384,N_6468);
and U6508 (N_6508,N_6399,N_6285);
or U6509 (N_6509,N_6420,N_6490);
nand U6510 (N_6510,N_6389,N_6457);
and U6511 (N_6511,N_6406,N_6370);
nor U6512 (N_6512,N_6337,N_6391);
nor U6513 (N_6513,N_6258,N_6273);
nand U6514 (N_6514,N_6404,N_6375);
xor U6515 (N_6515,N_6486,N_6449);
nand U6516 (N_6516,N_6477,N_6378);
and U6517 (N_6517,N_6435,N_6254);
nor U6518 (N_6518,N_6277,N_6329);
xor U6519 (N_6519,N_6400,N_6379);
or U6520 (N_6520,N_6321,N_6408);
or U6521 (N_6521,N_6283,N_6385);
xor U6522 (N_6522,N_6272,N_6482);
and U6523 (N_6523,N_6421,N_6314);
or U6524 (N_6524,N_6360,N_6495);
nand U6525 (N_6525,N_6434,N_6287);
nand U6526 (N_6526,N_6318,N_6419);
nor U6527 (N_6527,N_6412,N_6438);
xnor U6528 (N_6528,N_6439,N_6363);
xnor U6529 (N_6529,N_6344,N_6349);
nand U6530 (N_6530,N_6266,N_6356);
nand U6531 (N_6531,N_6393,N_6348);
nand U6532 (N_6532,N_6369,N_6403);
or U6533 (N_6533,N_6444,N_6425);
xor U6534 (N_6534,N_6289,N_6373);
and U6535 (N_6535,N_6250,N_6330);
xnor U6536 (N_6536,N_6487,N_6301);
and U6537 (N_6537,N_6261,N_6341);
and U6538 (N_6538,N_6417,N_6323);
or U6539 (N_6539,N_6343,N_6298);
nor U6540 (N_6540,N_6267,N_6331);
and U6541 (N_6541,N_6475,N_6332);
nand U6542 (N_6542,N_6358,N_6294);
xor U6543 (N_6543,N_6405,N_6462);
nor U6544 (N_6544,N_6480,N_6310);
xor U6545 (N_6545,N_6271,N_6265);
and U6546 (N_6546,N_6322,N_6422);
nor U6547 (N_6547,N_6325,N_6448);
and U6548 (N_6548,N_6453,N_6455);
nor U6549 (N_6549,N_6304,N_6276);
nand U6550 (N_6550,N_6368,N_6494);
nor U6551 (N_6551,N_6461,N_6432);
nand U6552 (N_6552,N_6488,N_6395);
nor U6553 (N_6553,N_6251,N_6383);
nand U6554 (N_6554,N_6317,N_6402);
and U6555 (N_6555,N_6396,N_6484);
nand U6556 (N_6556,N_6416,N_6352);
or U6557 (N_6557,N_6498,N_6253);
xor U6558 (N_6558,N_6284,N_6433);
nor U6559 (N_6559,N_6418,N_6442);
nor U6560 (N_6560,N_6320,N_6274);
nand U6561 (N_6561,N_6450,N_6296);
or U6562 (N_6562,N_6472,N_6324);
or U6563 (N_6563,N_6336,N_6374);
xnor U6564 (N_6564,N_6479,N_6460);
and U6565 (N_6565,N_6464,N_6454);
and U6566 (N_6566,N_6259,N_6353);
xnor U6567 (N_6567,N_6312,N_6492);
xnor U6568 (N_6568,N_6456,N_6292);
xor U6569 (N_6569,N_6280,N_6485);
xnor U6570 (N_6570,N_6409,N_6496);
xor U6571 (N_6571,N_6476,N_6387);
nor U6572 (N_6572,N_6365,N_6397);
nand U6573 (N_6573,N_6328,N_6380);
xor U6574 (N_6574,N_6263,N_6364);
xor U6575 (N_6575,N_6413,N_6446);
nand U6576 (N_6576,N_6445,N_6388);
nor U6577 (N_6577,N_6275,N_6361);
nor U6578 (N_6578,N_6255,N_6429);
xor U6579 (N_6579,N_6447,N_6407);
xnor U6580 (N_6580,N_6491,N_6346);
and U6581 (N_6581,N_6436,N_6291);
nand U6582 (N_6582,N_6398,N_6426);
xnor U6583 (N_6583,N_6288,N_6466);
and U6584 (N_6584,N_6308,N_6339);
nor U6585 (N_6585,N_6452,N_6410);
nor U6586 (N_6586,N_6281,N_6345);
nand U6587 (N_6587,N_6286,N_6300);
nor U6588 (N_6588,N_6302,N_6401);
or U6589 (N_6589,N_6430,N_6437);
nand U6590 (N_6590,N_6478,N_6376);
or U6591 (N_6591,N_6252,N_6355);
and U6592 (N_6592,N_6260,N_6351);
nor U6593 (N_6593,N_6390,N_6316);
xnor U6594 (N_6594,N_6414,N_6326);
or U6595 (N_6595,N_6362,N_6279);
and U6596 (N_6596,N_6471,N_6340);
or U6597 (N_6597,N_6411,N_6415);
or U6598 (N_6598,N_6270,N_6311);
and U6599 (N_6599,N_6290,N_6459);
and U6600 (N_6600,N_6473,N_6497);
nand U6601 (N_6601,N_6427,N_6469);
nor U6602 (N_6602,N_6467,N_6338);
nand U6603 (N_6603,N_6335,N_6257);
or U6604 (N_6604,N_6441,N_6443);
or U6605 (N_6605,N_6262,N_6458);
or U6606 (N_6606,N_6313,N_6297);
and U6607 (N_6607,N_6256,N_6303);
or U6608 (N_6608,N_6481,N_6367);
xnor U6609 (N_6609,N_6489,N_6382);
and U6610 (N_6610,N_6428,N_6293);
xor U6611 (N_6611,N_6392,N_6394);
xnor U6612 (N_6612,N_6278,N_6499);
nor U6613 (N_6613,N_6465,N_6423);
xnor U6614 (N_6614,N_6350,N_6327);
and U6615 (N_6615,N_6354,N_6371);
or U6616 (N_6616,N_6333,N_6377);
nor U6617 (N_6617,N_6381,N_6372);
nand U6618 (N_6618,N_6463,N_6493);
nor U6619 (N_6619,N_6424,N_6440);
nor U6620 (N_6620,N_6347,N_6334);
xnor U6621 (N_6621,N_6431,N_6315);
and U6622 (N_6622,N_6282,N_6264);
and U6623 (N_6623,N_6295,N_6357);
xnor U6624 (N_6624,N_6319,N_6386);
nor U6625 (N_6625,N_6327,N_6417);
xnor U6626 (N_6626,N_6270,N_6453);
nor U6627 (N_6627,N_6479,N_6491);
nor U6628 (N_6628,N_6428,N_6481);
or U6629 (N_6629,N_6310,N_6442);
and U6630 (N_6630,N_6482,N_6448);
nand U6631 (N_6631,N_6325,N_6417);
nor U6632 (N_6632,N_6321,N_6342);
nor U6633 (N_6633,N_6267,N_6376);
or U6634 (N_6634,N_6252,N_6380);
xor U6635 (N_6635,N_6305,N_6388);
xnor U6636 (N_6636,N_6336,N_6376);
nor U6637 (N_6637,N_6483,N_6369);
nand U6638 (N_6638,N_6394,N_6265);
nand U6639 (N_6639,N_6482,N_6389);
xnor U6640 (N_6640,N_6456,N_6490);
nor U6641 (N_6641,N_6284,N_6270);
xor U6642 (N_6642,N_6389,N_6315);
nor U6643 (N_6643,N_6387,N_6437);
and U6644 (N_6644,N_6441,N_6425);
nor U6645 (N_6645,N_6428,N_6251);
nor U6646 (N_6646,N_6277,N_6311);
or U6647 (N_6647,N_6478,N_6286);
or U6648 (N_6648,N_6393,N_6457);
or U6649 (N_6649,N_6469,N_6354);
and U6650 (N_6650,N_6429,N_6335);
and U6651 (N_6651,N_6380,N_6498);
xnor U6652 (N_6652,N_6466,N_6472);
xnor U6653 (N_6653,N_6357,N_6386);
and U6654 (N_6654,N_6286,N_6450);
and U6655 (N_6655,N_6317,N_6342);
and U6656 (N_6656,N_6274,N_6477);
nor U6657 (N_6657,N_6482,N_6352);
nor U6658 (N_6658,N_6420,N_6435);
nand U6659 (N_6659,N_6338,N_6420);
or U6660 (N_6660,N_6337,N_6417);
nor U6661 (N_6661,N_6255,N_6298);
xnor U6662 (N_6662,N_6367,N_6343);
nor U6663 (N_6663,N_6459,N_6434);
or U6664 (N_6664,N_6411,N_6251);
and U6665 (N_6665,N_6455,N_6482);
nand U6666 (N_6666,N_6478,N_6416);
xnor U6667 (N_6667,N_6420,N_6323);
xor U6668 (N_6668,N_6425,N_6341);
xnor U6669 (N_6669,N_6355,N_6445);
nand U6670 (N_6670,N_6478,N_6331);
and U6671 (N_6671,N_6262,N_6444);
xnor U6672 (N_6672,N_6300,N_6393);
nand U6673 (N_6673,N_6354,N_6331);
or U6674 (N_6674,N_6369,N_6450);
or U6675 (N_6675,N_6278,N_6428);
nand U6676 (N_6676,N_6284,N_6419);
xor U6677 (N_6677,N_6285,N_6280);
nand U6678 (N_6678,N_6382,N_6386);
xnor U6679 (N_6679,N_6404,N_6477);
and U6680 (N_6680,N_6348,N_6342);
nor U6681 (N_6681,N_6323,N_6358);
nor U6682 (N_6682,N_6280,N_6275);
nand U6683 (N_6683,N_6478,N_6441);
and U6684 (N_6684,N_6426,N_6364);
or U6685 (N_6685,N_6480,N_6349);
nand U6686 (N_6686,N_6476,N_6496);
or U6687 (N_6687,N_6296,N_6387);
xor U6688 (N_6688,N_6474,N_6454);
or U6689 (N_6689,N_6363,N_6279);
nand U6690 (N_6690,N_6489,N_6418);
or U6691 (N_6691,N_6329,N_6431);
nand U6692 (N_6692,N_6409,N_6455);
and U6693 (N_6693,N_6457,N_6352);
nand U6694 (N_6694,N_6360,N_6373);
and U6695 (N_6695,N_6388,N_6322);
or U6696 (N_6696,N_6426,N_6465);
and U6697 (N_6697,N_6266,N_6403);
or U6698 (N_6698,N_6373,N_6305);
or U6699 (N_6699,N_6390,N_6306);
and U6700 (N_6700,N_6302,N_6373);
nor U6701 (N_6701,N_6297,N_6437);
and U6702 (N_6702,N_6432,N_6264);
nor U6703 (N_6703,N_6432,N_6308);
xor U6704 (N_6704,N_6435,N_6380);
nand U6705 (N_6705,N_6348,N_6487);
nand U6706 (N_6706,N_6303,N_6395);
and U6707 (N_6707,N_6346,N_6381);
nor U6708 (N_6708,N_6421,N_6463);
xor U6709 (N_6709,N_6496,N_6325);
xor U6710 (N_6710,N_6332,N_6391);
or U6711 (N_6711,N_6271,N_6348);
nor U6712 (N_6712,N_6296,N_6452);
and U6713 (N_6713,N_6310,N_6272);
xnor U6714 (N_6714,N_6320,N_6389);
and U6715 (N_6715,N_6480,N_6447);
xnor U6716 (N_6716,N_6274,N_6485);
nand U6717 (N_6717,N_6404,N_6320);
or U6718 (N_6718,N_6365,N_6264);
nor U6719 (N_6719,N_6345,N_6318);
nor U6720 (N_6720,N_6459,N_6314);
nand U6721 (N_6721,N_6317,N_6269);
xnor U6722 (N_6722,N_6454,N_6484);
nand U6723 (N_6723,N_6483,N_6293);
nand U6724 (N_6724,N_6314,N_6388);
nor U6725 (N_6725,N_6394,N_6332);
or U6726 (N_6726,N_6414,N_6402);
xor U6727 (N_6727,N_6493,N_6375);
and U6728 (N_6728,N_6363,N_6299);
and U6729 (N_6729,N_6313,N_6353);
or U6730 (N_6730,N_6306,N_6343);
xnor U6731 (N_6731,N_6324,N_6432);
xnor U6732 (N_6732,N_6271,N_6276);
nor U6733 (N_6733,N_6375,N_6251);
or U6734 (N_6734,N_6417,N_6352);
and U6735 (N_6735,N_6329,N_6402);
nand U6736 (N_6736,N_6373,N_6295);
or U6737 (N_6737,N_6373,N_6276);
or U6738 (N_6738,N_6250,N_6473);
xor U6739 (N_6739,N_6317,N_6417);
and U6740 (N_6740,N_6280,N_6416);
xor U6741 (N_6741,N_6255,N_6438);
and U6742 (N_6742,N_6348,N_6460);
and U6743 (N_6743,N_6296,N_6341);
or U6744 (N_6744,N_6409,N_6357);
nand U6745 (N_6745,N_6352,N_6303);
xnor U6746 (N_6746,N_6307,N_6400);
xnor U6747 (N_6747,N_6356,N_6378);
or U6748 (N_6748,N_6352,N_6445);
nor U6749 (N_6749,N_6480,N_6498);
nor U6750 (N_6750,N_6705,N_6634);
or U6751 (N_6751,N_6571,N_6578);
nand U6752 (N_6752,N_6548,N_6504);
nand U6753 (N_6753,N_6597,N_6741);
xor U6754 (N_6754,N_6722,N_6606);
nor U6755 (N_6755,N_6556,N_6586);
nor U6756 (N_6756,N_6622,N_6584);
xor U6757 (N_6757,N_6544,N_6538);
nand U6758 (N_6758,N_6518,N_6532);
nor U6759 (N_6759,N_6585,N_6537);
and U6760 (N_6760,N_6596,N_6662);
nor U6761 (N_6761,N_6656,N_6620);
nand U6762 (N_6762,N_6539,N_6575);
nand U6763 (N_6763,N_6646,N_6581);
or U6764 (N_6764,N_6643,N_6639);
and U6765 (N_6765,N_6615,N_6589);
nand U6766 (N_6766,N_6691,N_6627);
nor U6767 (N_6767,N_6654,N_6702);
xnor U6768 (N_6768,N_6683,N_6524);
nand U6769 (N_6769,N_6647,N_6587);
nand U6770 (N_6770,N_6680,N_6673);
nand U6771 (N_6771,N_6607,N_6531);
xor U6772 (N_6772,N_6605,N_6667);
xnor U6773 (N_6773,N_6614,N_6602);
or U6774 (N_6774,N_6633,N_6552);
nand U6775 (N_6775,N_6540,N_6649);
nor U6776 (N_6776,N_6714,N_6671);
xnor U6777 (N_6777,N_6593,N_6618);
or U6778 (N_6778,N_6645,N_6572);
xor U6779 (N_6779,N_6557,N_6583);
nand U6780 (N_6780,N_6612,N_6638);
nor U6781 (N_6781,N_6555,N_6574);
nand U6782 (N_6782,N_6545,N_6536);
nand U6783 (N_6783,N_6610,N_6547);
and U6784 (N_6784,N_6500,N_6511);
xnor U6785 (N_6785,N_6554,N_6632);
and U6786 (N_6786,N_6515,N_6648);
nor U6787 (N_6787,N_6650,N_6601);
and U6788 (N_6788,N_6735,N_6655);
or U6789 (N_6789,N_6663,N_6718);
or U6790 (N_6790,N_6668,N_6579);
xnor U6791 (N_6791,N_6630,N_6534);
nor U6792 (N_6792,N_6651,N_6727);
xor U6793 (N_6793,N_6566,N_6682);
nand U6794 (N_6794,N_6636,N_6708);
and U6795 (N_6795,N_6559,N_6679);
and U6796 (N_6796,N_6635,N_6652);
xor U6797 (N_6797,N_6528,N_6573);
and U6798 (N_6798,N_6600,N_6724);
nor U6799 (N_6799,N_6717,N_6512);
nor U6800 (N_6800,N_6734,N_6603);
nand U6801 (N_6801,N_6563,N_6693);
xor U6802 (N_6802,N_6725,N_6553);
or U6803 (N_6803,N_6505,N_6733);
nor U6804 (N_6804,N_6526,N_6700);
nand U6805 (N_6805,N_6677,N_6684);
nor U6806 (N_6806,N_6501,N_6590);
or U6807 (N_6807,N_6529,N_6608);
or U6808 (N_6808,N_6506,N_6522);
or U6809 (N_6809,N_6523,N_6748);
or U6810 (N_6810,N_6686,N_6619);
or U6811 (N_6811,N_6582,N_6591);
and U6812 (N_6812,N_6687,N_6669);
xor U6813 (N_6813,N_6688,N_6704);
and U6814 (N_6814,N_6565,N_6517);
xor U6815 (N_6815,N_6699,N_6685);
or U6816 (N_6816,N_6541,N_6509);
nor U6817 (N_6817,N_6569,N_6550);
nand U6818 (N_6818,N_6535,N_6670);
or U6819 (N_6819,N_6576,N_6570);
and U6820 (N_6820,N_6599,N_6743);
nor U6821 (N_6821,N_6613,N_6661);
nor U6822 (N_6822,N_6623,N_6562);
nand U6823 (N_6823,N_6624,N_6527);
nor U6824 (N_6824,N_6715,N_6660);
nor U6825 (N_6825,N_6697,N_6598);
or U6826 (N_6826,N_6672,N_6592);
and U6827 (N_6827,N_6696,N_6626);
nor U6828 (N_6828,N_6510,N_6629);
and U6829 (N_6829,N_6701,N_6561);
nor U6830 (N_6830,N_6525,N_6681);
nor U6831 (N_6831,N_6674,N_6703);
nand U6832 (N_6832,N_6723,N_6716);
nor U6833 (N_6833,N_6665,N_6551);
or U6834 (N_6834,N_6709,N_6549);
nand U6835 (N_6835,N_6644,N_6503);
or U6836 (N_6836,N_6710,N_6625);
nand U6837 (N_6837,N_6731,N_6664);
xor U6838 (N_6838,N_6580,N_6659);
and U6839 (N_6839,N_6519,N_6508);
nand U6840 (N_6840,N_6631,N_6745);
and U6841 (N_6841,N_6533,N_6543);
nand U6842 (N_6842,N_6558,N_6595);
nor U6843 (N_6843,N_6694,N_6737);
xor U6844 (N_6844,N_6711,N_6692);
and U6845 (N_6845,N_6564,N_6719);
xor U6846 (N_6846,N_6726,N_6747);
nor U6847 (N_6847,N_6642,N_6713);
xor U6848 (N_6848,N_6730,N_6628);
nor U6849 (N_6849,N_6617,N_6738);
or U6850 (N_6850,N_6740,N_6749);
nor U6851 (N_6851,N_6502,N_6616);
or U6852 (N_6852,N_6530,N_6577);
nor U6853 (N_6853,N_6640,N_6594);
nand U6854 (N_6854,N_6729,N_6588);
nand U6855 (N_6855,N_6678,N_6721);
nor U6856 (N_6856,N_6604,N_6611);
xor U6857 (N_6857,N_6712,N_6567);
nor U6858 (N_6858,N_6689,N_6676);
nand U6859 (N_6859,N_6653,N_6513);
nand U6860 (N_6860,N_6657,N_6746);
nor U6861 (N_6861,N_6516,N_6720);
or U6862 (N_6862,N_6514,N_6521);
nor U6863 (N_6863,N_6706,N_6560);
nor U6864 (N_6864,N_6658,N_6621);
xnor U6865 (N_6865,N_6507,N_6641);
xor U6866 (N_6866,N_6568,N_6520);
xnor U6867 (N_6867,N_6698,N_6739);
and U6868 (N_6868,N_6728,N_6542);
and U6869 (N_6869,N_6666,N_6695);
nor U6870 (N_6870,N_6546,N_6736);
nand U6871 (N_6871,N_6690,N_6742);
and U6872 (N_6872,N_6637,N_6744);
nand U6873 (N_6873,N_6707,N_6609);
nand U6874 (N_6874,N_6675,N_6732);
xor U6875 (N_6875,N_6679,N_6706);
and U6876 (N_6876,N_6579,N_6607);
or U6877 (N_6877,N_6518,N_6710);
nand U6878 (N_6878,N_6541,N_6607);
or U6879 (N_6879,N_6563,N_6682);
or U6880 (N_6880,N_6649,N_6598);
and U6881 (N_6881,N_6723,N_6748);
nand U6882 (N_6882,N_6640,N_6722);
nand U6883 (N_6883,N_6611,N_6610);
xor U6884 (N_6884,N_6747,N_6583);
nor U6885 (N_6885,N_6527,N_6540);
xnor U6886 (N_6886,N_6591,N_6502);
nand U6887 (N_6887,N_6529,N_6735);
nand U6888 (N_6888,N_6749,N_6559);
or U6889 (N_6889,N_6623,N_6609);
nand U6890 (N_6890,N_6549,N_6569);
or U6891 (N_6891,N_6566,N_6536);
or U6892 (N_6892,N_6643,N_6584);
or U6893 (N_6893,N_6606,N_6590);
and U6894 (N_6894,N_6748,N_6630);
or U6895 (N_6895,N_6648,N_6615);
nand U6896 (N_6896,N_6737,N_6624);
and U6897 (N_6897,N_6550,N_6607);
or U6898 (N_6898,N_6663,N_6503);
or U6899 (N_6899,N_6731,N_6658);
nor U6900 (N_6900,N_6558,N_6555);
or U6901 (N_6901,N_6681,N_6560);
nand U6902 (N_6902,N_6649,N_6729);
nand U6903 (N_6903,N_6678,N_6734);
or U6904 (N_6904,N_6541,N_6537);
xnor U6905 (N_6905,N_6648,N_6717);
xor U6906 (N_6906,N_6594,N_6722);
nor U6907 (N_6907,N_6718,N_6694);
or U6908 (N_6908,N_6618,N_6704);
nor U6909 (N_6909,N_6708,N_6513);
or U6910 (N_6910,N_6627,N_6708);
and U6911 (N_6911,N_6598,N_6504);
or U6912 (N_6912,N_6684,N_6655);
and U6913 (N_6913,N_6571,N_6574);
xor U6914 (N_6914,N_6560,N_6692);
nor U6915 (N_6915,N_6677,N_6668);
nor U6916 (N_6916,N_6592,N_6720);
nand U6917 (N_6917,N_6698,N_6692);
xor U6918 (N_6918,N_6637,N_6732);
or U6919 (N_6919,N_6504,N_6735);
and U6920 (N_6920,N_6502,N_6578);
xor U6921 (N_6921,N_6586,N_6502);
nand U6922 (N_6922,N_6558,N_6718);
or U6923 (N_6923,N_6585,N_6629);
xor U6924 (N_6924,N_6541,N_6639);
nor U6925 (N_6925,N_6658,N_6515);
and U6926 (N_6926,N_6605,N_6684);
or U6927 (N_6927,N_6651,N_6517);
nand U6928 (N_6928,N_6678,N_6634);
nand U6929 (N_6929,N_6731,N_6631);
nor U6930 (N_6930,N_6622,N_6697);
or U6931 (N_6931,N_6516,N_6653);
nor U6932 (N_6932,N_6636,N_6589);
nor U6933 (N_6933,N_6579,N_6613);
xnor U6934 (N_6934,N_6708,N_6506);
and U6935 (N_6935,N_6570,N_6535);
xor U6936 (N_6936,N_6537,N_6611);
and U6937 (N_6937,N_6627,N_6503);
xnor U6938 (N_6938,N_6646,N_6510);
xor U6939 (N_6939,N_6572,N_6632);
nand U6940 (N_6940,N_6710,N_6551);
nand U6941 (N_6941,N_6534,N_6523);
or U6942 (N_6942,N_6683,N_6694);
or U6943 (N_6943,N_6686,N_6572);
or U6944 (N_6944,N_6527,N_6531);
nor U6945 (N_6945,N_6629,N_6662);
and U6946 (N_6946,N_6578,N_6707);
nor U6947 (N_6947,N_6521,N_6572);
or U6948 (N_6948,N_6644,N_6690);
or U6949 (N_6949,N_6647,N_6506);
or U6950 (N_6950,N_6698,N_6691);
and U6951 (N_6951,N_6615,N_6624);
nand U6952 (N_6952,N_6606,N_6596);
nor U6953 (N_6953,N_6660,N_6699);
and U6954 (N_6954,N_6741,N_6567);
nand U6955 (N_6955,N_6515,N_6611);
nand U6956 (N_6956,N_6711,N_6548);
and U6957 (N_6957,N_6523,N_6744);
xor U6958 (N_6958,N_6714,N_6527);
nand U6959 (N_6959,N_6699,N_6567);
xor U6960 (N_6960,N_6666,N_6508);
or U6961 (N_6961,N_6726,N_6722);
or U6962 (N_6962,N_6582,N_6568);
and U6963 (N_6963,N_6715,N_6695);
nor U6964 (N_6964,N_6501,N_6656);
or U6965 (N_6965,N_6530,N_6725);
and U6966 (N_6966,N_6654,N_6625);
xnor U6967 (N_6967,N_6586,N_6671);
nor U6968 (N_6968,N_6711,N_6667);
nand U6969 (N_6969,N_6749,N_6709);
or U6970 (N_6970,N_6523,N_6569);
or U6971 (N_6971,N_6679,N_6606);
xnor U6972 (N_6972,N_6644,N_6573);
nand U6973 (N_6973,N_6568,N_6740);
or U6974 (N_6974,N_6581,N_6622);
and U6975 (N_6975,N_6681,N_6537);
nor U6976 (N_6976,N_6739,N_6608);
nor U6977 (N_6977,N_6518,N_6576);
nor U6978 (N_6978,N_6543,N_6621);
xnor U6979 (N_6979,N_6657,N_6576);
nand U6980 (N_6980,N_6661,N_6627);
nor U6981 (N_6981,N_6692,N_6559);
xor U6982 (N_6982,N_6719,N_6607);
and U6983 (N_6983,N_6594,N_6510);
nor U6984 (N_6984,N_6601,N_6675);
nor U6985 (N_6985,N_6651,N_6697);
and U6986 (N_6986,N_6674,N_6746);
or U6987 (N_6987,N_6695,N_6673);
nor U6988 (N_6988,N_6614,N_6633);
or U6989 (N_6989,N_6711,N_6682);
nor U6990 (N_6990,N_6721,N_6555);
nand U6991 (N_6991,N_6626,N_6738);
nor U6992 (N_6992,N_6624,N_6594);
and U6993 (N_6993,N_6579,N_6530);
nor U6994 (N_6994,N_6575,N_6535);
nand U6995 (N_6995,N_6549,N_6658);
or U6996 (N_6996,N_6534,N_6642);
and U6997 (N_6997,N_6529,N_6671);
and U6998 (N_6998,N_6645,N_6506);
xnor U6999 (N_6999,N_6737,N_6617);
and U7000 (N_7000,N_6771,N_6940);
nor U7001 (N_7001,N_6807,N_6942);
nor U7002 (N_7002,N_6835,N_6890);
and U7003 (N_7003,N_6785,N_6880);
and U7004 (N_7004,N_6983,N_6897);
nand U7005 (N_7005,N_6887,N_6946);
xor U7006 (N_7006,N_6795,N_6803);
nand U7007 (N_7007,N_6924,N_6957);
and U7008 (N_7008,N_6896,N_6846);
nor U7009 (N_7009,N_6776,N_6796);
or U7010 (N_7010,N_6826,N_6763);
xnor U7011 (N_7011,N_6865,N_6971);
or U7012 (N_7012,N_6994,N_6939);
and U7013 (N_7013,N_6847,N_6851);
and U7014 (N_7014,N_6870,N_6884);
nand U7015 (N_7015,N_6817,N_6808);
xor U7016 (N_7016,N_6872,N_6955);
or U7017 (N_7017,N_6819,N_6873);
and U7018 (N_7018,N_6829,N_6798);
or U7019 (N_7019,N_6898,N_6838);
nand U7020 (N_7020,N_6828,N_6977);
nor U7021 (N_7021,N_6961,N_6783);
xnor U7022 (N_7022,N_6750,N_6938);
xnor U7023 (N_7023,N_6913,N_6877);
nor U7024 (N_7024,N_6858,N_6911);
and U7025 (N_7025,N_6947,N_6929);
nor U7026 (N_7026,N_6906,N_6967);
and U7027 (N_7027,N_6864,N_6770);
and U7028 (N_7028,N_6844,N_6821);
or U7029 (N_7029,N_6909,N_6927);
and U7030 (N_7030,N_6781,N_6894);
and U7031 (N_7031,N_6892,N_6822);
nand U7032 (N_7032,N_6901,N_6797);
nand U7033 (N_7033,N_6958,N_6790);
nor U7034 (N_7034,N_6834,N_6928);
nand U7035 (N_7035,N_6916,N_6923);
xnor U7036 (N_7036,N_6816,N_6786);
xnor U7037 (N_7037,N_6792,N_6879);
nand U7038 (N_7038,N_6841,N_6799);
or U7039 (N_7039,N_6878,N_6886);
nor U7040 (N_7040,N_6905,N_6926);
nor U7041 (N_7041,N_6860,N_6862);
xnor U7042 (N_7042,N_6809,N_6996);
xnor U7043 (N_7043,N_6831,N_6768);
and U7044 (N_7044,N_6780,N_6973);
and U7045 (N_7045,N_6999,N_6866);
nor U7046 (N_7046,N_6964,N_6986);
nand U7047 (N_7047,N_6793,N_6988);
nand U7048 (N_7048,N_6843,N_6992);
nor U7049 (N_7049,N_6993,N_6981);
nor U7050 (N_7050,N_6766,N_6899);
xnor U7051 (N_7051,N_6757,N_6802);
xor U7052 (N_7052,N_6871,N_6850);
nand U7053 (N_7053,N_6908,N_6918);
and U7054 (N_7054,N_6760,N_6811);
and U7055 (N_7055,N_6775,N_6839);
nor U7056 (N_7056,N_6920,N_6932);
nor U7057 (N_7057,N_6982,N_6936);
nor U7058 (N_7058,N_6985,N_6893);
nor U7059 (N_7059,N_6900,N_6840);
or U7060 (N_7060,N_6969,N_6823);
and U7061 (N_7061,N_6980,N_6922);
xnor U7062 (N_7062,N_6904,N_6945);
nand U7063 (N_7063,N_6959,N_6812);
and U7064 (N_7064,N_6842,N_6800);
nor U7065 (N_7065,N_6997,N_6859);
xnor U7066 (N_7066,N_6806,N_6875);
and U7067 (N_7067,N_6794,N_6810);
and U7068 (N_7068,N_6934,N_6805);
or U7069 (N_7069,N_6990,N_6944);
xor U7070 (N_7070,N_6857,N_6869);
xnor U7071 (N_7071,N_6965,N_6933);
nand U7072 (N_7072,N_6949,N_6998);
nand U7073 (N_7073,N_6778,N_6820);
and U7074 (N_7074,N_6902,N_6813);
and U7075 (N_7075,N_6975,N_6772);
nand U7076 (N_7076,N_6852,N_6764);
and U7077 (N_7077,N_6948,N_6951);
xnor U7078 (N_7078,N_6925,N_6848);
xnor U7079 (N_7079,N_6836,N_6950);
nand U7080 (N_7080,N_6931,N_6941);
nor U7081 (N_7081,N_6814,N_6773);
nand U7082 (N_7082,N_6789,N_6854);
xnor U7083 (N_7083,N_6943,N_6968);
xnor U7084 (N_7084,N_6930,N_6788);
xnor U7085 (N_7085,N_6818,N_6978);
xnor U7086 (N_7086,N_6759,N_6849);
xor U7087 (N_7087,N_6921,N_6863);
nor U7088 (N_7088,N_6991,N_6758);
nor U7089 (N_7089,N_6974,N_6882);
and U7090 (N_7090,N_6876,N_6867);
nor U7091 (N_7091,N_6755,N_6856);
nor U7092 (N_7092,N_6861,N_6787);
nor U7093 (N_7093,N_6966,N_6791);
and U7094 (N_7094,N_6976,N_6889);
or U7095 (N_7095,N_6804,N_6824);
or U7096 (N_7096,N_6917,N_6995);
xnor U7097 (N_7097,N_6832,N_6855);
and U7098 (N_7098,N_6753,N_6774);
nor U7099 (N_7099,N_6914,N_6912);
or U7100 (N_7100,N_6762,N_6972);
xor U7101 (N_7101,N_6767,N_6765);
nand U7102 (N_7102,N_6874,N_6782);
nand U7103 (N_7103,N_6888,N_6779);
xnor U7104 (N_7104,N_6987,N_6881);
xnor U7105 (N_7105,N_6907,N_6751);
xnor U7106 (N_7106,N_6895,N_6937);
or U7107 (N_7107,N_6935,N_6885);
nand U7108 (N_7108,N_6954,N_6956);
xor U7109 (N_7109,N_6784,N_6761);
nor U7110 (N_7110,N_6827,N_6845);
or U7111 (N_7111,N_6801,N_6853);
xor U7112 (N_7112,N_6970,N_6769);
nor U7113 (N_7113,N_6756,N_6979);
xnor U7114 (N_7114,N_6962,N_6915);
xor U7115 (N_7115,N_6883,N_6891);
and U7116 (N_7116,N_6868,N_6989);
xor U7117 (N_7117,N_6910,N_6837);
nand U7118 (N_7118,N_6903,N_6960);
or U7119 (N_7119,N_6777,N_6752);
xnor U7120 (N_7120,N_6984,N_6833);
nand U7121 (N_7121,N_6919,N_6825);
or U7122 (N_7122,N_6963,N_6830);
and U7123 (N_7123,N_6952,N_6754);
or U7124 (N_7124,N_6815,N_6953);
nand U7125 (N_7125,N_6960,N_6837);
nor U7126 (N_7126,N_6845,N_6788);
nand U7127 (N_7127,N_6865,N_6937);
or U7128 (N_7128,N_6757,N_6779);
and U7129 (N_7129,N_6972,N_6774);
nor U7130 (N_7130,N_6935,N_6939);
nor U7131 (N_7131,N_6910,N_6811);
and U7132 (N_7132,N_6953,N_6948);
and U7133 (N_7133,N_6904,N_6870);
nor U7134 (N_7134,N_6784,N_6966);
nand U7135 (N_7135,N_6859,N_6954);
and U7136 (N_7136,N_6816,N_6965);
xnor U7137 (N_7137,N_6956,N_6998);
or U7138 (N_7138,N_6834,N_6885);
nor U7139 (N_7139,N_6875,N_6883);
and U7140 (N_7140,N_6956,N_6986);
xnor U7141 (N_7141,N_6981,N_6959);
xor U7142 (N_7142,N_6888,N_6802);
xnor U7143 (N_7143,N_6774,N_6865);
and U7144 (N_7144,N_6806,N_6790);
or U7145 (N_7145,N_6750,N_6929);
xnor U7146 (N_7146,N_6789,N_6889);
or U7147 (N_7147,N_6776,N_6982);
and U7148 (N_7148,N_6915,N_6863);
nor U7149 (N_7149,N_6887,N_6779);
and U7150 (N_7150,N_6842,N_6971);
or U7151 (N_7151,N_6972,N_6965);
and U7152 (N_7152,N_6916,N_6917);
and U7153 (N_7153,N_6876,N_6956);
and U7154 (N_7154,N_6824,N_6759);
xor U7155 (N_7155,N_6778,N_6775);
nand U7156 (N_7156,N_6958,N_6898);
xnor U7157 (N_7157,N_6909,N_6892);
and U7158 (N_7158,N_6954,N_6863);
and U7159 (N_7159,N_6791,N_6771);
nand U7160 (N_7160,N_6804,N_6772);
nor U7161 (N_7161,N_6903,N_6885);
nor U7162 (N_7162,N_6910,N_6826);
nand U7163 (N_7163,N_6800,N_6912);
nand U7164 (N_7164,N_6812,N_6872);
and U7165 (N_7165,N_6810,N_6909);
and U7166 (N_7166,N_6765,N_6878);
nand U7167 (N_7167,N_6889,N_6982);
or U7168 (N_7168,N_6990,N_6986);
nor U7169 (N_7169,N_6836,N_6807);
and U7170 (N_7170,N_6777,N_6803);
and U7171 (N_7171,N_6901,N_6850);
nand U7172 (N_7172,N_6896,N_6759);
and U7173 (N_7173,N_6907,N_6821);
or U7174 (N_7174,N_6848,N_6980);
or U7175 (N_7175,N_6872,N_6795);
nor U7176 (N_7176,N_6899,N_6860);
and U7177 (N_7177,N_6930,N_6848);
nor U7178 (N_7178,N_6937,N_6799);
and U7179 (N_7179,N_6905,N_6891);
or U7180 (N_7180,N_6762,N_6920);
and U7181 (N_7181,N_6817,N_6907);
or U7182 (N_7182,N_6945,N_6931);
nor U7183 (N_7183,N_6816,N_6814);
and U7184 (N_7184,N_6834,N_6984);
or U7185 (N_7185,N_6993,N_6899);
and U7186 (N_7186,N_6847,N_6907);
nand U7187 (N_7187,N_6815,N_6897);
nor U7188 (N_7188,N_6904,N_6777);
or U7189 (N_7189,N_6796,N_6938);
and U7190 (N_7190,N_6798,N_6826);
nand U7191 (N_7191,N_6851,N_6861);
or U7192 (N_7192,N_6959,N_6790);
nor U7193 (N_7193,N_6966,N_6968);
nand U7194 (N_7194,N_6850,N_6817);
or U7195 (N_7195,N_6869,N_6942);
nand U7196 (N_7196,N_6795,N_6756);
nand U7197 (N_7197,N_6944,N_6843);
or U7198 (N_7198,N_6840,N_6858);
and U7199 (N_7199,N_6945,N_6955);
or U7200 (N_7200,N_6849,N_6831);
xor U7201 (N_7201,N_6870,N_6783);
or U7202 (N_7202,N_6926,N_6776);
nor U7203 (N_7203,N_6994,N_6775);
or U7204 (N_7204,N_6875,N_6831);
nor U7205 (N_7205,N_6770,N_6971);
or U7206 (N_7206,N_6786,N_6798);
nor U7207 (N_7207,N_6790,N_6774);
nor U7208 (N_7208,N_6815,N_6836);
or U7209 (N_7209,N_6825,N_6970);
xnor U7210 (N_7210,N_6915,N_6859);
or U7211 (N_7211,N_6881,N_6957);
or U7212 (N_7212,N_6767,N_6950);
nand U7213 (N_7213,N_6890,N_6985);
or U7214 (N_7214,N_6831,N_6903);
xor U7215 (N_7215,N_6814,N_6917);
xor U7216 (N_7216,N_6846,N_6833);
or U7217 (N_7217,N_6879,N_6915);
and U7218 (N_7218,N_6855,N_6753);
nor U7219 (N_7219,N_6815,N_6839);
nand U7220 (N_7220,N_6797,N_6818);
or U7221 (N_7221,N_6808,N_6818);
xnor U7222 (N_7222,N_6934,N_6816);
or U7223 (N_7223,N_6910,N_6981);
nand U7224 (N_7224,N_6757,N_6950);
xor U7225 (N_7225,N_6909,N_6966);
nor U7226 (N_7226,N_6952,N_6954);
nor U7227 (N_7227,N_6823,N_6816);
xnor U7228 (N_7228,N_6834,N_6764);
nor U7229 (N_7229,N_6859,N_6849);
nand U7230 (N_7230,N_6881,N_6767);
nor U7231 (N_7231,N_6994,N_6865);
and U7232 (N_7232,N_6886,N_6911);
nor U7233 (N_7233,N_6770,N_6995);
nand U7234 (N_7234,N_6838,N_6887);
xor U7235 (N_7235,N_6985,N_6950);
nor U7236 (N_7236,N_6798,N_6888);
xor U7237 (N_7237,N_6764,N_6775);
nand U7238 (N_7238,N_6877,N_6815);
nor U7239 (N_7239,N_6794,N_6966);
nand U7240 (N_7240,N_6867,N_6997);
or U7241 (N_7241,N_6847,N_6777);
nor U7242 (N_7242,N_6878,N_6984);
and U7243 (N_7243,N_6813,N_6948);
or U7244 (N_7244,N_6966,N_6904);
nand U7245 (N_7245,N_6960,N_6867);
nand U7246 (N_7246,N_6892,N_6761);
nand U7247 (N_7247,N_6984,N_6761);
nor U7248 (N_7248,N_6955,N_6905);
and U7249 (N_7249,N_6766,N_6832);
and U7250 (N_7250,N_7130,N_7203);
nand U7251 (N_7251,N_7072,N_7231);
and U7252 (N_7252,N_7189,N_7078);
and U7253 (N_7253,N_7191,N_7234);
and U7254 (N_7254,N_7031,N_7131);
xnor U7255 (N_7255,N_7220,N_7059);
nand U7256 (N_7256,N_7071,N_7018);
nor U7257 (N_7257,N_7110,N_7023);
nand U7258 (N_7258,N_7000,N_7217);
xor U7259 (N_7259,N_7202,N_7222);
and U7260 (N_7260,N_7032,N_7162);
xnor U7261 (N_7261,N_7185,N_7027);
nor U7262 (N_7262,N_7080,N_7103);
nand U7263 (N_7263,N_7124,N_7054);
xnor U7264 (N_7264,N_7092,N_7063);
nor U7265 (N_7265,N_7028,N_7168);
or U7266 (N_7266,N_7020,N_7187);
xor U7267 (N_7267,N_7226,N_7004);
and U7268 (N_7268,N_7184,N_7154);
and U7269 (N_7269,N_7113,N_7219);
nand U7270 (N_7270,N_7160,N_7003);
nor U7271 (N_7271,N_7206,N_7157);
xnor U7272 (N_7272,N_7211,N_7169);
xor U7273 (N_7273,N_7045,N_7002);
or U7274 (N_7274,N_7239,N_7114);
or U7275 (N_7275,N_7141,N_7161);
and U7276 (N_7276,N_7170,N_7196);
or U7277 (N_7277,N_7042,N_7193);
xnor U7278 (N_7278,N_7188,N_7121);
nand U7279 (N_7279,N_7177,N_7145);
or U7280 (N_7280,N_7129,N_7224);
nand U7281 (N_7281,N_7104,N_7225);
and U7282 (N_7282,N_7052,N_7127);
xnor U7283 (N_7283,N_7182,N_7136);
nor U7284 (N_7284,N_7172,N_7164);
nor U7285 (N_7285,N_7134,N_7137);
nor U7286 (N_7286,N_7039,N_7019);
nor U7287 (N_7287,N_7135,N_7246);
or U7288 (N_7288,N_7171,N_7061);
and U7289 (N_7289,N_7095,N_7144);
nor U7290 (N_7290,N_7088,N_7001);
nor U7291 (N_7291,N_7090,N_7093);
nand U7292 (N_7292,N_7146,N_7006);
nand U7293 (N_7293,N_7152,N_7083);
or U7294 (N_7294,N_7047,N_7087);
nand U7295 (N_7295,N_7174,N_7012);
nor U7296 (N_7296,N_7118,N_7100);
nor U7297 (N_7297,N_7033,N_7183);
xnor U7298 (N_7298,N_7076,N_7163);
nor U7299 (N_7299,N_7201,N_7214);
and U7300 (N_7300,N_7107,N_7073);
or U7301 (N_7301,N_7051,N_7109);
xor U7302 (N_7302,N_7212,N_7053);
nor U7303 (N_7303,N_7165,N_7204);
and U7304 (N_7304,N_7082,N_7035);
nand U7305 (N_7305,N_7086,N_7194);
nand U7306 (N_7306,N_7240,N_7067);
or U7307 (N_7307,N_7247,N_7243);
xor U7308 (N_7308,N_7123,N_7149);
nor U7309 (N_7309,N_7156,N_7116);
or U7310 (N_7310,N_7017,N_7148);
xor U7311 (N_7311,N_7044,N_7106);
or U7312 (N_7312,N_7005,N_7102);
and U7313 (N_7313,N_7014,N_7112);
nor U7314 (N_7314,N_7040,N_7158);
nand U7315 (N_7315,N_7151,N_7101);
nor U7316 (N_7316,N_7208,N_7179);
or U7317 (N_7317,N_7128,N_7105);
and U7318 (N_7318,N_7108,N_7167);
or U7319 (N_7319,N_7132,N_7230);
and U7320 (N_7320,N_7062,N_7064);
nor U7321 (N_7321,N_7022,N_7021);
xnor U7322 (N_7322,N_7024,N_7173);
or U7323 (N_7323,N_7126,N_7155);
nand U7324 (N_7324,N_7248,N_7120);
or U7325 (N_7325,N_7069,N_7150);
nand U7326 (N_7326,N_7070,N_7046);
nand U7327 (N_7327,N_7180,N_7016);
and U7328 (N_7328,N_7210,N_7115);
nand U7329 (N_7329,N_7192,N_7015);
or U7330 (N_7330,N_7235,N_7068);
xor U7331 (N_7331,N_7249,N_7209);
xor U7332 (N_7332,N_7013,N_7111);
nand U7333 (N_7333,N_7049,N_7181);
or U7334 (N_7334,N_7175,N_7138);
xor U7335 (N_7335,N_7176,N_7099);
nand U7336 (N_7336,N_7057,N_7081);
xor U7337 (N_7337,N_7228,N_7195);
xnor U7338 (N_7338,N_7213,N_7238);
or U7339 (N_7339,N_7216,N_7050);
nand U7340 (N_7340,N_7242,N_7207);
nand U7341 (N_7341,N_7097,N_7029);
nor U7342 (N_7342,N_7009,N_7122);
nor U7343 (N_7343,N_7056,N_7159);
or U7344 (N_7344,N_7232,N_7244);
nand U7345 (N_7345,N_7025,N_7048);
or U7346 (N_7346,N_7236,N_7077);
or U7347 (N_7347,N_7223,N_7200);
nand U7348 (N_7348,N_7007,N_7089);
xnor U7349 (N_7349,N_7055,N_7084);
xor U7350 (N_7350,N_7037,N_7066);
or U7351 (N_7351,N_7036,N_7178);
or U7352 (N_7352,N_7142,N_7218);
or U7353 (N_7353,N_7119,N_7166);
and U7354 (N_7354,N_7030,N_7125);
and U7355 (N_7355,N_7140,N_7241);
or U7356 (N_7356,N_7038,N_7215);
xor U7357 (N_7357,N_7147,N_7085);
and U7358 (N_7358,N_7117,N_7098);
nor U7359 (N_7359,N_7074,N_7010);
and U7360 (N_7360,N_7233,N_7237);
and U7361 (N_7361,N_7043,N_7245);
and U7362 (N_7362,N_7041,N_7096);
or U7363 (N_7363,N_7060,N_7091);
or U7364 (N_7364,N_7075,N_7034);
or U7365 (N_7365,N_7229,N_7221);
and U7366 (N_7366,N_7197,N_7058);
xor U7367 (N_7367,N_7026,N_7190);
nand U7368 (N_7368,N_7139,N_7186);
xor U7369 (N_7369,N_7065,N_7079);
xnor U7370 (N_7370,N_7133,N_7199);
xor U7371 (N_7371,N_7008,N_7227);
xnor U7372 (N_7372,N_7143,N_7011);
xnor U7373 (N_7373,N_7205,N_7153);
nand U7374 (N_7374,N_7094,N_7198);
nor U7375 (N_7375,N_7042,N_7030);
nor U7376 (N_7376,N_7153,N_7037);
nand U7377 (N_7377,N_7132,N_7129);
and U7378 (N_7378,N_7054,N_7098);
xor U7379 (N_7379,N_7091,N_7048);
nor U7380 (N_7380,N_7213,N_7066);
nor U7381 (N_7381,N_7049,N_7083);
xnor U7382 (N_7382,N_7220,N_7156);
and U7383 (N_7383,N_7156,N_7109);
or U7384 (N_7384,N_7143,N_7241);
nand U7385 (N_7385,N_7067,N_7125);
nand U7386 (N_7386,N_7224,N_7236);
nor U7387 (N_7387,N_7091,N_7155);
or U7388 (N_7388,N_7126,N_7003);
nand U7389 (N_7389,N_7040,N_7130);
nand U7390 (N_7390,N_7188,N_7131);
xnor U7391 (N_7391,N_7248,N_7061);
nand U7392 (N_7392,N_7190,N_7020);
xor U7393 (N_7393,N_7017,N_7227);
and U7394 (N_7394,N_7117,N_7110);
xor U7395 (N_7395,N_7013,N_7088);
nor U7396 (N_7396,N_7203,N_7200);
or U7397 (N_7397,N_7174,N_7043);
and U7398 (N_7398,N_7020,N_7013);
xnor U7399 (N_7399,N_7157,N_7148);
xor U7400 (N_7400,N_7167,N_7026);
nand U7401 (N_7401,N_7220,N_7050);
nand U7402 (N_7402,N_7057,N_7192);
nor U7403 (N_7403,N_7031,N_7085);
and U7404 (N_7404,N_7106,N_7008);
xor U7405 (N_7405,N_7187,N_7006);
nor U7406 (N_7406,N_7127,N_7155);
and U7407 (N_7407,N_7230,N_7162);
or U7408 (N_7408,N_7212,N_7030);
nand U7409 (N_7409,N_7238,N_7127);
nand U7410 (N_7410,N_7186,N_7098);
nand U7411 (N_7411,N_7016,N_7146);
or U7412 (N_7412,N_7009,N_7022);
and U7413 (N_7413,N_7012,N_7054);
and U7414 (N_7414,N_7143,N_7150);
nand U7415 (N_7415,N_7041,N_7072);
nand U7416 (N_7416,N_7194,N_7189);
or U7417 (N_7417,N_7039,N_7051);
and U7418 (N_7418,N_7140,N_7080);
nand U7419 (N_7419,N_7066,N_7174);
xor U7420 (N_7420,N_7125,N_7199);
and U7421 (N_7421,N_7211,N_7019);
xor U7422 (N_7422,N_7210,N_7204);
or U7423 (N_7423,N_7176,N_7056);
or U7424 (N_7424,N_7173,N_7053);
and U7425 (N_7425,N_7051,N_7097);
nor U7426 (N_7426,N_7187,N_7130);
xor U7427 (N_7427,N_7100,N_7148);
nand U7428 (N_7428,N_7001,N_7147);
nor U7429 (N_7429,N_7040,N_7030);
xor U7430 (N_7430,N_7002,N_7184);
xor U7431 (N_7431,N_7210,N_7045);
nand U7432 (N_7432,N_7087,N_7199);
xor U7433 (N_7433,N_7016,N_7058);
or U7434 (N_7434,N_7058,N_7201);
nor U7435 (N_7435,N_7086,N_7135);
nor U7436 (N_7436,N_7004,N_7208);
or U7437 (N_7437,N_7088,N_7032);
nor U7438 (N_7438,N_7229,N_7117);
nor U7439 (N_7439,N_7139,N_7095);
nand U7440 (N_7440,N_7181,N_7226);
nand U7441 (N_7441,N_7199,N_7244);
nor U7442 (N_7442,N_7132,N_7177);
nand U7443 (N_7443,N_7244,N_7111);
xor U7444 (N_7444,N_7113,N_7005);
nand U7445 (N_7445,N_7005,N_7206);
or U7446 (N_7446,N_7085,N_7209);
nand U7447 (N_7447,N_7052,N_7017);
xnor U7448 (N_7448,N_7099,N_7200);
or U7449 (N_7449,N_7029,N_7153);
and U7450 (N_7450,N_7249,N_7037);
nand U7451 (N_7451,N_7223,N_7174);
xnor U7452 (N_7452,N_7238,N_7235);
nand U7453 (N_7453,N_7149,N_7237);
and U7454 (N_7454,N_7169,N_7016);
nor U7455 (N_7455,N_7202,N_7191);
nor U7456 (N_7456,N_7123,N_7033);
nor U7457 (N_7457,N_7156,N_7191);
nor U7458 (N_7458,N_7036,N_7006);
xor U7459 (N_7459,N_7099,N_7059);
nand U7460 (N_7460,N_7103,N_7168);
xor U7461 (N_7461,N_7030,N_7208);
nor U7462 (N_7462,N_7157,N_7139);
nor U7463 (N_7463,N_7079,N_7239);
nor U7464 (N_7464,N_7014,N_7105);
nand U7465 (N_7465,N_7163,N_7207);
xor U7466 (N_7466,N_7207,N_7216);
xnor U7467 (N_7467,N_7145,N_7042);
nor U7468 (N_7468,N_7224,N_7185);
and U7469 (N_7469,N_7071,N_7151);
xnor U7470 (N_7470,N_7141,N_7136);
or U7471 (N_7471,N_7150,N_7170);
nor U7472 (N_7472,N_7187,N_7226);
nand U7473 (N_7473,N_7012,N_7080);
or U7474 (N_7474,N_7036,N_7240);
nor U7475 (N_7475,N_7088,N_7094);
and U7476 (N_7476,N_7234,N_7156);
nand U7477 (N_7477,N_7036,N_7040);
and U7478 (N_7478,N_7123,N_7166);
nor U7479 (N_7479,N_7127,N_7038);
nor U7480 (N_7480,N_7115,N_7006);
and U7481 (N_7481,N_7173,N_7103);
nand U7482 (N_7482,N_7183,N_7244);
xor U7483 (N_7483,N_7172,N_7182);
xnor U7484 (N_7484,N_7187,N_7166);
or U7485 (N_7485,N_7059,N_7222);
nand U7486 (N_7486,N_7032,N_7000);
or U7487 (N_7487,N_7015,N_7077);
nand U7488 (N_7488,N_7065,N_7013);
nand U7489 (N_7489,N_7019,N_7033);
and U7490 (N_7490,N_7112,N_7067);
and U7491 (N_7491,N_7087,N_7237);
nand U7492 (N_7492,N_7216,N_7111);
nor U7493 (N_7493,N_7210,N_7142);
nor U7494 (N_7494,N_7055,N_7030);
nand U7495 (N_7495,N_7179,N_7093);
xnor U7496 (N_7496,N_7066,N_7053);
or U7497 (N_7497,N_7009,N_7235);
nor U7498 (N_7498,N_7176,N_7197);
xnor U7499 (N_7499,N_7196,N_7102);
or U7500 (N_7500,N_7456,N_7361);
nor U7501 (N_7501,N_7292,N_7419);
and U7502 (N_7502,N_7260,N_7314);
and U7503 (N_7503,N_7278,N_7411);
or U7504 (N_7504,N_7284,N_7305);
and U7505 (N_7505,N_7420,N_7453);
or U7506 (N_7506,N_7319,N_7328);
and U7507 (N_7507,N_7477,N_7359);
xor U7508 (N_7508,N_7255,N_7499);
and U7509 (N_7509,N_7426,N_7400);
nand U7510 (N_7510,N_7395,N_7437);
and U7511 (N_7511,N_7300,N_7414);
nand U7512 (N_7512,N_7330,N_7262);
or U7513 (N_7513,N_7270,N_7341);
nor U7514 (N_7514,N_7277,N_7408);
nand U7515 (N_7515,N_7257,N_7498);
xor U7516 (N_7516,N_7464,N_7324);
nor U7517 (N_7517,N_7433,N_7335);
nand U7518 (N_7518,N_7273,N_7308);
and U7519 (N_7519,N_7457,N_7332);
nand U7520 (N_7520,N_7415,N_7425);
nand U7521 (N_7521,N_7288,N_7475);
or U7522 (N_7522,N_7274,N_7362);
nor U7523 (N_7523,N_7383,N_7470);
xor U7524 (N_7524,N_7418,N_7369);
and U7525 (N_7525,N_7334,N_7391);
xnor U7526 (N_7526,N_7476,N_7430);
nor U7527 (N_7527,N_7303,N_7325);
nor U7528 (N_7528,N_7482,N_7434);
xnor U7529 (N_7529,N_7312,N_7337);
and U7530 (N_7530,N_7250,N_7364);
or U7531 (N_7531,N_7340,N_7298);
nand U7532 (N_7532,N_7465,N_7385);
xnor U7533 (N_7533,N_7387,N_7342);
nand U7534 (N_7534,N_7377,N_7368);
xnor U7535 (N_7535,N_7406,N_7279);
or U7536 (N_7536,N_7469,N_7458);
nand U7537 (N_7537,N_7331,N_7378);
or U7538 (N_7538,N_7269,N_7263);
xnor U7539 (N_7539,N_7344,N_7353);
xnor U7540 (N_7540,N_7490,N_7450);
xnor U7541 (N_7541,N_7393,N_7253);
nor U7542 (N_7542,N_7407,N_7259);
xor U7543 (N_7543,N_7297,N_7311);
nor U7544 (N_7544,N_7268,N_7461);
nor U7545 (N_7545,N_7296,N_7401);
nand U7546 (N_7546,N_7290,N_7496);
nand U7547 (N_7547,N_7294,N_7447);
nand U7548 (N_7548,N_7375,N_7322);
xnor U7549 (N_7549,N_7439,N_7355);
xor U7550 (N_7550,N_7388,N_7301);
nand U7551 (N_7551,N_7380,N_7316);
xnor U7552 (N_7552,N_7452,N_7267);
and U7553 (N_7553,N_7487,N_7405);
nand U7554 (N_7554,N_7363,N_7497);
nand U7555 (N_7555,N_7356,N_7409);
xor U7556 (N_7556,N_7462,N_7379);
nor U7557 (N_7557,N_7373,N_7351);
nor U7558 (N_7558,N_7390,N_7365);
xor U7559 (N_7559,N_7327,N_7360);
and U7560 (N_7560,N_7317,N_7323);
nor U7561 (N_7561,N_7252,N_7310);
and U7562 (N_7562,N_7329,N_7424);
nand U7563 (N_7563,N_7333,N_7371);
nor U7564 (N_7564,N_7438,N_7471);
and U7565 (N_7565,N_7402,N_7285);
xnor U7566 (N_7566,N_7441,N_7302);
xnor U7567 (N_7567,N_7473,N_7442);
xnor U7568 (N_7568,N_7386,N_7480);
and U7569 (N_7569,N_7410,N_7306);
nor U7570 (N_7570,N_7384,N_7404);
nand U7571 (N_7571,N_7397,N_7256);
xor U7572 (N_7572,N_7454,N_7449);
xor U7573 (N_7573,N_7428,N_7478);
or U7574 (N_7574,N_7488,N_7336);
xnor U7575 (N_7575,N_7343,N_7304);
xor U7576 (N_7576,N_7354,N_7416);
nor U7577 (N_7577,N_7276,N_7339);
nor U7578 (N_7578,N_7318,N_7350);
nand U7579 (N_7579,N_7491,N_7287);
and U7580 (N_7580,N_7352,N_7467);
nand U7581 (N_7581,N_7423,N_7348);
or U7582 (N_7582,N_7264,N_7429);
or U7583 (N_7583,N_7398,N_7271);
xnor U7584 (N_7584,N_7315,N_7466);
nand U7585 (N_7585,N_7486,N_7421);
and U7586 (N_7586,N_7459,N_7258);
and U7587 (N_7587,N_7448,N_7484);
nand U7588 (N_7588,N_7338,N_7394);
nor U7589 (N_7589,N_7474,N_7254);
or U7590 (N_7590,N_7451,N_7345);
nand U7591 (N_7591,N_7280,N_7366);
nand U7592 (N_7592,N_7445,N_7396);
or U7593 (N_7593,N_7265,N_7320);
nand U7594 (N_7594,N_7436,N_7309);
and U7595 (N_7595,N_7389,N_7489);
or U7596 (N_7596,N_7349,N_7293);
or U7597 (N_7597,N_7376,N_7272);
nand U7598 (N_7598,N_7494,N_7346);
and U7599 (N_7599,N_7291,N_7275);
nor U7600 (N_7600,N_7463,N_7326);
and U7601 (N_7601,N_7431,N_7468);
nand U7602 (N_7602,N_7372,N_7367);
and U7603 (N_7603,N_7281,N_7321);
xor U7604 (N_7604,N_7446,N_7392);
nand U7605 (N_7605,N_7370,N_7417);
xor U7606 (N_7606,N_7495,N_7266);
nand U7607 (N_7607,N_7382,N_7251);
or U7608 (N_7608,N_7381,N_7460);
nor U7609 (N_7609,N_7295,N_7283);
and U7610 (N_7610,N_7357,N_7261);
or U7611 (N_7611,N_7412,N_7479);
and U7612 (N_7612,N_7313,N_7347);
or U7613 (N_7613,N_7427,N_7422);
or U7614 (N_7614,N_7483,N_7443);
xnor U7615 (N_7615,N_7358,N_7435);
nand U7616 (N_7616,N_7472,N_7485);
or U7617 (N_7617,N_7289,N_7440);
nor U7618 (N_7618,N_7413,N_7481);
and U7619 (N_7619,N_7299,N_7403);
nand U7620 (N_7620,N_7307,N_7492);
xor U7621 (N_7621,N_7286,N_7374);
or U7622 (N_7622,N_7432,N_7455);
nor U7623 (N_7623,N_7493,N_7444);
xnor U7624 (N_7624,N_7282,N_7399);
xnor U7625 (N_7625,N_7388,N_7487);
nor U7626 (N_7626,N_7328,N_7305);
nor U7627 (N_7627,N_7497,N_7378);
nand U7628 (N_7628,N_7392,N_7471);
nor U7629 (N_7629,N_7405,N_7262);
and U7630 (N_7630,N_7440,N_7265);
xnor U7631 (N_7631,N_7443,N_7473);
or U7632 (N_7632,N_7419,N_7484);
nand U7633 (N_7633,N_7416,N_7495);
and U7634 (N_7634,N_7292,N_7331);
or U7635 (N_7635,N_7327,N_7316);
xnor U7636 (N_7636,N_7406,N_7468);
nor U7637 (N_7637,N_7476,N_7379);
xnor U7638 (N_7638,N_7447,N_7316);
xor U7639 (N_7639,N_7398,N_7479);
and U7640 (N_7640,N_7335,N_7291);
xor U7641 (N_7641,N_7374,N_7297);
xnor U7642 (N_7642,N_7341,N_7328);
and U7643 (N_7643,N_7357,N_7480);
and U7644 (N_7644,N_7284,N_7378);
and U7645 (N_7645,N_7325,N_7354);
xor U7646 (N_7646,N_7438,N_7291);
nor U7647 (N_7647,N_7396,N_7303);
nand U7648 (N_7648,N_7381,N_7387);
nand U7649 (N_7649,N_7358,N_7339);
and U7650 (N_7650,N_7283,N_7461);
nand U7651 (N_7651,N_7408,N_7357);
xnor U7652 (N_7652,N_7351,N_7439);
nor U7653 (N_7653,N_7329,N_7339);
and U7654 (N_7654,N_7370,N_7255);
or U7655 (N_7655,N_7404,N_7268);
xor U7656 (N_7656,N_7428,N_7489);
nand U7657 (N_7657,N_7396,N_7315);
nand U7658 (N_7658,N_7332,N_7433);
nand U7659 (N_7659,N_7260,N_7272);
xnor U7660 (N_7660,N_7352,N_7487);
and U7661 (N_7661,N_7492,N_7355);
and U7662 (N_7662,N_7460,N_7308);
nand U7663 (N_7663,N_7474,N_7272);
xor U7664 (N_7664,N_7388,N_7491);
nor U7665 (N_7665,N_7271,N_7419);
nand U7666 (N_7666,N_7499,N_7448);
and U7667 (N_7667,N_7256,N_7483);
nor U7668 (N_7668,N_7436,N_7339);
nand U7669 (N_7669,N_7272,N_7353);
xor U7670 (N_7670,N_7444,N_7282);
and U7671 (N_7671,N_7286,N_7381);
nand U7672 (N_7672,N_7279,N_7477);
or U7673 (N_7673,N_7367,N_7270);
or U7674 (N_7674,N_7387,N_7368);
and U7675 (N_7675,N_7475,N_7412);
and U7676 (N_7676,N_7427,N_7461);
and U7677 (N_7677,N_7486,N_7368);
nand U7678 (N_7678,N_7402,N_7345);
and U7679 (N_7679,N_7277,N_7435);
or U7680 (N_7680,N_7368,N_7472);
nor U7681 (N_7681,N_7488,N_7485);
or U7682 (N_7682,N_7477,N_7310);
xor U7683 (N_7683,N_7349,N_7289);
and U7684 (N_7684,N_7271,N_7255);
and U7685 (N_7685,N_7495,N_7448);
or U7686 (N_7686,N_7408,N_7450);
and U7687 (N_7687,N_7394,N_7382);
and U7688 (N_7688,N_7352,N_7438);
and U7689 (N_7689,N_7359,N_7412);
nor U7690 (N_7690,N_7390,N_7477);
xnor U7691 (N_7691,N_7441,N_7466);
xnor U7692 (N_7692,N_7329,N_7294);
nand U7693 (N_7693,N_7337,N_7438);
and U7694 (N_7694,N_7476,N_7492);
nor U7695 (N_7695,N_7296,N_7482);
and U7696 (N_7696,N_7325,N_7290);
nand U7697 (N_7697,N_7256,N_7357);
nand U7698 (N_7698,N_7359,N_7438);
xor U7699 (N_7699,N_7480,N_7269);
nand U7700 (N_7700,N_7365,N_7445);
or U7701 (N_7701,N_7282,N_7456);
nand U7702 (N_7702,N_7348,N_7337);
and U7703 (N_7703,N_7499,N_7268);
and U7704 (N_7704,N_7422,N_7278);
nand U7705 (N_7705,N_7335,N_7372);
nor U7706 (N_7706,N_7335,N_7329);
and U7707 (N_7707,N_7344,N_7447);
nor U7708 (N_7708,N_7330,N_7386);
xor U7709 (N_7709,N_7336,N_7455);
xor U7710 (N_7710,N_7452,N_7435);
and U7711 (N_7711,N_7411,N_7310);
xor U7712 (N_7712,N_7264,N_7450);
or U7713 (N_7713,N_7413,N_7476);
and U7714 (N_7714,N_7480,N_7388);
nor U7715 (N_7715,N_7273,N_7327);
and U7716 (N_7716,N_7279,N_7422);
nor U7717 (N_7717,N_7304,N_7336);
and U7718 (N_7718,N_7337,N_7266);
nor U7719 (N_7719,N_7254,N_7347);
or U7720 (N_7720,N_7324,N_7468);
and U7721 (N_7721,N_7322,N_7474);
nor U7722 (N_7722,N_7384,N_7296);
xnor U7723 (N_7723,N_7387,N_7448);
or U7724 (N_7724,N_7487,N_7282);
xor U7725 (N_7725,N_7464,N_7431);
nor U7726 (N_7726,N_7486,N_7308);
and U7727 (N_7727,N_7414,N_7404);
xnor U7728 (N_7728,N_7420,N_7337);
nor U7729 (N_7729,N_7392,N_7435);
nand U7730 (N_7730,N_7465,N_7482);
nand U7731 (N_7731,N_7380,N_7405);
or U7732 (N_7732,N_7436,N_7356);
and U7733 (N_7733,N_7450,N_7432);
nor U7734 (N_7734,N_7434,N_7331);
or U7735 (N_7735,N_7252,N_7286);
nand U7736 (N_7736,N_7455,N_7321);
or U7737 (N_7737,N_7266,N_7412);
nand U7738 (N_7738,N_7350,N_7484);
xor U7739 (N_7739,N_7438,N_7301);
nand U7740 (N_7740,N_7448,N_7462);
and U7741 (N_7741,N_7386,N_7407);
or U7742 (N_7742,N_7416,N_7396);
and U7743 (N_7743,N_7461,N_7394);
and U7744 (N_7744,N_7386,N_7318);
nor U7745 (N_7745,N_7381,N_7453);
and U7746 (N_7746,N_7444,N_7325);
xor U7747 (N_7747,N_7363,N_7255);
and U7748 (N_7748,N_7370,N_7294);
nor U7749 (N_7749,N_7359,N_7293);
nor U7750 (N_7750,N_7726,N_7694);
and U7751 (N_7751,N_7669,N_7698);
xnor U7752 (N_7752,N_7520,N_7574);
or U7753 (N_7753,N_7730,N_7558);
nor U7754 (N_7754,N_7582,N_7637);
or U7755 (N_7755,N_7618,N_7608);
or U7756 (N_7756,N_7510,N_7530);
xor U7757 (N_7757,N_7549,N_7681);
or U7758 (N_7758,N_7528,N_7629);
nor U7759 (N_7759,N_7733,N_7553);
xor U7760 (N_7760,N_7704,N_7740);
or U7761 (N_7761,N_7573,N_7602);
or U7762 (N_7762,N_7588,N_7655);
and U7763 (N_7763,N_7557,N_7531);
or U7764 (N_7764,N_7601,N_7703);
or U7765 (N_7765,N_7554,N_7591);
and U7766 (N_7766,N_7643,N_7693);
and U7767 (N_7767,N_7578,N_7514);
xor U7768 (N_7768,N_7718,N_7749);
xor U7769 (N_7769,N_7671,N_7529);
and U7770 (N_7770,N_7536,N_7640);
or U7771 (N_7771,N_7533,N_7515);
or U7772 (N_7772,N_7727,N_7571);
xnor U7773 (N_7773,N_7567,N_7663);
or U7774 (N_7774,N_7611,N_7562);
nand U7775 (N_7775,N_7638,N_7662);
xnor U7776 (N_7776,N_7687,N_7737);
and U7777 (N_7777,N_7508,N_7566);
and U7778 (N_7778,N_7517,N_7524);
or U7779 (N_7779,N_7604,N_7595);
or U7780 (N_7780,N_7700,N_7642);
nand U7781 (N_7781,N_7501,N_7555);
xor U7782 (N_7782,N_7587,N_7691);
or U7783 (N_7783,N_7584,N_7542);
xnor U7784 (N_7784,N_7717,N_7610);
nor U7785 (N_7785,N_7725,N_7634);
and U7786 (N_7786,N_7736,N_7516);
nor U7787 (N_7787,N_7722,N_7563);
xor U7788 (N_7788,N_7512,N_7678);
xor U7789 (N_7789,N_7504,N_7556);
nand U7790 (N_7790,N_7713,N_7652);
or U7791 (N_7791,N_7551,N_7645);
xor U7792 (N_7792,N_7589,N_7715);
xor U7793 (N_7793,N_7646,N_7711);
nor U7794 (N_7794,N_7689,N_7626);
and U7795 (N_7795,N_7699,N_7561);
or U7796 (N_7796,N_7621,N_7630);
and U7797 (N_7797,N_7500,N_7743);
nor U7798 (N_7798,N_7709,N_7522);
nand U7799 (N_7799,N_7633,N_7649);
nor U7800 (N_7800,N_7635,N_7632);
or U7801 (N_7801,N_7503,N_7619);
xnor U7802 (N_7802,N_7732,N_7576);
nand U7803 (N_7803,N_7534,N_7661);
xnor U7804 (N_7804,N_7653,N_7712);
or U7805 (N_7805,N_7540,N_7721);
or U7806 (N_7806,N_7741,N_7716);
xor U7807 (N_7807,N_7507,N_7747);
or U7808 (N_7808,N_7575,N_7731);
or U7809 (N_7809,N_7547,N_7583);
nand U7810 (N_7810,N_7523,N_7586);
nor U7811 (N_7811,N_7541,N_7739);
xnor U7812 (N_7812,N_7624,N_7605);
xnor U7813 (N_7813,N_7603,N_7692);
nand U7814 (N_7814,N_7525,N_7686);
and U7815 (N_7815,N_7690,N_7639);
nand U7816 (N_7816,N_7746,N_7532);
or U7817 (N_7817,N_7666,N_7647);
or U7818 (N_7818,N_7674,N_7545);
nor U7819 (N_7819,N_7723,N_7565);
xor U7820 (N_7820,N_7615,N_7577);
and U7821 (N_7821,N_7708,N_7641);
xor U7822 (N_7822,N_7654,N_7735);
nand U7823 (N_7823,N_7585,N_7535);
nand U7824 (N_7824,N_7707,N_7623);
xor U7825 (N_7825,N_7506,N_7617);
or U7826 (N_7826,N_7527,N_7616);
nor U7827 (N_7827,N_7680,N_7636);
xor U7828 (N_7828,N_7590,N_7609);
nand U7829 (N_7829,N_7676,N_7648);
xor U7830 (N_7830,N_7673,N_7580);
nor U7831 (N_7831,N_7606,N_7569);
or U7832 (N_7832,N_7724,N_7656);
nand U7833 (N_7833,N_7612,N_7683);
xor U7834 (N_7834,N_7706,N_7650);
nand U7835 (N_7835,N_7742,N_7701);
nand U7836 (N_7836,N_7657,N_7519);
or U7837 (N_7837,N_7684,N_7744);
nand U7838 (N_7838,N_7631,N_7627);
nand U7839 (N_7839,N_7596,N_7625);
nor U7840 (N_7840,N_7594,N_7719);
nor U7841 (N_7841,N_7564,N_7728);
or U7842 (N_7842,N_7570,N_7695);
xor U7843 (N_7843,N_7672,N_7548);
xnor U7844 (N_7844,N_7600,N_7720);
nand U7845 (N_7845,N_7607,N_7651);
nor U7846 (N_7846,N_7592,N_7659);
and U7847 (N_7847,N_7622,N_7729);
and U7848 (N_7848,N_7660,N_7521);
and U7849 (N_7849,N_7544,N_7710);
and U7850 (N_7850,N_7675,N_7513);
and U7851 (N_7851,N_7559,N_7579);
xnor U7852 (N_7852,N_7679,N_7518);
and U7853 (N_7853,N_7682,N_7658);
nor U7854 (N_7854,N_7664,N_7668);
nor U7855 (N_7855,N_7511,N_7734);
and U7856 (N_7856,N_7597,N_7526);
or U7857 (N_7857,N_7546,N_7745);
xnor U7858 (N_7858,N_7614,N_7644);
nor U7859 (N_7859,N_7543,N_7677);
nand U7860 (N_7860,N_7560,N_7581);
xnor U7861 (N_7861,N_7613,N_7502);
nand U7862 (N_7862,N_7685,N_7599);
and U7863 (N_7863,N_7552,N_7665);
nand U7864 (N_7864,N_7620,N_7670);
or U7865 (N_7865,N_7550,N_7705);
and U7866 (N_7866,N_7568,N_7539);
xnor U7867 (N_7867,N_7593,N_7509);
xor U7868 (N_7868,N_7667,N_7714);
and U7869 (N_7869,N_7628,N_7572);
and U7870 (N_7870,N_7696,N_7538);
and U7871 (N_7871,N_7702,N_7738);
nand U7872 (N_7872,N_7748,N_7598);
nor U7873 (N_7873,N_7697,N_7505);
or U7874 (N_7874,N_7537,N_7688);
nand U7875 (N_7875,N_7506,N_7551);
and U7876 (N_7876,N_7591,N_7517);
nor U7877 (N_7877,N_7595,N_7519);
xor U7878 (N_7878,N_7594,N_7722);
xnor U7879 (N_7879,N_7720,N_7703);
and U7880 (N_7880,N_7520,N_7611);
and U7881 (N_7881,N_7619,N_7701);
and U7882 (N_7882,N_7693,N_7559);
nand U7883 (N_7883,N_7584,N_7564);
and U7884 (N_7884,N_7551,N_7684);
and U7885 (N_7885,N_7617,N_7703);
nor U7886 (N_7886,N_7660,N_7549);
and U7887 (N_7887,N_7617,N_7566);
or U7888 (N_7888,N_7642,N_7633);
nand U7889 (N_7889,N_7561,N_7574);
nand U7890 (N_7890,N_7658,N_7695);
nor U7891 (N_7891,N_7631,N_7641);
and U7892 (N_7892,N_7599,N_7735);
and U7893 (N_7893,N_7541,N_7711);
xor U7894 (N_7894,N_7542,N_7686);
xnor U7895 (N_7895,N_7625,N_7735);
xor U7896 (N_7896,N_7502,N_7525);
nand U7897 (N_7897,N_7534,N_7584);
or U7898 (N_7898,N_7646,N_7631);
or U7899 (N_7899,N_7516,N_7744);
nor U7900 (N_7900,N_7563,N_7537);
and U7901 (N_7901,N_7521,N_7578);
xnor U7902 (N_7902,N_7703,N_7740);
or U7903 (N_7903,N_7676,N_7634);
and U7904 (N_7904,N_7741,N_7506);
and U7905 (N_7905,N_7566,N_7540);
nand U7906 (N_7906,N_7652,N_7638);
or U7907 (N_7907,N_7529,N_7598);
and U7908 (N_7908,N_7594,N_7696);
xor U7909 (N_7909,N_7628,N_7578);
xor U7910 (N_7910,N_7524,N_7609);
or U7911 (N_7911,N_7610,N_7564);
and U7912 (N_7912,N_7555,N_7614);
nand U7913 (N_7913,N_7630,N_7736);
nor U7914 (N_7914,N_7525,N_7643);
and U7915 (N_7915,N_7695,N_7726);
nand U7916 (N_7916,N_7645,N_7608);
or U7917 (N_7917,N_7576,N_7606);
nor U7918 (N_7918,N_7643,N_7719);
xor U7919 (N_7919,N_7711,N_7517);
xor U7920 (N_7920,N_7515,N_7547);
nand U7921 (N_7921,N_7546,N_7744);
nor U7922 (N_7922,N_7542,N_7611);
and U7923 (N_7923,N_7670,N_7720);
nand U7924 (N_7924,N_7564,N_7683);
xor U7925 (N_7925,N_7611,N_7710);
nor U7926 (N_7926,N_7725,N_7501);
and U7927 (N_7927,N_7735,N_7586);
xor U7928 (N_7928,N_7743,N_7622);
or U7929 (N_7929,N_7704,N_7521);
and U7930 (N_7930,N_7744,N_7691);
and U7931 (N_7931,N_7508,N_7646);
xor U7932 (N_7932,N_7501,N_7706);
or U7933 (N_7933,N_7566,N_7568);
nand U7934 (N_7934,N_7529,N_7710);
nor U7935 (N_7935,N_7606,N_7660);
nor U7936 (N_7936,N_7735,N_7557);
nand U7937 (N_7937,N_7688,N_7576);
nand U7938 (N_7938,N_7578,N_7725);
xnor U7939 (N_7939,N_7659,N_7529);
or U7940 (N_7940,N_7744,N_7550);
xnor U7941 (N_7941,N_7670,N_7730);
xor U7942 (N_7942,N_7661,N_7678);
xor U7943 (N_7943,N_7590,N_7639);
and U7944 (N_7944,N_7709,N_7590);
xnor U7945 (N_7945,N_7506,N_7646);
nor U7946 (N_7946,N_7647,N_7702);
nand U7947 (N_7947,N_7541,N_7599);
nor U7948 (N_7948,N_7537,N_7632);
or U7949 (N_7949,N_7689,N_7722);
or U7950 (N_7950,N_7576,N_7600);
nand U7951 (N_7951,N_7531,N_7682);
nand U7952 (N_7952,N_7620,N_7549);
or U7953 (N_7953,N_7651,N_7598);
nor U7954 (N_7954,N_7584,N_7525);
xor U7955 (N_7955,N_7680,N_7527);
and U7956 (N_7956,N_7641,N_7571);
nor U7957 (N_7957,N_7544,N_7590);
and U7958 (N_7958,N_7528,N_7744);
and U7959 (N_7959,N_7545,N_7682);
xor U7960 (N_7960,N_7721,N_7511);
or U7961 (N_7961,N_7546,N_7608);
nor U7962 (N_7962,N_7671,N_7558);
nor U7963 (N_7963,N_7527,N_7557);
xnor U7964 (N_7964,N_7558,N_7695);
and U7965 (N_7965,N_7540,N_7503);
xor U7966 (N_7966,N_7531,N_7637);
or U7967 (N_7967,N_7741,N_7573);
or U7968 (N_7968,N_7702,N_7605);
xnor U7969 (N_7969,N_7701,N_7571);
and U7970 (N_7970,N_7697,N_7511);
and U7971 (N_7971,N_7747,N_7619);
and U7972 (N_7972,N_7665,N_7706);
and U7973 (N_7973,N_7653,N_7525);
nand U7974 (N_7974,N_7501,N_7656);
or U7975 (N_7975,N_7516,N_7660);
nand U7976 (N_7976,N_7589,N_7562);
xor U7977 (N_7977,N_7525,N_7504);
xnor U7978 (N_7978,N_7537,N_7518);
xor U7979 (N_7979,N_7684,N_7715);
xnor U7980 (N_7980,N_7535,N_7696);
and U7981 (N_7981,N_7552,N_7673);
or U7982 (N_7982,N_7725,N_7685);
nand U7983 (N_7983,N_7544,N_7674);
nor U7984 (N_7984,N_7524,N_7506);
xor U7985 (N_7985,N_7636,N_7731);
or U7986 (N_7986,N_7714,N_7541);
xnor U7987 (N_7987,N_7500,N_7627);
and U7988 (N_7988,N_7679,N_7620);
xor U7989 (N_7989,N_7633,N_7529);
nor U7990 (N_7990,N_7658,N_7713);
xor U7991 (N_7991,N_7745,N_7594);
and U7992 (N_7992,N_7555,N_7730);
and U7993 (N_7993,N_7732,N_7579);
nor U7994 (N_7994,N_7614,N_7735);
or U7995 (N_7995,N_7745,N_7625);
and U7996 (N_7996,N_7599,N_7618);
xnor U7997 (N_7997,N_7586,N_7673);
nand U7998 (N_7998,N_7667,N_7525);
or U7999 (N_7999,N_7623,N_7629);
xnor U8000 (N_8000,N_7785,N_7954);
or U8001 (N_8001,N_7826,N_7771);
xor U8002 (N_8002,N_7788,N_7829);
xor U8003 (N_8003,N_7979,N_7922);
and U8004 (N_8004,N_7989,N_7834);
and U8005 (N_8005,N_7844,N_7816);
nor U8006 (N_8006,N_7876,N_7973);
xor U8007 (N_8007,N_7787,N_7934);
and U8008 (N_8008,N_7755,N_7839);
xor U8009 (N_8009,N_7814,N_7808);
and U8010 (N_8010,N_7982,N_7843);
nand U8011 (N_8011,N_7978,N_7825);
or U8012 (N_8012,N_7789,N_7828);
nor U8013 (N_8013,N_7772,N_7952);
or U8014 (N_8014,N_7965,N_7991);
and U8015 (N_8015,N_7783,N_7900);
and U8016 (N_8016,N_7903,N_7907);
xor U8017 (N_8017,N_7767,N_7792);
or U8018 (N_8018,N_7803,N_7842);
nand U8019 (N_8019,N_7925,N_7874);
and U8020 (N_8020,N_7894,N_7906);
and U8021 (N_8021,N_7750,N_7801);
nand U8022 (N_8022,N_7985,N_7854);
and U8023 (N_8023,N_7951,N_7780);
xnor U8024 (N_8024,N_7984,N_7879);
xor U8025 (N_8025,N_7940,N_7892);
xor U8026 (N_8026,N_7917,N_7975);
nor U8027 (N_8027,N_7941,N_7912);
nor U8028 (N_8028,N_7840,N_7970);
xor U8029 (N_8029,N_7977,N_7891);
or U8030 (N_8030,N_7966,N_7926);
and U8031 (N_8031,N_7774,N_7886);
nor U8032 (N_8032,N_7857,N_7797);
and U8033 (N_8033,N_7962,N_7953);
xor U8034 (N_8034,N_7847,N_7961);
and U8035 (N_8035,N_7918,N_7986);
nor U8036 (N_8036,N_7791,N_7763);
nand U8037 (N_8037,N_7761,N_7893);
or U8038 (N_8038,N_7956,N_7849);
and U8039 (N_8039,N_7770,N_7905);
nor U8040 (N_8040,N_7818,N_7924);
nand U8041 (N_8041,N_7853,N_7964);
and U8042 (N_8042,N_7841,N_7757);
nor U8043 (N_8043,N_7974,N_7884);
nor U8044 (N_8044,N_7784,N_7887);
or U8045 (N_8045,N_7996,N_7890);
nand U8046 (N_8046,N_7959,N_7766);
xor U8047 (N_8047,N_7931,N_7983);
and U8048 (N_8048,N_7759,N_7955);
and U8049 (N_8049,N_7981,N_7895);
nand U8050 (N_8050,N_7942,N_7756);
nand U8051 (N_8051,N_7773,N_7846);
nand U8052 (N_8052,N_7938,N_7870);
nand U8053 (N_8053,N_7995,N_7776);
nor U8054 (N_8054,N_7817,N_7960);
nand U8055 (N_8055,N_7883,N_7999);
xnor U8056 (N_8056,N_7968,N_7899);
or U8057 (N_8057,N_7762,N_7832);
nor U8058 (N_8058,N_7971,N_7921);
nand U8059 (N_8059,N_7898,N_7781);
or U8060 (N_8060,N_7889,N_7980);
or U8061 (N_8061,N_7793,N_7831);
nor U8062 (N_8062,N_7993,N_7782);
and U8063 (N_8063,N_7779,N_7976);
nor U8064 (N_8064,N_7805,N_7822);
nor U8065 (N_8065,N_7919,N_7939);
nand U8066 (N_8066,N_7848,N_7753);
or U8067 (N_8067,N_7928,N_7888);
nor U8068 (N_8068,N_7752,N_7927);
and U8069 (N_8069,N_7865,N_7804);
or U8070 (N_8070,N_7881,N_7972);
or U8071 (N_8071,N_7994,N_7858);
xnor U8072 (N_8072,N_7944,N_7778);
and U8073 (N_8073,N_7824,N_7910);
or U8074 (N_8074,N_7802,N_7998);
nor U8075 (N_8075,N_7769,N_7947);
nand U8076 (N_8076,N_7811,N_7904);
or U8077 (N_8077,N_7936,N_7836);
nor U8078 (N_8078,N_7902,N_7815);
nand U8079 (N_8079,N_7862,N_7850);
and U8080 (N_8080,N_7914,N_7819);
nand U8081 (N_8081,N_7877,N_7861);
nor U8082 (N_8082,N_7997,N_7885);
nand U8083 (N_8083,N_7930,N_7794);
and U8084 (N_8084,N_7799,N_7880);
nor U8085 (N_8085,N_7790,N_7909);
xor U8086 (N_8086,N_7957,N_7963);
and U8087 (N_8087,N_7935,N_7923);
or U8088 (N_8088,N_7845,N_7777);
and U8089 (N_8089,N_7911,N_7946);
nand U8090 (N_8090,N_7810,N_7775);
and U8091 (N_8091,N_7988,N_7855);
nor U8092 (N_8092,N_7937,N_7837);
nor U8093 (N_8093,N_7765,N_7798);
and U8094 (N_8094,N_7807,N_7851);
and U8095 (N_8095,N_7916,N_7827);
and U8096 (N_8096,N_7920,N_7967);
nor U8097 (N_8097,N_7866,N_7913);
nor U8098 (N_8098,N_7950,N_7878);
and U8099 (N_8099,N_7949,N_7882);
nand U8100 (N_8100,N_7754,N_7856);
or U8101 (N_8101,N_7751,N_7820);
or U8102 (N_8102,N_7786,N_7863);
and U8103 (N_8103,N_7821,N_7867);
or U8104 (N_8104,N_7812,N_7908);
nor U8105 (N_8105,N_7932,N_7795);
or U8106 (N_8106,N_7760,N_7933);
or U8107 (N_8107,N_7869,N_7896);
or U8108 (N_8108,N_7852,N_7764);
and U8109 (N_8109,N_7809,N_7875);
and U8110 (N_8110,N_7958,N_7929);
nand U8111 (N_8111,N_7987,N_7823);
nor U8112 (N_8112,N_7897,N_7796);
xor U8113 (N_8113,N_7864,N_7768);
nor U8114 (N_8114,N_7838,N_7860);
nor U8115 (N_8115,N_7948,N_7833);
or U8116 (N_8116,N_7871,N_7830);
and U8117 (N_8117,N_7859,N_7813);
and U8118 (N_8118,N_7806,N_7943);
or U8119 (N_8119,N_7969,N_7915);
xnor U8120 (N_8120,N_7868,N_7901);
and U8121 (N_8121,N_7872,N_7835);
nor U8122 (N_8122,N_7945,N_7873);
nor U8123 (N_8123,N_7800,N_7992);
nor U8124 (N_8124,N_7990,N_7758);
xor U8125 (N_8125,N_7982,N_7789);
or U8126 (N_8126,N_7942,N_7864);
nand U8127 (N_8127,N_7980,N_7807);
or U8128 (N_8128,N_7752,N_7998);
or U8129 (N_8129,N_7953,N_7945);
xor U8130 (N_8130,N_7896,N_7774);
xnor U8131 (N_8131,N_7952,N_7822);
and U8132 (N_8132,N_7891,N_7846);
nor U8133 (N_8133,N_7768,N_7805);
or U8134 (N_8134,N_7907,N_7773);
or U8135 (N_8135,N_7798,N_7767);
nand U8136 (N_8136,N_7873,N_7808);
nand U8137 (N_8137,N_7763,N_7754);
nor U8138 (N_8138,N_7901,N_7959);
nor U8139 (N_8139,N_7876,N_7872);
nor U8140 (N_8140,N_7961,N_7780);
or U8141 (N_8141,N_7946,N_7814);
or U8142 (N_8142,N_7790,N_7770);
nand U8143 (N_8143,N_7772,N_7996);
or U8144 (N_8144,N_7850,N_7941);
and U8145 (N_8145,N_7771,N_7818);
nand U8146 (N_8146,N_7828,N_7889);
and U8147 (N_8147,N_7855,N_7823);
and U8148 (N_8148,N_7959,N_7845);
or U8149 (N_8149,N_7782,N_7760);
xor U8150 (N_8150,N_7826,N_7995);
or U8151 (N_8151,N_7803,N_7787);
and U8152 (N_8152,N_7758,N_7913);
nand U8153 (N_8153,N_7842,N_7956);
or U8154 (N_8154,N_7868,N_7937);
xnor U8155 (N_8155,N_7764,N_7867);
nand U8156 (N_8156,N_7827,N_7884);
or U8157 (N_8157,N_7767,N_7850);
or U8158 (N_8158,N_7853,N_7966);
and U8159 (N_8159,N_7925,N_7894);
nand U8160 (N_8160,N_7918,N_7820);
nor U8161 (N_8161,N_7805,N_7867);
xnor U8162 (N_8162,N_7921,N_7877);
nor U8163 (N_8163,N_7763,N_7773);
xnor U8164 (N_8164,N_7967,N_7758);
xnor U8165 (N_8165,N_7948,N_7785);
or U8166 (N_8166,N_7784,N_7816);
nand U8167 (N_8167,N_7912,N_7800);
xnor U8168 (N_8168,N_7876,N_7815);
or U8169 (N_8169,N_7800,N_7943);
and U8170 (N_8170,N_7888,N_7966);
and U8171 (N_8171,N_7845,N_7854);
nor U8172 (N_8172,N_7856,N_7829);
and U8173 (N_8173,N_7961,N_7815);
or U8174 (N_8174,N_7847,N_7974);
nand U8175 (N_8175,N_7992,N_7926);
nor U8176 (N_8176,N_7788,N_7766);
xor U8177 (N_8177,N_7754,N_7979);
nand U8178 (N_8178,N_7824,N_7868);
nor U8179 (N_8179,N_7817,N_7962);
nor U8180 (N_8180,N_7898,N_7807);
or U8181 (N_8181,N_7876,N_7914);
nor U8182 (N_8182,N_7948,N_7975);
nor U8183 (N_8183,N_7758,N_7854);
or U8184 (N_8184,N_7810,N_7866);
and U8185 (N_8185,N_7821,N_7883);
and U8186 (N_8186,N_7822,N_7956);
nor U8187 (N_8187,N_7802,N_7980);
nand U8188 (N_8188,N_7949,N_7792);
nor U8189 (N_8189,N_7842,N_7872);
and U8190 (N_8190,N_7828,N_7824);
and U8191 (N_8191,N_7827,N_7777);
nor U8192 (N_8192,N_7850,N_7887);
nor U8193 (N_8193,N_7918,N_7783);
and U8194 (N_8194,N_7849,N_7787);
and U8195 (N_8195,N_7862,N_7869);
or U8196 (N_8196,N_7821,N_7791);
and U8197 (N_8197,N_7840,N_7868);
xnor U8198 (N_8198,N_7839,N_7799);
nand U8199 (N_8199,N_7905,N_7941);
and U8200 (N_8200,N_7832,N_7837);
or U8201 (N_8201,N_7754,N_7995);
or U8202 (N_8202,N_7974,N_7767);
nor U8203 (N_8203,N_7859,N_7865);
xor U8204 (N_8204,N_7759,N_7983);
xor U8205 (N_8205,N_7975,N_7782);
nand U8206 (N_8206,N_7766,N_7988);
xnor U8207 (N_8207,N_7790,N_7825);
or U8208 (N_8208,N_7935,N_7912);
or U8209 (N_8209,N_7996,N_7799);
xnor U8210 (N_8210,N_7773,N_7936);
xnor U8211 (N_8211,N_7752,N_7861);
nand U8212 (N_8212,N_7893,N_7804);
or U8213 (N_8213,N_7997,N_7937);
nand U8214 (N_8214,N_7867,N_7755);
nor U8215 (N_8215,N_7945,N_7909);
xnor U8216 (N_8216,N_7942,N_7912);
and U8217 (N_8217,N_7980,N_7982);
and U8218 (N_8218,N_7954,N_7750);
and U8219 (N_8219,N_7854,N_7822);
xor U8220 (N_8220,N_7816,N_7924);
xor U8221 (N_8221,N_7836,N_7939);
nor U8222 (N_8222,N_7997,N_7982);
and U8223 (N_8223,N_7938,N_7795);
nand U8224 (N_8224,N_7883,N_7811);
nor U8225 (N_8225,N_7924,N_7991);
xnor U8226 (N_8226,N_7902,N_7851);
nand U8227 (N_8227,N_7802,N_7797);
or U8228 (N_8228,N_7946,N_7938);
xor U8229 (N_8229,N_7782,N_7873);
and U8230 (N_8230,N_7984,N_7790);
and U8231 (N_8231,N_7766,N_7974);
or U8232 (N_8232,N_7973,N_7922);
nor U8233 (N_8233,N_7830,N_7985);
xor U8234 (N_8234,N_7883,N_7788);
nand U8235 (N_8235,N_7776,N_7770);
and U8236 (N_8236,N_7941,N_7790);
or U8237 (N_8237,N_7925,N_7990);
xnor U8238 (N_8238,N_7775,N_7876);
xor U8239 (N_8239,N_7975,N_7786);
nor U8240 (N_8240,N_7777,N_7808);
and U8241 (N_8241,N_7935,N_7821);
nand U8242 (N_8242,N_7923,N_7920);
xor U8243 (N_8243,N_7757,N_7937);
nand U8244 (N_8244,N_7988,N_7903);
xnor U8245 (N_8245,N_7953,N_7815);
nor U8246 (N_8246,N_7916,N_7796);
xor U8247 (N_8247,N_7913,N_7887);
nor U8248 (N_8248,N_7857,N_7787);
nor U8249 (N_8249,N_7833,N_7805);
nand U8250 (N_8250,N_8062,N_8016);
and U8251 (N_8251,N_8012,N_8236);
and U8252 (N_8252,N_8222,N_8014);
nand U8253 (N_8253,N_8110,N_8146);
and U8254 (N_8254,N_8203,N_8249);
nor U8255 (N_8255,N_8165,N_8172);
nor U8256 (N_8256,N_8247,N_8186);
or U8257 (N_8257,N_8230,N_8160);
nand U8258 (N_8258,N_8064,N_8041);
nand U8259 (N_8259,N_8215,N_8117);
nand U8260 (N_8260,N_8218,N_8109);
nor U8261 (N_8261,N_8126,N_8105);
nand U8262 (N_8262,N_8031,N_8025);
xnor U8263 (N_8263,N_8161,N_8189);
nand U8264 (N_8264,N_8140,N_8211);
xnor U8265 (N_8265,N_8106,N_8077);
or U8266 (N_8266,N_8086,N_8131);
xnor U8267 (N_8267,N_8061,N_8089);
nor U8268 (N_8268,N_8133,N_8036);
xor U8269 (N_8269,N_8214,N_8123);
or U8270 (N_8270,N_8134,N_8093);
or U8271 (N_8271,N_8150,N_8038);
nand U8272 (N_8272,N_8095,N_8141);
nand U8273 (N_8273,N_8022,N_8159);
nand U8274 (N_8274,N_8180,N_8166);
nand U8275 (N_8275,N_8048,N_8034);
or U8276 (N_8276,N_8010,N_8020);
and U8277 (N_8277,N_8050,N_8137);
nand U8278 (N_8278,N_8130,N_8055);
or U8279 (N_8279,N_8081,N_8088);
and U8280 (N_8280,N_8018,N_8071);
nor U8281 (N_8281,N_8009,N_8212);
nor U8282 (N_8282,N_8181,N_8192);
and U8283 (N_8283,N_8128,N_8051);
nor U8284 (N_8284,N_8135,N_8239);
nor U8285 (N_8285,N_8224,N_8188);
nor U8286 (N_8286,N_8007,N_8175);
nor U8287 (N_8287,N_8210,N_8205);
nor U8288 (N_8288,N_8248,N_8138);
nor U8289 (N_8289,N_8111,N_8120);
nor U8290 (N_8290,N_8059,N_8001);
nand U8291 (N_8291,N_8094,N_8057);
or U8292 (N_8292,N_8082,N_8080);
and U8293 (N_8293,N_8087,N_8127);
xnor U8294 (N_8294,N_8201,N_8092);
xnor U8295 (N_8295,N_8073,N_8169);
and U8296 (N_8296,N_8244,N_8151);
xnor U8297 (N_8297,N_8090,N_8200);
or U8298 (N_8298,N_8220,N_8155);
or U8299 (N_8299,N_8074,N_8217);
xnor U8300 (N_8300,N_8047,N_8216);
and U8301 (N_8301,N_8191,N_8079);
and U8302 (N_8302,N_8174,N_8225);
nand U8303 (N_8303,N_8043,N_8167);
nor U8304 (N_8304,N_8008,N_8119);
xor U8305 (N_8305,N_8037,N_8237);
xor U8306 (N_8306,N_8234,N_8058);
nand U8307 (N_8307,N_8164,N_8158);
nor U8308 (N_8308,N_8195,N_8013);
and U8309 (N_8309,N_8136,N_8084);
xor U8310 (N_8310,N_8170,N_8207);
xnor U8311 (N_8311,N_8149,N_8070);
and U8312 (N_8312,N_8091,N_8098);
xor U8313 (N_8313,N_8190,N_8102);
or U8314 (N_8314,N_8024,N_8197);
xnor U8315 (N_8315,N_8227,N_8011);
or U8316 (N_8316,N_8053,N_8046);
nor U8317 (N_8317,N_8017,N_8000);
nand U8318 (N_8318,N_8152,N_8100);
nor U8319 (N_8319,N_8142,N_8107);
nor U8320 (N_8320,N_8063,N_8246);
or U8321 (N_8321,N_8231,N_8209);
or U8322 (N_8322,N_8067,N_8101);
and U8323 (N_8323,N_8033,N_8068);
nand U8324 (N_8324,N_8039,N_8143);
xnor U8325 (N_8325,N_8085,N_8173);
nand U8326 (N_8326,N_8183,N_8005);
or U8327 (N_8327,N_8199,N_8006);
xnor U8328 (N_8328,N_8178,N_8238);
xor U8329 (N_8329,N_8213,N_8066);
or U8330 (N_8330,N_8121,N_8103);
and U8331 (N_8331,N_8198,N_8153);
and U8332 (N_8332,N_8196,N_8240);
nor U8333 (N_8333,N_8163,N_8118);
nor U8334 (N_8334,N_8054,N_8023);
xor U8335 (N_8335,N_8148,N_8113);
or U8336 (N_8336,N_8122,N_8182);
or U8337 (N_8337,N_8096,N_8108);
and U8338 (N_8338,N_8147,N_8114);
and U8339 (N_8339,N_8132,N_8056);
nor U8340 (N_8340,N_8221,N_8243);
nor U8341 (N_8341,N_8002,N_8029);
and U8342 (N_8342,N_8219,N_8003);
or U8343 (N_8343,N_8226,N_8116);
or U8344 (N_8344,N_8233,N_8099);
nand U8345 (N_8345,N_8245,N_8179);
or U8346 (N_8346,N_8028,N_8075);
nand U8347 (N_8347,N_8242,N_8019);
xnor U8348 (N_8348,N_8078,N_8194);
or U8349 (N_8349,N_8241,N_8144);
xor U8350 (N_8350,N_8115,N_8139);
nor U8351 (N_8351,N_8223,N_8045);
or U8352 (N_8352,N_8156,N_8044);
and U8353 (N_8353,N_8021,N_8032);
nand U8354 (N_8354,N_8228,N_8168);
nand U8355 (N_8355,N_8124,N_8027);
or U8356 (N_8356,N_8040,N_8177);
nand U8357 (N_8357,N_8026,N_8112);
nor U8358 (N_8358,N_8185,N_8235);
nand U8359 (N_8359,N_8076,N_8052);
xor U8360 (N_8360,N_8104,N_8208);
nor U8361 (N_8361,N_8229,N_8065);
xnor U8362 (N_8362,N_8125,N_8035);
nor U8363 (N_8363,N_8145,N_8193);
nand U8364 (N_8364,N_8184,N_8157);
and U8365 (N_8365,N_8202,N_8069);
nand U8366 (N_8366,N_8083,N_8206);
nor U8367 (N_8367,N_8004,N_8176);
and U8368 (N_8368,N_8049,N_8171);
nand U8369 (N_8369,N_8154,N_8097);
nor U8370 (N_8370,N_8042,N_8129);
nor U8371 (N_8371,N_8015,N_8162);
nand U8372 (N_8372,N_8187,N_8204);
nand U8373 (N_8373,N_8030,N_8060);
and U8374 (N_8374,N_8232,N_8072);
xnor U8375 (N_8375,N_8140,N_8117);
nand U8376 (N_8376,N_8004,N_8238);
or U8377 (N_8377,N_8051,N_8037);
and U8378 (N_8378,N_8204,N_8020);
and U8379 (N_8379,N_8162,N_8185);
nor U8380 (N_8380,N_8184,N_8230);
and U8381 (N_8381,N_8007,N_8038);
or U8382 (N_8382,N_8038,N_8196);
xnor U8383 (N_8383,N_8102,N_8116);
or U8384 (N_8384,N_8065,N_8179);
xnor U8385 (N_8385,N_8097,N_8000);
or U8386 (N_8386,N_8062,N_8097);
xor U8387 (N_8387,N_8205,N_8045);
xnor U8388 (N_8388,N_8145,N_8222);
or U8389 (N_8389,N_8165,N_8115);
or U8390 (N_8390,N_8048,N_8064);
nand U8391 (N_8391,N_8231,N_8193);
nor U8392 (N_8392,N_8246,N_8151);
nand U8393 (N_8393,N_8063,N_8092);
xor U8394 (N_8394,N_8020,N_8106);
nor U8395 (N_8395,N_8147,N_8215);
or U8396 (N_8396,N_8158,N_8081);
nand U8397 (N_8397,N_8150,N_8216);
or U8398 (N_8398,N_8002,N_8154);
or U8399 (N_8399,N_8072,N_8027);
nor U8400 (N_8400,N_8097,N_8151);
nor U8401 (N_8401,N_8143,N_8053);
nor U8402 (N_8402,N_8240,N_8062);
and U8403 (N_8403,N_8009,N_8184);
and U8404 (N_8404,N_8016,N_8024);
nor U8405 (N_8405,N_8139,N_8100);
and U8406 (N_8406,N_8092,N_8193);
or U8407 (N_8407,N_8119,N_8174);
nand U8408 (N_8408,N_8005,N_8114);
nor U8409 (N_8409,N_8078,N_8212);
and U8410 (N_8410,N_8081,N_8023);
or U8411 (N_8411,N_8007,N_8212);
or U8412 (N_8412,N_8144,N_8174);
nand U8413 (N_8413,N_8198,N_8066);
or U8414 (N_8414,N_8038,N_8057);
nand U8415 (N_8415,N_8209,N_8133);
nor U8416 (N_8416,N_8067,N_8001);
nand U8417 (N_8417,N_8210,N_8191);
and U8418 (N_8418,N_8047,N_8086);
xor U8419 (N_8419,N_8035,N_8113);
and U8420 (N_8420,N_8172,N_8187);
nand U8421 (N_8421,N_8042,N_8010);
nand U8422 (N_8422,N_8060,N_8092);
nor U8423 (N_8423,N_8034,N_8166);
nor U8424 (N_8424,N_8181,N_8089);
and U8425 (N_8425,N_8086,N_8197);
nand U8426 (N_8426,N_8104,N_8002);
nor U8427 (N_8427,N_8164,N_8044);
and U8428 (N_8428,N_8214,N_8109);
nand U8429 (N_8429,N_8133,N_8005);
nand U8430 (N_8430,N_8103,N_8054);
and U8431 (N_8431,N_8016,N_8063);
nor U8432 (N_8432,N_8176,N_8049);
or U8433 (N_8433,N_8217,N_8246);
and U8434 (N_8434,N_8169,N_8181);
and U8435 (N_8435,N_8174,N_8198);
or U8436 (N_8436,N_8173,N_8034);
or U8437 (N_8437,N_8210,N_8033);
and U8438 (N_8438,N_8008,N_8249);
nand U8439 (N_8439,N_8008,N_8093);
or U8440 (N_8440,N_8153,N_8137);
or U8441 (N_8441,N_8100,N_8044);
nand U8442 (N_8442,N_8147,N_8000);
nor U8443 (N_8443,N_8118,N_8039);
nor U8444 (N_8444,N_8049,N_8027);
xor U8445 (N_8445,N_8207,N_8139);
nand U8446 (N_8446,N_8242,N_8031);
nor U8447 (N_8447,N_8129,N_8049);
xnor U8448 (N_8448,N_8034,N_8194);
nor U8449 (N_8449,N_8012,N_8082);
or U8450 (N_8450,N_8065,N_8049);
nand U8451 (N_8451,N_8211,N_8019);
nor U8452 (N_8452,N_8035,N_8108);
or U8453 (N_8453,N_8024,N_8096);
xnor U8454 (N_8454,N_8135,N_8212);
xor U8455 (N_8455,N_8217,N_8037);
xnor U8456 (N_8456,N_8221,N_8174);
or U8457 (N_8457,N_8057,N_8018);
nor U8458 (N_8458,N_8063,N_8062);
nor U8459 (N_8459,N_8172,N_8204);
xnor U8460 (N_8460,N_8235,N_8152);
or U8461 (N_8461,N_8160,N_8106);
and U8462 (N_8462,N_8105,N_8115);
nand U8463 (N_8463,N_8037,N_8092);
nor U8464 (N_8464,N_8213,N_8033);
xor U8465 (N_8465,N_8144,N_8086);
nand U8466 (N_8466,N_8016,N_8107);
and U8467 (N_8467,N_8194,N_8180);
nor U8468 (N_8468,N_8037,N_8210);
nor U8469 (N_8469,N_8215,N_8216);
nand U8470 (N_8470,N_8206,N_8152);
nand U8471 (N_8471,N_8058,N_8108);
xor U8472 (N_8472,N_8145,N_8122);
nor U8473 (N_8473,N_8036,N_8063);
nand U8474 (N_8474,N_8170,N_8153);
and U8475 (N_8475,N_8017,N_8025);
nor U8476 (N_8476,N_8233,N_8057);
nor U8477 (N_8477,N_8087,N_8016);
and U8478 (N_8478,N_8136,N_8193);
xnor U8479 (N_8479,N_8203,N_8201);
and U8480 (N_8480,N_8114,N_8038);
nand U8481 (N_8481,N_8132,N_8009);
and U8482 (N_8482,N_8154,N_8133);
and U8483 (N_8483,N_8145,N_8207);
and U8484 (N_8484,N_8035,N_8249);
nor U8485 (N_8485,N_8001,N_8109);
nand U8486 (N_8486,N_8087,N_8140);
nand U8487 (N_8487,N_8082,N_8001);
and U8488 (N_8488,N_8033,N_8112);
nand U8489 (N_8489,N_8061,N_8022);
nand U8490 (N_8490,N_8117,N_8179);
nand U8491 (N_8491,N_8019,N_8007);
xnor U8492 (N_8492,N_8194,N_8240);
xnor U8493 (N_8493,N_8076,N_8202);
nand U8494 (N_8494,N_8207,N_8094);
xor U8495 (N_8495,N_8130,N_8082);
nor U8496 (N_8496,N_8018,N_8148);
nand U8497 (N_8497,N_8023,N_8009);
xnor U8498 (N_8498,N_8042,N_8214);
xor U8499 (N_8499,N_8070,N_8026);
nor U8500 (N_8500,N_8290,N_8470);
nand U8501 (N_8501,N_8458,N_8253);
nand U8502 (N_8502,N_8269,N_8292);
and U8503 (N_8503,N_8284,N_8319);
and U8504 (N_8504,N_8429,N_8497);
nor U8505 (N_8505,N_8341,N_8484);
nor U8506 (N_8506,N_8279,N_8351);
nand U8507 (N_8507,N_8428,N_8260);
and U8508 (N_8508,N_8337,N_8409);
or U8509 (N_8509,N_8286,N_8391);
nand U8510 (N_8510,N_8482,N_8465);
or U8511 (N_8511,N_8311,N_8339);
nand U8512 (N_8512,N_8417,N_8298);
nor U8513 (N_8513,N_8464,N_8383);
nand U8514 (N_8514,N_8262,N_8375);
and U8515 (N_8515,N_8338,N_8363);
xnor U8516 (N_8516,N_8282,N_8435);
nor U8517 (N_8517,N_8361,N_8291);
and U8518 (N_8518,N_8461,N_8350);
xor U8519 (N_8519,N_8400,N_8296);
xor U8520 (N_8520,N_8270,N_8408);
or U8521 (N_8521,N_8432,N_8295);
nor U8522 (N_8522,N_8475,N_8445);
or U8523 (N_8523,N_8425,N_8406);
xnor U8524 (N_8524,N_8380,N_8471);
or U8525 (N_8525,N_8437,N_8402);
nand U8526 (N_8526,N_8394,N_8301);
xor U8527 (N_8527,N_8404,N_8343);
nand U8528 (N_8528,N_8362,N_8324);
nand U8529 (N_8529,N_8422,N_8359);
nand U8530 (N_8530,N_8313,N_8459);
or U8531 (N_8531,N_8411,N_8345);
or U8532 (N_8532,N_8336,N_8306);
nand U8533 (N_8533,N_8352,N_8257);
and U8534 (N_8534,N_8367,N_8259);
or U8535 (N_8535,N_8283,N_8430);
xnor U8536 (N_8536,N_8423,N_8381);
or U8537 (N_8537,N_8302,N_8366);
nand U8538 (N_8538,N_8491,N_8390);
xor U8539 (N_8539,N_8316,N_8255);
nor U8540 (N_8540,N_8440,N_8405);
nand U8541 (N_8541,N_8307,N_8321);
nor U8542 (N_8542,N_8463,N_8309);
or U8543 (N_8543,N_8310,N_8261);
or U8544 (N_8544,N_8370,N_8293);
nand U8545 (N_8545,N_8489,N_8444);
or U8546 (N_8546,N_8399,N_8469);
and U8547 (N_8547,N_8446,N_8396);
and U8548 (N_8548,N_8304,N_8377);
or U8549 (N_8549,N_8490,N_8481);
and U8550 (N_8550,N_8300,N_8492);
nand U8551 (N_8551,N_8340,N_8384);
or U8552 (N_8552,N_8267,N_8467);
and U8553 (N_8553,N_8498,N_8280);
nor U8554 (N_8554,N_8397,N_8288);
nand U8555 (N_8555,N_8483,N_8456);
or U8556 (N_8556,N_8389,N_8407);
nor U8557 (N_8557,N_8495,N_8438);
xnor U8558 (N_8558,N_8276,N_8289);
nor U8559 (N_8559,N_8424,N_8305);
or U8560 (N_8560,N_8354,N_8335);
nor U8561 (N_8561,N_8256,N_8455);
xnor U8562 (N_8562,N_8254,N_8393);
and U8563 (N_8563,N_8453,N_8488);
nor U8564 (N_8564,N_8472,N_8251);
nand U8565 (N_8565,N_8285,N_8374);
nor U8566 (N_8566,N_8266,N_8487);
nor U8567 (N_8567,N_8353,N_8378);
or U8568 (N_8568,N_8330,N_8454);
xor U8569 (N_8569,N_8348,N_8312);
nand U8570 (N_8570,N_8272,N_8443);
and U8571 (N_8571,N_8371,N_8277);
nand U8572 (N_8572,N_8358,N_8449);
or U8573 (N_8573,N_8331,N_8476);
xor U8574 (N_8574,N_8480,N_8431);
nand U8575 (N_8575,N_8379,N_8264);
nand U8576 (N_8576,N_8332,N_8436);
and U8577 (N_8577,N_8479,N_8442);
nor U8578 (N_8578,N_8448,N_8493);
nor U8579 (N_8579,N_8368,N_8252);
nor U8580 (N_8580,N_8323,N_8486);
and U8581 (N_8581,N_8496,N_8357);
or U8582 (N_8582,N_8320,N_8268);
or U8583 (N_8583,N_8403,N_8314);
nor U8584 (N_8584,N_8326,N_8473);
or U8585 (N_8585,N_8439,N_8494);
nor U8586 (N_8586,N_8278,N_8434);
xor U8587 (N_8587,N_8369,N_8395);
nand U8588 (N_8588,N_8349,N_8274);
nor U8589 (N_8589,N_8451,N_8347);
xnor U8590 (N_8590,N_8426,N_8328);
xnor U8591 (N_8591,N_8478,N_8364);
and U8592 (N_8592,N_8466,N_8388);
nor U8593 (N_8593,N_8299,N_8452);
nand U8594 (N_8594,N_8499,N_8382);
nor U8595 (N_8595,N_8346,N_8412);
and U8596 (N_8596,N_8271,N_8329);
or U8597 (N_8597,N_8477,N_8457);
nand U8598 (N_8598,N_8419,N_8474);
and U8599 (N_8599,N_8485,N_8421);
nand U8600 (N_8600,N_8258,N_8373);
nor U8601 (N_8601,N_8294,N_8297);
and U8602 (N_8602,N_8355,N_8325);
or U8603 (N_8603,N_8334,N_8398);
and U8604 (N_8604,N_8250,N_8418);
nand U8605 (N_8605,N_8460,N_8327);
nand U8606 (N_8606,N_8287,N_8308);
and U8607 (N_8607,N_8416,N_8365);
xnor U8608 (N_8608,N_8385,N_8387);
nor U8609 (N_8609,N_8303,N_8433);
xnor U8610 (N_8610,N_8441,N_8275);
or U8611 (N_8611,N_8392,N_8413);
xnor U8612 (N_8612,N_8427,N_8386);
nand U8613 (N_8613,N_8317,N_8356);
or U8614 (N_8614,N_8333,N_8344);
or U8615 (N_8615,N_8420,N_8410);
xnor U8616 (N_8616,N_8415,N_8376);
nor U8617 (N_8617,N_8462,N_8263);
or U8618 (N_8618,N_8450,N_8322);
or U8619 (N_8619,N_8447,N_8315);
nand U8620 (N_8620,N_8401,N_8468);
nand U8621 (N_8621,N_8360,N_8265);
and U8622 (N_8622,N_8372,N_8318);
xor U8623 (N_8623,N_8281,N_8273);
or U8624 (N_8624,N_8414,N_8342);
nor U8625 (N_8625,N_8280,N_8459);
or U8626 (N_8626,N_8447,N_8394);
nor U8627 (N_8627,N_8396,N_8463);
xnor U8628 (N_8628,N_8416,N_8393);
xor U8629 (N_8629,N_8352,N_8364);
and U8630 (N_8630,N_8327,N_8346);
and U8631 (N_8631,N_8322,N_8401);
xor U8632 (N_8632,N_8287,N_8286);
or U8633 (N_8633,N_8341,N_8287);
or U8634 (N_8634,N_8402,N_8256);
xnor U8635 (N_8635,N_8420,N_8461);
or U8636 (N_8636,N_8351,N_8386);
nand U8637 (N_8637,N_8425,N_8287);
nand U8638 (N_8638,N_8281,N_8313);
or U8639 (N_8639,N_8456,N_8323);
or U8640 (N_8640,N_8469,N_8316);
nand U8641 (N_8641,N_8457,N_8345);
and U8642 (N_8642,N_8374,N_8375);
nand U8643 (N_8643,N_8363,N_8281);
nand U8644 (N_8644,N_8458,N_8368);
xnor U8645 (N_8645,N_8495,N_8250);
nand U8646 (N_8646,N_8340,N_8493);
and U8647 (N_8647,N_8276,N_8461);
or U8648 (N_8648,N_8283,N_8349);
nor U8649 (N_8649,N_8360,N_8482);
nor U8650 (N_8650,N_8468,N_8424);
and U8651 (N_8651,N_8298,N_8270);
or U8652 (N_8652,N_8282,N_8256);
xnor U8653 (N_8653,N_8486,N_8427);
nor U8654 (N_8654,N_8332,N_8489);
and U8655 (N_8655,N_8484,N_8401);
nand U8656 (N_8656,N_8263,N_8369);
xnor U8657 (N_8657,N_8350,N_8438);
xor U8658 (N_8658,N_8316,N_8337);
xor U8659 (N_8659,N_8351,N_8422);
xor U8660 (N_8660,N_8384,N_8403);
xnor U8661 (N_8661,N_8295,N_8259);
or U8662 (N_8662,N_8334,N_8449);
nand U8663 (N_8663,N_8352,N_8467);
or U8664 (N_8664,N_8444,N_8343);
xor U8665 (N_8665,N_8281,N_8348);
xnor U8666 (N_8666,N_8387,N_8494);
nand U8667 (N_8667,N_8444,N_8267);
or U8668 (N_8668,N_8421,N_8381);
or U8669 (N_8669,N_8473,N_8399);
or U8670 (N_8670,N_8307,N_8301);
nand U8671 (N_8671,N_8451,N_8497);
and U8672 (N_8672,N_8304,N_8480);
and U8673 (N_8673,N_8265,N_8272);
nand U8674 (N_8674,N_8253,N_8323);
nor U8675 (N_8675,N_8272,N_8274);
nor U8676 (N_8676,N_8447,N_8267);
and U8677 (N_8677,N_8277,N_8343);
nand U8678 (N_8678,N_8274,N_8307);
or U8679 (N_8679,N_8296,N_8364);
and U8680 (N_8680,N_8490,N_8324);
and U8681 (N_8681,N_8332,N_8337);
nand U8682 (N_8682,N_8273,N_8393);
nand U8683 (N_8683,N_8395,N_8472);
or U8684 (N_8684,N_8329,N_8383);
xnor U8685 (N_8685,N_8323,N_8321);
and U8686 (N_8686,N_8409,N_8440);
or U8687 (N_8687,N_8474,N_8329);
and U8688 (N_8688,N_8489,N_8430);
nor U8689 (N_8689,N_8498,N_8457);
nand U8690 (N_8690,N_8483,N_8450);
and U8691 (N_8691,N_8334,N_8442);
and U8692 (N_8692,N_8421,N_8309);
xnor U8693 (N_8693,N_8455,N_8381);
and U8694 (N_8694,N_8450,N_8488);
or U8695 (N_8695,N_8365,N_8335);
or U8696 (N_8696,N_8281,N_8365);
or U8697 (N_8697,N_8254,N_8423);
nor U8698 (N_8698,N_8350,N_8382);
nor U8699 (N_8699,N_8350,N_8325);
nor U8700 (N_8700,N_8484,N_8374);
nand U8701 (N_8701,N_8441,N_8322);
or U8702 (N_8702,N_8345,N_8396);
nand U8703 (N_8703,N_8477,N_8400);
or U8704 (N_8704,N_8439,N_8459);
nor U8705 (N_8705,N_8302,N_8420);
and U8706 (N_8706,N_8290,N_8351);
and U8707 (N_8707,N_8424,N_8278);
nor U8708 (N_8708,N_8447,N_8287);
or U8709 (N_8709,N_8390,N_8471);
or U8710 (N_8710,N_8417,N_8288);
nor U8711 (N_8711,N_8271,N_8429);
and U8712 (N_8712,N_8458,N_8468);
xor U8713 (N_8713,N_8399,N_8302);
nand U8714 (N_8714,N_8329,N_8473);
or U8715 (N_8715,N_8491,N_8260);
nand U8716 (N_8716,N_8490,N_8355);
or U8717 (N_8717,N_8410,N_8393);
nand U8718 (N_8718,N_8398,N_8474);
nor U8719 (N_8719,N_8486,N_8301);
or U8720 (N_8720,N_8431,N_8386);
nor U8721 (N_8721,N_8344,N_8395);
and U8722 (N_8722,N_8280,N_8250);
or U8723 (N_8723,N_8494,N_8488);
nor U8724 (N_8724,N_8382,N_8395);
xnor U8725 (N_8725,N_8372,N_8259);
or U8726 (N_8726,N_8367,N_8387);
nor U8727 (N_8727,N_8336,N_8361);
xor U8728 (N_8728,N_8305,N_8434);
nor U8729 (N_8729,N_8482,N_8485);
xor U8730 (N_8730,N_8260,N_8326);
nand U8731 (N_8731,N_8319,N_8376);
nor U8732 (N_8732,N_8496,N_8332);
nor U8733 (N_8733,N_8474,N_8468);
nand U8734 (N_8734,N_8485,N_8306);
nor U8735 (N_8735,N_8258,N_8431);
and U8736 (N_8736,N_8253,N_8328);
and U8737 (N_8737,N_8391,N_8269);
nor U8738 (N_8738,N_8414,N_8355);
nor U8739 (N_8739,N_8394,N_8488);
and U8740 (N_8740,N_8271,N_8316);
or U8741 (N_8741,N_8390,N_8444);
nor U8742 (N_8742,N_8476,N_8491);
or U8743 (N_8743,N_8484,N_8290);
nor U8744 (N_8744,N_8333,N_8391);
and U8745 (N_8745,N_8381,N_8410);
xnor U8746 (N_8746,N_8485,N_8481);
nor U8747 (N_8747,N_8251,N_8445);
nor U8748 (N_8748,N_8315,N_8394);
nand U8749 (N_8749,N_8326,N_8457);
nand U8750 (N_8750,N_8658,N_8518);
or U8751 (N_8751,N_8559,N_8701);
xor U8752 (N_8752,N_8500,N_8536);
xor U8753 (N_8753,N_8625,N_8671);
or U8754 (N_8754,N_8520,N_8618);
or U8755 (N_8755,N_8713,N_8655);
xnor U8756 (N_8756,N_8545,N_8634);
and U8757 (N_8757,N_8633,N_8630);
xor U8758 (N_8758,N_8694,N_8653);
or U8759 (N_8759,N_8531,N_8605);
nand U8760 (N_8760,N_8728,N_8506);
nand U8761 (N_8761,N_8639,N_8687);
or U8762 (N_8762,N_8538,N_8646);
nand U8763 (N_8763,N_8729,N_8503);
nor U8764 (N_8764,N_8548,N_8534);
xnor U8765 (N_8765,N_8617,N_8711);
nand U8766 (N_8766,N_8680,N_8693);
nand U8767 (N_8767,N_8684,N_8527);
nand U8768 (N_8768,N_8681,N_8741);
nand U8769 (N_8769,N_8676,N_8575);
nor U8770 (N_8770,N_8674,N_8665);
and U8771 (N_8771,N_8673,N_8517);
or U8772 (N_8772,N_8513,N_8696);
or U8773 (N_8773,N_8567,N_8542);
and U8774 (N_8774,N_8648,N_8739);
or U8775 (N_8775,N_8704,N_8710);
nand U8776 (N_8776,N_8734,N_8637);
nor U8777 (N_8777,N_8510,N_8712);
or U8778 (N_8778,N_8582,N_8622);
xor U8779 (N_8779,N_8533,N_8511);
or U8780 (N_8780,N_8677,N_8643);
xnor U8781 (N_8781,N_8656,N_8579);
nor U8782 (N_8782,N_8565,N_8636);
and U8783 (N_8783,N_8547,N_8661);
nor U8784 (N_8784,N_8612,N_8587);
nand U8785 (N_8785,N_8716,N_8645);
and U8786 (N_8786,N_8599,N_8718);
nor U8787 (N_8787,N_8574,N_8621);
xor U8788 (N_8788,N_8686,N_8738);
and U8789 (N_8789,N_8535,N_8679);
and U8790 (N_8790,N_8588,N_8737);
nand U8791 (N_8791,N_8508,N_8723);
or U8792 (N_8792,N_8721,N_8589);
xor U8793 (N_8793,N_8744,N_8730);
or U8794 (N_8794,N_8584,N_8551);
nand U8795 (N_8795,N_8600,N_8539);
xor U8796 (N_8796,N_8745,N_8546);
nand U8797 (N_8797,N_8735,N_8623);
or U8798 (N_8798,N_8550,N_8652);
or U8799 (N_8799,N_8719,N_8613);
xnor U8800 (N_8800,N_8557,N_8591);
xor U8801 (N_8801,N_8660,N_8705);
nand U8802 (N_8802,N_8644,N_8666);
and U8803 (N_8803,N_8595,N_8543);
nor U8804 (N_8804,N_8553,N_8561);
and U8805 (N_8805,N_8736,N_8624);
and U8806 (N_8806,N_8727,N_8523);
nand U8807 (N_8807,N_8628,N_8558);
xnor U8808 (N_8808,N_8609,N_8732);
or U8809 (N_8809,N_8749,N_8702);
nor U8810 (N_8810,N_8649,N_8549);
xnor U8811 (N_8811,N_8554,N_8640);
or U8812 (N_8812,N_8703,N_8733);
nor U8813 (N_8813,N_8602,N_8583);
xnor U8814 (N_8814,N_8578,N_8570);
nand U8815 (N_8815,N_8626,N_8509);
and U8816 (N_8816,N_8743,N_8678);
or U8817 (N_8817,N_8581,N_8715);
nand U8818 (N_8818,N_8706,N_8585);
xnor U8819 (N_8819,N_8619,N_8638);
and U8820 (N_8820,N_8627,N_8620);
and U8821 (N_8821,N_8748,N_8651);
or U8822 (N_8822,N_8530,N_8522);
xnor U8823 (N_8823,N_8722,N_8708);
xnor U8824 (N_8824,N_8515,N_8695);
nand U8825 (N_8825,N_8501,N_8566);
and U8826 (N_8826,N_8675,N_8569);
xor U8827 (N_8827,N_8593,N_8725);
nand U8828 (N_8828,N_8664,N_8699);
and U8829 (N_8829,N_8720,N_8629);
xor U8830 (N_8830,N_8608,N_8726);
nor U8831 (N_8831,N_8601,N_8592);
xor U8832 (N_8832,N_8697,N_8504);
and U8833 (N_8833,N_8717,N_8632);
xnor U8834 (N_8834,N_8505,N_8709);
xnor U8835 (N_8835,N_8514,N_8747);
xor U8836 (N_8836,N_8586,N_8685);
nand U8837 (N_8837,N_8532,N_8663);
xor U8838 (N_8838,N_8576,N_8683);
nand U8839 (N_8839,N_8698,N_8654);
nor U8840 (N_8840,N_8571,N_8552);
or U8841 (N_8841,N_8541,N_8596);
nand U8842 (N_8842,N_8642,N_8690);
xnor U8843 (N_8843,N_8597,N_8573);
and U8844 (N_8844,N_8610,N_8604);
and U8845 (N_8845,N_8691,N_8672);
nor U8846 (N_8846,N_8714,N_8521);
nand U8847 (N_8847,N_8635,N_8537);
and U8848 (N_8848,N_8700,N_8659);
and U8849 (N_8849,N_8615,N_8682);
or U8850 (N_8850,N_8540,N_8502);
and U8851 (N_8851,N_8526,N_8507);
and U8852 (N_8852,N_8603,N_8562);
or U8853 (N_8853,N_8647,N_8524);
nand U8854 (N_8854,N_8731,N_8555);
xnor U8855 (N_8855,N_8564,N_8641);
or U8856 (N_8856,N_8740,N_8657);
nand U8857 (N_8857,N_8631,N_8616);
or U8858 (N_8858,N_8742,N_8650);
and U8859 (N_8859,N_8667,N_8670);
nand U8860 (N_8860,N_8529,N_8611);
nand U8861 (N_8861,N_8607,N_8568);
xor U8862 (N_8862,N_8662,N_8563);
and U8863 (N_8863,N_8580,N_8556);
xor U8864 (N_8864,N_8519,N_8614);
and U8865 (N_8865,N_8512,N_8572);
nor U8866 (N_8866,N_8707,N_8724);
and U8867 (N_8867,N_8544,N_8525);
or U8868 (N_8868,N_8528,N_8746);
nand U8869 (N_8869,N_8598,N_8594);
nor U8870 (N_8870,N_8590,N_8606);
nor U8871 (N_8871,N_8692,N_8669);
and U8872 (N_8872,N_8577,N_8668);
or U8873 (N_8873,N_8516,N_8689);
nor U8874 (N_8874,N_8688,N_8560);
nand U8875 (N_8875,N_8697,N_8514);
or U8876 (N_8876,N_8711,N_8504);
nand U8877 (N_8877,N_8512,N_8684);
and U8878 (N_8878,N_8728,N_8529);
or U8879 (N_8879,N_8601,N_8501);
nor U8880 (N_8880,N_8739,N_8554);
nand U8881 (N_8881,N_8602,N_8562);
nand U8882 (N_8882,N_8746,N_8530);
nor U8883 (N_8883,N_8507,N_8580);
xnor U8884 (N_8884,N_8718,N_8637);
nand U8885 (N_8885,N_8573,N_8723);
xor U8886 (N_8886,N_8700,N_8515);
nor U8887 (N_8887,N_8521,N_8612);
and U8888 (N_8888,N_8518,N_8530);
nor U8889 (N_8889,N_8547,N_8586);
nand U8890 (N_8890,N_8729,N_8660);
nand U8891 (N_8891,N_8710,N_8695);
nand U8892 (N_8892,N_8562,N_8613);
xor U8893 (N_8893,N_8736,N_8703);
and U8894 (N_8894,N_8632,N_8608);
and U8895 (N_8895,N_8685,N_8508);
or U8896 (N_8896,N_8729,N_8556);
and U8897 (N_8897,N_8619,N_8594);
nand U8898 (N_8898,N_8503,N_8618);
xor U8899 (N_8899,N_8558,N_8634);
xor U8900 (N_8900,N_8600,N_8587);
nor U8901 (N_8901,N_8696,N_8624);
nand U8902 (N_8902,N_8687,N_8538);
nand U8903 (N_8903,N_8675,N_8576);
and U8904 (N_8904,N_8557,N_8570);
xnor U8905 (N_8905,N_8737,N_8623);
or U8906 (N_8906,N_8555,N_8583);
xor U8907 (N_8907,N_8551,N_8649);
nand U8908 (N_8908,N_8734,N_8615);
and U8909 (N_8909,N_8582,N_8719);
nor U8910 (N_8910,N_8505,N_8542);
nor U8911 (N_8911,N_8655,N_8606);
and U8912 (N_8912,N_8705,N_8516);
or U8913 (N_8913,N_8562,N_8660);
or U8914 (N_8914,N_8549,N_8713);
xor U8915 (N_8915,N_8596,N_8588);
or U8916 (N_8916,N_8708,N_8517);
xnor U8917 (N_8917,N_8655,N_8570);
and U8918 (N_8918,N_8528,N_8734);
nor U8919 (N_8919,N_8551,N_8581);
and U8920 (N_8920,N_8519,N_8691);
nand U8921 (N_8921,N_8579,N_8669);
or U8922 (N_8922,N_8540,N_8529);
nand U8923 (N_8923,N_8585,N_8730);
nor U8924 (N_8924,N_8563,N_8593);
nor U8925 (N_8925,N_8609,N_8720);
nand U8926 (N_8926,N_8642,N_8551);
or U8927 (N_8927,N_8518,N_8696);
nand U8928 (N_8928,N_8546,N_8686);
nor U8929 (N_8929,N_8560,N_8655);
or U8930 (N_8930,N_8677,N_8605);
or U8931 (N_8931,N_8717,N_8531);
and U8932 (N_8932,N_8700,N_8672);
nor U8933 (N_8933,N_8709,N_8686);
nand U8934 (N_8934,N_8725,N_8688);
nand U8935 (N_8935,N_8649,N_8658);
or U8936 (N_8936,N_8584,N_8720);
or U8937 (N_8937,N_8723,N_8528);
or U8938 (N_8938,N_8527,N_8641);
nor U8939 (N_8939,N_8689,N_8639);
xor U8940 (N_8940,N_8561,N_8634);
nand U8941 (N_8941,N_8602,N_8705);
xor U8942 (N_8942,N_8629,N_8730);
nand U8943 (N_8943,N_8611,N_8570);
nand U8944 (N_8944,N_8663,N_8569);
and U8945 (N_8945,N_8545,N_8614);
and U8946 (N_8946,N_8566,N_8608);
xnor U8947 (N_8947,N_8638,N_8622);
nand U8948 (N_8948,N_8570,N_8654);
and U8949 (N_8949,N_8556,N_8517);
or U8950 (N_8950,N_8736,N_8642);
or U8951 (N_8951,N_8703,N_8731);
or U8952 (N_8952,N_8529,N_8640);
and U8953 (N_8953,N_8739,N_8573);
xnor U8954 (N_8954,N_8659,N_8521);
xor U8955 (N_8955,N_8579,N_8520);
or U8956 (N_8956,N_8643,N_8685);
and U8957 (N_8957,N_8736,N_8622);
or U8958 (N_8958,N_8662,N_8527);
xor U8959 (N_8959,N_8593,N_8518);
or U8960 (N_8960,N_8627,N_8579);
and U8961 (N_8961,N_8672,N_8645);
xor U8962 (N_8962,N_8731,N_8514);
xnor U8963 (N_8963,N_8689,N_8733);
nand U8964 (N_8964,N_8577,N_8597);
xnor U8965 (N_8965,N_8570,N_8559);
nand U8966 (N_8966,N_8566,N_8543);
nor U8967 (N_8967,N_8649,N_8612);
xor U8968 (N_8968,N_8714,N_8677);
and U8969 (N_8969,N_8523,N_8648);
xnor U8970 (N_8970,N_8729,N_8740);
and U8971 (N_8971,N_8697,N_8575);
nor U8972 (N_8972,N_8704,N_8532);
xnor U8973 (N_8973,N_8667,N_8618);
nand U8974 (N_8974,N_8726,N_8616);
nand U8975 (N_8975,N_8692,N_8704);
nor U8976 (N_8976,N_8513,N_8739);
or U8977 (N_8977,N_8539,N_8725);
nor U8978 (N_8978,N_8669,N_8513);
xor U8979 (N_8979,N_8719,N_8635);
xnor U8980 (N_8980,N_8648,N_8696);
nor U8981 (N_8981,N_8577,N_8622);
nor U8982 (N_8982,N_8708,N_8539);
nor U8983 (N_8983,N_8643,N_8505);
nor U8984 (N_8984,N_8716,N_8736);
nor U8985 (N_8985,N_8737,N_8508);
nor U8986 (N_8986,N_8743,N_8663);
nand U8987 (N_8987,N_8503,N_8588);
nor U8988 (N_8988,N_8634,N_8697);
nand U8989 (N_8989,N_8721,N_8576);
nand U8990 (N_8990,N_8605,N_8712);
and U8991 (N_8991,N_8663,N_8713);
and U8992 (N_8992,N_8725,N_8534);
xnor U8993 (N_8993,N_8746,N_8579);
or U8994 (N_8994,N_8602,N_8701);
nand U8995 (N_8995,N_8723,N_8665);
or U8996 (N_8996,N_8596,N_8551);
or U8997 (N_8997,N_8548,N_8539);
nand U8998 (N_8998,N_8515,N_8676);
xnor U8999 (N_8999,N_8698,N_8681);
xnor U9000 (N_9000,N_8773,N_8999);
and U9001 (N_9001,N_8812,N_8863);
xor U9002 (N_9002,N_8894,N_8989);
xnor U9003 (N_9003,N_8798,N_8913);
or U9004 (N_9004,N_8957,N_8998);
nor U9005 (N_9005,N_8907,N_8800);
or U9006 (N_9006,N_8891,N_8853);
xnor U9007 (N_9007,N_8940,N_8946);
or U9008 (N_9008,N_8920,N_8987);
xor U9009 (N_9009,N_8779,N_8846);
and U9010 (N_9010,N_8844,N_8964);
and U9011 (N_9011,N_8758,N_8935);
and U9012 (N_9012,N_8971,N_8928);
xnor U9013 (N_9013,N_8823,N_8792);
and U9014 (N_9014,N_8807,N_8764);
nand U9015 (N_9015,N_8840,N_8910);
or U9016 (N_9016,N_8790,N_8967);
nor U9017 (N_9017,N_8917,N_8828);
nand U9018 (N_9018,N_8951,N_8939);
nand U9019 (N_9019,N_8919,N_8845);
or U9020 (N_9020,N_8995,N_8841);
nand U9021 (N_9021,N_8756,N_8769);
nand U9022 (N_9022,N_8912,N_8780);
and U9023 (N_9023,N_8821,N_8945);
and U9024 (N_9024,N_8778,N_8947);
nand U9025 (N_9025,N_8905,N_8753);
nand U9026 (N_9026,N_8864,N_8783);
xnor U9027 (N_9027,N_8897,N_8956);
xor U9028 (N_9028,N_8880,N_8752);
and U9029 (N_9029,N_8819,N_8761);
xnor U9030 (N_9030,N_8953,N_8930);
or U9031 (N_9031,N_8992,N_8958);
and U9032 (N_9032,N_8784,N_8826);
nor U9033 (N_9033,N_8899,N_8755);
and U9034 (N_9034,N_8955,N_8867);
nor U9035 (N_9035,N_8994,N_8911);
and U9036 (N_9036,N_8921,N_8815);
and U9037 (N_9037,N_8873,N_8776);
or U9038 (N_9038,N_8974,N_8789);
xor U9039 (N_9039,N_8916,N_8918);
nor U9040 (N_9040,N_8825,N_8952);
nor U9041 (N_9041,N_8996,N_8877);
or U9042 (N_9042,N_8962,N_8865);
xor U9043 (N_9043,N_8931,N_8885);
xnor U9044 (N_9044,N_8855,N_8811);
or U9045 (N_9045,N_8806,N_8791);
xor U9046 (N_9046,N_8925,N_8796);
or U9047 (N_9047,N_8858,N_8802);
or U9048 (N_9048,N_8793,N_8808);
and U9049 (N_9049,N_8878,N_8978);
and U9050 (N_9050,N_8927,N_8866);
and U9051 (N_9051,N_8856,N_8909);
nor U9052 (N_9052,N_8751,N_8852);
or U9053 (N_9053,N_8972,N_8850);
and U9054 (N_9054,N_8991,N_8861);
xnor U9055 (N_9055,N_8963,N_8810);
nor U9056 (N_9056,N_8893,N_8906);
xnor U9057 (N_9057,N_8805,N_8882);
and U9058 (N_9058,N_8914,N_8782);
and U9059 (N_9059,N_8981,N_8838);
and U9060 (N_9060,N_8997,N_8970);
and U9061 (N_9061,N_8944,N_8831);
and U9062 (N_9062,N_8879,N_8772);
nor U9063 (N_9063,N_8932,N_8869);
or U9064 (N_9064,N_8982,N_8874);
xnor U9065 (N_9065,N_8775,N_8872);
xor U9066 (N_9066,N_8993,N_8923);
xor U9067 (N_9067,N_8820,N_8943);
xnor U9068 (N_9068,N_8848,N_8937);
xor U9069 (N_9069,N_8774,N_8760);
nor U9070 (N_9070,N_8915,N_8767);
xor U9071 (N_9071,N_8851,N_8871);
nand U9072 (N_9072,N_8979,N_8794);
or U9073 (N_9073,N_8849,N_8942);
and U9074 (N_9074,N_8883,N_8797);
and U9075 (N_9075,N_8834,N_8754);
or U9076 (N_9076,N_8857,N_8949);
nor U9077 (N_9077,N_8777,N_8762);
nor U9078 (N_9078,N_8892,N_8990);
and U9079 (N_9079,N_8816,N_8973);
nor U9080 (N_9080,N_8827,N_8771);
nor U9081 (N_9081,N_8896,N_8975);
xnor U9082 (N_9082,N_8924,N_8960);
and U9083 (N_9083,N_8890,N_8922);
nand U9084 (N_9084,N_8759,N_8842);
xnor U9085 (N_9085,N_8954,N_8766);
and U9086 (N_9086,N_8830,N_8985);
nand U9087 (N_9087,N_8847,N_8824);
nand U9088 (N_9088,N_8876,N_8862);
nor U9089 (N_9089,N_8948,N_8832);
and U9090 (N_9090,N_8926,N_8936);
nor U9091 (N_9091,N_8763,N_8898);
nor U9092 (N_9092,N_8785,N_8750);
xor U9093 (N_9093,N_8968,N_8884);
and U9094 (N_9094,N_8980,N_8984);
xor U9095 (N_9095,N_8795,N_8904);
and U9096 (N_9096,N_8854,N_8901);
xor U9097 (N_9097,N_8934,N_8817);
nand U9098 (N_9098,N_8903,N_8868);
or U9099 (N_9099,N_8961,N_8965);
nand U9100 (N_9100,N_8768,N_8833);
nand U9101 (N_9101,N_8757,N_8938);
nand U9102 (N_9102,N_8870,N_8839);
nand U9103 (N_9103,N_8765,N_8803);
and U9104 (N_9104,N_8781,N_8986);
xor U9105 (N_9105,N_8818,N_8895);
nand U9106 (N_9106,N_8966,N_8835);
and U9107 (N_9107,N_8929,N_8983);
xor U9108 (N_9108,N_8786,N_8814);
or U9109 (N_9109,N_8977,N_8801);
xnor U9110 (N_9110,N_8988,N_8799);
or U9111 (N_9111,N_8788,N_8886);
nor U9112 (N_9112,N_8829,N_8933);
or U9113 (N_9113,N_8859,N_8875);
or U9114 (N_9114,N_8837,N_8941);
xnor U9115 (N_9115,N_8950,N_8902);
and U9116 (N_9116,N_8888,N_8887);
and U9117 (N_9117,N_8843,N_8813);
and U9118 (N_9118,N_8770,N_8804);
nand U9119 (N_9119,N_8881,N_8860);
nor U9120 (N_9120,N_8809,N_8959);
xor U9121 (N_9121,N_8889,N_8787);
nor U9122 (N_9122,N_8822,N_8908);
and U9123 (N_9123,N_8836,N_8976);
and U9124 (N_9124,N_8900,N_8969);
nand U9125 (N_9125,N_8967,N_8759);
or U9126 (N_9126,N_8996,N_8807);
nand U9127 (N_9127,N_8967,N_8885);
xnor U9128 (N_9128,N_8911,N_8921);
nor U9129 (N_9129,N_8996,N_8969);
nand U9130 (N_9130,N_8933,N_8999);
or U9131 (N_9131,N_8904,N_8978);
xor U9132 (N_9132,N_8972,N_8928);
and U9133 (N_9133,N_8755,N_8819);
xnor U9134 (N_9134,N_8830,N_8875);
nand U9135 (N_9135,N_8795,N_8889);
or U9136 (N_9136,N_8891,N_8815);
nor U9137 (N_9137,N_8773,N_8780);
and U9138 (N_9138,N_8914,N_8908);
nand U9139 (N_9139,N_8778,N_8904);
xor U9140 (N_9140,N_8858,N_8849);
and U9141 (N_9141,N_8929,N_8868);
xor U9142 (N_9142,N_8940,N_8904);
nor U9143 (N_9143,N_8797,N_8840);
and U9144 (N_9144,N_8993,N_8986);
nand U9145 (N_9145,N_8755,N_8818);
nor U9146 (N_9146,N_8967,N_8976);
nand U9147 (N_9147,N_8905,N_8871);
nor U9148 (N_9148,N_8918,N_8950);
xnor U9149 (N_9149,N_8778,N_8843);
and U9150 (N_9150,N_8959,N_8884);
nand U9151 (N_9151,N_8807,N_8850);
xnor U9152 (N_9152,N_8789,N_8882);
xor U9153 (N_9153,N_8866,N_8967);
or U9154 (N_9154,N_8758,N_8805);
nand U9155 (N_9155,N_8842,N_8970);
nor U9156 (N_9156,N_8932,N_8884);
xor U9157 (N_9157,N_8987,N_8823);
and U9158 (N_9158,N_8804,N_8928);
and U9159 (N_9159,N_8982,N_8767);
and U9160 (N_9160,N_8983,N_8959);
xor U9161 (N_9161,N_8969,N_8823);
and U9162 (N_9162,N_8790,N_8925);
and U9163 (N_9163,N_8930,N_8784);
nand U9164 (N_9164,N_8757,N_8811);
or U9165 (N_9165,N_8872,N_8904);
or U9166 (N_9166,N_8765,N_8763);
nand U9167 (N_9167,N_8772,N_8781);
nand U9168 (N_9168,N_8866,N_8832);
nand U9169 (N_9169,N_8966,N_8922);
or U9170 (N_9170,N_8785,N_8861);
or U9171 (N_9171,N_8795,N_8916);
nand U9172 (N_9172,N_8945,N_8815);
nor U9173 (N_9173,N_8982,N_8777);
and U9174 (N_9174,N_8866,N_8854);
nor U9175 (N_9175,N_8884,N_8881);
and U9176 (N_9176,N_8835,N_8848);
xor U9177 (N_9177,N_8757,N_8845);
nand U9178 (N_9178,N_8986,N_8770);
nand U9179 (N_9179,N_8888,N_8823);
or U9180 (N_9180,N_8811,N_8906);
and U9181 (N_9181,N_8946,N_8895);
and U9182 (N_9182,N_8956,N_8905);
xor U9183 (N_9183,N_8865,N_8836);
and U9184 (N_9184,N_8950,N_8872);
nor U9185 (N_9185,N_8983,N_8787);
nor U9186 (N_9186,N_8781,N_8975);
and U9187 (N_9187,N_8992,N_8836);
xor U9188 (N_9188,N_8878,N_8784);
xnor U9189 (N_9189,N_8811,N_8908);
and U9190 (N_9190,N_8751,N_8906);
nand U9191 (N_9191,N_8917,N_8786);
and U9192 (N_9192,N_8939,N_8830);
or U9193 (N_9193,N_8925,N_8907);
nand U9194 (N_9194,N_8944,N_8916);
or U9195 (N_9195,N_8844,N_8941);
xor U9196 (N_9196,N_8856,N_8805);
nand U9197 (N_9197,N_8863,N_8776);
or U9198 (N_9198,N_8869,N_8760);
nand U9199 (N_9199,N_8822,N_8836);
xor U9200 (N_9200,N_8772,N_8800);
and U9201 (N_9201,N_8904,N_8790);
or U9202 (N_9202,N_8891,N_8818);
nand U9203 (N_9203,N_8811,N_8964);
nand U9204 (N_9204,N_8904,N_8847);
or U9205 (N_9205,N_8831,N_8868);
and U9206 (N_9206,N_8954,N_8860);
xor U9207 (N_9207,N_8984,N_8853);
or U9208 (N_9208,N_8996,N_8918);
nand U9209 (N_9209,N_8812,N_8793);
and U9210 (N_9210,N_8883,N_8972);
nand U9211 (N_9211,N_8817,N_8804);
nor U9212 (N_9212,N_8989,N_8959);
nand U9213 (N_9213,N_8759,N_8855);
nor U9214 (N_9214,N_8853,N_8800);
nand U9215 (N_9215,N_8833,N_8858);
and U9216 (N_9216,N_8824,N_8798);
and U9217 (N_9217,N_8828,N_8810);
nand U9218 (N_9218,N_8984,N_8898);
nor U9219 (N_9219,N_8753,N_8985);
nor U9220 (N_9220,N_8914,N_8753);
xor U9221 (N_9221,N_8782,N_8856);
nand U9222 (N_9222,N_8950,N_8908);
nor U9223 (N_9223,N_8833,N_8980);
nand U9224 (N_9224,N_8867,N_8849);
nor U9225 (N_9225,N_8804,N_8920);
nand U9226 (N_9226,N_8805,N_8975);
or U9227 (N_9227,N_8850,N_8846);
nand U9228 (N_9228,N_8863,N_8961);
nor U9229 (N_9229,N_8806,N_8990);
xnor U9230 (N_9230,N_8781,N_8928);
or U9231 (N_9231,N_8956,N_8774);
and U9232 (N_9232,N_8770,N_8996);
or U9233 (N_9233,N_8832,N_8921);
nor U9234 (N_9234,N_8835,N_8977);
xor U9235 (N_9235,N_8780,N_8782);
or U9236 (N_9236,N_8891,N_8856);
nor U9237 (N_9237,N_8947,N_8836);
or U9238 (N_9238,N_8954,N_8936);
or U9239 (N_9239,N_8859,N_8783);
and U9240 (N_9240,N_8937,N_8919);
and U9241 (N_9241,N_8961,N_8920);
xnor U9242 (N_9242,N_8775,N_8836);
and U9243 (N_9243,N_8943,N_8826);
nand U9244 (N_9244,N_8874,N_8956);
xnor U9245 (N_9245,N_8777,N_8792);
nand U9246 (N_9246,N_8940,N_8817);
and U9247 (N_9247,N_8991,N_8886);
or U9248 (N_9248,N_8999,N_8910);
and U9249 (N_9249,N_8778,N_8761);
nor U9250 (N_9250,N_9136,N_9245);
nor U9251 (N_9251,N_9209,N_9173);
and U9252 (N_9252,N_9117,N_9214);
or U9253 (N_9253,N_9015,N_9029);
nand U9254 (N_9254,N_9002,N_9140);
nand U9255 (N_9255,N_9189,N_9167);
nand U9256 (N_9256,N_9203,N_9206);
xor U9257 (N_9257,N_9187,N_9014);
and U9258 (N_9258,N_9126,N_9229);
nand U9259 (N_9259,N_9218,N_9048);
xnor U9260 (N_9260,N_9095,N_9121);
or U9261 (N_9261,N_9194,N_9240);
nor U9262 (N_9262,N_9088,N_9078);
xnor U9263 (N_9263,N_9163,N_9197);
and U9264 (N_9264,N_9112,N_9177);
nor U9265 (N_9265,N_9059,N_9246);
or U9266 (N_9266,N_9020,N_9032);
xnor U9267 (N_9267,N_9198,N_9151);
nand U9268 (N_9268,N_9181,N_9075);
and U9269 (N_9269,N_9208,N_9129);
xor U9270 (N_9270,N_9232,N_9047);
and U9271 (N_9271,N_9133,N_9216);
xor U9272 (N_9272,N_9186,N_9195);
or U9273 (N_9273,N_9179,N_9217);
and U9274 (N_9274,N_9104,N_9144);
xnor U9275 (N_9275,N_9161,N_9239);
xor U9276 (N_9276,N_9238,N_9164);
nor U9277 (N_9277,N_9087,N_9099);
nor U9278 (N_9278,N_9006,N_9065);
nor U9279 (N_9279,N_9130,N_9124);
or U9280 (N_9280,N_9084,N_9150);
and U9281 (N_9281,N_9023,N_9007);
nand U9282 (N_9282,N_9019,N_9086);
or U9283 (N_9283,N_9131,N_9158);
nand U9284 (N_9284,N_9021,N_9040);
or U9285 (N_9285,N_9068,N_9009);
nand U9286 (N_9286,N_9123,N_9118);
nor U9287 (N_9287,N_9051,N_9185);
nand U9288 (N_9288,N_9119,N_9026);
nand U9289 (N_9289,N_9005,N_9225);
xnor U9290 (N_9290,N_9132,N_9241);
nor U9291 (N_9291,N_9157,N_9204);
xnor U9292 (N_9292,N_9137,N_9063);
nor U9293 (N_9293,N_9011,N_9235);
or U9294 (N_9294,N_9028,N_9142);
xor U9295 (N_9295,N_9069,N_9052);
nor U9296 (N_9296,N_9000,N_9033);
or U9297 (N_9297,N_9156,N_9091);
nand U9298 (N_9298,N_9237,N_9146);
nor U9299 (N_9299,N_9192,N_9012);
xnor U9300 (N_9300,N_9101,N_9223);
xor U9301 (N_9301,N_9178,N_9108);
nand U9302 (N_9302,N_9058,N_9188);
xor U9303 (N_9303,N_9045,N_9122);
nor U9304 (N_9304,N_9202,N_9175);
xor U9305 (N_9305,N_9227,N_9074);
or U9306 (N_9306,N_9176,N_9024);
nor U9307 (N_9307,N_9172,N_9145);
nand U9308 (N_9308,N_9042,N_9125);
nand U9309 (N_9309,N_9138,N_9134);
or U9310 (N_9310,N_9022,N_9107);
or U9311 (N_9311,N_9010,N_9160);
nand U9312 (N_9312,N_9062,N_9030);
nor U9313 (N_9313,N_9228,N_9139);
nor U9314 (N_9314,N_9085,N_9098);
and U9315 (N_9315,N_9248,N_9061);
nand U9316 (N_9316,N_9220,N_9105);
and U9317 (N_9317,N_9190,N_9018);
and U9318 (N_9318,N_9182,N_9111);
and U9319 (N_9319,N_9004,N_9102);
xnor U9320 (N_9320,N_9056,N_9219);
and U9321 (N_9321,N_9044,N_9097);
xnor U9322 (N_9322,N_9128,N_9116);
nor U9323 (N_9323,N_9115,N_9222);
and U9324 (N_9324,N_9171,N_9073);
and U9325 (N_9325,N_9155,N_9221);
or U9326 (N_9326,N_9143,N_9162);
or U9327 (N_9327,N_9038,N_9013);
nand U9328 (N_9328,N_9039,N_9081);
nand U9329 (N_9329,N_9233,N_9174);
nor U9330 (N_9330,N_9183,N_9050);
nand U9331 (N_9331,N_9025,N_9120);
nor U9332 (N_9332,N_9031,N_9090);
xor U9333 (N_9333,N_9113,N_9096);
xor U9334 (N_9334,N_9082,N_9114);
or U9335 (N_9335,N_9207,N_9234);
nor U9336 (N_9336,N_9154,N_9149);
nor U9337 (N_9337,N_9064,N_9147);
and U9338 (N_9338,N_9094,N_9166);
nand U9339 (N_9339,N_9016,N_9055);
nand U9340 (N_9340,N_9215,N_9001);
or U9341 (N_9341,N_9027,N_9169);
or U9342 (N_9342,N_9212,N_9083);
or U9343 (N_9343,N_9247,N_9076);
xor U9344 (N_9344,N_9127,N_9205);
and U9345 (N_9345,N_9067,N_9041);
or U9346 (N_9346,N_9148,N_9153);
and U9347 (N_9347,N_9200,N_9017);
nor U9348 (N_9348,N_9230,N_9191);
nor U9349 (N_9349,N_9077,N_9231);
or U9350 (N_9350,N_9035,N_9184);
or U9351 (N_9351,N_9236,N_9249);
nor U9352 (N_9352,N_9224,N_9057);
nor U9353 (N_9353,N_9210,N_9199);
nor U9354 (N_9354,N_9211,N_9110);
or U9355 (N_9355,N_9165,N_9243);
nand U9356 (N_9356,N_9066,N_9070);
nand U9357 (N_9357,N_9049,N_9226);
nor U9358 (N_9358,N_9180,N_9092);
or U9359 (N_9359,N_9079,N_9043);
nor U9360 (N_9360,N_9036,N_9093);
nor U9361 (N_9361,N_9072,N_9213);
nor U9362 (N_9362,N_9244,N_9168);
nand U9363 (N_9363,N_9109,N_9152);
nand U9364 (N_9364,N_9100,N_9037);
nor U9365 (N_9365,N_9089,N_9060);
or U9366 (N_9366,N_9053,N_9071);
nand U9367 (N_9367,N_9008,N_9054);
nor U9368 (N_9368,N_9196,N_9135);
nand U9369 (N_9369,N_9080,N_9159);
xnor U9370 (N_9370,N_9193,N_9242);
nor U9371 (N_9371,N_9034,N_9103);
and U9372 (N_9372,N_9046,N_9141);
nor U9373 (N_9373,N_9170,N_9106);
xnor U9374 (N_9374,N_9201,N_9003);
nor U9375 (N_9375,N_9084,N_9028);
nor U9376 (N_9376,N_9115,N_9192);
xor U9377 (N_9377,N_9006,N_9058);
and U9378 (N_9378,N_9170,N_9005);
and U9379 (N_9379,N_9131,N_9138);
or U9380 (N_9380,N_9156,N_9215);
nand U9381 (N_9381,N_9162,N_9172);
or U9382 (N_9382,N_9229,N_9067);
nand U9383 (N_9383,N_9176,N_9090);
nand U9384 (N_9384,N_9006,N_9063);
or U9385 (N_9385,N_9109,N_9170);
nor U9386 (N_9386,N_9129,N_9100);
xor U9387 (N_9387,N_9143,N_9133);
nor U9388 (N_9388,N_9017,N_9132);
nor U9389 (N_9389,N_9188,N_9222);
nand U9390 (N_9390,N_9126,N_9081);
xnor U9391 (N_9391,N_9084,N_9202);
or U9392 (N_9392,N_9119,N_9168);
nor U9393 (N_9393,N_9234,N_9094);
nor U9394 (N_9394,N_9081,N_9017);
nand U9395 (N_9395,N_9205,N_9130);
nand U9396 (N_9396,N_9135,N_9074);
xor U9397 (N_9397,N_9040,N_9102);
or U9398 (N_9398,N_9087,N_9150);
and U9399 (N_9399,N_9193,N_9210);
or U9400 (N_9400,N_9108,N_9185);
and U9401 (N_9401,N_9166,N_9051);
or U9402 (N_9402,N_9180,N_9001);
or U9403 (N_9403,N_9077,N_9190);
nor U9404 (N_9404,N_9149,N_9244);
nand U9405 (N_9405,N_9160,N_9182);
and U9406 (N_9406,N_9224,N_9102);
nand U9407 (N_9407,N_9092,N_9124);
and U9408 (N_9408,N_9121,N_9070);
and U9409 (N_9409,N_9113,N_9074);
nor U9410 (N_9410,N_9072,N_9245);
xor U9411 (N_9411,N_9123,N_9210);
and U9412 (N_9412,N_9223,N_9025);
or U9413 (N_9413,N_9099,N_9145);
nand U9414 (N_9414,N_9082,N_9008);
or U9415 (N_9415,N_9155,N_9004);
nand U9416 (N_9416,N_9116,N_9195);
nand U9417 (N_9417,N_9172,N_9022);
and U9418 (N_9418,N_9161,N_9015);
nand U9419 (N_9419,N_9144,N_9075);
nand U9420 (N_9420,N_9215,N_9068);
and U9421 (N_9421,N_9090,N_9215);
xnor U9422 (N_9422,N_9172,N_9006);
nand U9423 (N_9423,N_9119,N_9060);
xor U9424 (N_9424,N_9242,N_9224);
nor U9425 (N_9425,N_9218,N_9159);
or U9426 (N_9426,N_9010,N_9063);
nor U9427 (N_9427,N_9007,N_9201);
nand U9428 (N_9428,N_9095,N_9223);
nor U9429 (N_9429,N_9127,N_9149);
nor U9430 (N_9430,N_9141,N_9227);
nor U9431 (N_9431,N_9235,N_9100);
and U9432 (N_9432,N_9069,N_9086);
nand U9433 (N_9433,N_9187,N_9027);
nor U9434 (N_9434,N_9147,N_9080);
xor U9435 (N_9435,N_9061,N_9063);
xor U9436 (N_9436,N_9177,N_9196);
nand U9437 (N_9437,N_9018,N_9231);
nand U9438 (N_9438,N_9079,N_9083);
xnor U9439 (N_9439,N_9237,N_9097);
xnor U9440 (N_9440,N_9127,N_9160);
xnor U9441 (N_9441,N_9222,N_9175);
or U9442 (N_9442,N_9078,N_9113);
nand U9443 (N_9443,N_9022,N_9170);
xnor U9444 (N_9444,N_9113,N_9205);
or U9445 (N_9445,N_9192,N_9028);
nor U9446 (N_9446,N_9230,N_9032);
xor U9447 (N_9447,N_9107,N_9051);
xor U9448 (N_9448,N_9178,N_9124);
xor U9449 (N_9449,N_9184,N_9100);
nand U9450 (N_9450,N_9075,N_9196);
and U9451 (N_9451,N_9166,N_9148);
and U9452 (N_9452,N_9039,N_9164);
nor U9453 (N_9453,N_9103,N_9173);
nor U9454 (N_9454,N_9091,N_9102);
or U9455 (N_9455,N_9135,N_9018);
nor U9456 (N_9456,N_9020,N_9209);
nand U9457 (N_9457,N_9036,N_9070);
xor U9458 (N_9458,N_9018,N_9211);
and U9459 (N_9459,N_9149,N_9236);
xnor U9460 (N_9460,N_9116,N_9223);
nor U9461 (N_9461,N_9005,N_9032);
and U9462 (N_9462,N_9222,N_9235);
nand U9463 (N_9463,N_9238,N_9222);
or U9464 (N_9464,N_9133,N_9240);
and U9465 (N_9465,N_9041,N_9075);
nor U9466 (N_9466,N_9122,N_9100);
or U9467 (N_9467,N_9168,N_9038);
and U9468 (N_9468,N_9237,N_9081);
or U9469 (N_9469,N_9014,N_9176);
or U9470 (N_9470,N_9104,N_9109);
or U9471 (N_9471,N_9085,N_9206);
nand U9472 (N_9472,N_9193,N_9054);
nor U9473 (N_9473,N_9176,N_9077);
nor U9474 (N_9474,N_9065,N_9183);
nor U9475 (N_9475,N_9141,N_9122);
or U9476 (N_9476,N_9087,N_9024);
xnor U9477 (N_9477,N_9174,N_9114);
or U9478 (N_9478,N_9185,N_9193);
nor U9479 (N_9479,N_9005,N_9041);
and U9480 (N_9480,N_9101,N_9149);
and U9481 (N_9481,N_9205,N_9143);
nor U9482 (N_9482,N_9041,N_9095);
nand U9483 (N_9483,N_9232,N_9000);
nor U9484 (N_9484,N_9182,N_9149);
nand U9485 (N_9485,N_9150,N_9174);
and U9486 (N_9486,N_9055,N_9108);
or U9487 (N_9487,N_9092,N_9211);
nand U9488 (N_9488,N_9171,N_9174);
and U9489 (N_9489,N_9011,N_9134);
nand U9490 (N_9490,N_9242,N_9192);
or U9491 (N_9491,N_9062,N_9198);
xor U9492 (N_9492,N_9173,N_9002);
nand U9493 (N_9493,N_9188,N_9164);
xnor U9494 (N_9494,N_9000,N_9248);
or U9495 (N_9495,N_9053,N_9108);
and U9496 (N_9496,N_9051,N_9119);
xor U9497 (N_9497,N_9240,N_9203);
xnor U9498 (N_9498,N_9107,N_9067);
or U9499 (N_9499,N_9047,N_9243);
xor U9500 (N_9500,N_9262,N_9363);
and U9501 (N_9501,N_9352,N_9407);
or U9502 (N_9502,N_9449,N_9459);
and U9503 (N_9503,N_9487,N_9364);
nand U9504 (N_9504,N_9312,N_9499);
nor U9505 (N_9505,N_9446,N_9304);
or U9506 (N_9506,N_9464,N_9329);
or U9507 (N_9507,N_9265,N_9466);
or U9508 (N_9508,N_9256,N_9368);
and U9509 (N_9509,N_9340,N_9257);
nor U9510 (N_9510,N_9461,N_9467);
or U9511 (N_9511,N_9331,N_9382);
and U9512 (N_9512,N_9403,N_9444);
nand U9513 (N_9513,N_9404,N_9405);
or U9514 (N_9514,N_9384,N_9313);
xnor U9515 (N_9515,N_9337,N_9290);
nand U9516 (N_9516,N_9317,N_9438);
nor U9517 (N_9517,N_9483,N_9310);
or U9518 (N_9518,N_9372,N_9434);
nand U9519 (N_9519,N_9359,N_9396);
nor U9520 (N_9520,N_9472,N_9264);
xor U9521 (N_9521,N_9356,N_9482);
and U9522 (N_9522,N_9383,N_9360);
and U9523 (N_9523,N_9453,N_9498);
nor U9524 (N_9524,N_9377,N_9366);
and U9525 (N_9525,N_9333,N_9254);
xnor U9526 (N_9526,N_9454,N_9282);
xor U9527 (N_9527,N_9490,N_9489);
nand U9528 (N_9528,N_9495,N_9432);
nand U9529 (N_9529,N_9277,N_9378);
and U9530 (N_9530,N_9379,N_9494);
nand U9531 (N_9531,N_9381,N_9347);
nor U9532 (N_9532,N_9465,N_9392);
nand U9533 (N_9533,N_9485,N_9278);
and U9534 (N_9534,N_9270,N_9341);
and U9535 (N_9535,N_9354,N_9321);
or U9536 (N_9536,N_9477,N_9408);
xor U9537 (N_9537,N_9420,N_9339);
nor U9538 (N_9538,N_9258,N_9425);
nand U9539 (N_9539,N_9322,N_9394);
and U9540 (N_9540,N_9428,N_9348);
or U9541 (N_9541,N_9338,N_9463);
xnor U9542 (N_9542,N_9447,N_9388);
nor U9543 (N_9543,N_9301,N_9323);
and U9544 (N_9544,N_9296,N_9299);
nor U9545 (N_9545,N_9390,N_9402);
and U9546 (N_9546,N_9426,N_9441);
nand U9547 (N_9547,N_9288,N_9385);
or U9548 (N_9548,N_9488,N_9315);
or U9549 (N_9549,N_9484,N_9266);
and U9550 (N_9550,N_9255,N_9389);
and U9551 (N_9551,N_9344,N_9260);
nor U9552 (N_9552,N_9279,N_9320);
or U9553 (N_9553,N_9429,N_9410);
and U9554 (N_9554,N_9330,N_9401);
or U9555 (N_9555,N_9411,N_9274);
xnor U9556 (N_9556,N_9427,N_9305);
xnor U9557 (N_9557,N_9457,N_9286);
or U9558 (N_9558,N_9253,N_9335);
nor U9559 (N_9559,N_9480,N_9287);
nand U9560 (N_9560,N_9285,N_9291);
or U9561 (N_9561,N_9311,N_9462);
xnor U9562 (N_9562,N_9294,N_9450);
xor U9563 (N_9563,N_9439,N_9324);
nor U9564 (N_9564,N_9442,N_9493);
xor U9565 (N_9565,N_9433,N_9268);
or U9566 (N_9566,N_9496,N_9292);
or U9567 (N_9567,N_9267,N_9458);
xnor U9568 (N_9568,N_9460,N_9275);
nor U9569 (N_9569,N_9351,N_9471);
nor U9570 (N_9570,N_9309,N_9334);
xnor U9571 (N_9571,N_9400,N_9343);
or U9572 (N_9572,N_9328,N_9424);
nand U9573 (N_9573,N_9355,N_9478);
xnor U9574 (N_9574,N_9371,N_9362);
or U9575 (N_9575,N_9409,N_9468);
xor U9576 (N_9576,N_9297,N_9492);
nand U9577 (N_9577,N_9399,N_9370);
nor U9578 (N_9578,N_9276,N_9491);
nor U9579 (N_9579,N_9263,N_9397);
nor U9580 (N_9580,N_9289,N_9452);
and U9581 (N_9581,N_9436,N_9252);
and U9582 (N_9582,N_9481,N_9308);
and U9583 (N_9583,N_9393,N_9314);
xor U9584 (N_9584,N_9353,N_9415);
nand U9585 (N_9585,N_9373,N_9295);
xnor U9586 (N_9586,N_9261,N_9349);
and U9587 (N_9587,N_9479,N_9435);
xnor U9588 (N_9588,N_9251,N_9280);
nand U9589 (N_9589,N_9451,N_9273);
nor U9590 (N_9590,N_9306,N_9325);
nor U9591 (N_9591,N_9469,N_9327);
or U9592 (N_9592,N_9298,N_9423);
xnor U9593 (N_9593,N_9430,N_9475);
nand U9594 (N_9594,N_9300,N_9342);
and U9595 (N_9595,N_9412,N_9473);
and U9596 (N_9596,N_9332,N_9307);
xor U9597 (N_9597,N_9419,N_9345);
xor U9598 (N_9598,N_9418,N_9367);
and U9599 (N_9599,N_9281,N_9272);
and U9600 (N_9600,N_9414,N_9455);
xnor U9601 (N_9601,N_9476,N_9250);
or U9602 (N_9602,N_9376,N_9445);
xor U9603 (N_9603,N_9387,N_9486);
nand U9604 (N_9604,N_9319,N_9375);
nor U9605 (N_9605,N_9284,N_9316);
or U9606 (N_9606,N_9303,N_9259);
or U9607 (N_9607,N_9440,N_9361);
nor U9608 (N_9608,N_9497,N_9456);
nor U9609 (N_9609,N_9269,N_9391);
nor U9610 (N_9610,N_9271,N_9380);
xnor U9611 (N_9611,N_9302,N_9413);
and U9612 (N_9612,N_9416,N_9474);
xnor U9613 (N_9613,N_9350,N_9437);
xnor U9614 (N_9614,N_9357,N_9336);
xor U9615 (N_9615,N_9421,N_9358);
nand U9616 (N_9616,N_9422,N_9374);
nor U9617 (N_9617,N_9395,N_9443);
nand U9618 (N_9618,N_9318,N_9470);
nor U9619 (N_9619,N_9431,N_9326);
xnor U9620 (N_9620,N_9406,N_9369);
or U9621 (N_9621,N_9398,N_9346);
and U9622 (N_9622,N_9365,N_9417);
nor U9623 (N_9623,N_9293,N_9448);
nand U9624 (N_9624,N_9386,N_9283);
xnor U9625 (N_9625,N_9334,N_9431);
nand U9626 (N_9626,N_9261,N_9393);
or U9627 (N_9627,N_9301,N_9413);
nor U9628 (N_9628,N_9409,N_9334);
or U9629 (N_9629,N_9419,N_9370);
and U9630 (N_9630,N_9499,N_9311);
or U9631 (N_9631,N_9442,N_9399);
or U9632 (N_9632,N_9282,N_9275);
xnor U9633 (N_9633,N_9437,N_9285);
nor U9634 (N_9634,N_9267,N_9378);
or U9635 (N_9635,N_9295,N_9275);
nor U9636 (N_9636,N_9442,N_9286);
and U9637 (N_9637,N_9470,N_9463);
nor U9638 (N_9638,N_9488,N_9448);
and U9639 (N_9639,N_9262,N_9387);
nor U9640 (N_9640,N_9450,N_9444);
or U9641 (N_9641,N_9419,N_9352);
or U9642 (N_9642,N_9362,N_9286);
or U9643 (N_9643,N_9349,N_9267);
and U9644 (N_9644,N_9347,N_9259);
xnor U9645 (N_9645,N_9293,N_9429);
xor U9646 (N_9646,N_9282,N_9498);
or U9647 (N_9647,N_9387,N_9451);
and U9648 (N_9648,N_9311,N_9260);
nor U9649 (N_9649,N_9475,N_9324);
nor U9650 (N_9650,N_9461,N_9277);
nor U9651 (N_9651,N_9254,N_9343);
nand U9652 (N_9652,N_9383,N_9259);
nand U9653 (N_9653,N_9473,N_9447);
xor U9654 (N_9654,N_9373,N_9377);
or U9655 (N_9655,N_9401,N_9374);
nand U9656 (N_9656,N_9310,N_9407);
xnor U9657 (N_9657,N_9276,N_9292);
and U9658 (N_9658,N_9304,N_9367);
nor U9659 (N_9659,N_9256,N_9378);
or U9660 (N_9660,N_9435,N_9334);
xnor U9661 (N_9661,N_9457,N_9394);
nand U9662 (N_9662,N_9340,N_9322);
nor U9663 (N_9663,N_9337,N_9499);
nand U9664 (N_9664,N_9344,N_9419);
nand U9665 (N_9665,N_9282,N_9488);
nor U9666 (N_9666,N_9406,N_9265);
xnor U9667 (N_9667,N_9416,N_9339);
nand U9668 (N_9668,N_9420,N_9475);
nand U9669 (N_9669,N_9436,N_9359);
or U9670 (N_9670,N_9386,N_9401);
nor U9671 (N_9671,N_9452,N_9262);
xnor U9672 (N_9672,N_9307,N_9465);
and U9673 (N_9673,N_9499,N_9275);
and U9674 (N_9674,N_9336,N_9405);
and U9675 (N_9675,N_9424,N_9472);
nor U9676 (N_9676,N_9483,N_9427);
xnor U9677 (N_9677,N_9480,N_9278);
nor U9678 (N_9678,N_9415,N_9362);
xor U9679 (N_9679,N_9497,N_9381);
or U9680 (N_9680,N_9395,N_9402);
and U9681 (N_9681,N_9277,N_9293);
xnor U9682 (N_9682,N_9313,N_9275);
and U9683 (N_9683,N_9472,N_9274);
and U9684 (N_9684,N_9303,N_9291);
nand U9685 (N_9685,N_9319,N_9256);
nand U9686 (N_9686,N_9484,N_9292);
or U9687 (N_9687,N_9427,N_9375);
xnor U9688 (N_9688,N_9441,N_9437);
xnor U9689 (N_9689,N_9408,N_9499);
nor U9690 (N_9690,N_9441,N_9477);
and U9691 (N_9691,N_9364,N_9454);
or U9692 (N_9692,N_9292,N_9449);
nor U9693 (N_9693,N_9292,N_9423);
nor U9694 (N_9694,N_9454,N_9325);
or U9695 (N_9695,N_9388,N_9265);
nor U9696 (N_9696,N_9291,N_9373);
or U9697 (N_9697,N_9444,N_9460);
nand U9698 (N_9698,N_9316,N_9354);
nor U9699 (N_9699,N_9356,N_9403);
and U9700 (N_9700,N_9371,N_9285);
or U9701 (N_9701,N_9317,N_9377);
or U9702 (N_9702,N_9390,N_9479);
and U9703 (N_9703,N_9417,N_9474);
and U9704 (N_9704,N_9359,N_9320);
nand U9705 (N_9705,N_9289,N_9430);
xnor U9706 (N_9706,N_9409,N_9288);
nand U9707 (N_9707,N_9386,N_9426);
nor U9708 (N_9708,N_9287,N_9271);
and U9709 (N_9709,N_9262,N_9492);
nand U9710 (N_9710,N_9488,N_9351);
xor U9711 (N_9711,N_9495,N_9342);
and U9712 (N_9712,N_9252,N_9392);
nor U9713 (N_9713,N_9325,N_9260);
and U9714 (N_9714,N_9271,N_9360);
nor U9715 (N_9715,N_9307,N_9394);
nand U9716 (N_9716,N_9496,N_9493);
nor U9717 (N_9717,N_9378,N_9465);
and U9718 (N_9718,N_9388,N_9449);
nor U9719 (N_9719,N_9475,N_9374);
nor U9720 (N_9720,N_9395,N_9424);
nor U9721 (N_9721,N_9430,N_9448);
xnor U9722 (N_9722,N_9449,N_9445);
nand U9723 (N_9723,N_9371,N_9280);
xor U9724 (N_9724,N_9388,N_9471);
and U9725 (N_9725,N_9421,N_9430);
nand U9726 (N_9726,N_9282,N_9405);
nand U9727 (N_9727,N_9318,N_9364);
and U9728 (N_9728,N_9421,N_9425);
nor U9729 (N_9729,N_9313,N_9429);
xor U9730 (N_9730,N_9391,N_9255);
and U9731 (N_9731,N_9371,N_9335);
or U9732 (N_9732,N_9333,N_9497);
nand U9733 (N_9733,N_9481,N_9318);
and U9734 (N_9734,N_9485,N_9459);
or U9735 (N_9735,N_9375,N_9370);
xnor U9736 (N_9736,N_9364,N_9493);
nand U9737 (N_9737,N_9436,N_9352);
or U9738 (N_9738,N_9296,N_9308);
nand U9739 (N_9739,N_9418,N_9333);
and U9740 (N_9740,N_9297,N_9262);
nor U9741 (N_9741,N_9346,N_9426);
nand U9742 (N_9742,N_9496,N_9355);
and U9743 (N_9743,N_9428,N_9334);
nor U9744 (N_9744,N_9434,N_9307);
xnor U9745 (N_9745,N_9313,N_9377);
or U9746 (N_9746,N_9284,N_9398);
xor U9747 (N_9747,N_9387,N_9353);
nand U9748 (N_9748,N_9485,N_9303);
nand U9749 (N_9749,N_9462,N_9333);
and U9750 (N_9750,N_9724,N_9529);
nand U9751 (N_9751,N_9503,N_9715);
nor U9752 (N_9752,N_9543,N_9571);
nor U9753 (N_9753,N_9727,N_9520);
nand U9754 (N_9754,N_9680,N_9653);
nor U9755 (N_9755,N_9592,N_9588);
and U9756 (N_9756,N_9746,N_9615);
or U9757 (N_9757,N_9515,N_9623);
or U9758 (N_9758,N_9514,N_9531);
nor U9759 (N_9759,N_9532,N_9572);
xnor U9760 (N_9760,N_9641,N_9707);
or U9761 (N_9761,N_9675,N_9664);
and U9762 (N_9762,N_9647,N_9679);
and U9763 (N_9763,N_9749,N_9690);
nor U9764 (N_9764,N_9577,N_9534);
nor U9765 (N_9765,N_9671,N_9578);
nand U9766 (N_9766,N_9564,N_9669);
nand U9767 (N_9767,N_9622,N_9716);
and U9768 (N_9768,N_9734,N_9616);
nand U9769 (N_9769,N_9652,N_9639);
nand U9770 (N_9770,N_9747,N_9689);
and U9771 (N_9771,N_9637,N_9657);
and U9772 (N_9772,N_9740,N_9567);
xnor U9773 (N_9773,N_9708,N_9599);
nand U9774 (N_9774,N_9633,N_9674);
nand U9775 (N_9775,N_9553,N_9714);
xor U9776 (N_9776,N_9551,N_9505);
and U9777 (N_9777,N_9518,N_9525);
and U9778 (N_9778,N_9739,N_9663);
and U9779 (N_9779,N_9506,N_9646);
xnor U9780 (N_9780,N_9598,N_9594);
nor U9781 (N_9781,N_9721,N_9603);
or U9782 (N_9782,N_9713,N_9596);
xor U9783 (N_9783,N_9700,N_9711);
and U9784 (N_9784,N_9651,N_9738);
nor U9785 (N_9785,N_9628,N_9557);
nand U9786 (N_9786,N_9648,N_9545);
or U9787 (N_9787,N_9654,N_9565);
nand U9788 (N_9788,N_9683,N_9576);
xor U9789 (N_9789,N_9579,N_9722);
nand U9790 (N_9790,N_9611,N_9587);
nand U9791 (N_9791,N_9613,N_9546);
or U9792 (N_9792,N_9712,N_9600);
xor U9793 (N_9793,N_9575,N_9692);
or U9794 (N_9794,N_9530,N_9619);
nor U9795 (N_9795,N_9582,N_9629);
nand U9796 (N_9796,N_9562,N_9649);
nor U9797 (N_9797,N_9583,N_9549);
or U9798 (N_9798,N_9695,N_9535);
nor U9799 (N_9799,N_9741,N_9642);
or U9800 (N_9800,N_9504,N_9558);
xor U9801 (N_9801,N_9609,N_9574);
or U9802 (N_9802,N_9511,N_9697);
and U9803 (N_9803,N_9590,N_9559);
nand U9804 (N_9804,N_9507,N_9569);
nand U9805 (N_9805,N_9573,N_9635);
xor U9806 (N_9806,N_9659,N_9709);
xnor U9807 (N_9807,N_9729,N_9644);
and U9808 (N_9808,N_9720,N_9580);
and U9809 (N_9809,N_9526,N_9607);
xor U9810 (N_9810,N_9550,N_9684);
and U9811 (N_9811,N_9634,N_9560);
nor U9812 (N_9812,N_9718,N_9547);
nor U9813 (N_9813,N_9627,N_9593);
nor U9814 (N_9814,N_9521,N_9737);
and U9815 (N_9815,N_9661,N_9608);
and U9816 (N_9816,N_9640,N_9702);
nor U9817 (N_9817,N_9730,N_9527);
and U9818 (N_9818,N_9673,N_9732);
or U9819 (N_9819,N_9660,N_9698);
or U9820 (N_9820,N_9510,N_9541);
or U9821 (N_9821,N_9602,N_9589);
nand U9822 (N_9822,N_9668,N_9536);
and U9823 (N_9823,N_9509,N_9605);
or U9824 (N_9824,N_9524,N_9672);
and U9825 (N_9825,N_9706,N_9745);
nor U9826 (N_9826,N_9743,N_9665);
xor U9827 (N_9827,N_9705,N_9617);
nand U9828 (N_9828,N_9687,N_9555);
nor U9829 (N_9829,N_9638,N_9537);
or U9830 (N_9830,N_9523,N_9658);
nor U9831 (N_9831,N_9696,N_9500);
and U9832 (N_9832,N_9614,N_9744);
and U9833 (N_9833,N_9563,N_9552);
and U9834 (N_9834,N_9533,N_9542);
xor U9835 (N_9835,N_9725,N_9694);
xnor U9836 (N_9836,N_9544,N_9726);
nand U9837 (N_9837,N_9517,N_9540);
xnor U9838 (N_9838,N_9606,N_9512);
and U9839 (N_9839,N_9670,N_9701);
nor U9840 (N_9840,N_9561,N_9568);
xor U9841 (N_9841,N_9585,N_9597);
nand U9842 (N_9842,N_9630,N_9501);
and U9843 (N_9843,N_9636,N_9667);
nor U9844 (N_9844,N_9612,N_9581);
and U9845 (N_9845,N_9554,N_9621);
nand U9846 (N_9846,N_9570,N_9650);
xnor U9847 (N_9847,N_9685,N_9688);
nor U9848 (N_9848,N_9691,N_9735);
nor U9849 (N_9849,N_9566,N_9699);
and U9850 (N_9850,N_9513,N_9645);
nand U9851 (N_9851,N_9516,N_9704);
and U9852 (N_9852,N_9742,N_9643);
xnor U9853 (N_9853,N_9682,N_9519);
and U9854 (N_9854,N_9662,N_9719);
and U9855 (N_9855,N_9631,N_9548);
nand U9856 (N_9856,N_9731,N_9522);
and U9857 (N_9857,N_9655,N_9666);
and U9858 (N_9858,N_9710,N_9624);
nor U9859 (N_9859,N_9717,N_9686);
nor U9860 (N_9860,N_9584,N_9736);
xor U9861 (N_9861,N_9539,N_9677);
and U9862 (N_9862,N_9703,N_9604);
xnor U9863 (N_9863,N_9556,N_9656);
xnor U9864 (N_9864,N_9748,N_9528);
nor U9865 (N_9865,N_9625,N_9601);
and U9866 (N_9866,N_9595,N_9618);
xor U9867 (N_9867,N_9586,N_9626);
and U9868 (N_9868,N_9591,N_9502);
or U9869 (N_9869,N_9620,N_9728);
nor U9870 (N_9870,N_9676,N_9508);
and U9871 (N_9871,N_9681,N_9610);
xnor U9872 (N_9872,N_9723,N_9693);
nand U9873 (N_9873,N_9632,N_9538);
and U9874 (N_9874,N_9733,N_9678);
and U9875 (N_9875,N_9630,N_9675);
nand U9876 (N_9876,N_9637,N_9653);
xnor U9877 (N_9877,N_9582,N_9707);
or U9878 (N_9878,N_9530,N_9535);
or U9879 (N_9879,N_9596,N_9585);
nor U9880 (N_9880,N_9574,N_9554);
nor U9881 (N_9881,N_9547,N_9613);
nor U9882 (N_9882,N_9741,N_9560);
xor U9883 (N_9883,N_9551,N_9702);
nor U9884 (N_9884,N_9717,N_9684);
xor U9885 (N_9885,N_9683,N_9737);
nor U9886 (N_9886,N_9553,N_9581);
and U9887 (N_9887,N_9600,N_9710);
nor U9888 (N_9888,N_9501,N_9693);
nor U9889 (N_9889,N_9712,N_9569);
and U9890 (N_9890,N_9714,N_9727);
or U9891 (N_9891,N_9674,N_9517);
and U9892 (N_9892,N_9556,N_9566);
xnor U9893 (N_9893,N_9635,N_9706);
nand U9894 (N_9894,N_9541,N_9709);
nor U9895 (N_9895,N_9697,N_9548);
nand U9896 (N_9896,N_9649,N_9709);
and U9897 (N_9897,N_9515,N_9565);
and U9898 (N_9898,N_9550,N_9630);
or U9899 (N_9899,N_9741,N_9746);
nand U9900 (N_9900,N_9640,N_9740);
or U9901 (N_9901,N_9556,N_9584);
or U9902 (N_9902,N_9742,N_9652);
xor U9903 (N_9903,N_9690,N_9606);
or U9904 (N_9904,N_9725,N_9711);
and U9905 (N_9905,N_9682,N_9677);
and U9906 (N_9906,N_9550,N_9731);
nand U9907 (N_9907,N_9658,N_9668);
or U9908 (N_9908,N_9656,N_9669);
and U9909 (N_9909,N_9554,N_9612);
nand U9910 (N_9910,N_9531,N_9532);
or U9911 (N_9911,N_9682,N_9727);
nand U9912 (N_9912,N_9536,N_9596);
nand U9913 (N_9913,N_9705,N_9535);
or U9914 (N_9914,N_9567,N_9557);
and U9915 (N_9915,N_9717,N_9707);
and U9916 (N_9916,N_9667,N_9650);
or U9917 (N_9917,N_9587,N_9560);
and U9918 (N_9918,N_9630,N_9722);
xor U9919 (N_9919,N_9708,N_9686);
and U9920 (N_9920,N_9588,N_9605);
xor U9921 (N_9921,N_9526,N_9554);
and U9922 (N_9922,N_9571,N_9676);
nand U9923 (N_9923,N_9622,N_9747);
or U9924 (N_9924,N_9525,N_9542);
nor U9925 (N_9925,N_9544,N_9534);
nand U9926 (N_9926,N_9574,N_9607);
and U9927 (N_9927,N_9736,N_9516);
nand U9928 (N_9928,N_9685,N_9621);
and U9929 (N_9929,N_9561,N_9662);
nor U9930 (N_9930,N_9640,N_9649);
or U9931 (N_9931,N_9588,N_9511);
nor U9932 (N_9932,N_9507,N_9724);
nor U9933 (N_9933,N_9711,N_9591);
nor U9934 (N_9934,N_9516,N_9545);
or U9935 (N_9935,N_9728,N_9661);
and U9936 (N_9936,N_9537,N_9517);
nand U9937 (N_9937,N_9713,N_9588);
nor U9938 (N_9938,N_9500,N_9666);
and U9939 (N_9939,N_9548,N_9647);
nand U9940 (N_9940,N_9606,N_9501);
nor U9941 (N_9941,N_9672,N_9617);
and U9942 (N_9942,N_9573,N_9534);
and U9943 (N_9943,N_9743,N_9631);
xor U9944 (N_9944,N_9571,N_9748);
and U9945 (N_9945,N_9601,N_9612);
and U9946 (N_9946,N_9713,N_9748);
and U9947 (N_9947,N_9516,N_9638);
nor U9948 (N_9948,N_9620,N_9667);
or U9949 (N_9949,N_9696,N_9608);
nor U9950 (N_9950,N_9557,N_9688);
nand U9951 (N_9951,N_9503,N_9742);
nand U9952 (N_9952,N_9588,N_9597);
nand U9953 (N_9953,N_9664,N_9602);
xor U9954 (N_9954,N_9635,N_9596);
nand U9955 (N_9955,N_9500,N_9695);
nor U9956 (N_9956,N_9684,N_9688);
and U9957 (N_9957,N_9656,N_9623);
nor U9958 (N_9958,N_9671,N_9507);
or U9959 (N_9959,N_9566,N_9537);
and U9960 (N_9960,N_9598,N_9698);
nor U9961 (N_9961,N_9597,N_9672);
or U9962 (N_9962,N_9695,N_9561);
xnor U9963 (N_9963,N_9621,N_9665);
or U9964 (N_9964,N_9686,N_9694);
nor U9965 (N_9965,N_9735,N_9682);
and U9966 (N_9966,N_9598,N_9516);
nor U9967 (N_9967,N_9623,N_9683);
and U9968 (N_9968,N_9602,N_9614);
and U9969 (N_9969,N_9598,N_9730);
or U9970 (N_9970,N_9628,N_9522);
nor U9971 (N_9971,N_9558,N_9625);
nand U9972 (N_9972,N_9677,N_9684);
nor U9973 (N_9973,N_9548,N_9547);
and U9974 (N_9974,N_9736,N_9643);
or U9975 (N_9975,N_9517,N_9659);
or U9976 (N_9976,N_9694,N_9710);
or U9977 (N_9977,N_9571,N_9530);
nor U9978 (N_9978,N_9652,N_9662);
nor U9979 (N_9979,N_9580,N_9749);
and U9980 (N_9980,N_9511,N_9551);
nor U9981 (N_9981,N_9747,N_9683);
nand U9982 (N_9982,N_9527,N_9742);
and U9983 (N_9983,N_9509,N_9550);
nand U9984 (N_9984,N_9749,N_9659);
nand U9985 (N_9985,N_9612,N_9591);
and U9986 (N_9986,N_9615,N_9697);
xor U9987 (N_9987,N_9666,N_9527);
nand U9988 (N_9988,N_9535,N_9508);
nand U9989 (N_9989,N_9537,N_9611);
and U9990 (N_9990,N_9563,N_9539);
xnor U9991 (N_9991,N_9620,N_9699);
nand U9992 (N_9992,N_9546,N_9634);
or U9993 (N_9993,N_9634,N_9547);
and U9994 (N_9994,N_9729,N_9741);
or U9995 (N_9995,N_9646,N_9503);
or U9996 (N_9996,N_9676,N_9585);
and U9997 (N_9997,N_9674,N_9529);
and U9998 (N_9998,N_9669,N_9648);
xnor U9999 (N_9999,N_9719,N_9509);
and U10000 (N_10000,N_9936,N_9846);
xnor U10001 (N_10001,N_9770,N_9979);
xnor U10002 (N_10002,N_9808,N_9918);
nor U10003 (N_10003,N_9791,N_9914);
nand U10004 (N_10004,N_9804,N_9815);
nor U10005 (N_10005,N_9952,N_9935);
or U10006 (N_10006,N_9887,N_9903);
xnor U10007 (N_10007,N_9776,N_9839);
or U10008 (N_10008,N_9906,N_9872);
nor U10009 (N_10009,N_9995,N_9809);
or U10010 (N_10010,N_9897,N_9997);
or U10011 (N_10011,N_9949,N_9852);
xnor U10012 (N_10012,N_9807,N_9834);
nand U10013 (N_10013,N_9948,N_9963);
or U10014 (N_10014,N_9898,N_9976);
nand U10015 (N_10015,N_9837,N_9970);
nor U10016 (N_10016,N_9891,N_9858);
and U10017 (N_10017,N_9845,N_9781);
xor U10018 (N_10018,N_9971,N_9895);
and U10019 (N_10019,N_9962,N_9864);
and U10020 (N_10020,N_9853,N_9783);
nor U10021 (N_10021,N_9944,N_9857);
nand U10022 (N_10022,N_9925,N_9802);
nor U10023 (N_10023,N_9828,N_9848);
xor U10024 (N_10024,N_9987,N_9803);
nor U10025 (N_10025,N_9762,N_9819);
nand U10026 (N_10026,N_9978,N_9821);
xnor U10027 (N_10027,N_9943,N_9933);
nor U10028 (N_10028,N_9830,N_9827);
xor U10029 (N_10029,N_9939,N_9924);
and U10030 (N_10030,N_9896,N_9875);
xor U10031 (N_10031,N_9940,N_9928);
or U10032 (N_10032,N_9879,N_9871);
and U10033 (N_10033,N_9765,N_9905);
nand U10034 (N_10034,N_9934,N_9882);
nand U10035 (N_10035,N_9812,N_9790);
or U10036 (N_10036,N_9958,N_9824);
nand U10037 (N_10037,N_9868,N_9767);
or U10038 (N_10038,N_9913,N_9937);
and U10039 (N_10039,N_9922,N_9794);
and U10040 (N_10040,N_9917,N_9910);
xor U10041 (N_10041,N_9855,N_9793);
nand U10042 (N_10042,N_9880,N_9862);
xor U10043 (N_10043,N_9780,N_9873);
and U10044 (N_10044,N_9960,N_9863);
nor U10045 (N_10045,N_9769,N_9929);
nand U10046 (N_10046,N_9972,N_9854);
nand U10047 (N_10047,N_9957,N_9801);
and U10048 (N_10048,N_9805,N_9763);
or U10049 (N_10049,N_9760,N_9982);
nor U10050 (N_10050,N_9799,N_9822);
and U10051 (N_10051,N_9927,N_9994);
and U10052 (N_10052,N_9867,N_9959);
xnor U10053 (N_10053,N_9876,N_9985);
xor U10054 (N_10054,N_9861,N_9849);
nand U10055 (N_10055,N_9814,N_9768);
nor U10056 (N_10056,N_9823,N_9993);
xor U10057 (N_10057,N_9850,N_9986);
nand U10058 (N_10058,N_9788,N_9946);
nor U10059 (N_10059,N_9800,N_9974);
nand U10060 (N_10060,N_9990,N_9992);
xnor U10061 (N_10061,N_9953,N_9885);
nand U10062 (N_10062,N_9832,N_9980);
nand U10063 (N_10063,N_9789,N_9916);
nor U10064 (N_10064,N_9865,N_9951);
nand U10065 (N_10065,N_9878,N_9966);
nand U10066 (N_10066,N_9899,N_9919);
nor U10067 (N_10067,N_9969,N_9838);
xor U10068 (N_10068,N_9842,N_9900);
nand U10069 (N_10069,N_9818,N_9826);
nand U10070 (N_10070,N_9816,N_9908);
xnor U10071 (N_10071,N_9947,N_9806);
or U10072 (N_10072,N_9920,N_9792);
xor U10073 (N_10073,N_9941,N_9923);
nand U10074 (N_10074,N_9964,N_9938);
nand U10075 (N_10075,N_9890,N_9989);
nor U10076 (N_10076,N_9798,N_9844);
or U10077 (N_10077,N_9945,N_9911);
nand U10078 (N_10078,N_9831,N_9870);
nand U10079 (N_10079,N_9775,N_9886);
and U10080 (N_10080,N_9753,N_9983);
nand U10081 (N_10081,N_9892,N_9786);
nand U10082 (N_10082,N_9764,N_9965);
nand U10083 (N_10083,N_9778,N_9881);
and U10084 (N_10084,N_9796,N_9766);
or U10085 (N_10085,N_9785,N_9784);
xnor U10086 (N_10086,N_9755,N_9893);
and U10087 (N_10087,N_9884,N_9869);
and U10088 (N_10088,N_9926,N_9930);
and U10089 (N_10089,N_9988,N_9797);
nand U10090 (N_10090,N_9759,N_9779);
and U10091 (N_10091,N_9757,N_9968);
nand U10092 (N_10092,N_9782,N_9889);
nor U10093 (N_10093,N_9975,N_9902);
xor U10094 (N_10094,N_9756,N_9977);
nor U10095 (N_10095,N_9811,N_9847);
nor U10096 (N_10096,N_9904,N_9877);
xor U10097 (N_10097,N_9973,N_9829);
and U10098 (N_10098,N_9909,N_9866);
nor U10099 (N_10099,N_9773,N_9754);
or U10100 (N_10100,N_9901,N_9888);
nand U10101 (N_10101,N_9984,N_9774);
or U10102 (N_10102,N_9915,N_9955);
and U10103 (N_10103,N_9825,N_9787);
nor U10104 (N_10104,N_9750,N_9956);
or U10105 (N_10105,N_9772,N_9981);
nand U10106 (N_10106,N_9967,N_9777);
nor U10107 (N_10107,N_9840,N_9996);
nor U10108 (N_10108,N_9836,N_9931);
and U10109 (N_10109,N_9856,N_9795);
nand U10110 (N_10110,N_9833,N_9961);
and U10111 (N_10111,N_9841,N_9813);
nand U10112 (N_10112,N_9810,N_9907);
nand U10113 (N_10113,N_9758,N_9942);
nand U10114 (N_10114,N_9874,N_9843);
nor U10115 (N_10115,N_9991,N_9859);
xnor U10116 (N_10116,N_9912,N_9752);
or U10117 (N_10117,N_9820,N_9998);
nand U10118 (N_10118,N_9954,N_9921);
xnor U10119 (N_10119,N_9771,N_9851);
and U10120 (N_10120,N_9932,N_9817);
or U10121 (N_10121,N_9751,N_9950);
nand U10122 (N_10122,N_9860,N_9883);
xnor U10123 (N_10123,N_9894,N_9999);
or U10124 (N_10124,N_9761,N_9835);
xor U10125 (N_10125,N_9972,N_9975);
xor U10126 (N_10126,N_9920,N_9817);
nor U10127 (N_10127,N_9950,N_9958);
nor U10128 (N_10128,N_9941,N_9959);
nand U10129 (N_10129,N_9949,N_9820);
and U10130 (N_10130,N_9819,N_9889);
nand U10131 (N_10131,N_9829,N_9957);
and U10132 (N_10132,N_9895,N_9821);
nor U10133 (N_10133,N_9980,N_9970);
or U10134 (N_10134,N_9975,N_9838);
xnor U10135 (N_10135,N_9919,N_9786);
and U10136 (N_10136,N_9925,N_9929);
and U10137 (N_10137,N_9781,N_9864);
and U10138 (N_10138,N_9814,N_9974);
nand U10139 (N_10139,N_9814,N_9812);
or U10140 (N_10140,N_9836,N_9950);
nor U10141 (N_10141,N_9984,N_9772);
nand U10142 (N_10142,N_9899,N_9838);
xor U10143 (N_10143,N_9936,N_9780);
and U10144 (N_10144,N_9911,N_9822);
or U10145 (N_10145,N_9970,N_9806);
nand U10146 (N_10146,N_9973,N_9800);
xnor U10147 (N_10147,N_9853,N_9978);
nor U10148 (N_10148,N_9809,N_9871);
or U10149 (N_10149,N_9786,N_9918);
nor U10150 (N_10150,N_9954,N_9750);
xor U10151 (N_10151,N_9765,N_9773);
nand U10152 (N_10152,N_9786,N_9981);
or U10153 (N_10153,N_9815,N_9886);
or U10154 (N_10154,N_9982,N_9833);
and U10155 (N_10155,N_9840,N_9879);
nand U10156 (N_10156,N_9915,N_9902);
or U10157 (N_10157,N_9839,N_9842);
nand U10158 (N_10158,N_9758,N_9872);
nor U10159 (N_10159,N_9855,N_9945);
xnor U10160 (N_10160,N_9795,N_9756);
xnor U10161 (N_10161,N_9931,N_9887);
nand U10162 (N_10162,N_9968,N_9987);
xor U10163 (N_10163,N_9871,N_9948);
nand U10164 (N_10164,N_9831,N_9840);
nand U10165 (N_10165,N_9857,N_9760);
and U10166 (N_10166,N_9793,N_9816);
xor U10167 (N_10167,N_9910,N_9919);
nand U10168 (N_10168,N_9921,N_9807);
xnor U10169 (N_10169,N_9922,N_9957);
nand U10170 (N_10170,N_9782,N_9801);
or U10171 (N_10171,N_9828,N_9904);
and U10172 (N_10172,N_9843,N_9888);
or U10173 (N_10173,N_9903,N_9985);
nand U10174 (N_10174,N_9797,N_9765);
nand U10175 (N_10175,N_9805,N_9966);
or U10176 (N_10176,N_9982,N_9875);
xnor U10177 (N_10177,N_9946,N_9876);
nor U10178 (N_10178,N_9785,N_9781);
or U10179 (N_10179,N_9925,N_9958);
xnor U10180 (N_10180,N_9948,N_9866);
xor U10181 (N_10181,N_9973,N_9772);
xor U10182 (N_10182,N_9779,N_9910);
and U10183 (N_10183,N_9775,N_9801);
xor U10184 (N_10184,N_9791,N_9886);
xnor U10185 (N_10185,N_9912,N_9952);
nand U10186 (N_10186,N_9981,N_9939);
xor U10187 (N_10187,N_9995,N_9874);
nand U10188 (N_10188,N_9979,N_9793);
and U10189 (N_10189,N_9953,N_9900);
and U10190 (N_10190,N_9859,N_9861);
xor U10191 (N_10191,N_9780,N_9852);
and U10192 (N_10192,N_9825,N_9754);
and U10193 (N_10193,N_9873,N_9958);
xnor U10194 (N_10194,N_9932,N_9888);
nor U10195 (N_10195,N_9996,N_9990);
nand U10196 (N_10196,N_9750,N_9829);
nand U10197 (N_10197,N_9890,N_9835);
nor U10198 (N_10198,N_9902,N_9865);
and U10199 (N_10199,N_9781,N_9916);
nand U10200 (N_10200,N_9935,N_9884);
nand U10201 (N_10201,N_9765,N_9911);
or U10202 (N_10202,N_9951,N_9891);
and U10203 (N_10203,N_9962,N_9937);
or U10204 (N_10204,N_9966,N_9983);
xnor U10205 (N_10205,N_9800,N_9781);
xnor U10206 (N_10206,N_9992,N_9778);
or U10207 (N_10207,N_9752,N_9850);
nand U10208 (N_10208,N_9950,N_9839);
and U10209 (N_10209,N_9775,N_9875);
or U10210 (N_10210,N_9792,N_9981);
nand U10211 (N_10211,N_9887,N_9872);
nor U10212 (N_10212,N_9869,N_9825);
xor U10213 (N_10213,N_9919,N_9969);
and U10214 (N_10214,N_9875,N_9953);
and U10215 (N_10215,N_9860,N_9888);
nor U10216 (N_10216,N_9995,N_9864);
nor U10217 (N_10217,N_9844,N_9931);
or U10218 (N_10218,N_9867,N_9892);
and U10219 (N_10219,N_9951,N_9977);
or U10220 (N_10220,N_9971,N_9841);
xnor U10221 (N_10221,N_9961,N_9854);
or U10222 (N_10222,N_9970,N_9790);
nor U10223 (N_10223,N_9772,N_9853);
or U10224 (N_10224,N_9901,N_9967);
xnor U10225 (N_10225,N_9760,N_9751);
nand U10226 (N_10226,N_9765,N_9866);
nor U10227 (N_10227,N_9935,N_9888);
xnor U10228 (N_10228,N_9980,N_9814);
and U10229 (N_10229,N_9906,N_9827);
nor U10230 (N_10230,N_9864,N_9791);
nand U10231 (N_10231,N_9991,N_9795);
xor U10232 (N_10232,N_9785,N_9823);
nor U10233 (N_10233,N_9950,N_9846);
nand U10234 (N_10234,N_9945,N_9878);
xor U10235 (N_10235,N_9889,N_9954);
or U10236 (N_10236,N_9853,N_9863);
xor U10237 (N_10237,N_9825,N_9867);
nor U10238 (N_10238,N_9853,N_9813);
and U10239 (N_10239,N_9941,N_9878);
nand U10240 (N_10240,N_9981,N_9751);
xor U10241 (N_10241,N_9981,N_9754);
nand U10242 (N_10242,N_9927,N_9824);
nor U10243 (N_10243,N_9974,N_9781);
and U10244 (N_10244,N_9861,N_9979);
or U10245 (N_10245,N_9893,N_9971);
or U10246 (N_10246,N_9979,N_9987);
nor U10247 (N_10247,N_9967,N_9948);
nor U10248 (N_10248,N_9772,N_9827);
or U10249 (N_10249,N_9859,N_9968);
xor U10250 (N_10250,N_10218,N_10053);
and U10251 (N_10251,N_10066,N_10247);
nand U10252 (N_10252,N_10123,N_10051);
xnor U10253 (N_10253,N_10194,N_10141);
nand U10254 (N_10254,N_10032,N_10006);
or U10255 (N_10255,N_10188,N_10169);
nand U10256 (N_10256,N_10087,N_10225);
nor U10257 (N_10257,N_10039,N_10146);
or U10258 (N_10258,N_10115,N_10208);
nor U10259 (N_10259,N_10185,N_10048);
or U10260 (N_10260,N_10090,N_10160);
or U10261 (N_10261,N_10096,N_10076);
nand U10262 (N_10262,N_10065,N_10178);
or U10263 (N_10263,N_10072,N_10157);
and U10264 (N_10264,N_10224,N_10055);
xor U10265 (N_10265,N_10081,N_10068);
nor U10266 (N_10266,N_10176,N_10173);
or U10267 (N_10267,N_10165,N_10223);
and U10268 (N_10268,N_10153,N_10029);
or U10269 (N_10269,N_10004,N_10159);
and U10270 (N_10270,N_10212,N_10041);
nand U10271 (N_10271,N_10040,N_10246);
nor U10272 (N_10272,N_10136,N_10080);
or U10273 (N_10273,N_10104,N_10062);
nor U10274 (N_10274,N_10018,N_10144);
or U10275 (N_10275,N_10163,N_10181);
nor U10276 (N_10276,N_10150,N_10149);
xor U10277 (N_10277,N_10139,N_10003);
or U10278 (N_10278,N_10238,N_10005);
nor U10279 (N_10279,N_10120,N_10151);
and U10280 (N_10280,N_10046,N_10043);
nand U10281 (N_10281,N_10241,N_10024);
nand U10282 (N_10282,N_10098,N_10064);
and U10283 (N_10283,N_10113,N_10045);
nor U10284 (N_10284,N_10199,N_10170);
or U10285 (N_10285,N_10002,N_10112);
nor U10286 (N_10286,N_10110,N_10122);
xnor U10287 (N_10287,N_10240,N_10059);
or U10288 (N_10288,N_10226,N_10017);
xor U10289 (N_10289,N_10000,N_10042);
or U10290 (N_10290,N_10184,N_10130);
nor U10291 (N_10291,N_10128,N_10154);
nand U10292 (N_10292,N_10237,N_10177);
nand U10293 (N_10293,N_10044,N_10101);
xor U10294 (N_10294,N_10027,N_10008);
and U10295 (N_10295,N_10099,N_10058);
nand U10296 (N_10296,N_10168,N_10093);
nor U10297 (N_10297,N_10155,N_10033);
nor U10298 (N_10298,N_10019,N_10190);
xor U10299 (N_10299,N_10119,N_10095);
nor U10300 (N_10300,N_10228,N_10158);
xnor U10301 (N_10301,N_10227,N_10232);
xnor U10302 (N_10302,N_10147,N_10083);
or U10303 (N_10303,N_10105,N_10001);
xnor U10304 (N_10304,N_10013,N_10089);
and U10305 (N_10305,N_10152,N_10088);
and U10306 (N_10306,N_10200,N_10061);
or U10307 (N_10307,N_10197,N_10242);
nor U10308 (N_10308,N_10100,N_10191);
and U10309 (N_10309,N_10107,N_10217);
nand U10310 (N_10310,N_10245,N_10121);
nor U10311 (N_10311,N_10162,N_10057);
nand U10312 (N_10312,N_10063,N_10210);
nand U10313 (N_10313,N_10108,N_10180);
nor U10314 (N_10314,N_10067,N_10209);
xnor U10315 (N_10315,N_10140,N_10243);
and U10316 (N_10316,N_10114,N_10195);
nor U10317 (N_10317,N_10248,N_10126);
and U10318 (N_10318,N_10131,N_10175);
nor U10319 (N_10319,N_10049,N_10117);
xor U10320 (N_10320,N_10182,N_10164);
xor U10321 (N_10321,N_10030,N_10085);
nor U10322 (N_10322,N_10103,N_10235);
and U10323 (N_10323,N_10229,N_10127);
or U10324 (N_10324,N_10023,N_10097);
xor U10325 (N_10325,N_10236,N_10193);
and U10326 (N_10326,N_10054,N_10021);
or U10327 (N_10327,N_10198,N_10221);
nand U10328 (N_10328,N_10034,N_10028);
and U10329 (N_10329,N_10213,N_10074);
nor U10330 (N_10330,N_10204,N_10222);
nand U10331 (N_10331,N_10125,N_10206);
nand U10332 (N_10332,N_10082,N_10249);
xor U10333 (N_10333,N_10143,N_10022);
nor U10334 (N_10334,N_10137,N_10145);
xnor U10335 (N_10335,N_10075,N_10202);
nor U10336 (N_10336,N_10201,N_10025);
and U10337 (N_10337,N_10133,N_10069);
xnor U10338 (N_10338,N_10038,N_10186);
and U10339 (N_10339,N_10047,N_10205);
or U10340 (N_10340,N_10239,N_10091);
xor U10341 (N_10341,N_10070,N_10118);
xnor U10342 (N_10342,N_10031,N_10134);
nor U10343 (N_10343,N_10060,N_10015);
or U10344 (N_10344,N_10215,N_10124);
xnor U10345 (N_10345,N_10092,N_10189);
or U10346 (N_10346,N_10230,N_10037);
nand U10347 (N_10347,N_10231,N_10116);
or U10348 (N_10348,N_10010,N_10196);
nand U10349 (N_10349,N_10129,N_10148);
nand U10350 (N_10350,N_10161,N_10174);
xnor U10351 (N_10351,N_10179,N_10079);
or U10352 (N_10352,N_10167,N_10211);
or U10353 (N_10353,N_10172,N_10102);
nand U10354 (N_10354,N_10012,N_10214);
nor U10355 (N_10355,N_10166,N_10106);
nand U10356 (N_10356,N_10035,N_10156);
and U10357 (N_10357,N_10207,N_10183);
and U10358 (N_10358,N_10135,N_10220);
xor U10359 (N_10359,N_10234,N_10016);
xor U10360 (N_10360,N_10219,N_10084);
nand U10361 (N_10361,N_10036,N_10111);
or U10362 (N_10362,N_10109,N_10014);
nor U10363 (N_10363,N_10009,N_10138);
nand U10364 (N_10364,N_10026,N_10052);
or U10365 (N_10365,N_10007,N_10086);
nor U10366 (N_10366,N_10203,N_10142);
or U10367 (N_10367,N_10132,N_10071);
nand U10368 (N_10368,N_10171,N_10233);
nand U10369 (N_10369,N_10077,N_10187);
xnor U10370 (N_10370,N_10011,N_10020);
nor U10371 (N_10371,N_10078,N_10073);
xor U10372 (N_10372,N_10056,N_10216);
nor U10373 (N_10373,N_10192,N_10050);
xor U10374 (N_10374,N_10094,N_10244);
nand U10375 (N_10375,N_10191,N_10016);
or U10376 (N_10376,N_10107,N_10221);
xnor U10377 (N_10377,N_10001,N_10057);
or U10378 (N_10378,N_10139,N_10193);
nor U10379 (N_10379,N_10217,N_10167);
xor U10380 (N_10380,N_10145,N_10174);
xor U10381 (N_10381,N_10139,N_10024);
or U10382 (N_10382,N_10088,N_10033);
nor U10383 (N_10383,N_10173,N_10079);
xnor U10384 (N_10384,N_10231,N_10019);
and U10385 (N_10385,N_10161,N_10188);
and U10386 (N_10386,N_10050,N_10122);
or U10387 (N_10387,N_10217,N_10188);
nor U10388 (N_10388,N_10242,N_10210);
nand U10389 (N_10389,N_10208,N_10170);
or U10390 (N_10390,N_10004,N_10216);
nand U10391 (N_10391,N_10041,N_10000);
and U10392 (N_10392,N_10120,N_10006);
and U10393 (N_10393,N_10206,N_10245);
and U10394 (N_10394,N_10078,N_10238);
xor U10395 (N_10395,N_10117,N_10047);
or U10396 (N_10396,N_10165,N_10073);
and U10397 (N_10397,N_10190,N_10088);
xor U10398 (N_10398,N_10086,N_10064);
xor U10399 (N_10399,N_10086,N_10054);
or U10400 (N_10400,N_10094,N_10114);
nand U10401 (N_10401,N_10201,N_10233);
or U10402 (N_10402,N_10210,N_10115);
xnor U10403 (N_10403,N_10200,N_10231);
nand U10404 (N_10404,N_10006,N_10138);
and U10405 (N_10405,N_10029,N_10179);
nand U10406 (N_10406,N_10001,N_10084);
xnor U10407 (N_10407,N_10052,N_10161);
xnor U10408 (N_10408,N_10242,N_10158);
or U10409 (N_10409,N_10173,N_10139);
and U10410 (N_10410,N_10128,N_10001);
xor U10411 (N_10411,N_10040,N_10209);
xnor U10412 (N_10412,N_10032,N_10179);
or U10413 (N_10413,N_10222,N_10003);
nor U10414 (N_10414,N_10035,N_10217);
xnor U10415 (N_10415,N_10074,N_10244);
and U10416 (N_10416,N_10083,N_10128);
nor U10417 (N_10417,N_10117,N_10143);
nand U10418 (N_10418,N_10082,N_10221);
xnor U10419 (N_10419,N_10229,N_10126);
xnor U10420 (N_10420,N_10028,N_10039);
or U10421 (N_10421,N_10029,N_10245);
nor U10422 (N_10422,N_10245,N_10085);
xnor U10423 (N_10423,N_10203,N_10055);
nor U10424 (N_10424,N_10063,N_10064);
nand U10425 (N_10425,N_10060,N_10211);
nor U10426 (N_10426,N_10005,N_10249);
nor U10427 (N_10427,N_10079,N_10101);
and U10428 (N_10428,N_10240,N_10205);
xnor U10429 (N_10429,N_10059,N_10188);
nor U10430 (N_10430,N_10026,N_10091);
and U10431 (N_10431,N_10040,N_10162);
or U10432 (N_10432,N_10133,N_10181);
and U10433 (N_10433,N_10175,N_10129);
and U10434 (N_10434,N_10029,N_10189);
xnor U10435 (N_10435,N_10249,N_10154);
nand U10436 (N_10436,N_10211,N_10058);
or U10437 (N_10437,N_10055,N_10052);
and U10438 (N_10438,N_10168,N_10049);
xor U10439 (N_10439,N_10114,N_10115);
and U10440 (N_10440,N_10214,N_10186);
and U10441 (N_10441,N_10155,N_10211);
xnor U10442 (N_10442,N_10177,N_10155);
nor U10443 (N_10443,N_10089,N_10150);
or U10444 (N_10444,N_10136,N_10219);
nor U10445 (N_10445,N_10134,N_10162);
xnor U10446 (N_10446,N_10169,N_10178);
xnor U10447 (N_10447,N_10246,N_10086);
or U10448 (N_10448,N_10056,N_10117);
nor U10449 (N_10449,N_10218,N_10104);
or U10450 (N_10450,N_10244,N_10053);
or U10451 (N_10451,N_10038,N_10008);
or U10452 (N_10452,N_10233,N_10048);
nor U10453 (N_10453,N_10131,N_10009);
xnor U10454 (N_10454,N_10208,N_10182);
nor U10455 (N_10455,N_10083,N_10177);
nand U10456 (N_10456,N_10070,N_10056);
xnor U10457 (N_10457,N_10155,N_10066);
nor U10458 (N_10458,N_10050,N_10013);
or U10459 (N_10459,N_10111,N_10162);
and U10460 (N_10460,N_10146,N_10022);
or U10461 (N_10461,N_10064,N_10215);
nand U10462 (N_10462,N_10073,N_10076);
nand U10463 (N_10463,N_10128,N_10103);
xor U10464 (N_10464,N_10128,N_10032);
xor U10465 (N_10465,N_10168,N_10134);
and U10466 (N_10466,N_10163,N_10081);
or U10467 (N_10467,N_10143,N_10041);
or U10468 (N_10468,N_10235,N_10220);
and U10469 (N_10469,N_10136,N_10009);
and U10470 (N_10470,N_10246,N_10024);
nor U10471 (N_10471,N_10000,N_10220);
or U10472 (N_10472,N_10056,N_10069);
or U10473 (N_10473,N_10049,N_10183);
nor U10474 (N_10474,N_10170,N_10248);
xor U10475 (N_10475,N_10215,N_10079);
nor U10476 (N_10476,N_10018,N_10172);
and U10477 (N_10477,N_10094,N_10034);
xor U10478 (N_10478,N_10057,N_10237);
or U10479 (N_10479,N_10144,N_10057);
xor U10480 (N_10480,N_10126,N_10079);
nand U10481 (N_10481,N_10228,N_10202);
nand U10482 (N_10482,N_10168,N_10174);
xor U10483 (N_10483,N_10129,N_10146);
or U10484 (N_10484,N_10153,N_10071);
nand U10485 (N_10485,N_10118,N_10093);
nand U10486 (N_10486,N_10154,N_10000);
nor U10487 (N_10487,N_10237,N_10145);
nand U10488 (N_10488,N_10062,N_10219);
or U10489 (N_10489,N_10013,N_10072);
nor U10490 (N_10490,N_10065,N_10224);
xor U10491 (N_10491,N_10172,N_10014);
nand U10492 (N_10492,N_10125,N_10247);
nor U10493 (N_10493,N_10000,N_10162);
and U10494 (N_10494,N_10074,N_10006);
or U10495 (N_10495,N_10228,N_10168);
and U10496 (N_10496,N_10045,N_10165);
or U10497 (N_10497,N_10032,N_10068);
nor U10498 (N_10498,N_10095,N_10173);
or U10499 (N_10499,N_10231,N_10044);
and U10500 (N_10500,N_10457,N_10480);
or U10501 (N_10501,N_10445,N_10436);
or U10502 (N_10502,N_10491,N_10268);
xnor U10503 (N_10503,N_10287,N_10282);
or U10504 (N_10504,N_10418,N_10252);
or U10505 (N_10505,N_10396,N_10384);
nor U10506 (N_10506,N_10309,N_10322);
xor U10507 (N_10507,N_10275,N_10332);
nor U10508 (N_10508,N_10378,N_10336);
nand U10509 (N_10509,N_10493,N_10297);
xor U10510 (N_10510,N_10355,N_10345);
nand U10511 (N_10511,N_10293,N_10284);
nand U10512 (N_10512,N_10385,N_10476);
or U10513 (N_10513,N_10393,N_10485);
or U10514 (N_10514,N_10292,N_10419);
nor U10515 (N_10515,N_10352,N_10375);
or U10516 (N_10516,N_10438,N_10269);
nand U10517 (N_10517,N_10306,N_10323);
xor U10518 (N_10518,N_10456,N_10435);
or U10519 (N_10519,N_10363,N_10424);
or U10520 (N_10520,N_10423,N_10390);
nand U10521 (N_10521,N_10434,N_10343);
xnor U10522 (N_10522,N_10443,N_10466);
nor U10523 (N_10523,N_10326,N_10404);
xnor U10524 (N_10524,N_10462,N_10260);
nor U10525 (N_10525,N_10376,N_10356);
nand U10526 (N_10526,N_10471,N_10362);
and U10527 (N_10527,N_10474,N_10380);
nor U10528 (N_10528,N_10458,N_10486);
or U10529 (N_10529,N_10450,N_10351);
nor U10530 (N_10530,N_10431,N_10420);
nand U10531 (N_10531,N_10400,N_10488);
nor U10532 (N_10532,N_10310,N_10273);
nand U10533 (N_10533,N_10461,N_10330);
nor U10534 (N_10534,N_10300,N_10286);
and U10535 (N_10535,N_10394,N_10426);
nand U10536 (N_10536,N_10366,N_10428);
xor U10537 (N_10537,N_10421,N_10283);
and U10538 (N_10538,N_10379,N_10319);
nand U10539 (N_10539,N_10484,N_10329);
xor U10540 (N_10540,N_10274,N_10392);
or U10541 (N_10541,N_10361,N_10251);
nor U10542 (N_10542,N_10307,N_10279);
nand U10543 (N_10543,N_10311,N_10403);
nor U10544 (N_10544,N_10453,N_10441);
and U10545 (N_10545,N_10440,N_10409);
xnor U10546 (N_10546,N_10401,N_10406);
xor U10547 (N_10547,N_10398,N_10377);
nor U10548 (N_10548,N_10271,N_10359);
or U10549 (N_10549,N_10315,N_10328);
nand U10550 (N_10550,N_10254,N_10460);
nand U10551 (N_10551,N_10371,N_10342);
nand U10552 (N_10552,N_10285,N_10391);
nand U10553 (N_10553,N_10429,N_10439);
nor U10554 (N_10554,N_10427,N_10302);
and U10555 (N_10555,N_10316,N_10369);
or U10556 (N_10556,N_10447,N_10314);
or U10557 (N_10557,N_10432,N_10313);
nor U10558 (N_10558,N_10477,N_10270);
or U10559 (N_10559,N_10280,N_10259);
nand U10560 (N_10560,N_10386,N_10367);
or U10561 (N_10561,N_10261,N_10290);
xor U10562 (N_10562,N_10444,N_10495);
and U10563 (N_10563,N_10478,N_10305);
nor U10564 (N_10564,N_10492,N_10463);
nand U10565 (N_10565,N_10276,N_10320);
nand U10566 (N_10566,N_10494,N_10483);
nand U10567 (N_10567,N_10372,N_10324);
nor U10568 (N_10568,N_10277,N_10451);
or U10569 (N_10569,N_10469,N_10364);
nor U10570 (N_10570,N_10365,N_10317);
and U10571 (N_10571,N_10454,N_10373);
nor U10572 (N_10572,N_10383,N_10308);
and U10573 (N_10573,N_10425,N_10301);
and U10574 (N_10574,N_10250,N_10387);
or U10575 (N_10575,N_10449,N_10422);
nor U10576 (N_10576,N_10470,N_10312);
nor U10577 (N_10577,N_10294,N_10490);
or U10578 (N_10578,N_10331,N_10341);
and U10579 (N_10579,N_10253,N_10459);
nand U10580 (N_10580,N_10263,N_10498);
xnor U10581 (N_10581,N_10281,N_10472);
and U10582 (N_10582,N_10481,N_10338);
nor U10583 (N_10583,N_10412,N_10414);
xor U10584 (N_10584,N_10448,N_10321);
or U10585 (N_10585,N_10468,N_10257);
nor U10586 (N_10586,N_10304,N_10357);
or U10587 (N_10587,N_10416,N_10405);
nand U10588 (N_10588,N_10295,N_10399);
or U10589 (N_10589,N_10267,N_10303);
nand U10590 (N_10590,N_10288,N_10397);
xnor U10591 (N_10591,N_10415,N_10289);
or U10592 (N_10592,N_10467,N_10354);
and U10593 (N_10593,N_10446,N_10382);
xnor U10594 (N_10594,N_10465,N_10347);
nor U10595 (N_10595,N_10299,N_10255);
xnor U10596 (N_10596,N_10346,N_10497);
or U10597 (N_10597,N_10370,N_10442);
nand U10598 (N_10598,N_10298,N_10487);
nor U10599 (N_10599,N_10475,N_10411);
xnor U10600 (N_10600,N_10407,N_10413);
nand U10601 (N_10601,N_10258,N_10464);
xnor U10602 (N_10602,N_10395,N_10499);
and U10603 (N_10603,N_10344,N_10374);
and U10604 (N_10604,N_10318,N_10430);
xnor U10605 (N_10605,N_10262,N_10272);
xnor U10606 (N_10606,N_10381,N_10339);
and U10607 (N_10607,N_10489,N_10340);
and U10608 (N_10608,N_10433,N_10350);
and U10609 (N_10609,N_10353,N_10388);
nor U10610 (N_10610,N_10325,N_10264);
nand U10611 (N_10611,N_10335,N_10473);
nor U10612 (N_10612,N_10437,N_10389);
xnor U10613 (N_10613,N_10296,N_10452);
and U10614 (N_10614,N_10496,N_10358);
nor U10615 (N_10615,N_10256,N_10265);
or U10616 (N_10616,N_10278,N_10402);
nor U10617 (N_10617,N_10417,N_10482);
or U10618 (N_10618,N_10349,N_10291);
nand U10619 (N_10619,N_10333,N_10368);
or U10620 (N_10620,N_10337,N_10360);
nor U10621 (N_10621,N_10455,N_10408);
nor U10622 (N_10622,N_10479,N_10266);
xnor U10623 (N_10623,N_10334,N_10348);
and U10624 (N_10624,N_10327,N_10410);
and U10625 (N_10625,N_10332,N_10495);
xor U10626 (N_10626,N_10338,N_10381);
nand U10627 (N_10627,N_10266,N_10466);
nor U10628 (N_10628,N_10349,N_10254);
nand U10629 (N_10629,N_10414,N_10386);
nand U10630 (N_10630,N_10310,N_10399);
or U10631 (N_10631,N_10301,N_10283);
xor U10632 (N_10632,N_10484,N_10405);
nand U10633 (N_10633,N_10442,N_10361);
nand U10634 (N_10634,N_10475,N_10400);
xor U10635 (N_10635,N_10469,N_10276);
nor U10636 (N_10636,N_10296,N_10390);
or U10637 (N_10637,N_10498,N_10437);
or U10638 (N_10638,N_10383,N_10418);
xnor U10639 (N_10639,N_10258,N_10256);
and U10640 (N_10640,N_10258,N_10445);
or U10641 (N_10641,N_10391,N_10367);
nor U10642 (N_10642,N_10312,N_10414);
nand U10643 (N_10643,N_10310,N_10394);
nand U10644 (N_10644,N_10303,N_10461);
xor U10645 (N_10645,N_10389,N_10349);
nor U10646 (N_10646,N_10475,N_10279);
xnor U10647 (N_10647,N_10372,N_10333);
nor U10648 (N_10648,N_10387,N_10459);
nor U10649 (N_10649,N_10329,N_10322);
or U10650 (N_10650,N_10362,N_10309);
and U10651 (N_10651,N_10309,N_10471);
xor U10652 (N_10652,N_10259,N_10463);
and U10653 (N_10653,N_10415,N_10382);
and U10654 (N_10654,N_10435,N_10406);
xor U10655 (N_10655,N_10485,N_10301);
nor U10656 (N_10656,N_10414,N_10433);
xor U10657 (N_10657,N_10409,N_10372);
or U10658 (N_10658,N_10499,N_10469);
and U10659 (N_10659,N_10387,N_10363);
and U10660 (N_10660,N_10478,N_10336);
and U10661 (N_10661,N_10283,N_10468);
nand U10662 (N_10662,N_10442,N_10484);
or U10663 (N_10663,N_10466,N_10337);
xor U10664 (N_10664,N_10435,N_10356);
xnor U10665 (N_10665,N_10467,N_10393);
and U10666 (N_10666,N_10277,N_10350);
nor U10667 (N_10667,N_10288,N_10339);
xor U10668 (N_10668,N_10309,N_10269);
and U10669 (N_10669,N_10494,N_10433);
nand U10670 (N_10670,N_10358,N_10321);
and U10671 (N_10671,N_10299,N_10365);
and U10672 (N_10672,N_10437,N_10335);
xnor U10673 (N_10673,N_10392,N_10301);
nand U10674 (N_10674,N_10281,N_10456);
or U10675 (N_10675,N_10353,N_10260);
or U10676 (N_10676,N_10404,N_10337);
nor U10677 (N_10677,N_10373,N_10426);
xnor U10678 (N_10678,N_10260,N_10474);
xor U10679 (N_10679,N_10374,N_10251);
or U10680 (N_10680,N_10429,N_10317);
and U10681 (N_10681,N_10376,N_10462);
and U10682 (N_10682,N_10275,N_10304);
nand U10683 (N_10683,N_10470,N_10412);
and U10684 (N_10684,N_10273,N_10356);
nand U10685 (N_10685,N_10466,N_10276);
or U10686 (N_10686,N_10461,N_10365);
or U10687 (N_10687,N_10282,N_10400);
xnor U10688 (N_10688,N_10275,N_10411);
xor U10689 (N_10689,N_10493,N_10401);
and U10690 (N_10690,N_10288,N_10382);
or U10691 (N_10691,N_10269,N_10489);
nor U10692 (N_10692,N_10384,N_10439);
and U10693 (N_10693,N_10382,N_10358);
xor U10694 (N_10694,N_10410,N_10390);
nor U10695 (N_10695,N_10312,N_10323);
xnor U10696 (N_10696,N_10362,N_10405);
nand U10697 (N_10697,N_10300,N_10285);
nand U10698 (N_10698,N_10360,N_10406);
and U10699 (N_10699,N_10333,N_10453);
nor U10700 (N_10700,N_10285,N_10443);
nor U10701 (N_10701,N_10402,N_10374);
nand U10702 (N_10702,N_10359,N_10431);
or U10703 (N_10703,N_10495,N_10263);
xnor U10704 (N_10704,N_10422,N_10404);
nand U10705 (N_10705,N_10456,N_10419);
xnor U10706 (N_10706,N_10393,N_10480);
and U10707 (N_10707,N_10374,N_10407);
nor U10708 (N_10708,N_10368,N_10482);
nor U10709 (N_10709,N_10352,N_10353);
or U10710 (N_10710,N_10475,N_10493);
nand U10711 (N_10711,N_10258,N_10347);
nor U10712 (N_10712,N_10454,N_10307);
nor U10713 (N_10713,N_10294,N_10356);
nor U10714 (N_10714,N_10434,N_10332);
nor U10715 (N_10715,N_10424,N_10478);
nor U10716 (N_10716,N_10488,N_10443);
xor U10717 (N_10717,N_10386,N_10498);
and U10718 (N_10718,N_10475,N_10393);
xnor U10719 (N_10719,N_10402,N_10408);
nand U10720 (N_10720,N_10484,N_10354);
nand U10721 (N_10721,N_10336,N_10357);
and U10722 (N_10722,N_10402,N_10443);
and U10723 (N_10723,N_10376,N_10377);
or U10724 (N_10724,N_10318,N_10264);
nor U10725 (N_10725,N_10457,N_10428);
xnor U10726 (N_10726,N_10352,N_10312);
and U10727 (N_10727,N_10250,N_10479);
xor U10728 (N_10728,N_10491,N_10381);
xor U10729 (N_10729,N_10253,N_10353);
nor U10730 (N_10730,N_10302,N_10289);
or U10731 (N_10731,N_10265,N_10312);
nor U10732 (N_10732,N_10489,N_10256);
nor U10733 (N_10733,N_10372,N_10433);
xnor U10734 (N_10734,N_10418,N_10265);
xor U10735 (N_10735,N_10350,N_10429);
and U10736 (N_10736,N_10479,N_10301);
nand U10737 (N_10737,N_10492,N_10254);
nor U10738 (N_10738,N_10291,N_10486);
nand U10739 (N_10739,N_10342,N_10489);
and U10740 (N_10740,N_10353,N_10351);
or U10741 (N_10741,N_10404,N_10270);
xor U10742 (N_10742,N_10301,N_10302);
nand U10743 (N_10743,N_10359,N_10252);
or U10744 (N_10744,N_10339,N_10313);
or U10745 (N_10745,N_10443,N_10280);
xnor U10746 (N_10746,N_10404,N_10477);
nand U10747 (N_10747,N_10454,N_10319);
and U10748 (N_10748,N_10413,N_10298);
or U10749 (N_10749,N_10455,N_10459);
xor U10750 (N_10750,N_10613,N_10680);
and U10751 (N_10751,N_10685,N_10590);
nor U10752 (N_10752,N_10711,N_10654);
nand U10753 (N_10753,N_10732,N_10672);
xor U10754 (N_10754,N_10655,N_10589);
xor U10755 (N_10755,N_10551,N_10548);
nor U10756 (N_10756,N_10625,N_10521);
and U10757 (N_10757,N_10631,N_10679);
nor U10758 (N_10758,N_10695,N_10620);
nor U10759 (N_10759,N_10530,N_10678);
nand U10760 (N_10760,N_10571,N_10673);
and U10761 (N_10761,N_10607,N_10684);
and U10762 (N_10762,N_10581,N_10504);
nand U10763 (N_10763,N_10708,N_10526);
xor U10764 (N_10764,N_10611,N_10618);
and U10765 (N_10765,N_10587,N_10597);
nand U10766 (N_10766,N_10682,N_10698);
and U10767 (N_10767,N_10591,N_10586);
and U10768 (N_10768,N_10520,N_10659);
or U10769 (N_10769,N_10668,N_10709);
and U10770 (N_10770,N_10585,N_10535);
xnor U10771 (N_10771,N_10693,N_10675);
nand U10772 (N_10772,N_10663,N_10576);
nor U10773 (N_10773,N_10734,N_10578);
nand U10774 (N_10774,N_10536,N_10588);
xor U10775 (N_10775,N_10544,N_10584);
nor U10776 (N_10776,N_10700,N_10735);
and U10777 (N_10777,N_10593,N_10603);
or U10778 (N_10778,N_10653,N_10543);
or U10779 (N_10779,N_10583,N_10564);
or U10780 (N_10780,N_10533,N_10748);
or U10781 (N_10781,N_10612,N_10624);
xnor U10782 (N_10782,N_10633,N_10522);
xnor U10783 (N_10783,N_10649,N_10537);
or U10784 (N_10784,N_10572,N_10691);
xnor U10785 (N_10785,N_10740,N_10729);
nor U10786 (N_10786,N_10517,N_10651);
or U10787 (N_10787,N_10547,N_10558);
or U10788 (N_10788,N_10745,N_10686);
nand U10789 (N_10789,N_10630,N_10639);
nand U10790 (N_10790,N_10565,N_10688);
or U10791 (N_10791,N_10519,N_10608);
or U10792 (N_10792,N_10738,N_10502);
and U10793 (N_10793,N_10515,N_10637);
xor U10794 (N_10794,N_10616,N_10661);
or U10795 (N_10795,N_10542,N_10665);
xor U10796 (N_10796,N_10614,N_10666);
nand U10797 (N_10797,N_10710,N_10712);
and U10798 (N_10798,N_10531,N_10501);
or U10799 (N_10799,N_10622,N_10638);
or U10800 (N_10800,N_10539,N_10619);
and U10801 (N_10801,N_10636,N_10528);
and U10802 (N_10802,N_10677,N_10648);
and U10803 (N_10803,N_10557,N_10697);
nand U10804 (N_10804,N_10687,N_10561);
xnor U10805 (N_10805,N_10609,N_10601);
and U10806 (N_10806,N_10525,N_10615);
and U10807 (N_10807,N_10541,N_10580);
xor U10808 (N_10808,N_10599,N_10706);
nand U10809 (N_10809,N_10643,N_10594);
nand U10810 (N_10810,N_10634,N_10570);
and U10811 (N_10811,N_10715,N_10716);
or U10812 (N_10812,N_10721,N_10598);
xor U10813 (N_10813,N_10646,N_10546);
and U10814 (N_10814,N_10555,N_10644);
nand U10815 (N_10815,N_10577,N_10562);
nand U10816 (N_10816,N_10699,N_10600);
xnor U10817 (N_10817,N_10736,N_10647);
and U10818 (N_10818,N_10746,N_10662);
or U10819 (N_10819,N_10725,N_10730);
nor U10820 (N_10820,N_10742,N_10690);
or U10821 (N_10821,N_10595,N_10642);
or U10822 (N_10822,N_10670,N_10617);
nor U10823 (N_10823,N_10556,N_10575);
nand U10824 (N_10824,N_10726,N_10683);
or U10825 (N_10825,N_10605,N_10692);
nor U10826 (N_10826,N_10724,N_10568);
nor U10827 (N_10827,N_10705,N_10579);
xnor U10828 (N_10828,N_10563,N_10744);
nor U10829 (N_10829,N_10566,N_10731);
or U10830 (N_10830,N_10719,N_10534);
nor U10831 (N_10831,N_10669,N_10714);
nand U10832 (N_10832,N_10658,N_10552);
and U10833 (N_10833,N_10626,N_10505);
or U10834 (N_10834,N_10507,N_10553);
nor U10835 (N_10835,N_10733,N_10723);
xor U10836 (N_10836,N_10676,N_10627);
xor U10837 (N_10837,N_10529,N_10737);
xor U10838 (N_10838,N_10720,N_10703);
nand U10839 (N_10839,N_10621,N_10549);
nor U10840 (N_10840,N_10518,N_10704);
nor U10841 (N_10841,N_10569,N_10508);
xnor U10842 (N_10842,N_10727,N_10606);
nor U10843 (N_10843,N_10524,N_10689);
and U10844 (N_10844,N_10671,N_10660);
and U10845 (N_10845,N_10667,N_10510);
or U10846 (N_10846,N_10527,N_10707);
nand U10847 (N_10847,N_10604,N_10645);
nand U10848 (N_10848,N_10538,N_10717);
or U10849 (N_10849,N_10596,N_10506);
nand U10850 (N_10850,N_10623,N_10500);
nand U10851 (N_10851,N_10523,N_10657);
and U10852 (N_10852,N_10629,N_10503);
and U10853 (N_10853,N_10674,N_10514);
nor U10854 (N_10854,N_10532,N_10664);
xor U10855 (N_10855,N_10739,N_10610);
xor U10856 (N_10856,N_10545,N_10747);
xor U10857 (N_10857,N_10513,N_10702);
nor U10858 (N_10858,N_10641,N_10722);
and U10859 (N_10859,N_10635,N_10602);
and U10860 (N_10860,N_10516,N_10554);
or U10861 (N_10861,N_10582,N_10749);
xnor U10862 (N_10862,N_10560,N_10640);
nand U10863 (N_10863,N_10573,N_10741);
and U10864 (N_10864,N_10743,N_10511);
or U10865 (N_10865,N_10540,N_10550);
or U10866 (N_10866,N_10701,N_10574);
or U10867 (N_10867,N_10650,N_10728);
or U10868 (N_10868,N_10696,N_10718);
nor U10869 (N_10869,N_10713,N_10512);
nor U10870 (N_10870,N_10656,N_10652);
nor U10871 (N_10871,N_10628,N_10592);
xor U10872 (N_10872,N_10632,N_10559);
xnor U10873 (N_10873,N_10567,N_10694);
or U10874 (N_10874,N_10509,N_10681);
and U10875 (N_10875,N_10566,N_10522);
nand U10876 (N_10876,N_10590,N_10581);
or U10877 (N_10877,N_10525,N_10705);
xnor U10878 (N_10878,N_10660,N_10632);
nor U10879 (N_10879,N_10733,N_10510);
xnor U10880 (N_10880,N_10579,N_10643);
nand U10881 (N_10881,N_10578,N_10733);
nand U10882 (N_10882,N_10710,N_10733);
nand U10883 (N_10883,N_10548,N_10722);
or U10884 (N_10884,N_10502,N_10636);
or U10885 (N_10885,N_10503,N_10618);
or U10886 (N_10886,N_10610,N_10700);
and U10887 (N_10887,N_10711,N_10638);
nor U10888 (N_10888,N_10532,N_10602);
or U10889 (N_10889,N_10525,N_10702);
xnor U10890 (N_10890,N_10538,N_10746);
nand U10891 (N_10891,N_10586,N_10538);
nand U10892 (N_10892,N_10728,N_10711);
nor U10893 (N_10893,N_10618,N_10699);
nor U10894 (N_10894,N_10611,N_10664);
or U10895 (N_10895,N_10520,N_10563);
nand U10896 (N_10896,N_10513,N_10549);
xnor U10897 (N_10897,N_10663,N_10580);
xor U10898 (N_10898,N_10713,N_10741);
xor U10899 (N_10899,N_10509,N_10678);
and U10900 (N_10900,N_10669,N_10696);
or U10901 (N_10901,N_10638,N_10606);
nand U10902 (N_10902,N_10545,N_10714);
xor U10903 (N_10903,N_10653,N_10673);
or U10904 (N_10904,N_10734,N_10714);
nand U10905 (N_10905,N_10507,N_10669);
and U10906 (N_10906,N_10524,N_10528);
nand U10907 (N_10907,N_10557,N_10532);
nor U10908 (N_10908,N_10716,N_10694);
nor U10909 (N_10909,N_10538,N_10527);
nor U10910 (N_10910,N_10537,N_10531);
or U10911 (N_10911,N_10612,N_10656);
nor U10912 (N_10912,N_10601,N_10552);
and U10913 (N_10913,N_10641,N_10665);
or U10914 (N_10914,N_10735,N_10571);
and U10915 (N_10915,N_10670,N_10735);
xor U10916 (N_10916,N_10693,N_10511);
nor U10917 (N_10917,N_10724,N_10627);
xnor U10918 (N_10918,N_10677,N_10744);
and U10919 (N_10919,N_10626,N_10724);
xnor U10920 (N_10920,N_10536,N_10504);
or U10921 (N_10921,N_10626,N_10586);
xnor U10922 (N_10922,N_10503,N_10738);
xor U10923 (N_10923,N_10620,N_10503);
or U10924 (N_10924,N_10614,N_10678);
xor U10925 (N_10925,N_10675,N_10649);
nand U10926 (N_10926,N_10718,N_10554);
xnor U10927 (N_10927,N_10568,N_10599);
and U10928 (N_10928,N_10721,N_10594);
or U10929 (N_10929,N_10643,N_10641);
or U10930 (N_10930,N_10608,N_10543);
nor U10931 (N_10931,N_10717,N_10588);
nand U10932 (N_10932,N_10566,N_10654);
or U10933 (N_10933,N_10693,N_10564);
nor U10934 (N_10934,N_10573,N_10716);
xor U10935 (N_10935,N_10507,N_10668);
and U10936 (N_10936,N_10540,N_10580);
nand U10937 (N_10937,N_10616,N_10685);
or U10938 (N_10938,N_10740,N_10693);
and U10939 (N_10939,N_10693,N_10526);
and U10940 (N_10940,N_10530,N_10726);
or U10941 (N_10941,N_10741,N_10735);
nor U10942 (N_10942,N_10713,N_10538);
nor U10943 (N_10943,N_10527,N_10617);
nand U10944 (N_10944,N_10679,N_10613);
and U10945 (N_10945,N_10500,N_10712);
xnor U10946 (N_10946,N_10554,N_10734);
xor U10947 (N_10947,N_10678,N_10551);
or U10948 (N_10948,N_10511,N_10512);
nor U10949 (N_10949,N_10600,N_10712);
or U10950 (N_10950,N_10607,N_10545);
nor U10951 (N_10951,N_10703,N_10745);
or U10952 (N_10952,N_10650,N_10577);
nand U10953 (N_10953,N_10692,N_10705);
xnor U10954 (N_10954,N_10565,N_10620);
or U10955 (N_10955,N_10560,N_10672);
and U10956 (N_10956,N_10545,N_10647);
xor U10957 (N_10957,N_10616,N_10720);
xor U10958 (N_10958,N_10655,N_10624);
nor U10959 (N_10959,N_10518,N_10664);
or U10960 (N_10960,N_10733,N_10703);
nand U10961 (N_10961,N_10602,N_10607);
nor U10962 (N_10962,N_10603,N_10601);
nand U10963 (N_10963,N_10692,N_10524);
xnor U10964 (N_10964,N_10630,N_10685);
and U10965 (N_10965,N_10744,N_10653);
nand U10966 (N_10966,N_10665,N_10654);
xnor U10967 (N_10967,N_10646,N_10573);
nand U10968 (N_10968,N_10638,N_10661);
and U10969 (N_10969,N_10686,N_10671);
nor U10970 (N_10970,N_10670,N_10534);
and U10971 (N_10971,N_10555,N_10665);
and U10972 (N_10972,N_10579,N_10731);
nand U10973 (N_10973,N_10749,N_10604);
and U10974 (N_10974,N_10678,N_10616);
nand U10975 (N_10975,N_10513,N_10644);
xnor U10976 (N_10976,N_10707,N_10616);
nor U10977 (N_10977,N_10582,N_10536);
xnor U10978 (N_10978,N_10514,N_10570);
xnor U10979 (N_10979,N_10562,N_10518);
or U10980 (N_10980,N_10676,N_10603);
xor U10981 (N_10981,N_10567,N_10661);
or U10982 (N_10982,N_10573,N_10723);
nor U10983 (N_10983,N_10613,N_10558);
nand U10984 (N_10984,N_10596,N_10658);
nor U10985 (N_10985,N_10579,N_10672);
xor U10986 (N_10986,N_10626,N_10649);
xnor U10987 (N_10987,N_10555,N_10659);
or U10988 (N_10988,N_10717,N_10562);
nor U10989 (N_10989,N_10741,N_10698);
and U10990 (N_10990,N_10693,N_10664);
or U10991 (N_10991,N_10652,N_10543);
or U10992 (N_10992,N_10707,N_10629);
or U10993 (N_10993,N_10629,N_10738);
or U10994 (N_10994,N_10622,N_10587);
and U10995 (N_10995,N_10581,N_10707);
or U10996 (N_10996,N_10529,N_10690);
or U10997 (N_10997,N_10706,N_10620);
nand U10998 (N_10998,N_10669,N_10736);
xnor U10999 (N_10999,N_10611,N_10621);
xnor U11000 (N_11000,N_10809,N_10887);
or U11001 (N_11001,N_10935,N_10995);
nor U11002 (N_11002,N_10855,N_10997);
xor U11003 (N_11003,N_10974,N_10802);
nor U11004 (N_11004,N_10996,N_10991);
xor U11005 (N_11005,N_10852,N_10756);
or U11006 (N_11006,N_10897,N_10786);
and U11007 (N_11007,N_10955,N_10796);
nand U11008 (N_11008,N_10872,N_10947);
xor U11009 (N_11009,N_10779,N_10854);
nor U11010 (N_11010,N_10839,N_10797);
nor U11011 (N_11011,N_10999,N_10882);
and U11012 (N_11012,N_10994,N_10856);
nor U11013 (N_11013,N_10965,N_10903);
nand U11014 (N_11014,N_10926,N_10795);
nor U11015 (N_11015,N_10895,N_10884);
and U11016 (N_11016,N_10777,N_10964);
or U11017 (N_11017,N_10859,N_10820);
nor U11018 (N_11018,N_10973,N_10932);
and U11019 (N_11019,N_10939,N_10837);
nor U11020 (N_11020,N_10845,N_10780);
xnor U11021 (N_11021,N_10771,N_10773);
nor U11022 (N_11022,N_10946,N_10883);
or U11023 (N_11023,N_10767,N_10826);
nand U11024 (N_11024,N_10900,N_10823);
xor U11025 (N_11025,N_10967,N_10979);
nand U11026 (N_11026,N_10908,N_10987);
nor U11027 (N_11027,N_10805,N_10891);
nand U11028 (N_11028,N_10817,N_10831);
nand U11029 (N_11029,N_10940,N_10954);
nor U11030 (N_11030,N_10869,N_10880);
nand U11031 (N_11031,N_10915,N_10844);
nand U11032 (N_11032,N_10772,N_10770);
nand U11033 (N_11033,N_10933,N_10972);
nor U11034 (N_11034,N_10789,N_10881);
and U11035 (N_11035,N_10899,N_10835);
nor U11036 (N_11036,N_10792,N_10936);
and U11037 (N_11037,N_10788,N_10815);
or U11038 (N_11038,N_10998,N_10871);
or U11039 (N_11039,N_10879,N_10941);
and U11040 (N_11040,N_10866,N_10948);
and U11041 (N_11041,N_10867,N_10912);
nand U11042 (N_11042,N_10898,N_10864);
or U11043 (N_11043,N_10827,N_10982);
or U11044 (N_11044,N_10878,N_10976);
or U11045 (N_11045,N_10853,N_10988);
xor U11046 (N_11046,N_10757,N_10759);
xor U11047 (N_11047,N_10916,N_10752);
nor U11048 (N_11048,N_10896,N_10834);
xnor U11049 (N_11049,N_10787,N_10782);
and U11050 (N_11050,N_10840,N_10841);
and U11051 (N_11051,N_10793,N_10975);
nand U11052 (N_11052,N_10818,N_10848);
nand U11053 (N_11053,N_10930,N_10825);
or U11054 (N_11054,N_10813,N_10894);
xor U11055 (N_11055,N_10924,N_10901);
and U11056 (N_11056,N_10763,N_10775);
nor U11057 (N_11057,N_10784,N_10816);
or U11058 (N_11058,N_10931,N_10798);
or U11059 (N_11059,N_10806,N_10846);
nor U11060 (N_11060,N_10785,N_10914);
nor U11061 (N_11061,N_10937,N_10783);
nand U11062 (N_11062,N_10918,N_10943);
nand U11063 (N_11063,N_10858,N_10873);
and U11064 (N_11064,N_10919,N_10790);
xor U11065 (N_11065,N_10934,N_10968);
and U11066 (N_11066,N_10870,N_10944);
nor U11067 (N_11067,N_10923,N_10851);
nor U11068 (N_11068,N_10992,N_10925);
xnor U11069 (N_11069,N_10857,N_10875);
and U11070 (N_11070,N_10833,N_10886);
or U11071 (N_11071,N_10760,N_10910);
nor U11072 (N_11072,N_10978,N_10791);
nand U11073 (N_11073,N_10989,N_10830);
nand U11074 (N_11074,N_10832,N_10913);
xnor U11075 (N_11075,N_10893,N_10753);
nand U11076 (N_11076,N_10774,N_10981);
or U11077 (N_11077,N_10980,N_10849);
and U11078 (N_11078,N_10765,N_10890);
or U11079 (N_11079,N_10807,N_10824);
nand U11080 (N_11080,N_10768,N_10750);
or U11081 (N_11081,N_10889,N_10838);
nand U11082 (N_11082,N_10874,N_10755);
and U11083 (N_11083,N_10892,N_10960);
xor U11084 (N_11084,N_10794,N_10909);
nor U11085 (N_11085,N_10758,N_10984);
xor U11086 (N_11086,N_10819,N_10761);
xor U11087 (N_11087,N_10904,N_10938);
and U11088 (N_11088,N_10956,N_10842);
and U11089 (N_11089,N_10917,N_10971);
nor U11090 (N_11090,N_10958,N_10993);
nor U11091 (N_11091,N_10906,N_10804);
xnor U11092 (N_11092,N_10754,N_10862);
nor U11093 (N_11093,N_10990,N_10865);
nor U11094 (N_11094,N_10877,N_10762);
or U11095 (N_11095,N_10843,N_10850);
or U11096 (N_11096,N_10902,N_10907);
or U11097 (N_11097,N_10966,N_10921);
or U11098 (N_11098,N_10814,N_10985);
or U11099 (N_11099,N_10952,N_10847);
xnor U11100 (N_11100,N_10927,N_10969);
xor U11101 (N_11101,N_10829,N_10778);
nand U11102 (N_11102,N_10953,N_10803);
nand U11103 (N_11103,N_10959,N_10957);
and U11104 (N_11104,N_10800,N_10970);
xor U11105 (N_11105,N_10861,N_10950);
xnor U11106 (N_11106,N_10885,N_10822);
nand U11107 (N_11107,N_10799,N_10836);
nand U11108 (N_11108,N_10828,N_10977);
nor U11109 (N_11109,N_10801,N_10945);
nand U11110 (N_11110,N_10983,N_10942);
nor U11111 (N_11111,N_10920,N_10769);
xnor U11112 (N_11112,N_10821,N_10808);
or U11113 (N_11113,N_10949,N_10911);
and U11114 (N_11114,N_10810,N_10922);
nand U11115 (N_11115,N_10961,N_10951);
nor U11116 (N_11116,N_10929,N_10928);
nor U11117 (N_11117,N_10811,N_10766);
xnor U11118 (N_11118,N_10888,N_10963);
nor U11119 (N_11119,N_10781,N_10986);
nand U11120 (N_11120,N_10863,N_10812);
nor U11121 (N_11121,N_10751,N_10764);
xnor U11122 (N_11122,N_10876,N_10776);
nor U11123 (N_11123,N_10868,N_10860);
xnor U11124 (N_11124,N_10905,N_10962);
nand U11125 (N_11125,N_10768,N_10966);
xnor U11126 (N_11126,N_10817,N_10833);
xor U11127 (N_11127,N_10812,N_10963);
or U11128 (N_11128,N_10819,N_10812);
and U11129 (N_11129,N_10789,N_10893);
and U11130 (N_11130,N_10901,N_10917);
xnor U11131 (N_11131,N_10877,N_10898);
nor U11132 (N_11132,N_10992,N_10947);
xnor U11133 (N_11133,N_10771,N_10941);
nor U11134 (N_11134,N_10887,N_10976);
nand U11135 (N_11135,N_10759,N_10788);
xor U11136 (N_11136,N_10987,N_10993);
or U11137 (N_11137,N_10798,N_10823);
or U11138 (N_11138,N_10805,N_10866);
nand U11139 (N_11139,N_10752,N_10796);
nand U11140 (N_11140,N_10865,N_10756);
or U11141 (N_11141,N_10778,N_10756);
xnor U11142 (N_11142,N_10878,N_10771);
nand U11143 (N_11143,N_10938,N_10762);
or U11144 (N_11144,N_10942,N_10879);
or U11145 (N_11145,N_10770,N_10757);
or U11146 (N_11146,N_10937,N_10775);
nor U11147 (N_11147,N_10812,N_10826);
xnor U11148 (N_11148,N_10940,N_10760);
xor U11149 (N_11149,N_10968,N_10837);
xor U11150 (N_11150,N_10767,N_10995);
or U11151 (N_11151,N_10836,N_10813);
nand U11152 (N_11152,N_10949,N_10756);
xnor U11153 (N_11153,N_10828,N_10832);
nand U11154 (N_11154,N_10781,N_10774);
and U11155 (N_11155,N_10932,N_10924);
or U11156 (N_11156,N_10755,N_10939);
xor U11157 (N_11157,N_10871,N_10795);
or U11158 (N_11158,N_10892,N_10753);
or U11159 (N_11159,N_10905,N_10954);
or U11160 (N_11160,N_10906,N_10831);
or U11161 (N_11161,N_10831,N_10913);
or U11162 (N_11162,N_10792,N_10935);
xor U11163 (N_11163,N_10784,N_10910);
or U11164 (N_11164,N_10996,N_10976);
or U11165 (N_11165,N_10964,N_10986);
nor U11166 (N_11166,N_10884,N_10830);
and U11167 (N_11167,N_10967,N_10939);
xnor U11168 (N_11168,N_10890,N_10920);
nand U11169 (N_11169,N_10828,N_10844);
or U11170 (N_11170,N_10813,N_10775);
and U11171 (N_11171,N_10896,N_10855);
xnor U11172 (N_11172,N_10823,N_10961);
xnor U11173 (N_11173,N_10899,N_10938);
xor U11174 (N_11174,N_10812,N_10906);
and U11175 (N_11175,N_10761,N_10965);
xor U11176 (N_11176,N_10839,N_10942);
nor U11177 (N_11177,N_10844,N_10767);
nand U11178 (N_11178,N_10870,N_10958);
nand U11179 (N_11179,N_10804,N_10963);
and U11180 (N_11180,N_10943,N_10755);
nand U11181 (N_11181,N_10889,N_10983);
nand U11182 (N_11182,N_10861,N_10850);
or U11183 (N_11183,N_10790,N_10955);
and U11184 (N_11184,N_10878,N_10992);
and U11185 (N_11185,N_10986,N_10963);
nor U11186 (N_11186,N_10847,N_10823);
nand U11187 (N_11187,N_10876,N_10832);
and U11188 (N_11188,N_10966,N_10916);
xnor U11189 (N_11189,N_10973,N_10869);
nand U11190 (N_11190,N_10752,N_10925);
xor U11191 (N_11191,N_10945,N_10980);
nand U11192 (N_11192,N_10925,N_10761);
nand U11193 (N_11193,N_10897,N_10957);
nor U11194 (N_11194,N_10841,N_10797);
nand U11195 (N_11195,N_10775,N_10906);
or U11196 (N_11196,N_10896,N_10774);
and U11197 (N_11197,N_10801,N_10792);
nor U11198 (N_11198,N_10999,N_10994);
nand U11199 (N_11199,N_10837,N_10993);
nand U11200 (N_11200,N_10977,N_10861);
or U11201 (N_11201,N_10925,N_10756);
nor U11202 (N_11202,N_10792,N_10901);
and U11203 (N_11203,N_10770,N_10968);
and U11204 (N_11204,N_10970,N_10960);
or U11205 (N_11205,N_10776,N_10836);
xnor U11206 (N_11206,N_10914,N_10884);
or U11207 (N_11207,N_10891,N_10924);
and U11208 (N_11208,N_10816,N_10846);
xor U11209 (N_11209,N_10926,N_10791);
xnor U11210 (N_11210,N_10897,N_10995);
xor U11211 (N_11211,N_10971,N_10968);
nand U11212 (N_11212,N_10907,N_10994);
nand U11213 (N_11213,N_10935,N_10967);
and U11214 (N_11214,N_10918,N_10891);
and U11215 (N_11215,N_10888,N_10951);
nand U11216 (N_11216,N_10874,N_10927);
nand U11217 (N_11217,N_10885,N_10888);
and U11218 (N_11218,N_10896,N_10756);
or U11219 (N_11219,N_10756,N_10810);
nand U11220 (N_11220,N_10831,N_10807);
and U11221 (N_11221,N_10878,N_10889);
nand U11222 (N_11222,N_10917,N_10923);
nor U11223 (N_11223,N_10814,N_10912);
xnor U11224 (N_11224,N_10857,N_10918);
xnor U11225 (N_11225,N_10755,N_10863);
nor U11226 (N_11226,N_10810,N_10953);
nand U11227 (N_11227,N_10882,N_10963);
xnor U11228 (N_11228,N_10895,N_10832);
or U11229 (N_11229,N_10787,N_10808);
or U11230 (N_11230,N_10951,N_10857);
nand U11231 (N_11231,N_10905,N_10977);
xor U11232 (N_11232,N_10859,N_10808);
xor U11233 (N_11233,N_10898,N_10938);
and U11234 (N_11234,N_10977,N_10884);
nor U11235 (N_11235,N_10790,N_10922);
nor U11236 (N_11236,N_10828,N_10917);
xor U11237 (N_11237,N_10814,N_10836);
or U11238 (N_11238,N_10996,N_10899);
nand U11239 (N_11239,N_10871,N_10858);
or U11240 (N_11240,N_10780,N_10781);
xor U11241 (N_11241,N_10896,N_10929);
or U11242 (N_11242,N_10983,N_10805);
or U11243 (N_11243,N_10759,N_10824);
nand U11244 (N_11244,N_10865,N_10889);
or U11245 (N_11245,N_10829,N_10960);
xor U11246 (N_11246,N_10761,N_10842);
and U11247 (N_11247,N_10961,N_10842);
nor U11248 (N_11248,N_10928,N_10876);
nand U11249 (N_11249,N_10896,N_10768);
xor U11250 (N_11250,N_11248,N_11215);
nor U11251 (N_11251,N_11245,N_11121);
or U11252 (N_11252,N_11075,N_11012);
xor U11253 (N_11253,N_11080,N_11065);
and U11254 (N_11254,N_11182,N_11064);
xnor U11255 (N_11255,N_11137,N_11060);
and U11256 (N_11256,N_11239,N_11123);
xor U11257 (N_11257,N_11050,N_11092);
or U11258 (N_11258,N_11247,N_11026);
xor U11259 (N_11259,N_11113,N_11188);
and U11260 (N_11260,N_11218,N_11073);
or U11261 (N_11261,N_11184,N_11224);
xnor U11262 (N_11262,N_11093,N_11104);
or U11263 (N_11263,N_11020,N_11095);
nor U11264 (N_11264,N_11109,N_11046);
xor U11265 (N_11265,N_11070,N_11030);
xnor U11266 (N_11266,N_11015,N_11219);
nand U11267 (N_11267,N_11003,N_11047);
nand U11268 (N_11268,N_11209,N_11086);
xnor U11269 (N_11269,N_11194,N_11161);
xnor U11270 (N_11270,N_11119,N_11189);
nor U11271 (N_11271,N_11227,N_11231);
and U11272 (N_11272,N_11179,N_11134);
nand U11273 (N_11273,N_11208,N_11053);
or U11274 (N_11274,N_11001,N_11027);
nand U11275 (N_11275,N_11101,N_11203);
or U11276 (N_11276,N_11116,N_11160);
nand U11277 (N_11277,N_11005,N_11082);
nor U11278 (N_11278,N_11112,N_11062);
or U11279 (N_11279,N_11089,N_11130);
nor U11280 (N_11280,N_11202,N_11229);
nand U11281 (N_11281,N_11057,N_11055);
xnor U11282 (N_11282,N_11226,N_11139);
nor U11283 (N_11283,N_11185,N_11138);
nand U11284 (N_11284,N_11158,N_11187);
nand U11285 (N_11285,N_11155,N_11083);
or U11286 (N_11286,N_11122,N_11151);
and U11287 (N_11287,N_11129,N_11036);
xnor U11288 (N_11288,N_11141,N_11156);
nor U11289 (N_11289,N_11240,N_11068);
or U11290 (N_11290,N_11197,N_11178);
or U11291 (N_11291,N_11222,N_11180);
xnor U11292 (N_11292,N_11132,N_11225);
and U11293 (N_11293,N_11033,N_11107);
nand U11294 (N_11294,N_11214,N_11085);
or U11295 (N_11295,N_11166,N_11096);
xnor U11296 (N_11296,N_11090,N_11002);
or U11297 (N_11297,N_11131,N_11106);
nor U11298 (N_11298,N_11169,N_11146);
nor U11299 (N_11299,N_11198,N_11152);
xnor U11300 (N_11300,N_11031,N_11032);
nor U11301 (N_11301,N_11220,N_11011);
and U11302 (N_11302,N_11223,N_11014);
or U11303 (N_11303,N_11099,N_11034);
and U11304 (N_11304,N_11111,N_11142);
xor U11305 (N_11305,N_11058,N_11038);
nand U11306 (N_11306,N_11079,N_11066);
xnor U11307 (N_11307,N_11084,N_11196);
and U11308 (N_11308,N_11174,N_11230);
nand U11309 (N_11309,N_11041,N_11199);
or U11310 (N_11310,N_11241,N_11087);
nor U11311 (N_11311,N_11069,N_11035);
xnor U11312 (N_11312,N_11204,N_11242);
nor U11313 (N_11313,N_11018,N_11024);
and U11314 (N_11314,N_11195,N_11023);
xnor U11315 (N_11315,N_11192,N_11052);
nand U11316 (N_11316,N_11000,N_11249);
xor U11317 (N_11317,N_11044,N_11171);
or U11318 (N_11318,N_11211,N_11213);
nand U11319 (N_11319,N_11097,N_11008);
or U11320 (N_11320,N_11098,N_11217);
nor U11321 (N_11321,N_11110,N_11067);
or U11322 (N_11322,N_11105,N_11128);
or U11323 (N_11323,N_11193,N_11173);
xnor U11324 (N_11324,N_11124,N_11071);
nor U11325 (N_11325,N_11135,N_11010);
xnor U11326 (N_11326,N_11072,N_11061);
or U11327 (N_11327,N_11232,N_11118);
and U11328 (N_11328,N_11022,N_11170);
or U11329 (N_11329,N_11117,N_11054);
or U11330 (N_11330,N_11207,N_11043);
nor U11331 (N_11331,N_11228,N_11191);
xor U11332 (N_11332,N_11186,N_11039);
nor U11333 (N_11333,N_11235,N_11019);
xor U11334 (N_11334,N_11221,N_11094);
or U11335 (N_11335,N_11009,N_11016);
or U11336 (N_11336,N_11243,N_11074);
nand U11337 (N_11337,N_11051,N_11076);
nand U11338 (N_11338,N_11127,N_11167);
and U11339 (N_11339,N_11153,N_11201);
nor U11340 (N_11340,N_11059,N_11088);
xor U11341 (N_11341,N_11234,N_11017);
or U11342 (N_11342,N_11233,N_11103);
and U11343 (N_11343,N_11029,N_11007);
xor U11344 (N_11344,N_11181,N_11206);
nor U11345 (N_11345,N_11164,N_11147);
or U11346 (N_11346,N_11143,N_11216);
or U11347 (N_11347,N_11145,N_11100);
or U11348 (N_11348,N_11120,N_11246);
nand U11349 (N_11349,N_11205,N_11028);
xor U11350 (N_11350,N_11165,N_11154);
nor U11351 (N_11351,N_11157,N_11091);
or U11352 (N_11352,N_11021,N_11172);
nor U11353 (N_11353,N_11140,N_11133);
nand U11354 (N_11354,N_11150,N_11136);
nand U11355 (N_11355,N_11162,N_11108);
and U11356 (N_11356,N_11063,N_11056);
and U11357 (N_11357,N_11159,N_11144);
and U11358 (N_11358,N_11125,N_11212);
nand U11359 (N_11359,N_11176,N_11081);
or U11360 (N_11360,N_11210,N_11148);
or U11361 (N_11361,N_11115,N_11025);
and U11362 (N_11362,N_11049,N_11183);
nor U11363 (N_11363,N_11200,N_11040);
nor U11364 (N_11364,N_11048,N_11237);
nand U11365 (N_11365,N_11006,N_11037);
xor U11366 (N_11366,N_11045,N_11078);
xor U11367 (N_11367,N_11042,N_11004);
xnor U11368 (N_11368,N_11149,N_11177);
and U11369 (N_11369,N_11190,N_11102);
and U11370 (N_11370,N_11013,N_11244);
nand U11371 (N_11371,N_11236,N_11168);
and U11372 (N_11372,N_11175,N_11238);
xnor U11373 (N_11373,N_11163,N_11114);
and U11374 (N_11374,N_11126,N_11077);
nor U11375 (N_11375,N_11001,N_11134);
xor U11376 (N_11376,N_11058,N_11188);
nor U11377 (N_11377,N_11068,N_11177);
and U11378 (N_11378,N_11055,N_11198);
nor U11379 (N_11379,N_11047,N_11009);
nor U11380 (N_11380,N_11065,N_11155);
xnor U11381 (N_11381,N_11203,N_11016);
xor U11382 (N_11382,N_11002,N_11019);
xnor U11383 (N_11383,N_11140,N_11167);
nor U11384 (N_11384,N_11088,N_11194);
or U11385 (N_11385,N_11073,N_11199);
nand U11386 (N_11386,N_11195,N_11010);
and U11387 (N_11387,N_11000,N_11201);
nor U11388 (N_11388,N_11027,N_11215);
or U11389 (N_11389,N_11233,N_11069);
or U11390 (N_11390,N_11025,N_11169);
and U11391 (N_11391,N_11021,N_11148);
xor U11392 (N_11392,N_11126,N_11104);
nor U11393 (N_11393,N_11187,N_11171);
nand U11394 (N_11394,N_11052,N_11197);
nor U11395 (N_11395,N_11218,N_11108);
or U11396 (N_11396,N_11098,N_11066);
and U11397 (N_11397,N_11116,N_11152);
xor U11398 (N_11398,N_11036,N_11144);
and U11399 (N_11399,N_11195,N_11104);
nand U11400 (N_11400,N_11104,N_11158);
or U11401 (N_11401,N_11183,N_11203);
or U11402 (N_11402,N_11182,N_11037);
or U11403 (N_11403,N_11248,N_11153);
nor U11404 (N_11404,N_11037,N_11062);
xor U11405 (N_11405,N_11027,N_11103);
xnor U11406 (N_11406,N_11173,N_11107);
nand U11407 (N_11407,N_11153,N_11212);
xor U11408 (N_11408,N_11040,N_11186);
nand U11409 (N_11409,N_11168,N_11084);
and U11410 (N_11410,N_11013,N_11185);
and U11411 (N_11411,N_11014,N_11158);
and U11412 (N_11412,N_11014,N_11049);
and U11413 (N_11413,N_11104,N_11044);
nand U11414 (N_11414,N_11225,N_11119);
xor U11415 (N_11415,N_11095,N_11091);
nand U11416 (N_11416,N_11130,N_11063);
nor U11417 (N_11417,N_11080,N_11220);
xor U11418 (N_11418,N_11174,N_11156);
and U11419 (N_11419,N_11053,N_11154);
and U11420 (N_11420,N_11030,N_11230);
nor U11421 (N_11421,N_11164,N_11191);
nor U11422 (N_11422,N_11103,N_11113);
nand U11423 (N_11423,N_11213,N_11215);
nor U11424 (N_11424,N_11121,N_11097);
xor U11425 (N_11425,N_11067,N_11116);
xor U11426 (N_11426,N_11212,N_11163);
and U11427 (N_11427,N_11124,N_11008);
or U11428 (N_11428,N_11111,N_11222);
xnor U11429 (N_11429,N_11054,N_11185);
nand U11430 (N_11430,N_11148,N_11104);
nand U11431 (N_11431,N_11193,N_11059);
xor U11432 (N_11432,N_11019,N_11132);
or U11433 (N_11433,N_11133,N_11126);
nor U11434 (N_11434,N_11012,N_11163);
xnor U11435 (N_11435,N_11090,N_11028);
xnor U11436 (N_11436,N_11234,N_11071);
xnor U11437 (N_11437,N_11015,N_11064);
nand U11438 (N_11438,N_11219,N_11198);
xnor U11439 (N_11439,N_11065,N_11189);
or U11440 (N_11440,N_11242,N_11245);
and U11441 (N_11441,N_11033,N_11028);
and U11442 (N_11442,N_11108,N_11014);
or U11443 (N_11443,N_11161,N_11115);
and U11444 (N_11444,N_11087,N_11236);
and U11445 (N_11445,N_11212,N_11199);
and U11446 (N_11446,N_11183,N_11135);
and U11447 (N_11447,N_11119,N_11200);
or U11448 (N_11448,N_11065,N_11114);
and U11449 (N_11449,N_11176,N_11071);
nor U11450 (N_11450,N_11182,N_11004);
nor U11451 (N_11451,N_11093,N_11193);
or U11452 (N_11452,N_11002,N_11111);
nand U11453 (N_11453,N_11191,N_11231);
or U11454 (N_11454,N_11181,N_11187);
and U11455 (N_11455,N_11054,N_11038);
xnor U11456 (N_11456,N_11097,N_11141);
or U11457 (N_11457,N_11163,N_11216);
nor U11458 (N_11458,N_11015,N_11120);
or U11459 (N_11459,N_11129,N_11224);
nand U11460 (N_11460,N_11148,N_11036);
and U11461 (N_11461,N_11174,N_11107);
nor U11462 (N_11462,N_11236,N_11173);
and U11463 (N_11463,N_11142,N_11200);
or U11464 (N_11464,N_11163,N_11037);
and U11465 (N_11465,N_11186,N_11219);
nand U11466 (N_11466,N_11225,N_11105);
nor U11467 (N_11467,N_11120,N_11224);
nand U11468 (N_11468,N_11149,N_11013);
nor U11469 (N_11469,N_11143,N_11174);
and U11470 (N_11470,N_11150,N_11245);
nor U11471 (N_11471,N_11088,N_11070);
or U11472 (N_11472,N_11152,N_11127);
xor U11473 (N_11473,N_11080,N_11108);
or U11474 (N_11474,N_11196,N_11107);
nand U11475 (N_11475,N_11032,N_11027);
nor U11476 (N_11476,N_11004,N_11209);
or U11477 (N_11477,N_11124,N_11028);
nand U11478 (N_11478,N_11025,N_11209);
or U11479 (N_11479,N_11153,N_11069);
nand U11480 (N_11480,N_11135,N_11112);
and U11481 (N_11481,N_11140,N_11150);
xnor U11482 (N_11482,N_11176,N_11004);
nor U11483 (N_11483,N_11103,N_11063);
nor U11484 (N_11484,N_11028,N_11223);
or U11485 (N_11485,N_11086,N_11212);
xor U11486 (N_11486,N_11075,N_11243);
and U11487 (N_11487,N_11133,N_11004);
nor U11488 (N_11488,N_11235,N_11045);
or U11489 (N_11489,N_11123,N_11055);
nand U11490 (N_11490,N_11165,N_11176);
nor U11491 (N_11491,N_11200,N_11113);
or U11492 (N_11492,N_11017,N_11159);
nor U11493 (N_11493,N_11073,N_11191);
or U11494 (N_11494,N_11176,N_11184);
and U11495 (N_11495,N_11110,N_11040);
nor U11496 (N_11496,N_11226,N_11218);
xnor U11497 (N_11497,N_11091,N_11066);
nand U11498 (N_11498,N_11035,N_11158);
xnor U11499 (N_11499,N_11241,N_11237);
nand U11500 (N_11500,N_11296,N_11307);
nand U11501 (N_11501,N_11291,N_11304);
or U11502 (N_11502,N_11358,N_11422);
or U11503 (N_11503,N_11395,N_11499);
and U11504 (N_11504,N_11365,N_11494);
or U11505 (N_11505,N_11392,N_11278);
nor U11506 (N_11506,N_11279,N_11355);
nor U11507 (N_11507,N_11418,N_11491);
xor U11508 (N_11508,N_11288,N_11300);
xor U11509 (N_11509,N_11469,N_11368);
xnor U11510 (N_11510,N_11330,N_11322);
xnor U11511 (N_11511,N_11261,N_11464);
nor U11512 (N_11512,N_11462,N_11460);
nand U11513 (N_11513,N_11301,N_11430);
nand U11514 (N_11514,N_11425,N_11305);
nor U11515 (N_11515,N_11447,N_11335);
nand U11516 (N_11516,N_11428,N_11394);
or U11517 (N_11517,N_11391,N_11281);
and U11518 (N_11518,N_11276,N_11269);
or U11519 (N_11519,N_11334,N_11496);
nand U11520 (N_11520,N_11381,N_11433);
and U11521 (N_11521,N_11492,N_11495);
and U11522 (N_11522,N_11407,N_11378);
or U11523 (N_11523,N_11316,N_11376);
nor U11524 (N_11524,N_11331,N_11252);
nor U11525 (N_11525,N_11478,N_11454);
or U11526 (N_11526,N_11293,N_11292);
nor U11527 (N_11527,N_11280,N_11324);
or U11528 (N_11528,N_11497,N_11317);
nand U11529 (N_11529,N_11493,N_11306);
or U11530 (N_11530,N_11277,N_11397);
or U11531 (N_11531,N_11406,N_11314);
nor U11532 (N_11532,N_11452,N_11318);
and U11533 (N_11533,N_11268,N_11339);
nor U11534 (N_11534,N_11337,N_11251);
nand U11535 (N_11535,N_11442,N_11253);
nor U11536 (N_11536,N_11383,N_11264);
or U11537 (N_11537,N_11362,N_11364);
or U11538 (N_11538,N_11284,N_11417);
xor U11539 (N_11539,N_11267,N_11434);
xor U11540 (N_11540,N_11479,N_11333);
nand U11541 (N_11541,N_11379,N_11256);
nand U11542 (N_11542,N_11321,N_11275);
nand U11543 (N_11543,N_11312,N_11467);
and U11544 (N_11544,N_11262,N_11257);
nor U11545 (N_11545,N_11265,N_11295);
or U11546 (N_11546,N_11471,N_11429);
xor U11547 (N_11547,N_11352,N_11308);
nor U11548 (N_11548,N_11328,N_11481);
nor U11549 (N_11549,N_11488,N_11375);
nor U11550 (N_11550,N_11413,N_11448);
nand U11551 (N_11551,N_11455,N_11270);
and U11552 (N_11552,N_11289,N_11332);
nand U11553 (N_11553,N_11426,N_11311);
or U11554 (N_11554,N_11282,N_11370);
or U11555 (N_11555,N_11389,N_11483);
and U11556 (N_11556,N_11439,N_11357);
nor U11557 (N_11557,N_11440,N_11273);
nand U11558 (N_11558,N_11287,N_11470);
and U11559 (N_11559,N_11393,N_11423);
or U11560 (N_11560,N_11411,N_11450);
or U11561 (N_11561,N_11346,N_11345);
nand U11562 (N_11562,N_11310,N_11309);
nand U11563 (N_11563,N_11298,N_11427);
nand U11564 (N_11564,N_11415,N_11286);
nand U11565 (N_11565,N_11336,N_11482);
nor U11566 (N_11566,N_11441,N_11432);
nand U11567 (N_11567,N_11353,N_11402);
xor U11568 (N_11568,N_11258,N_11473);
nand U11569 (N_11569,N_11315,N_11329);
xnor U11570 (N_11570,N_11377,N_11387);
xnor U11571 (N_11571,N_11272,N_11359);
xnor U11572 (N_11572,N_11484,N_11369);
and U11573 (N_11573,N_11366,N_11347);
and U11574 (N_11574,N_11323,N_11356);
nand U11575 (N_11575,N_11348,N_11461);
xor U11576 (N_11576,N_11476,N_11283);
and U11577 (N_11577,N_11319,N_11340);
xnor U11578 (N_11578,N_11285,N_11326);
nand U11579 (N_11579,N_11255,N_11403);
nor U11580 (N_11580,N_11463,N_11435);
or U11581 (N_11581,N_11421,N_11468);
and U11582 (N_11582,N_11374,N_11480);
nor U11583 (N_11583,N_11343,N_11416);
and U11584 (N_11584,N_11475,N_11487);
nor U11585 (N_11585,N_11390,N_11371);
nor U11586 (N_11586,N_11490,N_11438);
nor U11587 (N_11587,N_11354,N_11360);
nor U11588 (N_11588,N_11456,N_11266);
xnor U11589 (N_11589,N_11299,N_11342);
nand U11590 (N_11590,N_11250,N_11414);
or U11591 (N_11591,N_11404,N_11458);
or U11592 (N_11592,N_11271,N_11408);
nor U11593 (N_11593,N_11373,N_11274);
xor U11594 (N_11594,N_11401,N_11325);
and U11595 (N_11595,N_11486,N_11382);
xnor U11596 (N_11596,N_11449,N_11294);
nand U11597 (N_11597,N_11412,N_11443);
or U11598 (N_11598,N_11320,N_11341);
xnor U11599 (N_11599,N_11372,N_11344);
nor U11600 (N_11600,N_11431,N_11446);
or U11601 (N_11601,N_11457,N_11489);
and U11602 (N_11602,N_11405,N_11297);
nand U11603 (N_11603,N_11465,N_11444);
or U11604 (N_11604,N_11327,N_11396);
or U11605 (N_11605,N_11367,N_11349);
or U11606 (N_11606,N_11388,N_11386);
xnor U11607 (N_11607,N_11399,N_11385);
xor U11608 (N_11608,N_11453,N_11419);
and U11609 (N_11609,N_11459,N_11472);
or U11610 (N_11610,N_11398,N_11498);
nor U11611 (N_11611,N_11485,N_11380);
or U11612 (N_11612,N_11303,N_11420);
or U11613 (N_11613,N_11437,N_11338);
nor U11614 (N_11614,N_11477,N_11410);
or U11615 (N_11615,N_11351,N_11466);
or U11616 (N_11616,N_11254,N_11409);
and U11617 (N_11617,N_11350,N_11445);
and U11618 (N_11618,N_11302,N_11290);
nand U11619 (N_11619,N_11260,N_11361);
and U11620 (N_11620,N_11259,N_11424);
nand U11621 (N_11621,N_11451,N_11363);
xnor U11622 (N_11622,N_11474,N_11436);
and U11623 (N_11623,N_11400,N_11263);
and U11624 (N_11624,N_11384,N_11313);
nand U11625 (N_11625,N_11285,N_11408);
or U11626 (N_11626,N_11412,N_11310);
or U11627 (N_11627,N_11336,N_11294);
xor U11628 (N_11628,N_11499,N_11314);
xnor U11629 (N_11629,N_11294,N_11306);
or U11630 (N_11630,N_11377,N_11459);
nor U11631 (N_11631,N_11446,N_11382);
xor U11632 (N_11632,N_11250,N_11417);
and U11633 (N_11633,N_11493,N_11362);
and U11634 (N_11634,N_11464,N_11494);
nor U11635 (N_11635,N_11472,N_11429);
xor U11636 (N_11636,N_11265,N_11292);
nor U11637 (N_11637,N_11327,N_11451);
or U11638 (N_11638,N_11420,N_11262);
and U11639 (N_11639,N_11365,N_11374);
nor U11640 (N_11640,N_11498,N_11437);
xnor U11641 (N_11641,N_11422,N_11466);
or U11642 (N_11642,N_11470,N_11400);
nand U11643 (N_11643,N_11454,N_11309);
xnor U11644 (N_11644,N_11427,N_11293);
xnor U11645 (N_11645,N_11279,N_11490);
nand U11646 (N_11646,N_11299,N_11384);
nand U11647 (N_11647,N_11410,N_11435);
nor U11648 (N_11648,N_11274,N_11421);
nand U11649 (N_11649,N_11402,N_11429);
or U11650 (N_11650,N_11452,N_11368);
or U11651 (N_11651,N_11403,N_11416);
xor U11652 (N_11652,N_11353,N_11280);
xnor U11653 (N_11653,N_11495,N_11432);
xnor U11654 (N_11654,N_11260,N_11327);
nor U11655 (N_11655,N_11420,N_11488);
and U11656 (N_11656,N_11365,N_11320);
nor U11657 (N_11657,N_11485,N_11355);
or U11658 (N_11658,N_11461,N_11408);
nor U11659 (N_11659,N_11474,N_11308);
nor U11660 (N_11660,N_11331,N_11352);
and U11661 (N_11661,N_11269,N_11450);
xor U11662 (N_11662,N_11344,N_11342);
or U11663 (N_11663,N_11468,N_11472);
xor U11664 (N_11664,N_11295,N_11349);
or U11665 (N_11665,N_11333,N_11323);
nand U11666 (N_11666,N_11313,N_11414);
or U11667 (N_11667,N_11285,N_11268);
nor U11668 (N_11668,N_11463,N_11310);
or U11669 (N_11669,N_11443,N_11418);
and U11670 (N_11670,N_11255,N_11481);
nand U11671 (N_11671,N_11326,N_11496);
nor U11672 (N_11672,N_11280,N_11447);
xor U11673 (N_11673,N_11289,N_11378);
nor U11674 (N_11674,N_11250,N_11498);
or U11675 (N_11675,N_11321,N_11259);
and U11676 (N_11676,N_11472,N_11381);
or U11677 (N_11677,N_11373,N_11366);
nor U11678 (N_11678,N_11269,N_11474);
and U11679 (N_11679,N_11461,N_11310);
and U11680 (N_11680,N_11275,N_11395);
and U11681 (N_11681,N_11319,N_11349);
nor U11682 (N_11682,N_11446,N_11282);
xnor U11683 (N_11683,N_11487,N_11351);
or U11684 (N_11684,N_11330,N_11299);
nand U11685 (N_11685,N_11328,N_11366);
or U11686 (N_11686,N_11455,N_11411);
and U11687 (N_11687,N_11360,N_11381);
nand U11688 (N_11688,N_11358,N_11311);
xnor U11689 (N_11689,N_11261,N_11449);
or U11690 (N_11690,N_11273,N_11343);
xnor U11691 (N_11691,N_11346,N_11302);
or U11692 (N_11692,N_11454,N_11386);
nor U11693 (N_11693,N_11482,N_11276);
or U11694 (N_11694,N_11449,N_11435);
and U11695 (N_11695,N_11271,N_11498);
nand U11696 (N_11696,N_11378,N_11314);
nor U11697 (N_11697,N_11369,N_11314);
xor U11698 (N_11698,N_11454,N_11379);
xnor U11699 (N_11699,N_11469,N_11384);
nand U11700 (N_11700,N_11368,N_11402);
nand U11701 (N_11701,N_11469,N_11340);
and U11702 (N_11702,N_11349,N_11409);
xor U11703 (N_11703,N_11278,N_11268);
or U11704 (N_11704,N_11316,N_11300);
nor U11705 (N_11705,N_11420,N_11474);
nor U11706 (N_11706,N_11484,N_11403);
nor U11707 (N_11707,N_11296,N_11370);
xnor U11708 (N_11708,N_11285,N_11382);
nor U11709 (N_11709,N_11432,N_11354);
nor U11710 (N_11710,N_11451,N_11292);
xnor U11711 (N_11711,N_11474,N_11276);
nand U11712 (N_11712,N_11442,N_11353);
nor U11713 (N_11713,N_11444,N_11294);
nor U11714 (N_11714,N_11452,N_11466);
nor U11715 (N_11715,N_11419,N_11341);
nand U11716 (N_11716,N_11469,N_11289);
and U11717 (N_11717,N_11317,N_11258);
or U11718 (N_11718,N_11257,N_11470);
nor U11719 (N_11719,N_11480,N_11353);
or U11720 (N_11720,N_11455,N_11313);
xnor U11721 (N_11721,N_11394,N_11278);
xnor U11722 (N_11722,N_11406,N_11309);
and U11723 (N_11723,N_11301,N_11279);
xor U11724 (N_11724,N_11400,N_11370);
nor U11725 (N_11725,N_11318,N_11437);
nor U11726 (N_11726,N_11296,N_11376);
xor U11727 (N_11727,N_11493,N_11483);
nand U11728 (N_11728,N_11365,N_11385);
or U11729 (N_11729,N_11448,N_11347);
nand U11730 (N_11730,N_11401,N_11382);
nand U11731 (N_11731,N_11349,N_11452);
nor U11732 (N_11732,N_11257,N_11394);
or U11733 (N_11733,N_11466,N_11378);
xnor U11734 (N_11734,N_11407,N_11318);
nor U11735 (N_11735,N_11328,N_11475);
xnor U11736 (N_11736,N_11394,N_11308);
nand U11737 (N_11737,N_11352,N_11410);
xnor U11738 (N_11738,N_11403,N_11317);
nand U11739 (N_11739,N_11314,N_11432);
xor U11740 (N_11740,N_11361,N_11434);
and U11741 (N_11741,N_11414,N_11445);
and U11742 (N_11742,N_11378,N_11339);
nand U11743 (N_11743,N_11380,N_11335);
or U11744 (N_11744,N_11339,N_11452);
nand U11745 (N_11745,N_11411,N_11345);
nor U11746 (N_11746,N_11258,N_11494);
nor U11747 (N_11747,N_11486,N_11404);
nor U11748 (N_11748,N_11408,N_11400);
nand U11749 (N_11749,N_11304,N_11303);
or U11750 (N_11750,N_11593,N_11539);
xor U11751 (N_11751,N_11502,N_11611);
nor U11752 (N_11752,N_11607,N_11556);
nor U11753 (N_11753,N_11632,N_11585);
and U11754 (N_11754,N_11722,N_11622);
xnor U11755 (N_11755,N_11626,N_11586);
and U11756 (N_11756,N_11725,N_11583);
or U11757 (N_11757,N_11741,N_11679);
nor U11758 (N_11758,N_11678,N_11548);
nor U11759 (N_11759,N_11706,N_11653);
nand U11760 (N_11760,N_11567,N_11691);
xnor U11761 (N_11761,N_11528,N_11541);
nor U11762 (N_11762,N_11547,N_11553);
or U11763 (N_11763,N_11596,N_11545);
or U11764 (N_11764,N_11538,N_11625);
nand U11765 (N_11765,N_11578,N_11619);
xor U11766 (N_11766,N_11521,N_11638);
or U11767 (N_11767,N_11623,N_11637);
xor U11768 (N_11768,N_11517,N_11514);
nand U11769 (N_11769,N_11627,N_11674);
or U11770 (N_11770,N_11672,N_11647);
xnor U11771 (N_11771,N_11654,N_11579);
xnor U11772 (N_11772,N_11608,N_11577);
nor U11773 (N_11773,N_11644,N_11661);
nor U11774 (N_11774,N_11718,N_11742);
and U11775 (N_11775,N_11512,N_11649);
nor U11776 (N_11776,N_11666,N_11564);
and U11777 (N_11777,N_11501,N_11677);
and U11778 (N_11778,N_11519,N_11524);
or U11779 (N_11779,N_11575,N_11552);
and U11780 (N_11780,N_11656,N_11709);
or U11781 (N_11781,N_11581,N_11689);
or U11782 (N_11782,N_11712,N_11588);
or U11783 (N_11783,N_11702,N_11744);
nand U11784 (N_11784,N_11582,N_11614);
nor U11785 (N_11785,N_11694,N_11682);
or U11786 (N_11786,N_11565,N_11738);
nand U11787 (N_11787,N_11642,N_11600);
xor U11788 (N_11788,N_11518,N_11597);
xnor U11789 (N_11789,N_11748,N_11745);
xnor U11790 (N_11790,N_11606,N_11536);
and U11791 (N_11791,N_11729,N_11735);
nand U11792 (N_11792,N_11639,N_11715);
nand U11793 (N_11793,N_11568,N_11673);
xor U11794 (N_11794,N_11646,N_11605);
nor U11795 (N_11795,N_11714,N_11676);
nand U11796 (N_11796,N_11665,N_11736);
xor U11797 (N_11797,N_11680,N_11713);
or U11798 (N_11798,N_11511,N_11520);
nor U11799 (N_11799,N_11658,N_11563);
xnor U11800 (N_11800,N_11739,N_11645);
xor U11801 (N_11801,N_11560,N_11590);
or U11802 (N_11802,N_11719,N_11531);
and U11803 (N_11803,N_11584,N_11724);
xor U11804 (N_11804,N_11610,N_11526);
or U11805 (N_11805,N_11570,N_11576);
or U11806 (N_11806,N_11613,N_11746);
and U11807 (N_11807,N_11500,N_11508);
or U11808 (N_11808,N_11651,N_11657);
and U11809 (N_11809,N_11617,N_11603);
xnor U11810 (N_11810,N_11717,N_11635);
nor U11811 (N_11811,N_11628,N_11703);
nand U11812 (N_11812,N_11532,N_11660);
xor U11813 (N_11813,N_11509,N_11542);
nor U11814 (N_11814,N_11507,N_11684);
or U11815 (N_11815,N_11624,N_11631);
nand U11816 (N_11816,N_11599,N_11515);
or U11817 (N_11817,N_11700,N_11602);
nand U11818 (N_11818,N_11527,N_11523);
nor U11819 (N_11819,N_11634,N_11731);
or U11820 (N_11820,N_11609,N_11723);
nand U11821 (N_11821,N_11696,N_11534);
or U11822 (N_11822,N_11506,N_11683);
xnor U11823 (N_11823,N_11557,N_11566);
nor U11824 (N_11824,N_11640,N_11716);
or U11825 (N_11825,N_11690,N_11551);
xnor U11826 (N_11826,N_11734,N_11733);
nand U11827 (N_11827,N_11572,N_11643);
nand U11828 (N_11828,N_11668,N_11699);
xor U11829 (N_11829,N_11562,N_11503);
xor U11830 (N_11830,N_11747,N_11561);
and U11831 (N_11831,N_11670,N_11681);
nand U11832 (N_11832,N_11720,N_11697);
nand U11833 (N_11833,N_11663,N_11510);
nor U11834 (N_11834,N_11554,N_11569);
or U11835 (N_11835,N_11727,N_11749);
and U11836 (N_11836,N_11662,N_11701);
nand U11837 (N_11837,N_11705,N_11505);
nand U11838 (N_11838,N_11549,N_11522);
xnor U11839 (N_11839,N_11740,N_11621);
nor U11840 (N_11840,N_11648,N_11629);
xnor U11841 (N_11841,N_11571,N_11544);
nand U11842 (N_11842,N_11559,N_11550);
nor U11843 (N_11843,N_11595,N_11667);
xor U11844 (N_11844,N_11555,N_11636);
xnor U11845 (N_11845,N_11687,N_11693);
xor U11846 (N_11846,N_11671,N_11732);
nor U11847 (N_11847,N_11601,N_11591);
and U11848 (N_11848,N_11598,N_11574);
and U11849 (N_11849,N_11686,N_11688);
and U11850 (N_11850,N_11558,N_11533);
or U11851 (N_11851,N_11540,N_11685);
or U11852 (N_11852,N_11708,N_11707);
and U11853 (N_11853,N_11504,N_11710);
and U11854 (N_11854,N_11612,N_11633);
or U11855 (N_11855,N_11513,N_11618);
and U11856 (N_11856,N_11737,N_11616);
nand U11857 (N_11857,N_11704,N_11730);
nand U11858 (N_11858,N_11652,N_11641);
and U11859 (N_11859,N_11692,N_11726);
nand U11860 (N_11860,N_11620,N_11711);
xor U11861 (N_11861,N_11543,N_11615);
xor U11862 (N_11862,N_11516,N_11580);
xnor U11863 (N_11863,N_11669,N_11537);
and U11864 (N_11864,N_11530,N_11698);
or U11865 (N_11865,N_11728,N_11655);
and U11866 (N_11866,N_11525,N_11650);
nand U11867 (N_11867,N_11743,N_11529);
or U11868 (N_11868,N_11594,N_11573);
or U11869 (N_11869,N_11630,N_11589);
nand U11870 (N_11870,N_11535,N_11675);
or U11871 (N_11871,N_11592,N_11546);
nor U11872 (N_11872,N_11721,N_11604);
or U11873 (N_11873,N_11664,N_11659);
and U11874 (N_11874,N_11695,N_11587);
and U11875 (N_11875,N_11639,N_11610);
and U11876 (N_11876,N_11635,N_11657);
and U11877 (N_11877,N_11589,N_11609);
nand U11878 (N_11878,N_11745,N_11621);
and U11879 (N_11879,N_11655,N_11550);
and U11880 (N_11880,N_11518,N_11512);
and U11881 (N_11881,N_11570,N_11732);
nand U11882 (N_11882,N_11629,N_11716);
or U11883 (N_11883,N_11642,N_11588);
nand U11884 (N_11884,N_11554,N_11583);
xnor U11885 (N_11885,N_11552,N_11546);
nor U11886 (N_11886,N_11615,N_11504);
or U11887 (N_11887,N_11529,N_11537);
nand U11888 (N_11888,N_11555,N_11519);
nor U11889 (N_11889,N_11592,N_11741);
nor U11890 (N_11890,N_11508,N_11639);
nor U11891 (N_11891,N_11608,N_11545);
nand U11892 (N_11892,N_11524,N_11560);
or U11893 (N_11893,N_11656,N_11743);
or U11894 (N_11894,N_11625,N_11606);
nand U11895 (N_11895,N_11740,N_11669);
xor U11896 (N_11896,N_11667,N_11531);
and U11897 (N_11897,N_11689,N_11613);
nand U11898 (N_11898,N_11571,N_11711);
nor U11899 (N_11899,N_11612,N_11519);
nand U11900 (N_11900,N_11643,N_11652);
xor U11901 (N_11901,N_11624,N_11542);
or U11902 (N_11902,N_11501,N_11670);
nor U11903 (N_11903,N_11574,N_11720);
nand U11904 (N_11904,N_11549,N_11519);
nand U11905 (N_11905,N_11605,N_11723);
xor U11906 (N_11906,N_11582,N_11723);
nor U11907 (N_11907,N_11574,N_11722);
nand U11908 (N_11908,N_11529,N_11623);
nand U11909 (N_11909,N_11517,N_11598);
nand U11910 (N_11910,N_11640,N_11611);
or U11911 (N_11911,N_11604,N_11526);
nand U11912 (N_11912,N_11739,N_11729);
xor U11913 (N_11913,N_11615,N_11735);
or U11914 (N_11914,N_11587,N_11545);
or U11915 (N_11915,N_11590,N_11576);
nor U11916 (N_11916,N_11700,N_11665);
xnor U11917 (N_11917,N_11701,N_11535);
nor U11918 (N_11918,N_11649,N_11618);
xor U11919 (N_11919,N_11560,N_11612);
and U11920 (N_11920,N_11651,N_11573);
and U11921 (N_11921,N_11629,N_11719);
nand U11922 (N_11922,N_11677,N_11620);
and U11923 (N_11923,N_11702,N_11578);
nand U11924 (N_11924,N_11532,N_11687);
nand U11925 (N_11925,N_11640,N_11583);
nand U11926 (N_11926,N_11617,N_11570);
nor U11927 (N_11927,N_11569,N_11575);
or U11928 (N_11928,N_11566,N_11657);
xnor U11929 (N_11929,N_11559,N_11708);
or U11930 (N_11930,N_11581,N_11532);
nand U11931 (N_11931,N_11613,N_11728);
nor U11932 (N_11932,N_11623,N_11739);
nor U11933 (N_11933,N_11652,N_11735);
and U11934 (N_11934,N_11639,N_11501);
or U11935 (N_11935,N_11651,N_11712);
nor U11936 (N_11936,N_11544,N_11518);
xnor U11937 (N_11937,N_11636,N_11651);
or U11938 (N_11938,N_11688,N_11624);
xnor U11939 (N_11939,N_11627,N_11661);
nand U11940 (N_11940,N_11563,N_11727);
xor U11941 (N_11941,N_11617,N_11518);
nor U11942 (N_11942,N_11633,N_11701);
and U11943 (N_11943,N_11684,N_11679);
or U11944 (N_11944,N_11587,N_11732);
xor U11945 (N_11945,N_11712,N_11611);
or U11946 (N_11946,N_11719,N_11677);
and U11947 (N_11947,N_11532,N_11673);
xor U11948 (N_11948,N_11628,N_11539);
and U11949 (N_11949,N_11655,N_11697);
nor U11950 (N_11950,N_11661,N_11527);
xor U11951 (N_11951,N_11689,N_11621);
xnor U11952 (N_11952,N_11553,N_11718);
xnor U11953 (N_11953,N_11699,N_11541);
nand U11954 (N_11954,N_11664,N_11592);
xnor U11955 (N_11955,N_11501,N_11547);
nand U11956 (N_11956,N_11558,N_11701);
or U11957 (N_11957,N_11556,N_11727);
nand U11958 (N_11958,N_11712,N_11638);
nand U11959 (N_11959,N_11587,N_11592);
and U11960 (N_11960,N_11567,N_11719);
nand U11961 (N_11961,N_11551,N_11563);
and U11962 (N_11962,N_11697,N_11547);
or U11963 (N_11963,N_11709,N_11710);
or U11964 (N_11964,N_11711,N_11707);
and U11965 (N_11965,N_11532,N_11500);
nor U11966 (N_11966,N_11570,N_11698);
nand U11967 (N_11967,N_11552,N_11557);
and U11968 (N_11968,N_11691,N_11655);
nand U11969 (N_11969,N_11566,N_11588);
xnor U11970 (N_11970,N_11562,N_11645);
nand U11971 (N_11971,N_11734,N_11619);
xnor U11972 (N_11972,N_11716,N_11524);
nor U11973 (N_11973,N_11664,N_11641);
nor U11974 (N_11974,N_11707,N_11606);
nand U11975 (N_11975,N_11695,N_11595);
and U11976 (N_11976,N_11599,N_11615);
nand U11977 (N_11977,N_11518,N_11527);
and U11978 (N_11978,N_11577,N_11658);
nor U11979 (N_11979,N_11718,N_11645);
xnor U11980 (N_11980,N_11632,N_11572);
and U11981 (N_11981,N_11664,N_11607);
or U11982 (N_11982,N_11566,N_11704);
nor U11983 (N_11983,N_11575,N_11518);
or U11984 (N_11984,N_11585,N_11507);
nand U11985 (N_11985,N_11603,N_11503);
xnor U11986 (N_11986,N_11729,N_11620);
xor U11987 (N_11987,N_11522,N_11737);
nor U11988 (N_11988,N_11714,N_11642);
and U11989 (N_11989,N_11607,N_11577);
nand U11990 (N_11990,N_11541,N_11644);
or U11991 (N_11991,N_11668,N_11691);
nor U11992 (N_11992,N_11704,N_11699);
or U11993 (N_11993,N_11573,N_11730);
xor U11994 (N_11994,N_11646,N_11714);
nor U11995 (N_11995,N_11669,N_11569);
xnor U11996 (N_11996,N_11697,N_11702);
nand U11997 (N_11997,N_11626,N_11538);
xor U11998 (N_11998,N_11715,N_11713);
xnor U11999 (N_11999,N_11531,N_11633);
nor U12000 (N_12000,N_11751,N_11854);
and U12001 (N_12001,N_11974,N_11859);
or U12002 (N_12002,N_11798,N_11965);
nor U12003 (N_12003,N_11954,N_11957);
xnor U12004 (N_12004,N_11875,N_11899);
and U12005 (N_12005,N_11858,N_11977);
nor U12006 (N_12006,N_11786,N_11849);
xor U12007 (N_12007,N_11860,N_11955);
or U12008 (N_12008,N_11837,N_11753);
or U12009 (N_12009,N_11873,N_11807);
xor U12010 (N_12010,N_11769,N_11795);
nor U12011 (N_12011,N_11821,N_11937);
or U12012 (N_12012,N_11862,N_11797);
nand U12013 (N_12013,N_11861,N_11811);
nand U12014 (N_12014,N_11764,N_11757);
xnor U12015 (N_12015,N_11758,N_11902);
nor U12016 (N_12016,N_11922,N_11832);
nand U12017 (N_12017,N_11770,N_11936);
and U12018 (N_12018,N_11956,N_11999);
or U12019 (N_12019,N_11782,N_11890);
nand U12020 (N_12020,N_11962,N_11935);
xor U12021 (N_12021,N_11793,N_11768);
xnor U12022 (N_12022,N_11947,N_11976);
and U12023 (N_12023,N_11896,N_11830);
nand U12024 (N_12024,N_11750,N_11978);
or U12025 (N_12025,N_11819,N_11825);
nor U12026 (N_12026,N_11848,N_11929);
xor U12027 (N_12027,N_11765,N_11767);
xnor U12028 (N_12028,N_11771,N_11833);
and U12029 (N_12029,N_11993,N_11763);
nor U12030 (N_12030,N_11949,N_11989);
nand U12031 (N_12031,N_11824,N_11778);
xnor U12032 (N_12032,N_11943,N_11953);
or U12033 (N_12033,N_11790,N_11996);
nand U12034 (N_12034,N_11970,N_11844);
nand U12035 (N_12035,N_11988,N_11952);
nor U12036 (N_12036,N_11879,N_11923);
xnor U12037 (N_12037,N_11846,N_11963);
or U12038 (N_12038,N_11818,N_11853);
nor U12039 (N_12039,N_11912,N_11838);
xor U12040 (N_12040,N_11983,N_11900);
xnor U12041 (N_12041,N_11813,N_11759);
xnor U12042 (N_12042,N_11775,N_11968);
xnor U12043 (N_12043,N_11967,N_11752);
nand U12044 (N_12044,N_11754,N_11883);
nor U12045 (N_12045,N_11841,N_11831);
and U12046 (N_12046,N_11945,N_11780);
xor U12047 (N_12047,N_11939,N_11930);
nand U12048 (N_12048,N_11938,N_11920);
nand U12049 (N_12049,N_11834,N_11785);
xor U12050 (N_12050,N_11906,N_11823);
nor U12051 (N_12051,N_11919,N_11975);
and U12052 (N_12052,N_11864,N_11980);
nand U12053 (N_12053,N_11942,N_11924);
xor U12054 (N_12054,N_11842,N_11991);
or U12055 (N_12055,N_11966,N_11982);
or U12056 (N_12056,N_11760,N_11761);
xor U12057 (N_12057,N_11788,N_11792);
nand U12058 (N_12058,N_11884,N_11969);
or U12059 (N_12059,N_11845,N_11791);
and U12060 (N_12060,N_11866,N_11876);
xnor U12061 (N_12061,N_11971,N_11863);
nor U12062 (N_12062,N_11784,N_11928);
and U12063 (N_12063,N_11891,N_11997);
or U12064 (N_12064,N_11941,N_11893);
xor U12065 (N_12065,N_11892,N_11774);
or U12066 (N_12066,N_11762,N_11926);
nor U12067 (N_12067,N_11925,N_11918);
or U12068 (N_12068,N_11828,N_11856);
or U12069 (N_12069,N_11802,N_11933);
and U12070 (N_12070,N_11852,N_11872);
xor U12071 (N_12071,N_11855,N_11794);
nor U12072 (N_12072,N_11911,N_11783);
nor U12073 (N_12073,N_11914,N_11800);
xnor U12074 (N_12074,N_11755,N_11889);
nor U12075 (N_12075,N_11960,N_11973);
or U12076 (N_12076,N_11882,N_11885);
and U12077 (N_12077,N_11972,N_11979);
nor U12078 (N_12078,N_11817,N_11756);
xnor U12079 (N_12079,N_11836,N_11870);
nand U12080 (N_12080,N_11804,N_11895);
and U12081 (N_12081,N_11905,N_11984);
and U12082 (N_12082,N_11816,N_11809);
nand U12083 (N_12083,N_11874,N_11917);
nor U12084 (N_12084,N_11847,N_11829);
nand U12085 (N_12085,N_11995,N_11931);
xnor U12086 (N_12086,N_11808,N_11909);
and U12087 (N_12087,N_11867,N_11881);
and U12088 (N_12088,N_11773,N_11789);
xnor U12089 (N_12089,N_11986,N_11787);
or U12090 (N_12090,N_11887,N_11994);
and U12091 (N_12091,N_11903,N_11915);
xor U12092 (N_12092,N_11806,N_11958);
nand U12093 (N_12093,N_11921,N_11799);
nor U12094 (N_12094,N_11850,N_11990);
nand U12095 (N_12095,N_11897,N_11766);
nand U12096 (N_12096,N_11877,N_11946);
nand U12097 (N_12097,N_11835,N_11810);
and U12098 (N_12098,N_11964,N_11803);
xnor U12099 (N_12099,N_11948,N_11781);
nand U12100 (N_12100,N_11812,N_11839);
nand U12101 (N_12101,N_11908,N_11871);
and U12102 (N_12102,N_11772,N_11826);
xor U12103 (N_12103,N_11927,N_11776);
and U12104 (N_12104,N_11878,N_11998);
nor U12105 (N_12105,N_11907,N_11940);
xnor U12106 (N_12106,N_11985,N_11843);
and U12107 (N_12107,N_11910,N_11894);
nand U12108 (N_12108,N_11801,N_11951);
nand U12109 (N_12109,N_11779,N_11886);
or U12110 (N_12110,N_11815,N_11857);
nor U12111 (N_12111,N_11944,N_11880);
nor U12112 (N_12112,N_11904,N_11827);
and U12113 (N_12113,N_11898,N_11961);
xor U12114 (N_12114,N_11888,N_11959);
and U12115 (N_12115,N_11869,N_11987);
and U12116 (N_12116,N_11913,N_11865);
and U12117 (N_12117,N_11840,N_11868);
and U12118 (N_12118,N_11814,N_11901);
nor U12119 (N_12119,N_11822,N_11796);
or U12120 (N_12120,N_11820,N_11934);
nand U12121 (N_12121,N_11992,N_11981);
nand U12122 (N_12122,N_11916,N_11805);
xnor U12123 (N_12123,N_11851,N_11950);
and U12124 (N_12124,N_11777,N_11932);
nor U12125 (N_12125,N_11760,N_11832);
nor U12126 (N_12126,N_11909,N_11968);
xnor U12127 (N_12127,N_11970,N_11830);
xnor U12128 (N_12128,N_11983,N_11870);
and U12129 (N_12129,N_11751,N_11978);
and U12130 (N_12130,N_11960,N_11889);
xor U12131 (N_12131,N_11992,N_11904);
nand U12132 (N_12132,N_11787,N_11770);
nand U12133 (N_12133,N_11842,N_11833);
nand U12134 (N_12134,N_11792,N_11924);
and U12135 (N_12135,N_11823,N_11760);
or U12136 (N_12136,N_11934,N_11754);
or U12137 (N_12137,N_11861,N_11953);
nand U12138 (N_12138,N_11874,N_11895);
or U12139 (N_12139,N_11889,N_11789);
nand U12140 (N_12140,N_11781,N_11986);
nand U12141 (N_12141,N_11775,N_11919);
xor U12142 (N_12142,N_11761,N_11914);
and U12143 (N_12143,N_11977,N_11854);
nor U12144 (N_12144,N_11845,N_11927);
or U12145 (N_12145,N_11960,N_11930);
xor U12146 (N_12146,N_11767,N_11993);
xnor U12147 (N_12147,N_11870,N_11919);
and U12148 (N_12148,N_11930,N_11800);
and U12149 (N_12149,N_11837,N_11872);
nor U12150 (N_12150,N_11951,N_11996);
or U12151 (N_12151,N_11986,N_11771);
or U12152 (N_12152,N_11946,N_11763);
and U12153 (N_12153,N_11781,N_11800);
or U12154 (N_12154,N_11943,N_11865);
nand U12155 (N_12155,N_11995,N_11813);
xnor U12156 (N_12156,N_11804,N_11809);
and U12157 (N_12157,N_11894,N_11770);
xor U12158 (N_12158,N_11992,N_11909);
nor U12159 (N_12159,N_11760,N_11923);
xor U12160 (N_12160,N_11911,N_11752);
nor U12161 (N_12161,N_11839,N_11757);
xor U12162 (N_12162,N_11946,N_11874);
nand U12163 (N_12163,N_11752,N_11925);
and U12164 (N_12164,N_11756,N_11856);
and U12165 (N_12165,N_11751,N_11828);
nor U12166 (N_12166,N_11896,N_11763);
or U12167 (N_12167,N_11985,N_11998);
nand U12168 (N_12168,N_11761,N_11843);
and U12169 (N_12169,N_11836,N_11764);
and U12170 (N_12170,N_11906,N_11947);
xor U12171 (N_12171,N_11915,N_11863);
and U12172 (N_12172,N_11822,N_11772);
xor U12173 (N_12173,N_11767,N_11797);
nand U12174 (N_12174,N_11852,N_11916);
nor U12175 (N_12175,N_11754,N_11867);
nor U12176 (N_12176,N_11753,N_11897);
nor U12177 (N_12177,N_11958,N_11775);
xor U12178 (N_12178,N_11792,N_11873);
and U12179 (N_12179,N_11818,N_11753);
nor U12180 (N_12180,N_11893,N_11828);
nand U12181 (N_12181,N_11952,N_11921);
and U12182 (N_12182,N_11999,N_11787);
or U12183 (N_12183,N_11955,N_11875);
nor U12184 (N_12184,N_11909,N_11790);
nand U12185 (N_12185,N_11959,N_11785);
or U12186 (N_12186,N_11980,N_11935);
nor U12187 (N_12187,N_11991,N_11944);
xnor U12188 (N_12188,N_11822,N_11992);
nor U12189 (N_12189,N_11903,N_11868);
nand U12190 (N_12190,N_11978,N_11971);
nand U12191 (N_12191,N_11908,N_11772);
and U12192 (N_12192,N_11838,N_11970);
nand U12193 (N_12193,N_11894,N_11962);
or U12194 (N_12194,N_11928,N_11822);
xnor U12195 (N_12195,N_11985,N_11847);
nand U12196 (N_12196,N_11993,N_11860);
or U12197 (N_12197,N_11925,N_11908);
and U12198 (N_12198,N_11865,N_11764);
nor U12199 (N_12199,N_11966,N_11772);
xor U12200 (N_12200,N_11983,N_11970);
nor U12201 (N_12201,N_11827,N_11927);
nand U12202 (N_12202,N_11939,N_11993);
nand U12203 (N_12203,N_11818,N_11939);
and U12204 (N_12204,N_11967,N_11780);
or U12205 (N_12205,N_11933,N_11973);
nand U12206 (N_12206,N_11914,N_11962);
nor U12207 (N_12207,N_11884,N_11771);
xnor U12208 (N_12208,N_11752,N_11870);
xnor U12209 (N_12209,N_11983,N_11971);
or U12210 (N_12210,N_11812,N_11813);
and U12211 (N_12211,N_11937,N_11822);
xnor U12212 (N_12212,N_11978,N_11795);
or U12213 (N_12213,N_11794,N_11919);
xor U12214 (N_12214,N_11947,N_11999);
nor U12215 (N_12215,N_11955,N_11973);
xor U12216 (N_12216,N_11794,N_11816);
nor U12217 (N_12217,N_11953,N_11850);
nand U12218 (N_12218,N_11958,N_11832);
xnor U12219 (N_12219,N_11946,N_11966);
nand U12220 (N_12220,N_11794,N_11896);
or U12221 (N_12221,N_11865,N_11985);
xor U12222 (N_12222,N_11939,N_11897);
xor U12223 (N_12223,N_11968,N_11929);
xnor U12224 (N_12224,N_11882,N_11871);
and U12225 (N_12225,N_11818,N_11966);
xor U12226 (N_12226,N_11955,N_11784);
or U12227 (N_12227,N_11931,N_11953);
nor U12228 (N_12228,N_11965,N_11896);
nor U12229 (N_12229,N_11913,N_11837);
xor U12230 (N_12230,N_11867,N_11929);
or U12231 (N_12231,N_11841,N_11919);
nand U12232 (N_12232,N_11919,N_11998);
or U12233 (N_12233,N_11955,N_11838);
xor U12234 (N_12234,N_11906,N_11822);
and U12235 (N_12235,N_11855,N_11788);
xor U12236 (N_12236,N_11990,N_11755);
nor U12237 (N_12237,N_11907,N_11816);
nor U12238 (N_12238,N_11786,N_11828);
nand U12239 (N_12239,N_11770,N_11873);
xnor U12240 (N_12240,N_11869,N_11778);
xnor U12241 (N_12241,N_11823,N_11933);
nor U12242 (N_12242,N_11983,N_11824);
or U12243 (N_12243,N_11837,N_11993);
xor U12244 (N_12244,N_11906,N_11764);
xor U12245 (N_12245,N_11910,N_11852);
nor U12246 (N_12246,N_11996,N_11915);
xor U12247 (N_12247,N_11769,N_11925);
or U12248 (N_12248,N_11821,N_11853);
and U12249 (N_12249,N_11788,N_11805);
nor U12250 (N_12250,N_12105,N_12113);
nand U12251 (N_12251,N_12156,N_12110);
and U12252 (N_12252,N_12198,N_12210);
nand U12253 (N_12253,N_12245,N_12218);
nand U12254 (N_12254,N_12169,N_12197);
xor U12255 (N_12255,N_12171,N_12058);
nand U12256 (N_12256,N_12075,N_12200);
nand U12257 (N_12257,N_12001,N_12055);
nor U12258 (N_12258,N_12117,N_12107);
xnor U12259 (N_12259,N_12042,N_12209);
and U12260 (N_12260,N_12114,N_12219);
xnor U12261 (N_12261,N_12004,N_12237);
xor U12262 (N_12262,N_12181,N_12191);
or U12263 (N_12263,N_12227,N_12241);
or U12264 (N_12264,N_12080,N_12024);
xor U12265 (N_12265,N_12231,N_12192);
and U12266 (N_12266,N_12036,N_12230);
or U12267 (N_12267,N_12053,N_12244);
or U12268 (N_12268,N_12132,N_12205);
nand U12269 (N_12269,N_12246,N_12170);
or U12270 (N_12270,N_12025,N_12070);
or U12271 (N_12271,N_12199,N_12222);
or U12272 (N_12272,N_12161,N_12130);
xnor U12273 (N_12273,N_12081,N_12176);
or U12274 (N_12274,N_12060,N_12138);
nand U12275 (N_12275,N_12018,N_12248);
nand U12276 (N_12276,N_12046,N_12247);
or U12277 (N_12277,N_12163,N_12229);
nand U12278 (N_12278,N_12011,N_12065);
xor U12279 (N_12279,N_12103,N_12104);
or U12280 (N_12280,N_12097,N_12196);
and U12281 (N_12281,N_12056,N_12108);
nor U12282 (N_12282,N_12158,N_12094);
and U12283 (N_12283,N_12189,N_12021);
xnor U12284 (N_12284,N_12002,N_12249);
xor U12285 (N_12285,N_12096,N_12214);
xnor U12286 (N_12286,N_12217,N_12016);
nand U12287 (N_12287,N_12050,N_12185);
nor U12288 (N_12288,N_12093,N_12022);
nand U12289 (N_12289,N_12092,N_12008);
or U12290 (N_12290,N_12146,N_12121);
and U12291 (N_12291,N_12013,N_12137);
and U12292 (N_12292,N_12115,N_12051);
xnor U12293 (N_12293,N_12165,N_12076);
and U12294 (N_12294,N_12236,N_12220);
and U12295 (N_12295,N_12005,N_12116);
and U12296 (N_12296,N_12153,N_12187);
and U12297 (N_12297,N_12106,N_12045);
and U12298 (N_12298,N_12054,N_12135);
nand U12299 (N_12299,N_12172,N_12186);
nand U12300 (N_12300,N_12047,N_12149);
or U12301 (N_12301,N_12071,N_12086);
nand U12302 (N_12302,N_12202,N_12152);
or U12303 (N_12303,N_12240,N_12059);
nand U12304 (N_12304,N_12033,N_12133);
nor U12305 (N_12305,N_12194,N_12098);
xor U12306 (N_12306,N_12029,N_12041);
xor U12307 (N_12307,N_12141,N_12061);
xnor U12308 (N_12308,N_12213,N_12083);
nand U12309 (N_12309,N_12111,N_12216);
nor U12310 (N_12310,N_12040,N_12073);
xor U12311 (N_12311,N_12228,N_12195);
nor U12312 (N_12312,N_12118,N_12147);
or U12313 (N_12313,N_12234,N_12242);
xnor U12314 (N_12314,N_12221,N_12090);
nor U12315 (N_12315,N_12188,N_12159);
and U12316 (N_12316,N_12078,N_12072);
and U12317 (N_12317,N_12067,N_12112);
nand U12318 (N_12318,N_12063,N_12175);
xor U12319 (N_12319,N_12035,N_12123);
xor U12320 (N_12320,N_12007,N_12150);
or U12321 (N_12321,N_12140,N_12155);
and U12322 (N_12322,N_12226,N_12183);
nand U12323 (N_12323,N_12032,N_12085);
xor U12324 (N_12324,N_12026,N_12157);
nor U12325 (N_12325,N_12206,N_12239);
or U12326 (N_12326,N_12243,N_12139);
xor U12327 (N_12327,N_12162,N_12212);
and U12328 (N_12328,N_12109,N_12144);
xnor U12329 (N_12329,N_12173,N_12142);
and U12330 (N_12330,N_12148,N_12178);
nor U12331 (N_12331,N_12120,N_12174);
or U12332 (N_12332,N_12020,N_12037);
nor U12333 (N_12333,N_12043,N_12126);
or U12334 (N_12334,N_12238,N_12203);
xnor U12335 (N_12335,N_12034,N_12164);
or U12336 (N_12336,N_12128,N_12100);
nand U12337 (N_12337,N_12160,N_12048);
nor U12338 (N_12338,N_12136,N_12177);
nand U12339 (N_12339,N_12014,N_12211);
or U12340 (N_12340,N_12235,N_12028);
xor U12341 (N_12341,N_12204,N_12030);
xnor U12342 (N_12342,N_12180,N_12038);
xnor U12343 (N_12343,N_12124,N_12031);
nor U12344 (N_12344,N_12077,N_12062);
nor U12345 (N_12345,N_12134,N_12215);
nor U12346 (N_12346,N_12099,N_12145);
nand U12347 (N_12347,N_12015,N_12232);
nor U12348 (N_12348,N_12208,N_12207);
xor U12349 (N_12349,N_12131,N_12088);
xor U12350 (N_12350,N_12066,N_12010);
and U12351 (N_12351,N_12069,N_12023);
or U12352 (N_12352,N_12068,N_12052);
and U12353 (N_12353,N_12087,N_12074);
nor U12354 (N_12354,N_12057,N_12019);
nor U12355 (N_12355,N_12039,N_12223);
nand U12356 (N_12356,N_12224,N_12000);
xor U12357 (N_12357,N_12184,N_12166);
xnor U12358 (N_12358,N_12084,N_12179);
and U12359 (N_12359,N_12091,N_12017);
and U12360 (N_12360,N_12102,N_12044);
and U12361 (N_12361,N_12129,N_12095);
nor U12362 (N_12362,N_12201,N_12233);
nand U12363 (N_12363,N_12143,N_12167);
xnor U12364 (N_12364,N_12027,N_12127);
nor U12365 (N_12365,N_12193,N_12182);
nand U12366 (N_12366,N_12009,N_12079);
and U12367 (N_12367,N_12154,N_12049);
or U12368 (N_12368,N_12168,N_12003);
nand U12369 (N_12369,N_12125,N_12012);
and U12370 (N_12370,N_12101,N_12082);
nor U12371 (N_12371,N_12064,N_12089);
xnor U12372 (N_12372,N_12151,N_12225);
and U12373 (N_12373,N_12119,N_12190);
nor U12374 (N_12374,N_12122,N_12006);
nand U12375 (N_12375,N_12235,N_12213);
and U12376 (N_12376,N_12038,N_12055);
nand U12377 (N_12377,N_12169,N_12221);
nor U12378 (N_12378,N_12151,N_12156);
and U12379 (N_12379,N_12078,N_12013);
and U12380 (N_12380,N_12051,N_12089);
nand U12381 (N_12381,N_12066,N_12157);
nand U12382 (N_12382,N_12192,N_12108);
xor U12383 (N_12383,N_12056,N_12212);
nand U12384 (N_12384,N_12093,N_12206);
and U12385 (N_12385,N_12132,N_12202);
and U12386 (N_12386,N_12037,N_12003);
xnor U12387 (N_12387,N_12088,N_12184);
nand U12388 (N_12388,N_12119,N_12242);
xnor U12389 (N_12389,N_12140,N_12222);
and U12390 (N_12390,N_12072,N_12017);
and U12391 (N_12391,N_12228,N_12246);
nor U12392 (N_12392,N_12004,N_12215);
nand U12393 (N_12393,N_12100,N_12094);
or U12394 (N_12394,N_12178,N_12010);
nor U12395 (N_12395,N_12156,N_12194);
or U12396 (N_12396,N_12101,N_12091);
nor U12397 (N_12397,N_12073,N_12162);
nand U12398 (N_12398,N_12240,N_12152);
or U12399 (N_12399,N_12100,N_12189);
or U12400 (N_12400,N_12236,N_12222);
xor U12401 (N_12401,N_12036,N_12185);
nor U12402 (N_12402,N_12102,N_12001);
xor U12403 (N_12403,N_12181,N_12167);
xnor U12404 (N_12404,N_12151,N_12236);
or U12405 (N_12405,N_12031,N_12042);
or U12406 (N_12406,N_12042,N_12196);
or U12407 (N_12407,N_12056,N_12038);
xor U12408 (N_12408,N_12086,N_12229);
or U12409 (N_12409,N_12052,N_12166);
nand U12410 (N_12410,N_12005,N_12147);
nor U12411 (N_12411,N_12235,N_12132);
nand U12412 (N_12412,N_12046,N_12157);
and U12413 (N_12413,N_12013,N_12241);
or U12414 (N_12414,N_12148,N_12135);
nand U12415 (N_12415,N_12012,N_12124);
nand U12416 (N_12416,N_12218,N_12150);
nand U12417 (N_12417,N_12249,N_12084);
nand U12418 (N_12418,N_12156,N_12154);
nand U12419 (N_12419,N_12162,N_12238);
or U12420 (N_12420,N_12216,N_12039);
xor U12421 (N_12421,N_12248,N_12176);
or U12422 (N_12422,N_12175,N_12033);
or U12423 (N_12423,N_12243,N_12052);
xnor U12424 (N_12424,N_12019,N_12091);
or U12425 (N_12425,N_12066,N_12131);
or U12426 (N_12426,N_12230,N_12136);
xor U12427 (N_12427,N_12007,N_12136);
and U12428 (N_12428,N_12090,N_12227);
nand U12429 (N_12429,N_12161,N_12200);
or U12430 (N_12430,N_12063,N_12043);
nand U12431 (N_12431,N_12214,N_12083);
or U12432 (N_12432,N_12170,N_12228);
nor U12433 (N_12433,N_12135,N_12068);
or U12434 (N_12434,N_12139,N_12125);
and U12435 (N_12435,N_12171,N_12121);
or U12436 (N_12436,N_12113,N_12074);
nor U12437 (N_12437,N_12101,N_12025);
and U12438 (N_12438,N_12211,N_12176);
nor U12439 (N_12439,N_12172,N_12214);
nor U12440 (N_12440,N_12150,N_12219);
xnor U12441 (N_12441,N_12176,N_12011);
and U12442 (N_12442,N_12121,N_12091);
or U12443 (N_12443,N_12194,N_12202);
xnor U12444 (N_12444,N_12231,N_12012);
nor U12445 (N_12445,N_12206,N_12079);
and U12446 (N_12446,N_12154,N_12054);
nor U12447 (N_12447,N_12167,N_12032);
xor U12448 (N_12448,N_12031,N_12115);
nor U12449 (N_12449,N_12155,N_12239);
xnor U12450 (N_12450,N_12094,N_12231);
nor U12451 (N_12451,N_12136,N_12061);
xor U12452 (N_12452,N_12154,N_12221);
or U12453 (N_12453,N_12101,N_12113);
nand U12454 (N_12454,N_12144,N_12056);
or U12455 (N_12455,N_12111,N_12026);
and U12456 (N_12456,N_12116,N_12213);
nand U12457 (N_12457,N_12176,N_12094);
nand U12458 (N_12458,N_12187,N_12123);
or U12459 (N_12459,N_12232,N_12192);
or U12460 (N_12460,N_12008,N_12024);
nand U12461 (N_12461,N_12233,N_12020);
nor U12462 (N_12462,N_12244,N_12227);
and U12463 (N_12463,N_12218,N_12222);
and U12464 (N_12464,N_12068,N_12059);
and U12465 (N_12465,N_12071,N_12025);
nand U12466 (N_12466,N_12230,N_12219);
xor U12467 (N_12467,N_12060,N_12220);
nand U12468 (N_12468,N_12168,N_12162);
xor U12469 (N_12469,N_12059,N_12030);
nand U12470 (N_12470,N_12035,N_12040);
or U12471 (N_12471,N_12218,N_12091);
nor U12472 (N_12472,N_12214,N_12193);
nand U12473 (N_12473,N_12098,N_12153);
or U12474 (N_12474,N_12086,N_12161);
or U12475 (N_12475,N_12249,N_12123);
nand U12476 (N_12476,N_12227,N_12169);
or U12477 (N_12477,N_12151,N_12120);
or U12478 (N_12478,N_12101,N_12075);
or U12479 (N_12479,N_12099,N_12188);
nand U12480 (N_12480,N_12048,N_12248);
and U12481 (N_12481,N_12215,N_12095);
nand U12482 (N_12482,N_12024,N_12104);
nor U12483 (N_12483,N_12054,N_12079);
or U12484 (N_12484,N_12040,N_12110);
nor U12485 (N_12485,N_12075,N_12073);
xnor U12486 (N_12486,N_12006,N_12028);
xnor U12487 (N_12487,N_12099,N_12212);
and U12488 (N_12488,N_12108,N_12244);
or U12489 (N_12489,N_12085,N_12114);
or U12490 (N_12490,N_12226,N_12175);
xnor U12491 (N_12491,N_12070,N_12077);
or U12492 (N_12492,N_12068,N_12192);
or U12493 (N_12493,N_12062,N_12113);
nor U12494 (N_12494,N_12018,N_12150);
nand U12495 (N_12495,N_12167,N_12182);
nand U12496 (N_12496,N_12201,N_12118);
nand U12497 (N_12497,N_12104,N_12071);
or U12498 (N_12498,N_12085,N_12003);
nor U12499 (N_12499,N_12084,N_12003);
or U12500 (N_12500,N_12420,N_12427);
nand U12501 (N_12501,N_12251,N_12412);
nor U12502 (N_12502,N_12293,N_12326);
nor U12503 (N_12503,N_12265,N_12305);
or U12504 (N_12504,N_12463,N_12466);
xor U12505 (N_12505,N_12302,N_12409);
or U12506 (N_12506,N_12378,N_12276);
xor U12507 (N_12507,N_12356,N_12289);
or U12508 (N_12508,N_12348,N_12454);
nor U12509 (N_12509,N_12382,N_12380);
or U12510 (N_12510,N_12373,N_12390);
nor U12511 (N_12511,N_12467,N_12465);
nor U12512 (N_12512,N_12271,N_12440);
xnor U12513 (N_12513,N_12284,N_12333);
nand U12514 (N_12514,N_12350,N_12272);
or U12515 (N_12515,N_12482,N_12349);
or U12516 (N_12516,N_12419,N_12285);
nor U12517 (N_12517,N_12343,N_12258);
nand U12518 (N_12518,N_12321,N_12329);
nor U12519 (N_12519,N_12376,N_12460);
and U12520 (N_12520,N_12307,N_12354);
nand U12521 (N_12521,N_12352,N_12328);
nand U12522 (N_12522,N_12297,N_12404);
nand U12523 (N_12523,N_12322,N_12336);
nor U12524 (N_12524,N_12488,N_12264);
nor U12525 (N_12525,N_12342,N_12282);
or U12526 (N_12526,N_12447,N_12345);
nor U12527 (N_12527,N_12439,N_12372);
and U12528 (N_12528,N_12444,N_12394);
and U12529 (N_12529,N_12387,N_12499);
or U12530 (N_12530,N_12263,N_12492);
nor U12531 (N_12531,N_12250,N_12386);
nor U12532 (N_12532,N_12381,N_12323);
and U12533 (N_12533,N_12410,N_12429);
nor U12534 (N_12534,N_12461,N_12411);
or U12535 (N_12535,N_12291,N_12423);
xor U12536 (N_12536,N_12455,N_12487);
nor U12537 (N_12537,N_12457,N_12298);
and U12538 (N_12538,N_12421,N_12320);
xor U12539 (N_12539,N_12377,N_12344);
or U12540 (N_12540,N_12490,N_12474);
or U12541 (N_12541,N_12456,N_12355);
nor U12542 (N_12542,N_12464,N_12395);
nand U12543 (N_12543,N_12443,N_12473);
or U12544 (N_12544,N_12300,N_12310);
nand U12545 (N_12545,N_12476,N_12366);
nor U12546 (N_12546,N_12277,N_12491);
and U12547 (N_12547,N_12257,N_12294);
nand U12548 (N_12548,N_12485,N_12253);
nand U12549 (N_12549,N_12475,N_12256);
or U12550 (N_12550,N_12296,N_12498);
or U12551 (N_12551,N_12311,N_12408);
xor U12552 (N_12552,N_12288,N_12406);
nor U12553 (N_12553,N_12340,N_12337);
xnor U12554 (N_12554,N_12434,N_12259);
or U12555 (N_12555,N_12332,N_12339);
xnor U12556 (N_12556,N_12407,N_12325);
xnor U12557 (N_12557,N_12384,N_12270);
and U12558 (N_12558,N_12433,N_12252);
or U12559 (N_12559,N_12334,N_12260);
nand U12560 (N_12560,N_12292,N_12335);
and U12561 (N_12561,N_12458,N_12414);
nand U12562 (N_12562,N_12254,N_12255);
nor U12563 (N_12563,N_12317,N_12379);
nor U12564 (N_12564,N_12315,N_12309);
nor U12565 (N_12565,N_12301,N_12306);
nor U12566 (N_12566,N_12481,N_12383);
or U12567 (N_12567,N_12389,N_12459);
or U12568 (N_12568,N_12374,N_12451);
and U12569 (N_12569,N_12478,N_12484);
nor U12570 (N_12570,N_12422,N_12330);
or U12571 (N_12571,N_12338,N_12278);
nand U12572 (N_12572,N_12331,N_12393);
or U12573 (N_12573,N_12425,N_12341);
nor U12574 (N_12574,N_12452,N_12415);
or U12575 (N_12575,N_12402,N_12369);
nor U12576 (N_12576,N_12364,N_12483);
nor U12577 (N_12577,N_12426,N_12280);
or U12578 (N_12578,N_12391,N_12290);
nor U12579 (N_12579,N_12432,N_12400);
and U12580 (N_12580,N_12442,N_12324);
nand U12581 (N_12581,N_12262,N_12281);
nor U12582 (N_12582,N_12267,N_12497);
nand U12583 (N_12583,N_12295,N_12495);
and U12584 (N_12584,N_12362,N_12441);
xor U12585 (N_12585,N_12449,N_12494);
and U12586 (N_12586,N_12275,N_12357);
xor U12587 (N_12587,N_12359,N_12268);
xor U12588 (N_12588,N_12279,N_12468);
and U12589 (N_12589,N_12477,N_12417);
and U12590 (N_12590,N_12450,N_12388);
and U12591 (N_12591,N_12418,N_12453);
nand U12592 (N_12592,N_12399,N_12401);
or U12593 (N_12593,N_12486,N_12318);
nand U12594 (N_12594,N_12435,N_12431);
or U12595 (N_12595,N_12358,N_12385);
xnor U12596 (N_12596,N_12303,N_12375);
nand U12597 (N_12597,N_12286,N_12405);
nand U12598 (N_12598,N_12313,N_12274);
xnor U12599 (N_12599,N_12496,N_12308);
nor U12600 (N_12600,N_12283,N_12438);
xnor U12601 (N_12601,N_12365,N_12446);
nand U12602 (N_12602,N_12370,N_12469);
xnor U12603 (N_12603,N_12430,N_12493);
or U12604 (N_12604,N_12368,N_12304);
and U12605 (N_12605,N_12360,N_12269);
nand U12606 (N_12606,N_12428,N_12489);
or U12607 (N_12607,N_12445,N_12448);
nand U12608 (N_12608,N_12397,N_12437);
nor U12609 (N_12609,N_12312,N_12462);
nand U12610 (N_12610,N_12371,N_12363);
xor U12611 (N_12611,N_12479,N_12480);
or U12612 (N_12612,N_12351,N_12471);
nand U12613 (N_12613,N_12319,N_12299);
and U12614 (N_12614,N_12413,N_12314);
nand U12615 (N_12615,N_12273,N_12346);
xnor U12616 (N_12616,N_12392,N_12472);
xnor U12617 (N_12617,N_12347,N_12266);
and U12618 (N_12618,N_12287,N_12367);
nor U12619 (N_12619,N_12396,N_12361);
and U12620 (N_12620,N_12316,N_12436);
xnor U12621 (N_12621,N_12327,N_12398);
nor U12622 (N_12622,N_12424,N_12353);
or U12623 (N_12623,N_12261,N_12470);
nor U12624 (N_12624,N_12416,N_12403);
xor U12625 (N_12625,N_12407,N_12438);
xnor U12626 (N_12626,N_12394,N_12253);
and U12627 (N_12627,N_12496,N_12325);
xnor U12628 (N_12628,N_12409,N_12438);
or U12629 (N_12629,N_12363,N_12268);
nand U12630 (N_12630,N_12263,N_12316);
or U12631 (N_12631,N_12492,N_12435);
or U12632 (N_12632,N_12464,N_12390);
nor U12633 (N_12633,N_12309,N_12256);
and U12634 (N_12634,N_12491,N_12467);
and U12635 (N_12635,N_12276,N_12368);
and U12636 (N_12636,N_12323,N_12387);
and U12637 (N_12637,N_12369,N_12401);
nor U12638 (N_12638,N_12385,N_12499);
and U12639 (N_12639,N_12256,N_12499);
and U12640 (N_12640,N_12431,N_12400);
xor U12641 (N_12641,N_12254,N_12306);
nand U12642 (N_12642,N_12465,N_12417);
or U12643 (N_12643,N_12459,N_12303);
nor U12644 (N_12644,N_12250,N_12453);
nand U12645 (N_12645,N_12484,N_12326);
or U12646 (N_12646,N_12306,N_12366);
or U12647 (N_12647,N_12342,N_12268);
nor U12648 (N_12648,N_12326,N_12289);
or U12649 (N_12649,N_12327,N_12385);
and U12650 (N_12650,N_12470,N_12279);
or U12651 (N_12651,N_12372,N_12369);
or U12652 (N_12652,N_12324,N_12322);
xnor U12653 (N_12653,N_12268,N_12334);
nor U12654 (N_12654,N_12470,N_12296);
or U12655 (N_12655,N_12290,N_12464);
xor U12656 (N_12656,N_12450,N_12387);
and U12657 (N_12657,N_12424,N_12301);
nor U12658 (N_12658,N_12295,N_12329);
xnor U12659 (N_12659,N_12471,N_12274);
and U12660 (N_12660,N_12405,N_12437);
or U12661 (N_12661,N_12371,N_12332);
nand U12662 (N_12662,N_12359,N_12315);
or U12663 (N_12663,N_12400,N_12375);
and U12664 (N_12664,N_12483,N_12281);
nor U12665 (N_12665,N_12275,N_12397);
nand U12666 (N_12666,N_12267,N_12340);
xnor U12667 (N_12667,N_12450,N_12331);
nor U12668 (N_12668,N_12478,N_12440);
nor U12669 (N_12669,N_12388,N_12310);
nor U12670 (N_12670,N_12358,N_12493);
or U12671 (N_12671,N_12392,N_12262);
xor U12672 (N_12672,N_12358,N_12337);
nor U12673 (N_12673,N_12426,N_12421);
xor U12674 (N_12674,N_12315,N_12431);
xor U12675 (N_12675,N_12393,N_12463);
and U12676 (N_12676,N_12444,N_12385);
nor U12677 (N_12677,N_12326,N_12367);
xnor U12678 (N_12678,N_12267,N_12399);
nor U12679 (N_12679,N_12413,N_12280);
nand U12680 (N_12680,N_12490,N_12499);
nand U12681 (N_12681,N_12474,N_12292);
nand U12682 (N_12682,N_12467,N_12356);
nand U12683 (N_12683,N_12317,N_12275);
nand U12684 (N_12684,N_12467,N_12442);
nand U12685 (N_12685,N_12410,N_12467);
nor U12686 (N_12686,N_12332,N_12375);
nand U12687 (N_12687,N_12424,N_12398);
xor U12688 (N_12688,N_12276,N_12324);
nor U12689 (N_12689,N_12325,N_12323);
and U12690 (N_12690,N_12379,N_12441);
and U12691 (N_12691,N_12410,N_12469);
nor U12692 (N_12692,N_12325,N_12255);
or U12693 (N_12693,N_12363,N_12401);
and U12694 (N_12694,N_12424,N_12346);
and U12695 (N_12695,N_12497,N_12395);
or U12696 (N_12696,N_12485,N_12438);
and U12697 (N_12697,N_12314,N_12291);
nand U12698 (N_12698,N_12469,N_12355);
or U12699 (N_12699,N_12497,N_12490);
or U12700 (N_12700,N_12277,N_12408);
xnor U12701 (N_12701,N_12304,N_12425);
or U12702 (N_12702,N_12436,N_12327);
nor U12703 (N_12703,N_12268,N_12432);
xor U12704 (N_12704,N_12315,N_12403);
or U12705 (N_12705,N_12416,N_12261);
xnor U12706 (N_12706,N_12492,N_12290);
nor U12707 (N_12707,N_12286,N_12309);
and U12708 (N_12708,N_12310,N_12332);
xor U12709 (N_12709,N_12324,N_12289);
and U12710 (N_12710,N_12421,N_12377);
xor U12711 (N_12711,N_12273,N_12345);
xnor U12712 (N_12712,N_12331,N_12484);
and U12713 (N_12713,N_12331,N_12347);
nand U12714 (N_12714,N_12272,N_12354);
nor U12715 (N_12715,N_12269,N_12321);
nand U12716 (N_12716,N_12286,N_12380);
or U12717 (N_12717,N_12456,N_12350);
and U12718 (N_12718,N_12474,N_12395);
nand U12719 (N_12719,N_12397,N_12444);
and U12720 (N_12720,N_12412,N_12277);
xnor U12721 (N_12721,N_12301,N_12494);
nor U12722 (N_12722,N_12452,N_12397);
xor U12723 (N_12723,N_12276,N_12263);
xor U12724 (N_12724,N_12342,N_12402);
or U12725 (N_12725,N_12433,N_12423);
xor U12726 (N_12726,N_12474,N_12302);
xnor U12727 (N_12727,N_12299,N_12284);
or U12728 (N_12728,N_12364,N_12343);
xnor U12729 (N_12729,N_12257,N_12490);
nand U12730 (N_12730,N_12407,N_12301);
nor U12731 (N_12731,N_12342,N_12397);
or U12732 (N_12732,N_12300,N_12376);
nor U12733 (N_12733,N_12306,N_12278);
nor U12734 (N_12734,N_12402,N_12394);
and U12735 (N_12735,N_12458,N_12431);
and U12736 (N_12736,N_12415,N_12332);
and U12737 (N_12737,N_12346,N_12423);
and U12738 (N_12738,N_12253,N_12415);
xnor U12739 (N_12739,N_12398,N_12415);
or U12740 (N_12740,N_12371,N_12309);
or U12741 (N_12741,N_12495,N_12381);
and U12742 (N_12742,N_12329,N_12263);
xor U12743 (N_12743,N_12297,N_12357);
nand U12744 (N_12744,N_12310,N_12351);
or U12745 (N_12745,N_12398,N_12270);
and U12746 (N_12746,N_12476,N_12372);
and U12747 (N_12747,N_12268,N_12310);
and U12748 (N_12748,N_12343,N_12422);
and U12749 (N_12749,N_12402,N_12344);
nor U12750 (N_12750,N_12500,N_12654);
nand U12751 (N_12751,N_12560,N_12684);
nand U12752 (N_12752,N_12715,N_12539);
nor U12753 (N_12753,N_12723,N_12698);
nand U12754 (N_12754,N_12600,N_12669);
xnor U12755 (N_12755,N_12635,N_12542);
and U12756 (N_12756,N_12555,N_12725);
and U12757 (N_12757,N_12601,N_12716);
or U12758 (N_12758,N_12507,N_12605);
or U12759 (N_12759,N_12590,N_12674);
xnor U12760 (N_12760,N_12556,N_12672);
nand U12761 (N_12761,N_12705,N_12623);
nand U12762 (N_12762,N_12610,N_12718);
xnor U12763 (N_12763,N_12522,N_12594);
nand U12764 (N_12764,N_12593,N_12614);
or U12765 (N_12765,N_12652,N_12563);
nand U12766 (N_12766,N_12648,N_12588);
nand U12767 (N_12767,N_12641,N_12526);
xor U12768 (N_12768,N_12587,N_12671);
or U12769 (N_12769,N_12683,N_12565);
or U12770 (N_12770,N_12537,N_12509);
and U12771 (N_12771,N_12735,N_12711);
nand U12772 (N_12772,N_12746,N_12665);
nand U12773 (N_12773,N_12659,N_12679);
and U12774 (N_12774,N_12704,N_12667);
xor U12775 (N_12775,N_12739,N_12714);
xor U12776 (N_12776,N_12620,N_12632);
or U12777 (N_12777,N_12708,N_12727);
or U12778 (N_12778,N_12651,N_12677);
nor U12779 (N_12779,N_12567,N_12645);
nor U12780 (N_12780,N_12628,N_12685);
or U12781 (N_12781,N_12637,N_12657);
nand U12782 (N_12782,N_12630,N_12535);
or U12783 (N_12783,N_12569,N_12707);
nand U12784 (N_12784,N_12749,N_12599);
or U12785 (N_12785,N_12661,N_12547);
or U12786 (N_12786,N_12639,N_12688);
and U12787 (N_12787,N_12607,N_12673);
or U12788 (N_12788,N_12681,N_12619);
nor U12789 (N_12789,N_12602,N_12742);
nor U12790 (N_12790,N_12622,N_12655);
xor U12791 (N_12791,N_12699,N_12616);
nor U12792 (N_12792,N_12670,N_12734);
nor U12793 (N_12793,N_12695,N_12540);
nor U12794 (N_12794,N_12702,N_12501);
nor U12795 (N_12795,N_12516,N_12611);
nor U12796 (N_12796,N_12730,N_12524);
nor U12797 (N_12797,N_12576,N_12744);
or U12798 (N_12798,N_12731,N_12517);
xnor U12799 (N_12799,N_12544,N_12696);
nor U12800 (N_12800,N_12738,N_12710);
and U12801 (N_12801,N_12643,N_12553);
and U12802 (N_12802,N_12728,N_12658);
and U12803 (N_12803,N_12687,N_12678);
xor U12804 (N_12804,N_12660,N_12519);
nor U12805 (N_12805,N_12512,N_12724);
nor U12806 (N_12806,N_12558,N_12546);
nand U12807 (N_12807,N_12664,N_12515);
and U12808 (N_12808,N_12656,N_12733);
nor U12809 (N_12809,N_12533,N_12634);
xor U12810 (N_12810,N_12580,N_12548);
nor U12811 (N_12811,N_12729,N_12649);
nand U12812 (N_12812,N_12668,N_12653);
xnor U12813 (N_12813,N_12529,N_12748);
nand U12814 (N_12814,N_12527,N_12726);
or U12815 (N_12815,N_12518,N_12712);
and U12816 (N_12816,N_12609,N_12709);
and U12817 (N_12817,N_12650,N_12581);
xnor U12818 (N_12818,N_12640,N_12525);
or U12819 (N_12819,N_12638,N_12564);
xnor U12820 (N_12820,N_12736,N_12692);
or U12821 (N_12821,N_12502,N_12575);
xor U12822 (N_12822,N_12644,N_12545);
nand U12823 (N_12823,N_12720,N_12552);
nor U12824 (N_12824,N_12697,N_12597);
xor U12825 (N_12825,N_12586,N_12625);
xor U12826 (N_12826,N_12603,N_12561);
or U12827 (N_12827,N_12506,N_12618);
nor U12828 (N_12828,N_12520,N_12570);
nor U12829 (N_12829,N_12680,N_12617);
nand U12830 (N_12830,N_12568,N_12740);
and U12831 (N_12831,N_12737,N_12666);
xor U12832 (N_12832,N_12528,N_12574);
and U12833 (N_12833,N_12557,N_12589);
and U12834 (N_12834,N_12510,N_12689);
nand U12835 (N_12835,N_12534,N_12741);
nand U12836 (N_12836,N_12703,N_12538);
nor U12837 (N_12837,N_12722,N_12541);
nor U12838 (N_12838,N_12682,N_12700);
nor U12839 (N_12839,N_12503,N_12584);
nand U12840 (N_12840,N_12579,N_12615);
or U12841 (N_12841,N_12591,N_12662);
and U12842 (N_12842,N_12642,N_12554);
nor U12843 (N_12843,N_12571,N_12612);
nor U12844 (N_12844,N_12631,N_12585);
xor U12845 (N_12845,N_12536,N_12592);
nand U12846 (N_12846,N_12549,N_12573);
nor U12847 (N_12847,N_12691,N_12531);
nand U12848 (N_12848,N_12606,N_12627);
nand U12849 (N_12849,N_12747,N_12604);
xnor U12850 (N_12850,N_12636,N_12582);
and U12851 (N_12851,N_12523,N_12717);
and U12852 (N_12852,N_12513,N_12694);
and U12853 (N_12853,N_12583,N_12701);
xor U12854 (N_12854,N_12596,N_12732);
nand U12855 (N_12855,N_12504,N_12647);
and U12856 (N_12856,N_12562,N_12508);
nand U12857 (N_12857,N_12663,N_12543);
nand U12858 (N_12858,N_12721,N_12706);
xnor U12859 (N_12859,N_12745,N_12646);
xor U12860 (N_12860,N_12505,N_12690);
xor U12861 (N_12861,N_12613,N_12514);
or U12862 (N_12862,N_12566,N_12511);
and U12863 (N_12863,N_12693,N_12572);
xor U12864 (N_12864,N_12621,N_12578);
nand U12865 (N_12865,N_12577,N_12550);
and U12866 (N_12866,N_12598,N_12713);
xnor U12867 (N_12867,N_12532,N_12559);
or U12868 (N_12868,N_12551,N_12675);
and U12869 (N_12869,N_12624,N_12676);
or U12870 (N_12870,N_12629,N_12595);
nand U12871 (N_12871,N_12608,N_12743);
nand U12872 (N_12872,N_12686,N_12626);
nand U12873 (N_12873,N_12530,N_12633);
nand U12874 (N_12874,N_12719,N_12521);
or U12875 (N_12875,N_12591,N_12689);
or U12876 (N_12876,N_12607,N_12682);
and U12877 (N_12877,N_12696,N_12580);
and U12878 (N_12878,N_12633,N_12678);
nand U12879 (N_12879,N_12634,N_12611);
nor U12880 (N_12880,N_12725,N_12744);
xnor U12881 (N_12881,N_12535,N_12698);
nor U12882 (N_12882,N_12583,N_12634);
xnor U12883 (N_12883,N_12723,N_12550);
xnor U12884 (N_12884,N_12593,N_12697);
and U12885 (N_12885,N_12652,N_12608);
xnor U12886 (N_12886,N_12585,N_12525);
xnor U12887 (N_12887,N_12517,N_12519);
or U12888 (N_12888,N_12511,N_12728);
nand U12889 (N_12889,N_12664,N_12529);
or U12890 (N_12890,N_12721,N_12711);
and U12891 (N_12891,N_12627,N_12659);
nand U12892 (N_12892,N_12558,N_12656);
or U12893 (N_12893,N_12651,N_12639);
xor U12894 (N_12894,N_12604,N_12697);
and U12895 (N_12895,N_12683,N_12534);
nand U12896 (N_12896,N_12721,N_12730);
nand U12897 (N_12897,N_12671,N_12731);
nor U12898 (N_12898,N_12696,N_12510);
nor U12899 (N_12899,N_12537,N_12647);
or U12900 (N_12900,N_12735,N_12596);
nor U12901 (N_12901,N_12634,N_12500);
xnor U12902 (N_12902,N_12556,N_12666);
or U12903 (N_12903,N_12654,N_12525);
or U12904 (N_12904,N_12734,N_12710);
nor U12905 (N_12905,N_12572,N_12729);
nand U12906 (N_12906,N_12739,N_12677);
xnor U12907 (N_12907,N_12649,N_12739);
nor U12908 (N_12908,N_12701,N_12652);
xnor U12909 (N_12909,N_12719,N_12637);
xor U12910 (N_12910,N_12541,N_12659);
xnor U12911 (N_12911,N_12528,N_12604);
xor U12912 (N_12912,N_12575,N_12619);
nor U12913 (N_12913,N_12693,N_12652);
or U12914 (N_12914,N_12621,N_12675);
nor U12915 (N_12915,N_12742,N_12583);
nand U12916 (N_12916,N_12513,N_12673);
and U12917 (N_12917,N_12710,N_12611);
and U12918 (N_12918,N_12664,N_12506);
xnor U12919 (N_12919,N_12549,N_12594);
or U12920 (N_12920,N_12624,N_12640);
and U12921 (N_12921,N_12550,N_12691);
nand U12922 (N_12922,N_12564,N_12510);
nor U12923 (N_12923,N_12501,N_12695);
and U12924 (N_12924,N_12683,N_12572);
nor U12925 (N_12925,N_12518,N_12553);
or U12926 (N_12926,N_12683,N_12555);
xor U12927 (N_12927,N_12599,N_12720);
and U12928 (N_12928,N_12512,N_12672);
xnor U12929 (N_12929,N_12656,N_12653);
nand U12930 (N_12930,N_12593,N_12625);
nor U12931 (N_12931,N_12524,N_12663);
and U12932 (N_12932,N_12533,N_12531);
nor U12933 (N_12933,N_12725,N_12575);
xnor U12934 (N_12934,N_12740,N_12564);
xor U12935 (N_12935,N_12509,N_12618);
or U12936 (N_12936,N_12587,N_12502);
nand U12937 (N_12937,N_12676,N_12636);
or U12938 (N_12938,N_12704,N_12545);
nor U12939 (N_12939,N_12748,N_12729);
and U12940 (N_12940,N_12680,N_12716);
nand U12941 (N_12941,N_12510,N_12618);
and U12942 (N_12942,N_12603,N_12638);
and U12943 (N_12943,N_12590,N_12669);
or U12944 (N_12944,N_12712,N_12701);
xor U12945 (N_12945,N_12664,N_12582);
nor U12946 (N_12946,N_12521,N_12641);
xnor U12947 (N_12947,N_12500,N_12741);
or U12948 (N_12948,N_12581,N_12605);
xor U12949 (N_12949,N_12647,N_12584);
or U12950 (N_12950,N_12596,N_12744);
or U12951 (N_12951,N_12503,N_12541);
or U12952 (N_12952,N_12621,N_12721);
xnor U12953 (N_12953,N_12541,N_12674);
nor U12954 (N_12954,N_12643,N_12681);
or U12955 (N_12955,N_12510,N_12507);
and U12956 (N_12956,N_12576,N_12603);
nand U12957 (N_12957,N_12644,N_12710);
xnor U12958 (N_12958,N_12639,N_12608);
xnor U12959 (N_12959,N_12615,N_12705);
and U12960 (N_12960,N_12733,N_12699);
and U12961 (N_12961,N_12578,N_12611);
and U12962 (N_12962,N_12567,N_12545);
xnor U12963 (N_12963,N_12502,N_12535);
and U12964 (N_12964,N_12681,N_12536);
or U12965 (N_12965,N_12653,N_12677);
nor U12966 (N_12966,N_12709,N_12693);
nand U12967 (N_12967,N_12749,N_12748);
and U12968 (N_12968,N_12518,N_12521);
and U12969 (N_12969,N_12566,N_12738);
or U12970 (N_12970,N_12645,N_12719);
and U12971 (N_12971,N_12633,N_12718);
nor U12972 (N_12972,N_12566,N_12635);
nor U12973 (N_12973,N_12549,N_12512);
xnor U12974 (N_12974,N_12738,N_12659);
nor U12975 (N_12975,N_12580,N_12666);
xor U12976 (N_12976,N_12629,N_12505);
and U12977 (N_12977,N_12679,N_12698);
or U12978 (N_12978,N_12505,N_12710);
xnor U12979 (N_12979,N_12549,N_12532);
and U12980 (N_12980,N_12540,N_12595);
and U12981 (N_12981,N_12536,N_12523);
and U12982 (N_12982,N_12699,N_12553);
nor U12983 (N_12983,N_12614,N_12520);
xor U12984 (N_12984,N_12734,N_12723);
or U12985 (N_12985,N_12596,N_12581);
nand U12986 (N_12986,N_12503,N_12640);
and U12987 (N_12987,N_12728,N_12513);
nand U12988 (N_12988,N_12616,N_12544);
or U12989 (N_12989,N_12547,N_12677);
and U12990 (N_12990,N_12652,N_12658);
nor U12991 (N_12991,N_12611,N_12555);
nand U12992 (N_12992,N_12518,N_12622);
nand U12993 (N_12993,N_12742,N_12570);
xnor U12994 (N_12994,N_12577,N_12537);
or U12995 (N_12995,N_12738,N_12608);
or U12996 (N_12996,N_12735,N_12558);
and U12997 (N_12997,N_12710,N_12672);
nand U12998 (N_12998,N_12684,N_12654);
or U12999 (N_12999,N_12523,N_12749);
xor U13000 (N_13000,N_12761,N_12849);
xnor U13001 (N_13001,N_12962,N_12878);
and U13002 (N_13002,N_12846,N_12908);
or U13003 (N_13003,N_12756,N_12996);
and U13004 (N_13004,N_12824,N_12780);
or U13005 (N_13005,N_12788,N_12791);
and U13006 (N_13006,N_12966,N_12776);
nand U13007 (N_13007,N_12880,N_12903);
xor U13008 (N_13008,N_12939,N_12924);
or U13009 (N_13009,N_12796,N_12909);
nor U13010 (N_13010,N_12990,N_12921);
nor U13011 (N_13011,N_12840,N_12844);
or U13012 (N_13012,N_12853,N_12787);
nand U13013 (N_13013,N_12879,N_12792);
nand U13014 (N_13014,N_12960,N_12752);
xnor U13015 (N_13015,N_12816,N_12959);
nand U13016 (N_13016,N_12781,N_12976);
nor U13017 (N_13017,N_12968,N_12957);
nand U13018 (N_13018,N_12891,N_12809);
nor U13019 (N_13019,N_12907,N_12889);
nor U13020 (N_13020,N_12997,N_12805);
nor U13021 (N_13021,N_12902,N_12782);
xnor U13022 (N_13022,N_12911,N_12868);
xor U13023 (N_13023,N_12854,N_12810);
or U13024 (N_13024,N_12870,N_12825);
xnor U13025 (N_13025,N_12819,N_12794);
or U13026 (N_13026,N_12858,N_12926);
and U13027 (N_13027,N_12750,N_12951);
nand U13028 (N_13028,N_12998,N_12917);
or U13029 (N_13029,N_12871,N_12777);
nor U13030 (N_13030,N_12783,N_12949);
and U13031 (N_13031,N_12979,N_12847);
nand U13032 (N_13032,N_12892,N_12842);
and U13033 (N_13033,N_12835,N_12764);
nor U13034 (N_13034,N_12937,N_12793);
xor U13035 (N_13035,N_12839,N_12867);
xnor U13036 (N_13036,N_12888,N_12821);
nor U13037 (N_13037,N_12778,N_12934);
nand U13038 (N_13038,N_12947,N_12986);
or U13039 (N_13039,N_12914,N_12904);
and U13040 (N_13040,N_12789,N_12905);
or U13041 (N_13041,N_12807,N_12980);
nand U13042 (N_13042,N_12857,N_12940);
or U13043 (N_13043,N_12988,N_12884);
nor U13044 (N_13044,N_12872,N_12852);
nand U13045 (N_13045,N_12952,N_12762);
or U13046 (N_13046,N_12785,N_12804);
or U13047 (N_13047,N_12806,N_12763);
and U13048 (N_13048,N_12965,N_12987);
nand U13049 (N_13049,N_12895,N_12992);
xor U13050 (N_13050,N_12881,N_12850);
or U13051 (N_13051,N_12887,N_12898);
or U13052 (N_13052,N_12931,N_12938);
xor U13053 (N_13053,N_12877,N_12873);
nand U13054 (N_13054,N_12827,N_12760);
nor U13055 (N_13055,N_12860,N_12955);
or U13056 (N_13056,N_12795,N_12862);
nor U13057 (N_13057,N_12834,N_12919);
or U13058 (N_13058,N_12841,N_12983);
or U13059 (N_13059,N_12896,N_12882);
nand U13060 (N_13060,N_12808,N_12875);
xor U13061 (N_13061,N_12830,N_12843);
nand U13062 (N_13062,N_12797,N_12784);
xnor U13063 (N_13063,N_12993,N_12768);
and U13064 (N_13064,N_12751,N_12942);
xnor U13065 (N_13065,N_12933,N_12771);
xor U13066 (N_13066,N_12769,N_12774);
xor U13067 (N_13067,N_12901,N_12829);
nand U13068 (N_13068,N_12989,N_12773);
xnor U13069 (N_13069,N_12865,N_12984);
or U13070 (N_13070,N_12946,N_12802);
nor U13071 (N_13071,N_12831,N_12972);
nor U13072 (N_13072,N_12803,N_12967);
nand U13073 (N_13073,N_12923,N_12823);
nand U13074 (N_13074,N_12855,N_12925);
xor U13075 (N_13075,N_12978,N_12812);
and U13076 (N_13076,N_12876,N_12848);
and U13077 (N_13077,N_12950,N_12906);
and U13078 (N_13078,N_12765,N_12943);
nand U13079 (N_13079,N_12856,N_12836);
nor U13080 (N_13080,N_12837,N_12929);
or U13081 (N_13081,N_12786,N_12910);
nor U13082 (N_13082,N_12948,N_12818);
or U13083 (N_13083,N_12958,N_12963);
nor U13084 (N_13084,N_12995,N_12920);
and U13085 (N_13085,N_12981,N_12935);
or U13086 (N_13086,N_12944,N_12832);
xor U13087 (N_13087,N_12969,N_12866);
or U13088 (N_13088,N_12845,N_12759);
and U13089 (N_13089,N_12864,N_12956);
nand U13090 (N_13090,N_12930,N_12953);
and U13091 (N_13091,N_12815,N_12912);
nand U13092 (N_13092,N_12822,N_12894);
and U13093 (N_13093,N_12964,N_12994);
xor U13094 (N_13094,N_12915,N_12755);
or U13095 (N_13095,N_12799,N_12820);
nor U13096 (N_13096,N_12753,N_12922);
or U13097 (N_13097,N_12811,N_12985);
and U13098 (N_13098,N_12817,N_12885);
or U13099 (N_13099,N_12772,N_12833);
or U13100 (N_13100,N_12801,N_12916);
or U13101 (N_13101,N_12861,N_12991);
xor U13102 (N_13102,N_12970,N_12838);
and U13103 (N_13103,N_12800,N_12913);
or U13104 (N_13104,N_12766,N_12869);
xnor U13105 (N_13105,N_12790,N_12897);
nor U13106 (N_13106,N_12770,N_12757);
nand U13107 (N_13107,N_12927,N_12900);
and U13108 (N_13108,N_12893,N_12851);
or U13109 (N_13109,N_12961,N_12999);
or U13110 (N_13110,N_12758,N_12982);
xnor U13111 (N_13111,N_12977,N_12775);
nor U13112 (N_13112,N_12813,N_12971);
nor U13113 (N_13113,N_12936,N_12863);
xnor U13114 (N_13114,N_12779,N_12859);
nor U13115 (N_13115,N_12767,N_12754);
nor U13116 (N_13116,N_12973,N_12954);
or U13117 (N_13117,N_12918,N_12828);
nor U13118 (N_13118,N_12941,N_12826);
or U13119 (N_13119,N_12974,N_12874);
and U13120 (N_13120,N_12890,N_12798);
nand U13121 (N_13121,N_12814,N_12883);
xor U13122 (N_13122,N_12932,N_12899);
or U13123 (N_13123,N_12945,N_12928);
nor U13124 (N_13124,N_12886,N_12975);
xor U13125 (N_13125,N_12864,N_12779);
or U13126 (N_13126,N_12957,N_12803);
and U13127 (N_13127,N_12901,N_12825);
xnor U13128 (N_13128,N_12955,N_12750);
nor U13129 (N_13129,N_12816,N_12793);
and U13130 (N_13130,N_12795,N_12926);
nor U13131 (N_13131,N_12860,N_12852);
and U13132 (N_13132,N_12870,N_12890);
xor U13133 (N_13133,N_12959,N_12857);
nand U13134 (N_13134,N_12932,N_12875);
and U13135 (N_13135,N_12786,N_12880);
nand U13136 (N_13136,N_12836,N_12946);
nor U13137 (N_13137,N_12768,N_12976);
and U13138 (N_13138,N_12955,N_12775);
or U13139 (N_13139,N_12959,N_12834);
nor U13140 (N_13140,N_12958,N_12876);
nand U13141 (N_13141,N_12989,N_12984);
nor U13142 (N_13142,N_12823,N_12833);
and U13143 (N_13143,N_12963,N_12982);
or U13144 (N_13144,N_12813,N_12994);
and U13145 (N_13145,N_12970,N_12787);
or U13146 (N_13146,N_12812,N_12854);
xor U13147 (N_13147,N_12875,N_12820);
nor U13148 (N_13148,N_12833,N_12801);
nor U13149 (N_13149,N_12757,N_12762);
nand U13150 (N_13150,N_12778,N_12941);
nand U13151 (N_13151,N_12999,N_12804);
xnor U13152 (N_13152,N_12987,N_12837);
and U13153 (N_13153,N_12953,N_12762);
nand U13154 (N_13154,N_12767,N_12841);
nor U13155 (N_13155,N_12856,N_12958);
and U13156 (N_13156,N_12873,N_12762);
and U13157 (N_13157,N_12990,N_12813);
xor U13158 (N_13158,N_12794,N_12910);
nand U13159 (N_13159,N_12788,N_12849);
nand U13160 (N_13160,N_12800,N_12862);
nor U13161 (N_13161,N_12882,N_12932);
nor U13162 (N_13162,N_12951,N_12934);
nor U13163 (N_13163,N_12876,N_12870);
or U13164 (N_13164,N_12873,N_12781);
and U13165 (N_13165,N_12856,N_12940);
and U13166 (N_13166,N_12906,N_12799);
nand U13167 (N_13167,N_12882,N_12987);
or U13168 (N_13168,N_12862,N_12831);
nor U13169 (N_13169,N_12824,N_12924);
and U13170 (N_13170,N_12762,N_12978);
or U13171 (N_13171,N_12816,N_12788);
nor U13172 (N_13172,N_12918,N_12965);
nand U13173 (N_13173,N_12973,N_12828);
xnor U13174 (N_13174,N_12975,N_12931);
or U13175 (N_13175,N_12769,N_12785);
or U13176 (N_13176,N_12925,N_12760);
and U13177 (N_13177,N_12885,N_12873);
xor U13178 (N_13178,N_12983,N_12790);
or U13179 (N_13179,N_12818,N_12815);
or U13180 (N_13180,N_12809,N_12869);
nor U13181 (N_13181,N_12904,N_12959);
xnor U13182 (N_13182,N_12901,N_12926);
nand U13183 (N_13183,N_12778,N_12791);
nor U13184 (N_13184,N_12802,N_12968);
nor U13185 (N_13185,N_12861,N_12839);
or U13186 (N_13186,N_12977,N_12832);
xor U13187 (N_13187,N_12958,N_12805);
nor U13188 (N_13188,N_12894,N_12939);
xnor U13189 (N_13189,N_12882,N_12866);
nor U13190 (N_13190,N_12832,N_12804);
and U13191 (N_13191,N_12946,N_12760);
and U13192 (N_13192,N_12957,N_12868);
nor U13193 (N_13193,N_12886,N_12855);
xnor U13194 (N_13194,N_12781,N_12949);
nor U13195 (N_13195,N_12880,N_12932);
nor U13196 (N_13196,N_12954,N_12831);
nor U13197 (N_13197,N_12873,N_12798);
nand U13198 (N_13198,N_12931,N_12936);
nor U13199 (N_13199,N_12940,N_12800);
nor U13200 (N_13200,N_12804,N_12759);
xnor U13201 (N_13201,N_12784,N_12849);
or U13202 (N_13202,N_12856,N_12793);
nand U13203 (N_13203,N_12804,N_12892);
xnor U13204 (N_13204,N_12825,N_12766);
or U13205 (N_13205,N_12966,N_12774);
nor U13206 (N_13206,N_12794,N_12956);
xor U13207 (N_13207,N_12909,N_12856);
xor U13208 (N_13208,N_12940,N_12989);
or U13209 (N_13209,N_12767,N_12915);
nand U13210 (N_13210,N_12872,N_12931);
nand U13211 (N_13211,N_12914,N_12751);
nor U13212 (N_13212,N_12758,N_12963);
or U13213 (N_13213,N_12996,N_12871);
or U13214 (N_13214,N_12805,N_12909);
nand U13215 (N_13215,N_12813,N_12916);
nand U13216 (N_13216,N_12920,N_12974);
nand U13217 (N_13217,N_12949,N_12860);
and U13218 (N_13218,N_12758,N_12861);
nor U13219 (N_13219,N_12857,N_12964);
xnor U13220 (N_13220,N_12761,N_12997);
xor U13221 (N_13221,N_12964,N_12943);
or U13222 (N_13222,N_12828,N_12771);
nor U13223 (N_13223,N_12872,N_12867);
and U13224 (N_13224,N_12858,N_12876);
xor U13225 (N_13225,N_12927,N_12862);
and U13226 (N_13226,N_12963,N_12857);
xnor U13227 (N_13227,N_12928,N_12782);
xor U13228 (N_13228,N_12987,N_12905);
or U13229 (N_13229,N_12995,N_12981);
nor U13230 (N_13230,N_12878,N_12779);
and U13231 (N_13231,N_12776,N_12760);
nor U13232 (N_13232,N_12998,N_12974);
nand U13233 (N_13233,N_12760,N_12929);
xnor U13234 (N_13234,N_12954,N_12852);
xor U13235 (N_13235,N_12935,N_12919);
nand U13236 (N_13236,N_12952,N_12751);
xor U13237 (N_13237,N_12958,N_12801);
and U13238 (N_13238,N_12840,N_12883);
nor U13239 (N_13239,N_12866,N_12750);
nor U13240 (N_13240,N_12989,N_12866);
nand U13241 (N_13241,N_12772,N_12837);
nor U13242 (N_13242,N_12992,N_12877);
nor U13243 (N_13243,N_12949,N_12931);
xor U13244 (N_13244,N_12893,N_12781);
xnor U13245 (N_13245,N_12787,N_12768);
or U13246 (N_13246,N_12796,N_12885);
or U13247 (N_13247,N_12772,N_12898);
nand U13248 (N_13248,N_12836,N_12892);
and U13249 (N_13249,N_12863,N_12902);
nand U13250 (N_13250,N_13096,N_13205);
or U13251 (N_13251,N_13245,N_13231);
nand U13252 (N_13252,N_13058,N_13072);
and U13253 (N_13253,N_13005,N_13095);
or U13254 (N_13254,N_13022,N_13079);
or U13255 (N_13255,N_13093,N_13221);
nor U13256 (N_13256,N_13220,N_13047);
nand U13257 (N_13257,N_13163,N_13004);
nand U13258 (N_13258,N_13199,N_13131);
or U13259 (N_13259,N_13158,N_13101);
nand U13260 (N_13260,N_13025,N_13232);
and U13261 (N_13261,N_13204,N_13110);
or U13262 (N_13262,N_13184,N_13238);
or U13263 (N_13263,N_13170,N_13020);
or U13264 (N_13264,N_13078,N_13111);
or U13265 (N_13265,N_13212,N_13210);
and U13266 (N_13266,N_13179,N_13227);
nor U13267 (N_13267,N_13139,N_13133);
or U13268 (N_13268,N_13087,N_13026);
nor U13269 (N_13269,N_13146,N_13161);
nor U13270 (N_13270,N_13243,N_13070);
nand U13271 (N_13271,N_13136,N_13211);
or U13272 (N_13272,N_13157,N_13197);
nand U13273 (N_13273,N_13202,N_13102);
and U13274 (N_13274,N_13048,N_13040);
nor U13275 (N_13275,N_13099,N_13010);
nand U13276 (N_13276,N_13144,N_13105);
xnor U13277 (N_13277,N_13084,N_13107);
xnor U13278 (N_13278,N_13246,N_13066);
or U13279 (N_13279,N_13014,N_13222);
or U13280 (N_13280,N_13094,N_13226);
xnor U13281 (N_13281,N_13098,N_13162);
xnor U13282 (N_13282,N_13086,N_13115);
xnor U13283 (N_13283,N_13153,N_13037);
nor U13284 (N_13284,N_13074,N_13008);
xnor U13285 (N_13285,N_13062,N_13035);
xor U13286 (N_13286,N_13126,N_13082);
nor U13287 (N_13287,N_13104,N_13130);
nor U13288 (N_13288,N_13174,N_13239);
nand U13289 (N_13289,N_13063,N_13194);
nand U13290 (N_13290,N_13106,N_13241);
and U13291 (N_13291,N_13043,N_13006);
or U13292 (N_13292,N_13100,N_13120);
and U13293 (N_13293,N_13019,N_13223);
or U13294 (N_13294,N_13219,N_13012);
xnor U13295 (N_13295,N_13032,N_13121);
or U13296 (N_13296,N_13039,N_13054);
and U13297 (N_13297,N_13209,N_13189);
nand U13298 (N_13298,N_13206,N_13112);
or U13299 (N_13299,N_13148,N_13081);
and U13300 (N_13300,N_13135,N_13141);
nor U13301 (N_13301,N_13090,N_13059);
and U13302 (N_13302,N_13108,N_13237);
nor U13303 (N_13303,N_13214,N_13218);
xor U13304 (N_13304,N_13142,N_13000);
nand U13305 (N_13305,N_13233,N_13200);
xor U13306 (N_13306,N_13071,N_13134);
nor U13307 (N_13307,N_13064,N_13155);
nand U13308 (N_13308,N_13242,N_13244);
xor U13309 (N_13309,N_13143,N_13127);
and U13310 (N_13310,N_13196,N_13080);
or U13311 (N_13311,N_13177,N_13016);
and U13312 (N_13312,N_13113,N_13181);
or U13313 (N_13313,N_13169,N_13151);
xnor U13314 (N_13314,N_13249,N_13156);
nor U13315 (N_13315,N_13191,N_13027);
nor U13316 (N_13316,N_13088,N_13201);
and U13317 (N_13317,N_13217,N_13234);
or U13318 (N_13318,N_13018,N_13017);
and U13319 (N_13319,N_13092,N_13152);
or U13320 (N_13320,N_13248,N_13188);
nand U13321 (N_13321,N_13216,N_13122);
xor U13322 (N_13322,N_13077,N_13075);
xnor U13323 (N_13323,N_13045,N_13109);
xnor U13324 (N_13324,N_13068,N_13028);
nor U13325 (N_13325,N_13215,N_13235);
or U13326 (N_13326,N_13085,N_13147);
or U13327 (N_13327,N_13103,N_13138);
nor U13328 (N_13328,N_13060,N_13076);
nand U13329 (N_13329,N_13007,N_13159);
nor U13330 (N_13330,N_13023,N_13050);
nor U13331 (N_13331,N_13145,N_13228);
and U13332 (N_13332,N_13224,N_13240);
nand U13333 (N_13333,N_13117,N_13044);
nor U13334 (N_13334,N_13187,N_13061);
nand U13335 (N_13335,N_13089,N_13097);
nor U13336 (N_13336,N_13198,N_13069);
nor U13337 (N_13337,N_13229,N_13067);
nor U13338 (N_13338,N_13021,N_13185);
nand U13339 (N_13339,N_13015,N_13013);
nand U13340 (N_13340,N_13150,N_13168);
and U13341 (N_13341,N_13029,N_13046);
and U13342 (N_13342,N_13171,N_13034);
and U13343 (N_13343,N_13057,N_13230);
or U13344 (N_13344,N_13175,N_13213);
xor U13345 (N_13345,N_13172,N_13207);
nand U13346 (N_13346,N_13119,N_13116);
or U13347 (N_13347,N_13052,N_13195);
or U13348 (N_13348,N_13190,N_13160);
nor U13349 (N_13349,N_13003,N_13149);
nand U13350 (N_13350,N_13049,N_13114);
or U13351 (N_13351,N_13173,N_13036);
nand U13352 (N_13352,N_13176,N_13051);
or U13353 (N_13353,N_13002,N_13073);
nor U13354 (N_13354,N_13041,N_13154);
nor U13355 (N_13355,N_13236,N_13033);
and U13356 (N_13356,N_13164,N_13192);
nand U13357 (N_13357,N_13186,N_13208);
and U13358 (N_13358,N_13166,N_13123);
nand U13359 (N_13359,N_13193,N_13183);
nand U13360 (N_13360,N_13165,N_13225);
xor U13361 (N_13361,N_13247,N_13024);
nor U13362 (N_13362,N_13001,N_13118);
nor U13363 (N_13363,N_13031,N_13180);
nand U13364 (N_13364,N_13203,N_13065);
and U13365 (N_13365,N_13030,N_13140);
or U13366 (N_13366,N_13056,N_13091);
and U13367 (N_13367,N_13128,N_13129);
nor U13368 (N_13368,N_13132,N_13124);
xor U13369 (N_13369,N_13167,N_13178);
nand U13370 (N_13370,N_13137,N_13055);
or U13371 (N_13371,N_13038,N_13009);
and U13372 (N_13372,N_13125,N_13083);
nand U13373 (N_13373,N_13182,N_13053);
nor U13374 (N_13374,N_13042,N_13011);
and U13375 (N_13375,N_13100,N_13090);
xnor U13376 (N_13376,N_13012,N_13153);
and U13377 (N_13377,N_13097,N_13016);
and U13378 (N_13378,N_13058,N_13041);
or U13379 (N_13379,N_13173,N_13182);
or U13380 (N_13380,N_13214,N_13007);
nand U13381 (N_13381,N_13185,N_13206);
nor U13382 (N_13382,N_13005,N_13064);
nand U13383 (N_13383,N_13242,N_13106);
nor U13384 (N_13384,N_13224,N_13021);
nand U13385 (N_13385,N_13197,N_13062);
xor U13386 (N_13386,N_13049,N_13023);
or U13387 (N_13387,N_13076,N_13089);
nand U13388 (N_13388,N_13104,N_13008);
and U13389 (N_13389,N_13040,N_13131);
and U13390 (N_13390,N_13061,N_13162);
xor U13391 (N_13391,N_13086,N_13183);
nor U13392 (N_13392,N_13103,N_13071);
xor U13393 (N_13393,N_13180,N_13033);
nand U13394 (N_13394,N_13032,N_13243);
nand U13395 (N_13395,N_13217,N_13218);
or U13396 (N_13396,N_13180,N_13236);
xor U13397 (N_13397,N_13240,N_13246);
nor U13398 (N_13398,N_13240,N_13223);
and U13399 (N_13399,N_13239,N_13185);
and U13400 (N_13400,N_13213,N_13169);
nand U13401 (N_13401,N_13127,N_13196);
xor U13402 (N_13402,N_13240,N_13168);
or U13403 (N_13403,N_13017,N_13205);
and U13404 (N_13404,N_13140,N_13054);
and U13405 (N_13405,N_13119,N_13120);
xnor U13406 (N_13406,N_13210,N_13128);
xor U13407 (N_13407,N_13178,N_13195);
and U13408 (N_13408,N_13084,N_13060);
and U13409 (N_13409,N_13155,N_13166);
and U13410 (N_13410,N_13065,N_13052);
or U13411 (N_13411,N_13032,N_13073);
nand U13412 (N_13412,N_13010,N_13089);
nor U13413 (N_13413,N_13057,N_13221);
nand U13414 (N_13414,N_13155,N_13050);
nand U13415 (N_13415,N_13235,N_13232);
and U13416 (N_13416,N_13188,N_13226);
xor U13417 (N_13417,N_13215,N_13244);
nand U13418 (N_13418,N_13217,N_13022);
and U13419 (N_13419,N_13050,N_13137);
nor U13420 (N_13420,N_13190,N_13104);
xor U13421 (N_13421,N_13044,N_13065);
or U13422 (N_13422,N_13241,N_13041);
or U13423 (N_13423,N_13043,N_13129);
xnor U13424 (N_13424,N_13194,N_13145);
and U13425 (N_13425,N_13198,N_13162);
xnor U13426 (N_13426,N_13225,N_13021);
and U13427 (N_13427,N_13175,N_13152);
xor U13428 (N_13428,N_13142,N_13154);
and U13429 (N_13429,N_13072,N_13165);
nor U13430 (N_13430,N_13060,N_13019);
xor U13431 (N_13431,N_13025,N_13170);
nor U13432 (N_13432,N_13194,N_13090);
or U13433 (N_13433,N_13161,N_13086);
nor U13434 (N_13434,N_13087,N_13221);
nand U13435 (N_13435,N_13233,N_13124);
or U13436 (N_13436,N_13155,N_13034);
nand U13437 (N_13437,N_13043,N_13133);
xor U13438 (N_13438,N_13074,N_13153);
nand U13439 (N_13439,N_13047,N_13051);
nand U13440 (N_13440,N_13216,N_13025);
xnor U13441 (N_13441,N_13132,N_13078);
or U13442 (N_13442,N_13143,N_13232);
nor U13443 (N_13443,N_13000,N_13198);
and U13444 (N_13444,N_13039,N_13056);
or U13445 (N_13445,N_13228,N_13217);
nand U13446 (N_13446,N_13037,N_13246);
xor U13447 (N_13447,N_13096,N_13152);
xnor U13448 (N_13448,N_13178,N_13050);
nor U13449 (N_13449,N_13243,N_13136);
xor U13450 (N_13450,N_13221,N_13208);
or U13451 (N_13451,N_13101,N_13225);
and U13452 (N_13452,N_13224,N_13047);
xor U13453 (N_13453,N_13053,N_13067);
nand U13454 (N_13454,N_13182,N_13242);
and U13455 (N_13455,N_13055,N_13089);
xor U13456 (N_13456,N_13067,N_13135);
nor U13457 (N_13457,N_13244,N_13153);
and U13458 (N_13458,N_13168,N_13016);
xor U13459 (N_13459,N_13112,N_13229);
xor U13460 (N_13460,N_13131,N_13125);
nor U13461 (N_13461,N_13111,N_13105);
nor U13462 (N_13462,N_13014,N_13210);
nor U13463 (N_13463,N_13118,N_13017);
xor U13464 (N_13464,N_13165,N_13142);
nor U13465 (N_13465,N_13000,N_13212);
xnor U13466 (N_13466,N_13053,N_13168);
xnor U13467 (N_13467,N_13016,N_13094);
xor U13468 (N_13468,N_13072,N_13173);
or U13469 (N_13469,N_13122,N_13113);
nand U13470 (N_13470,N_13013,N_13151);
nor U13471 (N_13471,N_13073,N_13213);
nand U13472 (N_13472,N_13163,N_13043);
or U13473 (N_13473,N_13127,N_13185);
nand U13474 (N_13474,N_13010,N_13130);
and U13475 (N_13475,N_13217,N_13131);
nand U13476 (N_13476,N_13086,N_13095);
xnor U13477 (N_13477,N_13245,N_13084);
or U13478 (N_13478,N_13071,N_13079);
nand U13479 (N_13479,N_13086,N_13034);
nor U13480 (N_13480,N_13000,N_13170);
nor U13481 (N_13481,N_13244,N_13078);
and U13482 (N_13482,N_13135,N_13205);
nor U13483 (N_13483,N_13036,N_13236);
nor U13484 (N_13484,N_13228,N_13027);
xor U13485 (N_13485,N_13203,N_13084);
xnor U13486 (N_13486,N_13045,N_13040);
nor U13487 (N_13487,N_13232,N_13021);
nand U13488 (N_13488,N_13046,N_13213);
xor U13489 (N_13489,N_13245,N_13163);
and U13490 (N_13490,N_13007,N_13230);
and U13491 (N_13491,N_13178,N_13125);
xnor U13492 (N_13492,N_13181,N_13246);
xor U13493 (N_13493,N_13105,N_13136);
xor U13494 (N_13494,N_13189,N_13195);
nor U13495 (N_13495,N_13113,N_13224);
nand U13496 (N_13496,N_13061,N_13206);
nor U13497 (N_13497,N_13065,N_13213);
nand U13498 (N_13498,N_13169,N_13070);
and U13499 (N_13499,N_13150,N_13247);
or U13500 (N_13500,N_13329,N_13287);
or U13501 (N_13501,N_13301,N_13413);
nand U13502 (N_13502,N_13345,N_13321);
nand U13503 (N_13503,N_13350,N_13403);
and U13504 (N_13504,N_13470,N_13351);
xnor U13505 (N_13505,N_13475,N_13252);
and U13506 (N_13506,N_13455,N_13383);
nor U13507 (N_13507,N_13299,N_13333);
xnor U13508 (N_13508,N_13311,N_13479);
xor U13509 (N_13509,N_13493,N_13378);
nor U13510 (N_13510,N_13336,N_13457);
xnor U13511 (N_13511,N_13354,N_13335);
and U13512 (N_13512,N_13273,N_13255);
nor U13513 (N_13513,N_13466,N_13411);
xor U13514 (N_13514,N_13290,N_13313);
xnor U13515 (N_13515,N_13414,N_13469);
or U13516 (N_13516,N_13492,N_13305);
and U13517 (N_13517,N_13284,N_13282);
xor U13518 (N_13518,N_13300,N_13484);
nor U13519 (N_13519,N_13454,N_13490);
and U13520 (N_13520,N_13265,N_13314);
nor U13521 (N_13521,N_13434,N_13286);
nand U13522 (N_13522,N_13369,N_13291);
or U13523 (N_13523,N_13447,N_13362);
nor U13524 (N_13524,N_13306,N_13302);
xnor U13525 (N_13525,N_13483,N_13464);
xnor U13526 (N_13526,N_13281,N_13393);
nand U13527 (N_13527,N_13485,N_13331);
xnor U13528 (N_13528,N_13380,N_13285);
or U13529 (N_13529,N_13275,N_13296);
nor U13530 (N_13530,N_13445,N_13416);
or U13531 (N_13531,N_13385,N_13297);
nor U13532 (N_13532,N_13423,N_13478);
nor U13533 (N_13533,N_13330,N_13259);
or U13534 (N_13534,N_13417,N_13359);
xnor U13535 (N_13535,N_13352,N_13420);
and U13536 (N_13536,N_13357,N_13332);
and U13537 (N_13537,N_13394,N_13461);
xor U13538 (N_13538,N_13446,N_13381);
nand U13539 (N_13539,N_13459,N_13495);
nand U13540 (N_13540,N_13346,N_13316);
xnor U13541 (N_13541,N_13427,N_13395);
xor U13542 (N_13542,N_13268,N_13327);
xnor U13543 (N_13543,N_13408,N_13410);
nand U13544 (N_13544,N_13384,N_13367);
and U13545 (N_13545,N_13298,N_13254);
and U13546 (N_13546,N_13486,N_13477);
nand U13547 (N_13547,N_13437,N_13386);
xnor U13548 (N_13548,N_13365,N_13375);
and U13549 (N_13549,N_13338,N_13419);
nor U13550 (N_13550,N_13438,N_13366);
nor U13551 (N_13551,N_13371,N_13409);
or U13552 (N_13552,N_13401,N_13278);
or U13553 (N_13553,N_13473,N_13439);
and U13554 (N_13554,N_13435,N_13271);
nand U13555 (N_13555,N_13382,N_13289);
or U13556 (N_13556,N_13463,N_13356);
and U13557 (N_13557,N_13295,N_13266);
and U13558 (N_13558,N_13426,N_13431);
xor U13559 (N_13559,N_13342,N_13355);
nor U13560 (N_13560,N_13322,N_13280);
nand U13561 (N_13561,N_13480,N_13468);
and U13562 (N_13562,N_13253,N_13277);
nand U13563 (N_13563,N_13433,N_13308);
nand U13564 (N_13564,N_13353,N_13407);
xor U13565 (N_13565,N_13274,N_13474);
nor U13566 (N_13566,N_13261,N_13467);
nor U13567 (N_13567,N_13312,N_13405);
nor U13568 (N_13568,N_13272,N_13317);
nand U13569 (N_13569,N_13347,N_13462);
or U13570 (N_13570,N_13499,N_13488);
xor U13571 (N_13571,N_13315,N_13458);
nand U13572 (N_13572,N_13448,N_13397);
or U13573 (N_13573,N_13497,N_13418);
xor U13574 (N_13574,N_13341,N_13404);
xnor U13575 (N_13575,N_13422,N_13349);
nand U13576 (N_13576,N_13482,N_13443);
nor U13577 (N_13577,N_13376,N_13340);
nor U13578 (N_13578,N_13440,N_13264);
xor U13579 (N_13579,N_13251,N_13372);
and U13580 (N_13580,N_13487,N_13326);
nand U13581 (N_13581,N_13460,N_13262);
xnor U13582 (N_13582,N_13391,N_13343);
and U13583 (N_13583,N_13368,N_13364);
nor U13584 (N_13584,N_13304,N_13392);
xor U13585 (N_13585,N_13318,N_13276);
nor U13586 (N_13586,N_13258,N_13450);
nand U13587 (N_13587,N_13279,N_13406);
and U13588 (N_13588,N_13430,N_13292);
nand U13589 (N_13589,N_13396,N_13432);
nor U13590 (N_13590,N_13379,N_13476);
nand U13591 (N_13591,N_13402,N_13400);
nor U13592 (N_13592,N_13449,N_13373);
xnor U13593 (N_13593,N_13325,N_13303);
or U13594 (N_13594,N_13456,N_13494);
xnor U13595 (N_13595,N_13337,N_13421);
nand U13596 (N_13596,N_13307,N_13472);
and U13597 (N_13597,N_13328,N_13309);
or U13598 (N_13598,N_13260,N_13377);
xnor U13599 (N_13599,N_13334,N_13398);
or U13600 (N_13600,N_13441,N_13471);
and U13601 (N_13601,N_13358,N_13263);
xnor U13602 (N_13602,N_13412,N_13361);
or U13603 (N_13603,N_13390,N_13348);
xor U13604 (N_13604,N_13360,N_13250);
xor U13605 (N_13605,N_13288,N_13429);
and U13606 (N_13606,N_13451,N_13256);
nor U13607 (N_13607,N_13363,N_13269);
and U13608 (N_13608,N_13270,N_13320);
nor U13609 (N_13609,N_13424,N_13453);
and U13610 (N_13610,N_13267,N_13481);
nor U13611 (N_13611,N_13452,N_13489);
xor U13612 (N_13612,N_13387,N_13323);
nor U13613 (N_13613,N_13324,N_13491);
and U13614 (N_13614,N_13293,N_13294);
xor U13615 (N_13615,N_13310,N_13428);
and U13616 (N_13616,N_13339,N_13496);
or U13617 (N_13617,N_13283,N_13388);
and U13618 (N_13618,N_13442,N_13425);
and U13619 (N_13619,N_13370,N_13498);
xor U13620 (N_13620,N_13257,N_13374);
and U13621 (N_13621,N_13399,N_13319);
nand U13622 (N_13622,N_13444,N_13465);
nand U13623 (N_13623,N_13415,N_13344);
nand U13624 (N_13624,N_13389,N_13436);
and U13625 (N_13625,N_13365,N_13288);
xor U13626 (N_13626,N_13314,N_13254);
or U13627 (N_13627,N_13387,N_13394);
nand U13628 (N_13628,N_13280,N_13449);
nand U13629 (N_13629,N_13409,N_13454);
nor U13630 (N_13630,N_13465,N_13454);
and U13631 (N_13631,N_13390,N_13439);
or U13632 (N_13632,N_13473,N_13418);
and U13633 (N_13633,N_13429,N_13278);
nor U13634 (N_13634,N_13257,N_13459);
nor U13635 (N_13635,N_13480,N_13487);
nand U13636 (N_13636,N_13300,N_13365);
nor U13637 (N_13637,N_13304,N_13419);
nand U13638 (N_13638,N_13406,N_13353);
nand U13639 (N_13639,N_13268,N_13415);
nor U13640 (N_13640,N_13347,N_13476);
and U13641 (N_13641,N_13494,N_13484);
nand U13642 (N_13642,N_13408,N_13412);
nand U13643 (N_13643,N_13442,N_13381);
and U13644 (N_13644,N_13483,N_13478);
or U13645 (N_13645,N_13336,N_13308);
or U13646 (N_13646,N_13426,N_13381);
and U13647 (N_13647,N_13290,N_13333);
and U13648 (N_13648,N_13295,N_13353);
or U13649 (N_13649,N_13254,N_13353);
nand U13650 (N_13650,N_13489,N_13312);
nand U13651 (N_13651,N_13287,N_13259);
nor U13652 (N_13652,N_13488,N_13474);
nor U13653 (N_13653,N_13417,N_13416);
and U13654 (N_13654,N_13444,N_13433);
nor U13655 (N_13655,N_13416,N_13449);
nor U13656 (N_13656,N_13307,N_13450);
or U13657 (N_13657,N_13412,N_13312);
xnor U13658 (N_13658,N_13485,N_13364);
nand U13659 (N_13659,N_13496,N_13419);
xnor U13660 (N_13660,N_13498,N_13406);
or U13661 (N_13661,N_13376,N_13489);
nand U13662 (N_13662,N_13265,N_13378);
or U13663 (N_13663,N_13340,N_13390);
and U13664 (N_13664,N_13371,N_13472);
nand U13665 (N_13665,N_13335,N_13282);
and U13666 (N_13666,N_13377,N_13464);
nand U13667 (N_13667,N_13289,N_13342);
xnor U13668 (N_13668,N_13292,N_13320);
nand U13669 (N_13669,N_13253,N_13317);
nand U13670 (N_13670,N_13322,N_13347);
nand U13671 (N_13671,N_13410,N_13441);
nand U13672 (N_13672,N_13410,N_13280);
nand U13673 (N_13673,N_13279,N_13381);
nand U13674 (N_13674,N_13449,N_13288);
and U13675 (N_13675,N_13315,N_13480);
xor U13676 (N_13676,N_13452,N_13407);
xnor U13677 (N_13677,N_13252,N_13491);
or U13678 (N_13678,N_13328,N_13315);
nor U13679 (N_13679,N_13485,N_13313);
nand U13680 (N_13680,N_13441,N_13275);
nor U13681 (N_13681,N_13357,N_13276);
xor U13682 (N_13682,N_13493,N_13457);
nor U13683 (N_13683,N_13382,N_13413);
nand U13684 (N_13684,N_13295,N_13364);
xor U13685 (N_13685,N_13303,N_13283);
xnor U13686 (N_13686,N_13497,N_13277);
or U13687 (N_13687,N_13495,N_13350);
or U13688 (N_13688,N_13492,N_13444);
xnor U13689 (N_13689,N_13321,N_13398);
nand U13690 (N_13690,N_13490,N_13300);
nor U13691 (N_13691,N_13303,N_13390);
or U13692 (N_13692,N_13478,N_13451);
xnor U13693 (N_13693,N_13322,N_13420);
nor U13694 (N_13694,N_13420,N_13267);
xnor U13695 (N_13695,N_13390,N_13345);
nor U13696 (N_13696,N_13306,N_13466);
nor U13697 (N_13697,N_13286,N_13273);
nand U13698 (N_13698,N_13265,N_13441);
nand U13699 (N_13699,N_13355,N_13424);
and U13700 (N_13700,N_13376,N_13394);
xnor U13701 (N_13701,N_13265,N_13261);
and U13702 (N_13702,N_13412,N_13347);
and U13703 (N_13703,N_13312,N_13497);
nand U13704 (N_13704,N_13406,N_13458);
nand U13705 (N_13705,N_13377,N_13356);
and U13706 (N_13706,N_13417,N_13492);
and U13707 (N_13707,N_13484,N_13254);
nor U13708 (N_13708,N_13494,N_13363);
and U13709 (N_13709,N_13464,N_13436);
xnor U13710 (N_13710,N_13478,N_13297);
nor U13711 (N_13711,N_13253,N_13450);
nor U13712 (N_13712,N_13269,N_13447);
xnor U13713 (N_13713,N_13260,N_13401);
or U13714 (N_13714,N_13427,N_13408);
and U13715 (N_13715,N_13415,N_13260);
and U13716 (N_13716,N_13475,N_13495);
xnor U13717 (N_13717,N_13290,N_13393);
nand U13718 (N_13718,N_13440,N_13360);
nor U13719 (N_13719,N_13304,N_13322);
nand U13720 (N_13720,N_13333,N_13475);
or U13721 (N_13721,N_13304,N_13481);
nand U13722 (N_13722,N_13400,N_13309);
xnor U13723 (N_13723,N_13276,N_13352);
nand U13724 (N_13724,N_13376,N_13435);
nand U13725 (N_13725,N_13271,N_13400);
xnor U13726 (N_13726,N_13341,N_13448);
and U13727 (N_13727,N_13295,N_13451);
and U13728 (N_13728,N_13326,N_13493);
nor U13729 (N_13729,N_13368,N_13452);
or U13730 (N_13730,N_13335,N_13276);
or U13731 (N_13731,N_13407,N_13369);
nor U13732 (N_13732,N_13309,N_13343);
or U13733 (N_13733,N_13457,N_13361);
and U13734 (N_13734,N_13304,N_13458);
xnor U13735 (N_13735,N_13380,N_13260);
xor U13736 (N_13736,N_13377,N_13467);
nand U13737 (N_13737,N_13328,N_13281);
and U13738 (N_13738,N_13460,N_13437);
and U13739 (N_13739,N_13275,N_13339);
nor U13740 (N_13740,N_13457,N_13317);
xor U13741 (N_13741,N_13400,N_13274);
or U13742 (N_13742,N_13380,N_13476);
or U13743 (N_13743,N_13473,N_13317);
xor U13744 (N_13744,N_13300,N_13451);
nand U13745 (N_13745,N_13434,N_13364);
and U13746 (N_13746,N_13390,N_13433);
or U13747 (N_13747,N_13411,N_13347);
xor U13748 (N_13748,N_13412,N_13317);
xor U13749 (N_13749,N_13425,N_13457);
xnor U13750 (N_13750,N_13587,N_13700);
and U13751 (N_13751,N_13517,N_13569);
nor U13752 (N_13752,N_13733,N_13683);
nand U13753 (N_13753,N_13542,N_13556);
and U13754 (N_13754,N_13502,N_13548);
nor U13755 (N_13755,N_13592,N_13703);
nor U13756 (N_13756,N_13748,N_13538);
nor U13757 (N_13757,N_13554,N_13680);
nor U13758 (N_13758,N_13627,N_13581);
or U13759 (N_13759,N_13615,N_13524);
xor U13760 (N_13760,N_13543,N_13686);
xor U13761 (N_13761,N_13726,N_13589);
nand U13762 (N_13762,N_13614,N_13642);
and U13763 (N_13763,N_13591,N_13722);
and U13764 (N_13764,N_13622,N_13578);
or U13765 (N_13765,N_13718,N_13712);
and U13766 (N_13766,N_13738,N_13546);
nand U13767 (N_13767,N_13661,N_13590);
or U13768 (N_13768,N_13678,N_13744);
xor U13769 (N_13769,N_13646,N_13629);
nor U13770 (N_13770,N_13709,N_13514);
nor U13771 (N_13771,N_13663,N_13645);
nand U13772 (N_13772,N_13525,N_13552);
and U13773 (N_13773,N_13582,N_13594);
nand U13774 (N_13774,N_13567,N_13721);
xor U13775 (N_13775,N_13739,N_13530);
xnor U13776 (N_13776,N_13638,N_13707);
and U13777 (N_13777,N_13656,N_13536);
and U13778 (N_13778,N_13518,N_13605);
or U13779 (N_13779,N_13557,N_13508);
and U13780 (N_13780,N_13540,N_13708);
and U13781 (N_13781,N_13521,N_13580);
or U13782 (N_13782,N_13544,N_13681);
nor U13783 (N_13783,N_13644,N_13549);
nor U13784 (N_13784,N_13639,N_13746);
nand U13785 (N_13785,N_13631,N_13635);
nand U13786 (N_13786,N_13720,N_13640);
and U13787 (N_13787,N_13724,N_13526);
or U13788 (N_13788,N_13507,N_13672);
nor U13789 (N_13789,N_13611,N_13562);
and U13790 (N_13790,N_13692,N_13725);
nand U13791 (N_13791,N_13673,N_13513);
and U13792 (N_13792,N_13694,N_13565);
xor U13793 (N_13793,N_13714,N_13547);
and U13794 (N_13794,N_13685,N_13519);
xor U13795 (N_13795,N_13667,N_13660);
nand U13796 (N_13796,N_13583,N_13597);
nor U13797 (N_13797,N_13595,N_13734);
or U13798 (N_13798,N_13603,N_13558);
and U13799 (N_13799,N_13649,N_13743);
nand U13800 (N_13800,N_13702,N_13527);
and U13801 (N_13801,N_13529,N_13636);
and U13802 (N_13802,N_13600,N_13500);
or U13803 (N_13803,N_13617,N_13577);
nand U13804 (N_13804,N_13684,N_13670);
xor U13805 (N_13805,N_13728,N_13699);
and U13806 (N_13806,N_13659,N_13564);
and U13807 (N_13807,N_13599,N_13607);
xor U13808 (N_13808,N_13576,N_13501);
and U13809 (N_13809,N_13588,N_13658);
xnor U13810 (N_13810,N_13559,N_13665);
nand U13811 (N_13811,N_13510,N_13669);
nand U13812 (N_13812,N_13747,N_13641);
xnor U13813 (N_13813,N_13650,N_13676);
nor U13814 (N_13814,N_13719,N_13652);
or U13815 (N_13815,N_13677,N_13624);
and U13816 (N_13816,N_13654,N_13691);
nand U13817 (N_13817,N_13553,N_13632);
and U13818 (N_13818,N_13533,N_13602);
and U13819 (N_13819,N_13742,N_13723);
nor U13820 (N_13820,N_13740,N_13705);
or U13821 (N_13821,N_13571,N_13522);
nor U13822 (N_13822,N_13647,N_13633);
xor U13823 (N_13823,N_13630,N_13745);
or U13824 (N_13824,N_13610,N_13623);
and U13825 (N_13825,N_13651,N_13563);
xor U13826 (N_13826,N_13637,N_13609);
and U13827 (N_13827,N_13717,N_13568);
and U13828 (N_13828,N_13619,N_13666);
nor U13829 (N_13829,N_13706,N_13545);
xnor U13830 (N_13830,N_13573,N_13596);
nand U13831 (N_13831,N_13698,N_13730);
nor U13832 (N_13832,N_13523,N_13749);
or U13833 (N_13833,N_13731,N_13537);
or U13834 (N_13834,N_13535,N_13593);
xnor U13835 (N_13835,N_13531,N_13503);
xnor U13836 (N_13836,N_13675,N_13628);
nor U13837 (N_13837,N_13566,N_13570);
nor U13838 (N_13838,N_13606,N_13693);
nor U13839 (N_13839,N_13621,N_13732);
and U13840 (N_13840,N_13511,N_13575);
or U13841 (N_13841,N_13579,N_13697);
and U13842 (N_13842,N_13584,N_13539);
and U13843 (N_13843,N_13551,N_13668);
and U13844 (N_13844,N_13689,N_13608);
nor U13845 (N_13845,N_13679,N_13505);
xnor U13846 (N_13846,N_13572,N_13648);
or U13847 (N_13847,N_13601,N_13710);
and U13848 (N_13848,N_13506,N_13613);
nor U13849 (N_13849,N_13515,N_13520);
xor U13850 (N_13850,N_13713,N_13715);
xor U13851 (N_13851,N_13664,N_13737);
xnor U13852 (N_13852,N_13727,N_13682);
nor U13853 (N_13853,N_13585,N_13687);
nor U13854 (N_13854,N_13512,N_13671);
or U13855 (N_13855,N_13704,N_13532);
and U13856 (N_13856,N_13618,N_13662);
and U13857 (N_13857,N_13695,N_13574);
nand U13858 (N_13858,N_13674,N_13729);
or U13859 (N_13859,N_13716,N_13643);
or U13860 (N_13860,N_13560,N_13528);
nor U13861 (N_13861,N_13711,N_13541);
or U13862 (N_13862,N_13616,N_13653);
and U13863 (N_13863,N_13735,N_13696);
xnor U13864 (N_13864,N_13634,N_13586);
and U13865 (N_13865,N_13620,N_13688);
or U13866 (N_13866,N_13555,N_13550);
nor U13867 (N_13867,N_13657,N_13604);
xor U13868 (N_13868,N_13741,N_13626);
and U13869 (N_13869,N_13516,N_13561);
nor U13870 (N_13870,N_13598,N_13504);
xor U13871 (N_13871,N_13534,N_13655);
xor U13872 (N_13872,N_13509,N_13612);
nor U13873 (N_13873,N_13701,N_13625);
nand U13874 (N_13874,N_13690,N_13736);
or U13875 (N_13875,N_13550,N_13618);
xor U13876 (N_13876,N_13747,N_13699);
nand U13877 (N_13877,N_13576,N_13645);
nand U13878 (N_13878,N_13517,N_13573);
or U13879 (N_13879,N_13515,N_13709);
or U13880 (N_13880,N_13689,N_13539);
nor U13881 (N_13881,N_13669,N_13505);
nand U13882 (N_13882,N_13705,N_13569);
xor U13883 (N_13883,N_13581,N_13616);
nor U13884 (N_13884,N_13620,N_13696);
nor U13885 (N_13885,N_13579,N_13629);
and U13886 (N_13886,N_13749,N_13621);
or U13887 (N_13887,N_13661,N_13705);
nand U13888 (N_13888,N_13713,N_13508);
nor U13889 (N_13889,N_13586,N_13671);
or U13890 (N_13890,N_13696,N_13653);
and U13891 (N_13891,N_13570,N_13674);
or U13892 (N_13892,N_13734,N_13720);
xor U13893 (N_13893,N_13702,N_13727);
xnor U13894 (N_13894,N_13673,N_13537);
and U13895 (N_13895,N_13616,N_13514);
or U13896 (N_13896,N_13690,N_13704);
nor U13897 (N_13897,N_13502,N_13632);
and U13898 (N_13898,N_13592,N_13670);
nand U13899 (N_13899,N_13558,N_13733);
nand U13900 (N_13900,N_13548,N_13636);
xor U13901 (N_13901,N_13703,N_13632);
and U13902 (N_13902,N_13582,N_13728);
or U13903 (N_13903,N_13575,N_13659);
or U13904 (N_13904,N_13517,N_13695);
and U13905 (N_13905,N_13746,N_13625);
xnor U13906 (N_13906,N_13540,N_13522);
and U13907 (N_13907,N_13674,N_13624);
or U13908 (N_13908,N_13689,N_13697);
xnor U13909 (N_13909,N_13547,N_13644);
and U13910 (N_13910,N_13709,N_13533);
nor U13911 (N_13911,N_13740,N_13516);
and U13912 (N_13912,N_13505,N_13687);
or U13913 (N_13913,N_13715,N_13695);
nand U13914 (N_13914,N_13558,N_13527);
nor U13915 (N_13915,N_13655,N_13634);
nor U13916 (N_13916,N_13550,N_13578);
nor U13917 (N_13917,N_13525,N_13619);
nor U13918 (N_13918,N_13566,N_13624);
or U13919 (N_13919,N_13600,N_13580);
and U13920 (N_13920,N_13522,N_13695);
xor U13921 (N_13921,N_13508,N_13710);
nand U13922 (N_13922,N_13612,N_13667);
nand U13923 (N_13923,N_13639,N_13627);
or U13924 (N_13924,N_13611,N_13669);
and U13925 (N_13925,N_13565,N_13703);
nor U13926 (N_13926,N_13697,N_13507);
and U13927 (N_13927,N_13746,N_13587);
nand U13928 (N_13928,N_13703,N_13549);
nor U13929 (N_13929,N_13537,N_13609);
xnor U13930 (N_13930,N_13641,N_13685);
and U13931 (N_13931,N_13527,N_13704);
nor U13932 (N_13932,N_13565,N_13704);
nor U13933 (N_13933,N_13630,N_13612);
nor U13934 (N_13934,N_13562,N_13652);
or U13935 (N_13935,N_13644,N_13679);
and U13936 (N_13936,N_13567,N_13581);
and U13937 (N_13937,N_13580,N_13641);
or U13938 (N_13938,N_13673,N_13571);
nor U13939 (N_13939,N_13503,N_13538);
nor U13940 (N_13940,N_13685,N_13599);
nand U13941 (N_13941,N_13610,N_13711);
and U13942 (N_13942,N_13571,N_13746);
nor U13943 (N_13943,N_13688,N_13686);
and U13944 (N_13944,N_13582,N_13724);
nand U13945 (N_13945,N_13712,N_13724);
or U13946 (N_13946,N_13694,N_13618);
and U13947 (N_13947,N_13584,N_13538);
nor U13948 (N_13948,N_13541,N_13625);
nand U13949 (N_13949,N_13639,N_13668);
nand U13950 (N_13950,N_13741,N_13632);
nor U13951 (N_13951,N_13744,N_13736);
nand U13952 (N_13952,N_13723,N_13569);
and U13953 (N_13953,N_13614,N_13646);
nor U13954 (N_13954,N_13545,N_13526);
xor U13955 (N_13955,N_13612,N_13506);
and U13956 (N_13956,N_13549,N_13566);
xnor U13957 (N_13957,N_13652,N_13558);
nor U13958 (N_13958,N_13564,N_13567);
nor U13959 (N_13959,N_13591,N_13647);
or U13960 (N_13960,N_13639,N_13505);
nand U13961 (N_13961,N_13685,N_13738);
or U13962 (N_13962,N_13545,N_13619);
nand U13963 (N_13963,N_13543,N_13701);
and U13964 (N_13964,N_13642,N_13617);
xnor U13965 (N_13965,N_13652,N_13722);
nand U13966 (N_13966,N_13574,N_13657);
nand U13967 (N_13967,N_13553,N_13613);
xor U13968 (N_13968,N_13606,N_13556);
or U13969 (N_13969,N_13570,N_13689);
and U13970 (N_13970,N_13659,N_13694);
or U13971 (N_13971,N_13707,N_13723);
or U13972 (N_13972,N_13600,N_13709);
xnor U13973 (N_13973,N_13725,N_13601);
nand U13974 (N_13974,N_13634,N_13622);
and U13975 (N_13975,N_13644,N_13533);
xnor U13976 (N_13976,N_13504,N_13730);
and U13977 (N_13977,N_13547,N_13638);
and U13978 (N_13978,N_13610,N_13582);
or U13979 (N_13979,N_13593,N_13743);
or U13980 (N_13980,N_13708,N_13649);
nor U13981 (N_13981,N_13628,N_13664);
xnor U13982 (N_13982,N_13549,N_13695);
nor U13983 (N_13983,N_13741,N_13563);
nand U13984 (N_13984,N_13516,N_13515);
and U13985 (N_13985,N_13530,N_13554);
nor U13986 (N_13986,N_13731,N_13628);
nand U13987 (N_13987,N_13698,N_13582);
and U13988 (N_13988,N_13593,N_13649);
nor U13989 (N_13989,N_13624,N_13555);
or U13990 (N_13990,N_13702,N_13636);
or U13991 (N_13991,N_13537,N_13551);
nor U13992 (N_13992,N_13731,N_13528);
or U13993 (N_13993,N_13642,N_13612);
nand U13994 (N_13994,N_13666,N_13726);
xor U13995 (N_13995,N_13626,N_13673);
and U13996 (N_13996,N_13664,N_13530);
nand U13997 (N_13997,N_13597,N_13520);
nand U13998 (N_13998,N_13637,N_13582);
nor U13999 (N_13999,N_13663,N_13705);
nor U14000 (N_14000,N_13948,N_13849);
or U14001 (N_14001,N_13875,N_13773);
xor U14002 (N_14002,N_13775,N_13898);
xor U14003 (N_14003,N_13820,N_13764);
nor U14004 (N_14004,N_13823,N_13783);
and U14005 (N_14005,N_13761,N_13767);
xnor U14006 (N_14006,N_13950,N_13928);
nand U14007 (N_14007,N_13754,N_13834);
or U14008 (N_14008,N_13765,N_13944);
xnor U14009 (N_14009,N_13779,N_13983);
xnor U14010 (N_14010,N_13840,N_13871);
nand U14011 (N_14011,N_13794,N_13947);
and U14012 (N_14012,N_13795,N_13770);
nor U14013 (N_14013,N_13828,N_13908);
xnor U14014 (N_14014,N_13774,N_13857);
nand U14015 (N_14015,N_13762,N_13866);
and U14016 (N_14016,N_13917,N_13913);
or U14017 (N_14017,N_13972,N_13781);
or U14018 (N_14018,N_13780,N_13812);
nor U14019 (N_14019,N_13964,N_13938);
nand U14020 (N_14020,N_13921,N_13895);
or U14021 (N_14021,N_13933,N_13784);
nor U14022 (N_14022,N_13778,N_13776);
or U14023 (N_14023,N_13988,N_13982);
xnor U14024 (N_14024,N_13924,N_13769);
or U14025 (N_14025,N_13884,N_13854);
xnor U14026 (N_14026,N_13966,N_13961);
xor U14027 (N_14027,N_13905,N_13865);
or U14028 (N_14028,N_13886,N_13827);
nand U14029 (N_14029,N_13887,N_13850);
nor U14030 (N_14030,N_13977,N_13830);
or U14031 (N_14031,N_13971,N_13806);
xor U14032 (N_14032,N_13943,N_13757);
xor U14033 (N_14033,N_13996,N_13911);
nor U14034 (N_14034,N_13959,N_13890);
and U14035 (N_14035,N_13804,N_13897);
xnor U14036 (N_14036,N_13906,N_13949);
xnor U14037 (N_14037,N_13867,N_13758);
nor U14038 (N_14038,N_13766,N_13907);
or U14039 (N_14039,N_13946,N_13880);
nand U14040 (N_14040,N_13892,N_13851);
and U14041 (N_14041,N_13914,N_13909);
or U14042 (N_14042,N_13863,N_13912);
nand U14043 (N_14043,N_13878,N_13787);
and U14044 (N_14044,N_13956,N_13796);
nor U14045 (N_14045,N_13888,N_13979);
xnor U14046 (N_14046,N_13902,N_13940);
or U14047 (N_14047,N_13965,N_13874);
and U14048 (N_14048,N_13922,N_13893);
xnor U14049 (N_14049,N_13882,N_13957);
and U14050 (N_14050,N_13879,N_13984);
nand U14051 (N_14051,N_13894,N_13763);
xor U14052 (N_14052,N_13899,N_13997);
nand U14053 (N_14053,N_13829,N_13861);
or U14054 (N_14054,N_13808,N_13927);
and U14055 (N_14055,N_13992,N_13817);
and U14056 (N_14056,N_13752,N_13836);
nand U14057 (N_14057,N_13864,N_13995);
nor U14058 (N_14058,N_13855,N_13807);
nand U14059 (N_14059,N_13993,N_13968);
and U14060 (N_14060,N_13797,N_13990);
nand U14061 (N_14061,N_13805,N_13788);
xnor U14062 (N_14062,N_13841,N_13809);
nand U14063 (N_14063,N_13816,N_13802);
or U14064 (N_14064,N_13777,N_13881);
xor U14065 (N_14065,N_13824,N_13852);
nand U14066 (N_14066,N_13853,N_13791);
nor U14067 (N_14067,N_13792,N_13785);
nand U14068 (N_14068,N_13953,N_13937);
xor U14069 (N_14069,N_13793,N_13955);
nand U14070 (N_14070,N_13985,N_13870);
or U14071 (N_14071,N_13932,N_13991);
nand U14072 (N_14072,N_13942,N_13837);
nand U14073 (N_14073,N_13903,N_13969);
nand U14074 (N_14074,N_13869,N_13960);
or U14075 (N_14075,N_13821,N_13926);
nor U14076 (N_14076,N_13930,N_13848);
nand U14077 (N_14077,N_13939,N_13974);
nor U14078 (N_14078,N_13856,N_13962);
and U14079 (N_14079,N_13825,N_13831);
and U14080 (N_14080,N_13973,N_13981);
nand U14081 (N_14081,N_13967,N_13919);
or U14082 (N_14082,N_13916,N_13786);
xor U14083 (N_14083,N_13904,N_13835);
or U14084 (N_14084,N_13790,N_13954);
nor U14085 (N_14085,N_13900,N_13929);
nor U14086 (N_14086,N_13803,N_13789);
and U14087 (N_14087,N_13891,N_13759);
and U14088 (N_14088,N_13975,N_13818);
or U14089 (N_14089,N_13842,N_13935);
and U14090 (N_14090,N_13994,N_13896);
nor U14091 (N_14091,N_13751,N_13883);
nand U14092 (N_14092,N_13800,N_13976);
xnor U14093 (N_14093,N_13999,N_13868);
xor U14094 (N_14094,N_13859,N_13755);
or U14095 (N_14095,N_13920,N_13782);
or U14096 (N_14096,N_13819,N_13877);
nor U14097 (N_14097,N_13798,N_13862);
and U14098 (N_14098,N_13945,N_13941);
nand U14099 (N_14099,N_13970,N_13858);
and U14100 (N_14100,N_13799,N_13915);
xor U14101 (N_14101,N_13872,N_13980);
or U14102 (N_14102,N_13814,N_13952);
nor U14103 (N_14103,N_13987,N_13844);
and U14104 (N_14104,N_13958,N_13936);
nand U14105 (N_14105,N_13815,N_13832);
xor U14106 (N_14106,N_13873,N_13918);
xor U14107 (N_14107,N_13925,N_13951);
nand U14108 (N_14108,N_13826,N_13813);
and U14109 (N_14109,N_13901,N_13750);
nand U14110 (N_14110,N_13998,N_13771);
nand U14111 (N_14111,N_13923,N_13833);
or U14112 (N_14112,N_13845,N_13989);
or U14113 (N_14113,N_13810,N_13822);
nor U14114 (N_14114,N_13963,N_13934);
or U14115 (N_14115,N_13839,N_13838);
nor U14116 (N_14116,N_13860,N_13986);
nand U14117 (N_14117,N_13811,N_13847);
nor U14118 (N_14118,N_13843,N_13768);
nor U14119 (N_14119,N_13978,N_13756);
xnor U14120 (N_14120,N_13889,N_13760);
xnor U14121 (N_14121,N_13772,N_13910);
or U14122 (N_14122,N_13885,N_13753);
and U14123 (N_14123,N_13846,N_13801);
and U14124 (N_14124,N_13876,N_13931);
or U14125 (N_14125,N_13797,N_13957);
xnor U14126 (N_14126,N_13803,N_13765);
nor U14127 (N_14127,N_13828,N_13903);
xor U14128 (N_14128,N_13897,N_13954);
nor U14129 (N_14129,N_13805,N_13943);
nor U14130 (N_14130,N_13840,N_13861);
or U14131 (N_14131,N_13940,N_13990);
nand U14132 (N_14132,N_13867,N_13989);
nor U14133 (N_14133,N_13943,N_13888);
xnor U14134 (N_14134,N_13967,N_13861);
and U14135 (N_14135,N_13767,N_13855);
nand U14136 (N_14136,N_13772,N_13904);
and U14137 (N_14137,N_13919,N_13831);
and U14138 (N_14138,N_13792,N_13959);
nor U14139 (N_14139,N_13949,N_13852);
xnor U14140 (N_14140,N_13782,N_13850);
nand U14141 (N_14141,N_13790,N_13967);
and U14142 (N_14142,N_13877,N_13776);
and U14143 (N_14143,N_13799,N_13996);
nand U14144 (N_14144,N_13838,N_13958);
and U14145 (N_14145,N_13869,N_13817);
nand U14146 (N_14146,N_13981,N_13922);
xnor U14147 (N_14147,N_13796,N_13808);
nor U14148 (N_14148,N_13828,N_13829);
or U14149 (N_14149,N_13800,N_13888);
or U14150 (N_14150,N_13883,N_13761);
or U14151 (N_14151,N_13822,N_13904);
and U14152 (N_14152,N_13856,N_13924);
and U14153 (N_14153,N_13829,N_13865);
or U14154 (N_14154,N_13796,N_13963);
nor U14155 (N_14155,N_13926,N_13825);
nand U14156 (N_14156,N_13865,N_13836);
and U14157 (N_14157,N_13918,N_13796);
xor U14158 (N_14158,N_13820,N_13811);
nand U14159 (N_14159,N_13968,N_13961);
nor U14160 (N_14160,N_13977,N_13824);
xor U14161 (N_14161,N_13924,N_13836);
nor U14162 (N_14162,N_13982,N_13858);
and U14163 (N_14163,N_13946,N_13958);
xor U14164 (N_14164,N_13890,N_13942);
nor U14165 (N_14165,N_13952,N_13755);
nand U14166 (N_14166,N_13903,N_13751);
or U14167 (N_14167,N_13938,N_13913);
nor U14168 (N_14168,N_13938,N_13825);
xor U14169 (N_14169,N_13771,N_13789);
or U14170 (N_14170,N_13998,N_13808);
nor U14171 (N_14171,N_13803,N_13947);
and U14172 (N_14172,N_13842,N_13852);
xor U14173 (N_14173,N_13935,N_13876);
and U14174 (N_14174,N_13845,N_13947);
nand U14175 (N_14175,N_13799,N_13807);
nand U14176 (N_14176,N_13765,N_13863);
and U14177 (N_14177,N_13879,N_13992);
and U14178 (N_14178,N_13842,N_13937);
or U14179 (N_14179,N_13896,N_13946);
and U14180 (N_14180,N_13976,N_13901);
and U14181 (N_14181,N_13806,N_13854);
or U14182 (N_14182,N_13927,N_13923);
or U14183 (N_14183,N_13950,N_13831);
nor U14184 (N_14184,N_13864,N_13921);
and U14185 (N_14185,N_13899,N_13772);
or U14186 (N_14186,N_13906,N_13847);
xor U14187 (N_14187,N_13997,N_13972);
or U14188 (N_14188,N_13999,N_13967);
xnor U14189 (N_14189,N_13855,N_13809);
and U14190 (N_14190,N_13836,N_13937);
xor U14191 (N_14191,N_13813,N_13873);
and U14192 (N_14192,N_13824,N_13966);
nor U14193 (N_14193,N_13759,N_13827);
and U14194 (N_14194,N_13803,N_13881);
nor U14195 (N_14195,N_13802,N_13915);
and U14196 (N_14196,N_13935,N_13840);
and U14197 (N_14197,N_13837,N_13990);
nand U14198 (N_14198,N_13768,N_13902);
nand U14199 (N_14199,N_13941,N_13827);
nor U14200 (N_14200,N_13851,N_13971);
xor U14201 (N_14201,N_13802,N_13885);
or U14202 (N_14202,N_13949,N_13966);
nor U14203 (N_14203,N_13782,N_13772);
nor U14204 (N_14204,N_13793,N_13995);
xnor U14205 (N_14205,N_13939,N_13923);
xor U14206 (N_14206,N_13753,N_13870);
and U14207 (N_14207,N_13886,N_13774);
nand U14208 (N_14208,N_13835,N_13879);
nor U14209 (N_14209,N_13760,N_13757);
xnor U14210 (N_14210,N_13813,N_13871);
nand U14211 (N_14211,N_13833,N_13827);
nor U14212 (N_14212,N_13876,N_13831);
xor U14213 (N_14213,N_13845,N_13805);
and U14214 (N_14214,N_13841,N_13760);
nand U14215 (N_14215,N_13811,N_13910);
xnor U14216 (N_14216,N_13832,N_13836);
nand U14217 (N_14217,N_13818,N_13775);
xnor U14218 (N_14218,N_13783,N_13931);
nor U14219 (N_14219,N_13759,N_13922);
nand U14220 (N_14220,N_13782,N_13938);
or U14221 (N_14221,N_13934,N_13937);
or U14222 (N_14222,N_13768,N_13983);
xnor U14223 (N_14223,N_13879,N_13823);
or U14224 (N_14224,N_13872,N_13830);
or U14225 (N_14225,N_13823,N_13907);
and U14226 (N_14226,N_13932,N_13848);
or U14227 (N_14227,N_13931,N_13865);
xnor U14228 (N_14228,N_13851,N_13816);
xor U14229 (N_14229,N_13802,N_13910);
nand U14230 (N_14230,N_13984,N_13883);
or U14231 (N_14231,N_13931,N_13764);
nor U14232 (N_14232,N_13783,N_13851);
and U14233 (N_14233,N_13816,N_13877);
nand U14234 (N_14234,N_13875,N_13819);
or U14235 (N_14235,N_13991,N_13966);
and U14236 (N_14236,N_13769,N_13970);
nand U14237 (N_14237,N_13874,N_13773);
nand U14238 (N_14238,N_13823,N_13899);
nor U14239 (N_14239,N_13814,N_13972);
and U14240 (N_14240,N_13987,N_13897);
nand U14241 (N_14241,N_13918,N_13807);
xnor U14242 (N_14242,N_13872,N_13852);
or U14243 (N_14243,N_13905,N_13761);
nand U14244 (N_14244,N_13909,N_13901);
or U14245 (N_14245,N_13975,N_13952);
xnor U14246 (N_14246,N_13899,N_13767);
nand U14247 (N_14247,N_13785,N_13760);
nor U14248 (N_14248,N_13761,N_13819);
xor U14249 (N_14249,N_13808,N_13859);
nand U14250 (N_14250,N_14127,N_14017);
nand U14251 (N_14251,N_14161,N_14086);
and U14252 (N_14252,N_14095,N_14003);
and U14253 (N_14253,N_14000,N_14122);
nor U14254 (N_14254,N_14205,N_14227);
nor U14255 (N_14255,N_14045,N_14190);
nor U14256 (N_14256,N_14139,N_14005);
and U14257 (N_14257,N_14211,N_14200);
xnor U14258 (N_14258,N_14133,N_14018);
and U14259 (N_14259,N_14060,N_14083);
and U14260 (N_14260,N_14091,N_14144);
nand U14261 (N_14261,N_14110,N_14080);
nand U14262 (N_14262,N_14111,N_14062);
nor U14263 (N_14263,N_14103,N_14069);
and U14264 (N_14264,N_14226,N_14006);
nor U14265 (N_14265,N_14021,N_14100);
and U14266 (N_14266,N_14240,N_14028);
nand U14267 (N_14267,N_14037,N_14019);
xor U14268 (N_14268,N_14189,N_14158);
or U14269 (N_14269,N_14206,N_14112);
or U14270 (N_14270,N_14081,N_14027);
xor U14271 (N_14271,N_14098,N_14185);
nand U14272 (N_14272,N_14076,N_14214);
and U14273 (N_14273,N_14188,N_14044);
nor U14274 (N_14274,N_14136,N_14038);
and U14275 (N_14275,N_14047,N_14030);
nand U14276 (N_14276,N_14223,N_14154);
xnor U14277 (N_14277,N_14014,N_14164);
nand U14278 (N_14278,N_14070,N_14106);
nand U14279 (N_14279,N_14124,N_14064);
nor U14280 (N_14280,N_14007,N_14011);
nor U14281 (N_14281,N_14013,N_14043);
nand U14282 (N_14282,N_14022,N_14036);
and U14283 (N_14283,N_14169,N_14094);
nor U14284 (N_14284,N_14002,N_14101);
and U14285 (N_14285,N_14152,N_14222);
and U14286 (N_14286,N_14221,N_14247);
xnor U14287 (N_14287,N_14046,N_14059);
nand U14288 (N_14288,N_14207,N_14004);
and U14289 (N_14289,N_14160,N_14029);
xnor U14290 (N_14290,N_14239,N_14143);
nor U14291 (N_14291,N_14042,N_14114);
and U14292 (N_14292,N_14132,N_14151);
xnor U14293 (N_14293,N_14097,N_14031);
xnor U14294 (N_14294,N_14148,N_14129);
nor U14295 (N_14295,N_14054,N_14196);
xor U14296 (N_14296,N_14245,N_14096);
and U14297 (N_14297,N_14232,N_14192);
xnor U14298 (N_14298,N_14179,N_14071);
or U14299 (N_14299,N_14033,N_14118);
nand U14300 (N_14300,N_14170,N_14012);
and U14301 (N_14301,N_14116,N_14215);
or U14302 (N_14302,N_14180,N_14078);
nand U14303 (N_14303,N_14236,N_14153);
nor U14304 (N_14304,N_14246,N_14177);
and U14305 (N_14305,N_14218,N_14165);
or U14306 (N_14306,N_14168,N_14150);
nor U14307 (N_14307,N_14121,N_14008);
or U14308 (N_14308,N_14217,N_14079);
nand U14309 (N_14309,N_14066,N_14141);
and U14310 (N_14310,N_14204,N_14191);
nor U14311 (N_14311,N_14082,N_14203);
xnor U14312 (N_14312,N_14175,N_14210);
and U14313 (N_14313,N_14052,N_14182);
or U14314 (N_14314,N_14237,N_14209);
nand U14315 (N_14315,N_14041,N_14113);
and U14316 (N_14316,N_14193,N_14202);
xnor U14317 (N_14317,N_14194,N_14174);
or U14318 (N_14318,N_14099,N_14163);
xor U14319 (N_14319,N_14092,N_14142);
nand U14320 (N_14320,N_14183,N_14159);
nand U14321 (N_14321,N_14093,N_14199);
and U14322 (N_14322,N_14087,N_14072);
nand U14323 (N_14323,N_14224,N_14230);
nand U14324 (N_14324,N_14241,N_14181);
xnor U14325 (N_14325,N_14024,N_14137);
xor U14326 (N_14326,N_14249,N_14243);
and U14327 (N_14327,N_14140,N_14147);
or U14328 (N_14328,N_14228,N_14178);
nand U14329 (N_14329,N_14242,N_14089);
nor U14330 (N_14330,N_14120,N_14049);
xnor U14331 (N_14331,N_14172,N_14010);
and U14332 (N_14332,N_14119,N_14219);
or U14333 (N_14333,N_14023,N_14195);
and U14334 (N_14334,N_14171,N_14051);
nor U14335 (N_14335,N_14234,N_14048);
xor U14336 (N_14336,N_14088,N_14220);
nand U14337 (N_14337,N_14117,N_14084);
or U14338 (N_14338,N_14156,N_14032);
nor U14339 (N_14339,N_14131,N_14216);
nand U14340 (N_14340,N_14149,N_14248);
nor U14341 (N_14341,N_14102,N_14025);
nor U14342 (N_14342,N_14238,N_14001);
and U14343 (N_14343,N_14115,N_14055);
or U14344 (N_14344,N_14077,N_14128);
and U14345 (N_14345,N_14184,N_14105);
and U14346 (N_14346,N_14073,N_14186);
nand U14347 (N_14347,N_14157,N_14075);
or U14348 (N_14348,N_14212,N_14126);
nand U14349 (N_14349,N_14090,N_14067);
nor U14350 (N_14350,N_14229,N_14166);
or U14351 (N_14351,N_14058,N_14040);
or U14352 (N_14352,N_14063,N_14225);
or U14353 (N_14353,N_14016,N_14173);
or U14354 (N_14354,N_14056,N_14085);
or U14355 (N_14355,N_14020,N_14015);
or U14356 (N_14356,N_14035,N_14125);
or U14357 (N_14357,N_14109,N_14123);
nand U14358 (N_14358,N_14145,N_14034);
and U14359 (N_14359,N_14208,N_14068);
nor U14360 (N_14360,N_14201,N_14135);
nor U14361 (N_14361,N_14138,N_14162);
and U14362 (N_14362,N_14057,N_14213);
nor U14363 (N_14363,N_14167,N_14155);
xor U14364 (N_14364,N_14244,N_14039);
and U14365 (N_14365,N_14104,N_14146);
and U14366 (N_14366,N_14107,N_14074);
and U14367 (N_14367,N_14065,N_14187);
and U14368 (N_14368,N_14050,N_14053);
nor U14369 (N_14369,N_14130,N_14009);
and U14370 (N_14370,N_14176,N_14197);
or U14371 (N_14371,N_14026,N_14061);
xnor U14372 (N_14372,N_14233,N_14235);
nor U14373 (N_14373,N_14198,N_14108);
xor U14374 (N_14374,N_14134,N_14231);
or U14375 (N_14375,N_14141,N_14099);
xor U14376 (N_14376,N_14073,N_14062);
and U14377 (N_14377,N_14066,N_14124);
and U14378 (N_14378,N_14194,N_14081);
nand U14379 (N_14379,N_14129,N_14031);
or U14380 (N_14380,N_14112,N_14218);
nand U14381 (N_14381,N_14148,N_14087);
or U14382 (N_14382,N_14003,N_14249);
or U14383 (N_14383,N_14241,N_14005);
nor U14384 (N_14384,N_14116,N_14203);
nor U14385 (N_14385,N_14076,N_14113);
nor U14386 (N_14386,N_14241,N_14171);
nor U14387 (N_14387,N_14194,N_14061);
and U14388 (N_14388,N_14196,N_14078);
nand U14389 (N_14389,N_14059,N_14159);
or U14390 (N_14390,N_14117,N_14247);
and U14391 (N_14391,N_14043,N_14170);
and U14392 (N_14392,N_14187,N_14047);
and U14393 (N_14393,N_14232,N_14210);
or U14394 (N_14394,N_14240,N_14004);
xor U14395 (N_14395,N_14001,N_14149);
nor U14396 (N_14396,N_14021,N_14105);
nor U14397 (N_14397,N_14246,N_14060);
and U14398 (N_14398,N_14135,N_14218);
and U14399 (N_14399,N_14233,N_14094);
xor U14400 (N_14400,N_14237,N_14116);
or U14401 (N_14401,N_14132,N_14226);
nand U14402 (N_14402,N_14105,N_14013);
nand U14403 (N_14403,N_14070,N_14147);
nor U14404 (N_14404,N_14141,N_14244);
or U14405 (N_14405,N_14182,N_14017);
xnor U14406 (N_14406,N_14029,N_14106);
or U14407 (N_14407,N_14066,N_14222);
or U14408 (N_14408,N_14162,N_14050);
xnor U14409 (N_14409,N_14098,N_14193);
nand U14410 (N_14410,N_14059,N_14004);
nor U14411 (N_14411,N_14155,N_14222);
nor U14412 (N_14412,N_14074,N_14236);
xor U14413 (N_14413,N_14035,N_14060);
and U14414 (N_14414,N_14186,N_14154);
xnor U14415 (N_14415,N_14019,N_14116);
and U14416 (N_14416,N_14058,N_14172);
nor U14417 (N_14417,N_14066,N_14054);
xnor U14418 (N_14418,N_14053,N_14009);
or U14419 (N_14419,N_14249,N_14101);
or U14420 (N_14420,N_14184,N_14063);
nand U14421 (N_14421,N_14222,N_14143);
or U14422 (N_14422,N_14150,N_14060);
or U14423 (N_14423,N_14050,N_14176);
and U14424 (N_14424,N_14130,N_14170);
or U14425 (N_14425,N_14036,N_14192);
and U14426 (N_14426,N_14117,N_14095);
and U14427 (N_14427,N_14154,N_14191);
nand U14428 (N_14428,N_14097,N_14198);
and U14429 (N_14429,N_14220,N_14032);
and U14430 (N_14430,N_14171,N_14120);
or U14431 (N_14431,N_14221,N_14007);
nand U14432 (N_14432,N_14048,N_14012);
or U14433 (N_14433,N_14003,N_14073);
nand U14434 (N_14434,N_14085,N_14111);
nand U14435 (N_14435,N_14030,N_14157);
nand U14436 (N_14436,N_14134,N_14131);
xnor U14437 (N_14437,N_14209,N_14049);
and U14438 (N_14438,N_14042,N_14049);
nand U14439 (N_14439,N_14060,N_14106);
xor U14440 (N_14440,N_14225,N_14110);
nand U14441 (N_14441,N_14217,N_14205);
and U14442 (N_14442,N_14119,N_14091);
nand U14443 (N_14443,N_14096,N_14042);
nand U14444 (N_14444,N_14141,N_14097);
or U14445 (N_14445,N_14165,N_14115);
nor U14446 (N_14446,N_14220,N_14109);
xnor U14447 (N_14447,N_14028,N_14076);
and U14448 (N_14448,N_14078,N_14245);
and U14449 (N_14449,N_14116,N_14064);
or U14450 (N_14450,N_14164,N_14219);
and U14451 (N_14451,N_14030,N_14112);
or U14452 (N_14452,N_14226,N_14022);
and U14453 (N_14453,N_14153,N_14019);
nand U14454 (N_14454,N_14047,N_14057);
or U14455 (N_14455,N_14212,N_14194);
nand U14456 (N_14456,N_14176,N_14124);
nor U14457 (N_14457,N_14096,N_14105);
and U14458 (N_14458,N_14190,N_14148);
nor U14459 (N_14459,N_14071,N_14079);
xor U14460 (N_14460,N_14189,N_14013);
or U14461 (N_14461,N_14051,N_14077);
or U14462 (N_14462,N_14004,N_14154);
xnor U14463 (N_14463,N_14123,N_14097);
nand U14464 (N_14464,N_14004,N_14229);
xnor U14465 (N_14465,N_14171,N_14231);
and U14466 (N_14466,N_14182,N_14066);
xnor U14467 (N_14467,N_14000,N_14220);
and U14468 (N_14468,N_14220,N_14132);
xor U14469 (N_14469,N_14144,N_14176);
or U14470 (N_14470,N_14244,N_14126);
nor U14471 (N_14471,N_14197,N_14057);
and U14472 (N_14472,N_14218,N_14245);
xnor U14473 (N_14473,N_14248,N_14187);
nand U14474 (N_14474,N_14150,N_14040);
nand U14475 (N_14475,N_14077,N_14035);
nor U14476 (N_14476,N_14133,N_14236);
nor U14477 (N_14477,N_14169,N_14204);
nor U14478 (N_14478,N_14136,N_14117);
nand U14479 (N_14479,N_14146,N_14206);
xnor U14480 (N_14480,N_14199,N_14083);
xor U14481 (N_14481,N_14077,N_14049);
xor U14482 (N_14482,N_14188,N_14022);
nor U14483 (N_14483,N_14247,N_14096);
and U14484 (N_14484,N_14247,N_14052);
xor U14485 (N_14485,N_14234,N_14129);
xor U14486 (N_14486,N_14199,N_14212);
or U14487 (N_14487,N_14178,N_14052);
nand U14488 (N_14488,N_14111,N_14168);
or U14489 (N_14489,N_14012,N_14049);
and U14490 (N_14490,N_14188,N_14119);
nor U14491 (N_14491,N_14064,N_14011);
or U14492 (N_14492,N_14100,N_14104);
or U14493 (N_14493,N_14226,N_14204);
and U14494 (N_14494,N_14017,N_14168);
nor U14495 (N_14495,N_14047,N_14202);
and U14496 (N_14496,N_14163,N_14168);
and U14497 (N_14497,N_14206,N_14102);
and U14498 (N_14498,N_14009,N_14124);
xnor U14499 (N_14499,N_14121,N_14189);
xnor U14500 (N_14500,N_14425,N_14286);
or U14501 (N_14501,N_14334,N_14284);
xnor U14502 (N_14502,N_14441,N_14408);
nand U14503 (N_14503,N_14363,N_14456);
or U14504 (N_14504,N_14279,N_14494);
nor U14505 (N_14505,N_14342,N_14454);
nor U14506 (N_14506,N_14319,N_14267);
or U14507 (N_14507,N_14305,N_14476);
nand U14508 (N_14508,N_14432,N_14352);
nor U14509 (N_14509,N_14429,N_14440);
and U14510 (N_14510,N_14424,N_14426);
nor U14511 (N_14511,N_14478,N_14451);
xnor U14512 (N_14512,N_14472,N_14262);
xor U14513 (N_14513,N_14459,N_14396);
nand U14514 (N_14514,N_14416,N_14350);
xnor U14515 (N_14515,N_14268,N_14353);
and U14516 (N_14516,N_14477,N_14392);
xor U14517 (N_14517,N_14292,N_14447);
nor U14518 (N_14518,N_14266,N_14475);
or U14519 (N_14519,N_14322,N_14498);
or U14520 (N_14520,N_14274,N_14313);
xor U14521 (N_14521,N_14341,N_14483);
nand U14522 (N_14522,N_14330,N_14436);
nand U14523 (N_14523,N_14395,N_14273);
or U14524 (N_14524,N_14321,N_14259);
nor U14525 (N_14525,N_14470,N_14423);
and U14526 (N_14526,N_14455,N_14289);
nand U14527 (N_14527,N_14439,N_14324);
nand U14528 (N_14528,N_14466,N_14445);
nor U14529 (N_14529,N_14347,N_14453);
nor U14530 (N_14530,N_14378,N_14356);
and U14531 (N_14531,N_14474,N_14282);
or U14532 (N_14532,N_14291,N_14487);
or U14533 (N_14533,N_14278,N_14308);
or U14534 (N_14534,N_14302,N_14486);
nand U14535 (N_14535,N_14258,N_14370);
nand U14536 (N_14536,N_14371,N_14269);
nor U14537 (N_14537,N_14435,N_14419);
or U14538 (N_14538,N_14318,N_14479);
xor U14539 (N_14539,N_14387,N_14462);
and U14540 (N_14540,N_14407,N_14499);
and U14541 (N_14541,N_14288,N_14281);
or U14542 (N_14542,N_14303,N_14368);
nand U14543 (N_14543,N_14484,N_14343);
nand U14544 (N_14544,N_14250,N_14492);
nand U14545 (N_14545,N_14497,N_14427);
or U14546 (N_14546,N_14400,N_14351);
nand U14547 (N_14547,N_14490,N_14434);
nor U14548 (N_14548,N_14257,N_14422);
and U14549 (N_14549,N_14331,N_14276);
nor U14550 (N_14550,N_14287,N_14421);
nor U14551 (N_14551,N_14359,N_14468);
xor U14552 (N_14552,N_14409,N_14309);
nand U14553 (N_14553,N_14335,N_14296);
nor U14554 (N_14554,N_14391,N_14283);
nand U14555 (N_14555,N_14323,N_14297);
nand U14556 (N_14556,N_14448,N_14355);
and U14557 (N_14557,N_14430,N_14493);
xnor U14558 (N_14558,N_14326,N_14383);
nand U14559 (N_14559,N_14307,N_14443);
or U14560 (N_14560,N_14294,N_14491);
xnor U14561 (N_14561,N_14373,N_14329);
xnor U14562 (N_14562,N_14364,N_14405);
and U14563 (N_14563,N_14415,N_14338);
xnor U14564 (N_14564,N_14457,N_14315);
and U14565 (N_14565,N_14310,N_14385);
xor U14566 (N_14566,N_14300,N_14403);
nor U14567 (N_14567,N_14265,N_14253);
nand U14568 (N_14568,N_14280,N_14290);
xor U14569 (N_14569,N_14399,N_14384);
nor U14570 (N_14570,N_14366,N_14428);
nand U14571 (N_14571,N_14304,N_14374);
nor U14572 (N_14572,N_14485,N_14301);
or U14573 (N_14573,N_14376,N_14255);
xnor U14574 (N_14574,N_14260,N_14412);
or U14575 (N_14575,N_14452,N_14261);
xnor U14576 (N_14576,N_14460,N_14404);
xor U14577 (N_14577,N_14489,N_14339);
nor U14578 (N_14578,N_14438,N_14377);
xor U14579 (N_14579,N_14410,N_14314);
nor U14580 (N_14580,N_14348,N_14327);
nor U14581 (N_14581,N_14442,N_14437);
and U14582 (N_14582,N_14357,N_14433);
nand U14583 (N_14583,N_14369,N_14345);
nand U14584 (N_14584,N_14496,N_14293);
and U14585 (N_14585,N_14256,N_14458);
xnor U14586 (N_14586,N_14320,N_14482);
or U14587 (N_14587,N_14461,N_14311);
or U14588 (N_14588,N_14271,N_14463);
nand U14589 (N_14589,N_14340,N_14375);
xnor U14590 (N_14590,N_14411,N_14495);
or U14591 (N_14591,N_14480,N_14372);
nor U14592 (N_14592,N_14354,N_14381);
or U14593 (N_14593,N_14316,N_14344);
nand U14594 (N_14594,N_14365,N_14277);
nand U14595 (N_14595,N_14252,N_14469);
and U14596 (N_14596,N_14379,N_14312);
nand U14597 (N_14597,N_14362,N_14481);
nand U14598 (N_14598,N_14471,N_14299);
xnor U14599 (N_14599,N_14473,N_14417);
and U14600 (N_14600,N_14390,N_14251);
and U14601 (N_14601,N_14361,N_14254);
and U14602 (N_14602,N_14488,N_14325);
or U14603 (N_14603,N_14401,N_14336);
and U14604 (N_14604,N_14389,N_14270);
and U14605 (N_14605,N_14380,N_14337);
or U14606 (N_14606,N_14328,N_14446);
nand U14607 (N_14607,N_14386,N_14317);
xor U14608 (N_14608,N_14295,N_14397);
nor U14609 (N_14609,N_14272,N_14467);
nor U14610 (N_14610,N_14420,N_14398);
xor U14611 (N_14611,N_14431,N_14464);
nand U14612 (N_14612,N_14465,N_14444);
nand U14613 (N_14613,N_14418,N_14358);
or U14614 (N_14614,N_14367,N_14450);
nand U14615 (N_14615,N_14264,N_14388);
nand U14616 (N_14616,N_14298,N_14394);
xor U14617 (N_14617,N_14333,N_14382);
nor U14618 (N_14618,N_14406,N_14414);
nor U14619 (N_14619,N_14285,N_14402);
or U14620 (N_14620,N_14263,N_14413);
nand U14621 (N_14621,N_14346,N_14349);
xnor U14622 (N_14622,N_14306,N_14449);
nor U14623 (N_14623,N_14393,N_14332);
and U14624 (N_14624,N_14275,N_14360);
or U14625 (N_14625,N_14260,N_14257);
nand U14626 (N_14626,N_14267,N_14485);
xor U14627 (N_14627,N_14256,N_14461);
nand U14628 (N_14628,N_14297,N_14388);
and U14629 (N_14629,N_14303,N_14362);
xnor U14630 (N_14630,N_14267,N_14471);
nor U14631 (N_14631,N_14441,N_14389);
or U14632 (N_14632,N_14263,N_14424);
nand U14633 (N_14633,N_14400,N_14497);
nor U14634 (N_14634,N_14334,N_14434);
nand U14635 (N_14635,N_14357,N_14452);
nand U14636 (N_14636,N_14274,N_14266);
or U14637 (N_14637,N_14487,N_14409);
or U14638 (N_14638,N_14339,N_14458);
and U14639 (N_14639,N_14405,N_14260);
xor U14640 (N_14640,N_14403,N_14430);
nand U14641 (N_14641,N_14411,N_14406);
or U14642 (N_14642,N_14362,N_14254);
xnor U14643 (N_14643,N_14299,N_14275);
xor U14644 (N_14644,N_14364,N_14325);
and U14645 (N_14645,N_14385,N_14391);
and U14646 (N_14646,N_14264,N_14440);
nand U14647 (N_14647,N_14311,N_14306);
xnor U14648 (N_14648,N_14336,N_14345);
and U14649 (N_14649,N_14264,N_14425);
xor U14650 (N_14650,N_14385,N_14324);
nor U14651 (N_14651,N_14370,N_14279);
xnor U14652 (N_14652,N_14494,N_14368);
and U14653 (N_14653,N_14425,N_14253);
xor U14654 (N_14654,N_14300,N_14309);
xor U14655 (N_14655,N_14376,N_14299);
nand U14656 (N_14656,N_14399,N_14462);
nor U14657 (N_14657,N_14377,N_14437);
xor U14658 (N_14658,N_14368,N_14398);
or U14659 (N_14659,N_14409,N_14418);
nor U14660 (N_14660,N_14488,N_14472);
nand U14661 (N_14661,N_14395,N_14434);
and U14662 (N_14662,N_14294,N_14426);
nand U14663 (N_14663,N_14350,N_14361);
or U14664 (N_14664,N_14338,N_14378);
nor U14665 (N_14665,N_14348,N_14472);
nand U14666 (N_14666,N_14368,N_14302);
xnor U14667 (N_14667,N_14257,N_14452);
nand U14668 (N_14668,N_14299,N_14331);
or U14669 (N_14669,N_14304,N_14356);
nand U14670 (N_14670,N_14278,N_14434);
and U14671 (N_14671,N_14469,N_14470);
nor U14672 (N_14672,N_14418,N_14275);
xnor U14673 (N_14673,N_14491,N_14375);
nor U14674 (N_14674,N_14300,N_14297);
or U14675 (N_14675,N_14491,N_14340);
and U14676 (N_14676,N_14285,N_14441);
or U14677 (N_14677,N_14318,N_14449);
nand U14678 (N_14678,N_14351,N_14257);
xnor U14679 (N_14679,N_14488,N_14297);
nor U14680 (N_14680,N_14491,N_14478);
xor U14681 (N_14681,N_14290,N_14312);
xnor U14682 (N_14682,N_14444,N_14323);
or U14683 (N_14683,N_14463,N_14441);
and U14684 (N_14684,N_14475,N_14426);
and U14685 (N_14685,N_14265,N_14323);
or U14686 (N_14686,N_14420,N_14263);
and U14687 (N_14687,N_14305,N_14477);
nand U14688 (N_14688,N_14407,N_14392);
and U14689 (N_14689,N_14472,N_14269);
nor U14690 (N_14690,N_14420,N_14476);
or U14691 (N_14691,N_14311,N_14370);
and U14692 (N_14692,N_14321,N_14427);
and U14693 (N_14693,N_14317,N_14316);
and U14694 (N_14694,N_14365,N_14303);
nand U14695 (N_14695,N_14464,N_14330);
nand U14696 (N_14696,N_14383,N_14347);
nor U14697 (N_14697,N_14486,N_14424);
nand U14698 (N_14698,N_14398,N_14460);
or U14699 (N_14699,N_14435,N_14308);
nand U14700 (N_14700,N_14400,N_14256);
nor U14701 (N_14701,N_14328,N_14387);
xor U14702 (N_14702,N_14487,N_14432);
and U14703 (N_14703,N_14316,N_14393);
xor U14704 (N_14704,N_14446,N_14374);
xor U14705 (N_14705,N_14256,N_14296);
xor U14706 (N_14706,N_14474,N_14367);
nand U14707 (N_14707,N_14485,N_14333);
nor U14708 (N_14708,N_14345,N_14268);
and U14709 (N_14709,N_14462,N_14461);
xnor U14710 (N_14710,N_14300,N_14417);
nor U14711 (N_14711,N_14259,N_14272);
nor U14712 (N_14712,N_14286,N_14277);
nand U14713 (N_14713,N_14396,N_14378);
or U14714 (N_14714,N_14468,N_14252);
nand U14715 (N_14715,N_14489,N_14449);
xor U14716 (N_14716,N_14327,N_14253);
and U14717 (N_14717,N_14369,N_14362);
xnor U14718 (N_14718,N_14460,N_14440);
xor U14719 (N_14719,N_14319,N_14339);
nor U14720 (N_14720,N_14322,N_14303);
or U14721 (N_14721,N_14340,N_14498);
xnor U14722 (N_14722,N_14402,N_14302);
nor U14723 (N_14723,N_14482,N_14483);
and U14724 (N_14724,N_14271,N_14339);
and U14725 (N_14725,N_14452,N_14414);
or U14726 (N_14726,N_14341,N_14359);
nor U14727 (N_14727,N_14406,N_14472);
and U14728 (N_14728,N_14315,N_14257);
or U14729 (N_14729,N_14313,N_14463);
xnor U14730 (N_14730,N_14255,N_14487);
nand U14731 (N_14731,N_14349,N_14406);
or U14732 (N_14732,N_14321,N_14312);
and U14733 (N_14733,N_14305,N_14422);
nor U14734 (N_14734,N_14257,N_14409);
nor U14735 (N_14735,N_14443,N_14334);
xor U14736 (N_14736,N_14329,N_14352);
and U14737 (N_14737,N_14424,N_14314);
or U14738 (N_14738,N_14493,N_14484);
or U14739 (N_14739,N_14420,N_14366);
nor U14740 (N_14740,N_14269,N_14387);
and U14741 (N_14741,N_14336,N_14332);
or U14742 (N_14742,N_14321,N_14496);
xnor U14743 (N_14743,N_14439,N_14387);
nand U14744 (N_14744,N_14336,N_14331);
and U14745 (N_14745,N_14425,N_14369);
nor U14746 (N_14746,N_14385,N_14406);
xor U14747 (N_14747,N_14314,N_14477);
nor U14748 (N_14748,N_14270,N_14294);
nand U14749 (N_14749,N_14268,N_14415);
nand U14750 (N_14750,N_14533,N_14657);
and U14751 (N_14751,N_14716,N_14596);
and U14752 (N_14752,N_14565,N_14524);
nor U14753 (N_14753,N_14514,N_14679);
or U14754 (N_14754,N_14665,N_14503);
nor U14755 (N_14755,N_14710,N_14559);
and U14756 (N_14756,N_14660,N_14674);
nand U14757 (N_14757,N_14702,N_14672);
nand U14758 (N_14758,N_14521,N_14637);
nand U14759 (N_14759,N_14719,N_14612);
xor U14760 (N_14760,N_14595,N_14537);
xnor U14761 (N_14761,N_14592,N_14510);
or U14762 (N_14762,N_14518,N_14544);
or U14763 (N_14763,N_14547,N_14636);
nand U14764 (N_14764,N_14585,N_14711);
nor U14765 (N_14765,N_14566,N_14737);
xnor U14766 (N_14766,N_14568,N_14605);
nor U14767 (N_14767,N_14651,N_14581);
nand U14768 (N_14768,N_14691,N_14707);
xnor U14769 (N_14769,N_14602,N_14517);
xor U14770 (N_14770,N_14527,N_14747);
xnor U14771 (N_14771,N_14735,N_14722);
nor U14772 (N_14772,N_14617,N_14626);
nor U14773 (N_14773,N_14678,N_14628);
nor U14774 (N_14774,N_14574,N_14616);
or U14775 (N_14775,N_14744,N_14604);
nand U14776 (N_14776,N_14690,N_14646);
or U14777 (N_14777,N_14745,N_14733);
nor U14778 (N_14778,N_14530,N_14557);
xor U14779 (N_14779,N_14538,N_14546);
or U14780 (N_14780,N_14578,N_14587);
and U14781 (N_14781,N_14586,N_14590);
xnor U14782 (N_14782,N_14624,N_14705);
nor U14783 (N_14783,N_14526,N_14562);
nand U14784 (N_14784,N_14550,N_14508);
and U14785 (N_14785,N_14622,N_14593);
or U14786 (N_14786,N_14642,N_14576);
nor U14787 (N_14787,N_14536,N_14502);
nand U14788 (N_14788,N_14531,N_14728);
or U14789 (N_14789,N_14555,N_14714);
nand U14790 (N_14790,N_14696,N_14573);
and U14791 (N_14791,N_14731,N_14726);
xnor U14792 (N_14792,N_14712,N_14720);
nand U14793 (N_14793,N_14706,N_14570);
or U14794 (N_14794,N_14746,N_14654);
or U14795 (N_14795,N_14741,N_14695);
and U14796 (N_14796,N_14739,N_14623);
nor U14797 (N_14797,N_14629,N_14564);
nor U14798 (N_14798,N_14619,N_14529);
xor U14799 (N_14799,N_14615,N_14644);
and U14800 (N_14800,N_14643,N_14727);
nor U14801 (N_14801,N_14507,N_14513);
nor U14802 (N_14802,N_14682,N_14692);
and U14803 (N_14803,N_14600,N_14631);
xnor U14804 (N_14804,N_14650,N_14667);
nand U14805 (N_14805,N_14662,N_14681);
or U14806 (N_14806,N_14670,N_14648);
and U14807 (N_14807,N_14621,N_14668);
or U14808 (N_14808,N_14666,N_14694);
and U14809 (N_14809,N_14689,N_14625);
and U14810 (N_14810,N_14743,N_14511);
or U14811 (N_14811,N_14700,N_14606);
or U14812 (N_14812,N_14532,N_14703);
and U14813 (N_14813,N_14515,N_14675);
or U14814 (N_14814,N_14724,N_14542);
nor U14815 (N_14815,N_14618,N_14734);
or U14816 (N_14816,N_14638,N_14554);
nor U14817 (N_14817,N_14699,N_14601);
xnor U14818 (N_14818,N_14540,N_14609);
nand U14819 (N_14819,N_14528,N_14543);
and U14820 (N_14820,N_14582,N_14556);
xor U14821 (N_14821,N_14680,N_14520);
nor U14822 (N_14822,N_14545,N_14505);
or U14823 (N_14823,N_14561,N_14738);
nor U14824 (N_14824,N_14676,N_14656);
nand U14825 (N_14825,N_14688,N_14693);
nand U14826 (N_14826,N_14649,N_14603);
xnor U14827 (N_14827,N_14580,N_14641);
xnor U14828 (N_14828,N_14658,N_14718);
or U14829 (N_14829,N_14611,N_14599);
nor U14830 (N_14830,N_14610,N_14558);
xnor U14831 (N_14831,N_14652,N_14740);
and U14832 (N_14832,N_14572,N_14639);
nor U14833 (N_14833,N_14630,N_14749);
nand U14834 (N_14834,N_14685,N_14549);
or U14835 (N_14835,N_14584,N_14725);
or U14836 (N_14836,N_14575,N_14598);
nor U14837 (N_14837,N_14519,N_14506);
or U14838 (N_14838,N_14567,N_14664);
or U14839 (N_14839,N_14589,N_14686);
nand U14840 (N_14840,N_14591,N_14500);
and U14841 (N_14841,N_14563,N_14683);
and U14842 (N_14842,N_14512,N_14541);
and U14843 (N_14843,N_14535,N_14551);
nor U14844 (N_14844,N_14653,N_14539);
nand U14845 (N_14845,N_14552,N_14501);
nor U14846 (N_14846,N_14742,N_14697);
nand U14847 (N_14847,N_14687,N_14583);
and U14848 (N_14848,N_14729,N_14560);
or U14849 (N_14849,N_14730,N_14577);
xnor U14850 (N_14850,N_14671,N_14579);
or U14851 (N_14851,N_14548,N_14717);
xor U14852 (N_14852,N_14597,N_14627);
or U14853 (N_14853,N_14522,N_14669);
xnor U14854 (N_14854,N_14516,N_14736);
nor U14855 (N_14855,N_14709,N_14713);
nand U14856 (N_14856,N_14613,N_14640);
nor U14857 (N_14857,N_14553,N_14608);
nand U14858 (N_14858,N_14647,N_14635);
xor U14859 (N_14859,N_14645,N_14594);
nand U14860 (N_14860,N_14634,N_14721);
nand U14861 (N_14861,N_14715,N_14684);
nand U14862 (N_14862,N_14661,N_14534);
xnor U14863 (N_14863,N_14523,N_14708);
or U14864 (N_14864,N_14663,N_14632);
nand U14865 (N_14865,N_14614,N_14571);
nor U14866 (N_14866,N_14701,N_14748);
or U14867 (N_14867,N_14620,N_14588);
nand U14868 (N_14868,N_14607,N_14723);
and U14869 (N_14869,N_14504,N_14655);
nor U14870 (N_14870,N_14509,N_14704);
xor U14871 (N_14871,N_14677,N_14673);
xnor U14872 (N_14872,N_14525,N_14569);
or U14873 (N_14873,N_14732,N_14659);
and U14874 (N_14874,N_14698,N_14633);
nand U14875 (N_14875,N_14691,N_14583);
and U14876 (N_14876,N_14520,N_14653);
xor U14877 (N_14877,N_14714,N_14598);
xor U14878 (N_14878,N_14741,N_14627);
nor U14879 (N_14879,N_14605,N_14689);
nand U14880 (N_14880,N_14673,N_14736);
and U14881 (N_14881,N_14656,N_14680);
nand U14882 (N_14882,N_14723,N_14731);
nand U14883 (N_14883,N_14595,N_14626);
xor U14884 (N_14884,N_14539,N_14571);
nor U14885 (N_14885,N_14568,N_14554);
or U14886 (N_14886,N_14601,N_14744);
nor U14887 (N_14887,N_14617,N_14551);
or U14888 (N_14888,N_14664,N_14696);
or U14889 (N_14889,N_14502,N_14556);
xnor U14890 (N_14890,N_14725,N_14661);
or U14891 (N_14891,N_14616,N_14582);
or U14892 (N_14892,N_14614,N_14542);
nor U14893 (N_14893,N_14668,N_14736);
xnor U14894 (N_14894,N_14686,N_14561);
nand U14895 (N_14895,N_14579,N_14643);
and U14896 (N_14896,N_14692,N_14589);
or U14897 (N_14897,N_14604,N_14728);
and U14898 (N_14898,N_14592,N_14589);
nand U14899 (N_14899,N_14687,N_14657);
nor U14900 (N_14900,N_14557,N_14735);
and U14901 (N_14901,N_14629,N_14702);
xnor U14902 (N_14902,N_14733,N_14727);
nand U14903 (N_14903,N_14723,N_14734);
nand U14904 (N_14904,N_14532,N_14596);
nand U14905 (N_14905,N_14724,N_14596);
xnor U14906 (N_14906,N_14642,N_14643);
or U14907 (N_14907,N_14618,N_14591);
nor U14908 (N_14908,N_14576,N_14673);
nand U14909 (N_14909,N_14572,N_14694);
xnor U14910 (N_14910,N_14510,N_14612);
or U14911 (N_14911,N_14592,N_14717);
or U14912 (N_14912,N_14524,N_14598);
or U14913 (N_14913,N_14530,N_14504);
nor U14914 (N_14914,N_14519,N_14648);
nor U14915 (N_14915,N_14624,N_14696);
nor U14916 (N_14916,N_14669,N_14589);
or U14917 (N_14917,N_14503,N_14722);
and U14918 (N_14918,N_14603,N_14665);
or U14919 (N_14919,N_14679,N_14675);
and U14920 (N_14920,N_14610,N_14633);
or U14921 (N_14921,N_14617,N_14619);
xnor U14922 (N_14922,N_14659,N_14547);
and U14923 (N_14923,N_14693,N_14515);
and U14924 (N_14924,N_14690,N_14730);
or U14925 (N_14925,N_14559,N_14601);
nor U14926 (N_14926,N_14577,N_14571);
nor U14927 (N_14927,N_14745,N_14646);
and U14928 (N_14928,N_14635,N_14571);
and U14929 (N_14929,N_14649,N_14535);
nor U14930 (N_14930,N_14693,N_14597);
nor U14931 (N_14931,N_14694,N_14636);
or U14932 (N_14932,N_14744,N_14559);
or U14933 (N_14933,N_14735,N_14665);
and U14934 (N_14934,N_14667,N_14525);
nand U14935 (N_14935,N_14525,N_14709);
or U14936 (N_14936,N_14678,N_14685);
and U14937 (N_14937,N_14686,N_14645);
nand U14938 (N_14938,N_14659,N_14711);
nor U14939 (N_14939,N_14643,N_14721);
or U14940 (N_14940,N_14749,N_14675);
nor U14941 (N_14941,N_14684,N_14601);
and U14942 (N_14942,N_14677,N_14575);
nand U14943 (N_14943,N_14620,N_14652);
and U14944 (N_14944,N_14655,N_14570);
nand U14945 (N_14945,N_14705,N_14546);
xor U14946 (N_14946,N_14711,N_14704);
and U14947 (N_14947,N_14542,N_14697);
or U14948 (N_14948,N_14672,N_14602);
xnor U14949 (N_14949,N_14626,N_14710);
nor U14950 (N_14950,N_14531,N_14565);
nor U14951 (N_14951,N_14510,N_14633);
nor U14952 (N_14952,N_14649,N_14546);
xnor U14953 (N_14953,N_14629,N_14507);
nor U14954 (N_14954,N_14650,N_14505);
nor U14955 (N_14955,N_14638,N_14689);
nor U14956 (N_14956,N_14560,N_14736);
and U14957 (N_14957,N_14569,N_14590);
and U14958 (N_14958,N_14748,N_14724);
or U14959 (N_14959,N_14730,N_14500);
or U14960 (N_14960,N_14544,N_14736);
or U14961 (N_14961,N_14592,N_14697);
nor U14962 (N_14962,N_14630,N_14540);
and U14963 (N_14963,N_14745,N_14618);
or U14964 (N_14964,N_14573,N_14621);
and U14965 (N_14965,N_14556,N_14615);
or U14966 (N_14966,N_14658,N_14651);
and U14967 (N_14967,N_14706,N_14519);
and U14968 (N_14968,N_14614,N_14610);
or U14969 (N_14969,N_14565,N_14619);
nand U14970 (N_14970,N_14607,N_14581);
xor U14971 (N_14971,N_14618,N_14708);
xnor U14972 (N_14972,N_14529,N_14725);
nand U14973 (N_14973,N_14574,N_14501);
xor U14974 (N_14974,N_14719,N_14534);
and U14975 (N_14975,N_14734,N_14556);
or U14976 (N_14976,N_14707,N_14543);
or U14977 (N_14977,N_14632,N_14741);
nand U14978 (N_14978,N_14544,N_14636);
nor U14979 (N_14979,N_14733,N_14716);
and U14980 (N_14980,N_14640,N_14600);
xor U14981 (N_14981,N_14576,N_14712);
xor U14982 (N_14982,N_14603,N_14673);
xor U14983 (N_14983,N_14747,N_14627);
or U14984 (N_14984,N_14545,N_14621);
or U14985 (N_14985,N_14703,N_14560);
nand U14986 (N_14986,N_14731,N_14708);
nand U14987 (N_14987,N_14653,N_14584);
and U14988 (N_14988,N_14534,N_14697);
and U14989 (N_14989,N_14536,N_14573);
or U14990 (N_14990,N_14640,N_14561);
nor U14991 (N_14991,N_14595,N_14633);
and U14992 (N_14992,N_14574,N_14504);
nor U14993 (N_14993,N_14677,N_14724);
nand U14994 (N_14994,N_14534,N_14607);
nor U14995 (N_14995,N_14536,N_14510);
and U14996 (N_14996,N_14695,N_14640);
nor U14997 (N_14997,N_14671,N_14632);
xor U14998 (N_14998,N_14735,N_14501);
nor U14999 (N_14999,N_14689,N_14683);
or U15000 (N_15000,N_14905,N_14894);
nor U15001 (N_15001,N_14795,N_14834);
nand U15002 (N_15002,N_14941,N_14986);
and U15003 (N_15003,N_14843,N_14818);
and U15004 (N_15004,N_14861,N_14985);
nor U15005 (N_15005,N_14934,N_14997);
or U15006 (N_15006,N_14767,N_14891);
and U15007 (N_15007,N_14946,N_14979);
or U15008 (N_15008,N_14824,N_14760);
nand U15009 (N_15009,N_14812,N_14860);
nor U15010 (N_15010,N_14902,N_14836);
and U15011 (N_15011,N_14810,N_14845);
nand U15012 (N_15012,N_14922,N_14947);
or U15013 (N_15013,N_14917,N_14775);
xor U15014 (N_15014,N_14859,N_14751);
nand U15015 (N_15015,N_14973,N_14950);
or U15016 (N_15016,N_14958,N_14821);
nand U15017 (N_15017,N_14808,N_14964);
and U15018 (N_15018,N_14753,N_14781);
nor U15019 (N_15019,N_14755,N_14980);
or U15020 (N_15020,N_14939,N_14960);
and U15021 (N_15021,N_14855,N_14884);
nor U15022 (N_15022,N_14995,N_14926);
nor U15023 (N_15023,N_14954,N_14910);
xor U15024 (N_15024,N_14952,N_14969);
nand U15025 (N_15025,N_14937,N_14813);
xor U15026 (N_15026,N_14970,N_14957);
xor U15027 (N_15027,N_14908,N_14907);
or U15028 (N_15028,N_14815,N_14787);
nand U15029 (N_15029,N_14779,N_14802);
nor U15030 (N_15030,N_14993,N_14768);
nor U15031 (N_15031,N_14974,N_14967);
nor U15032 (N_15032,N_14889,N_14992);
xnor U15033 (N_15033,N_14752,N_14971);
nor U15034 (N_15034,N_14948,N_14949);
nor U15035 (N_15035,N_14919,N_14975);
or U15036 (N_15036,N_14842,N_14841);
or U15037 (N_15037,N_14844,N_14772);
nand U15038 (N_15038,N_14887,N_14798);
xor U15039 (N_15039,N_14785,N_14858);
or U15040 (N_15040,N_14840,N_14763);
nand U15041 (N_15041,N_14929,N_14807);
nand U15042 (N_15042,N_14849,N_14953);
or U15043 (N_15043,N_14893,N_14942);
and U15044 (N_15044,N_14883,N_14898);
and U15045 (N_15045,N_14904,N_14863);
xnor U15046 (N_15046,N_14783,N_14959);
nand U15047 (N_15047,N_14984,N_14771);
nor U15048 (N_15048,N_14924,N_14761);
or U15049 (N_15049,N_14987,N_14923);
nor U15050 (N_15050,N_14820,N_14900);
or U15051 (N_15051,N_14892,N_14873);
and U15052 (N_15052,N_14876,N_14945);
xor U15053 (N_15053,N_14879,N_14872);
xor U15054 (N_15054,N_14912,N_14996);
xnor U15055 (N_15055,N_14827,N_14990);
nand U15056 (N_15056,N_14853,N_14822);
nand U15057 (N_15057,N_14916,N_14878);
nor U15058 (N_15058,N_14811,N_14799);
xnor U15059 (N_15059,N_14831,N_14773);
nand U15060 (N_15060,N_14899,N_14847);
nor U15061 (N_15061,N_14851,N_14870);
or U15062 (N_15062,N_14758,N_14852);
and U15063 (N_15063,N_14756,N_14790);
nand U15064 (N_15064,N_14956,N_14998);
xnor U15065 (N_15065,N_14774,N_14793);
nand U15066 (N_15066,N_14886,N_14982);
nor U15067 (N_15067,N_14875,N_14814);
and U15068 (N_15068,N_14911,N_14944);
xnor U15069 (N_15069,N_14806,N_14965);
nand U15070 (N_15070,N_14963,N_14750);
nand U15071 (N_15071,N_14867,N_14830);
nor U15072 (N_15072,N_14933,N_14931);
and U15073 (N_15073,N_14981,N_14961);
nand U15074 (N_15074,N_14936,N_14817);
nor U15075 (N_15075,N_14885,N_14782);
nor U15076 (N_15076,N_14826,N_14977);
xnor U15077 (N_15077,N_14951,N_14829);
or U15078 (N_15078,N_14932,N_14788);
or U15079 (N_15079,N_14809,N_14784);
and U15080 (N_15080,N_14994,N_14930);
nor U15081 (N_15081,N_14976,N_14777);
or U15082 (N_15082,N_14869,N_14819);
nand U15083 (N_15083,N_14918,N_14903);
and U15084 (N_15084,N_14914,N_14797);
and U15085 (N_15085,N_14759,N_14780);
and U15086 (N_15086,N_14943,N_14856);
and U15087 (N_15087,N_14915,N_14805);
nand U15088 (N_15088,N_14881,N_14989);
and U15089 (N_15089,N_14864,N_14764);
nand U15090 (N_15090,N_14833,N_14938);
nor U15091 (N_15091,N_14928,N_14823);
or U15092 (N_15092,N_14865,N_14972);
nand U15093 (N_15093,N_14882,N_14804);
nor U15094 (N_15094,N_14791,N_14897);
or U15095 (N_15095,N_14955,N_14801);
or U15096 (N_15096,N_14966,N_14757);
and U15097 (N_15097,N_14999,N_14800);
xor U15098 (N_15098,N_14754,N_14803);
nor U15099 (N_15099,N_14854,N_14837);
nor U15100 (N_15100,N_14848,N_14794);
nand U15101 (N_15101,N_14762,N_14906);
and U15102 (N_15102,N_14770,N_14839);
xor U15103 (N_15103,N_14789,N_14792);
and U15104 (N_15104,N_14935,N_14778);
nand U15105 (N_15105,N_14925,N_14927);
xnor U15106 (N_15106,N_14896,N_14838);
nor U15107 (N_15107,N_14765,N_14835);
xor U15108 (N_15108,N_14868,N_14962);
xor U15109 (N_15109,N_14940,N_14796);
and U15110 (N_15110,N_14909,N_14866);
nor U15111 (N_15111,N_14913,N_14862);
or U15112 (N_15112,N_14832,N_14786);
nor U15113 (N_15113,N_14816,N_14888);
and U15114 (N_15114,N_14850,N_14874);
nand U15115 (N_15115,N_14871,N_14988);
xor U15116 (N_15116,N_14769,N_14766);
nor U15117 (N_15117,N_14921,N_14890);
nand U15118 (N_15118,N_14983,N_14920);
and U15119 (N_15119,N_14776,N_14880);
or U15120 (N_15120,N_14978,N_14846);
nor U15121 (N_15121,N_14901,N_14828);
and U15122 (N_15122,N_14877,N_14968);
nand U15123 (N_15123,N_14825,N_14895);
xnor U15124 (N_15124,N_14857,N_14991);
or U15125 (N_15125,N_14897,N_14852);
or U15126 (N_15126,N_14960,N_14993);
nor U15127 (N_15127,N_14923,N_14901);
nand U15128 (N_15128,N_14954,N_14970);
nor U15129 (N_15129,N_14793,N_14900);
nor U15130 (N_15130,N_14779,N_14928);
and U15131 (N_15131,N_14802,N_14813);
nor U15132 (N_15132,N_14846,N_14913);
nand U15133 (N_15133,N_14875,N_14940);
xnor U15134 (N_15134,N_14843,N_14862);
nand U15135 (N_15135,N_14845,N_14907);
xnor U15136 (N_15136,N_14975,N_14773);
nor U15137 (N_15137,N_14977,N_14965);
nand U15138 (N_15138,N_14988,N_14879);
or U15139 (N_15139,N_14908,N_14763);
or U15140 (N_15140,N_14845,N_14858);
or U15141 (N_15141,N_14813,N_14892);
and U15142 (N_15142,N_14764,N_14871);
or U15143 (N_15143,N_14907,N_14869);
xor U15144 (N_15144,N_14944,N_14938);
xor U15145 (N_15145,N_14944,N_14934);
nor U15146 (N_15146,N_14859,N_14988);
nor U15147 (N_15147,N_14835,N_14794);
nor U15148 (N_15148,N_14783,N_14769);
nand U15149 (N_15149,N_14827,N_14776);
or U15150 (N_15150,N_14934,N_14921);
nor U15151 (N_15151,N_14999,N_14870);
nand U15152 (N_15152,N_14920,N_14925);
nand U15153 (N_15153,N_14867,N_14801);
nor U15154 (N_15154,N_14770,N_14780);
xnor U15155 (N_15155,N_14838,N_14879);
nor U15156 (N_15156,N_14976,N_14809);
nand U15157 (N_15157,N_14989,N_14968);
nand U15158 (N_15158,N_14806,N_14863);
xnor U15159 (N_15159,N_14969,N_14770);
xor U15160 (N_15160,N_14985,N_14919);
xnor U15161 (N_15161,N_14922,N_14869);
nor U15162 (N_15162,N_14790,N_14758);
and U15163 (N_15163,N_14828,N_14812);
nand U15164 (N_15164,N_14880,N_14909);
or U15165 (N_15165,N_14840,N_14990);
and U15166 (N_15166,N_14767,N_14905);
xor U15167 (N_15167,N_14787,N_14846);
or U15168 (N_15168,N_14841,N_14789);
xnor U15169 (N_15169,N_14948,N_14904);
nor U15170 (N_15170,N_14847,N_14799);
nor U15171 (N_15171,N_14797,N_14934);
nor U15172 (N_15172,N_14992,N_14857);
nand U15173 (N_15173,N_14786,N_14974);
and U15174 (N_15174,N_14884,N_14783);
nand U15175 (N_15175,N_14882,N_14965);
xnor U15176 (N_15176,N_14756,N_14872);
xor U15177 (N_15177,N_14754,N_14890);
nand U15178 (N_15178,N_14897,N_14803);
or U15179 (N_15179,N_14763,N_14947);
or U15180 (N_15180,N_14882,N_14897);
or U15181 (N_15181,N_14906,N_14807);
nand U15182 (N_15182,N_14814,N_14863);
or U15183 (N_15183,N_14785,N_14992);
xnor U15184 (N_15184,N_14957,N_14801);
nand U15185 (N_15185,N_14851,N_14845);
xor U15186 (N_15186,N_14964,N_14858);
or U15187 (N_15187,N_14871,N_14840);
and U15188 (N_15188,N_14952,N_14768);
and U15189 (N_15189,N_14859,N_14822);
xnor U15190 (N_15190,N_14939,N_14956);
nand U15191 (N_15191,N_14916,N_14853);
nor U15192 (N_15192,N_14886,N_14835);
xor U15193 (N_15193,N_14979,N_14770);
nor U15194 (N_15194,N_14799,N_14967);
and U15195 (N_15195,N_14786,N_14926);
and U15196 (N_15196,N_14875,N_14932);
or U15197 (N_15197,N_14814,N_14771);
xor U15198 (N_15198,N_14897,N_14865);
nor U15199 (N_15199,N_14925,N_14871);
nor U15200 (N_15200,N_14793,N_14977);
nand U15201 (N_15201,N_14861,N_14968);
and U15202 (N_15202,N_14951,N_14799);
xor U15203 (N_15203,N_14858,N_14890);
and U15204 (N_15204,N_14908,N_14926);
xnor U15205 (N_15205,N_14793,N_14989);
xnor U15206 (N_15206,N_14832,N_14800);
nand U15207 (N_15207,N_14768,N_14837);
nand U15208 (N_15208,N_14868,N_14950);
and U15209 (N_15209,N_14900,N_14944);
or U15210 (N_15210,N_14766,N_14795);
xor U15211 (N_15211,N_14886,N_14913);
xor U15212 (N_15212,N_14803,N_14896);
and U15213 (N_15213,N_14779,N_14980);
and U15214 (N_15214,N_14912,N_14898);
and U15215 (N_15215,N_14903,N_14885);
nand U15216 (N_15216,N_14963,N_14972);
xnor U15217 (N_15217,N_14796,N_14810);
nor U15218 (N_15218,N_14876,N_14916);
or U15219 (N_15219,N_14966,N_14975);
or U15220 (N_15220,N_14925,N_14827);
nor U15221 (N_15221,N_14987,N_14931);
nand U15222 (N_15222,N_14994,N_14972);
nand U15223 (N_15223,N_14777,N_14857);
xor U15224 (N_15224,N_14908,N_14871);
nor U15225 (N_15225,N_14796,N_14750);
or U15226 (N_15226,N_14852,N_14815);
xor U15227 (N_15227,N_14994,N_14773);
or U15228 (N_15228,N_14854,N_14772);
nor U15229 (N_15229,N_14838,N_14827);
nor U15230 (N_15230,N_14903,N_14853);
nor U15231 (N_15231,N_14879,N_14962);
nand U15232 (N_15232,N_14761,N_14864);
or U15233 (N_15233,N_14984,N_14950);
xnor U15234 (N_15234,N_14818,N_14906);
nor U15235 (N_15235,N_14790,N_14794);
and U15236 (N_15236,N_14992,N_14983);
xnor U15237 (N_15237,N_14911,N_14752);
and U15238 (N_15238,N_14802,N_14884);
nor U15239 (N_15239,N_14838,N_14864);
nor U15240 (N_15240,N_14965,N_14912);
or U15241 (N_15241,N_14843,N_14823);
nor U15242 (N_15242,N_14959,N_14990);
nand U15243 (N_15243,N_14805,N_14971);
or U15244 (N_15244,N_14784,N_14791);
or U15245 (N_15245,N_14837,N_14949);
xor U15246 (N_15246,N_14976,N_14877);
xnor U15247 (N_15247,N_14938,N_14789);
nand U15248 (N_15248,N_14855,N_14791);
nor U15249 (N_15249,N_14874,N_14768);
nand U15250 (N_15250,N_15204,N_15136);
or U15251 (N_15251,N_15225,N_15190);
xor U15252 (N_15252,N_15063,N_15202);
nand U15253 (N_15253,N_15167,N_15068);
and U15254 (N_15254,N_15232,N_15050);
and U15255 (N_15255,N_15193,N_15168);
or U15256 (N_15256,N_15183,N_15084);
nand U15257 (N_15257,N_15065,N_15201);
and U15258 (N_15258,N_15214,N_15109);
nor U15259 (N_15259,N_15011,N_15037);
nor U15260 (N_15260,N_15041,N_15161);
nand U15261 (N_15261,N_15110,N_15241);
nor U15262 (N_15262,N_15114,N_15036);
or U15263 (N_15263,N_15179,N_15249);
or U15264 (N_15264,N_15003,N_15053);
or U15265 (N_15265,N_15012,N_15196);
xor U15266 (N_15266,N_15197,N_15023);
nand U15267 (N_15267,N_15090,N_15020);
xor U15268 (N_15268,N_15058,N_15206);
or U15269 (N_15269,N_15205,N_15215);
and U15270 (N_15270,N_15240,N_15115);
xor U15271 (N_15271,N_15072,N_15075);
or U15272 (N_15272,N_15130,N_15047);
and U15273 (N_15273,N_15009,N_15247);
and U15274 (N_15274,N_15085,N_15242);
and U15275 (N_15275,N_15015,N_15106);
xor U15276 (N_15276,N_15028,N_15001);
and U15277 (N_15277,N_15024,N_15022);
and U15278 (N_15278,N_15119,N_15044);
xnor U15279 (N_15279,N_15010,N_15139);
nand U15280 (N_15280,N_15094,N_15078);
nor U15281 (N_15281,N_15025,N_15149);
and U15282 (N_15282,N_15019,N_15134);
nor U15283 (N_15283,N_15128,N_15112);
nor U15284 (N_15284,N_15228,N_15154);
xor U15285 (N_15285,N_15040,N_15016);
nand U15286 (N_15286,N_15049,N_15048);
nor U15287 (N_15287,N_15033,N_15055);
xor U15288 (N_15288,N_15234,N_15120);
or U15289 (N_15289,N_15054,N_15220);
nor U15290 (N_15290,N_15147,N_15081);
nand U15291 (N_15291,N_15144,N_15117);
nand U15292 (N_15292,N_15188,N_15164);
or U15293 (N_15293,N_15122,N_15180);
and U15294 (N_15294,N_15175,N_15069);
or U15295 (N_15295,N_15177,N_15199);
nand U15296 (N_15296,N_15231,N_15089);
nand U15297 (N_15297,N_15185,N_15108);
xor U15298 (N_15298,N_15039,N_15192);
xor U15299 (N_15299,N_15176,N_15006);
and U15300 (N_15300,N_15035,N_15145);
or U15301 (N_15301,N_15026,N_15057);
and U15302 (N_15302,N_15027,N_15098);
and U15303 (N_15303,N_15042,N_15034);
nand U15304 (N_15304,N_15248,N_15152);
and U15305 (N_15305,N_15123,N_15212);
and U15306 (N_15306,N_15159,N_15187);
or U15307 (N_15307,N_15173,N_15163);
nand U15308 (N_15308,N_15061,N_15194);
or U15309 (N_15309,N_15017,N_15138);
nand U15310 (N_15310,N_15153,N_15029);
and U15311 (N_15311,N_15079,N_15101);
xor U15312 (N_15312,N_15124,N_15107);
xnor U15313 (N_15313,N_15235,N_15021);
nand U15314 (N_15314,N_15046,N_15129);
nor U15315 (N_15315,N_15140,N_15002);
or U15316 (N_15316,N_15243,N_15246);
and U15317 (N_15317,N_15137,N_15142);
nor U15318 (N_15318,N_15051,N_15091);
or U15319 (N_15319,N_15071,N_15038);
nor U15320 (N_15320,N_15083,N_15174);
and U15321 (N_15321,N_15237,N_15062);
nor U15322 (N_15322,N_15158,N_15169);
xnor U15323 (N_15323,N_15171,N_15116);
or U15324 (N_15324,N_15076,N_15233);
and U15325 (N_15325,N_15151,N_15082);
xor U15326 (N_15326,N_15133,N_15184);
nand U15327 (N_15327,N_15067,N_15172);
xor U15328 (N_15328,N_15100,N_15077);
xor U15329 (N_15329,N_15096,N_15005);
or U15330 (N_15330,N_15236,N_15059);
xor U15331 (N_15331,N_15239,N_15229);
nand U15332 (N_15332,N_15103,N_15007);
nand U15333 (N_15333,N_15031,N_15238);
nor U15334 (N_15334,N_15030,N_15104);
or U15335 (N_15335,N_15143,N_15224);
or U15336 (N_15336,N_15052,N_15127);
nor U15337 (N_15337,N_15203,N_15073);
nor U15338 (N_15338,N_15198,N_15226);
or U15339 (N_15339,N_15157,N_15102);
xnor U15340 (N_15340,N_15219,N_15125);
or U15341 (N_15341,N_15191,N_15064);
xnor U15342 (N_15342,N_15111,N_15182);
nand U15343 (N_15343,N_15244,N_15221);
or U15344 (N_15344,N_15087,N_15018);
or U15345 (N_15345,N_15141,N_15216);
or U15346 (N_15346,N_15132,N_15146);
or U15347 (N_15347,N_15223,N_15209);
nor U15348 (N_15348,N_15135,N_15118);
and U15349 (N_15349,N_15060,N_15066);
nand U15350 (N_15350,N_15008,N_15166);
or U15351 (N_15351,N_15160,N_15099);
xor U15352 (N_15352,N_15043,N_15207);
nor U15353 (N_15353,N_15208,N_15165);
nor U15354 (N_15354,N_15162,N_15092);
and U15355 (N_15355,N_15056,N_15032);
nand U15356 (N_15356,N_15227,N_15245);
xnor U15357 (N_15357,N_15013,N_15150);
or U15358 (N_15358,N_15097,N_15222);
xor U15359 (N_15359,N_15113,N_15210);
xor U15360 (N_15360,N_15126,N_15088);
xor U15361 (N_15361,N_15200,N_15086);
or U15362 (N_15362,N_15080,N_15105);
nand U15363 (N_15363,N_15148,N_15195);
xor U15364 (N_15364,N_15045,N_15156);
or U15365 (N_15365,N_15213,N_15155);
or U15366 (N_15366,N_15189,N_15014);
nor U15367 (N_15367,N_15230,N_15178);
or U15368 (N_15368,N_15070,N_15121);
xor U15369 (N_15369,N_15218,N_15181);
nor U15370 (N_15370,N_15074,N_15095);
and U15371 (N_15371,N_15170,N_15093);
nor U15372 (N_15372,N_15211,N_15000);
nor U15373 (N_15373,N_15004,N_15217);
or U15374 (N_15374,N_15186,N_15131);
nand U15375 (N_15375,N_15228,N_15193);
and U15376 (N_15376,N_15082,N_15203);
nor U15377 (N_15377,N_15114,N_15179);
nor U15378 (N_15378,N_15195,N_15129);
nor U15379 (N_15379,N_15158,N_15117);
nor U15380 (N_15380,N_15211,N_15153);
or U15381 (N_15381,N_15062,N_15206);
xor U15382 (N_15382,N_15202,N_15091);
and U15383 (N_15383,N_15076,N_15071);
nor U15384 (N_15384,N_15074,N_15200);
nor U15385 (N_15385,N_15021,N_15166);
or U15386 (N_15386,N_15230,N_15133);
nand U15387 (N_15387,N_15082,N_15075);
nand U15388 (N_15388,N_15107,N_15224);
xnor U15389 (N_15389,N_15006,N_15190);
or U15390 (N_15390,N_15010,N_15119);
xor U15391 (N_15391,N_15110,N_15162);
nand U15392 (N_15392,N_15163,N_15084);
and U15393 (N_15393,N_15230,N_15160);
xnor U15394 (N_15394,N_15145,N_15210);
xor U15395 (N_15395,N_15124,N_15042);
xnor U15396 (N_15396,N_15230,N_15150);
nor U15397 (N_15397,N_15181,N_15000);
nor U15398 (N_15398,N_15135,N_15039);
xor U15399 (N_15399,N_15127,N_15159);
nor U15400 (N_15400,N_15239,N_15181);
nor U15401 (N_15401,N_15241,N_15122);
or U15402 (N_15402,N_15110,N_15127);
and U15403 (N_15403,N_15208,N_15089);
nor U15404 (N_15404,N_15034,N_15076);
nor U15405 (N_15405,N_15126,N_15080);
or U15406 (N_15406,N_15016,N_15174);
nor U15407 (N_15407,N_15196,N_15086);
nor U15408 (N_15408,N_15024,N_15236);
xor U15409 (N_15409,N_15002,N_15172);
or U15410 (N_15410,N_15115,N_15220);
nor U15411 (N_15411,N_15128,N_15101);
nand U15412 (N_15412,N_15027,N_15210);
nor U15413 (N_15413,N_15195,N_15051);
and U15414 (N_15414,N_15046,N_15199);
nor U15415 (N_15415,N_15220,N_15004);
xnor U15416 (N_15416,N_15065,N_15238);
and U15417 (N_15417,N_15147,N_15046);
nor U15418 (N_15418,N_15138,N_15038);
xor U15419 (N_15419,N_15228,N_15215);
nand U15420 (N_15420,N_15151,N_15109);
xnor U15421 (N_15421,N_15030,N_15031);
and U15422 (N_15422,N_15121,N_15068);
xor U15423 (N_15423,N_15049,N_15126);
xor U15424 (N_15424,N_15171,N_15167);
nand U15425 (N_15425,N_15049,N_15233);
xnor U15426 (N_15426,N_15092,N_15170);
nand U15427 (N_15427,N_15182,N_15035);
nand U15428 (N_15428,N_15103,N_15183);
xnor U15429 (N_15429,N_15061,N_15111);
and U15430 (N_15430,N_15172,N_15205);
xor U15431 (N_15431,N_15142,N_15242);
nand U15432 (N_15432,N_15175,N_15184);
nand U15433 (N_15433,N_15183,N_15203);
xor U15434 (N_15434,N_15248,N_15044);
or U15435 (N_15435,N_15177,N_15236);
nand U15436 (N_15436,N_15005,N_15207);
xnor U15437 (N_15437,N_15140,N_15047);
or U15438 (N_15438,N_15220,N_15131);
or U15439 (N_15439,N_15106,N_15184);
nand U15440 (N_15440,N_15001,N_15024);
nand U15441 (N_15441,N_15100,N_15037);
and U15442 (N_15442,N_15079,N_15233);
nand U15443 (N_15443,N_15123,N_15160);
nor U15444 (N_15444,N_15134,N_15039);
and U15445 (N_15445,N_15233,N_15064);
nand U15446 (N_15446,N_15031,N_15089);
xor U15447 (N_15447,N_15048,N_15091);
or U15448 (N_15448,N_15144,N_15169);
and U15449 (N_15449,N_15221,N_15024);
nor U15450 (N_15450,N_15089,N_15079);
nand U15451 (N_15451,N_15022,N_15153);
and U15452 (N_15452,N_15109,N_15030);
nand U15453 (N_15453,N_15150,N_15000);
xor U15454 (N_15454,N_15142,N_15114);
nand U15455 (N_15455,N_15061,N_15169);
nor U15456 (N_15456,N_15095,N_15166);
or U15457 (N_15457,N_15170,N_15065);
nor U15458 (N_15458,N_15022,N_15158);
xnor U15459 (N_15459,N_15032,N_15055);
nand U15460 (N_15460,N_15154,N_15051);
nand U15461 (N_15461,N_15011,N_15023);
or U15462 (N_15462,N_15181,N_15071);
nand U15463 (N_15463,N_15245,N_15158);
nand U15464 (N_15464,N_15026,N_15229);
nand U15465 (N_15465,N_15060,N_15163);
xnor U15466 (N_15466,N_15048,N_15008);
and U15467 (N_15467,N_15152,N_15237);
xnor U15468 (N_15468,N_15082,N_15035);
or U15469 (N_15469,N_15249,N_15122);
and U15470 (N_15470,N_15130,N_15040);
and U15471 (N_15471,N_15194,N_15128);
or U15472 (N_15472,N_15240,N_15105);
and U15473 (N_15473,N_15217,N_15005);
or U15474 (N_15474,N_15027,N_15139);
xnor U15475 (N_15475,N_15119,N_15208);
or U15476 (N_15476,N_15059,N_15044);
nand U15477 (N_15477,N_15158,N_15043);
and U15478 (N_15478,N_15071,N_15184);
nor U15479 (N_15479,N_15099,N_15110);
nand U15480 (N_15480,N_15139,N_15186);
and U15481 (N_15481,N_15074,N_15154);
xnor U15482 (N_15482,N_15018,N_15185);
and U15483 (N_15483,N_15117,N_15080);
or U15484 (N_15484,N_15111,N_15007);
xor U15485 (N_15485,N_15056,N_15113);
nor U15486 (N_15486,N_15179,N_15074);
xnor U15487 (N_15487,N_15009,N_15023);
and U15488 (N_15488,N_15151,N_15150);
or U15489 (N_15489,N_15023,N_15028);
nand U15490 (N_15490,N_15245,N_15018);
or U15491 (N_15491,N_15055,N_15072);
and U15492 (N_15492,N_15074,N_15033);
and U15493 (N_15493,N_15126,N_15144);
nor U15494 (N_15494,N_15188,N_15075);
or U15495 (N_15495,N_15039,N_15027);
nand U15496 (N_15496,N_15145,N_15225);
nand U15497 (N_15497,N_15061,N_15248);
nand U15498 (N_15498,N_15082,N_15055);
or U15499 (N_15499,N_15150,N_15192);
and U15500 (N_15500,N_15465,N_15410);
nor U15501 (N_15501,N_15384,N_15342);
xnor U15502 (N_15502,N_15413,N_15320);
nor U15503 (N_15503,N_15253,N_15314);
xor U15504 (N_15504,N_15363,N_15414);
and U15505 (N_15505,N_15458,N_15310);
nor U15506 (N_15506,N_15294,N_15438);
xnor U15507 (N_15507,N_15443,N_15255);
nand U15508 (N_15508,N_15337,N_15276);
or U15509 (N_15509,N_15453,N_15386);
and U15510 (N_15510,N_15457,N_15358);
and U15511 (N_15511,N_15442,N_15390);
and U15512 (N_15512,N_15370,N_15365);
nand U15513 (N_15513,N_15331,N_15425);
or U15514 (N_15514,N_15389,N_15278);
nor U15515 (N_15515,N_15251,N_15270);
xor U15516 (N_15516,N_15351,N_15329);
nand U15517 (N_15517,N_15494,N_15355);
nor U15518 (N_15518,N_15266,N_15480);
nand U15519 (N_15519,N_15293,N_15466);
xor U15520 (N_15520,N_15268,N_15335);
nand U15521 (N_15521,N_15327,N_15429);
nor U15522 (N_15522,N_15419,N_15279);
or U15523 (N_15523,N_15256,N_15492);
nor U15524 (N_15524,N_15322,N_15452);
and U15525 (N_15525,N_15372,N_15393);
nor U15526 (N_15526,N_15269,N_15485);
xnor U15527 (N_15527,N_15397,N_15490);
nor U15528 (N_15528,N_15292,N_15489);
nand U15529 (N_15529,N_15343,N_15291);
or U15530 (N_15530,N_15298,N_15282);
nor U15531 (N_15531,N_15339,N_15347);
nor U15532 (N_15532,N_15395,N_15421);
and U15533 (N_15533,N_15454,N_15496);
nor U15534 (N_15534,N_15433,N_15262);
nor U15535 (N_15535,N_15368,N_15328);
nand U15536 (N_15536,N_15264,N_15426);
nor U15537 (N_15537,N_15261,N_15402);
nor U15538 (N_15538,N_15472,N_15283);
and U15539 (N_15539,N_15364,N_15290);
nand U15540 (N_15540,N_15271,N_15306);
or U15541 (N_15541,N_15478,N_15275);
or U15542 (N_15542,N_15378,N_15341);
xnor U15543 (N_15543,N_15318,N_15469);
or U15544 (N_15544,N_15313,N_15354);
or U15545 (N_15545,N_15493,N_15317);
nor U15546 (N_15546,N_15312,N_15332);
nand U15547 (N_15547,N_15444,N_15422);
nor U15548 (N_15548,N_15250,N_15445);
nor U15549 (N_15549,N_15399,N_15359);
nor U15550 (N_15550,N_15280,N_15449);
xor U15551 (N_15551,N_15477,N_15455);
nand U15552 (N_15552,N_15420,N_15288);
nor U15553 (N_15553,N_15416,N_15428);
nor U15554 (N_15554,N_15304,N_15481);
nand U15555 (N_15555,N_15473,N_15305);
and U15556 (N_15556,N_15299,N_15408);
and U15557 (N_15557,N_15324,N_15498);
and U15558 (N_15558,N_15349,N_15285);
or U15559 (N_15559,N_15450,N_15303);
and U15560 (N_15560,N_15432,N_15391);
xor U15561 (N_15561,N_15350,N_15259);
nor U15562 (N_15562,N_15487,N_15418);
and U15563 (N_15563,N_15441,N_15330);
or U15564 (N_15564,N_15459,N_15281);
xnor U15565 (N_15565,N_15286,N_15417);
and U15566 (N_15566,N_15265,N_15315);
nor U15567 (N_15567,N_15474,N_15321);
nand U15568 (N_15568,N_15439,N_15333);
and U15569 (N_15569,N_15382,N_15289);
nand U15570 (N_15570,N_15352,N_15277);
and U15571 (N_15571,N_15468,N_15369);
and U15572 (N_15572,N_15375,N_15260);
nor U15573 (N_15573,N_15302,N_15464);
nand U15574 (N_15574,N_15486,N_15427);
and U15575 (N_15575,N_15373,N_15470);
and U15576 (N_15576,N_15311,N_15398);
and U15577 (N_15577,N_15360,N_15404);
nor U15578 (N_15578,N_15499,N_15267);
and U15579 (N_15579,N_15462,N_15258);
or U15580 (N_15580,N_15379,N_15476);
xnor U15581 (N_15581,N_15345,N_15254);
xnor U15582 (N_15582,N_15273,N_15407);
or U15583 (N_15583,N_15353,N_15301);
or U15584 (N_15584,N_15388,N_15415);
and U15585 (N_15585,N_15396,N_15257);
nor U15586 (N_15586,N_15463,N_15309);
nand U15587 (N_15587,N_15479,N_15381);
nand U15588 (N_15588,N_15387,N_15401);
xnor U15589 (N_15589,N_15340,N_15471);
and U15590 (N_15590,N_15252,N_15263);
xnor U15591 (N_15591,N_15300,N_15497);
nand U15592 (N_15592,N_15274,N_15316);
nand U15593 (N_15593,N_15380,N_15326);
nand U15594 (N_15594,N_15475,N_15287);
or U15595 (N_15595,N_15367,N_15295);
xor U15596 (N_15596,N_15334,N_15371);
and U15597 (N_15597,N_15406,N_15431);
xor U15598 (N_15598,N_15376,N_15361);
nor U15599 (N_15599,N_15356,N_15284);
nand U15600 (N_15600,N_15346,N_15403);
xor U15601 (N_15601,N_15400,N_15483);
or U15602 (N_15602,N_15484,N_15467);
nand U15603 (N_15603,N_15392,N_15446);
and U15604 (N_15604,N_15366,N_15362);
nor U15605 (N_15605,N_15461,N_15411);
nor U15606 (N_15606,N_15383,N_15434);
and U15607 (N_15607,N_15436,N_15272);
nor U15608 (N_15608,N_15385,N_15377);
and U15609 (N_15609,N_15308,N_15409);
or U15610 (N_15610,N_15348,N_15336);
and U15611 (N_15611,N_15325,N_15338);
nor U15612 (N_15612,N_15488,N_15435);
or U15613 (N_15613,N_15448,N_15447);
xor U15614 (N_15614,N_15491,N_15451);
or U15615 (N_15615,N_15482,N_15405);
nor U15616 (N_15616,N_15297,N_15495);
and U15617 (N_15617,N_15307,N_15319);
nor U15618 (N_15618,N_15430,N_15357);
or U15619 (N_15619,N_15456,N_15374);
or U15620 (N_15620,N_15460,N_15423);
and U15621 (N_15621,N_15424,N_15440);
nor U15622 (N_15622,N_15394,N_15344);
or U15623 (N_15623,N_15323,N_15412);
or U15624 (N_15624,N_15296,N_15437);
nand U15625 (N_15625,N_15435,N_15336);
nand U15626 (N_15626,N_15285,N_15398);
nand U15627 (N_15627,N_15360,N_15486);
or U15628 (N_15628,N_15336,N_15319);
or U15629 (N_15629,N_15470,N_15462);
xor U15630 (N_15630,N_15287,N_15250);
or U15631 (N_15631,N_15314,N_15383);
nand U15632 (N_15632,N_15438,N_15387);
xnor U15633 (N_15633,N_15445,N_15458);
nand U15634 (N_15634,N_15326,N_15344);
nor U15635 (N_15635,N_15439,N_15342);
or U15636 (N_15636,N_15475,N_15410);
and U15637 (N_15637,N_15371,N_15470);
xnor U15638 (N_15638,N_15290,N_15356);
xor U15639 (N_15639,N_15413,N_15360);
nand U15640 (N_15640,N_15340,N_15441);
xor U15641 (N_15641,N_15325,N_15406);
nor U15642 (N_15642,N_15295,N_15481);
xnor U15643 (N_15643,N_15498,N_15400);
nand U15644 (N_15644,N_15443,N_15335);
xnor U15645 (N_15645,N_15388,N_15414);
or U15646 (N_15646,N_15293,N_15369);
nor U15647 (N_15647,N_15414,N_15373);
and U15648 (N_15648,N_15494,N_15419);
nand U15649 (N_15649,N_15452,N_15266);
xor U15650 (N_15650,N_15309,N_15289);
nor U15651 (N_15651,N_15493,N_15429);
or U15652 (N_15652,N_15428,N_15356);
nand U15653 (N_15653,N_15470,N_15318);
or U15654 (N_15654,N_15401,N_15424);
nand U15655 (N_15655,N_15376,N_15489);
xor U15656 (N_15656,N_15398,N_15250);
and U15657 (N_15657,N_15290,N_15450);
nor U15658 (N_15658,N_15488,N_15353);
nor U15659 (N_15659,N_15380,N_15279);
and U15660 (N_15660,N_15410,N_15473);
nand U15661 (N_15661,N_15457,N_15335);
and U15662 (N_15662,N_15433,N_15296);
or U15663 (N_15663,N_15300,N_15284);
or U15664 (N_15664,N_15417,N_15261);
and U15665 (N_15665,N_15406,N_15316);
or U15666 (N_15666,N_15437,N_15357);
or U15667 (N_15667,N_15278,N_15367);
xor U15668 (N_15668,N_15417,N_15407);
or U15669 (N_15669,N_15290,N_15427);
nor U15670 (N_15670,N_15319,N_15343);
and U15671 (N_15671,N_15285,N_15450);
and U15672 (N_15672,N_15391,N_15499);
nor U15673 (N_15673,N_15276,N_15301);
or U15674 (N_15674,N_15455,N_15452);
nor U15675 (N_15675,N_15400,N_15429);
xnor U15676 (N_15676,N_15487,N_15346);
or U15677 (N_15677,N_15328,N_15397);
and U15678 (N_15678,N_15402,N_15355);
xor U15679 (N_15679,N_15432,N_15251);
or U15680 (N_15680,N_15488,N_15335);
and U15681 (N_15681,N_15331,N_15260);
and U15682 (N_15682,N_15458,N_15273);
nand U15683 (N_15683,N_15351,N_15480);
xor U15684 (N_15684,N_15390,N_15432);
or U15685 (N_15685,N_15433,N_15467);
xor U15686 (N_15686,N_15401,N_15314);
xor U15687 (N_15687,N_15488,N_15377);
or U15688 (N_15688,N_15466,N_15321);
nand U15689 (N_15689,N_15278,N_15260);
nand U15690 (N_15690,N_15463,N_15451);
nand U15691 (N_15691,N_15278,N_15286);
nor U15692 (N_15692,N_15345,N_15376);
nor U15693 (N_15693,N_15288,N_15372);
and U15694 (N_15694,N_15312,N_15377);
xnor U15695 (N_15695,N_15274,N_15381);
and U15696 (N_15696,N_15343,N_15440);
nor U15697 (N_15697,N_15400,N_15386);
xnor U15698 (N_15698,N_15403,N_15316);
and U15699 (N_15699,N_15346,N_15310);
and U15700 (N_15700,N_15250,N_15494);
nor U15701 (N_15701,N_15357,N_15395);
nand U15702 (N_15702,N_15261,N_15251);
and U15703 (N_15703,N_15292,N_15275);
nor U15704 (N_15704,N_15286,N_15416);
or U15705 (N_15705,N_15389,N_15290);
nand U15706 (N_15706,N_15256,N_15493);
nand U15707 (N_15707,N_15486,N_15315);
or U15708 (N_15708,N_15306,N_15279);
xor U15709 (N_15709,N_15325,N_15396);
nor U15710 (N_15710,N_15479,N_15412);
xnor U15711 (N_15711,N_15456,N_15356);
xnor U15712 (N_15712,N_15481,N_15261);
nor U15713 (N_15713,N_15383,N_15373);
and U15714 (N_15714,N_15461,N_15344);
or U15715 (N_15715,N_15377,N_15434);
or U15716 (N_15716,N_15270,N_15312);
and U15717 (N_15717,N_15421,N_15326);
nand U15718 (N_15718,N_15313,N_15346);
nor U15719 (N_15719,N_15436,N_15369);
and U15720 (N_15720,N_15434,N_15301);
or U15721 (N_15721,N_15303,N_15322);
nor U15722 (N_15722,N_15491,N_15257);
nor U15723 (N_15723,N_15347,N_15366);
nor U15724 (N_15724,N_15461,N_15474);
or U15725 (N_15725,N_15356,N_15409);
xor U15726 (N_15726,N_15333,N_15408);
or U15727 (N_15727,N_15319,N_15438);
or U15728 (N_15728,N_15277,N_15440);
nand U15729 (N_15729,N_15421,N_15411);
nor U15730 (N_15730,N_15393,N_15327);
xnor U15731 (N_15731,N_15416,N_15493);
and U15732 (N_15732,N_15475,N_15290);
nor U15733 (N_15733,N_15256,N_15393);
xnor U15734 (N_15734,N_15322,N_15384);
and U15735 (N_15735,N_15320,N_15368);
nand U15736 (N_15736,N_15457,N_15294);
or U15737 (N_15737,N_15389,N_15492);
nand U15738 (N_15738,N_15465,N_15369);
xnor U15739 (N_15739,N_15431,N_15320);
and U15740 (N_15740,N_15498,N_15372);
or U15741 (N_15741,N_15402,N_15264);
nand U15742 (N_15742,N_15458,N_15496);
and U15743 (N_15743,N_15378,N_15474);
xnor U15744 (N_15744,N_15468,N_15415);
or U15745 (N_15745,N_15498,N_15454);
nand U15746 (N_15746,N_15499,N_15304);
nor U15747 (N_15747,N_15438,N_15275);
nand U15748 (N_15748,N_15421,N_15262);
and U15749 (N_15749,N_15370,N_15466);
or U15750 (N_15750,N_15680,N_15565);
xnor U15751 (N_15751,N_15587,N_15664);
and U15752 (N_15752,N_15700,N_15655);
nor U15753 (N_15753,N_15528,N_15682);
or U15754 (N_15754,N_15585,N_15639);
nor U15755 (N_15755,N_15558,N_15714);
nor U15756 (N_15756,N_15689,N_15578);
xor U15757 (N_15757,N_15582,N_15660);
nor U15758 (N_15758,N_15686,N_15509);
xor U15759 (N_15759,N_15525,N_15653);
and U15760 (N_15760,N_15707,N_15600);
nand U15761 (N_15761,N_15554,N_15531);
or U15762 (N_15762,N_15698,N_15599);
nand U15763 (N_15763,N_15575,N_15584);
and U15764 (N_15764,N_15651,N_15515);
nor U15765 (N_15765,N_15577,N_15538);
and U15766 (N_15766,N_15597,N_15697);
nor U15767 (N_15767,N_15734,N_15636);
xnor U15768 (N_15768,N_15716,N_15556);
or U15769 (N_15769,N_15654,N_15625);
nand U15770 (N_15770,N_15683,N_15648);
and U15771 (N_15771,N_15665,N_15541);
and U15772 (N_15772,N_15604,N_15504);
and U15773 (N_15773,N_15657,N_15720);
or U15774 (N_15774,N_15743,N_15562);
or U15775 (N_15775,N_15514,N_15696);
and U15776 (N_15776,N_15638,N_15679);
or U15777 (N_15777,N_15678,N_15540);
and U15778 (N_15778,N_15711,N_15631);
nand U15779 (N_15779,N_15737,N_15746);
and U15780 (N_15780,N_15559,N_15690);
xnor U15781 (N_15781,N_15548,N_15503);
and U15782 (N_15782,N_15622,N_15675);
or U15783 (N_15783,N_15693,N_15641);
or U15784 (N_15784,N_15742,N_15672);
xnor U15785 (N_15785,N_15703,N_15522);
xnor U15786 (N_15786,N_15702,N_15581);
xor U15787 (N_15787,N_15688,N_15603);
nor U15788 (N_15788,N_15573,N_15637);
nor U15789 (N_15789,N_15727,N_15738);
and U15790 (N_15790,N_15586,N_15607);
xnor U15791 (N_15791,N_15701,N_15687);
nor U15792 (N_15792,N_15535,N_15719);
or U15793 (N_15793,N_15721,N_15588);
or U15794 (N_15794,N_15695,N_15523);
or U15795 (N_15795,N_15744,N_15512);
xor U15796 (N_15796,N_15506,N_15671);
nand U15797 (N_15797,N_15644,N_15574);
and U15798 (N_15798,N_15609,N_15610);
nor U15799 (N_15799,N_15659,N_15534);
xnor U15800 (N_15800,N_15708,N_15666);
nor U15801 (N_15801,N_15567,N_15723);
or U15802 (N_15802,N_15537,N_15741);
nor U15803 (N_15803,N_15544,N_15634);
nand U15804 (N_15804,N_15736,N_15517);
or U15805 (N_15805,N_15533,N_15612);
xor U15806 (N_15806,N_15501,N_15685);
xor U15807 (N_15807,N_15557,N_15626);
nand U15808 (N_15808,N_15589,N_15623);
nor U15809 (N_15809,N_15550,N_15661);
nand U15810 (N_15810,N_15621,N_15619);
or U15811 (N_15811,N_15731,N_15553);
nand U15812 (N_15812,N_15520,N_15510);
nor U15813 (N_15813,N_15642,N_15705);
nor U15814 (N_15814,N_15618,N_15712);
and U15815 (N_15815,N_15532,N_15605);
and U15816 (N_15816,N_15594,N_15724);
and U15817 (N_15817,N_15593,N_15595);
and U15818 (N_15818,N_15722,N_15733);
nand U15819 (N_15819,N_15627,N_15704);
nor U15820 (N_15820,N_15674,N_15692);
and U15821 (N_15821,N_15606,N_15576);
or U15822 (N_15822,N_15662,N_15563);
nor U15823 (N_15823,N_15656,N_15635);
xnor U15824 (N_15824,N_15616,N_15564);
nand U15825 (N_15825,N_15668,N_15518);
nand U15826 (N_15826,N_15749,N_15524);
or U15827 (N_15827,N_15545,N_15740);
xnor U15828 (N_15828,N_15725,N_15650);
and U15829 (N_15829,N_15511,N_15658);
xor U15830 (N_15830,N_15519,N_15728);
nor U15831 (N_15831,N_15630,N_15526);
or U15832 (N_15832,N_15560,N_15583);
nor U15833 (N_15833,N_15676,N_15549);
nor U15834 (N_15834,N_15516,N_15633);
or U15835 (N_15835,N_15670,N_15713);
nor U15836 (N_15836,N_15669,N_15645);
and U15837 (N_15837,N_15543,N_15569);
or U15838 (N_15838,N_15566,N_15748);
nand U15839 (N_15839,N_15629,N_15555);
or U15840 (N_15840,N_15632,N_15717);
and U15841 (N_15841,N_15551,N_15694);
nand U15842 (N_15842,N_15505,N_15570);
nand U15843 (N_15843,N_15691,N_15614);
nand U15844 (N_15844,N_15580,N_15590);
nand U15845 (N_15845,N_15611,N_15527);
nor U15846 (N_15846,N_15718,N_15715);
nor U15847 (N_15847,N_15732,N_15649);
nor U15848 (N_15848,N_15539,N_15730);
and U15849 (N_15849,N_15530,N_15521);
or U15850 (N_15850,N_15529,N_15613);
and U15851 (N_15851,N_15739,N_15568);
xor U15852 (N_15852,N_15647,N_15640);
xor U15853 (N_15853,N_15507,N_15536);
xor U15854 (N_15854,N_15673,N_15500);
xnor U15855 (N_15855,N_15684,N_15546);
nor U15856 (N_15856,N_15572,N_15601);
nand U15857 (N_15857,N_15735,N_15747);
nor U15858 (N_15858,N_15579,N_15726);
xnor U15859 (N_15859,N_15596,N_15552);
nand U15860 (N_15860,N_15620,N_15561);
xor U15861 (N_15861,N_15542,N_15643);
xor U15862 (N_15862,N_15628,N_15591);
and U15863 (N_15863,N_15709,N_15681);
and U15864 (N_15864,N_15745,N_15615);
nand U15865 (N_15865,N_15663,N_15699);
or U15866 (N_15866,N_15513,N_15508);
nand U15867 (N_15867,N_15652,N_15502);
and U15868 (N_15868,N_15598,N_15624);
and U15869 (N_15869,N_15617,N_15729);
nand U15870 (N_15870,N_15571,N_15592);
or U15871 (N_15871,N_15602,N_15677);
or U15872 (N_15872,N_15667,N_15710);
or U15873 (N_15873,N_15608,N_15547);
xnor U15874 (N_15874,N_15646,N_15706);
or U15875 (N_15875,N_15529,N_15565);
and U15876 (N_15876,N_15729,N_15748);
nor U15877 (N_15877,N_15628,N_15729);
nor U15878 (N_15878,N_15529,N_15556);
or U15879 (N_15879,N_15665,N_15738);
nor U15880 (N_15880,N_15580,N_15714);
xnor U15881 (N_15881,N_15702,N_15677);
or U15882 (N_15882,N_15629,N_15519);
nor U15883 (N_15883,N_15546,N_15522);
and U15884 (N_15884,N_15710,N_15503);
and U15885 (N_15885,N_15729,N_15648);
and U15886 (N_15886,N_15679,N_15670);
xnor U15887 (N_15887,N_15566,N_15602);
nand U15888 (N_15888,N_15538,N_15724);
nor U15889 (N_15889,N_15704,N_15608);
or U15890 (N_15890,N_15595,N_15687);
nor U15891 (N_15891,N_15533,N_15746);
or U15892 (N_15892,N_15715,N_15665);
nor U15893 (N_15893,N_15709,N_15739);
or U15894 (N_15894,N_15679,N_15693);
nand U15895 (N_15895,N_15628,N_15502);
and U15896 (N_15896,N_15656,N_15690);
and U15897 (N_15897,N_15541,N_15747);
nor U15898 (N_15898,N_15589,N_15695);
nand U15899 (N_15899,N_15729,N_15636);
and U15900 (N_15900,N_15630,N_15560);
xnor U15901 (N_15901,N_15731,N_15635);
nor U15902 (N_15902,N_15738,N_15549);
or U15903 (N_15903,N_15526,N_15568);
or U15904 (N_15904,N_15642,N_15665);
xor U15905 (N_15905,N_15741,N_15707);
or U15906 (N_15906,N_15515,N_15612);
and U15907 (N_15907,N_15632,N_15638);
and U15908 (N_15908,N_15511,N_15546);
xnor U15909 (N_15909,N_15627,N_15657);
nand U15910 (N_15910,N_15614,N_15506);
xor U15911 (N_15911,N_15735,N_15578);
nand U15912 (N_15912,N_15714,N_15566);
or U15913 (N_15913,N_15599,N_15725);
or U15914 (N_15914,N_15508,N_15536);
or U15915 (N_15915,N_15741,N_15611);
xnor U15916 (N_15916,N_15649,N_15689);
and U15917 (N_15917,N_15629,N_15593);
nor U15918 (N_15918,N_15521,N_15507);
nor U15919 (N_15919,N_15634,N_15622);
and U15920 (N_15920,N_15656,N_15566);
and U15921 (N_15921,N_15670,N_15533);
or U15922 (N_15922,N_15645,N_15741);
xnor U15923 (N_15923,N_15525,N_15599);
xnor U15924 (N_15924,N_15723,N_15683);
nand U15925 (N_15925,N_15655,N_15631);
and U15926 (N_15926,N_15710,N_15664);
nor U15927 (N_15927,N_15542,N_15728);
or U15928 (N_15928,N_15549,N_15705);
and U15929 (N_15929,N_15677,N_15645);
nand U15930 (N_15930,N_15530,N_15663);
and U15931 (N_15931,N_15747,N_15576);
xnor U15932 (N_15932,N_15614,N_15746);
xnor U15933 (N_15933,N_15689,N_15703);
nand U15934 (N_15934,N_15600,N_15523);
or U15935 (N_15935,N_15616,N_15688);
nor U15936 (N_15936,N_15668,N_15617);
xnor U15937 (N_15937,N_15626,N_15620);
and U15938 (N_15938,N_15694,N_15657);
nand U15939 (N_15939,N_15535,N_15558);
nand U15940 (N_15940,N_15662,N_15697);
nand U15941 (N_15941,N_15740,N_15615);
xnor U15942 (N_15942,N_15523,N_15661);
nand U15943 (N_15943,N_15599,N_15685);
or U15944 (N_15944,N_15723,N_15504);
nand U15945 (N_15945,N_15541,N_15629);
nor U15946 (N_15946,N_15520,N_15664);
or U15947 (N_15947,N_15574,N_15599);
nand U15948 (N_15948,N_15562,N_15605);
nor U15949 (N_15949,N_15552,N_15537);
nand U15950 (N_15950,N_15735,N_15658);
nor U15951 (N_15951,N_15591,N_15710);
or U15952 (N_15952,N_15513,N_15568);
and U15953 (N_15953,N_15705,N_15588);
and U15954 (N_15954,N_15501,N_15627);
or U15955 (N_15955,N_15717,N_15578);
or U15956 (N_15956,N_15617,N_15589);
or U15957 (N_15957,N_15566,N_15512);
nor U15958 (N_15958,N_15521,N_15600);
xor U15959 (N_15959,N_15562,N_15530);
xor U15960 (N_15960,N_15669,N_15703);
nor U15961 (N_15961,N_15563,N_15620);
or U15962 (N_15962,N_15726,N_15606);
and U15963 (N_15963,N_15609,N_15531);
xor U15964 (N_15964,N_15545,N_15543);
nor U15965 (N_15965,N_15741,N_15691);
and U15966 (N_15966,N_15633,N_15535);
nor U15967 (N_15967,N_15509,N_15640);
nor U15968 (N_15968,N_15571,N_15674);
nor U15969 (N_15969,N_15693,N_15682);
nand U15970 (N_15970,N_15525,N_15605);
or U15971 (N_15971,N_15746,N_15605);
nor U15972 (N_15972,N_15690,N_15744);
and U15973 (N_15973,N_15683,N_15700);
or U15974 (N_15974,N_15701,N_15673);
xnor U15975 (N_15975,N_15581,N_15591);
xnor U15976 (N_15976,N_15591,N_15519);
or U15977 (N_15977,N_15586,N_15529);
nand U15978 (N_15978,N_15722,N_15636);
nand U15979 (N_15979,N_15625,N_15621);
and U15980 (N_15980,N_15609,N_15744);
and U15981 (N_15981,N_15536,N_15747);
or U15982 (N_15982,N_15537,N_15716);
nand U15983 (N_15983,N_15584,N_15526);
xnor U15984 (N_15984,N_15556,N_15690);
xnor U15985 (N_15985,N_15703,N_15739);
and U15986 (N_15986,N_15679,N_15558);
nor U15987 (N_15987,N_15554,N_15503);
nand U15988 (N_15988,N_15530,N_15692);
xnor U15989 (N_15989,N_15588,N_15581);
nor U15990 (N_15990,N_15739,N_15593);
xor U15991 (N_15991,N_15522,N_15635);
nor U15992 (N_15992,N_15594,N_15670);
nand U15993 (N_15993,N_15726,N_15723);
nand U15994 (N_15994,N_15712,N_15542);
nor U15995 (N_15995,N_15546,N_15611);
xor U15996 (N_15996,N_15658,N_15725);
or U15997 (N_15997,N_15722,N_15676);
nor U15998 (N_15998,N_15674,N_15618);
and U15999 (N_15999,N_15642,N_15613);
and U16000 (N_16000,N_15819,N_15757);
xor U16001 (N_16001,N_15870,N_15924);
nor U16002 (N_16002,N_15808,N_15814);
nor U16003 (N_16003,N_15973,N_15985);
nor U16004 (N_16004,N_15824,N_15959);
and U16005 (N_16005,N_15986,N_15892);
nand U16006 (N_16006,N_15917,N_15775);
nor U16007 (N_16007,N_15825,N_15899);
nand U16008 (N_16008,N_15881,N_15956);
xnor U16009 (N_16009,N_15946,N_15805);
nor U16010 (N_16010,N_15800,N_15838);
nor U16011 (N_16011,N_15999,N_15906);
xor U16012 (N_16012,N_15789,N_15941);
or U16013 (N_16013,N_15823,N_15858);
or U16014 (N_16014,N_15774,N_15835);
xnor U16015 (N_16015,N_15836,N_15929);
or U16016 (N_16016,N_15850,N_15751);
nor U16017 (N_16017,N_15990,N_15813);
nor U16018 (N_16018,N_15908,N_15853);
or U16019 (N_16019,N_15770,N_15898);
and U16020 (N_16020,N_15977,N_15922);
nand U16021 (N_16021,N_15828,N_15916);
nor U16022 (N_16022,N_15937,N_15871);
xor U16023 (N_16023,N_15781,N_15829);
nor U16024 (N_16024,N_15764,N_15754);
xnor U16025 (N_16025,N_15880,N_15857);
nor U16026 (N_16026,N_15817,N_15914);
nand U16027 (N_16027,N_15833,N_15991);
or U16028 (N_16028,N_15890,N_15847);
or U16029 (N_16029,N_15983,N_15930);
nor U16030 (N_16030,N_15969,N_15927);
nor U16031 (N_16031,N_15773,N_15777);
or U16032 (N_16032,N_15998,N_15867);
xnor U16033 (N_16033,N_15887,N_15778);
or U16034 (N_16034,N_15976,N_15984);
and U16035 (N_16035,N_15962,N_15939);
nor U16036 (N_16036,N_15974,N_15830);
nor U16037 (N_16037,N_15905,N_15864);
nand U16038 (N_16038,N_15792,N_15957);
nand U16039 (N_16039,N_15963,N_15818);
or U16040 (N_16040,N_15869,N_15947);
nand U16041 (N_16041,N_15902,N_15921);
nor U16042 (N_16042,N_15938,N_15978);
nor U16043 (N_16043,N_15851,N_15782);
nor U16044 (N_16044,N_15812,N_15846);
and U16045 (N_16045,N_15893,N_15879);
nand U16046 (N_16046,N_15788,N_15882);
or U16047 (N_16047,N_15827,N_15750);
or U16048 (N_16048,N_15919,N_15840);
xor U16049 (N_16049,N_15960,N_15955);
nand U16050 (N_16050,N_15877,N_15903);
nor U16051 (N_16051,N_15854,N_15918);
or U16052 (N_16052,N_15756,N_15752);
xnor U16053 (N_16053,N_15943,N_15958);
xor U16054 (N_16054,N_15769,N_15761);
nand U16055 (N_16055,N_15992,N_15989);
nor U16056 (N_16056,N_15923,N_15994);
nor U16057 (N_16057,N_15860,N_15822);
or U16058 (N_16058,N_15886,N_15799);
nor U16059 (N_16059,N_15889,N_15925);
nand U16060 (N_16060,N_15873,N_15855);
nand U16061 (N_16061,N_15975,N_15896);
nand U16062 (N_16062,N_15856,N_15897);
and U16063 (N_16063,N_15894,N_15884);
and U16064 (N_16064,N_15791,N_15953);
xor U16065 (N_16065,N_15852,N_15785);
and U16066 (N_16066,N_15802,N_15913);
xnor U16067 (N_16067,N_15786,N_15971);
nand U16068 (N_16068,N_15876,N_15900);
and U16069 (N_16069,N_15763,N_15910);
xor U16070 (N_16070,N_15842,N_15936);
or U16071 (N_16071,N_15874,N_15888);
and U16072 (N_16072,N_15866,N_15796);
or U16073 (N_16073,N_15948,N_15932);
and U16074 (N_16074,N_15798,N_15891);
or U16075 (N_16075,N_15755,N_15935);
nor U16076 (N_16076,N_15972,N_15909);
xor U16077 (N_16077,N_15968,N_15807);
and U16078 (N_16078,N_15934,N_15895);
or U16079 (N_16079,N_15803,N_15753);
or U16080 (N_16080,N_15801,N_15945);
or U16081 (N_16081,N_15845,N_15861);
and U16082 (N_16082,N_15865,N_15816);
nand U16083 (N_16083,N_15804,N_15920);
and U16084 (N_16084,N_15848,N_15875);
xnor U16085 (N_16085,N_15787,N_15883);
nor U16086 (N_16086,N_15965,N_15988);
nor U16087 (N_16087,N_15815,N_15806);
nor U16088 (N_16088,N_15839,N_15964);
xor U16089 (N_16089,N_15926,N_15961);
or U16090 (N_16090,N_15772,N_15783);
or U16091 (N_16091,N_15970,N_15868);
nand U16092 (N_16092,N_15911,N_15954);
nor U16093 (N_16093,N_15834,N_15915);
nor U16094 (N_16094,N_15933,N_15849);
and U16095 (N_16095,N_15767,N_15809);
or U16096 (N_16096,N_15859,N_15776);
nand U16097 (N_16097,N_15794,N_15768);
and U16098 (N_16098,N_15950,N_15797);
and U16099 (N_16099,N_15949,N_15793);
nor U16100 (N_16100,N_15982,N_15997);
xnor U16101 (N_16101,N_15758,N_15995);
nor U16102 (N_16102,N_15901,N_15820);
and U16103 (N_16103,N_15904,N_15912);
xor U16104 (N_16104,N_15831,N_15759);
nand U16105 (N_16105,N_15795,N_15967);
nand U16106 (N_16106,N_15771,N_15832);
nand U16107 (N_16107,N_15765,N_15966);
nor U16108 (N_16108,N_15979,N_15790);
xnor U16109 (N_16109,N_15942,N_15821);
nor U16110 (N_16110,N_15996,N_15944);
nor U16111 (N_16111,N_15993,N_15931);
nor U16112 (N_16112,N_15863,N_15784);
nor U16113 (N_16113,N_15779,N_15862);
nor U16114 (N_16114,N_15907,N_15981);
nand U16115 (N_16115,N_15872,N_15951);
nor U16116 (N_16116,N_15980,N_15952);
nand U16117 (N_16117,N_15940,N_15844);
xnor U16118 (N_16118,N_15928,N_15837);
or U16119 (N_16119,N_15878,N_15841);
nand U16120 (N_16120,N_15987,N_15885);
nand U16121 (N_16121,N_15766,N_15780);
and U16122 (N_16122,N_15843,N_15762);
and U16123 (N_16123,N_15810,N_15826);
nand U16124 (N_16124,N_15811,N_15760);
nand U16125 (N_16125,N_15756,N_15813);
nor U16126 (N_16126,N_15891,N_15825);
xnor U16127 (N_16127,N_15923,N_15911);
nand U16128 (N_16128,N_15846,N_15867);
xnor U16129 (N_16129,N_15907,N_15753);
xor U16130 (N_16130,N_15770,N_15782);
nand U16131 (N_16131,N_15796,N_15931);
xor U16132 (N_16132,N_15796,N_15797);
or U16133 (N_16133,N_15916,N_15900);
nand U16134 (N_16134,N_15883,N_15798);
nand U16135 (N_16135,N_15857,N_15864);
nand U16136 (N_16136,N_15908,N_15760);
nand U16137 (N_16137,N_15780,N_15899);
nor U16138 (N_16138,N_15945,N_15852);
xor U16139 (N_16139,N_15985,N_15938);
xnor U16140 (N_16140,N_15978,N_15947);
xor U16141 (N_16141,N_15890,N_15916);
nor U16142 (N_16142,N_15788,N_15917);
and U16143 (N_16143,N_15994,N_15802);
nor U16144 (N_16144,N_15875,N_15774);
and U16145 (N_16145,N_15953,N_15908);
xor U16146 (N_16146,N_15901,N_15761);
or U16147 (N_16147,N_15933,N_15810);
and U16148 (N_16148,N_15885,N_15862);
xnor U16149 (N_16149,N_15880,N_15987);
nand U16150 (N_16150,N_15890,N_15880);
nor U16151 (N_16151,N_15979,N_15997);
nand U16152 (N_16152,N_15806,N_15862);
and U16153 (N_16153,N_15879,N_15979);
nand U16154 (N_16154,N_15785,N_15832);
nand U16155 (N_16155,N_15938,N_15851);
and U16156 (N_16156,N_15823,N_15962);
and U16157 (N_16157,N_15853,N_15820);
xor U16158 (N_16158,N_15773,N_15958);
nor U16159 (N_16159,N_15913,N_15755);
or U16160 (N_16160,N_15898,N_15897);
nand U16161 (N_16161,N_15897,N_15847);
xor U16162 (N_16162,N_15894,N_15792);
nor U16163 (N_16163,N_15971,N_15936);
or U16164 (N_16164,N_15857,N_15841);
or U16165 (N_16165,N_15985,N_15805);
or U16166 (N_16166,N_15898,N_15807);
or U16167 (N_16167,N_15913,N_15888);
or U16168 (N_16168,N_15821,N_15872);
nand U16169 (N_16169,N_15770,N_15868);
and U16170 (N_16170,N_15857,N_15997);
nor U16171 (N_16171,N_15785,N_15815);
nand U16172 (N_16172,N_15929,N_15954);
and U16173 (N_16173,N_15960,N_15818);
nand U16174 (N_16174,N_15835,N_15926);
xnor U16175 (N_16175,N_15808,N_15836);
nor U16176 (N_16176,N_15979,N_15794);
xnor U16177 (N_16177,N_15845,N_15801);
and U16178 (N_16178,N_15941,N_15975);
xor U16179 (N_16179,N_15850,N_15857);
or U16180 (N_16180,N_15977,N_15971);
and U16181 (N_16181,N_15811,N_15962);
nor U16182 (N_16182,N_15913,N_15838);
or U16183 (N_16183,N_15771,N_15958);
or U16184 (N_16184,N_15853,N_15781);
xor U16185 (N_16185,N_15966,N_15983);
and U16186 (N_16186,N_15820,N_15790);
and U16187 (N_16187,N_15907,N_15922);
and U16188 (N_16188,N_15993,N_15889);
and U16189 (N_16189,N_15899,N_15879);
nand U16190 (N_16190,N_15910,N_15987);
xnor U16191 (N_16191,N_15855,N_15982);
nor U16192 (N_16192,N_15864,N_15999);
nor U16193 (N_16193,N_15932,N_15910);
nor U16194 (N_16194,N_15830,N_15961);
and U16195 (N_16195,N_15918,N_15996);
nor U16196 (N_16196,N_15966,N_15888);
or U16197 (N_16197,N_15931,N_15891);
nand U16198 (N_16198,N_15973,N_15894);
nand U16199 (N_16199,N_15823,N_15987);
xnor U16200 (N_16200,N_15888,N_15997);
and U16201 (N_16201,N_15965,N_15945);
and U16202 (N_16202,N_15816,N_15876);
and U16203 (N_16203,N_15844,N_15843);
nand U16204 (N_16204,N_15910,N_15790);
nand U16205 (N_16205,N_15848,N_15853);
xnor U16206 (N_16206,N_15857,N_15835);
nor U16207 (N_16207,N_15905,N_15901);
nor U16208 (N_16208,N_15864,N_15975);
nand U16209 (N_16209,N_15813,N_15810);
and U16210 (N_16210,N_15951,N_15832);
xnor U16211 (N_16211,N_15964,N_15806);
and U16212 (N_16212,N_15904,N_15879);
and U16213 (N_16213,N_15830,N_15758);
nand U16214 (N_16214,N_15822,N_15959);
xor U16215 (N_16215,N_15893,N_15983);
and U16216 (N_16216,N_15908,N_15855);
nor U16217 (N_16217,N_15776,N_15807);
nand U16218 (N_16218,N_15872,N_15788);
nor U16219 (N_16219,N_15913,N_15901);
or U16220 (N_16220,N_15965,N_15833);
or U16221 (N_16221,N_15889,N_15867);
xnor U16222 (N_16222,N_15806,N_15849);
or U16223 (N_16223,N_15880,N_15922);
nor U16224 (N_16224,N_15779,N_15859);
xnor U16225 (N_16225,N_15893,N_15994);
nor U16226 (N_16226,N_15862,N_15959);
or U16227 (N_16227,N_15851,N_15947);
or U16228 (N_16228,N_15888,N_15860);
and U16229 (N_16229,N_15920,N_15985);
nand U16230 (N_16230,N_15808,N_15852);
nor U16231 (N_16231,N_15761,N_15984);
nor U16232 (N_16232,N_15900,N_15919);
and U16233 (N_16233,N_15899,N_15815);
and U16234 (N_16234,N_15910,N_15890);
nor U16235 (N_16235,N_15799,N_15806);
and U16236 (N_16236,N_15782,N_15890);
nand U16237 (N_16237,N_15751,N_15762);
xnor U16238 (N_16238,N_15918,N_15790);
nand U16239 (N_16239,N_15907,N_15987);
nand U16240 (N_16240,N_15777,N_15956);
xor U16241 (N_16241,N_15925,N_15938);
nand U16242 (N_16242,N_15903,N_15996);
and U16243 (N_16243,N_15859,N_15981);
nand U16244 (N_16244,N_15802,N_15974);
or U16245 (N_16245,N_15789,N_15953);
and U16246 (N_16246,N_15820,N_15904);
and U16247 (N_16247,N_15907,N_15812);
or U16248 (N_16248,N_15986,N_15860);
or U16249 (N_16249,N_15895,N_15755);
and U16250 (N_16250,N_16048,N_16143);
nand U16251 (N_16251,N_16237,N_16069);
nand U16252 (N_16252,N_16071,N_16134);
and U16253 (N_16253,N_16094,N_16200);
and U16254 (N_16254,N_16224,N_16093);
nand U16255 (N_16255,N_16183,N_16168);
and U16256 (N_16256,N_16004,N_16186);
nand U16257 (N_16257,N_16031,N_16214);
or U16258 (N_16258,N_16129,N_16121);
or U16259 (N_16259,N_16081,N_16023);
nand U16260 (N_16260,N_16162,N_16096);
xnor U16261 (N_16261,N_16032,N_16068);
xnor U16262 (N_16262,N_16054,N_16040);
or U16263 (N_16263,N_16243,N_16062);
nor U16264 (N_16264,N_16204,N_16212);
nor U16265 (N_16265,N_16242,N_16033);
xnor U16266 (N_16266,N_16110,N_16037);
nand U16267 (N_16267,N_16102,N_16114);
nand U16268 (N_16268,N_16160,N_16247);
and U16269 (N_16269,N_16026,N_16015);
nor U16270 (N_16270,N_16156,N_16169);
nand U16271 (N_16271,N_16058,N_16030);
xor U16272 (N_16272,N_16211,N_16007);
xnor U16273 (N_16273,N_16210,N_16187);
nand U16274 (N_16274,N_16227,N_16241);
nand U16275 (N_16275,N_16238,N_16053);
nand U16276 (N_16276,N_16085,N_16065);
or U16277 (N_16277,N_16146,N_16225);
nand U16278 (N_16278,N_16154,N_16017);
xor U16279 (N_16279,N_16099,N_16112);
xor U16280 (N_16280,N_16202,N_16052);
xor U16281 (N_16281,N_16235,N_16028);
or U16282 (N_16282,N_16232,N_16019);
and U16283 (N_16283,N_16008,N_16136);
xor U16284 (N_16284,N_16124,N_16185);
xor U16285 (N_16285,N_16066,N_16229);
xor U16286 (N_16286,N_16063,N_16117);
or U16287 (N_16287,N_16106,N_16181);
xor U16288 (N_16288,N_16043,N_16180);
and U16289 (N_16289,N_16190,N_16060);
xor U16290 (N_16290,N_16070,N_16199);
xor U16291 (N_16291,N_16098,N_16177);
and U16292 (N_16292,N_16233,N_16061);
and U16293 (N_16293,N_16105,N_16205);
and U16294 (N_16294,N_16158,N_16119);
xor U16295 (N_16295,N_16074,N_16024);
xnor U16296 (N_16296,N_16215,N_16127);
nor U16297 (N_16297,N_16239,N_16123);
nor U16298 (N_16298,N_16091,N_16223);
xor U16299 (N_16299,N_16115,N_16222);
nor U16300 (N_16300,N_16219,N_16050);
and U16301 (N_16301,N_16196,N_16072);
nor U16302 (N_16302,N_16100,N_16194);
xnor U16303 (N_16303,N_16109,N_16198);
nor U16304 (N_16304,N_16009,N_16145);
xor U16305 (N_16305,N_16001,N_16188);
nand U16306 (N_16306,N_16203,N_16178);
xor U16307 (N_16307,N_16064,N_16038);
or U16308 (N_16308,N_16151,N_16021);
nor U16309 (N_16309,N_16095,N_16059);
nand U16310 (N_16310,N_16116,N_16163);
nand U16311 (N_16311,N_16044,N_16216);
and U16312 (N_16312,N_16138,N_16122);
nand U16313 (N_16313,N_16039,N_16167);
and U16314 (N_16314,N_16249,N_16003);
nor U16315 (N_16315,N_16041,N_16155);
nand U16316 (N_16316,N_16171,N_16209);
xnor U16317 (N_16317,N_16049,N_16088);
or U16318 (N_16318,N_16213,N_16150);
nor U16319 (N_16319,N_16131,N_16228);
nor U16320 (N_16320,N_16148,N_16020);
or U16321 (N_16321,N_16079,N_16240);
or U16322 (N_16322,N_16226,N_16164);
or U16323 (N_16323,N_16104,N_16244);
nor U16324 (N_16324,N_16010,N_16236);
nand U16325 (N_16325,N_16182,N_16218);
or U16326 (N_16326,N_16108,N_16246);
and U16327 (N_16327,N_16016,N_16087);
xor U16328 (N_16328,N_16018,N_16221);
and U16329 (N_16329,N_16170,N_16002);
nor U16330 (N_16330,N_16137,N_16207);
xnor U16331 (N_16331,N_16152,N_16035);
nand U16332 (N_16332,N_16083,N_16084);
nor U16333 (N_16333,N_16147,N_16132);
nor U16334 (N_16334,N_16176,N_16184);
nand U16335 (N_16335,N_16092,N_16220);
nand U16336 (N_16336,N_16125,N_16245);
nor U16337 (N_16337,N_16042,N_16047);
nor U16338 (N_16338,N_16159,N_16142);
or U16339 (N_16339,N_16097,N_16101);
nand U16340 (N_16340,N_16130,N_16103);
or U16341 (N_16341,N_16165,N_16034);
nand U16342 (N_16342,N_16022,N_16166);
xnor U16343 (N_16343,N_16208,N_16161);
and U16344 (N_16344,N_16036,N_16128);
xnor U16345 (N_16345,N_16135,N_16014);
and U16346 (N_16346,N_16141,N_16089);
and U16347 (N_16347,N_16140,N_16057);
and U16348 (N_16348,N_16126,N_16012);
and U16349 (N_16349,N_16013,N_16230);
xnor U16350 (N_16350,N_16080,N_16113);
or U16351 (N_16351,N_16056,N_16111);
and U16352 (N_16352,N_16067,N_16120);
and U16353 (N_16353,N_16076,N_16000);
xnor U16354 (N_16354,N_16073,N_16051);
xnor U16355 (N_16355,N_16206,N_16173);
nand U16356 (N_16356,N_16149,N_16157);
nor U16357 (N_16357,N_16179,N_16086);
or U16358 (N_16358,N_16234,N_16248);
nor U16359 (N_16359,N_16077,N_16107);
and U16360 (N_16360,N_16046,N_16201);
and U16361 (N_16361,N_16144,N_16192);
nand U16362 (N_16362,N_16011,N_16191);
xor U16363 (N_16363,N_16197,N_16189);
or U16364 (N_16364,N_16025,N_16172);
nor U16365 (N_16365,N_16005,N_16175);
nand U16366 (N_16366,N_16055,N_16118);
nor U16367 (N_16367,N_16075,N_16139);
nor U16368 (N_16368,N_16153,N_16082);
or U16369 (N_16369,N_16231,N_16045);
nand U16370 (N_16370,N_16078,N_16174);
nand U16371 (N_16371,N_16193,N_16027);
nand U16372 (N_16372,N_16006,N_16090);
xor U16373 (N_16373,N_16133,N_16195);
nand U16374 (N_16374,N_16217,N_16029);
or U16375 (N_16375,N_16012,N_16232);
and U16376 (N_16376,N_16165,N_16033);
or U16377 (N_16377,N_16076,N_16085);
nand U16378 (N_16378,N_16115,N_16045);
nor U16379 (N_16379,N_16044,N_16046);
nor U16380 (N_16380,N_16063,N_16112);
and U16381 (N_16381,N_16239,N_16137);
nor U16382 (N_16382,N_16045,N_16062);
nand U16383 (N_16383,N_16098,N_16069);
and U16384 (N_16384,N_16239,N_16032);
xor U16385 (N_16385,N_16244,N_16161);
xor U16386 (N_16386,N_16179,N_16089);
nand U16387 (N_16387,N_16129,N_16125);
and U16388 (N_16388,N_16029,N_16202);
and U16389 (N_16389,N_16074,N_16153);
and U16390 (N_16390,N_16176,N_16141);
or U16391 (N_16391,N_16215,N_16102);
nand U16392 (N_16392,N_16053,N_16233);
nor U16393 (N_16393,N_16216,N_16110);
and U16394 (N_16394,N_16069,N_16060);
and U16395 (N_16395,N_16186,N_16048);
xor U16396 (N_16396,N_16191,N_16119);
xor U16397 (N_16397,N_16102,N_16157);
xor U16398 (N_16398,N_16114,N_16108);
and U16399 (N_16399,N_16070,N_16194);
nand U16400 (N_16400,N_16097,N_16013);
nand U16401 (N_16401,N_16235,N_16012);
or U16402 (N_16402,N_16117,N_16235);
nand U16403 (N_16403,N_16147,N_16089);
and U16404 (N_16404,N_16105,N_16064);
and U16405 (N_16405,N_16132,N_16115);
or U16406 (N_16406,N_16130,N_16234);
nor U16407 (N_16407,N_16244,N_16181);
nand U16408 (N_16408,N_16232,N_16226);
xnor U16409 (N_16409,N_16011,N_16091);
nor U16410 (N_16410,N_16165,N_16233);
or U16411 (N_16411,N_16248,N_16217);
or U16412 (N_16412,N_16114,N_16121);
and U16413 (N_16413,N_16041,N_16104);
or U16414 (N_16414,N_16167,N_16208);
xor U16415 (N_16415,N_16064,N_16146);
or U16416 (N_16416,N_16152,N_16098);
xnor U16417 (N_16417,N_16177,N_16116);
nor U16418 (N_16418,N_16085,N_16129);
and U16419 (N_16419,N_16188,N_16120);
xor U16420 (N_16420,N_16248,N_16118);
nand U16421 (N_16421,N_16046,N_16050);
nand U16422 (N_16422,N_16230,N_16223);
or U16423 (N_16423,N_16216,N_16063);
xnor U16424 (N_16424,N_16087,N_16190);
and U16425 (N_16425,N_16060,N_16103);
and U16426 (N_16426,N_16013,N_16034);
and U16427 (N_16427,N_16116,N_16049);
or U16428 (N_16428,N_16075,N_16083);
nor U16429 (N_16429,N_16019,N_16048);
nor U16430 (N_16430,N_16239,N_16183);
and U16431 (N_16431,N_16038,N_16167);
nor U16432 (N_16432,N_16234,N_16127);
nor U16433 (N_16433,N_16238,N_16017);
nand U16434 (N_16434,N_16204,N_16151);
or U16435 (N_16435,N_16174,N_16123);
or U16436 (N_16436,N_16204,N_16185);
and U16437 (N_16437,N_16162,N_16140);
and U16438 (N_16438,N_16006,N_16092);
xnor U16439 (N_16439,N_16101,N_16109);
or U16440 (N_16440,N_16070,N_16118);
nand U16441 (N_16441,N_16047,N_16101);
nor U16442 (N_16442,N_16012,N_16080);
or U16443 (N_16443,N_16105,N_16087);
nand U16444 (N_16444,N_16193,N_16239);
nor U16445 (N_16445,N_16154,N_16242);
xnor U16446 (N_16446,N_16169,N_16048);
and U16447 (N_16447,N_16178,N_16042);
nor U16448 (N_16448,N_16178,N_16241);
or U16449 (N_16449,N_16182,N_16064);
xor U16450 (N_16450,N_16173,N_16050);
nand U16451 (N_16451,N_16189,N_16242);
nand U16452 (N_16452,N_16107,N_16177);
nand U16453 (N_16453,N_16233,N_16032);
or U16454 (N_16454,N_16110,N_16068);
or U16455 (N_16455,N_16099,N_16014);
nand U16456 (N_16456,N_16241,N_16181);
and U16457 (N_16457,N_16026,N_16064);
nor U16458 (N_16458,N_16243,N_16190);
nor U16459 (N_16459,N_16122,N_16106);
nor U16460 (N_16460,N_16063,N_16092);
and U16461 (N_16461,N_16222,N_16192);
nor U16462 (N_16462,N_16007,N_16060);
nor U16463 (N_16463,N_16220,N_16213);
nand U16464 (N_16464,N_16238,N_16123);
nand U16465 (N_16465,N_16206,N_16183);
nand U16466 (N_16466,N_16150,N_16133);
xor U16467 (N_16467,N_16204,N_16112);
and U16468 (N_16468,N_16205,N_16104);
or U16469 (N_16469,N_16005,N_16001);
xor U16470 (N_16470,N_16135,N_16174);
and U16471 (N_16471,N_16074,N_16238);
or U16472 (N_16472,N_16172,N_16177);
xnor U16473 (N_16473,N_16119,N_16181);
and U16474 (N_16474,N_16009,N_16229);
or U16475 (N_16475,N_16016,N_16223);
xor U16476 (N_16476,N_16067,N_16058);
xor U16477 (N_16477,N_16100,N_16178);
xor U16478 (N_16478,N_16073,N_16149);
nor U16479 (N_16479,N_16010,N_16142);
xor U16480 (N_16480,N_16143,N_16096);
xor U16481 (N_16481,N_16140,N_16127);
or U16482 (N_16482,N_16041,N_16093);
and U16483 (N_16483,N_16051,N_16121);
nor U16484 (N_16484,N_16107,N_16032);
nand U16485 (N_16485,N_16033,N_16106);
and U16486 (N_16486,N_16139,N_16232);
or U16487 (N_16487,N_16045,N_16158);
xor U16488 (N_16488,N_16149,N_16101);
nand U16489 (N_16489,N_16005,N_16141);
or U16490 (N_16490,N_16155,N_16195);
nor U16491 (N_16491,N_16149,N_16199);
and U16492 (N_16492,N_16212,N_16090);
and U16493 (N_16493,N_16098,N_16247);
or U16494 (N_16494,N_16094,N_16003);
nor U16495 (N_16495,N_16242,N_16210);
xor U16496 (N_16496,N_16134,N_16205);
xor U16497 (N_16497,N_16082,N_16005);
or U16498 (N_16498,N_16203,N_16133);
xnor U16499 (N_16499,N_16188,N_16162);
or U16500 (N_16500,N_16331,N_16478);
or U16501 (N_16501,N_16253,N_16443);
nor U16502 (N_16502,N_16411,N_16303);
nor U16503 (N_16503,N_16435,N_16454);
and U16504 (N_16504,N_16315,N_16422);
xor U16505 (N_16505,N_16321,N_16417);
xor U16506 (N_16506,N_16346,N_16397);
and U16507 (N_16507,N_16440,N_16309);
or U16508 (N_16508,N_16258,N_16424);
xor U16509 (N_16509,N_16349,N_16415);
nor U16510 (N_16510,N_16353,N_16425);
or U16511 (N_16511,N_16280,N_16264);
nand U16512 (N_16512,N_16407,N_16496);
or U16513 (N_16513,N_16481,N_16398);
nor U16514 (N_16514,N_16328,N_16467);
xor U16515 (N_16515,N_16486,N_16271);
nor U16516 (N_16516,N_16493,N_16463);
nand U16517 (N_16517,N_16396,N_16325);
nor U16518 (N_16518,N_16433,N_16345);
and U16519 (N_16519,N_16497,N_16354);
and U16520 (N_16520,N_16394,N_16455);
or U16521 (N_16521,N_16342,N_16307);
nor U16522 (N_16522,N_16388,N_16360);
and U16523 (N_16523,N_16469,N_16372);
or U16524 (N_16524,N_16368,N_16423);
xnor U16525 (N_16525,N_16439,N_16350);
nor U16526 (N_16526,N_16337,N_16343);
nand U16527 (N_16527,N_16274,N_16319);
or U16528 (N_16528,N_16340,N_16299);
xor U16529 (N_16529,N_16428,N_16414);
and U16530 (N_16530,N_16359,N_16302);
or U16531 (N_16531,N_16498,N_16404);
nor U16532 (N_16532,N_16330,N_16326);
nor U16533 (N_16533,N_16399,N_16300);
xnor U16534 (N_16534,N_16301,N_16316);
nor U16535 (N_16535,N_16431,N_16445);
nand U16536 (N_16536,N_16357,N_16289);
or U16537 (N_16537,N_16489,N_16392);
nand U16538 (N_16538,N_16312,N_16421);
xnor U16539 (N_16539,N_16306,N_16441);
xnor U16540 (N_16540,N_16263,N_16487);
nand U16541 (N_16541,N_16281,N_16381);
and U16542 (N_16542,N_16288,N_16276);
or U16543 (N_16543,N_16362,N_16485);
xnor U16544 (N_16544,N_16255,N_16311);
xnor U16545 (N_16545,N_16484,N_16494);
xor U16546 (N_16546,N_16495,N_16291);
or U16547 (N_16547,N_16282,N_16283);
xnor U16548 (N_16548,N_16260,N_16450);
nand U16549 (N_16549,N_16279,N_16488);
nor U16550 (N_16550,N_16436,N_16416);
xor U16551 (N_16551,N_16338,N_16273);
xor U16552 (N_16552,N_16266,N_16389);
xnor U16553 (N_16553,N_16395,N_16472);
or U16554 (N_16554,N_16341,N_16332);
xnor U16555 (N_16555,N_16434,N_16476);
and U16556 (N_16556,N_16310,N_16387);
nor U16557 (N_16557,N_16275,N_16452);
nor U16558 (N_16558,N_16400,N_16317);
xor U16559 (N_16559,N_16297,N_16305);
nor U16560 (N_16560,N_16351,N_16418);
nor U16561 (N_16561,N_16430,N_16327);
and U16562 (N_16562,N_16278,N_16358);
and U16563 (N_16563,N_16401,N_16367);
and U16564 (N_16564,N_16470,N_16426);
or U16565 (N_16565,N_16479,N_16363);
and U16566 (N_16566,N_16313,N_16277);
and U16567 (N_16567,N_16406,N_16413);
xor U16568 (N_16568,N_16403,N_16322);
and U16569 (N_16569,N_16270,N_16268);
xor U16570 (N_16570,N_16444,N_16473);
and U16571 (N_16571,N_16456,N_16348);
xnor U16572 (N_16572,N_16465,N_16405);
or U16573 (N_16573,N_16390,N_16383);
and U16574 (N_16574,N_16457,N_16352);
and U16575 (N_16575,N_16458,N_16380);
nand U16576 (N_16576,N_16480,N_16371);
nand U16577 (N_16577,N_16471,N_16334);
xnor U16578 (N_16578,N_16369,N_16293);
and U16579 (N_16579,N_16462,N_16420);
nor U16580 (N_16580,N_16377,N_16296);
and U16581 (N_16581,N_16318,N_16460);
or U16582 (N_16582,N_16286,N_16290);
xnor U16583 (N_16583,N_16370,N_16329);
nand U16584 (N_16584,N_16308,N_16393);
or U16585 (N_16585,N_16298,N_16408);
nor U16586 (N_16586,N_16347,N_16442);
xnor U16587 (N_16587,N_16295,N_16385);
or U16588 (N_16588,N_16491,N_16335);
xnor U16589 (N_16589,N_16259,N_16429);
or U16590 (N_16590,N_16257,N_16451);
xor U16591 (N_16591,N_16323,N_16459);
xnor U16592 (N_16592,N_16386,N_16292);
or U16593 (N_16593,N_16468,N_16475);
or U16594 (N_16594,N_16254,N_16256);
and U16595 (N_16595,N_16265,N_16336);
xor U16596 (N_16596,N_16261,N_16250);
and U16597 (N_16597,N_16269,N_16447);
xor U16598 (N_16598,N_16361,N_16262);
xor U16599 (N_16599,N_16294,N_16382);
nand U16600 (N_16600,N_16437,N_16449);
nand U16601 (N_16601,N_16374,N_16375);
and U16602 (N_16602,N_16438,N_16376);
nor U16603 (N_16603,N_16344,N_16373);
and U16604 (N_16604,N_16419,N_16410);
or U16605 (N_16605,N_16466,N_16402);
and U16606 (N_16606,N_16324,N_16365);
nand U16607 (N_16607,N_16482,N_16314);
nand U16608 (N_16608,N_16499,N_16490);
xnor U16609 (N_16609,N_16391,N_16356);
xor U16610 (N_16610,N_16339,N_16464);
nand U16611 (N_16611,N_16304,N_16272);
or U16612 (N_16612,N_16483,N_16409);
and U16613 (N_16613,N_16378,N_16333);
and U16614 (N_16614,N_16427,N_16384);
or U16615 (N_16615,N_16492,N_16412);
xor U16616 (N_16616,N_16320,N_16379);
nand U16617 (N_16617,N_16446,N_16364);
nand U16618 (N_16618,N_16287,N_16267);
and U16619 (N_16619,N_16355,N_16453);
or U16620 (N_16620,N_16474,N_16285);
and U16621 (N_16621,N_16366,N_16251);
and U16622 (N_16622,N_16284,N_16252);
xor U16623 (N_16623,N_16448,N_16461);
nand U16624 (N_16624,N_16432,N_16477);
nor U16625 (N_16625,N_16311,N_16430);
and U16626 (N_16626,N_16381,N_16411);
and U16627 (N_16627,N_16369,N_16288);
nand U16628 (N_16628,N_16334,N_16301);
and U16629 (N_16629,N_16492,N_16397);
xor U16630 (N_16630,N_16435,N_16486);
or U16631 (N_16631,N_16345,N_16346);
nand U16632 (N_16632,N_16401,N_16263);
xnor U16633 (N_16633,N_16454,N_16310);
nand U16634 (N_16634,N_16274,N_16297);
nor U16635 (N_16635,N_16485,N_16391);
nor U16636 (N_16636,N_16306,N_16289);
nor U16637 (N_16637,N_16393,N_16406);
nand U16638 (N_16638,N_16366,N_16387);
xnor U16639 (N_16639,N_16427,N_16486);
nor U16640 (N_16640,N_16498,N_16418);
xor U16641 (N_16641,N_16428,N_16486);
xor U16642 (N_16642,N_16303,N_16483);
and U16643 (N_16643,N_16445,N_16291);
or U16644 (N_16644,N_16497,N_16468);
nor U16645 (N_16645,N_16362,N_16284);
nor U16646 (N_16646,N_16338,N_16488);
nor U16647 (N_16647,N_16471,N_16492);
xnor U16648 (N_16648,N_16323,N_16394);
nor U16649 (N_16649,N_16397,N_16410);
nand U16650 (N_16650,N_16338,N_16414);
xor U16651 (N_16651,N_16333,N_16367);
nand U16652 (N_16652,N_16481,N_16352);
or U16653 (N_16653,N_16335,N_16273);
nand U16654 (N_16654,N_16402,N_16285);
xnor U16655 (N_16655,N_16453,N_16312);
xnor U16656 (N_16656,N_16365,N_16478);
nor U16657 (N_16657,N_16408,N_16268);
nor U16658 (N_16658,N_16300,N_16416);
and U16659 (N_16659,N_16253,N_16402);
xor U16660 (N_16660,N_16339,N_16467);
nand U16661 (N_16661,N_16278,N_16258);
nor U16662 (N_16662,N_16442,N_16370);
xnor U16663 (N_16663,N_16323,N_16382);
nor U16664 (N_16664,N_16305,N_16482);
nand U16665 (N_16665,N_16485,N_16323);
xnor U16666 (N_16666,N_16307,N_16250);
xnor U16667 (N_16667,N_16394,N_16340);
xnor U16668 (N_16668,N_16344,N_16266);
nand U16669 (N_16669,N_16433,N_16471);
or U16670 (N_16670,N_16494,N_16451);
xnor U16671 (N_16671,N_16327,N_16417);
nand U16672 (N_16672,N_16292,N_16429);
nor U16673 (N_16673,N_16298,N_16336);
xor U16674 (N_16674,N_16494,N_16338);
nand U16675 (N_16675,N_16484,N_16451);
and U16676 (N_16676,N_16350,N_16307);
nor U16677 (N_16677,N_16429,N_16267);
nor U16678 (N_16678,N_16470,N_16360);
nand U16679 (N_16679,N_16462,N_16294);
and U16680 (N_16680,N_16408,N_16269);
nor U16681 (N_16681,N_16298,N_16379);
nand U16682 (N_16682,N_16443,N_16460);
and U16683 (N_16683,N_16429,N_16387);
nand U16684 (N_16684,N_16298,N_16398);
or U16685 (N_16685,N_16394,N_16414);
and U16686 (N_16686,N_16321,N_16437);
nor U16687 (N_16687,N_16309,N_16315);
and U16688 (N_16688,N_16456,N_16493);
nand U16689 (N_16689,N_16402,N_16350);
or U16690 (N_16690,N_16293,N_16357);
nand U16691 (N_16691,N_16428,N_16274);
and U16692 (N_16692,N_16459,N_16310);
and U16693 (N_16693,N_16362,N_16467);
xnor U16694 (N_16694,N_16421,N_16386);
or U16695 (N_16695,N_16440,N_16403);
nand U16696 (N_16696,N_16252,N_16459);
or U16697 (N_16697,N_16389,N_16302);
nor U16698 (N_16698,N_16255,N_16259);
or U16699 (N_16699,N_16378,N_16300);
and U16700 (N_16700,N_16452,N_16368);
or U16701 (N_16701,N_16286,N_16278);
or U16702 (N_16702,N_16452,N_16330);
or U16703 (N_16703,N_16492,N_16452);
or U16704 (N_16704,N_16360,N_16480);
and U16705 (N_16705,N_16478,N_16498);
xnor U16706 (N_16706,N_16405,N_16270);
nor U16707 (N_16707,N_16458,N_16274);
nand U16708 (N_16708,N_16315,N_16316);
xnor U16709 (N_16709,N_16276,N_16338);
xor U16710 (N_16710,N_16250,N_16339);
or U16711 (N_16711,N_16314,N_16375);
or U16712 (N_16712,N_16397,N_16343);
and U16713 (N_16713,N_16370,N_16331);
xor U16714 (N_16714,N_16453,N_16309);
and U16715 (N_16715,N_16479,N_16417);
nor U16716 (N_16716,N_16437,N_16264);
or U16717 (N_16717,N_16433,N_16486);
and U16718 (N_16718,N_16349,N_16342);
xnor U16719 (N_16719,N_16340,N_16364);
and U16720 (N_16720,N_16345,N_16307);
nor U16721 (N_16721,N_16458,N_16448);
or U16722 (N_16722,N_16252,N_16363);
or U16723 (N_16723,N_16478,N_16429);
nand U16724 (N_16724,N_16408,N_16295);
and U16725 (N_16725,N_16384,N_16459);
nor U16726 (N_16726,N_16322,N_16440);
nand U16727 (N_16727,N_16290,N_16430);
xnor U16728 (N_16728,N_16350,N_16333);
and U16729 (N_16729,N_16457,N_16395);
and U16730 (N_16730,N_16431,N_16318);
nand U16731 (N_16731,N_16324,N_16402);
or U16732 (N_16732,N_16480,N_16253);
and U16733 (N_16733,N_16264,N_16394);
nor U16734 (N_16734,N_16467,N_16436);
nand U16735 (N_16735,N_16444,N_16372);
nor U16736 (N_16736,N_16271,N_16345);
nor U16737 (N_16737,N_16448,N_16402);
nand U16738 (N_16738,N_16430,N_16307);
nand U16739 (N_16739,N_16497,N_16389);
xor U16740 (N_16740,N_16278,N_16339);
nor U16741 (N_16741,N_16334,N_16403);
nand U16742 (N_16742,N_16458,N_16445);
nand U16743 (N_16743,N_16338,N_16268);
nand U16744 (N_16744,N_16274,N_16363);
or U16745 (N_16745,N_16424,N_16430);
or U16746 (N_16746,N_16299,N_16488);
and U16747 (N_16747,N_16389,N_16414);
nand U16748 (N_16748,N_16292,N_16388);
xnor U16749 (N_16749,N_16274,N_16403);
and U16750 (N_16750,N_16544,N_16559);
or U16751 (N_16751,N_16678,N_16741);
xnor U16752 (N_16752,N_16686,N_16703);
or U16753 (N_16753,N_16645,N_16680);
or U16754 (N_16754,N_16724,N_16653);
nor U16755 (N_16755,N_16742,N_16743);
or U16756 (N_16756,N_16633,N_16608);
and U16757 (N_16757,N_16704,N_16650);
xor U16758 (N_16758,N_16710,N_16551);
and U16759 (N_16759,N_16589,N_16723);
nor U16760 (N_16760,N_16695,N_16727);
nand U16761 (N_16761,N_16513,N_16746);
and U16762 (N_16762,N_16581,N_16531);
and U16763 (N_16763,N_16639,N_16749);
nor U16764 (N_16764,N_16575,N_16655);
nor U16765 (N_16765,N_16651,N_16643);
nor U16766 (N_16766,N_16506,N_16698);
nor U16767 (N_16767,N_16640,N_16622);
nand U16768 (N_16768,N_16574,N_16524);
and U16769 (N_16769,N_16607,N_16595);
or U16770 (N_16770,N_16587,N_16736);
or U16771 (N_16771,N_16725,N_16648);
and U16772 (N_16772,N_16718,N_16500);
nand U16773 (N_16773,N_16674,N_16738);
xor U16774 (N_16774,N_16707,N_16702);
and U16775 (N_16775,N_16654,N_16629);
nand U16776 (N_16776,N_16526,N_16584);
nand U16777 (N_16777,N_16576,N_16693);
or U16778 (N_16778,N_16681,N_16549);
and U16779 (N_16779,N_16537,N_16519);
nand U16780 (N_16780,N_16522,N_16553);
xnor U16781 (N_16781,N_16730,N_16615);
nand U16782 (N_16782,N_16568,N_16744);
xnor U16783 (N_16783,N_16631,N_16700);
and U16784 (N_16784,N_16656,N_16572);
xor U16785 (N_16785,N_16600,N_16635);
and U16786 (N_16786,N_16632,N_16729);
or U16787 (N_16787,N_16660,N_16721);
xor U16788 (N_16788,N_16665,N_16542);
nand U16789 (N_16789,N_16592,N_16708);
nor U16790 (N_16790,N_16610,N_16566);
nand U16791 (N_16791,N_16521,N_16647);
or U16792 (N_16792,N_16518,N_16726);
or U16793 (N_16793,N_16605,N_16530);
or U16794 (N_16794,N_16617,N_16536);
xor U16795 (N_16795,N_16578,N_16685);
xnor U16796 (N_16796,N_16585,N_16565);
nor U16797 (N_16797,N_16720,N_16512);
nand U16798 (N_16798,N_16666,N_16560);
nand U16799 (N_16799,N_16667,N_16705);
xor U16800 (N_16800,N_16533,N_16508);
nor U16801 (N_16801,N_16555,N_16603);
and U16802 (N_16802,N_16613,N_16604);
or U16803 (N_16803,N_16675,N_16694);
nor U16804 (N_16804,N_16547,N_16642);
and U16805 (N_16805,N_16644,N_16599);
nor U16806 (N_16806,N_16534,N_16507);
nand U16807 (N_16807,N_16683,N_16696);
and U16808 (N_16808,N_16731,N_16535);
and U16809 (N_16809,N_16502,N_16571);
or U16810 (N_16810,N_16503,N_16596);
or U16811 (N_16811,N_16561,N_16541);
nor U16812 (N_16812,N_16658,N_16664);
or U16813 (N_16813,N_16557,N_16662);
and U16814 (N_16814,N_16601,N_16594);
xnor U16815 (N_16815,N_16583,N_16719);
xnor U16816 (N_16816,N_16509,N_16624);
nor U16817 (N_16817,N_16690,N_16563);
nor U16818 (N_16818,N_16668,N_16618);
xor U16819 (N_16819,N_16567,N_16735);
nor U16820 (N_16820,N_16593,N_16646);
nand U16821 (N_16821,N_16525,N_16616);
or U16822 (N_16822,N_16682,N_16649);
or U16823 (N_16823,N_16579,N_16562);
xor U16824 (N_16824,N_16699,N_16548);
nand U16825 (N_16825,N_16505,N_16523);
or U16826 (N_16826,N_16527,N_16625);
xnor U16827 (N_16827,N_16554,N_16545);
or U16828 (N_16828,N_16539,N_16728);
nand U16829 (N_16829,N_16709,N_16638);
nor U16830 (N_16830,N_16711,N_16620);
or U16831 (N_16831,N_16634,N_16689);
or U16832 (N_16832,N_16716,N_16715);
xnor U16833 (N_16833,N_16673,N_16598);
and U16834 (N_16834,N_16588,N_16687);
or U16835 (N_16835,N_16676,N_16684);
xnor U16836 (N_16836,N_16520,N_16661);
and U16837 (N_16837,N_16672,N_16546);
and U16838 (N_16838,N_16517,N_16669);
and U16839 (N_16839,N_16573,N_16627);
and U16840 (N_16840,N_16611,N_16543);
or U16841 (N_16841,N_16529,N_16657);
and U16842 (N_16842,N_16663,N_16670);
nand U16843 (N_16843,N_16582,N_16652);
nor U16844 (N_16844,N_16628,N_16734);
nor U16845 (N_16845,N_16590,N_16732);
and U16846 (N_16846,N_16597,N_16591);
xor U16847 (N_16847,N_16747,N_16733);
and U16848 (N_16848,N_16609,N_16740);
xnor U16849 (N_16849,N_16659,N_16714);
or U16850 (N_16850,N_16556,N_16745);
or U16851 (N_16851,N_16748,N_16552);
nand U16852 (N_16852,N_16739,N_16737);
xnor U16853 (N_16853,N_16612,N_16641);
or U16854 (N_16854,N_16671,N_16586);
nand U16855 (N_16855,N_16717,N_16692);
or U16856 (N_16856,N_16606,N_16619);
xor U16857 (N_16857,N_16688,N_16630);
or U16858 (N_16858,N_16722,N_16511);
and U16859 (N_16859,N_16679,N_16550);
xor U16860 (N_16860,N_16713,N_16538);
nor U16861 (N_16861,N_16602,N_16691);
or U16862 (N_16862,N_16637,N_16712);
or U16863 (N_16863,N_16614,N_16570);
or U16864 (N_16864,N_16558,N_16532);
and U16865 (N_16865,N_16504,N_16516);
and U16866 (N_16866,N_16636,N_16514);
xnor U16867 (N_16867,N_16540,N_16623);
nor U16868 (N_16868,N_16621,N_16515);
nor U16869 (N_16869,N_16701,N_16580);
nor U16870 (N_16870,N_16577,N_16510);
or U16871 (N_16871,N_16564,N_16569);
and U16872 (N_16872,N_16706,N_16677);
nand U16873 (N_16873,N_16697,N_16501);
xor U16874 (N_16874,N_16626,N_16528);
xnor U16875 (N_16875,N_16538,N_16565);
or U16876 (N_16876,N_16608,N_16626);
xnor U16877 (N_16877,N_16713,N_16720);
xor U16878 (N_16878,N_16544,N_16669);
and U16879 (N_16879,N_16744,N_16664);
and U16880 (N_16880,N_16544,N_16553);
and U16881 (N_16881,N_16654,N_16650);
nor U16882 (N_16882,N_16596,N_16566);
nor U16883 (N_16883,N_16522,N_16686);
and U16884 (N_16884,N_16650,N_16651);
and U16885 (N_16885,N_16724,N_16674);
nand U16886 (N_16886,N_16699,N_16614);
and U16887 (N_16887,N_16702,N_16619);
xnor U16888 (N_16888,N_16740,N_16565);
nand U16889 (N_16889,N_16590,N_16583);
nor U16890 (N_16890,N_16638,N_16526);
nand U16891 (N_16891,N_16556,N_16682);
nand U16892 (N_16892,N_16506,N_16720);
xnor U16893 (N_16893,N_16646,N_16558);
xnor U16894 (N_16894,N_16749,N_16657);
nand U16895 (N_16895,N_16706,N_16712);
nand U16896 (N_16896,N_16627,N_16647);
xnor U16897 (N_16897,N_16673,N_16555);
xnor U16898 (N_16898,N_16746,N_16684);
xnor U16899 (N_16899,N_16721,N_16632);
nor U16900 (N_16900,N_16559,N_16609);
nor U16901 (N_16901,N_16719,N_16701);
nor U16902 (N_16902,N_16633,N_16599);
nand U16903 (N_16903,N_16715,N_16532);
nand U16904 (N_16904,N_16636,N_16583);
nand U16905 (N_16905,N_16570,N_16586);
nand U16906 (N_16906,N_16529,N_16534);
and U16907 (N_16907,N_16658,N_16734);
or U16908 (N_16908,N_16569,N_16561);
and U16909 (N_16909,N_16567,N_16616);
nor U16910 (N_16910,N_16605,N_16744);
xnor U16911 (N_16911,N_16732,N_16665);
nand U16912 (N_16912,N_16611,N_16528);
nand U16913 (N_16913,N_16698,N_16737);
and U16914 (N_16914,N_16675,N_16648);
nand U16915 (N_16915,N_16523,N_16719);
xor U16916 (N_16916,N_16525,N_16647);
nor U16917 (N_16917,N_16744,N_16604);
and U16918 (N_16918,N_16728,N_16512);
xor U16919 (N_16919,N_16673,N_16735);
or U16920 (N_16920,N_16662,N_16695);
xnor U16921 (N_16921,N_16527,N_16684);
and U16922 (N_16922,N_16615,N_16529);
xnor U16923 (N_16923,N_16709,N_16692);
xnor U16924 (N_16924,N_16620,N_16624);
and U16925 (N_16925,N_16557,N_16550);
xnor U16926 (N_16926,N_16585,N_16534);
nor U16927 (N_16927,N_16705,N_16593);
nand U16928 (N_16928,N_16668,N_16729);
nor U16929 (N_16929,N_16712,N_16521);
nor U16930 (N_16930,N_16542,N_16596);
nor U16931 (N_16931,N_16545,N_16596);
or U16932 (N_16932,N_16706,N_16747);
nor U16933 (N_16933,N_16730,N_16561);
and U16934 (N_16934,N_16547,N_16649);
nor U16935 (N_16935,N_16507,N_16625);
xor U16936 (N_16936,N_16546,N_16556);
xor U16937 (N_16937,N_16526,N_16580);
and U16938 (N_16938,N_16581,N_16555);
nor U16939 (N_16939,N_16546,N_16736);
xor U16940 (N_16940,N_16652,N_16703);
nor U16941 (N_16941,N_16673,N_16611);
xor U16942 (N_16942,N_16630,N_16526);
or U16943 (N_16943,N_16555,N_16737);
and U16944 (N_16944,N_16679,N_16511);
or U16945 (N_16945,N_16581,N_16696);
and U16946 (N_16946,N_16601,N_16703);
xor U16947 (N_16947,N_16588,N_16640);
nor U16948 (N_16948,N_16513,N_16716);
xor U16949 (N_16949,N_16730,N_16518);
nor U16950 (N_16950,N_16639,N_16571);
or U16951 (N_16951,N_16705,N_16600);
xnor U16952 (N_16952,N_16596,N_16603);
xnor U16953 (N_16953,N_16587,N_16656);
and U16954 (N_16954,N_16663,N_16644);
nand U16955 (N_16955,N_16526,N_16569);
nor U16956 (N_16956,N_16586,N_16617);
nand U16957 (N_16957,N_16532,N_16702);
xnor U16958 (N_16958,N_16597,N_16580);
or U16959 (N_16959,N_16658,N_16652);
and U16960 (N_16960,N_16611,N_16591);
and U16961 (N_16961,N_16513,N_16736);
nand U16962 (N_16962,N_16680,N_16573);
and U16963 (N_16963,N_16614,N_16597);
nor U16964 (N_16964,N_16621,N_16663);
and U16965 (N_16965,N_16648,N_16613);
nand U16966 (N_16966,N_16676,N_16598);
nor U16967 (N_16967,N_16538,N_16671);
nor U16968 (N_16968,N_16631,N_16557);
nor U16969 (N_16969,N_16713,N_16749);
xor U16970 (N_16970,N_16664,N_16720);
xnor U16971 (N_16971,N_16622,N_16509);
nor U16972 (N_16972,N_16709,N_16717);
or U16973 (N_16973,N_16504,N_16636);
nand U16974 (N_16974,N_16682,N_16615);
and U16975 (N_16975,N_16665,N_16612);
and U16976 (N_16976,N_16729,N_16744);
or U16977 (N_16977,N_16708,N_16675);
nand U16978 (N_16978,N_16644,N_16695);
or U16979 (N_16979,N_16602,N_16595);
nor U16980 (N_16980,N_16640,N_16629);
nand U16981 (N_16981,N_16548,N_16535);
and U16982 (N_16982,N_16603,N_16675);
xnor U16983 (N_16983,N_16718,N_16522);
nand U16984 (N_16984,N_16726,N_16576);
nor U16985 (N_16985,N_16528,N_16502);
nand U16986 (N_16986,N_16627,N_16578);
nand U16987 (N_16987,N_16644,N_16676);
and U16988 (N_16988,N_16581,N_16747);
xor U16989 (N_16989,N_16675,N_16524);
nor U16990 (N_16990,N_16534,N_16505);
xor U16991 (N_16991,N_16650,N_16739);
nand U16992 (N_16992,N_16641,N_16539);
nand U16993 (N_16993,N_16697,N_16715);
xnor U16994 (N_16994,N_16656,N_16515);
and U16995 (N_16995,N_16711,N_16506);
nor U16996 (N_16996,N_16698,N_16586);
or U16997 (N_16997,N_16564,N_16706);
and U16998 (N_16998,N_16527,N_16697);
xnor U16999 (N_16999,N_16580,N_16716);
nand U17000 (N_17000,N_16845,N_16825);
xnor U17001 (N_17001,N_16802,N_16852);
or U17002 (N_17002,N_16887,N_16913);
xnor U17003 (N_17003,N_16991,N_16958);
and U17004 (N_17004,N_16933,N_16854);
xnor U17005 (N_17005,N_16899,N_16920);
or U17006 (N_17006,N_16773,N_16951);
and U17007 (N_17007,N_16925,N_16981);
or U17008 (N_17008,N_16890,N_16964);
nor U17009 (N_17009,N_16829,N_16885);
nand U17010 (N_17010,N_16918,N_16978);
xnor U17011 (N_17011,N_16774,N_16987);
or U17012 (N_17012,N_16752,N_16772);
or U17013 (N_17013,N_16908,N_16786);
and U17014 (N_17014,N_16777,N_16916);
nor U17015 (N_17015,N_16804,N_16841);
nor U17016 (N_17016,N_16873,N_16766);
and U17017 (N_17017,N_16901,N_16868);
nand U17018 (N_17018,N_16831,N_16930);
nand U17019 (N_17019,N_16986,N_16805);
and U17020 (N_17020,N_16988,N_16921);
and U17021 (N_17021,N_16932,N_16917);
and U17022 (N_17022,N_16946,N_16886);
or U17023 (N_17023,N_16803,N_16943);
or U17024 (N_17024,N_16770,N_16832);
and U17025 (N_17025,N_16843,N_16960);
nand U17026 (N_17026,N_16848,N_16827);
nor U17027 (N_17027,N_16788,N_16850);
and U17028 (N_17028,N_16993,N_16999);
xnor U17029 (N_17029,N_16979,N_16959);
xnor U17030 (N_17030,N_16900,N_16956);
nor U17031 (N_17031,N_16976,N_16775);
nor U17032 (N_17032,N_16792,N_16859);
nand U17033 (N_17033,N_16794,N_16838);
or U17034 (N_17034,N_16781,N_16862);
xnor U17035 (N_17035,N_16938,N_16814);
nand U17036 (N_17036,N_16799,N_16934);
xor U17037 (N_17037,N_16888,N_16973);
nand U17038 (N_17038,N_16871,N_16812);
xnor U17039 (N_17039,N_16961,N_16893);
nand U17040 (N_17040,N_16936,N_16904);
or U17041 (N_17041,N_16818,N_16785);
and U17042 (N_17042,N_16968,N_16911);
and U17043 (N_17043,N_16778,N_16791);
nor U17044 (N_17044,N_16974,N_16820);
nand U17045 (N_17045,N_16977,N_16758);
nor U17046 (N_17046,N_16753,N_16833);
xnor U17047 (N_17047,N_16881,N_16879);
or U17048 (N_17048,N_16878,N_16822);
nor U17049 (N_17049,N_16861,N_16909);
nor U17050 (N_17050,N_16947,N_16962);
and U17051 (N_17051,N_16903,N_16950);
and U17052 (N_17052,N_16857,N_16948);
nor U17053 (N_17053,N_16898,N_16839);
or U17054 (N_17054,N_16902,N_16755);
nor U17055 (N_17055,N_16905,N_16765);
and U17056 (N_17056,N_16874,N_16895);
xor U17057 (N_17057,N_16809,N_16860);
xor U17058 (N_17058,N_16894,N_16759);
nor U17059 (N_17059,N_16844,N_16761);
or U17060 (N_17060,N_16966,N_16883);
xnor U17061 (N_17061,N_16996,N_16750);
or U17062 (N_17062,N_16782,N_16880);
and U17063 (N_17063,N_16931,N_16944);
or U17064 (N_17064,N_16790,N_16823);
or U17065 (N_17065,N_16935,N_16965);
xor U17066 (N_17066,N_16937,N_16967);
or U17067 (N_17067,N_16897,N_16824);
and U17068 (N_17068,N_16789,N_16942);
nand U17069 (N_17069,N_16762,N_16807);
xor U17070 (N_17070,N_16754,N_16994);
nand U17071 (N_17071,N_16847,N_16858);
and U17072 (N_17072,N_16787,N_16940);
or U17073 (N_17073,N_16779,N_16983);
xnor U17074 (N_17074,N_16768,N_16853);
or U17075 (N_17075,N_16801,N_16896);
nor U17076 (N_17076,N_16776,N_16875);
xnor U17077 (N_17077,N_16828,N_16953);
or U17078 (N_17078,N_16813,N_16995);
or U17079 (N_17079,N_16760,N_16751);
xnor U17080 (N_17080,N_16798,N_16830);
and U17081 (N_17081,N_16949,N_16914);
nor U17082 (N_17082,N_16941,N_16855);
nand U17083 (N_17083,N_16876,N_16763);
or U17084 (N_17084,N_16926,N_16846);
nand U17085 (N_17085,N_16872,N_16797);
nand U17086 (N_17086,N_16923,N_16757);
nor U17087 (N_17087,N_16954,N_16984);
nor U17088 (N_17088,N_16919,N_16882);
xnor U17089 (N_17089,N_16769,N_16922);
nor U17090 (N_17090,N_16971,N_16834);
and U17091 (N_17091,N_16907,N_16836);
or U17092 (N_17092,N_16992,N_16819);
and U17093 (N_17093,N_16963,N_16815);
nor U17094 (N_17094,N_16800,N_16835);
or U17095 (N_17095,N_16945,N_16806);
or U17096 (N_17096,N_16877,N_16865);
or U17097 (N_17097,N_16884,N_16864);
nor U17098 (N_17098,N_16928,N_16891);
xnor U17099 (N_17099,N_16906,N_16793);
xor U17100 (N_17100,N_16811,N_16990);
nor U17101 (N_17101,N_16910,N_16851);
or U17102 (N_17102,N_16985,N_16816);
and U17103 (N_17103,N_16795,N_16970);
and U17104 (N_17104,N_16784,N_16771);
xnor U17105 (N_17105,N_16840,N_16808);
or U17106 (N_17106,N_16767,N_16764);
nor U17107 (N_17107,N_16927,N_16842);
nor U17108 (N_17108,N_16870,N_16939);
nor U17109 (N_17109,N_16892,N_16869);
or U17110 (N_17110,N_16780,N_16821);
nand U17111 (N_17111,N_16866,N_16783);
nor U17112 (N_17112,N_16826,N_16955);
nand U17113 (N_17113,N_16863,N_16989);
nand U17114 (N_17114,N_16912,N_16997);
nand U17115 (N_17115,N_16924,N_16756);
and U17116 (N_17116,N_16982,N_16952);
xor U17117 (N_17117,N_16915,N_16837);
nor U17118 (N_17118,N_16810,N_16969);
or U17119 (N_17119,N_16972,N_16998);
or U17120 (N_17120,N_16867,N_16817);
or U17121 (N_17121,N_16856,N_16980);
xnor U17122 (N_17122,N_16796,N_16849);
nor U17123 (N_17123,N_16975,N_16929);
nand U17124 (N_17124,N_16889,N_16957);
and U17125 (N_17125,N_16943,N_16902);
nor U17126 (N_17126,N_16936,N_16762);
or U17127 (N_17127,N_16919,N_16765);
xnor U17128 (N_17128,N_16827,N_16885);
nor U17129 (N_17129,N_16958,N_16961);
xnor U17130 (N_17130,N_16981,N_16783);
nand U17131 (N_17131,N_16977,N_16850);
nor U17132 (N_17132,N_16888,N_16883);
and U17133 (N_17133,N_16882,N_16868);
nand U17134 (N_17134,N_16956,N_16841);
nor U17135 (N_17135,N_16758,N_16871);
nand U17136 (N_17136,N_16984,N_16910);
and U17137 (N_17137,N_16841,N_16853);
nor U17138 (N_17138,N_16854,N_16877);
or U17139 (N_17139,N_16824,N_16868);
nand U17140 (N_17140,N_16849,N_16989);
and U17141 (N_17141,N_16973,N_16843);
nor U17142 (N_17142,N_16971,N_16810);
and U17143 (N_17143,N_16878,N_16869);
or U17144 (N_17144,N_16877,N_16812);
xnor U17145 (N_17145,N_16967,N_16872);
or U17146 (N_17146,N_16838,N_16922);
nor U17147 (N_17147,N_16988,N_16853);
or U17148 (N_17148,N_16955,N_16804);
xnor U17149 (N_17149,N_16755,N_16757);
nand U17150 (N_17150,N_16908,N_16886);
xor U17151 (N_17151,N_16936,N_16953);
xor U17152 (N_17152,N_16757,N_16937);
and U17153 (N_17153,N_16912,N_16821);
nor U17154 (N_17154,N_16818,N_16934);
xnor U17155 (N_17155,N_16935,N_16945);
nor U17156 (N_17156,N_16768,N_16914);
nor U17157 (N_17157,N_16826,N_16829);
or U17158 (N_17158,N_16910,N_16921);
and U17159 (N_17159,N_16811,N_16837);
and U17160 (N_17160,N_16902,N_16947);
nor U17161 (N_17161,N_16761,N_16770);
xor U17162 (N_17162,N_16909,N_16951);
nand U17163 (N_17163,N_16916,N_16849);
or U17164 (N_17164,N_16950,N_16817);
or U17165 (N_17165,N_16770,N_16986);
or U17166 (N_17166,N_16976,N_16867);
xor U17167 (N_17167,N_16946,N_16757);
or U17168 (N_17168,N_16771,N_16758);
nor U17169 (N_17169,N_16917,N_16887);
nand U17170 (N_17170,N_16811,N_16932);
nor U17171 (N_17171,N_16880,N_16779);
xor U17172 (N_17172,N_16851,N_16941);
or U17173 (N_17173,N_16915,N_16908);
nor U17174 (N_17174,N_16896,N_16829);
or U17175 (N_17175,N_16937,N_16859);
nor U17176 (N_17176,N_16838,N_16964);
or U17177 (N_17177,N_16888,N_16916);
or U17178 (N_17178,N_16928,N_16955);
and U17179 (N_17179,N_16880,N_16845);
xor U17180 (N_17180,N_16856,N_16913);
or U17181 (N_17181,N_16994,N_16758);
nor U17182 (N_17182,N_16915,N_16939);
nand U17183 (N_17183,N_16834,N_16963);
nand U17184 (N_17184,N_16978,N_16928);
xor U17185 (N_17185,N_16985,N_16836);
nor U17186 (N_17186,N_16851,N_16928);
or U17187 (N_17187,N_16849,N_16876);
nor U17188 (N_17188,N_16979,N_16756);
and U17189 (N_17189,N_16831,N_16960);
nand U17190 (N_17190,N_16751,N_16861);
xor U17191 (N_17191,N_16943,N_16842);
or U17192 (N_17192,N_16967,N_16809);
and U17193 (N_17193,N_16999,N_16786);
xnor U17194 (N_17194,N_16962,N_16973);
nand U17195 (N_17195,N_16912,N_16862);
xor U17196 (N_17196,N_16994,N_16995);
and U17197 (N_17197,N_16805,N_16763);
or U17198 (N_17198,N_16914,N_16826);
nor U17199 (N_17199,N_16951,N_16767);
nand U17200 (N_17200,N_16964,N_16919);
and U17201 (N_17201,N_16768,N_16844);
or U17202 (N_17202,N_16944,N_16887);
nand U17203 (N_17203,N_16985,N_16925);
and U17204 (N_17204,N_16886,N_16912);
nor U17205 (N_17205,N_16918,N_16776);
nand U17206 (N_17206,N_16946,N_16881);
nor U17207 (N_17207,N_16898,N_16913);
nor U17208 (N_17208,N_16957,N_16818);
nand U17209 (N_17209,N_16824,N_16864);
xnor U17210 (N_17210,N_16963,N_16914);
nor U17211 (N_17211,N_16833,N_16832);
nor U17212 (N_17212,N_16845,N_16820);
xnor U17213 (N_17213,N_16853,N_16774);
nand U17214 (N_17214,N_16918,N_16762);
nor U17215 (N_17215,N_16799,N_16960);
nor U17216 (N_17216,N_16950,N_16791);
nor U17217 (N_17217,N_16804,N_16871);
and U17218 (N_17218,N_16888,N_16831);
nor U17219 (N_17219,N_16899,N_16891);
and U17220 (N_17220,N_16967,N_16995);
or U17221 (N_17221,N_16966,N_16996);
and U17222 (N_17222,N_16905,N_16781);
or U17223 (N_17223,N_16897,N_16848);
xnor U17224 (N_17224,N_16929,N_16767);
xor U17225 (N_17225,N_16981,N_16988);
and U17226 (N_17226,N_16752,N_16807);
nor U17227 (N_17227,N_16878,N_16796);
nor U17228 (N_17228,N_16928,N_16939);
nor U17229 (N_17229,N_16840,N_16865);
and U17230 (N_17230,N_16860,N_16991);
nand U17231 (N_17231,N_16802,N_16879);
xor U17232 (N_17232,N_16892,N_16800);
nor U17233 (N_17233,N_16981,N_16894);
or U17234 (N_17234,N_16805,N_16785);
or U17235 (N_17235,N_16792,N_16797);
nand U17236 (N_17236,N_16911,N_16805);
or U17237 (N_17237,N_16779,N_16947);
and U17238 (N_17238,N_16943,N_16829);
and U17239 (N_17239,N_16973,N_16945);
and U17240 (N_17240,N_16814,N_16920);
or U17241 (N_17241,N_16941,N_16891);
nor U17242 (N_17242,N_16829,N_16854);
nor U17243 (N_17243,N_16884,N_16997);
xor U17244 (N_17244,N_16793,N_16761);
nor U17245 (N_17245,N_16750,N_16804);
nor U17246 (N_17246,N_16935,N_16757);
nor U17247 (N_17247,N_16832,N_16765);
nand U17248 (N_17248,N_16943,N_16912);
or U17249 (N_17249,N_16889,N_16766);
or U17250 (N_17250,N_17154,N_17135);
xor U17251 (N_17251,N_17189,N_17121);
and U17252 (N_17252,N_17194,N_17146);
xnor U17253 (N_17253,N_17045,N_17010);
nand U17254 (N_17254,N_17230,N_17148);
nand U17255 (N_17255,N_17171,N_17035);
and U17256 (N_17256,N_17072,N_17007);
nor U17257 (N_17257,N_17211,N_17044);
and U17258 (N_17258,N_17028,N_17206);
nand U17259 (N_17259,N_17084,N_17120);
nor U17260 (N_17260,N_17107,N_17223);
nor U17261 (N_17261,N_17021,N_17181);
nor U17262 (N_17262,N_17017,N_17060);
and U17263 (N_17263,N_17124,N_17221);
xnor U17264 (N_17264,N_17083,N_17052);
or U17265 (N_17265,N_17051,N_17064);
xor U17266 (N_17266,N_17094,N_17020);
xnor U17267 (N_17267,N_17100,N_17022);
and U17268 (N_17268,N_17165,N_17109);
nand U17269 (N_17269,N_17113,N_17208);
and U17270 (N_17270,N_17138,N_17011);
nand U17271 (N_17271,N_17000,N_17248);
or U17272 (N_17272,N_17136,N_17046);
and U17273 (N_17273,N_17015,N_17199);
and U17274 (N_17274,N_17106,N_17166);
or U17275 (N_17275,N_17085,N_17133);
xnor U17276 (N_17276,N_17229,N_17184);
xor U17277 (N_17277,N_17155,N_17246);
nand U17278 (N_17278,N_17188,N_17200);
and U17279 (N_17279,N_17212,N_17145);
or U17280 (N_17280,N_17164,N_17231);
xor U17281 (N_17281,N_17102,N_17070);
nand U17282 (N_17282,N_17243,N_17218);
nand U17283 (N_17283,N_17043,N_17012);
or U17284 (N_17284,N_17203,N_17047);
nand U17285 (N_17285,N_17003,N_17234);
xnor U17286 (N_17286,N_17233,N_17098);
or U17287 (N_17287,N_17095,N_17096);
nand U17288 (N_17288,N_17023,N_17108);
or U17289 (N_17289,N_17141,N_17013);
xor U17290 (N_17290,N_17071,N_17244);
nor U17291 (N_17291,N_17175,N_17116);
and U17292 (N_17292,N_17139,N_17160);
and U17293 (N_17293,N_17048,N_17176);
or U17294 (N_17294,N_17009,N_17073);
nand U17295 (N_17295,N_17127,N_17059);
nor U17296 (N_17296,N_17219,N_17092);
and U17297 (N_17297,N_17173,N_17152);
xor U17298 (N_17298,N_17032,N_17147);
nand U17299 (N_17299,N_17110,N_17215);
xor U17300 (N_17300,N_17119,N_17065);
or U17301 (N_17301,N_17174,N_17207);
xnor U17302 (N_17302,N_17226,N_17104);
nor U17303 (N_17303,N_17036,N_17132);
or U17304 (N_17304,N_17025,N_17190);
xnor U17305 (N_17305,N_17140,N_17042);
nor U17306 (N_17306,N_17056,N_17126);
xnor U17307 (N_17307,N_17187,N_17201);
or U17308 (N_17308,N_17205,N_17038);
and U17309 (N_17309,N_17074,N_17241);
nor U17310 (N_17310,N_17178,N_17237);
or U17311 (N_17311,N_17099,N_17128);
nand U17312 (N_17312,N_17118,N_17123);
nand U17313 (N_17313,N_17101,N_17058);
nand U17314 (N_17314,N_17076,N_17202);
and U17315 (N_17315,N_17090,N_17129);
nand U17316 (N_17316,N_17170,N_17180);
and U17317 (N_17317,N_17034,N_17182);
or U17318 (N_17318,N_17239,N_17004);
or U17319 (N_17319,N_17002,N_17087);
xnor U17320 (N_17320,N_17143,N_17050);
xnor U17321 (N_17321,N_17097,N_17213);
nand U17322 (N_17322,N_17049,N_17008);
or U17323 (N_17323,N_17069,N_17168);
nor U17324 (N_17324,N_17225,N_17169);
nor U17325 (N_17325,N_17209,N_17001);
nor U17326 (N_17326,N_17242,N_17112);
xnor U17327 (N_17327,N_17247,N_17193);
or U17328 (N_17328,N_17054,N_17019);
xor U17329 (N_17329,N_17066,N_17086);
nand U17330 (N_17330,N_17005,N_17158);
nor U17331 (N_17331,N_17068,N_17216);
or U17332 (N_17332,N_17024,N_17082);
nor U17333 (N_17333,N_17238,N_17142);
nand U17334 (N_17334,N_17183,N_17131);
and U17335 (N_17335,N_17220,N_17033);
nand U17336 (N_17336,N_17227,N_17204);
and U17337 (N_17337,N_17039,N_17186);
nor U17338 (N_17338,N_17079,N_17016);
nand U17339 (N_17339,N_17235,N_17157);
nand U17340 (N_17340,N_17197,N_17198);
nand U17341 (N_17341,N_17130,N_17114);
and U17342 (N_17342,N_17149,N_17093);
and U17343 (N_17343,N_17117,N_17026);
nor U17344 (N_17344,N_17177,N_17185);
and U17345 (N_17345,N_17228,N_17111);
or U17346 (N_17346,N_17195,N_17057);
and U17347 (N_17347,N_17192,N_17249);
and U17348 (N_17348,N_17089,N_17030);
and U17349 (N_17349,N_17103,N_17232);
and U17350 (N_17350,N_17217,N_17134);
nor U17351 (N_17351,N_17091,N_17063);
and U17352 (N_17352,N_17037,N_17159);
nor U17353 (N_17353,N_17115,N_17162);
xnor U17354 (N_17354,N_17027,N_17078);
xnor U17355 (N_17355,N_17014,N_17061);
and U17356 (N_17356,N_17053,N_17161);
nor U17357 (N_17357,N_17210,N_17041);
nand U17358 (N_17358,N_17075,N_17179);
and U17359 (N_17359,N_17125,N_17151);
nand U17360 (N_17360,N_17080,N_17167);
xnor U17361 (N_17361,N_17214,N_17018);
or U17362 (N_17362,N_17150,N_17236);
xnor U17363 (N_17363,N_17062,N_17067);
and U17364 (N_17364,N_17077,N_17122);
nand U17365 (N_17365,N_17031,N_17163);
or U17366 (N_17366,N_17222,N_17245);
nor U17367 (N_17367,N_17105,N_17137);
nor U17368 (N_17368,N_17224,N_17088);
nor U17369 (N_17369,N_17240,N_17081);
xor U17370 (N_17370,N_17191,N_17055);
and U17371 (N_17371,N_17156,N_17029);
and U17372 (N_17372,N_17040,N_17144);
nor U17373 (N_17373,N_17006,N_17172);
nor U17374 (N_17374,N_17153,N_17196);
or U17375 (N_17375,N_17126,N_17229);
or U17376 (N_17376,N_17058,N_17139);
xor U17377 (N_17377,N_17162,N_17106);
nand U17378 (N_17378,N_17052,N_17053);
nand U17379 (N_17379,N_17056,N_17017);
or U17380 (N_17380,N_17110,N_17227);
nand U17381 (N_17381,N_17142,N_17139);
nor U17382 (N_17382,N_17218,N_17231);
and U17383 (N_17383,N_17104,N_17092);
and U17384 (N_17384,N_17145,N_17120);
nor U17385 (N_17385,N_17055,N_17008);
and U17386 (N_17386,N_17120,N_17024);
nand U17387 (N_17387,N_17082,N_17225);
and U17388 (N_17388,N_17008,N_17186);
nand U17389 (N_17389,N_17040,N_17242);
or U17390 (N_17390,N_17108,N_17215);
nor U17391 (N_17391,N_17203,N_17075);
and U17392 (N_17392,N_17220,N_17083);
nand U17393 (N_17393,N_17133,N_17049);
nor U17394 (N_17394,N_17122,N_17034);
and U17395 (N_17395,N_17152,N_17120);
xor U17396 (N_17396,N_17161,N_17114);
and U17397 (N_17397,N_17099,N_17173);
or U17398 (N_17398,N_17246,N_17093);
or U17399 (N_17399,N_17231,N_17138);
nand U17400 (N_17400,N_17159,N_17176);
nor U17401 (N_17401,N_17010,N_17184);
or U17402 (N_17402,N_17090,N_17221);
or U17403 (N_17403,N_17238,N_17237);
nor U17404 (N_17404,N_17063,N_17213);
and U17405 (N_17405,N_17114,N_17050);
or U17406 (N_17406,N_17093,N_17193);
nand U17407 (N_17407,N_17219,N_17196);
nor U17408 (N_17408,N_17134,N_17192);
nand U17409 (N_17409,N_17196,N_17123);
or U17410 (N_17410,N_17238,N_17015);
and U17411 (N_17411,N_17050,N_17214);
and U17412 (N_17412,N_17176,N_17018);
nand U17413 (N_17413,N_17021,N_17141);
nor U17414 (N_17414,N_17202,N_17246);
xor U17415 (N_17415,N_17053,N_17014);
nor U17416 (N_17416,N_17080,N_17149);
nand U17417 (N_17417,N_17080,N_17179);
nor U17418 (N_17418,N_17147,N_17083);
nand U17419 (N_17419,N_17052,N_17213);
and U17420 (N_17420,N_17118,N_17139);
nand U17421 (N_17421,N_17122,N_17096);
or U17422 (N_17422,N_17035,N_17000);
xor U17423 (N_17423,N_17025,N_17006);
nand U17424 (N_17424,N_17040,N_17169);
or U17425 (N_17425,N_17129,N_17031);
nor U17426 (N_17426,N_17209,N_17181);
and U17427 (N_17427,N_17112,N_17233);
nand U17428 (N_17428,N_17163,N_17165);
xor U17429 (N_17429,N_17208,N_17134);
and U17430 (N_17430,N_17133,N_17022);
nand U17431 (N_17431,N_17135,N_17152);
nand U17432 (N_17432,N_17083,N_17010);
or U17433 (N_17433,N_17004,N_17206);
and U17434 (N_17434,N_17088,N_17185);
nand U17435 (N_17435,N_17073,N_17144);
xor U17436 (N_17436,N_17206,N_17084);
and U17437 (N_17437,N_17082,N_17006);
or U17438 (N_17438,N_17073,N_17139);
nand U17439 (N_17439,N_17173,N_17161);
xor U17440 (N_17440,N_17069,N_17064);
xnor U17441 (N_17441,N_17222,N_17157);
and U17442 (N_17442,N_17007,N_17099);
nor U17443 (N_17443,N_17007,N_17117);
and U17444 (N_17444,N_17109,N_17115);
or U17445 (N_17445,N_17232,N_17089);
nor U17446 (N_17446,N_17166,N_17129);
xor U17447 (N_17447,N_17219,N_17211);
and U17448 (N_17448,N_17119,N_17185);
xor U17449 (N_17449,N_17143,N_17136);
xnor U17450 (N_17450,N_17053,N_17201);
nor U17451 (N_17451,N_17160,N_17133);
nand U17452 (N_17452,N_17150,N_17049);
nand U17453 (N_17453,N_17042,N_17027);
and U17454 (N_17454,N_17085,N_17016);
or U17455 (N_17455,N_17231,N_17095);
or U17456 (N_17456,N_17229,N_17066);
xnor U17457 (N_17457,N_17013,N_17096);
xor U17458 (N_17458,N_17004,N_17176);
or U17459 (N_17459,N_17130,N_17017);
nand U17460 (N_17460,N_17073,N_17058);
xnor U17461 (N_17461,N_17244,N_17222);
and U17462 (N_17462,N_17144,N_17206);
nand U17463 (N_17463,N_17067,N_17057);
and U17464 (N_17464,N_17086,N_17007);
nand U17465 (N_17465,N_17199,N_17155);
and U17466 (N_17466,N_17031,N_17127);
and U17467 (N_17467,N_17174,N_17114);
xor U17468 (N_17468,N_17021,N_17228);
nand U17469 (N_17469,N_17057,N_17138);
and U17470 (N_17470,N_17242,N_17016);
xnor U17471 (N_17471,N_17213,N_17117);
nor U17472 (N_17472,N_17031,N_17083);
xnor U17473 (N_17473,N_17085,N_17243);
and U17474 (N_17474,N_17173,N_17182);
nand U17475 (N_17475,N_17182,N_17089);
and U17476 (N_17476,N_17237,N_17139);
xnor U17477 (N_17477,N_17109,N_17102);
or U17478 (N_17478,N_17022,N_17023);
nor U17479 (N_17479,N_17168,N_17102);
and U17480 (N_17480,N_17109,N_17200);
or U17481 (N_17481,N_17046,N_17069);
nand U17482 (N_17482,N_17197,N_17065);
nor U17483 (N_17483,N_17219,N_17086);
nand U17484 (N_17484,N_17241,N_17036);
and U17485 (N_17485,N_17109,N_17072);
nor U17486 (N_17486,N_17004,N_17085);
xor U17487 (N_17487,N_17104,N_17085);
nand U17488 (N_17488,N_17167,N_17115);
and U17489 (N_17489,N_17010,N_17091);
and U17490 (N_17490,N_17181,N_17001);
nand U17491 (N_17491,N_17111,N_17121);
or U17492 (N_17492,N_17238,N_17164);
or U17493 (N_17493,N_17137,N_17061);
nand U17494 (N_17494,N_17049,N_17016);
xnor U17495 (N_17495,N_17121,N_17155);
nor U17496 (N_17496,N_17063,N_17050);
xor U17497 (N_17497,N_17187,N_17197);
nor U17498 (N_17498,N_17072,N_17167);
xor U17499 (N_17499,N_17209,N_17190);
nand U17500 (N_17500,N_17363,N_17478);
xor U17501 (N_17501,N_17436,N_17379);
nand U17502 (N_17502,N_17450,N_17485);
or U17503 (N_17503,N_17497,N_17403);
and U17504 (N_17504,N_17285,N_17369);
or U17505 (N_17505,N_17417,N_17481);
and U17506 (N_17506,N_17418,N_17428);
and U17507 (N_17507,N_17374,N_17250);
and U17508 (N_17508,N_17288,N_17267);
and U17509 (N_17509,N_17471,N_17316);
xor U17510 (N_17510,N_17360,N_17333);
xnor U17511 (N_17511,N_17387,N_17454);
nor U17512 (N_17512,N_17272,N_17466);
and U17513 (N_17513,N_17282,N_17358);
or U17514 (N_17514,N_17266,N_17270);
nand U17515 (N_17515,N_17435,N_17364);
or U17516 (N_17516,N_17313,N_17396);
or U17517 (N_17517,N_17488,N_17355);
xor U17518 (N_17518,N_17460,N_17354);
nor U17519 (N_17519,N_17294,N_17440);
nand U17520 (N_17520,N_17477,N_17271);
and U17521 (N_17521,N_17377,N_17386);
nand U17522 (N_17522,N_17317,N_17468);
nor U17523 (N_17523,N_17397,N_17431);
nand U17524 (N_17524,N_17367,N_17342);
xnor U17525 (N_17525,N_17262,N_17498);
xnor U17526 (N_17526,N_17390,N_17305);
and U17527 (N_17527,N_17463,N_17320);
nand U17528 (N_17528,N_17456,N_17251);
and U17529 (N_17529,N_17307,N_17437);
nand U17530 (N_17530,N_17411,N_17395);
nand U17531 (N_17531,N_17323,N_17337);
and U17532 (N_17532,N_17274,N_17472);
xnor U17533 (N_17533,N_17489,N_17314);
nand U17534 (N_17534,N_17309,N_17448);
and U17535 (N_17535,N_17293,N_17301);
nor U17536 (N_17536,N_17325,N_17341);
or U17537 (N_17537,N_17365,N_17384);
xnor U17538 (N_17538,N_17493,N_17286);
and U17539 (N_17539,N_17302,N_17407);
nor U17540 (N_17540,N_17328,N_17308);
nand U17541 (N_17541,N_17289,N_17373);
nor U17542 (N_17542,N_17370,N_17495);
nand U17543 (N_17543,N_17453,N_17259);
nand U17544 (N_17544,N_17346,N_17296);
and U17545 (N_17545,N_17421,N_17359);
nor U17546 (N_17546,N_17290,N_17283);
and U17547 (N_17547,N_17393,N_17347);
and U17548 (N_17548,N_17414,N_17479);
nor U17549 (N_17549,N_17388,N_17258);
nor U17550 (N_17550,N_17327,N_17281);
or U17551 (N_17551,N_17280,N_17306);
nand U17552 (N_17552,N_17459,N_17398);
nor U17553 (N_17553,N_17315,N_17461);
nand U17554 (N_17554,N_17254,N_17394);
or U17555 (N_17555,N_17300,N_17438);
xor U17556 (N_17556,N_17442,N_17449);
nor U17557 (N_17557,N_17492,N_17462);
xnor U17558 (N_17558,N_17429,N_17380);
nand U17559 (N_17559,N_17298,N_17464);
and U17560 (N_17560,N_17439,N_17425);
xor U17561 (N_17561,N_17319,N_17279);
or U17562 (N_17562,N_17329,N_17265);
or U17563 (N_17563,N_17375,N_17484);
xor U17564 (N_17564,N_17292,N_17278);
xor U17565 (N_17565,N_17389,N_17295);
xor U17566 (N_17566,N_17352,N_17455);
and U17567 (N_17567,N_17297,N_17483);
nor U17568 (N_17568,N_17408,N_17322);
nor U17569 (N_17569,N_17392,N_17351);
or U17570 (N_17570,N_17255,N_17399);
and U17571 (N_17571,N_17423,N_17339);
or U17572 (N_17572,N_17496,N_17349);
and U17573 (N_17573,N_17366,N_17451);
nor U17574 (N_17574,N_17340,N_17268);
and U17575 (N_17575,N_17318,N_17264);
nand U17576 (N_17576,N_17304,N_17402);
nor U17577 (N_17577,N_17321,N_17273);
or U17578 (N_17578,N_17443,N_17330);
and U17579 (N_17579,N_17480,N_17311);
and U17580 (N_17580,N_17331,N_17332);
nand U17581 (N_17581,N_17263,N_17410);
xor U17582 (N_17582,N_17499,N_17382);
or U17583 (N_17583,N_17381,N_17412);
xnor U17584 (N_17584,N_17416,N_17470);
nor U17585 (N_17585,N_17474,N_17430);
nand U17586 (N_17586,N_17303,N_17345);
nor U17587 (N_17587,N_17487,N_17427);
and U17588 (N_17588,N_17269,N_17371);
and U17589 (N_17589,N_17362,N_17334);
nand U17590 (N_17590,N_17312,N_17275);
or U17591 (N_17591,N_17277,N_17383);
nand U17592 (N_17592,N_17446,N_17420);
xor U17593 (N_17593,N_17441,N_17256);
or U17594 (N_17594,N_17422,N_17465);
xor U17595 (N_17595,N_17434,N_17299);
and U17596 (N_17596,N_17473,N_17376);
and U17597 (N_17597,N_17494,N_17260);
and U17598 (N_17598,N_17257,N_17326);
xnor U17599 (N_17599,N_17424,N_17284);
and U17600 (N_17600,N_17291,N_17419);
or U17601 (N_17601,N_17490,N_17335);
or U17602 (N_17602,N_17336,N_17406);
nand U17603 (N_17603,N_17447,N_17324);
or U17604 (N_17604,N_17287,N_17445);
nand U17605 (N_17605,N_17458,N_17344);
nor U17606 (N_17606,N_17368,N_17432);
nand U17607 (N_17607,N_17253,N_17361);
nand U17608 (N_17608,N_17415,N_17353);
nand U17609 (N_17609,N_17476,N_17457);
or U17610 (N_17610,N_17404,N_17400);
nand U17611 (N_17611,N_17338,N_17350);
and U17612 (N_17612,N_17405,N_17475);
and U17613 (N_17613,N_17356,N_17252);
or U17614 (N_17614,N_17413,N_17469);
or U17615 (N_17615,N_17433,N_17378);
nand U17616 (N_17616,N_17276,N_17343);
and U17617 (N_17617,N_17385,N_17261);
nor U17618 (N_17618,N_17391,N_17444);
xnor U17619 (N_17619,N_17452,N_17486);
xnor U17620 (N_17620,N_17357,N_17348);
or U17621 (N_17621,N_17372,N_17426);
xnor U17622 (N_17622,N_17401,N_17491);
xor U17623 (N_17623,N_17409,N_17310);
nor U17624 (N_17624,N_17482,N_17467);
nor U17625 (N_17625,N_17322,N_17397);
nand U17626 (N_17626,N_17442,N_17391);
nand U17627 (N_17627,N_17356,N_17267);
nand U17628 (N_17628,N_17390,N_17256);
and U17629 (N_17629,N_17463,N_17348);
and U17630 (N_17630,N_17314,N_17343);
and U17631 (N_17631,N_17321,N_17421);
nand U17632 (N_17632,N_17338,N_17447);
nand U17633 (N_17633,N_17373,N_17341);
xor U17634 (N_17634,N_17396,N_17360);
nand U17635 (N_17635,N_17389,N_17414);
or U17636 (N_17636,N_17351,N_17298);
nor U17637 (N_17637,N_17379,N_17499);
or U17638 (N_17638,N_17266,N_17359);
nor U17639 (N_17639,N_17313,N_17376);
or U17640 (N_17640,N_17361,N_17337);
or U17641 (N_17641,N_17401,N_17422);
and U17642 (N_17642,N_17331,N_17453);
and U17643 (N_17643,N_17482,N_17393);
or U17644 (N_17644,N_17394,N_17392);
nor U17645 (N_17645,N_17319,N_17457);
nand U17646 (N_17646,N_17480,N_17448);
nand U17647 (N_17647,N_17374,N_17420);
or U17648 (N_17648,N_17388,N_17387);
nand U17649 (N_17649,N_17382,N_17440);
nand U17650 (N_17650,N_17394,N_17331);
nor U17651 (N_17651,N_17418,N_17354);
and U17652 (N_17652,N_17459,N_17253);
or U17653 (N_17653,N_17442,N_17334);
xnor U17654 (N_17654,N_17409,N_17450);
xor U17655 (N_17655,N_17366,N_17499);
nand U17656 (N_17656,N_17256,N_17338);
or U17657 (N_17657,N_17485,N_17346);
nand U17658 (N_17658,N_17427,N_17482);
nor U17659 (N_17659,N_17330,N_17360);
or U17660 (N_17660,N_17376,N_17315);
or U17661 (N_17661,N_17476,N_17478);
and U17662 (N_17662,N_17466,N_17343);
nor U17663 (N_17663,N_17479,N_17427);
xor U17664 (N_17664,N_17499,N_17472);
and U17665 (N_17665,N_17370,N_17361);
or U17666 (N_17666,N_17272,N_17351);
and U17667 (N_17667,N_17378,N_17493);
nor U17668 (N_17668,N_17490,N_17262);
or U17669 (N_17669,N_17333,N_17348);
or U17670 (N_17670,N_17263,N_17468);
and U17671 (N_17671,N_17304,N_17323);
and U17672 (N_17672,N_17403,N_17488);
nand U17673 (N_17673,N_17493,N_17447);
nand U17674 (N_17674,N_17361,N_17254);
nor U17675 (N_17675,N_17498,N_17449);
nand U17676 (N_17676,N_17271,N_17423);
or U17677 (N_17677,N_17479,N_17490);
nand U17678 (N_17678,N_17375,N_17323);
and U17679 (N_17679,N_17433,N_17434);
and U17680 (N_17680,N_17435,N_17292);
and U17681 (N_17681,N_17294,N_17407);
nor U17682 (N_17682,N_17334,N_17464);
nor U17683 (N_17683,N_17458,N_17363);
xnor U17684 (N_17684,N_17289,N_17323);
xnor U17685 (N_17685,N_17275,N_17336);
nand U17686 (N_17686,N_17404,N_17399);
nor U17687 (N_17687,N_17407,N_17273);
xor U17688 (N_17688,N_17483,N_17362);
xnor U17689 (N_17689,N_17412,N_17492);
and U17690 (N_17690,N_17332,N_17369);
or U17691 (N_17691,N_17415,N_17356);
nor U17692 (N_17692,N_17355,N_17347);
nand U17693 (N_17693,N_17368,N_17310);
nand U17694 (N_17694,N_17318,N_17377);
nor U17695 (N_17695,N_17253,N_17469);
or U17696 (N_17696,N_17372,N_17485);
xor U17697 (N_17697,N_17371,N_17344);
or U17698 (N_17698,N_17427,N_17495);
nand U17699 (N_17699,N_17305,N_17414);
and U17700 (N_17700,N_17416,N_17478);
xor U17701 (N_17701,N_17403,N_17401);
or U17702 (N_17702,N_17383,N_17338);
nor U17703 (N_17703,N_17394,N_17467);
nor U17704 (N_17704,N_17415,N_17306);
or U17705 (N_17705,N_17273,N_17259);
nand U17706 (N_17706,N_17496,N_17463);
nand U17707 (N_17707,N_17443,N_17334);
nor U17708 (N_17708,N_17295,N_17341);
nand U17709 (N_17709,N_17468,N_17453);
xor U17710 (N_17710,N_17498,N_17470);
xor U17711 (N_17711,N_17274,N_17269);
or U17712 (N_17712,N_17375,N_17315);
xnor U17713 (N_17713,N_17290,N_17301);
and U17714 (N_17714,N_17422,N_17308);
nand U17715 (N_17715,N_17450,N_17384);
xnor U17716 (N_17716,N_17438,N_17359);
or U17717 (N_17717,N_17338,N_17411);
and U17718 (N_17718,N_17489,N_17342);
nand U17719 (N_17719,N_17421,N_17354);
or U17720 (N_17720,N_17366,N_17278);
nor U17721 (N_17721,N_17444,N_17320);
nor U17722 (N_17722,N_17398,N_17332);
and U17723 (N_17723,N_17282,N_17269);
or U17724 (N_17724,N_17421,N_17378);
xnor U17725 (N_17725,N_17451,N_17483);
or U17726 (N_17726,N_17440,N_17271);
and U17727 (N_17727,N_17301,N_17410);
nor U17728 (N_17728,N_17495,N_17367);
or U17729 (N_17729,N_17363,N_17451);
nor U17730 (N_17730,N_17382,N_17497);
or U17731 (N_17731,N_17367,N_17289);
nand U17732 (N_17732,N_17296,N_17288);
and U17733 (N_17733,N_17437,N_17424);
xor U17734 (N_17734,N_17413,N_17268);
and U17735 (N_17735,N_17277,N_17439);
or U17736 (N_17736,N_17351,N_17442);
and U17737 (N_17737,N_17482,N_17270);
nor U17738 (N_17738,N_17424,N_17371);
nand U17739 (N_17739,N_17305,N_17410);
and U17740 (N_17740,N_17278,N_17401);
nor U17741 (N_17741,N_17307,N_17328);
xor U17742 (N_17742,N_17295,N_17461);
or U17743 (N_17743,N_17432,N_17403);
nor U17744 (N_17744,N_17266,N_17377);
nand U17745 (N_17745,N_17393,N_17277);
nor U17746 (N_17746,N_17441,N_17271);
nand U17747 (N_17747,N_17487,N_17252);
and U17748 (N_17748,N_17333,N_17479);
or U17749 (N_17749,N_17475,N_17348);
nand U17750 (N_17750,N_17641,N_17683);
nor U17751 (N_17751,N_17580,N_17688);
nand U17752 (N_17752,N_17560,N_17693);
and U17753 (N_17753,N_17749,N_17639);
xor U17754 (N_17754,N_17662,N_17674);
nand U17755 (N_17755,N_17739,N_17731);
and U17756 (N_17756,N_17540,N_17548);
nand U17757 (N_17757,N_17515,N_17655);
xnor U17758 (N_17758,N_17723,N_17546);
and U17759 (N_17759,N_17550,N_17737);
or U17760 (N_17760,N_17689,N_17503);
xor U17761 (N_17761,N_17627,N_17706);
nand U17762 (N_17762,N_17633,N_17525);
and U17763 (N_17763,N_17563,N_17623);
and U17764 (N_17764,N_17551,N_17680);
and U17765 (N_17765,N_17575,N_17556);
or U17766 (N_17766,N_17583,N_17602);
or U17767 (N_17767,N_17611,N_17539);
or U17768 (N_17768,N_17529,N_17507);
xor U17769 (N_17769,N_17506,N_17598);
xnor U17770 (N_17770,N_17610,N_17630);
nor U17771 (N_17771,N_17682,N_17678);
nand U17772 (N_17772,N_17606,N_17618);
nor U17773 (N_17773,N_17572,N_17586);
nand U17774 (N_17774,N_17660,N_17577);
nand U17775 (N_17775,N_17582,N_17579);
and U17776 (N_17776,N_17629,N_17526);
xnor U17777 (N_17777,N_17746,N_17576);
nor U17778 (N_17778,N_17535,N_17701);
or U17779 (N_17779,N_17700,N_17508);
or U17780 (N_17780,N_17541,N_17677);
xnor U17781 (N_17781,N_17542,N_17672);
or U17782 (N_17782,N_17523,N_17712);
xor U17783 (N_17783,N_17538,N_17621);
and U17784 (N_17784,N_17643,N_17620);
nor U17785 (N_17785,N_17511,N_17671);
or U17786 (N_17786,N_17645,N_17564);
xor U17787 (N_17787,N_17733,N_17686);
and U17788 (N_17788,N_17665,N_17625);
xnor U17789 (N_17789,N_17744,N_17636);
nor U17790 (N_17790,N_17615,N_17543);
nand U17791 (N_17791,N_17709,N_17527);
or U17792 (N_17792,N_17516,N_17567);
or U17793 (N_17793,N_17504,N_17510);
nor U17794 (N_17794,N_17715,N_17600);
nand U17795 (N_17795,N_17532,N_17558);
xnor U17796 (N_17796,N_17729,N_17631);
nor U17797 (N_17797,N_17666,N_17594);
and U17798 (N_17798,N_17726,N_17565);
nand U17799 (N_17799,N_17502,N_17617);
and U17800 (N_17800,N_17644,N_17705);
or U17801 (N_17801,N_17595,N_17584);
nand U17802 (N_17802,N_17651,N_17697);
nor U17803 (N_17803,N_17512,N_17696);
and U17804 (N_17804,N_17673,N_17652);
nor U17805 (N_17805,N_17741,N_17588);
xor U17806 (N_17806,N_17514,N_17509);
nor U17807 (N_17807,N_17581,N_17748);
xnor U17808 (N_17808,N_17647,N_17659);
and U17809 (N_17809,N_17518,N_17599);
nand U17810 (N_17810,N_17607,N_17690);
or U17811 (N_17811,N_17517,N_17533);
and U17812 (N_17812,N_17736,N_17707);
nor U17813 (N_17813,N_17691,N_17555);
nand U17814 (N_17814,N_17725,N_17520);
xnor U17815 (N_17815,N_17605,N_17613);
and U17816 (N_17816,N_17632,N_17571);
xor U17817 (N_17817,N_17521,N_17718);
nand U17818 (N_17818,N_17554,N_17717);
nand U17819 (N_17819,N_17708,N_17593);
and U17820 (N_17820,N_17528,N_17740);
or U17821 (N_17821,N_17663,N_17544);
nand U17822 (N_17822,N_17653,N_17640);
nand U17823 (N_17823,N_17537,N_17608);
or U17824 (N_17824,N_17743,N_17638);
nor U17825 (N_17825,N_17568,N_17679);
nand U17826 (N_17826,N_17648,N_17687);
or U17827 (N_17827,N_17658,N_17742);
xor U17828 (N_17828,N_17585,N_17616);
xor U17829 (N_17829,N_17724,N_17747);
xor U17830 (N_17830,N_17501,N_17698);
or U17831 (N_17831,N_17728,N_17668);
or U17832 (N_17832,N_17604,N_17552);
and U17833 (N_17833,N_17695,N_17589);
nor U17834 (N_17834,N_17549,N_17719);
xor U17835 (N_17835,N_17559,N_17553);
or U17836 (N_17836,N_17574,N_17675);
nor U17837 (N_17837,N_17745,N_17622);
nand U17838 (N_17838,N_17628,N_17557);
and U17839 (N_17839,N_17642,N_17650);
and U17840 (N_17840,N_17566,N_17596);
nor U17841 (N_17841,N_17505,N_17681);
and U17842 (N_17842,N_17614,N_17547);
and U17843 (N_17843,N_17624,N_17545);
or U17844 (N_17844,N_17626,N_17646);
nand U17845 (N_17845,N_17609,N_17722);
xnor U17846 (N_17846,N_17699,N_17710);
nor U17847 (N_17847,N_17587,N_17730);
nand U17848 (N_17848,N_17685,N_17735);
nor U17849 (N_17849,N_17694,N_17713);
nor U17850 (N_17850,N_17519,N_17714);
nand U17851 (N_17851,N_17601,N_17734);
nor U17852 (N_17852,N_17562,N_17654);
xor U17853 (N_17853,N_17603,N_17738);
xnor U17854 (N_17854,N_17570,N_17684);
nand U17855 (N_17855,N_17721,N_17561);
nor U17856 (N_17856,N_17513,N_17670);
nor U17857 (N_17857,N_17667,N_17711);
and U17858 (N_17858,N_17634,N_17656);
and U17859 (N_17859,N_17664,N_17703);
xor U17860 (N_17860,N_17569,N_17531);
xor U17861 (N_17861,N_17732,N_17524);
or U17862 (N_17862,N_17534,N_17676);
xor U17863 (N_17863,N_17720,N_17657);
or U17864 (N_17864,N_17635,N_17522);
xnor U17865 (N_17865,N_17573,N_17704);
nor U17866 (N_17866,N_17619,N_17702);
nand U17867 (N_17867,N_17536,N_17692);
and U17868 (N_17868,N_17637,N_17590);
and U17869 (N_17869,N_17500,N_17578);
nor U17870 (N_17870,N_17597,N_17592);
xor U17871 (N_17871,N_17669,N_17591);
and U17872 (N_17872,N_17649,N_17727);
nand U17873 (N_17873,N_17612,N_17661);
xor U17874 (N_17874,N_17716,N_17530);
xor U17875 (N_17875,N_17726,N_17635);
or U17876 (N_17876,N_17621,N_17540);
nor U17877 (N_17877,N_17600,N_17691);
nor U17878 (N_17878,N_17578,N_17692);
or U17879 (N_17879,N_17602,N_17701);
nand U17880 (N_17880,N_17654,N_17600);
or U17881 (N_17881,N_17552,N_17649);
and U17882 (N_17882,N_17540,N_17569);
nand U17883 (N_17883,N_17654,N_17724);
or U17884 (N_17884,N_17503,N_17731);
nand U17885 (N_17885,N_17731,N_17729);
nand U17886 (N_17886,N_17525,N_17686);
xnor U17887 (N_17887,N_17507,N_17637);
or U17888 (N_17888,N_17621,N_17602);
nor U17889 (N_17889,N_17535,N_17657);
and U17890 (N_17890,N_17719,N_17506);
nor U17891 (N_17891,N_17534,N_17511);
xnor U17892 (N_17892,N_17659,N_17731);
nor U17893 (N_17893,N_17707,N_17690);
nor U17894 (N_17894,N_17711,N_17624);
xor U17895 (N_17895,N_17529,N_17698);
nor U17896 (N_17896,N_17645,N_17573);
and U17897 (N_17897,N_17735,N_17617);
xor U17898 (N_17898,N_17643,N_17572);
or U17899 (N_17899,N_17680,N_17699);
xor U17900 (N_17900,N_17578,N_17511);
and U17901 (N_17901,N_17623,N_17564);
or U17902 (N_17902,N_17698,N_17604);
and U17903 (N_17903,N_17579,N_17721);
nand U17904 (N_17904,N_17541,N_17514);
xor U17905 (N_17905,N_17708,N_17637);
xor U17906 (N_17906,N_17532,N_17543);
and U17907 (N_17907,N_17528,N_17569);
xor U17908 (N_17908,N_17569,N_17678);
xor U17909 (N_17909,N_17546,N_17639);
and U17910 (N_17910,N_17685,N_17563);
nand U17911 (N_17911,N_17501,N_17541);
nor U17912 (N_17912,N_17625,N_17548);
nand U17913 (N_17913,N_17530,N_17721);
and U17914 (N_17914,N_17701,N_17507);
or U17915 (N_17915,N_17617,N_17555);
xnor U17916 (N_17916,N_17631,N_17516);
nor U17917 (N_17917,N_17505,N_17574);
nor U17918 (N_17918,N_17524,N_17694);
xnor U17919 (N_17919,N_17679,N_17646);
nor U17920 (N_17920,N_17692,N_17571);
xnor U17921 (N_17921,N_17717,N_17638);
or U17922 (N_17922,N_17654,N_17644);
and U17923 (N_17923,N_17731,N_17567);
and U17924 (N_17924,N_17680,N_17595);
and U17925 (N_17925,N_17565,N_17711);
or U17926 (N_17926,N_17585,N_17508);
or U17927 (N_17927,N_17704,N_17696);
nand U17928 (N_17928,N_17675,N_17636);
and U17929 (N_17929,N_17547,N_17559);
xnor U17930 (N_17930,N_17683,N_17508);
xnor U17931 (N_17931,N_17515,N_17536);
nor U17932 (N_17932,N_17517,N_17709);
nand U17933 (N_17933,N_17680,N_17591);
nand U17934 (N_17934,N_17650,N_17550);
nand U17935 (N_17935,N_17715,N_17671);
nor U17936 (N_17936,N_17683,N_17584);
nor U17937 (N_17937,N_17567,N_17730);
nand U17938 (N_17938,N_17552,N_17640);
nor U17939 (N_17939,N_17542,N_17728);
nor U17940 (N_17940,N_17604,N_17568);
nor U17941 (N_17941,N_17607,N_17747);
and U17942 (N_17942,N_17552,N_17713);
nor U17943 (N_17943,N_17632,N_17734);
nor U17944 (N_17944,N_17738,N_17727);
or U17945 (N_17945,N_17673,N_17707);
and U17946 (N_17946,N_17708,N_17728);
and U17947 (N_17947,N_17714,N_17606);
nor U17948 (N_17948,N_17566,N_17734);
xor U17949 (N_17949,N_17737,N_17573);
xor U17950 (N_17950,N_17705,N_17662);
or U17951 (N_17951,N_17540,N_17524);
xor U17952 (N_17952,N_17517,N_17551);
nor U17953 (N_17953,N_17732,N_17587);
nor U17954 (N_17954,N_17503,N_17571);
nand U17955 (N_17955,N_17573,N_17651);
nand U17956 (N_17956,N_17569,N_17625);
nor U17957 (N_17957,N_17623,N_17715);
nand U17958 (N_17958,N_17625,N_17526);
nor U17959 (N_17959,N_17552,N_17614);
and U17960 (N_17960,N_17565,N_17736);
xnor U17961 (N_17961,N_17615,N_17531);
xnor U17962 (N_17962,N_17583,N_17520);
xnor U17963 (N_17963,N_17746,N_17593);
and U17964 (N_17964,N_17622,N_17575);
nand U17965 (N_17965,N_17604,N_17539);
nor U17966 (N_17966,N_17662,N_17747);
or U17967 (N_17967,N_17624,N_17512);
or U17968 (N_17968,N_17509,N_17746);
nand U17969 (N_17969,N_17501,N_17727);
nand U17970 (N_17970,N_17652,N_17516);
nor U17971 (N_17971,N_17643,N_17691);
or U17972 (N_17972,N_17513,N_17688);
or U17973 (N_17973,N_17553,N_17629);
nor U17974 (N_17974,N_17600,N_17668);
nand U17975 (N_17975,N_17606,N_17599);
or U17976 (N_17976,N_17742,N_17688);
or U17977 (N_17977,N_17654,N_17608);
or U17978 (N_17978,N_17742,N_17508);
xnor U17979 (N_17979,N_17713,N_17733);
xor U17980 (N_17980,N_17520,N_17727);
and U17981 (N_17981,N_17629,N_17627);
nor U17982 (N_17982,N_17578,N_17517);
or U17983 (N_17983,N_17599,N_17649);
xnor U17984 (N_17984,N_17621,N_17713);
and U17985 (N_17985,N_17666,N_17654);
xnor U17986 (N_17986,N_17569,N_17697);
xor U17987 (N_17987,N_17684,N_17729);
nor U17988 (N_17988,N_17586,N_17512);
nand U17989 (N_17989,N_17718,N_17614);
nand U17990 (N_17990,N_17741,N_17509);
xnor U17991 (N_17991,N_17669,N_17746);
xor U17992 (N_17992,N_17584,N_17541);
xor U17993 (N_17993,N_17725,N_17630);
or U17994 (N_17994,N_17543,N_17644);
nor U17995 (N_17995,N_17501,N_17596);
nand U17996 (N_17996,N_17536,N_17721);
or U17997 (N_17997,N_17689,N_17502);
xnor U17998 (N_17998,N_17612,N_17543);
nor U17999 (N_17999,N_17572,N_17735);
nor U18000 (N_18000,N_17983,N_17780);
nand U18001 (N_18001,N_17908,N_17861);
nor U18002 (N_18002,N_17849,N_17797);
nor U18003 (N_18003,N_17787,N_17868);
or U18004 (N_18004,N_17781,N_17863);
nand U18005 (N_18005,N_17898,N_17977);
nand U18006 (N_18006,N_17967,N_17900);
and U18007 (N_18007,N_17776,N_17822);
or U18008 (N_18008,N_17915,N_17809);
or U18009 (N_18009,N_17974,N_17932);
nand U18010 (N_18010,N_17991,N_17790);
xor U18011 (N_18011,N_17812,N_17872);
nand U18012 (N_18012,N_17770,N_17938);
and U18013 (N_18013,N_17999,N_17876);
nor U18014 (N_18014,N_17851,N_17785);
and U18015 (N_18015,N_17981,N_17940);
nand U18016 (N_18016,N_17796,N_17950);
xor U18017 (N_18017,N_17802,N_17916);
nor U18018 (N_18018,N_17836,N_17899);
or U18019 (N_18019,N_17919,N_17995);
xnor U18020 (N_18020,N_17813,N_17841);
and U18021 (N_18021,N_17850,N_17779);
xnor U18022 (N_18022,N_17993,N_17988);
xnor U18023 (N_18023,N_17838,N_17910);
and U18024 (N_18024,N_17753,N_17979);
or U18025 (N_18025,N_17889,N_17829);
and U18026 (N_18026,N_17969,N_17904);
nand U18027 (N_18027,N_17965,N_17835);
nand U18028 (N_18028,N_17893,N_17807);
and U18029 (N_18029,N_17775,N_17754);
or U18030 (N_18030,N_17818,N_17973);
and U18031 (N_18031,N_17976,N_17852);
nor U18032 (N_18032,N_17857,N_17870);
nor U18033 (N_18033,N_17911,N_17824);
xor U18034 (N_18034,N_17843,N_17757);
xnor U18035 (N_18035,N_17946,N_17881);
nor U18036 (N_18036,N_17895,N_17992);
nand U18037 (N_18037,N_17806,N_17820);
xnor U18038 (N_18038,N_17817,N_17989);
nand U18039 (N_18039,N_17959,N_17941);
and U18040 (N_18040,N_17929,N_17943);
nor U18041 (N_18041,N_17887,N_17948);
xnor U18042 (N_18042,N_17846,N_17907);
xor U18043 (N_18043,N_17958,N_17833);
nand U18044 (N_18044,N_17853,N_17984);
nand U18045 (N_18045,N_17942,N_17926);
and U18046 (N_18046,N_17925,N_17762);
nor U18047 (N_18047,N_17971,N_17960);
nor U18048 (N_18048,N_17877,N_17874);
or U18049 (N_18049,N_17952,N_17772);
or U18050 (N_18050,N_17935,N_17882);
or U18051 (N_18051,N_17760,N_17901);
xor U18052 (N_18052,N_17964,N_17788);
xor U18053 (N_18053,N_17768,N_17801);
nand U18054 (N_18054,N_17982,N_17914);
nor U18055 (N_18055,N_17811,N_17860);
xnor U18056 (N_18056,N_17821,N_17842);
or U18057 (N_18057,N_17826,N_17962);
nand U18058 (N_18058,N_17786,N_17848);
nor U18059 (N_18059,N_17897,N_17830);
and U18060 (N_18060,N_17957,N_17794);
or U18061 (N_18061,N_17980,N_17771);
nand U18062 (N_18062,N_17751,N_17792);
xor U18063 (N_18063,N_17927,N_17905);
nand U18064 (N_18064,N_17782,N_17921);
or U18065 (N_18065,N_17875,N_17966);
xnor U18066 (N_18066,N_17756,N_17985);
or U18067 (N_18067,N_17918,N_17750);
and U18068 (N_18068,N_17862,N_17892);
nor U18069 (N_18069,N_17913,N_17855);
xnor U18070 (N_18070,N_17909,N_17944);
or U18071 (N_18071,N_17791,N_17945);
nor U18072 (N_18072,N_17752,N_17823);
and U18073 (N_18073,N_17784,N_17920);
and U18074 (N_18074,N_17924,N_17990);
or U18075 (N_18075,N_17890,N_17825);
and U18076 (N_18076,N_17922,N_17883);
nand U18077 (N_18077,N_17998,N_17769);
xnor U18078 (N_18078,N_17906,N_17902);
xor U18079 (N_18079,N_17814,N_17856);
xor U18080 (N_18080,N_17844,N_17763);
nor U18081 (N_18081,N_17759,N_17934);
xnor U18082 (N_18082,N_17947,N_17858);
and U18083 (N_18083,N_17956,N_17865);
xor U18084 (N_18084,N_17975,N_17903);
or U18085 (N_18085,N_17949,N_17837);
and U18086 (N_18086,N_17854,N_17933);
and U18087 (N_18087,N_17778,N_17783);
or U18088 (N_18088,N_17871,N_17972);
xnor U18089 (N_18089,N_17859,N_17799);
and U18090 (N_18090,N_17936,N_17832);
xnor U18091 (N_18091,N_17878,N_17994);
and U18092 (N_18092,N_17880,N_17758);
xnor U18093 (N_18093,N_17805,N_17886);
nor U18094 (N_18094,N_17867,N_17777);
nand U18095 (N_18095,N_17773,N_17831);
xnor U18096 (N_18096,N_17931,N_17978);
or U18097 (N_18097,N_17808,N_17798);
nand U18098 (N_18098,N_17970,N_17937);
and U18099 (N_18099,N_17839,N_17963);
nand U18100 (N_18100,N_17864,N_17986);
xor U18101 (N_18101,N_17793,N_17827);
or U18102 (N_18102,N_17939,N_17803);
or U18103 (N_18103,N_17996,N_17789);
or U18104 (N_18104,N_17928,N_17997);
nor U18105 (N_18105,N_17815,N_17800);
or U18106 (N_18106,N_17819,N_17896);
nor U18107 (N_18107,N_17884,N_17834);
xnor U18108 (N_18108,N_17894,N_17755);
nor U18109 (N_18109,N_17810,N_17767);
and U18110 (N_18110,N_17885,N_17774);
nor U18111 (N_18111,N_17873,N_17912);
nor U18112 (N_18112,N_17954,N_17845);
nand U18113 (N_18113,N_17761,N_17765);
nand U18114 (N_18114,N_17879,N_17968);
nor U18115 (N_18115,N_17930,N_17866);
nor U18116 (N_18116,N_17764,N_17953);
xor U18117 (N_18117,N_17888,N_17766);
nand U18118 (N_18118,N_17816,N_17955);
or U18119 (N_18119,N_17840,N_17987);
nand U18120 (N_18120,N_17828,N_17891);
and U18121 (N_18121,N_17795,N_17847);
and U18122 (N_18122,N_17961,N_17869);
xor U18123 (N_18123,N_17917,N_17951);
nor U18124 (N_18124,N_17923,N_17804);
nor U18125 (N_18125,N_17857,N_17916);
or U18126 (N_18126,N_17959,N_17798);
and U18127 (N_18127,N_17839,N_17779);
nand U18128 (N_18128,N_17828,N_17827);
xnor U18129 (N_18129,N_17975,N_17837);
nand U18130 (N_18130,N_17963,N_17954);
and U18131 (N_18131,N_17792,N_17847);
nand U18132 (N_18132,N_17970,N_17875);
nand U18133 (N_18133,N_17899,N_17830);
xor U18134 (N_18134,N_17853,N_17863);
nor U18135 (N_18135,N_17821,N_17827);
xor U18136 (N_18136,N_17820,N_17775);
and U18137 (N_18137,N_17801,N_17810);
and U18138 (N_18138,N_17837,N_17859);
nand U18139 (N_18139,N_17977,N_17961);
nand U18140 (N_18140,N_17947,N_17889);
nand U18141 (N_18141,N_17843,N_17839);
nand U18142 (N_18142,N_17836,N_17834);
or U18143 (N_18143,N_17965,N_17873);
xor U18144 (N_18144,N_17914,N_17768);
nor U18145 (N_18145,N_17771,N_17955);
or U18146 (N_18146,N_17796,N_17982);
xor U18147 (N_18147,N_17817,N_17901);
or U18148 (N_18148,N_17989,N_17924);
and U18149 (N_18149,N_17884,N_17918);
xor U18150 (N_18150,N_17784,N_17804);
nor U18151 (N_18151,N_17815,N_17982);
nand U18152 (N_18152,N_17842,N_17798);
nor U18153 (N_18153,N_17847,N_17773);
and U18154 (N_18154,N_17915,N_17752);
and U18155 (N_18155,N_17952,N_17756);
nor U18156 (N_18156,N_17808,N_17841);
and U18157 (N_18157,N_17864,N_17768);
xor U18158 (N_18158,N_17772,N_17861);
nand U18159 (N_18159,N_17875,N_17979);
or U18160 (N_18160,N_17974,N_17871);
xnor U18161 (N_18161,N_17858,N_17783);
nor U18162 (N_18162,N_17964,N_17889);
and U18163 (N_18163,N_17939,N_17762);
and U18164 (N_18164,N_17833,N_17917);
nor U18165 (N_18165,N_17808,N_17913);
xnor U18166 (N_18166,N_17972,N_17893);
or U18167 (N_18167,N_17976,N_17895);
or U18168 (N_18168,N_17791,N_17877);
nor U18169 (N_18169,N_17912,N_17816);
nor U18170 (N_18170,N_17934,N_17870);
nand U18171 (N_18171,N_17986,N_17800);
nor U18172 (N_18172,N_17817,N_17873);
xnor U18173 (N_18173,N_17766,N_17900);
or U18174 (N_18174,N_17856,N_17824);
nand U18175 (N_18175,N_17827,N_17826);
or U18176 (N_18176,N_17826,N_17940);
nor U18177 (N_18177,N_17796,N_17952);
or U18178 (N_18178,N_17873,N_17801);
or U18179 (N_18179,N_17818,N_17924);
nand U18180 (N_18180,N_17993,N_17974);
and U18181 (N_18181,N_17829,N_17934);
or U18182 (N_18182,N_17948,N_17760);
xnor U18183 (N_18183,N_17858,N_17878);
xor U18184 (N_18184,N_17889,N_17779);
or U18185 (N_18185,N_17953,N_17984);
and U18186 (N_18186,N_17773,N_17912);
and U18187 (N_18187,N_17763,N_17980);
xnor U18188 (N_18188,N_17917,N_17931);
nor U18189 (N_18189,N_17871,N_17885);
or U18190 (N_18190,N_17937,N_17941);
nand U18191 (N_18191,N_17952,N_17994);
nor U18192 (N_18192,N_17781,N_17771);
or U18193 (N_18193,N_17924,N_17782);
and U18194 (N_18194,N_17955,N_17981);
nor U18195 (N_18195,N_17993,N_17833);
or U18196 (N_18196,N_17948,N_17917);
xor U18197 (N_18197,N_17785,N_17965);
or U18198 (N_18198,N_17904,N_17756);
nand U18199 (N_18199,N_17830,N_17821);
and U18200 (N_18200,N_17904,N_17752);
nand U18201 (N_18201,N_17991,N_17750);
nor U18202 (N_18202,N_17909,N_17814);
nand U18203 (N_18203,N_17943,N_17908);
nor U18204 (N_18204,N_17943,N_17758);
or U18205 (N_18205,N_17890,N_17868);
xnor U18206 (N_18206,N_17950,N_17863);
nand U18207 (N_18207,N_17956,N_17887);
nor U18208 (N_18208,N_17785,N_17998);
or U18209 (N_18209,N_17989,N_17927);
or U18210 (N_18210,N_17779,N_17790);
nor U18211 (N_18211,N_17798,N_17904);
nor U18212 (N_18212,N_17993,N_17766);
or U18213 (N_18213,N_17862,N_17940);
nor U18214 (N_18214,N_17951,N_17878);
xor U18215 (N_18215,N_17850,N_17885);
xnor U18216 (N_18216,N_17781,N_17815);
nor U18217 (N_18217,N_17878,N_17947);
xnor U18218 (N_18218,N_17792,N_17892);
nor U18219 (N_18219,N_17921,N_17906);
xnor U18220 (N_18220,N_17949,N_17940);
or U18221 (N_18221,N_17841,N_17918);
xnor U18222 (N_18222,N_17797,N_17921);
xnor U18223 (N_18223,N_17970,N_17772);
nand U18224 (N_18224,N_17851,N_17853);
xnor U18225 (N_18225,N_17898,N_17802);
and U18226 (N_18226,N_17861,N_17986);
nor U18227 (N_18227,N_17939,N_17911);
nand U18228 (N_18228,N_17952,N_17813);
and U18229 (N_18229,N_17967,N_17910);
and U18230 (N_18230,N_17959,N_17913);
xnor U18231 (N_18231,N_17922,N_17812);
or U18232 (N_18232,N_17879,N_17958);
or U18233 (N_18233,N_17922,N_17890);
nand U18234 (N_18234,N_17849,N_17785);
and U18235 (N_18235,N_17898,N_17854);
or U18236 (N_18236,N_17929,N_17858);
and U18237 (N_18237,N_17964,N_17808);
nand U18238 (N_18238,N_17883,N_17888);
xor U18239 (N_18239,N_17760,N_17757);
and U18240 (N_18240,N_17880,N_17856);
xor U18241 (N_18241,N_17921,N_17761);
and U18242 (N_18242,N_17893,N_17815);
or U18243 (N_18243,N_17950,N_17960);
or U18244 (N_18244,N_17965,N_17894);
or U18245 (N_18245,N_17772,N_17808);
and U18246 (N_18246,N_17782,N_17937);
and U18247 (N_18247,N_17918,N_17752);
nor U18248 (N_18248,N_17891,N_17837);
xor U18249 (N_18249,N_17851,N_17761);
xnor U18250 (N_18250,N_18025,N_18036);
xor U18251 (N_18251,N_18143,N_18044);
or U18252 (N_18252,N_18165,N_18220);
and U18253 (N_18253,N_18139,N_18113);
or U18254 (N_18254,N_18146,N_18244);
nand U18255 (N_18255,N_18078,N_18156);
xnor U18256 (N_18256,N_18058,N_18248);
and U18257 (N_18257,N_18031,N_18116);
or U18258 (N_18258,N_18231,N_18006);
and U18259 (N_18259,N_18103,N_18134);
and U18260 (N_18260,N_18049,N_18135);
nor U18261 (N_18261,N_18069,N_18004);
or U18262 (N_18262,N_18083,N_18230);
and U18263 (N_18263,N_18092,N_18125);
nand U18264 (N_18264,N_18012,N_18182);
nand U18265 (N_18265,N_18054,N_18074);
and U18266 (N_18266,N_18038,N_18145);
xor U18267 (N_18267,N_18005,N_18216);
and U18268 (N_18268,N_18130,N_18114);
or U18269 (N_18269,N_18249,N_18105);
nor U18270 (N_18270,N_18077,N_18040);
nand U18271 (N_18271,N_18043,N_18007);
or U18272 (N_18272,N_18060,N_18093);
nor U18273 (N_18273,N_18213,N_18168);
nand U18274 (N_18274,N_18207,N_18067);
nor U18275 (N_18275,N_18023,N_18121);
nand U18276 (N_18276,N_18149,N_18141);
and U18277 (N_18277,N_18170,N_18097);
and U18278 (N_18278,N_18191,N_18172);
and U18279 (N_18279,N_18234,N_18064);
nand U18280 (N_18280,N_18223,N_18242);
nand U18281 (N_18281,N_18075,N_18238);
or U18282 (N_18282,N_18066,N_18022);
or U18283 (N_18283,N_18073,N_18072);
xor U18284 (N_18284,N_18164,N_18071);
and U18285 (N_18285,N_18039,N_18190);
and U18286 (N_18286,N_18112,N_18126);
and U18287 (N_18287,N_18186,N_18162);
nand U18288 (N_18288,N_18174,N_18118);
and U18289 (N_18289,N_18110,N_18133);
or U18290 (N_18290,N_18185,N_18026);
nor U18291 (N_18291,N_18035,N_18014);
xor U18292 (N_18292,N_18124,N_18193);
or U18293 (N_18293,N_18175,N_18240);
or U18294 (N_18294,N_18203,N_18001);
and U18295 (N_18295,N_18221,N_18048);
nand U18296 (N_18296,N_18153,N_18042);
xor U18297 (N_18297,N_18199,N_18187);
xor U18298 (N_18298,N_18120,N_18173);
nor U18299 (N_18299,N_18002,N_18087);
nor U18300 (N_18300,N_18089,N_18070);
nand U18301 (N_18301,N_18148,N_18013);
or U18302 (N_18302,N_18122,N_18151);
and U18303 (N_18303,N_18222,N_18056);
and U18304 (N_18304,N_18115,N_18102);
or U18305 (N_18305,N_18177,N_18217);
nor U18306 (N_18306,N_18018,N_18053);
nor U18307 (N_18307,N_18010,N_18076);
or U18308 (N_18308,N_18138,N_18119);
and U18309 (N_18309,N_18091,N_18210);
nor U18310 (N_18310,N_18196,N_18080);
xnor U18311 (N_18311,N_18226,N_18057);
xor U18312 (N_18312,N_18127,N_18107);
nor U18313 (N_18313,N_18198,N_18237);
and U18314 (N_18314,N_18033,N_18082);
nand U18315 (N_18315,N_18233,N_18243);
and U18316 (N_18316,N_18050,N_18009);
and U18317 (N_18317,N_18011,N_18161);
and U18318 (N_18318,N_18183,N_18157);
and U18319 (N_18319,N_18111,N_18239);
or U18320 (N_18320,N_18085,N_18000);
or U18321 (N_18321,N_18015,N_18051);
xor U18322 (N_18322,N_18128,N_18144);
or U18323 (N_18323,N_18142,N_18160);
nor U18324 (N_18324,N_18129,N_18189);
xnor U18325 (N_18325,N_18205,N_18181);
nand U18326 (N_18326,N_18154,N_18147);
xnor U18327 (N_18327,N_18108,N_18200);
nor U18328 (N_18328,N_18068,N_18098);
nor U18329 (N_18329,N_18099,N_18096);
xnor U18330 (N_18330,N_18109,N_18008);
nand U18331 (N_18331,N_18219,N_18045);
nand U18332 (N_18332,N_18034,N_18192);
xor U18333 (N_18333,N_18101,N_18188);
and U18334 (N_18334,N_18028,N_18204);
and U18335 (N_18335,N_18117,N_18061);
and U18336 (N_18336,N_18017,N_18224);
nand U18337 (N_18337,N_18159,N_18055);
xnor U18338 (N_18338,N_18041,N_18052);
or U18339 (N_18339,N_18194,N_18209);
xor U18340 (N_18340,N_18062,N_18245);
or U18341 (N_18341,N_18030,N_18016);
and U18342 (N_18342,N_18163,N_18197);
nor U18343 (N_18343,N_18167,N_18195);
and U18344 (N_18344,N_18024,N_18029);
nand U18345 (N_18345,N_18137,N_18140);
xnor U18346 (N_18346,N_18229,N_18178);
xor U18347 (N_18347,N_18247,N_18047);
nor U18348 (N_18348,N_18176,N_18106);
nand U18349 (N_18349,N_18027,N_18136);
xnor U18350 (N_18350,N_18208,N_18046);
nand U18351 (N_18351,N_18019,N_18150);
and U18352 (N_18352,N_18100,N_18084);
and U18353 (N_18353,N_18065,N_18132);
nor U18354 (N_18354,N_18131,N_18081);
or U18355 (N_18355,N_18225,N_18086);
or U18356 (N_18356,N_18228,N_18184);
and U18357 (N_18357,N_18090,N_18095);
and U18358 (N_18358,N_18155,N_18079);
or U18359 (N_18359,N_18235,N_18020);
nor U18360 (N_18360,N_18227,N_18094);
or U18361 (N_18361,N_18241,N_18063);
and U18362 (N_18362,N_18236,N_18201);
or U18363 (N_18363,N_18212,N_18021);
nor U18364 (N_18364,N_18104,N_18166);
nand U18365 (N_18365,N_18059,N_18246);
nor U18366 (N_18366,N_18179,N_18088);
nand U18367 (N_18367,N_18003,N_18169);
nand U18368 (N_18368,N_18206,N_18123);
nor U18369 (N_18369,N_18218,N_18214);
nand U18370 (N_18370,N_18158,N_18032);
and U18371 (N_18371,N_18152,N_18211);
and U18372 (N_18372,N_18171,N_18037);
nor U18373 (N_18373,N_18215,N_18202);
and U18374 (N_18374,N_18232,N_18180);
nand U18375 (N_18375,N_18109,N_18056);
or U18376 (N_18376,N_18078,N_18047);
nor U18377 (N_18377,N_18202,N_18119);
xnor U18378 (N_18378,N_18085,N_18005);
xor U18379 (N_18379,N_18059,N_18229);
or U18380 (N_18380,N_18029,N_18207);
nand U18381 (N_18381,N_18044,N_18061);
nand U18382 (N_18382,N_18170,N_18008);
nor U18383 (N_18383,N_18020,N_18196);
or U18384 (N_18384,N_18127,N_18060);
and U18385 (N_18385,N_18212,N_18081);
xor U18386 (N_18386,N_18152,N_18145);
nor U18387 (N_18387,N_18026,N_18146);
nand U18388 (N_18388,N_18142,N_18111);
or U18389 (N_18389,N_18205,N_18005);
or U18390 (N_18390,N_18178,N_18181);
and U18391 (N_18391,N_18218,N_18025);
or U18392 (N_18392,N_18194,N_18185);
nand U18393 (N_18393,N_18118,N_18237);
nor U18394 (N_18394,N_18019,N_18014);
or U18395 (N_18395,N_18197,N_18220);
or U18396 (N_18396,N_18120,N_18182);
and U18397 (N_18397,N_18015,N_18097);
xnor U18398 (N_18398,N_18222,N_18014);
and U18399 (N_18399,N_18150,N_18243);
xnor U18400 (N_18400,N_18113,N_18052);
and U18401 (N_18401,N_18083,N_18237);
nor U18402 (N_18402,N_18000,N_18132);
nor U18403 (N_18403,N_18221,N_18223);
xor U18404 (N_18404,N_18033,N_18159);
xnor U18405 (N_18405,N_18101,N_18080);
xor U18406 (N_18406,N_18170,N_18167);
or U18407 (N_18407,N_18232,N_18095);
xor U18408 (N_18408,N_18122,N_18201);
or U18409 (N_18409,N_18028,N_18121);
nand U18410 (N_18410,N_18009,N_18054);
nand U18411 (N_18411,N_18185,N_18110);
nor U18412 (N_18412,N_18065,N_18244);
nor U18413 (N_18413,N_18074,N_18239);
nor U18414 (N_18414,N_18091,N_18109);
nand U18415 (N_18415,N_18126,N_18206);
xor U18416 (N_18416,N_18007,N_18061);
and U18417 (N_18417,N_18013,N_18177);
and U18418 (N_18418,N_18154,N_18188);
or U18419 (N_18419,N_18216,N_18235);
and U18420 (N_18420,N_18163,N_18107);
and U18421 (N_18421,N_18038,N_18204);
xor U18422 (N_18422,N_18010,N_18214);
nor U18423 (N_18423,N_18155,N_18132);
nand U18424 (N_18424,N_18006,N_18060);
nand U18425 (N_18425,N_18218,N_18181);
and U18426 (N_18426,N_18245,N_18009);
nand U18427 (N_18427,N_18122,N_18213);
xor U18428 (N_18428,N_18228,N_18011);
and U18429 (N_18429,N_18088,N_18038);
or U18430 (N_18430,N_18052,N_18114);
or U18431 (N_18431,N_18216,N_18033);
nor U18432 (N_18432,N_18224,N_18028);
and U18433 (N_18433,N_18219,N_18200);
nand U18434 (N_18434,N_18152,N_18224);
nand U18435 (N_18435,N_18192,N_18190);
and U18436 (N_18436,N_18128,N_18227);
and U18437 (N_18437,N_18046,N_18012);
nor U18438 (N_18438,N_18168,N_18128);
or U18439 (N_18439,N_18034,N_18086);
and U18440 (N_18440,N_18048,N_18135);
xor U18441 (N_18441,N_18121,N_18122);
and U18442 (N_18442,N_18113,N_18119);
or U18443 (N_18443,N_18113,N_18179);
nor U18444 (N_18444,N_18034,N_18083);
nand U18445 (N_18445,N_18126,N_18123);
and U18446 (N_18446,N_18034,N_18082);
xor U18447 (N_18447,N_18243,N_18174);
or U18448 (N_18448,N_18224,N_18197);
nand U18449 (N_18449,N_18184,N_18216);
nand U18450 (N_18450,N_18172,N_18171);
nor U18451 (N_18451,N_18134,N_18018);
nor U18452 (N_18452,N_18037,N_18140);
and U18453 (N_18453,N_18116,N_18226);
nand U18454 (N_18454,N_18120,N_18059);
xor U18455 (N_18455,N_18059,N_18015);
nor U18456 (N_18456,N_18062,N_18249);
or U18457 (N_18457,N_18053,N_18087);
nand U18458 (N_18458,N_18188,N_18042);
or U18459 (N_18459,N_18036,N_18028);
nor U18460 (N_18460,N_18148,N_18072);
nand U18461 (N_18461,N_18172,N_18182);
nor U18462 (N_18462,N_18166,N_18192);
xnor U18463 (N_18463,N_18163,N_18041);
or U18464 (N_18464,N_18164,N_18037);
xnor U18465 (N_18465,N_18036,N_18074);
and U18466 (N_18466,N_18103,N_18149);
or U18467 (N_18467,N_18189,N_18048);
xor U18468 (N_18468,N_18224,N_18015);
nand U18469 (N_18469,N_18001,N_18054);
nand U18470 (N_18470,N_18044,N_18160);
nor U18471 (N_18471,N_18176,N_18140);
nor U18472 (N_18472,N_18181,N_18223);
nand U18473 (N_18473,N_18094,N_18128);
nor U18474 (N_18474,N_18247,N_18163);
or U18475 (N_18475,N_18220,N_18122);
or U18476 (N_18476,N_18027,N_18115);
nand U18477 (N_18477,N_18113,N_18051);
or U18478 (N_18478,N_18152,N_18066);
or U18479 (N_18479,N_18131,N_18039);
xnor U18480 (N_18480,N_18032,N_18089);
and U18481 (N_18481,N_18198,N_18178);
or U18482 (N_18482,N_18198,N_18076);
xor U18483 (N_18483,N_18242,N_18182);
or U18484 (N_18484,N_18045,N_18234);
and U18485 (N_18485,N_18017,N_18248);
and U18486 (N_18486,N_18212,N_18144);
nand U18487 (N_18487,N_18023,N_18132);
nor U18488 (N_18488,N_18082,N_18011);
and U18489 (N_18489,N_18008,N_18101);
nand U18490 (N_18490,N_18025,N_18020);
or U18491 (N_18491,N_18227,N_18141);
and U18492 (N_18492,N_18007,N_18169);
xnor U18493 (N_18493,N_18218,N_18115);
and U18494 (N_18494,N_18049,N_18198);
xor U18495 (N_18495,N_18062,N_18006);
or U18496 (N_18496,N_18182,N_18112);
xor U18497 (N_18497,N_18240,N_18062);
xor U18498 (N_18498,N_18093,N_18073);
and U18499 (N_18499,N_18034,N_18143);
nor U18500 (N_18500,N_18429,N_18327);
xnor U18501 (N_18501,N_18460,N_18380);
xor U18502 (N_18502,N_18370,N_18495);
and U18503 (N_18503,N_18413,N_18354);
or U18504 (N_18504,N_18387,N_18438);
xnor U18505 (N_18505,N_18353,N_18382);
nand U18506 (N_18506,N_18391,N_18477);
and U18507 (N_18507,N_18449,N_18462);
nor U18508 (N_18508,N_18260,N_18364);
xnor U18509 (N_18509,N_18344,N_18360);
nand U18510 (N_18510,N_18322,N_18346);
xnor U18511 (N_18511,N_18358,N_18420);
or U18512 (N_18512,N_18445,N_18279);
nand U18513 (N_18513,N_18266,N_18384);
xnor U18514 (N_18514,N_18252,N_18458);
xor U18515 (N_18515,N_18342,N_18411);
xnor U18516 (N_18516,N_18268,N_18457);
xnor U18517 (N_18517,N_18287,N_18406);
or U18518 (N_18518,N_18271,N_18465);
nand U18519 (N_18519,N_18483,N_18325);
xnor U18520 (N_18520,N_18434,N_18479);
xnor U18521 (N_18521,N_18398,N_18273);
or U18522 (N_18522,N_18447,N_18464);
and U18523 (N_18523,N_18362,N_18446);
nand U18524 (N_18524,N_18355,N_18454);
nor U18525 (N_18525,N_18472,N_18459);
xor U18526 (N_18526,N_18363,N_18421);
or U18527 (N_18527,N_18390,N_18359);
or U18528 (N_18528,N_18250,N_18461);
xnor U18529 (N_18529,N_18320,N_18395);
xor U18530 (N_18530,N_18361,N_18270);
xnor U18531 (N_18531,N_18432,N_18276);
nand U18532 (N_18532,N_18377,N_18478);
nor U18533 (N_18533,N_18452,N_18265);
xnor U18534 (N_18534,N_18453,N_18290);
nor U18535 (N_18535,N_18385,N_18407);
xor U18536 (N_18536,N_18326,N_18482);
nand U18537 (N_18537,N_18497,N_18475);
xnor U18538 (N_18538,N_18489,N_18401);
and U18539 (N_18539,N_18275,N_18254);
nand U18540 (N_18540,N_18402,N_18451);
nor U18541 (N_18541,N_18394,N_18272);
and U18542 (N_18542,N_18280,N_18357);
and U18543 (N_18543,N_18435,N_18296);
or U18544 (N_18544,N_18282,N_18318);
or U18545 (N_18545,N_18261,N_18339);
nand U18546 (N_18546,N_18373,N_18392);
xnor U18547 (N_18547,N_18412,N_18300);
xor U18548 (N_18548,N_18263,N_18337);
and U18549 (N_18549,N_18253,N_18316);
nand U18550 (N_18550,N_18443,N_18437);
or U18551 (N_18551,N_18468,N_18424);
nor U18552 (N_18552,N_18264,N_18348);
nand U18553 (N_18553,N_18471,N_18259);
xor U18554 (N_18554,N_18397,N_18288);
and U18555 (N_18555,N_18383,N_18433);
or U18556 (N_18556,N_18450,N_18303);
nor U18557 (N_18557,N_18409,N_18470);
xor U18558 (N_18558,N_18305,N_18352);
xnor U18559 (N_18559,N_18474,N_18405);
xnor U18560 (N_18560,N_18444,N_18313);
xnor U18561 (N_18561,N_18334,N_18256);
xor U18562 (N_18562,N_18415,N_18350);
nor U18563 (N_18563,N_18331,N_18369);
nand U18564 (N_18564,N_18374,N_18292);
or U18565 (N_18565,N_18492,N_18410);
nand U18566 (N_18566,N_18277,N_18498);
xor U18567 (N_18567,N_18343,N_18274);
or U18568 (N_18568,N_18289,N_18367);
xor U18569 (N_18569,N_18328,N_18487);
and U18570 (N_18570,N_18351,N_18321);
xor U18571 (N_18571,N_18293,N_18307);
or U18572 (N_18572,N_18340,N_18371);
xor U18573 (N_18573,N_18285,N_18430);
or U18574 (N_18574,N_18414,N_18258);
nor U18575 (N_18575,N_18312,N_18388);
nor U18576 (N_18576,N_18375,N_18330);
nor U18577 (N_18577,N_18349,N_18310);
or U18578 (N_18578,N_18448,N_18267);
nand U18579 (N_18579,N_18368,N_18376);
and U18580 (N_18580,N_18311,N_18319);
xnor U18581 (N_18581,N_18455,N_18416);
xnor U18582 (N_18582,N_18436,N_18393);
nor U18583 (N_18583,N_18297,N_18378);
or U18584 (N_18584,N_18308,N_18335);
nand U18585 (N_18585,N_18333,N_18491);
xor U18586 (N_18586,N_18473,N_18456);
nand U18587 (N_18587,N_18295,N_18299);
nor U18588 (N_18588,N_18255,N_18323);
and U18589 (N_18589,N_18372,N_18431);
xnor U18590 (N_18590,N_18417,N_18314);
nor U18591 (N_18591,N_18347,N_18251);
nor U18592 (N_18592,N_18356,N_18476);
nand U18593 (N_18593,N_18315,N_18493);
xor U18594 (N_18594,N_18400,N_18332);
and U18595 (N_18595,N_18423,N_18317);
or U18596 (N_18596,N_18463,N_18488);
nand U18597 (N_18597,N_18329,N_18338);
xor U18598 (N_18598,N_18403,N_18496);
nand U18599 (N_18599,N_18336,N_18499);
nand U18600 (N_18600,N_18439,N_18426);
and U18601 (N_18601,N_18278,N_18485);
and U18602 (N_18602,N_18427,N_18304);
nor U18603 (N_18603,N_18441,N_18428);
xnor U18604 (N_18604,N_18386,N_18341);
or U18605 (N_18605,N_18365,N_18486);
or U18606 (N_18606,N_18399,N_18418);
or U18607 (N_18607,N_18467,N_18494);
nor U18608 (N_18608,N_18425,N_18269);
xor U18609 (N_18609,N_18469,N_18324);
nor U18610 (N_18610,N_18345,N_18480);
xnor U18611 (N_18611,N_18301,N_18306);
nor U18612 (N_18612,N_18481,N_18408);
or U18613 (N_18613,N_18396,N_18440);
nand U18614 (N_18614,N_18419,N_18466);
xnor U18615 (N_18615,N_18442,N_18262);
and U18616 (N_18616,N_18291,N_18302);
nand U18617 (N_18617,N_18422,N_18379);
and U18618 (N_18618,N_18366,N_18294);
or U18619 (N_18619,N_18284,N_18257);
nand U18620 (N_18620,N_18381,N_18283);
nor U18621 (N_18621,N_18490,N_18309);
and U18622 (N_18622,N_18281,N_18298);
nand U18623 (N_18623,N_18286,N_18404);
and U18624 (N_18624,N_18484,N_18389);
xnor U18625 (N_18625,N_18386,N_18354);
nand U18626 (N_18626,N_18255,N_18260);
and U18627 (N_18627,N_18320,N_18469);
xor U18628 (N_18628,N_18291,N_18354);
nand U18629 (N_18629,N_18317,N_18400);
nor U18630 (N_18630,N_18484,N_18279);
and U18631 (N_18631,N_18395,N_18461);
and U18632 (N_18632,N_18296,N_18404);
xnor U18633 (N_18633,N_18348,N_18344);
nor U18634 (N_18634,N_18395,N_18467);
nand U18635 (N_18635,N_18418,N_18430);
nor U18636 (N_18636,N_18314,N_18433);
nor U18637 (N_18637,N_18306,N_18302);
nor U18638 (N_18638,N_18482,N_18331);
or U18639 (N_18639,N_18297,N_18262);
nand U18640 (N_18640,N_18443,N_18383);
nand U18641 (N_18641,N_18401,N_18279);
nand U18642 (N_18642,N_18495,N_18312);
xor U18643 (N_18643,N_18293,N_18340);
or U18644 (N_18644,N_18438,N_18345);
or U18645 (N_18645,N_18376,N_18319);
and U18646 (N_18646,N_18377,N_18448);
or U18647 (N_18647,N_18389,N_18255);
nor U18648 (N_18648,N_18285,N_18352);
or U18649 (N_18649,N_18482,N_18388);
nand U18650 (N_18650,N_18377,N_18414);
or U18651 (N_18651,N_18330,N_18315);
and U18652 (N_18652,N_18271,N_18356);
or U18653 (N_18653,N_18394,N_18269);
nand U18654 (N_18654,N_18454,N_18337);
nand U18655 (N_18655,N_18441,N_18410);
or U18656 (N_18656,N_18460,N_18348);
and U18657 (N_18657,N_18381,N_18397);
nor U18658 (N_18658,N_18403,N_18489);
xnor U18659 (N_18659,N_18461,N_18279);
nor U18660 (N_18660,N_18350,N_18495);
and U18661 (N_18661,N_18365,N_18415);
xnor U18662 (N_18662,N_18381,N_18302);
xnor U18663 (N_18663,N_18454,N_18272);
nand U18664 (N_18664,N_18321,N_18418);
nand U18665 (N_18665,N_18356,N_18459);
nand U18666 (N_18666,N_18316,N_18460);
nand U18667 (N_18667,N_18263,N_18480);
and U18668 (N_18668,N_18331,N_18253);
nor U18669 (N_18669,N_18273,N_18428);
xnor U18670 (N_18670,N_18335,N_18333);
and U18671 (N_18671,N_18308,N_18419);
and U18672 (N_18672,N_18299,N_18343);
nand U18673 (N_18673,N_18274,N_18300);
nand U18674 (N_18674,N_18289,N_18309);
or U18675 (N_18675,N_18443,N_18491);
nor U18676 (N_18676,N_18496,N_18368);
nand U18677 (N_18677,N_18319,N_18275);
or U18678 (N_18678,N_18449,N_18355);
or U18679 (N_18679,N_18407,N_18326);
nand U18680 (N_18680,N_18281,N_18332);
nand U18681 (N_18681,N_18275,N_18465);
nand U18682 (N_18682,N_18276,N_18352);
nor U18683 (N_18683,N_18321,N_18367);
nand U18684 (N_18684,N_18392,N_18263);
and U18685 (N_18685,N_18374,N_18303);
xor U18686 (N_18686,N_18425,N_18301);
xnor U18687 (N_18687,N_18268,N_18468);
nor U18688 (N_18688,N_18444,N_18269);
or U18689 (N_18689,N_18482,N_18256);
xnor U18690 (N_18690,N_18423,N_18443);
nor U18691 (N_18691,N_18360,N_18399);
nand U18692 (N_18692,N_18499,N_18322);
xnor U18693 (N_18693,N_18367,N_18281);
nand U18694 (N_18694,N_18389,N_18341);
xor U18695 (N_18695,N_18403,N_18406);
xor U18696 (N_18696,N_18353,N_18409);
nor U18697 (N_18697,N_18380,N_18381);
and U18698 (N_18698,N_18484,N_18485);
nand U18699 (N_18699,N_18310,N_18468);
and U18700 (N_18700,N_18428,N_18282);
nor U18701 (N_18701,N_18445,N_18269);
or U18702 (N_18702,N_18378,N_18423);
nor U18703 (N_18703,N_18434,N_18267);
xnor U18704 (N_18704,N_18300,N_18406);
or U18705 (N_18705,N_18441,N_18480);
nor U18706 (N_18706,N_18334,N_18490);
nor U18707 (N_18707,N_18374,N_18288);
or U18708 (N_18708,N_18278,N_18252);
nor U18709 (N_18709,N_18350,N_18484);
and U18710 (N_18710,N_18292,N_18313);
and U18711 (N_18711,N_18250,N_18313);
xnor U18712 (N_18712,N_18262,N_18400);
nand U18713 (N_18713,N_18400,N_18436);
or U18714 (N_18714,N_18402,N_18491);
nand U18715 (N_18715,N_18302,N_18404);
nor U18716 (N_18716,N_18437,N_18458);
and U18717 (N_18717,N_18271,N_18431);
xnor U18718 (N_18718,N_18356,N_18331);
nand U18719 (N_18719,N_18295,N_18289);
and U18720 (N_18720,N_18293,N_18406);
and U18721 (N_18721,N_18423,N_18365);
nor U18722 (N_18722,N_18320,N_18425);
and U18723 (N_18723,N_18324,N_18433);
nand U18724 (N_18724,N_18488,N_18383);
or U18725 (N_18725,N_18263,N_18307);
and U18726 (N_18726,N_18291,N_18482);
nand U18727 (N_18727,N_18395,N_18354);
nor U18728 (N_18728,N_18491,N_18315);
or U18729 (N_18729,N_18498,N_18332);
nor U18730 (N_18730,N_18275,N_18371);
xnor U18731 (N_18731,N_18391,N_18410);
nand U18732 (N_18732,N_18428,N_18408);
and U18733 (N_18733,N_18262,N_18458);
xor U18734 (N_18734,N_18332,N_18434);
or U18735 (N_18735,N_18499,N_18425);
nand U18736 (N_18736,N_18461,N_18314);
or U18737 (N_18737,N_18431,N_18407);
xor U18738 (N_18738,N_18368,N_18323);
or U18739 (N_18739,N_18367,N_18259);
nand U18740 (N_18740,N_18306,N_18470);
xor U18741 (N_18741,N_18372,N_18315);
and U18742 (N_18742,N_18458,N_18366);
or U18743 (N_18743,N_18447,N_18328);
and U18744 (N_18744,N_18262,N_18366);
or U18745 (N_18745,N_18357,N_18298);
xor U18746 (N_18746,N_18445,N_18438);
xor U18747 (N_18747,N_18320,N_18487);
and U18748 (N_18748,N_18436,N_18367);
xor U18749 (N_18749,N_18484,N_18412);
nand U18750 (N_18750,N_18612,N_18544);
nor U18751 (N_18751,N_18668,N_18686);
nand U18752 (N_18752,N_18545,N_18599);
xnor U18753 (N_18753,N_18598,N_18670);
or U18754 (N_18754,N_18549,N_18517);
nand U18755 (N_18755,N_18593,N_18640);
nand U18756 (N_18756,N_18644,N_18655);
nand U18757 (N_18757,N_18678,N_18737);
and U18758 (N_18758,N_18527,N_18660);
nor U18759 (N_18759,N_18533,N_18620);
and U18760 (N_18760,N_18747,N_18725);
xor U18761 (N_18761,N_18665,N_18591);
nand U18762 (N_18762,N_18741,N_18652);
and U18763 (N_18763,N_18687,N_18602);
nand U18764 (N_18764,N_18672,N_18711);
nand U18765 (N_18765,N_18634,N_18525);
and U18766 (N_18766,N_18623,N_18580);
nand U18767 (N_18767,N_18715,N_18691);
nor U18768 (N_18768,N_18651,N_18584);
xor U18769 (N_18769,N_18653,N_18556);
and U18770 (N_18770,N_18571,N_18749);
xor U18771 (N_18771,N_18663,N_18702);
xor U18772 (N_18772,N_18676,N_18698);
nor U18773 (N_18773,N_18743,N_18683);
nand U18774 (N_18774,N_18576,N_18566);
xor U18775 (N_18775,N_18709,N_18721);
or U18776 (N_18776,N_18546,N_18558);
xor U18777 (N_18777,N_18561,N_18699);
xor U18778 (N_18778,N_18536,N_18604);
and U18779 (N_18779,N_18514,N_18723);
or U18780 (N_18780,N_18650,N_18642);
xor U18781 (N_18781,N_18637,N_18564);
or U18782 (N_18782,N_18518,N_18532);
nand U18783 (N_18783,N_18645,N_18673);
nor U18784 (N_18784,N_18712,N_18734);
xnor U18785 (N_18785,N_18624,N_18722);
xnor U18786 (N_18786,N_18688,N_18562);
xnor U18787 (N_18787,N_18675,N_18577);
nand U18788 (N_18788,N_18504,N_18694);
or U18789 (N_18789,N_18745,N_18707);
xnor U18790 (N_18790,N_18628,N_18746);
or U18791 (N_18791,N_18587,N_18735);
nor U18792 (N_18792,N_18523,N_18729);
nand U18793 (N_18793,N_18718,N_18573);
and U18794 (N_18794,N_18727,N_18617);
nand U18795 (N_18795,N_18626,N_18714);
nand U18796 (N_18796,N_18716,N_18575);
xor U18797 (N_18797,N_18710,N_18596);
nor U18798 (N_18798,N_18703,N_18543);
nand U18799 (N_18799,N_18529,N_18554);
xnor U18800 (N_18800,N_18685,N_18541);
or U18801 (N_18801,N_18531,N_18552);
and U18802 (N_18802,N_18616,N_18540);
and U18803 (N_18803,N_18516,N_18693);
nor U18804 (N_18804,N_18553,N_18661);
or U18805 (N_18805,N_18601,N_18635);
nor U18806 (N_18806,N_18681,N_18647);
nor U18807 (N_18807,N_18732,N_18510);
nand U18808 (N_18808,N_18520,N_18501);
nor U18809 (N_18809,N_18701,N_18537);
nor U18810 (N_18810,N_18696,N_18530);
nand U18811 (N_18811,N_18684,N_18618);
nand U18812 (N_18812,N_18667,N_18717);
xnor U18813 (N_18813,N_18720,N_18568);
nor U18814 (N_18814,N_18572,N_18742);
xnor U18815 (N_18815,N_18619,N_18646);
nand U18816 (N_18816,N_18574,N_18567);
nand U18817 (N_18817,N_18595,N_18695);
nor U18818 (N_18818,N_18538,N_18597);
nand U18819 (N_18819,N_18594,N_18609);
nand U18820 (N_18820,N_18654,N_18512);
nand U18821 (N_18821,N_18502,N_18585);
xnor U18822 (N_18822,N_18606,N_18633);
nor U18823 (N_18823,N_18611,N_18590);
nand U18824 (N_18824,N_18682,N_18524);
or U18825 (N_18825,N_18583,N_18656);
nand U18826 (N_18826,N_18542,N_18563);
or U18827 (N_18827,N_18615,N_18690);
xor U18828 (N_18828,N_18600,N_18500);
and U18829 (N_18829,N_18679,N_18521);
or U18830 (N_18830,N_18700,N_18565);
or U18831 (N_18831,N_18713,N_18509);
nand U18832 (N_18832,N_18560,N_18614);
or U18833 (N_18833,N_18570,N_18674);
xnor U18834 (N_18834,N_18551,N_18592);
and U18835 (N_18835,N_18708,N_18515);
or U18836 (N_18836,N_18621,N_18578);
nor U18837 (N_18837,N_18582,N_18528);
nor U18838 (N_18838,N_18726,N_18503);
nand U18839 (N_18839,N_18744,N_18550);
nor U18840 (N_18840,N_18632,N_18511);
xnor U18841 (N_18841,N_18581,N_18719);
nand U18842 (N_18842,N_18522,N_18505);
nand U18843 (N_18843,N_18689,N_18603);
nor U18844 (N_18844,N_18738,N_18677);
and U18845 (N_18845,N_18748,N_18586);
or U18846 (N_18846,N_18724,N_18629);
nor U18847 (N_18847,N_18648,N_18630);
and U18848 (N_18848,N_18569,N_18662);
nand U18849 (N_18849,N_18680,N_18638);
or U18850 (N_18850,N_18526,N_18739);
nor U18851 (N_18851,N_18658,N_18608);
and U18852 (N_18852,N_18607,N_18508);
xnor U18853 (N_18853,N_18547,N_18733);
xnor U18854 (N_18854,N_18555,N_18657);
nand U18855 (N_18855,N_18506,N_18639);
nand U18856 (N_18856,N_18671,N_18631);
nand U18857 (N_18857,N_18605,N_18706);
nand U18858 (N_18858,N_18627,N_18557);
xnor U18859 (N_18859,N_18740,N_18588);
or U18860 (N_18860,N_18513,N_18643);
and U18861 (N_18861,N_18535,N_18636);
nor U18862 (N_18862,N_18704,N_18622);
xor U18863 (N_18863,N_18697,N_18507);
nor U18864 (N_18864,N_18692,N_18625);
nor U18865 (N_18865,N_18731,N_18579);
xor U18866 (N_18866,N_18664,N_18548);
and U18867 (N_18867,N_18613,N_18736);
or U18868 (N_18868,N_18641,N_18669);
and U18869 (N_18869,N_18705,N_18730);
xor U18870 (N_18870,N_18666,N_18589);
or U18871 (N_18871,N_18649,N_18539);
nor U18872 (N_18872,N_18659,N_18534);
xnor U18873 (N_18873,N_18559,N_18519);
and U18874 (N_18874,N_18728,N_18610);
or U18875 (N_18875,N_18528,N_18621);
or U18876 (N_18876,N_18539,N_18631);
xor U18877 (N_18877,N_18719,N_18540);
xnor U18878 (N_18878,N_18664,N_18702);
nand U18879 (N_18879,N_18502,N_18500);
xor U18880 (N_18880,N_18509,N_18697);
xnor U18881 (N_18881,N_18648,N_18667);
xnor U18882 (N_18882,N_18645,N_18716);
and U18883 (N_18883,N_18718,N_18534);
or U18884 (N_18884,N_18568,N_18533);
or U18885 (N_18885,N_18532,N_18587);
xnor U18886 (N_18886,N_18736,N_18666);
nor U18887 (N_18887,N_18629,N_18553);
xnor U18888 (N_18888,N_18620,N_18706);
nor U18889 (N_18889,N_18736,N_18551);
nor U18890 (N_18890,N_18742,N_18597);
nor U18891 (N_18891,N_18558,N_18717);
nor U18892 (N_18892,N_18577,N_18529);
or U18893 (N_18893,N_18548,N_18651);
or U18894 (N_18894,N_18505,N_18617);
and U18895 (N_18895,N_18575,N_18614);
and U18896 (N_18896,N_18554,N_18653);
xnor U18897 (N_18897,N_18561,N_18588);
nor U18898 (N_18898,N_18564,N_18678);
and U18899 (N_18899,N_18710,N_18708);
and U18900 (N_18900,N_18536,N_18586);
and U18901 (N_18901,N_18687,N_18645);
nand U18902 (N_18902,N_18630,N_18691);
and U18903 (N_18903,N_18640,N_18688);
nand U18904 (N_18904,N_18651,N_18526);
or U18905 (N_18905,N_18728,N_18559);
nor U18906 (N_18906,N_18642,N_18617);
or U18907 (N_18907,N_18676,N_18743);
or U18908 (N_18908,N_18566,N_18639);
and U18909 (N_18909,N_18686,N_18501);
or U18910 (N_18910,N_18546,N_18705);
nor U18911 (N_18911,N_18688,N_18676);
and U18912 (N_18912,N_18689,N_18691);
and U18913 (N_18913,N_18682,N_18587);
nand U18914 (N_18914,N_18567,N_18701);
xor U18915 (N_18915,N_18574,N_18634);
and U18916 (N_18916,N_18589,N_18720);
nor U18917 (N_18917,N_18631,N_18541);
nand U18918 (N_18918,N_18519,N_18708);
and U18919 (N_18919,N_18552,N_18530);
and U18920 (N_18920,N_18649,N_18575);
and U18921 (N_18921,N_18742,N_18635);
or U18922 (N_18922,N_18641,N_18501);
nand U18923 (N_18923,N_18568,N_18541);
xor U18924 (N_18924,N_18734,N_18595);
and U18925 (N_18925,N_18621,N_18500);
xnor U18926 (N_18926,N_18581,N_18709);
nor U18927 (N_18927,N_18575,N_18615);
xnor U18928 (N_18928,N_18543,N_18589);
or U18929 (N_18929,N_18549,N_18653);
nand U18930 (N_18930,N_18544,N_18583);
and U18931 (N_18931,N_18661,N_18691);
or U18932 (N_18932,N_18718,N_18702);
nand U18933 (N_18933,N_18551,N_18555);
xnor U18934 (N_18934,N_18542,N_18543);
nand U18935 (N_18935,N_18528,N_18518);
nand U18936 (N_18936,N_18577,N_18605);
nor U18937 (N_18937,N_18670,N_18686);
and U18938 (N_18938,N_18677,N_18564);
nand U18939 (N_18939,N_18699,N_18601);
xnor U18940 (N_18940,N_18743,N_18735);
nor U18941 (N_18941,N_18598,N_18692);
or U18942 (N_18942,N_18619,N_18524);
nand U18943 (N_18943,N_18540,N_18738);
or U18944 (N_18944,N_18543,N_18554);
and U18945 (N_18945,N_18520,N_18644);
nor U18946 (N_18946,N_18687,N_18587);
nor U18947 (N_18947,N_18658,N_18631);
and U18948 (N_18948,N_18625,N_18584);
xor U18949 (N_18949,N_18716,N_18520);
xor U18950 (N_18950,N_18512,N_18694);
xor U18951 (N_18951,N_18607,N_18618);
nor U18952 (N_18952,N_18522,N_18677);
or U18953 (N_18953,N_18693,N_18523);
xor U18954 (N_18954,N_18506,N_18528);
and U18955 (N_18955,N_18633,N_18603);
nor U18956 (N_18956,N_18656,N_18557);
xor U18957 (N_18957,N_18563,N_18685);
or U18958 (N_18958,N_18563,N_18722);
nor U18959 (N_18959,N_18739,N_18624);
and U18960 (N_18960,N_18686,N_18648);
or U18961 (N_18961,N_18591,N_18652);
xor U18962 (N_18962,N_18649,N_18735);
and U18963 (N_18963,N_18528,N_18622);
and U18964 (N_18964,N_18558,N_18665);
and U18965 (N_18965,N_18722,N_18714);
or U18966 (N_18966,N_18707,N_18580);
nand U18967 (N_18967,N_18598,N_18667);
and U18968 (N_18968,N_18739,N_18515);
nand U18969 (N_18969,N_18651,N_18505);
and U18970 (N_18970,N_18724,N_18696);
nor U18971 (N_18971,N_18695,N_18659);
nand U18972 (N_18972,N_18526,N_18555);
xnor U18973 (N_18973,N_18610,N_18532);
xor U18974 (N_18974,N_18636,N_18682);
xor U18975 (N_18975,N_18503,N_18525);
nor U18976 (N_18976,N_18506,N_18567);
xor U18977 (N_18977,N_18526,N_18649);
and U18978 (N_18978,N_18732,N_18749);
xnor U18979 (N_18979,N_18709,N_18556);
xor U18980 (N_18980,N_18747,N_18609);
nor U18981 (N_18981,N_18538,N_18717);
xnor U18982 (N_18982,N_18604,N_18594);
nand U18983 (N_18983,N_18631,N_18666);
or U18984 (N_18984,N_18661,N_18566);
or U18985 (N_18985,N_18656,N_18633);
or U18986 (N_18986,N_18642,N_18568);
xnor U18987 (N_18987,N_18713,N_18543);
nand U18988 (N_18988,N_18567,N_18523);
xor U18989 (N_18989,N_18520,N_18688);
xnor U18990 (N_18990,N_18617,N_18742);
nand U18991 (N_18991,N_18639,N_18585);
nor U18992 (N_18992,N_18635,N_18701);
and U18993 (N_18993,N_18563,N_18648);
xor U18994 (N_18994,N_18595,N_18660);
nor U18995 (N_18995,N_18672,N_18624);
xnor U18996 (N_18996,N_18650,N_18569);
and U18997 (N_18997,N_18708,N_18684);
or U18998 (N_18998,N_18709,N_18516);
xor U18999 (N_18999,N_18621,N_18554);
nand U19000 (N_19000,N_18783,N_18956);
nand U19001 (N_19001,N_18846,N_18830);
xor U19002 (N_19002,N_18942,N_18912);
and U19003 (N_19003,N_18941,N_18754);
xnor U19004 (N_19004,N_18898,N_18977);
nand U19005 (N_19005,N_18927,N_18960);
nor U19006 (N_19006,N_18862,N_18943);
or U19007 (N_19007,N_18961,N_18986);
nand U19008 (N_19008,N_18821,N_18966);
or U19009 (N_19009,N_18968,N_18831);
nand U19010 (N_19010,N_18923,N_18750);
nor U19011 (N_19011,N_18920,N_18985);
xor U19012 (N_19012,N_18905,N_18804);
xnor U19013 (N_19013,N_18870,N_18921);
nor U19014 (N_19014,N_18789,N_18962);
nand U19015 (N_19015,N_18872,N_18899);
xnor U19016 (N_19016,N_18932,N_18842);
nand U19017 (N_19017,N_18991,N_18980);
nor U19018 (N_19018,N_18827,N_18885);
nor U19019 (N_19019,N_18992,N_18918);
nor U19020 (N_19020,N_18857,N_18904);
xor U19021 (N_19021,N_18837,N_18843);
xor U19022 (N_19022,N_18996,N_18816);
nand U19023 (N_19023,N_18798,N_18934);
and U19024 (N_19024,N_18852,N_18903);
nand U19025 (N_19025,N_18790,N_18752);
nor U19026 (N_19026,N_18756,N_18832);
and U19027 (N_19027,N_18867,N_18836);
nand U19028 (N_19028,N_18981,N_18775);
xor U19029 (N_19029,N_18972,N_18999);
nand U19030 (N_19030,N_18791,N_18847);
nor U19031 (N_19031,N_18987,N_18990);
nor U19032 (N_19032,N_18967,N_18848);
or U19033 (N_19033,N_18861,N_18755);
nor U19034 (N_19034,N_18864,N_18771);
and U19035 (N_19035,N_18982,N_18763);
xor U19036 (N_19036,N_18853,N_18926);
or U19037 (N_19037,N_18875,N_18856);
and U19038 (N_19038,N_18955,N_18928);
and U19039 (N_19039,N_18845,N_18974);
xor U19040 (N_19040,N_18841,N_18777);
and U19041 (N_19041,N_18808,N_18768);
or U19042 (N_19042,N_18812,N_18902);
nor U19043 (N_19043,N_18963,N_18892);
nand U19044 (N_19044,N_18801,N_18829);
or U19045 (N_19045,N_18869,N_18976);
or U19046 (N_19046,N_18998,N_18809);
nand U19047 (N_19047,N_18973,N_18901);
nor U19048 (N_19048,N_18951,N_18924);
or U19049 (N_19049,N_18793,N_18938);
nand U19050 (N_19050,N_18880,N_18925);
or U19051 (N_19051,N_18954,N_18844);
nand U19052 (N_19052,N_18946,N_18959);
nor U19053 (N_19053,N_18994,N_18811);
xnor U19054 (N_19054,N_18820,N_18948);
xnor U19055 (N_19055,N_18947,N_18840);
nand U19056 (N_19056,N_18806,N_18807);
or U19057 (N_19057,N_18907,N_18970);
nor U19058 (N_19058,N_18826,N_18817);
or U19059 (N_19059,N_18819,N_18776);
or U19060 (N_19060,N_18860,N_18939);
or U19061 (N_19061,N_18865,N_18868);
xnor U19062 (N_19062,N_18803,N_18854);
nor U19063 (N_19063,N_18858,N_18873);
nand U19064 (N_19064,N_18751,N_18802);
nor U19065 (N_19065,N_18759,N_18879);
nor U19066 (N_19066,N_18773,N_18814);
nand U19067 (N_19067,N_18891,N_18889);
nand U19068 (N_19068,N_18893,N_18784);
nor U19069 (N_19069,N_18876,N_18953);
nor U19070 (N_19070,N_18993,N_18761);
or U19071 (N_19071,N_18952,N_18935);
and U19072 (N_19072,N_18795,N_18930);
xor U19073 (N_19073,N_18805,N_18969);
nor U19074 (N_19074,N_18786,N_18828);
and U19075 (N_19075,N_18871,N_18917);
xor U19076 (N_19076,N_18792,N_18878);
xor U19077 (N_19077,N_18958,N_18919);
xor U19078 (N_19078,N_18762,N_18979);
nand U19079 (N_19079,N_18911,N_18855);
or U19080 (N_19080,N_18913,N_18988);
xnor U19081 (N_19081,N_18813,N_18770);
nand U19082 (N_19082,N_18890,N_18818);
or U19083 (N_19083,N_18944,N_18863);
nand U19084 (N_19084,N_18800,N_18850);
and U19085 (N_19085,N_18883,N_18785);
nor U19086 (N_19086,N_18950,N_18910);
xnor U19087 (N_19087,N_18838,N_18887);
and U19088 (N_19088,N_18797,N_18894);
nand U19089 (N_19089,N_18758,N_18874);
and U19090 (N_19090,N_18866,N_18989);
xnor U19091 (N_19091,N_18881,N_18897);
or U19092 (N_19092,N_18965,N_18971);
nand U19093 (N_19093,N_18774,N_18886);
nand U19094 (N_19094,N_18908,N_18794);
nand U19095 (N_19095,N_18810,N_18900);
nand U19096 (N_19096,N_18915,N_18884);
xor U19097 (N_19097,N_18929,N_18769);
and U19098 (N_19098,N_18834,N_18839);
xnor U19099 (N_19099,N_18787,N_18984);
nand U19100 (N_19100,N_18888,N_18781);
nand U19101 (N_19101,N_18922,N_18906);
xor U19102 (N_19102,N_18916,N_18833);
nor U19103 (N_19103,N_18949,N_18772);
xor U19104 (N_19104,N_18995,N_18765);
xor U19105 (N_19105,N_18799,N_18796);
and U19106 (N_19106,N_18824,N_18766);
and U19107 (N_19107,N_18978,N_18753);
nor U19108 (N_19108,N_18936,N_18764);
nor U19109 (N_19109,N_18945,N_18964);
or U19110 (N_19110,N_18822,N_18851);
nand U19111 (N_19111,N_18760,N_18937);
nand U19112 (N_19112,N_18780,N_18779);
nor U19113 (N_19113,N_18877,N_18859);
or U19114 (N_19114,N_18909,N_18933);
xor U19115 (N_19115,N_18896,N_18757);
xnor U19116 (N_19116,N_18975,N_18957);
nor U19117 (N_19117,N_18778,N_18983);
and U19118 (N_19118,N_18940,N_18882);
or U19119 (N_19119,N_18825,N_18815);
or U19120 (N_19120,N_18788,N_18782);
nand U19121 (N_19121,N_18849,N_18823);
nor U19122 (N_19122,N_18997,N_18767);
nor U19123 (N_19123,N_18931,N_18895);
xor U19124 (N_19124,N_18835,N_18914);
or U19125 (N_19125,N_18976,N_18972);
nor U19126 (N_19126,N_18870,N_18869);
xnor U19127 (N_19127,N_18827,N_18995);
nand U19128 (N_19128,N_18940,N_18759);
xnor U19129 (N_19129,N_18965,N_18880);
nand U19130 (N_19130,N_18939,N_18824);
and U19131 (N_19131,N_18823,N_18755);
or U19132 (N_19132,N_18759,N_18893);
xnor U19133 (N_19133,N_18789,N_18870);
and U19134 (N_19134,N_18917,N_18765);
xor U19135 (N_19135,N_18877,N_18833);
nor U19136 (N_19136,N_18851,N_18854);
nor U19137 (N_19137,N_18780,N_18820);
xor U19138 (N_19138,N_18809,N_18967);
and U19139 (N_19139,N_18962,N_18884);
xor U19140 (N_19140,N_18986,N_18985);
or U19141 (N_19141,N_18819,N_18902);
or U19142 (N_19142,N_18798,N_18813);
nand U19143 (N_19143,N_18811,N_18911);
nor U19144 (N_19144,N_18825,N_18783);
and U19145 (N_19145,N_18916,N_18857);
nor U19146 (N_19146,N_18979,N_18753);
and U19147 (N_19147,N_18935,N_18830);
or U19148 (N_19148,N_18878,N_18873);
xor U19149 (N_19149,N_18847,N_18795);
nand U19150 (N_19150,N_18822,N_18981);
xor U19151 (N_19151,N_18957,N_18932);
and U19152 (N_19152,N_18841,N_18898);
nand U19153 (N_19153,N_18784,N_18955);
and U19154 (N_19154,N_18784,N_18929);
and U19155 (N_19155,N_18917,N_18924);
nand U19156 (N_19156,N_18794,N_18832);
nand U19157 (N_19157,N_18868,N_18792);
and U19158 (N_19158,N_18961,N_18947);
and U19159 (N_19159,N_18829,N_18782);
and U19160 (N_19160,N_18778,N_18935);
nand U19161 (N_19161,N_18880,N_18825);
nand U19162 (N_19162,N_18993,N_18757);
nor U19163 (N_19163,N_18911,N_18777);
or U19164 (N_19164,N_18949,N_18821);
and U19165 (N_19165,N_18965,N_18831);
or U19166 (N_19166,N_18881,N_18791);
nand U19167 (N_19167,N_18782,N_18845);
xnor U19168 (N_19168,N_18943,N_18826);
nand U19169 (N_19169,N_18877,N_18928);
nand U19170 (N_19170,N_18794,N_18921);
nand U19171 (N_19171,N_18758,N_18805);
or U19172 (N_19172,N_18875,N_18766);
and U19173 (N_19173,N_18759,N_18956);
and U19174 (N_19174,N_18818,N_18873);
and U19175 (N_19175,N_18815,N_18778);
and U19176 (N_19176,N_18895,N_18867);
nand U19177 (N_19177,N_18984,N_18890);
and U19178 (N_19178,N_18787,N_18769);
nor U19179 (N_19179,N_18803,N_18789);
nand U19180 (N_19180,N_18884,N_18938);
xor U19181 (N_19181,N_18777,N_18925);
nand U19182 (N_19182,N_18979,N_18871);
or U19183 (N_19183,N_18867,N_18762);
nor U19184 (N_19184,N_18980,N_18854);
and U19185 (N_19185,N_18906,N_18830);
nor U19186 (N_19186,N_18863,N_18809);
nand U19187 (N_19187,N_18998,N_18878);
and U19188 (N_19188,N_18876,N_18942);
or U19189 (N_19189,N_18829,N_18804);
nand U19190 (N_19190,N_18795,N_18798);
and U19191 (N_19191,N_18892,N_18853);
nor U19192 (N_19192,N_18912,N_18866);
nor U19193 (N_19193,N_18937,N_18876);
xnor U19194 (N_19194,N_18857,N_18873);
or U19195 (N_19195,N_18808,N_18754);
nor U19196 (N_19196,N_18968,N_18764);
or U19197 (N_19197,N_18948,N_18862);
nand U19198 (N_19198,N_18881,N_18831);
or U19199 (N_19199,N_18850,N_18965);
or U19200 (N_19200,N_18779,N_18845);
and U19201 (N_19201,N_18966,N_18933);
xor U19202 (N_19202,N_18971,N_18852);
nor U19203 (N_19203,N_18996,N_18931);
and U19204 (N_19204,N_18979,N_18830);
nor U19205 (N_19205,N_18866,N_18793);
nand U19206 (N_19206,N_18761,N_18985);
xnor U19207 (N_19207,N_18778,N_18863);
and U19208 (N_19208,N_18895,N_18932);
or U19209 (N_19209,N_18796,N_18772);
nor U19210 (N_19210,N_18822,N_18845);
nand U19211 (N_19211,N_18969,N_18887);
xnor U19212 (N_19212,N_18994,N_18927);
nor U19213 (N_19213,N_18774,N_18979);
xor U19214 (N_19214,N_18922,N_18965);
and U19215 (N_19215,N_18912,N_18842);
and U19216 (N_19216,N_18801,N_18884);
or U19217 (N_19217,N_18976,N_18833);
nor U19218 (N_19218,N_18821,N_18826);
nand U19219 (N_19219,N_18844,N_18766);
xor U19220 (N_19220,N_18990,N_18845);
nor U19221 (N_19221,N_18965,N_18815);
and U19222 (N_19222,N_18989,N_18920);
or U19223 (N_19223,N_18906,N_18958);
nand U19224 (N_19224,N_18934,N_18828);
or U19225 (N_19225,N_18820,N_18828);
nor U19226 (N_19226,N_18916,N_18820);
and U19227 (N_19227,N_18958,N_18922);
xnor U19228 (N_19228,N_18789,N_18801);
nand U19229 (N_19229,N_18888,N_18915);
or U19230 (N_19230,N_18821,N_18796);
nor U19231 (N_19231,N_18803,N_18837);
nand U19232 (N_19232,N_18958,N_18775);
nor U19233 (N_19233,N_18801,N_18972);
and U19234 (N_19234,N_18960,N_18807);
xnor U19235 (N_19235,N_18776,N_18882);
and U19236 (N_19236,N_18811,N_18998);
nor U19237 (N_19237,N_18836,N_18771);
or U19238 (N_19238,N_18997,N_18934);
xor U19239 (N_19239,N_18818,N_18911);
or U19240 (N_19240,N_18835,N_18962);
nand U19241 (N_19241,N_18788,N_18767);
and U19242 (N_19242,N_18827,N_18799);
xnor U19243 (N_19243,N_18981,N_18887);
nand U19244 (N_19244,N_18983,N_18973);
or U19245 (N_19245,N_18913,N_18959);
nor U19246 (N_19246,N_18895,N_18948);
or U19247 (N_19247,N_18806,N_18846);
xnor U19248 (N_19248,N_18761,N_18798);
xnor U19249 (N_19249,N_18996,N_18770);
xor U19250 (N_19250,N_19044,N_19068);
and U19251 (N_19251,N_19138,N_19054);
nand U19252 (N_19252,N_19158,N_19192);
xor U19253 (N_19253,N_19144,N_19186);
xor U19254 (N_19254,N_19011,N_19195);
xnor U19255 (N_19255,N_19225,N_19052);
or U19256 (N_19256,N_19160,N_19080);
nand U19257 (N_19257,N_19005,N_19117);
or U19258 (N_19258,N_19064,N_19175);
or U19259 (N_19259,N_19094,N_19016);
and U19260 (N_19260,N_19046,N_19084);
nand U19261 (N_19261,N_19010,N_19133);
nand U19262 (N_19262,N_19085,N_19164);
xor U19263 (N_19263,N_19100,N_19071);
or U19264 (N_19264,N_19041,N_19135);
nand U19265 (N_19265,N_19078,N_19157);
xnor U19266 (N_19266,N_19007,N_19063);
nand U19267 (N_19267,N_19112,N_19128);
and U19268 (N_19268,N_19076,N_19228);
and U19269 (N_19269,N_19248,N_19211);
or U19270 (N_19270,N_19176,N_19008);
xnor U19271 (N_19271,N_19139,N_19209);
or U19272 (N_19272,N_19103,N_19220);
xnor U19273 (N_19273,N_19045,N_19024);
and U19274 (N_19274,N_19058,N_19177);
or U19275 (N_19275,N_19077,N_19020);
nand U19276 (N_19276,N_19030,N_19124);
and U19277 (N_19277,N_19118,N_19150);
nor U19278 (N_19278,N_19090,N_19190);
xor U19279 (N_19279,N_19238,N_19185);
nand U19280 (N_19280,N_19126,N_19140);
nor U19281 (N_19281,N_19130,N_19232);
and U19282 (N_19282,N_19056,N_19104);
nor U19283 (N_19283,N_19042,N_19182);
xor U19284 (N_19284,N_19161,N_19121);
nand U19285 (N_19285,N_19106,N_19239);
or U19286 (N_19286,N_19205,N_19166);
nand U19287 (N_19287,N_19247,N_19039);
nand U19288 (N_19288,N_19061,N_19191);
or U19289 (N_19289,N_19137,N_19111);
or U19290 (N_19290,N_19123,N_19196);
xnor U19291 (N_19291,N_19216,N_19234);
nor U19292 (N_19292,N_19129,N_19212);
nor U19293 (N_19293,N_19214,N_19029);
nor U19294 (N_19294,N_19149,N_19241);
and U19295 (N_19295,N_19099,N_19155);
xnor U19296 (N_19296,N_19227,N_19116);
and U19297 (N_19297,N_19219,N_19197);
xor U19298 (N_19298,N_19067,N_19022);
nor U19299 (N_19299,N_19213,N_19057);
nand U19300 (N_19300,N_19110,N_19089);
or U19301 (N_19301,N_19184,N_19249);
and U19302 (N_19302,N_19156,N_19031);
or U19303 (N_19303,N_19229,N_19179);
nand U19304 (N_19304,N_19168,N_19086);
nor U19305 (N_19305,N_19218,N_19170);
nor U19306 (N_19306,N_19147,N_19189);
and U19307 (N_19307,N_19051,N_19180);
nor U19308 (N_19308,N_19003,N_19047);
or U19309 (N_19309,N_19231,N_19204);
and U19310 (N_19310,N_19171,N_19027);
xor U19311 (N_19311,N_19098,N_19079);
or U19312 (N_19312,N_19109,N_19115);
or U19313 (N_19313,N_19036,N_19183);
xnor U19314 (N_19314,N_19097,N_19159);
nor U19315 (N_19315,N_19198,N_19143);
nor U19316 (N_19316,N_19233,N_19049);
and U19317 (N_19317,N_19023,N_19242);
and U19318 (N_19318,N_19122,N_19028);
xor U19319 (N_19319,N_19194,N_19034);
or U19320 (N_19320,N_19217,N_19002);
nand U19321 (N_19321,N_19025,N_19000);
nor U19322 (N_19322,N_19221,N_19038);
and U19323 (N_19323,N_19001,N_19018);
and U19324 (N_19324,N_19141,N_19073);
xnor U19325 (N_19325,N_19173,N_19132);
and U19326 (N_19326,N_19222,N_19093);
or U19327 (N_19327,N_19037,N_19059);
nand U19328 (N_19328,N_19096,N_19230);
or U19329 (N_19329,N_19172,N_19095);
nor U19330 (N_19330,N_19120,N_19055);
nor U19331 (N_19331,N_19245,N_19012);
xnor U19332 (N_19332,N_19082,N_19014);
and U19333 (N_19333,N_19244,N_19060);
or U19334 (N_19334,N_19033,N_19050);
and U19335 (N_19335,N_19091,N_19201);
nor U19336 (N_19336,N_19026,N_19240);
nor U19337 (N_19337,N_19199,N_19134);
or U19338 (N_19338,N_19105,N_19146);
xnor U19339 (N_19339,N_19035,N_19148);
and U19340 (N_19340,N_19017,N_19187);
nor U19341 (N_19341,N_19004,N_19114);
and U19342 (N_19342,N_19165,N_19053);
nor U19343 (N_19343,N_19131,N_19043);
nor U19344 (N_19344,N_19092,N_19178);
and U19345 (N_19345,N_19006,N_19136);
nor U19346 (N_19346,N_19226,N_19167);
or U19347 (N_19347,N_19101,N_19069);
xnor U19348 (N_19348,N_19074,N_19021);
xnor U19349 (N_19349,N_19048,N_19200);
or U19350 (N_19350,N_19107,N_19088);
or U19351 (N_19351,N_19070,N_19040);
and U19352 (N_19352,N_19062,N_19108);
and U19353 (N_19353,N_19174,N_19206);
nand U19354 (N_19354,N_19127,N_19202);
nor U19355 (N_19355,N_19235,N_19208);
nand U19356 (N_19356,N_19125,N_19066);
nor U19357 (N_19357,N_19203,N_19032);
and U19358 (N_19358,N_19087,N_19075);
nor U19359 (N_19359,N_19102,N_19224);
and U19360 (N_19360,N_19210,N_19215);
and U19361 (N_19361,N_19162,N_19019);
or U19362 (N_19362,N_19207,N_19223);
xnor U19363 (N_19363,N_19169,N_19145);
xnor U19364 (N_19364,N_19009,N_19236);
and U19365 (N_19365,N_19243,N_19151);
and U19366 (N_19366,N_19154,N_19193);
or U19367 (N_19367,N_19083,N_19013);
nor U19368 (N_19368,N_19246,N_19142);
xor U19369 (N_19369,N_19152,N_19237);
or U19370 (N_19370,N_19072,N_19015);
nand U19371 (N_19371,N_19119,N_19163);
nand U19372 (N_19372,N_19113,N_19181);
nand U19373 (N_19373,N_19188,N_19065);
or U19374 (N_19374,N_19153,N_19081);
nor U19375 (N_19375,N_19143,N_19189);
and U19376 (N_19376,N_19006,N_19097);
xor U19377 (N_19377,N_19228,N_19024);
or U19378 (N_19378,N_19106,N_19237);
xnor U19379 (N_19379,N_19231,N_19064);
nor U19380 (N_19380,N_19029,N_19159);
and U19381 (N_19381,N_19029,N_19103);
nand U19382 (N_19382,N_19120,N_19017);
or U19383 (N_19383,N_19100,N_19153);
or U19384 (N_19384,N_19058,N_19140);
or U19385 (N_19385,N_19025,N_19177);
nand U19386 (N_19386,N_19216,N_19198);
and U19387 (N_19387,N_19228,N_19117);
xnor U19388 (N_19388,N_19126,N_19237);
and U19389 (N_19389,N_19025,N_19056);
xor U19390 (N_19390,N_19103,N_19248);
nor U19391 (N_19391,N_19121,N_19221);
xnor U19392 (N_19392,N_19198,N_19180);
nor U19393 (N_19393,N_19115,N_19199);
xor U19394 (N_19394,N_19143,N_19124);
xnor U19395 (N_19395,N_19129,N_19111);
nand U19396 (N_19396,N_19180,N_19015);
or U19397 (N_19397,N_19006,N_19003);
and U19398 (N_19398,N_19020,N_19181);
xnor U19399 (N_19399,N_19032,N_19043);
or U19400 (N_19400,N_19241,N_19109);
nor U19401 (N_19401,N_19067,N_19208);
nor U19402 (N_19402,N_19166,N_19069);
and U19403 (N_19403,N_19120,N_19127);
nor U19404 (N_19404,N_19156,N_19210);
nand U19405 (N_19405,N_19045,N_19035);
nand U19406 (N_19406,N_19202,N_19057);
xnor U19407 (N_19407,N_19029,N_19213);
xor U19408 (N_19408,N_19095,N_19075);
and U19409 (N_19409,N_19085,N_19175);
nand U19410 (N_19410,N_19176,N_19147);
nand U19411 (N_19411,N_19118,N_19131);
or U19412 (N_19412,N_19088,N_19181);
nand U19413 (N_19413,N_19152,N_19001);
nand U19414 (N_19414,N_19110,N_19202);
or U19415 (N_19415,N_19186,N_19075);
or U19416 (N_19416,N_19041,N_19242);
or U19417 (N_19417,N_19015,N_19039);
nand U19418 (N_19418,N_19225,N_19135);
nor U19419 (N_19419,N_19199,N_19021);
nor U19420 (N_19420,N_19188,N_19227);
or U19421 (N_19421,N_19112,N_19037);
and U19422 (N_19422,N_19206,N_19178);
and U19423 (N_19423,N_19186,N_19057);
xor U19424 (N_19424,N_19203,N_19149);
or U19425 (N_19425,N_19017,N_19157);
or U19426 (N_19426,N_19112,N_19125);
nand U19427 (N_19427,N_19111,N_19079);
nand U19428 (N_19428,N_19211,N_19203);
nand U19429 (N_19429,N_19074,N_19142);
and U19430 (N_19430,N_19074,N_19102);
nand U19431 (N_19431,N_19101,N_19091);
or U19432 (N_19432,N_19172,N_19022);
nor U19433 (N_19433,N_19077,N_19225);
xor U19434 (N_19434,N_19103,N_19013);
nand U19435 (N_19435,N_19205,N_19239);
or U19436 (N_19436,N_19054,N_19034);
xnor U19437 (N_19437,N_19153,N_19071);
and U19438 (N_19438,N_19128,N_19119);
nor U19439 (N_19439,N_19064,N_19016);
or U19440 (N_19440,N_19162,N_19098);
or U19441 (N_19441,N_19122,N_19023);
or U19442 (N_19442,N_19175,N_19105);
nor U19443 (N_19443,N_19111,N_19086);
xnor U19444 (N_19444,N_19100,N_19168);
and U19445 (N_19445,N_19196,N_19022);
and U19446 (N_19446,N_19008,N_19044);
and U19447 (N_19447,N_19201,N_19051);
nor U19448 (N_19448,N_19197,N_19118);
xor U19449 (N_19449,N_19154,N_19072);
and U19450 (N_19450,N_19138,N_19058);
nand U19451 (N_19451,N_19158,N_19156);
nand U19452 (N_19452,N_19013,N_19213);
xor U19453 (N_19453,N_19131,N_19117);
or U19454 (N_19454,N_19090,N_19026);
or U19455 (N_19455,N_19230,N_19244);
nor U19456 (N_19456,N_19004,N_19209);
nor U19457 (N_19457,N_19172,N_19209);
nand U19458 (N_19458,N_19142,N_19034);
or U19459 (N_19459,N_19199,N_19096);
or U19460 (N_19460,N_19108,N_19198);
nor U19461 (N_19461,N_19182,N_19065);
xor U19462 (N_19462,N_19117,N_19068);
nor U19463 (N_19463,N_19209,N_19237);
xor U19464 (N_19464,N_19221,N_19089);
or U19465 (N_19465,N_19156,N_19170);
nor U19466 (N_19466,N_19130,N_19025);
nor U19467 (N_19467,N_19115,N_19227);
nor U19468 (N_19468,N_19019,N_19018);
and U19469 (N_19469,N_19197,N_19164);
or U19470 (N_19470,N_19172,N_19079);
nand U19471 (N_19471,N_19082,N_19211);
and U19472 (N_19472,N_19223,N_19168);
xor U19473 (N_19473,N_19154,N_19118);
nand U19474 (N_19474,N_19001,N_19167);
nand U19475 (N_19475,N_19046,N_19137);
xnor U19476 (N_19476,N_19210,N_19214);
nor U19477 (N_19477,N_19098,N_19120);
nor U19478 (N_19478,N_19119,N_19240);
and U19479 (N_19479,N_19232,N_19108);
or U19480 (N_19480,N_19054,N_19083);
nor U19481 (N_19481,N_19132,N_19061);
nor U19482 (N_19482,N_19017,N_19006);
nor U19483 (N_19483,N_19109,N_19173);
nor U19484 (N_19484,N_19147,N_19006);
and U19485 (N_19485,N_19162,N_19023);
and U19486 (N_19486,N_19040,N_19140);
xnor U19487 (N_19487,N_19068,N_19217);
or U19488 (N_19488,N_19151,N_19234);
xor U19489 (N_19489,N_19151,N_19199);
nor U19490 (N_19490,N_19070,N_19156);
or U19491 (N_19491,N_19141,N_19128);
xnor U19492 (N_19492,N_19075,N_19243);
nor U19493 (N_19493,N_19168,N_19102);
xor U19494 (N_19494,N_19016,N_19240);
xnor U19495 (N_19495,N_19041,N_19180);
nand U19496 (N_19496,N_19130,N_19083);
or U19497 (N_19497,N_19245,N_19015);
xnor U19498 (N_19498,N_19180,N_19162);
nand U19499 (N_19499,N_19108,N_19003);
or U19500 (N_19500,N_19380,N_19404);
or U19501 (N_19501,N_19323,N_19407);
nor U19502 (N_19502,N_19257,N_19261);
or U19503 (N_19503,N_19405,N_19263);
and U19504 (N_19504,N_19436,N_19253);
and U19505 (N_19505,N_19367,N_19256);
or U19506 (N_19506,N_19417,N_19304);
nand U19507 (N_19507,N_19258,N_19430);
and U19508 (N_19508,N_19276,N_19411);
nand U19509 (N_19509,N_19271,N_19314);
nand U19510 (N_19510,N_19463,N_19279);
nand U19511 (N_19511,N_19477,N_19451);
nor U19512 (N_19512,N_19447,N_19471);
nor U19513 (N_19513,N_19265,N_19427);
nand U19514 (N_19514,N_19291,N_19371);
nand U19515 (N_19515,N_19292,N_19457);
xor U19516 (N_19516,N_19472,N_19348);
and U19517 (N_19517,N_19446,N_19342);
nand U19518 (N_19518,N_19432,N_19487);
nand U19519 (N_19519,N_19412,N_19382);
nand U19520 (N_19520,N_19293,N_19459);
and U19521 (N_19521,N_19486,N_19288);
xor U19522 (N_19522,N_19384,N_19460);
nor U19523 (N_19523,N_19422,N_19426);
nand U19524 (N_19524,N_19324,N_19482);
and U19525 (N_19525,N_19289,N_19421);
nor U19526 (N_19526,N_19343,N_19303);
nand U19527 (N_19527,N_19435,N_19360);
xor U19528 (N_19528,N_19373,N_19464);
nand U19529 (N_19529,N_19250,N_19310);
and U19530 (N_19530,N_19498,N_19285);
and U19531 (N_19531,N_19350,N_19390);
nand U19532 (N_19532,N_19375,N_19282);
xor U19533 (N_19533,N_19272,N_19496);
or U19534 (N_19534,N_19307,N_19366);
or U19535 (N_19535,N_19368,N_19488);
nor U19536 (N_19536,N_19281,N_19409);
and U19537 (N_19537,N_19251,N_19474);
or U19538 (N_19538,N_19420,N_19441);
nor U19539 (N_19539,N_19347,N_19468);
and U19540 (N_19540,N_19490,N_19315);
nor U19541 (N_19541,N_19294,N_19492);
or U19542 (N_19542,N_19356,N_19335);
xnor U19543 (N_19543,N_19444,N_19392);
nor U19544 (N_19544,N_19345,N_19332);
nand U19545 (N_19545,N_19453,N_19277);
nor U19546 (N_19546,N_19393,N_19341);
and U19547 (N_19547,N_19408,N_19445);
nor U19548 (N_19548,N_19467,N_19349);
nor U19549 (N_19549,N_19454,N_19317);
and U19550 (N_19550,N_19416,N_19280);
and U19551 (N_19551,N_19318,N_19287);
xnor U19552 (N_19552,N_19458,N_19481);
nand U19553 (N_19553,N_19494,N_19376);
xnor U19554 (N_19554,N_19329,N_19419);
xor U19555 (N_19555,N_19300,N_19320);
nand U19556 (N_19556,N_19312,N_19327);
nand U19557 (N_19557,N_19322,N_19346);
nand U19558 (N_19558,N_19295,N_19297);
xnor U19559 (N_19559,N_19495,N_19406);
and U19560 (N_19560,N_19316,N_19385);
and U19561 (N_19561,N_19440,N_19484);
nand U19562 (N_19562,N_19378,N_19479);
and U19563 (N_19563,N_19357,N_19308);
and U19564 (N_19564,N_19338,N_19399);
and U19565 (N_19565,N_19273,N_19344);
or U19566 (N_19566,N_19377,N_19267);
nor U19567 (N_19567,N_19355,N_19489);
xnor U19568 (N_19568,N_19443,N_19321);
nor U19569 (N_19569,N_19354,N_19306);
nor U19570 (N_19570,N_19359,N_19290);
xnor U19571 (N_19571,N_19470,N_19434);
nand U19572 (N_19572,N_19313,N_19264);
nand U19573 (N_19573,N_19372,N_19428);
nor U19574 (N_19574,N_19431,N_19352);
or U19575 (N_19575,N_19491,N_19395);
nand U19576 (N_19576,N_19284,N_19480);
xor U19577 (N_19577,N_19450,N_19437);
nand U19578 (N_19578,N_19418,N_19483);
nor U19579 (N_19579,N_19469,N_19333);
nand U19580 (N_19580,N_19305,N_19363);
nand U19581 (N_19581,N_19499,N_19286);
and U19582 (N_19582,N_19330,N_19462);
and U19583 (N_19583,N_19353,N_19334);
nand U19584 (N_19584,N_19401,N_19403);
xnor U19585 (N_19585,N_19336,N_19274);
or U19586 (N_19586,N_19298,N_19325);
xnor U19587 (N_19587,N_19328,N_19364);
or U19588 (N_19588,N_19299,N_19255);
nor U19589 (N_19589,N_19337,N_19398);
or U19590 (N_19590,N_19370,N_19268);
and U19591 (N_19591,N_19381,N_19461);
or U19592 (N_19592,N_19433,N_19358);
nor U19593 (N_19593,N_19389,N_19394);
nor U19594 (N_19594,N_19497,N_19275);
nor U19595 (N_19595,N_19478,N_19388);
nand U19596 (N_19596,N_19402,N_19423);
xor U19597 (N_19597,N_19476,N_19270);
or U19598 (N_19598,N_19319,N_19456);
nor U19599 (N_19599,N_19449,N_19302);
or U19600 (N_19600,N_19448,N_19379);
nor U19601 (N_19601,N_19311,N_19340);
and U19602 (N_19602,N_19391,N_19413);
and U19603 (N_19603,N_19259,N_19485);
or U19604 (N_19604,N_19465,N_19262);
nand U19605 (N_19605,N_19365,N_19455);
or U19606 (N_19606,N_19309,N_19301);
or U19607 (N_19607,N_19400,N_19414);
nor U19608 (N_19608,N_19266,N_19475);
nand U19609 (N_19609,N_19415,N_19374);
or U19610 (N_19610,N_19493,N_19425);
nor U19611 (N_19611,N_19396,N_19439);
nand U19612 (N_19612,N_19397,N_19369);
nand U19613 (N_19613,N_19283,N_19383);
and U19614 (N_19614,N_19326,N_19442);
or U19615 (N_19615,N_19452,N_19339);
nand U19616 (N_19616,N_19410,N_19438);
and U19617 (N_19617,N_19331,N_19424);
xor U19618 (N_19618,N_19351,N_19473);
nand U19619 (N_19619,N_19387,N_19362);
xor U19620 (N_19620,N_19260,N_19252);
nand U19621 (N_19621,N_19278,N_19296);
nand U19622 (N_19622,N_19429,N_19386);
and U19623 (N_19623,N_19466,N_19254);
or U19624 (N_19624,N_19361,N_19269);
nor U19625 (N_19625,N_19303,N_19289);
and U19626 (N_19626,N_19291,N_19391);
xnor U19627 (N_19627,N_19349,N_19298);
nand U19628 (N_19628,N_19341,N_19279);
or U19629 (N_19629,N_19456,N_19421);
xor U19630 (N_19630,N_19321,N_19381);
and U19631 (N_19631,N_19417,N_19448);
nand U19632 (N_19632,N_19396,N_19358);
nand U19633 (N_19633,N_19496,N_19347);
nor U19634 (N_19634,N_19426,N_19380);
or U19635 (N_19635,N_19489,N_19462);
and U19636 (N_19636,N_19294,N_19288);
xor U19637 (N_19637,N_19315,N_19354);
and U19638 (N_19638,N_19463,N_19406);
xnor U19639 (N_19639,N_19342,N_19275);
nor U19640 (N_19640,N_19339,N_19459);
xor U19641 (N_19641,N_19422,N_19399);
and U19642 (N_19642,N_19460,N_19372);
nor U19643 (N_19643,N_19308,N_19437);
or U19644 (N_19644,N_19400,N_19342);
nor U19645 (N_19645,N_19330,N_19312);
or U19646 (N_19646,N_19372,N_19303);
and U19647 (N_19647,N_19293,N_19382);
xnor U19648 (N_19648,N_19310,N_19385);
and U19649 (N_19649,N_19322,N_19360);
xor U19650 (N_19650,N_19308,N_19360);
xnor U19651 (N_19651,N_19478,N_19321);
or U19652 (N_19652,N_19265,N_19317);
or U19653 (N_19653,N_19494,N_19413);
nand U19654 (N_19654,N_19341,N_19371);
nor U19655 (N_19655,N_19477,N_19292);
nand U19656 (N_19656,N_19365,N_19463);
xor U19657 (N_19657,N_19402,N_19452);
xor U19658 (N_19658,N_19410,N_19492);
nand U19659 (N_19659,N_19338,N_19361);
or U19660 (N_19660,N_19498,N_19302);
nor U19661 (N_19661,N_19298,N_19281);
nand U19662 (N_19662,N_19292,N_19466);
and U19663 (N_19663,N_19308,N_19320);
xor U19664 (N_19664,N_19289,N_19399);
xor U19665 (N_19665,N_19424,N_19260);
and U19666 (N_19666,N_19274,N_19330);
nor U19667 (N_19667,N_19325,N_19429);
xnor U19668 (N_19668,N_19366,N_19357);
and U19669 (N_19669,N_19346,N_19436);
nor U19670 (N_19670,N_19418,N_19348);
or U19671 (N_19671,N_19424,N_19346);
or U19672 (N_19672,N_19329,N_19333);
or U19673 (N_19673,N_19450,N_19448);
nor U19674 (N_19674,N_19349,N_19326);
or U19675 (N_19675,N_19330,N_19445);
xor U19676 (N_19676,N_19356,N_19470);
and U19677 (N_19677,N_19309,N_19467);
and U19678 (N_19678,N_19349,N_19300);
xnor U19679 (N_19679,N_19276,N_19334);
nor U19680 (N_19680,N_19432,N_19488);
and U19681 (N_19681,N_19260,N_19453);
and U19682 (N_19682,N_19465,N_19283);
nor U19683 (N_19683,N_19271,N_19442);
or U19684 (N_19684,N_19324,N_19290);
xnor U19685 (N_19685,N_19337,N_19431);
and U19686 (N_19686,N_19402,N_19381);
nor U19687 (N_19687,N_19442,N_19373);
or U19688 (N_19688,N_19380,N_19436);
nand U19689 (N_19689,N_19437,N_19285);
nor U19690 (N_19690,N_19461,N_19437);
and U19691 (N_19691,N_19457,N_19338);
nor U19692 (N_19692,N_19443,N_19383);
xnor U19693 (N_19693,N_19476,N_19289);
and U19694 (N_19694,N_19297,N_19318);
or U19695 (N_19695,N_19280,N_19289);
nand U19696 (N_19696,N_19447,N_19430);
xor U19697 (N_19697,N_19465,N_19399);
nor U19698 (N_19698,N_19415,N_19286);
nand U19699 (N_19699,N_19497,N_19288);
or U19700 (N_19700,N_19392,N_19441);
or U19701 (N_19701,N_19422,N_19429);
or U19702 (N_19702,N_19354,N_19438);
nand U19703 (N_19703,N_19263,N_19443);
xor U19704 (N_19704,N_19448,N_19474);
nor U19705 (N_19705,N_19363,N_19496);
xor U19706 (N_19706,N_19388,N_19270);
nand U19707 (N_19707,N_19287,N_19400);
xor U19708 (N_19708,N_19421,N_19358);
xor U19709 (N_19709,N_19398,N_19434);
or U19710 (N_19710,N_19394,N_19478);
nor U19711 (N_19711,N_19425,N_19254);
or U19712 (N_19712,N_19492,N_19338);
xnor U19713 (N_19713,N_19470,N_19448);
nand U19714 (N_19714,N_19394,N_19311);
or U19715 (N_19715,N_19283,N_19391);
nand U19716 (N_19716,N_19323,N_19301);
nor U19717 (N_19717,N_19264,N_19411);
nand U19718 (N_19718,N_19298,N_19312);
nor U19719 (N_19719,N_19408,N_19256);
xor U19720 (N_19720,N_19457,N_19467);
nand U19721 (N_19721,N_19381,N_19266);
xnor U19722 (N_19722,N_19476,N_19461);
nor U19723 (N_19723,N_19270,N_19457);
nand U19724 (N_19724,N_19334,N_19452);
and U19725 (N_19725,N_19456,N_19271);
and U19726 (N_19726,N_19302,N_19304);
nor U19727 (N_19727,N_19496,N_19418);
nand U19728 (N_19728,N_19268,N_19419);
and U19729 (N_19729,N_19262,N_19368);
or U19730 (N_19730,N_19462,N_19404);
nand U19731 (N_19731,N_19354,N_19381);
and U19732 (N_19732,N_19470,N_19472);
and U19733 (N_19733,N_19334,N_19364);
and U19734 (N_19734,N_19447,N_19296);
nor U19735 (N_19735,N_19344,N_19281);
xor U19736 (N_19736,N_19471,N_19262);
nor U19737 (N_19737,N_19492,N_19279);
nand U19738 (N_19738,N_19338,N_19351);
nand U19739 (N_19739,N_19373,N_19310);
and U19740 (N_19740,N_19385,N_19322);
and U19741 (N_19741,N_19460,N_19436);
or U19742 (N_19742,N_19291,N_19450);
xnor U19743 (N_19743,N_19369,N_19336);
xor U19744 (N_19744,N_19414,N_19302);
nand U19745 (N_19745,N_19273,N_19480);
or U19746 (N_19746,N_19407,N_19431);
xor U19747 (N_19747,N_19348,N_19343);
and U19748 (N_19748,N_19336,N_19468);
nand U19749 (N_19749,N_19296,N_19449);
and U19750 (N_19750,N_19727,N_19528);
or U19751 (N_19751,N_19610,N_19672);
or U19752 (N_19752,N_19635,N_19578);
nor U19753 (N_19753,N_19518,N_19552);
nor U19754 (N_19754,N_19686,N_19576);
nor U19755 (N_19755,N_19730,N_19540);
and U19756 (N_19756,N_19705,N_19745);
or U19757 (N_19757,N_19563,N_19668);
or U19758 (N_19758,N_19514,N_19695);
nand U19759 (N_19759,N_19507,N_19503);
and U19760 (N_19760,N_19729,N_19621);
or U19761 (N_19761,N_19604,N_19502);
nor U19762 (N_19762,N_19532,N_19505);
nor U19763 (N_19763,N_19626,N_19746);
nand U19764 (N_19764,N_19506,N_19742);
or U19765 (N_19765,N_19543,N_19559);
and U19766 (N_19766,N_19657,N_19703);
and U19767 (N_19767,N_19740,N_19533);
nand U19768 (N_19768,N_19513,N_19651);
nand U19769 (N_19769,N_19662,N_19679);
nor U19770 (N_19770,N_19581,N_19556);
or U19771 (N_19771,N_19691,N_19720);
or U19772 (N_19772,N_19713,N_19515);
nor U19773 (N_19773,N_19516,N_19504);
nor U19774 (N_19774,N_19710,N_19625);
xnor U19775 (N_19775,N_19530,N_19572);
nand U19776 (N_19776,N_19707,N_19600);
and U19777 (N_19777,N_19612,N_19525);
xnor U19778 (N_19778,N_19709,N_19586);
nor U19779 (N_19779,N_19592,N_19582);
nor U19780 (N_19780,N_19573,N_19526);
nor U19781 (N_19781,N_19511,N_19589);
nand U19782 (N_19782,N_19676,N_19723);
and U19783 (N_19783,N_19697,N_19584);
nor U19784 (N_19784,N_19623,N_19569);
and U19785 (N_19785,N_19544,N_19732);
xnor U19786 (N_19786,N_19636,N_19591);
nand U19787 (N_19787,N_19598,N_19673);
or U19788 (N_19788,N_19666,N_19579);
or U19789 (N_19789,N_19701,N_19501);
and U19790 (N_19790,N_19646,N_19699);
or U19791 (N_19791,N_19541,N_19510);
and U19792 (N_19792,N_19637,N_19690);
nor U19793 (N_19793,N_19698,N_19549);
xor U19794 (N_19794,N_19570,N_19523);
or U19795 (N_19795,N_19733,N_19601);
nor U19796 (N_19796,N_19665,N_19674);
nand U19797 (N_19797,N_19588,N_19692);
nor U19798 (N_19798,N_19638,N_19749);
or U19799 (N_19799,N_19574,N_19652);
nand U19800 (N_19800,N_19554,N_19538);
or U19801 (N_19801,N_19630,N_19603);
or U19802 (N_19802,N_19688,N_19519);
and U19803 (N_19803,N_19696,N_19647);
nand U19804 (N_19804,N_19527,N_19550);
or U19805 (N_19805,N_19583,N_19640);
nand U19806 (N_19806,N_19689,N_19685);
xor U19807 (N_19807,N_19539,N_19711);
nor U19808 (N_19808,N_19509,N_19741);
or U19809 (N_19809,N_19680,N_19599);
or U19810 (N_19810,N_19634,N_19561);
and U19811 (N_19811,N_19667,N_19619);
and U19812 (N_19812,N_19517,N_19675);
and U19813 (N_19813,N_19567,N_19737);
or U19814 (N_19814,N_19564,N_19747);
or U19815 (N_19815,N_19687,N_19616);
or U19816 (N_19816,N_19655,N_19520);
or U19817 (N_19817,N_19717,N_19571);
xor U19818 (N_19818,N_19725,N_19605);
nand U19819 (N_19819,N_19560,N_19587);
or U19820 (N_19820,N_19620,N_19629);
and U19821 (N_19821,N_19649,N_19738);
xor U19822 (N_19822,N_19639,N_19508);
nor U19823 (N_19823,N_19669,N_19531);
nand U19824 (N_19824,N_19658,N_19670);
xnor U19825 (N_19825,N_19683,N_19693);
nand U19826 (N_19826,N_19708,N_19565);
nand U19827 (N_19827,N_19736,N_19536);
nand U19828 (N_19828,N_19615,N_19580);
and U19829 (N_19829,N_19546,N_19521);
and U19830 (N_19830,N_19716,N_19622);
nand U19831 (N_19831,N_19664,N_19631);
or U19832 (N_19832,N_19555,N_19643);
or U19833 (N_19833,N_19654,N_19656);
or U19834 (N_19834,N_19553,N_19577);
nor U19835 (N_19835,N_19661,N_19744);
or U19836 (N_19836,N_19714,N_19597);
and U19837 (N_19837,N_19735,N_19595);
and U19838 (N_19838,N_19704,N_19681);
nand U19839 (N_19839,N_19648,N_19608);
and U19840 (N_19840,N_19684,N_19613);
and U19841 (N_19841,N_19548,N_19534);
nand U19842 (N_19842,N_19522,N_19568);
nand U19843 (N_19843,N_19551,N_19535);
nand U19844 (N_19844,N_19734,N_19653);
and U19845 (N_19845,N_19739,N_19712);
nor U19846 (N_19846,N_19719,N_19500);
nand U19847 (N_19847,N_19529,N_19726);
xnor U19848 (N_19848,N_19617,N_19682);
xnor U19849 (N_19849,N_19537,N_19724);
nor U19850 (N_19850,N_19585,N_19602);
nor U19851 (N_19851,N_19557,N_19642);
nor U19852 (N_19852,N_19545,N_19694);
or U19853 (N_19853,N_19558,N_19644);
nor U19854 (N_19854,N_19728,N_19542);
and U19855 (N_19855,N_19677,N_19650);
nand U19856 (N_19856,N_19628,N_19645);
or U19857 (N_19857,N_19659,N_19607);
and U19858 (N_19858,N_19715,N_19512);
or U19859 (N_19859,N_19731,N_19660);
or U19860 (N_19860,N_19702,N_19614);
and U19861 (N_19861,N_19641,N_19671);
nand U19862 (N_19862,N_19606,N_19632);
and U19863 (N_19863,N_19748,N_19627);
nor U19864 (N_19864,N_19524,N_19678);
xnor U19865 (N_19865,N_19611,N_19593);
nand U19866 (N_19866,N_19743,N_19596);
nand U19867 (N_19867,N_19663,N_19718);
and U19868 (N_19868,N_19594,N_19722);
nor U19869 (N_19869,N_19618,N_19575);
nor U19870 (N_19870,N_19633,N_19566);
nand U19871 (N_19871,N_19562,N_19721);
and U19872 (N_19872,N_19624,N_19547);
and U19873 (N_19873,N_19700,N_19590);
or U19874 (N_19874,N_19609,N_19706);
and U19875 (N_19875,N_19516,N_19560);
nor U19876 (N_19876,N_19732,N_19690);
nand U19877 (N_19877,N_19717,N_19622);
nand U19878 (N_19878,N_19710,N_19680);
and U19879 (N_19879,N_19594,N_19638);
and U19880 (N_19880,N_19516,N_19682);
nand U19881 (N_19881,N_19571,N_19733);
and U19882 (N_19882,N_19636,N_19616);
nor U19883 (N_19883,N_19581,N_19742);
and U19884 (N_19884,N_19580,N_19722);
or U19885 (N_19885,N_19725,N_19658);
and U19886 (N_19886,N_19662,N_19623);
nor U19887 (N_19887,N_19748,N_19519);
xnor U19888 (N_19888,N_19732,N_19567);
xor U19889 (N_19889,N_19603,N_19505);
xnor U19890 (N_19890,N_19718,N_19662);
nor U19891 (N_19891,N_19722,N_19506);
or U19892 (N_19892,N_19520,N_19584);
nand U19893 (N_19893,N_19552,N_19516);
and U19894 (N_19894,N_19603,N_19531);
nor U19895 (N_19895,N_19676,N_19637);
nor U19896 (N_19896,N_19748,N_19635);
or U19897 (N_19897,N_19542,N_19696);
nand U19898 (N_19898,N_19626,N_19657);
nand U19899 (N_19899,N_19631,N_19646);
nor U19900 (N_19900,N_19654,N_19606);
or U19901 (N_19901,N_19630,N_19621);
and U19902 (N_19902,N_19517,N_19659);
nor U19903 (N_19903,N_19688,N_19730);
and U19904 (N_19904,N_19675,N_19705);
or U19905 (N_19905,N_19549,N_19748);
or U19906 (N_19906,N_19726,N_19720);
nor U19907 (N_19907,N_19540,N_19504);
nand U19908 (N_19908,N_19574,N_19627);
nor U19909 (N_19909,N_19717,N_19525);
nor U19910 (N_19910,N_19683,N_19571);
nand U19911 (N_19911,N_19700,N_19718);
or U19912 (N_19912,N_19529,N_19575);
nand U19913 (N_19913,N_19680,N_19589);
or U19914 (N_19914,N_19745,N_19527);
nand U19915 (N_19915,N_19570,N_19740);
xor U19916 (N_19916,N_19690,N_19706);
xor U19917 (N_19917,N_19563,N_19544);
or U19918 (N_19918,N_19670,N_19586);
or U19919 (N_19919,N_19570,N_19673);
or U19920 (N_19920,N_19553,N_19708);
nand U19921 (N_19921,N_19577,N_19614);
nor U19922 (N_19922,N_19588,N_19672);
or U19923 (N_19923,N_19615,N_19545);
or U19924 (N_19924,N_19544,N_19607);
or U19925 (N_19925,N_19604,N_19615);
or U19926 (N_19926,N_19661,N_19658);
or U19927 (N_19927,N_19562,N_19691);
nand U19928 (N_19928,N_19608,N_19743);
and U19929 (N_19929,N_19517,N_19564);
and U19930 (N_19930,N_19578,N_19709);
xor U19931 (N_19931,N_19664,N_19584);
nor U19932 (N_19932,N_19654,N_19674);
or U19933 (N_19933,N_19698,N_19591);
or U19934 (N_19934,N_19746,N_19552);
xnor U19935 (N_19935,N_19742,N_19666);
and U19936 (N_19936,N_19515,N_19726);
nor U19937 (N_19937,N_19688,N_19620);
xor U19938 (N_19938,N_19702,N_19570);
nand U19939 (N_19939,N_19697,N_19694);
or U19940 (N_19940,N_19743,N_19624);
and U19941 (N_19941,N_19695,N_19626);
and U19942 (N_19942,N_19645,N_19724);
and U19943 (N_19943,N_19593,N_19560);
or U19944 (N_19944,N_19587,N_19519);
or U19945 (N_19945,N_19717,N_19615);
and U19946 (N_19946,N_19678,N_19561);
xnor U19947 (N_19947,N_19644,N_19503);
xor U19948 (N_19948,N_19673,N_19710);
and U19949 (N_19949,N_19633,N_19516);
or U19950 (N_19950,N_19655,N_19558);
nor U19951 (N_19951,N_19699,N_19629);
xnor U19952 (N_19952,N_19622,N_19687);
or U19953 (N_19953,N_19540,N_19745);
or U19954 (N_19954,N_19560,N_19654);
and U19955 (N_19955,N_19717,N_19744);
and U19956 (N_19956,N_19724,N_19582);
and U19957 (N_19957,N_19501,N_19635);
nor U19958 (N_19958,N_19721,N_19515);
or U19959 (N_19959,N_19558,N_19569);
and U19960 (N_19960,N_19735,N_19715);
nand U19961 (N_19961,N_19739,N_19726);
or U19962 (N_19962,N_19552,N_19648);
nand U19963 (N_19963,N_19515,N_19739);
or U19964 (N_19964,N_19679,N_19671);
or U19965 (N_19965,N_19731,N_19682);
xor U19966 (N_19966,N_19709,N_19666);
and U19967 (N_19967,N_19747,N_19622);
xnor U19968 (N_19968,N_19587,N_19570);
nand U19969 (N_19969,N_19519,N_19705);
or U19970 (N_19970,N_19527,N_19513);
and U19971 (N_19971,N_19562,N_19674);
and U19972 (N_19972,N_19625,N_19706);
or U19973 (N_19973,N_19646,N_19664);
nand U19974 (N_19974,N_19708,N_19537);
nor U19975 (N_19975,N_19719,N_19597);
nand U19976 (N_19976,N_19592,N_19663);
xor U19977 (N_19977,N_19517,N_19506);
nand U19978 (N_19978,N_19669,N_19737);
or U19979 (N_19979,N_19505,N_19519);
or U19980 (N_19980,N_19583,N_19518);
nand U19981 (N_19981,N_19626,N_19594);
nand U19982 (N_19982,N_19514,N_19578);
xnor U19983 (N_19983,N_19623,N_19655);
or U19984 (N_19984,N_19509,N_19578);
nor U19985 (N_19985,N_19570,N_19671);
or U19986 (N_19986,N_19561,N_19579);
and U19987 (N_19987,N_19602,N_19633);
or U19988 (N_19988,N_19535,N_19675);
nor U19989 (N_19989,N_19613,N_19720);
nor U19990 (N_19990,N_19558,N_19508);
nand U19991 (N_19991,N_19738,N_19544);
nand U19992 (N_19992,N_19694,N_19565);
nor U19993 (N_19993,N_19630,N_19521);
nor U19994 (N_19994,N_19708,N_19734);
nor U19995 (N_19995,N_19551,N_19618);
xor U19996 (N_19996,N_19517,N_19706);
xnor U19997 (N_19997,N_19679,N_19582);
or U19998 (N_19998,N_19702,N_19699);
and U19999 (N_19999,N_19627,N_19557);
nand U20000 (N_20000,N_19979,N_19804);
or U20001 (N_20001,N_19808,N_19895);
and U20002 (N_20002,N_19883,N_19755);
nand U20003 (N_20003,N_19805,N_19904);
or U20004 (N_20004,N_19809,N_19955);
xnor U20005 (N_20005,N_19980,N_19932);
or U20006 (N_20006,N_19963,N_19996);
nand U20007 (N_20007,N_19941,N_19826);
xor U20008 (N_20008,N_19764,N_19854);
nor U20009 (N_20009,N_19972,N_19918);
xor U20010 (N_20010,N_19978,N_19959);
xnor U20011 (N_20011,N_19900,N_19853);
xor U20012 (N_20012,N_19943,N_19794);
xnor U20013 (N_20013,N_19820,N_19916);
nand U20014 (N_20014,N_19813,N_19757);
and U20015 (N_20015,N_19857,N_19850);
nand U20016 (N_20016,N_19924,N_19989);
nand U20017 (N_20017,N_19935,N_19837);
nor U20018 (N_20018,N_19763,N_19985);
and U20019 (N_20019,N_19872,N_19842);
nand U20020 (N_20020,N_19877,N_19823);
xnor U20021 (N_20021,N_19849,N_19832);
nor U20022 (N_20022,N_19915,N_19840);
xor U20023 (N_20023,N_19876,N_19863);
and U20024 (N_20024,N_19798,N_19843);
or U20025 (N_20025,N_19802,N_19998);
nand U20026 (N_20026,N_19868,N_19896);
or U20027 (N_20027,N_19846,N_19949);
xor U20028 (N_20028,N_19908,N_19881);
xor U20029 (N_20029,N_19884,N_19917);
xnor U20030 (N_20030,N_19759,N_19851);
xnor U20031 (N_20031,N_19889,N_19871);
and U20032 (N_20032,N_19782,N_19973);
xor U20033 (N_20033,N_19909,N_19762);
nand U20034 (N_20034,N_19905,N_19942);
and U20035 (N_20035,N_19761,N_19800);
and U20036 (N_20036,N_19780,N_19928);
and U20037 (N_20037,N_19838,N_19777);
and U20038 (N_20038,N_19776,N_19848);
xnor U20039 (N_20039,N_19930,N_19833);
nand U20040 (N_20040,N_19829,N_19841);
or U20041 (N_20041,N_19811,N_19927);
nor U20042 (N_20042,N_19769,N_19791);
nand U20043 (N_20043,N_19852,N_19903);
nor U20044 (N_20044,N_19750,N_19873);
nand U20045 (N_20045,N_19983,N_19882);
and U20046 (N_20046,N_19938,N_19925);
xor U20047 (N_20047,N_19799,N_19810);
or U20048 (N_20048,N_19987,N_19934);
nor U20049 (N_20049,N_19967,N_19931);
nand U20050 (N_20050,N_19960,N_19752);
and U20051 (N_20051,N_19890,N_19948);
xor U20052 (N_20052,N_19867,N_19806);
or U20053 (N_20053,N_19773,N_19919);
xor U20054 (N_20054,N_19962,N_19751);
nand U20055 (N_20055,N_19879,N_19844);
and U20056 (N_20056,N_19913,N_19830);
nor U20057 (N_20057,N_19785,N_19902);
xor U20058 (N_20058,N_19834,N_19807);
xor U20059 (N_20059,N_19986,N_19779);
nand U20060 (N_20060,N_19767,N_19774);
nor U20061 (N_20061,N_19760,N_19966);
nand U20062 (N_20062,N_19982,N_19910);
nand U20063 (N_20063,N_19961,N_19835);
and U20064 (N_20064,N_19891,N_19864);
or U20065 (N_20065,N_19885,N_19886);
nor U20066 (N_20066,N_19758,N_19839);
xnor U20067 (N_20067,N_19914,N_19944);
and U20068 (N_20068,N_19766,N_19888);
or U20069 (N_20069,N_19819,N_19869);
nand U20070 (N_20070,N_19793,N_19907);
nor U20071 (N_20071,N_19921,N_19906);
or U20072 (N_20072,N_19778,N_19898);
or U20073 (N_20073,N_19874,N_19816);
nand U20074 (N_20074,N_19781,N_19922);
nand U20075 (N_20075,N_19952,N_19964);
nand U20076 (N_20076,N_19754,N_19753);
nor U20077 (N_20077,N_19958,N_19965);
or U20078 (N_20078,N_19855,N_19878);
xor U20079 (N_20079,N_19926,N_19997);
nor U20080 (N_20080,N_19956,N_19920);
or U20081 (N_20081,N_19946,N_19999);
nand U20082 (N_20082,N_19814,N_19976);
nand U20083 (N_20083,N_19772,N_19950);
nor U20084 (N_20084,N_19817,N_19990);
and U20085 (N_20085,N_19975,N_19951);
xnor U20086 (N_20086,N_19968,N_19897);
nor U20087 (N_20087,N_19929,N_19875);
nand U20088 (N_20088,N_19893,N_19825);
and U20089 (N_20089,N_19861,N_19858);
or U20090 (N_20090,N_19933,N_19870);
and U20091 (N_20091,N_19827,N_19866);
or U20092 (N_20092,N_19783,N_19945);
nand U20093 (N_20093,N_19815,N_19912);
and U20094 (N_20094,N_19788,N_19862);
xor U20095 (N_20095,N_19865,N_19790);
nor U20096 (N_20096,N_19818,N_19957);
nand U20097 (N_20097,N_19824,N_19796);
nand U20098 (N_20098,N_19984,N_19981);
and U20099 (N_20099,N_19784,N_19847);
nand U20100 (N_20100,N_19977,N_19899);
nand U20101 (N_20101,N_19939,N_19937);
nor U20102 (N_20102,N_19995,N_19836);
or U20103 (N_20103,N_19993,N_19768);
and U20104 (N_20104,N_19795,N_19947);
xor U20105 (N_20105,N_19792,N_19994);
nand U20106 (N_20106,N_19770,N_19786);
nor U20107 (N_20107,N_19797,N_19765);
and U20108 (N_20108,N_19974,N_19803);
or U20109 (N_20109,N_19821,N_19901);
nand U20110 (N_20110,N_19923,N_19828);
nor U20111 (N_20111,N_19971,N_19940);
or U20112 (N_20112,N_19860,N_19991);
or U20113 (N_20113,N_19831,N_19988);
or U20114 (N_20114,N_19859,N_19954);
and U20115 (N_20115,N_19787,N_19880);
or U20116 (N_20116,N_19845,N_19775);
nand U20117 (N_20117,N_19801,N_19822);
nor U20118 (N_20118,N_19756,N_19992);
nor U20119 (N_20119,N_19970,N_19789);
nand U20120 (N_20120,N_19771,N_19887);
or U20121 (N_20121,N_19856,N_19812);
or U20122 (N_20122,N_19892,N_19953);
and U20123 (N_20123,N_19911,N_19894);
and U20124 (N_20124,N_19969,N_19936);
or U20125 (N_20125,N_19938,N_19891);
nand U20126 (N_20126,N_19855,N_19860);
nand U20127 (N_20127,N_19951,N_19874);
nor U20128 (N_20128,N_19932,N_19862);
nand U20129 (N_20129,N_19837,N_19958);
nand U20130 (N_20130,N_19933,N_19765);
nor U20131 (N_20131,N_19904,N_19854);
xor U20132 (N_20132,N_19963,N_19861);
xor U20133 (N_20133,N_19984,N_19818);
or U20134 (N_20134,N_19965,N_19897);
or U20135 (N_20135,N_19974,N_19908);
or U20136 (N_20136,N_19811,N_19765);
or U20137 (N_20137,N_19980,N_19899);
nand U20138 (N_20138,N_19862,N_19960);
xnor U20139 (N_20139,N_19859,N_19788);
and U20140 (N_20140,N_19864,N_19978);
nor U20141 (N_20141,N_19956,N_19806);
or U20142 (N_20142,N_19921,N_19907);
or U20143 (N_20143,N_19775,N_19934);
or U20144 (N_20144,N_19757,N_19853);
nor U20145 (N_20145,N_19979,N_19838);
nand U20146 (N_20146,N_19805,N_19810);
and U20147 (N_20147,N_19969,N_19889);
and U20148 (N_20148,N_19845,N_19866);
nand U20149 (N_20149,N_19834,N_19961);
nor U20150 (N_20150,N_19999,N_19857);
or U20151 (N_20151,N_19799,N_19821);
and U20152 (N_20152,N_19870,N_19763);
nor U20153 (N_20153,N_19943,N_19995);
nand U20154 (N_20154,N_19940,N_19859);
or U20155 (N_20155,N_19801,N_19839);
nand U20156 (N_20156,N_19834,N_19758);
xor U20157 (N_20157,N_19783,N_19901);
xnor U20158 (N_20158,N_19775,N_19831);
and U20159 (N_20159,N_19998,N_19774);
or U20160 (N_20160,N_19767,N_19971);
or U20161 (N_20161,N_19962,N_19848);
and U20162 (N_20162,N_19803,N_19865);
or U20163 (N_20163,N_19949,N_19959);
nor U20164 (N_20164,N_19887,N_19864);
xor U20165 (N_20165,N_19964,N_19885);
xnor U20166 (N_20166,N_19934,N_19763);
xor U20167 (N_20167,N_19858,N_19868);
and U20168 (N_20168,N_19855,N_19802);
or U20169 (N_20169,N_19919,N_19917);
nand U20170 (N_20170,N_19972,N_19907);
xnor U20171 (N_20171,N_19815,N_19772);
nand U20172 (N_20172,N_19959,N_19796);
xnor U20173 (N_20173,N_19964,N_19965);
and U20174 (N_20174,N_19865,N_19795);
nand U20175 (N_20175,N_19777,N_19866);
or U20176 (N_20176,N_19969,N_19771);
nand U20177 (N_20177,N_19900,N_19978);
xor U20178 (N_20178,N_19879,N_19961);
or U20179 (N_20179,N_19855,N_19974);
or U20180 (N_20180,N_19980,N_19979);
or U20181 (N_20181,N_19754,N_19984);
nor U20182 (N_20182,N_19994,N_19911);
or U20183 (N_20183,N_19978,N_19909);
and U20184 (N_20184,N_19951,N_19809);
or U20185 (N_20185,N_19825,N_19894);
nor U20186 (N_20186,N_19793,N_19811);
nand U20187 (N_20187,N_19786,N_19993);
nand U20188 (N_20188,N_19765,N_19938);
and U20189 (N_20189,N_19773,N_19995);
nor U20190 (N_20190,N_19901,N_19970);
or U20191 (N_20191,N_19910,N_19907);
nand U20192 (N_20192,N_19831,N_19803);
xor U20193 (N_20193,N_19772,N_19968);
xor U20194 (N_20194,N_19883,N_19822);
or U20195 (N_20195,N_19806,N_19788);
xor U20196 (N_20196,N_19930,N_19800);
or U20197 (N_20197,N_19840,N_19795);
nor U20198 (N_20198,N_19958,N_19992);
nor U20199 (N_20199,N_19759,N_19865);
or U20200 (N_20200,N_19930,N_19988);
and U20201 (N_20201,N_19770,N_19949);
or U20202 (N_20202,N_19895,N_19788);
or U20203 (N_20203,N_19956,N_19937);
xnor U20204 (N_20204,N_19757,N_19961);
nand U20205 (N_20205,N_19975,N_19987);
nor U20206 (N_20206,N_19830,N_19815);
nor U20207 (N_20207,N_19953,N_19933);
or U20208 (N_20208,N_19795,N_19992);
nor U20209 (N_20209,N_19883,N_19847);
and U20210 (N_20210,N_19909,N_19755);
nand U20211 (N_20211,N_19852,N_19932);
and U20212 (N_20212,N_19870,N_19900);
xnor U20213 (N_20213,N_19983,N_19814);
xnor U20214 (N_20214,N_19944,N_19864);
nand U20215 (N_20215,N_19942,N_19835);
nor U20216 (N_20216,N_19859,N_19808);
nand U20217 (N_20217,N_19928,N_19908);
nor U20218 (N_20218,N_19922,N_19981);
nor U20219 (N_20219,N_19808,N_19819);
xor U20220 (N_20220,N_19773,N_19756);
nand U20221 (N_20221,N_19751,N_19775);
or U20222 (N_20222,N_19899,N_19902);
nand U20223 (N_20223,N_19752,N_19841);
nand U20224 (N_20224,N_19858,N_19958);
and U20225 (N_20225,N_19877,N_19785);
and U20226 (N_20226,N_19922,N_19815);
or U20227 (N_20227,N_19956,N_19966);
and U20228 (N_20228,N_19862,N_19857);
nor U20229 (N_20229,N_19837,N_19797);
xor U20230 (N_20230,N_19861,N_19790);
or U20231 (N_20231,N_19844,N_19785);
xor U20232 (N_20232,N_19898,N_19970);
xnor U20233 (N_20233,N_19923,N_19805);
xnor U20234 (N_20234,N_19995,N_19790);
xnor U20235 (N_20235,N_19997,N_19883);
nor U20236 (N_20236,N_19764,N_19806);
and U20237 (N_20237,N_19859,N_19858);
nor U20238 (N_20238,N_19975,N_19991);
nand U20239 (N_20239,N_19940,N_19803);
nand U20240 (N_20240,N_19852,N_19842);
and U20241 (N_20241,N_19879,N_19913);
or U20242 (N_20242,N_19858,N_19902);
and U20243 (N_20243,N_19900,N_19915);
xnor U20244 (N_20244,N_19881,N_19826);
and U20245 (N_20245,N_19862,N_19863);
or U20246 (N_20246,N_19865,N_19871);
xor U20247 (N_20247,N_19824,N_19926);
xnor U20248 (N_20248,N_19969,N_19913);
nand U20249 (N_20249,N_19758,N_19938);
xnor U20250 (N_20250,N_20184,N_20123);
or U20251 (N_20251,N_20162,N_20023);
nor U20252 (N_20252,N_20066,N_20174);
xor U20253 (N_20253,N_20095,N_20075);
nor U20254 (N_20254,N_20031,N_20134);
and U20255 (N_20255,N_20070,N_20016);
nor U20256 (N_20256,N_20129,N_20247);
xor U20257 (N_20257,N_20244,N_20165);
or U20258 (N_20258,N_20214,N_20018);
nand U20259 (N_20259,N_20096,N_20013);
nor U20260 (N_20260,N_20086,N_20156);
nor U20261 (N_20261,N_20058,N_20012);
and U20262 (N_20262,N_20190,N_20201);
or U20263 (N_20263,N_20218,N_20039);
nor U20264 (N_20264,N_20178,N_20204);
nand U20265 (N_20265,N_20002,N_20232);
nor U20266 (N_20266,N_20087,N_20206);
nand U20267 (N_20267,N_20237,N_20091);
nor U20268 (N_20268,N_20110,N_20104);
nand U20269 (N_20269,N_20220,N_20215);
and U20270 (N_20270,N_20050,N_20153);
and U20271 (N_20271,N_20065,N_20188);
and U20272 (N_20272,N_20008,N_20005);
nor U20273 (N_20273,N_20027,N_20197);
xor U20274 (N_20274,N_20124,N_20192);
xnor U20275 (N_20275,N_20072,N_20077);
or U20276 (N_20276,N_20235,N_20117);
xor U20277 (N_20277,N_20248,N_20140);
nor U20278 (N_20278,N_20191,N_20239);
nand U20279 (N_20279,N_20047,N_20249);
or U20280 (N_20280,N_20099,N_20120);
nor U20281 (N_20281,N_20037,N_20195);
xor U20282 (N_20282,N_20240,N_20132);
nand U20283 (N_20283,N_20144,N_20126);
nand U20284 (N_20284,N_20207,N_20032);
xor U20285 (N_20285,N_20051,N_20138);
nand U20286 (N_20286,N_20045,N_20168);
nand U20287 (N_20287,N_20131,N_20015);
or U20288 (N_20288,N_20223,N_20097);
or U20289 (N_20289,N_20226,N_20200);
or U20290 (N_20290,N_20114,N_20154);
xnor U20291 (N_20291,N_20073,N_20135);
nand U20292 (N_20292,N_20054,N_20150);
and U20293 (N_20293,N_20147,N_20001);
nand U20294 (N_20294,N_20234,N_20062);
or U20295 (N_20295,N_20186,N_20090);
and U20296 (N_20296,N_20193,N_20042);
nand U20297 (N_20297,N_20143,N_20034);
or U20298 (N_20298,N_20033,N_20222);
or U20299 (N_20299,N_20089,N_20010);
nor U20300 (N_20300,N_20038,N_20189);
xnor U20301 (N_20301,N_20092,N_20020);
nor U20302 (N_20302,N_20246,N_20219);
nor U20303 (N_20303,N_20196,N_20229);
and U20304 (N_20304,N_20169,N_20181);
or U20305 (N_20305,N_20159,N_20171);
nand U20306 (N_20306,N_20083,N_20067);
nor U20307 (N_20307,N_20233,N_20179);
nor U20308 (N_20308,N_20017,N_20202);
or U20309 (N_20309,N_20101,N_20128);
xnor U20310 (N_20310,N_20009,N_20014);
nand U20311 (N_20311,N_20145,N_20216);
xor U20312 (N_20312,N_20228,N_20036);
and U20313 (N_20313,N_20213,N_20041);
and U20314 (N_20314,N_20203,N_20230);
xnor U20315 (N_20315,N_20231,N_20059);
xor U20316 (N_20316,N_20069,N_20113);
xor U20317 (N_20317,N_20139,N_20112);
and U20318 (N_20318,N_20149,N_20060);
nand U20319 (N_20319,N_20172,N_20004);
and U20320 (N_20320,N_20064,N_20071);
nor U20321 (N_20321,N_20238,N_20208);
nand U20322 (N_20322,N_20035,N_20105);
nand U20323 (N_20323,N_20000,N_20084);
xnor U20324 (N_20324,N_20127,N_20227);
xnor U20325 (N_20325,N_20019,N_20155);
nand U20326 (N_20326,N_20068,N_20079);
xor U20327 (N_20327,N_20146,N_20048);
nor U20328 (N_20328,N_20198,N_20103);
or U20329 (N_20329,N_20021,N_20245);
nand U20330 (N_20330,N_20176,N_20024);
and U20331 (N_20331,N_20163,N_20187);
nand U20332 (N_20332,N_20094,N_20183);
xor U20333 (N_20333,N_20107,N_20055);
nor U20334 (N_20334,N_20148,N_20209);
xor U20335 (N_20335,N_20081,N_20082);
or U20336 (N_20336,N_20007,N_20109);
nand U20337 (N_20337,N_20177,N_20056);
or U20338 (N_20338,N_20085,N_20093);
xor U20339 (N_20339,N_20243,N_20043);
and U20340 (N_20340,N_20052,N_20088);
nor U20341 (N_20341,N_20118,N_20166);
xnor U20342 (N_20342,N_20098,N_20011);
nor U20343 (N_20343,N_20063,N_20026);
nand U20344 (N_20344,N_20152,N_20157);
xor U20345 (N_20345,N_20133,N_20044);
nor U20346 (N_20346,N_20080,N_20242);
xnor U20347 (N_20347,N_20116,N_20057);
nor U20348 (N_20348,N_20158,N_20180);
xor U20349 (N_20349,N_20182,N_20211);
xor U20350 (N_20350,N_20210,N_20040);
xnor U20351 (N_20351,N_20161,N_20142);
xnor U20352 (N_20352,N_20061,N_20006);
and U20353 (N_20353,N_20074,N_20167);
nand U20354 (N_20354,N_20130,N_20022);
nand U20355 (N_20355,N_20122,N_20125);
nand U20356 (N_20356,N_20049,N_20108);
xnor U20357 (N_20357,N_20029,N_20225);
or U20358 (N_20358,N_20141,N_20185);
or U20359 (N_20359,N_20194,N_20170);
nand U20360 (N_20360,N_20028,N_20025);
xor U20361 (N_20361,N_20224,N_20030);
and U20362 (N_20362,N_20236,N_20119);
or U20363 (N_20363,N_20102,N_20053);
nor U20364 (N_20364,N_20046,N_20106);
and U20365 (N_20365,N_20199,N_20205);
xnor U20366 (N_20366,N_20221,N_20217);
xor U20367 (N_20367,N_20173,N_20136);
and U20368 (N_20368,N_20212,N_20111);
nand U20369 (N_20369,N_20175,N_20003);
nand U20370 (N_20370,N_20137,N_20078);
xnor U20371 (N_20371,N_20121,N_20115);
and U20372 (N_20372,N_20241,N_20151);
nor U20373 (N_20373,N_20164,N_20160);
xnor U20374 (N_20374,N_20100,N_20076);
and U20375 (N_20375,N_20205,N_20024);
xnor U20376 (N_20376,N_20060,N_20005);
nor U20377 (N_20377,N_20026,N_20145);
or U20378 (N_20378,N_20216,N_20058);
nor U20379 (N_20379,N_20214,N_20185);
and U20380 (N_20380,N_20155,N_20244);
nand U20381 (N_20381,N_20048,N_20057);
xor U20382 (N_20382,N_20156,N_20028);
nor U20383 (N_20383,N_20189,N_20188);
and U20384 (N_20384,N_20091,N_20197);
xor U20385 (N_20385,N_20025,N_20056);
nor U20386 (N_20386,N_20094,N_20006);
nor U20387 (N_20387,N_20004,N_20077);
nor U20388 (N_20388,N_20009,N_20105);
or U20389 (N_20389,N_20113,N_20240);
nor U20390 (N_20390,N_20194,N_20137);
and U20391 (N_20391,N_20072,N_20163);
xor U20392 (N_20392,N_20039,N_20191);
xnor U20393 (N_20393,N_20083,N_20032);
nor U20394 (N_20394,N_20205,N_20017);
nor U20395 (N_20395,N_20201,N_20216);
nand U20396 (N_20396,N_20173,N_20004);
xor U20397 (N_20397,N_20095,N_20194);
and U20398 (N_20398,N_20188,N_20023);
nor U20399 (N_20399,N_20141,N_20115);
xnor U20400 (N_20400,N_20096,N_20151);
xnor U20401 (N_20401,N_20192,N_20236);
xor U20402 (N_20402,N_20011,N_20170);
xnor U20403 (N_20403,N_20069,N_20127);
xnor U20404 (N_20404,N_20159,N_20223);
nor U20405 (N_20405,N_20067,N_20026);
and U20406 (N_20406,N_20151,N_20059);
nor U20407 (N_20407,N_20223,N_20241);
nor U20408 (N_20408,N_20056,N_20023);
or U20409 (N_20409,N_20241,N_20200);
and U20410 (N_20410,N_20191,N_20200);
xnor U20411 (N_20411,N_20109,N_20030);
nand U20412 (N_20412,N_20186,N_20041);
nand U20413 (N_20413,N_20231,N_20216);
or U20414 (N_20414,N_20156,N_20192);
nor U20415 (N_20415,N_20076,N_20138);
and U20416 (N_20416,N_20111,N_20107);
nor U20417 (N_20417,N_20097,N_20023);
and U20418 (N_20418,N_20053,N_20170);
and U20419 (N_20419,N_20128,N_20211);
or U20420 (N_20420,N_20077,N_20127);
and U20421 (N_20421,N_20070,N_20246);
nand U20422 (N_20422,N_20135,N_20036);
or U20423 (N_20423,N_20120,N_20111);
xnor U20424 (N_20424,N_20043,N_20011);
xor U20425 (N_20425,N_20186,N_20225);
nand U20426 (N_20426,N_20195,N_20209);
xnor U20427 (N_20427,N_20087,N_20200);
nor U20428 (N_20428,N_20041,N_20169);
xor U20429 (N_20429,N_20006,N_20114);
xnor U20430 (N_20430,N_20012,N_20187);
or U20431 (N_20431,N_20019,N_20076);
or U20432 (N_20432,N_20158,N_20061);
and U20433 (N_20433,N_20083,N_20239);
nor U20434 (N_20434,N_20074,N_20044);
xnor U20435 (N_20435,N_20145,N_20172);
nand U20436 (N_20436,N_20146,N_20009);
nand U20437 (N_20437,N_20066,N_20199);
nor U20438 (N_20438,N_20063,N_20104);
nor U20439 (N_20439,N_20129,N_20017);
nand U20440 (N_20440,N_20072,N_20145);
nor U20441 (N_20441,N_20147,N_20177);
xor U20442 (N_20442,N_20056,N_20026);
nand U20443 (N_20443,N_20026,N_20098);
nand U20444 (N_20444,N_20194,N_20037);
nor U20445 (N_20445,N_20073,N_20166);
or U20446 (N_20446,N_20053,N_20219);
or U20447 (N_20447,N_20040,N_20212);
and U20448 (N_20448,N_20188,N_20183);
and U20449 (N_20449,N_20237,N_20109);
nor U20450 (N_20450,N_20002,N_20209);
nor U20451 (N_20451,N_20132,N_20190);
nor U20452 (N_20452,N_20069,N_20200);
nand U20453 (N_20453,N_20137,N_20005);
xor U20454 (N_20454,N_20052,N_20132);
nand U20455 (N_20455,N_20156,N_20191);
xor U20456 (N_20456,N_20214,N_20213);
and U20457 (N_20457,N_20135,N_20035);
nand U20458 (N_20458,N_20049,N_20088);
or U20459 (N_20459,N_20187,N_20115);
and U20460 (N_20460,N_20218,N_20211);
xnor U20461 (N_20461,N_20058,N_20056);
nor U20462 (N_20462,N_20141,N_20072);
and U20463 (N_20463,N_20071,N_20044);
and U20464 (N_20464,N_20156,N_20221);
or U20465 (N_20465,N_20248,N_20078);
or U20466 (N_20466,N_20200,N_20013);
or U20467 (N_20467,N_20179,N_20144);
or U20468 (N_20468,N_20236,N_20163);
or U20469 (N_20469,N_20076,N_20027);
nor U20470 (N_20470,N_20180,N_20120);
xnor U20471 (N_20471,N_20170,N_20225);
or U20472 (N_20472,N_20143,N_20177);
nor U20473 (N_20473,N_20138,N_20238);
and U20474 (N_20474,N_20087,N_20042);
nor U20475 (N_20475,N_20086,N_20074);
and U20476 (N_20476,N_20081,N_20143);
or U20477 (N_20477,N_20073,N_20072);
and U20478 (N_20478,N_20106,N_20074);
nor U20479 (N_20479,N_20165,N_20119);
or U20480 (N_20480,N_20075,N_20089);
or U20481 (N_20481,N_20135,N_20157);
or U20482 (N_20482,N_20076,N_20242);
nand U20483 (N_20483,N_20054,N_20219);
or U20484 (N_20484,N_20213,N_20239);
or U20485 (N_20485,N_20033,N_20170);
and U20486 (N_20486,N_20061,N_20081);
and U20487 (N_20487,N_20194,N_20203);
or U20488 (N_20488,N_20087,N_20114);
or U20489 (N_20489,N_20051,N_20122);
and U20490 (N_20490,N_20243,N_20248);
nor U20491 (N_20491,N_20069,N_20111);
nand U20492 (N_20492,N_20241,N_20092);
and U20493 (N_20493,N_20088,N_20244);
or U20494 (N_20494,N_20093,N_20099);
xor U20495 (N_20495,N_20028,N_20034);
xnor U20496 (N_20496,N_20010,N_20227);
or U20497 (N_20497,N_20217,N_20048);
xnor U20498 (N_20498,N_20243,N_20169);
or U20499 (N_20499,N_20246,N_20083);
nor U20500 (N_20500,N_20334,N_20357);
nand U20501 (N_20501,N_20268,N_20387);
and U20502 (N_20502,N_20476,N_20296);
xnor U20503 (N_20503,N_20282,N_20408);
nand U20504 (N_20504,N_20265,N_20370);
or U20505 (N_20505,N_20270,N_20439);
or U20506 (N_20506,N_20393,N_20330);
or U20507 (N_20507,N_20478,N_20269);
nor U20508 (N_20508,N_20398,N_20451);
or U20509 (N_20509,N_20498,N_20454);
or U20510 (N_20510,N_20317,N_20493);
nand U20511 (N_20511,N_20427,N_20487);
or U20512 (N_20512,N_20436,N_20302);
and U20513 (N_20513,N_20336,N_20329);
nor U20514 (N_20514,N_20348,N_20466);
or U20515 (N_20515,N_20252,N_20327);
nor U20516 (N_20516,N_20338,N_20497);
or U20517 (N_20517,N_20346,N_20444);
or U20518 (N_20518,N_20422,N_20304);
xnor U20519 (N_20519,N_20312,N_20443);
nor U20520 (N_20520,N_20311,N_20409);
and U20521 (N_20521,N_20335,N_20486);
or U20522 (N_20522,N_20496,N_20288);
or U20523 (N_20523,N_20379,N_20449);
and U20524 (N_20524,N_20314,N_20353);
xor U20525 (N_20525,N_20301,N_20303);
nor U20526 (N_20526,N_20354,N_20435);
and U20527 (N_20527,N_20473,N_20331);
and U20528 (N_20528,N_20416,N_20445);
or U20529 (N_20529,N_20489,N_20448);
nor U20530 (N_20530,N_20321,N_20294);
nand U20531 (N_20531,N_20440,N_20446);
and U20532 (N_20532,N_20310,N_20428);
xnor U20533 (N_20533,N_20452,N_20433);
nand U20534 (N_20534,N_20365,N_20299);
and U20535 (N_20535,N_20319,N_20295);
and U20536 (N_20536,N_20350,N_20482);
and U20537 (N_20537,N_20495,N_20467);
xnor U20538 (N_20538,N_20341,N_20429);
and U20539 (N_20539,N_20332,N_20363);
or U20540 (N_20540,N_20279,N_20470);
nor U20541 (N_20541,N_20384,N_20391);
nand U20542 (N_20542,N_20257,N_20396);
xnor U20543 (N_20543,N_20281,N_20383);
xor U20544 (N_20544,N_20259,N_20456);
nand U20545 (N_20545,N_20277,N_20441);
and U20546 (N_20546,N_20455,N_20472);
nor U20547 (N_20547,N_20260,N_20380);
xnor U20548 (N_20548,N_20372,N_20479);
nor U20549 (N_20549,N_20438,N_20434);
nor U20550 (N_20550,N_20395,N_20460);
or U20551 (N_20551,N_20490,N_20300);
xnor U20552 (N_20552,N_20425,N_20392);
and U20553 (N_20553,N_20404,N_20366);
or U20554 (N_20554,N_20488,N_20356);
xnor U20555 (N_20555,N_20305,N_20307);
or U20556 (N_20556,N_20426,N_20377);
or U20557 (N_20557,N_20283,N_20458);
and U20558 (N_20558,N_20323,N_20275);
nor U20559 (N_20559,N_20287,N_20369);
nor U20560 (N_20560,N_20289,N_20273);
nor U20561 (N_20561,N_20390,N_20367);
xnor U20562 (N_20562,N_20388,N_20274);
xor U20563 (N_20563,N_20461,N_20264);
or U20564 (N_20564,N_20381,N_20421);
nand U20565 (N_20565,N_20320,N_20253);
xor U20566 (N_20566,N_20316,N_20293);
nand U20567 (N_20567,N_20278,N_20457);
nor U20568 (N_20568,N_20345,N_20328);
and U20569 (N_20569,N_20385,N_20415);
and U20570 (N_20570,N_20297,N_20453);
or U20571 (N_20571,N_20437,N_20306);
nor U20572 (N_20572,N_20250,N_20378);
and U20573 (N_20573,N_20399,N_20352);
or U20574 (N_20574,N_20373,N_20413);
or U20575 (N_20575,N_20462,N_20285);
nand U20576 (N_20576,N_20477,N_20412);
and U20577 (N_20577,N_20258,N_20469);
or U20578 (N_20578,N_20267,N_20480);
or U20579 (N_20579,N_20360,N_20405);
or U20580 (N_20580,N_20411,N_20255);
nand U20581 (N_20581,N_20344,N_20355);
and U20582 (N_20582,N_20464,N_20376);
xnor U20583 (N_20583,N_20263,N_20347);
or U20584 (N_20584,N_20397,N_20359);
nor U20585 (N_20585,N_20430,N_20484);
nor U20586 (N_20586,N_20271,N_20417);
nand U20587 (N_20587,N_20322,N_20400);
nor U20588 (N_20588,N_20483,N_20474);
and U20589 (N_20589,N_20292,N_20286);
nand U20590 (N_20590,N_20406,N_20368);
xor U20591 (N_20591,N_20342,N_20468);
nor U20592 (N_20592,N_20313,N_20272);
nor U20593 (N_20593,N_20308,N_20471);
nor U20594 (N_20594,N_20419,N_20326);
xor U20595 (N_20595,N_20485,N_20340);
or U20596 (N_20596,N_20339,N_20261);
and U20597 (N_20597,N_20315,N_20333);
and U20598 (N_20598,N_20499,N_20362);
nand U20599 (N_20599,N_20349,N_20343);
and U20600 (N_20600,N_20401,N_20491);
nor U20601 (N_20601,N_20254,N_20318);
xnor U20602 (N_20602,N_20459,N_20374);
nand U20603 (N_20603,N_20325,N_20291);
and U20604 (N_20604,N_20423,N_20337);
nand U20605 (N_20605,N_20402,N_20361);
nand U20606 (N_20606,N_20298,N_20442);
or U20607 (N_20607,N_20463,N_20410);
nor U20608 (N_20608,N_20280,N_20403);
and U20609 (N_20609,N_20432,N_20371);
xnor U20610 (N_20610,N_20389,N_20309);
and U20611 (N_20611,N_20358,N_20418);
nand U20612 (N_20612,N_20266,N_20494);
nand U20613 (N_20613,N_20382,N_20492);
and U20614 (N_20614,N_20256,N_20262);
and U20615 (N_20615,N_20431,N_20465);
or U20616 (N_20616,N_20447,N_20290);
and U20617 (N_20617,N_20284,N_20276);
and U20618 (N_20618,N_20450,N_20420);
nand U20619 (N_20619,N_20375,N_20251);
or U20620 (N_20620,N_20364,N_20407);
and U20621 (N_20621,N_20394,N_20475);
and U20622 (N_20622,N_20386,N_20414);
and U20623 (N_20623,N_20424,N_20351);
nor U20624 (N_20624,N_20324,N_20481);
or U20625 (N_20625,N_20390,N_20299);
and U20626 (N_20626,N_20415,N_20449);
or U20627 (N_20627,N_20350,N_20304);
nand U20628 (N_20628,N_20483,N_20256);
nor U20629 (N_20629,N_20452,N_20356);
nor U20630 (N_20630,N_20328,N_20257);
nand U20631 (N_20631,N_20259,N_20485);
xnor U20632 (N_20632,N_20409,N_20270);
and U20633 (N_20633,N_20344,N_20341);
nand U20634 (N_20634,N_20445,N_20303);
or U20635 (N_20635,N_20285,N_20459);
xnor U20636 (N_20636,N_20331,N_20374);
nand U20637 (N_20637,N_20441,N_20432);
nand U20638 (N_20638,N_20308,N_20438);
nor U20639 (N_20639,N_20430,N_20424);
and U20640 (N_20640,N_20275,N_20443);
xnor U20641 (N_20641,N_20465,N_20318);
nand U20642 (N_20642,N_20359,N_20408);
nor U20643 (N_20643,N_20302,N_20491);
nand U20644 (N_20644,N_20260,N_20367);
or U20645 (N_20645,N_20257,N_20283);
and U20646 (N_20646,N_20389,N_20283);
xnor U20647 (N_20647,N_20327,N_20291);
nand U20648 (N_20648,N_20261,N_20464);
xnor U20649 (N_20649,N_20387,N_20403);
nand U20650 (N_20650,N_20331,N_20319);
or U20651 (N_20651,N_20408,N_20431);
nor U20652 (N_20652,N_20358,N_20490);
or U20653 (N_20653,N_20366,N_20457);
nor U20654 (N_20654,N_20423,N_20474);
xnor U20655 (N_20655,N_20472,N_20417);
or U20656 (N_20656,N_20443,N_20436);
xnor U20657 (N_20657,N_20490,N_20408);
xnor U20658 (N_20658,N_20329,N_20404);
and U20659 (N_20659,N_20281,N_20480);
nor U20660 (N_20660,N_20431,N_20467);
nand U20661 (N_20661,N_20425,N_20372);
or U20662 (N_20662,N_20372,N_20349);
xor U20663 (N_20663,N_20499,N_20438);
or U20664 (N_20664,N_20456,N_20273);
nand U20665 (N_20665,N_20412,N_20265);
nand U20666 (N_20666,N_20276,N_20266);
nor U20667 (N_20667,N_20264,N_20274);
and U20668 (N_20668,N_20301,N_20264);
nor U20669 (N_20669,N_20261,N_20439);
and U20670 (N_20670,N_20378,N_20419);
nor U20671 (N_20671,N_20258,N_20459);
nor U20672 (N_20672,N_20250,N_20407);
nand U20673 (N_20673,N_20381,N_20440);
nor U20674 (N_20674,N_20298,N_20426);
nor U20675 (N_20675,N_20479,N_20476);
nor U20676 (N_20676,N_20264,N_20357);
and U20677 (N_20677,N_20334,N_20327);
and U20678 (N_20678,N_20498,N_20314);
nand U20679 (N_20679,N_20466,N_20373);
or U20680 (N_20680,N_20345,N_20305);
and U20681 (N_20681,N_20331,N_20477);
nand U20682 (N_20682,N_20441,N_20310);
nand U20683 (N_20683,N_20374,N_20466);
xnor U20684 (N_20684,N_20498,N_20364);
nand U20685 (N_20685,N_20433,N_20441);
xnor U20686 (N_20686,N_20284,N_20427);
nand U20687 (N_20687,N_20462,N_20269);
nand U20688 (N_20688,N_20258,N_20272);
or U20689 (N_20689,N_20363,N_20385);
xor U20690 (N_20690,N_20383,N_20390);
or U20691 (N_20691,N_20381,N_20480);
xor U20692 (N_20692,N_20286,N_20426);
and U20693 (N_20693,N_20476,N_20294);
xor U20694 (N_20694,N_20375,N_20294);
xor U20695 (N_20695,N_20372,N_20329);
and U20696 (N_20696,N_20389,N_20254);
nor U20697 (N_20697,N_20436,N_20318);
xnor U20698 (N_20698,N_20459,N_20325);
xor U20699 (N_20699,N_20288,N_20269);
and U20700 (N_20700,N_20283,N_20307);
and U20701 (N_20701,N_20271,N_20265);
xnor U20702 (N_20702,N_20488,N_20352);
or U20703 (N_20703,N_20366,N_20280);
and U20704 (N_20704,N_20398,N_20257);
nand U20705 (N_20705,N_20335,N_20290);
nand U20706 (N_20706,N_20388,N_20283);
nand U20707 (N_20707,N_20312,N_20355);
and U20708 (N_20708,N_20458,N_20492);
nand U20709 (N_20709,N_20311,N_20452);
and U20710 (N_20710,N_20337,N_20394);
nand U20711 (N_20711,N_20489,N_20301);
nand U20712 (N_20712,N_20430,N_20399);
nor U20713 (N_20713,N_20497,N_20392);
and U20714 (N_20714,N_20409,N_20360);
or U20715 (N_20715,N_20341,N_20269);
nand U20716 (N_20716,N_20293,N_20468);
nand U20717 (N_20717,N_20271,N_20277);
or U20718 (N_20718,N_20496,N_20457);
and U20719 (N_20719,N_20273,N_20436);
and U20720 (N_20720,N_20339,N_20438);
nor U20721 (N_20721,N_20307,N_20471);
and U20722 (N_20722,N_20315,N_20290);
or U20723 (N_20723,N_20423,N_20283);
nor U20724 (N_20724,N_20467,N_20394);
nand U20725 (N_20725,N_20452,N_20448);
nor U20726 (N_20726,N_20270,N_20407);
nor U20727 (N_20727,N_20387,N_20366);
nor U20728 (N_20728,N_20381,N_20303);
or U20729 (N_20729,N_20393,N_20407);
or U20730 (N_20730,N_20446,N_20291);
xnor U20731 (N_20731,N_20270,N_20319);
nand U20732 (N_20732,N_20331,N_20341);
or U20733 (N_20733,N_20286,N_20466);
nor U20734 (N_20734,N_20405,N_20335);
nor U20735 (N_20735,N_20416,N_20419);
nor U20736 (N_20736,N_20325,N_20490);
xor U20737 (N_20737,N_20274,N_20280);
or U20738 (N_20738,N_20448,N_20356);
or U20739 (N_20739,N_20383,N_20468);
xor U20740 (N_20740,N_20356,N_20446);
or U20741 (N_20741,N_20370,N_20472);
nor U20742 (N_20742,N_20354,N_20342);
nor U20743 (N_20743,N_20263,N_20264);
xor U20744 (N_20744,N_20357,N_20491);
xor U20745 (N_20745,N_20305,N_20431);
or U20746 (N_20746,N_20290,N_20363);
and U20747 (N_20747,N_20457,N_20312);
nand U20748 (N_20748,N_20369,N_20497);
or U20749 (N_20749,N_20427,N_20290);
or U20750 (N_20750,N_20686,N_20706);
nor U20751 (N_20751,N_20638,N_20612);
nand U20752 (N_20752,N_20684,N_20741);
nand U20753 (N_20753,N_20502,N_20565);
and U20754 (N_20754,N_20501,N_20649);
or U20755 (N_20755,N_20731,N_20717);
and U20756 (N_20756,N_20653,N_20722);
nor U20757 (N_20757,N_20572,N_20549);
xor U20758 (N_20758,N_20521,N_20512);
or U20759 (N_20759,N_20742,N_20744);
xor U20760 (N_20760,N_20506,N_20602);
nor U20761 (N_20761,N_20627,N_20635);
nor U20762 (N_20762,N_20743,N_20654);
nand U20763 (N_20763,N_20663,N_20678);
and U20764 (N_20764,N_20625,N_20724);
nor U20765 (N_20765,N_20639,N_20661);
and U20766 (N_20766,N_20631,N_20651);
nand U20767 (N_20767,N_20526,N_20548);
nand U20768 (N_20768,N_20746,N_20725);
xor U20769 (N_20769,N_20626,N_20566);
nand U20770 (N_20770,N_20593,N_20536);
and U20771 (N_20771,N_20504,N_20564);
nor U20772 (N_20772,N_20621,N_20718);
nor U20773 (N_20773,N_20580,N_20695);
or U20774 (N_20774,N_20587,N_20532);
nor U20775 (N_20775,N_20575,N_20543);
nor U20776 (N_20776,N_20640,N_20599);
or U20777 (N_20777,N_20540,N_20700);
or U20778 (N_20778,N_20614,N_20708);
xor U20779 (N_20779,N_20609,N_20582);
and U20780 (N_20780,N_20728,N_20520);
nand U20781 (N_20781,N_20545,N_20642);
xnor U20782 (N_20782,N_20527,N_20737);
nor U20783 (N_20783,N_20507,N_20542);
nor U20784 (N_20784,N_20522,N_20705);
xor U20785 (N_20785,N_20664,N_20616);
nand U20786 (N_20786,N_20714,N_20675);
and U20787 (N_20787,N_20607,N_20622);
nand U20788 (N_20788,N_20531,N_20538);
xnor U20789 (N_20789,N_20672,N_20516);
nand U20790 (N_20790,N_20608,N_20559);
xor U20791 (N_20791,N_20674,N_20689);
and U20792 (N_20792,N_20569,N_20681);
nor U20793 (N_20793,N_20628,N_20657);
nor U20794 (N_20794,N_20707,N_20665);
or U20795 (N_20795,N_20747,N_20552);
or U20796 (N_20796,N_20676,N_20513);
nand U20797 (N_20797,N_20690,N_20603);
nor U20798 (N_20798,N_20732,N_20528);
and U20799 (N_20799,N_20636,N_20594);
nand U20800 (N_20800,N_20656,N_20685);
and U20801 (N_20801,N_20601,N_20604);
or U20802 (N_20802,N_20697,N_20534);
and U20803 (N_20803,N_20720,N_20605);
xnor U20804 (N_20804,N_20677,N_20630);
xor U20805 (N_20805,N_20620,N_20694);
nand U20806 (N_20806,N_20586,N_20592);
or U20807 (N_20807,N_20632,N_20735);
or U20808 (N_20808,N_20734,N_20597);
or U20809 (N_20809,N_20644,N_20711);
xor U20810 (N_20810,N_20733,N_20698);
nand U20811 (N_20811,N_20629,N_20637);
nand U20812 (N_20812,N_20576,N_20558);
or U20813 (N_20813,N_20633,N_20519);
nand U20814 (N_20814,N_20573,N_20693);
nor U20815 (N_20815,N_20500,N_20583);
nand U20816 (N_20816,N_20715,N_20748);
nor U20817 (N_20817,N_20702,N_20557);
xor U20818 (N_20818,N_20589,N_20659);
and U20819 (N_20819,N_20551,N_20567);
and U20820 (N_20820,N_20688,N_20683);
and U20821 (N_20821,N_20739,N_20666);
or U20822 (N_20822,N_20553,N_20525);
nor U20823 (N_20823,N_20648,N_20547);
nand U20824 (N_20824,N_20533,N_20703);
nor U20825 (N_20825,N_20515,N_20562);
nand U20826 (N_20826,N_20669,N_20709);
nor U20827 (N_20827,N_20544,N_20554);
nand U20828 (N_20828,N_20726,N_20730);
or U20829 (N_20829,N_20598,N_20568);
nand U20830 (N_20830,N_20618,N_20574);
xor U20831 (N_20831,N_20518,N_20736);
nand U20832 (N_20832,N_20643,N_20523);
nand U20833 (N_20833,N_20541,N_20530);
nand U20834 (N_20834,N_20712,N_20581);
nand U20835 (N_20835,N_20606,N_20670);
xnor U20836 (N_20836,N_20671,N_20723);
or U20837 (N_20837,N_20591,N_20660);
and U20838 (N_20838,N_20577,N_20539);
and U20839 (N_20839,N_20578,N_20641);
and U20840 (N_20840,N_20595,N_20655);
and U20841 (N_20841,N_20619,N_20563);
and U20842 (N_20842,N_20550,N_20613);
xor U20843 (N_20843,N_20687,N_20647);
and U20844 (N_20844,N_20571,N_20679);
xnor U20845 (N_20845,N_20509,N_20588);
nor U20846 (N_20846,N_20652,N_20645);
or U20847 (N_20847,N_20727,N_20740);
and U20848 (N_20848,N_20600,N_20617);
or U20849 (N_20849,N_20611,N_20503);
and U20850 (N_20850,N_20555,N_20721);
or U20851 (N_20851,N_20658,N_20745);
xnor U20852 (N_20852,N_20529,N_20535);
xnor U20853 (N_20853,N_20710,N_20514);
nand U20854 (N_20854,N_20624,N_20680);
nor U20855 (N_20855,N_20570,N_20713);
xnor U20856 (N_20856,N_20738,N_20623);
nand U20857 (N_20857,N_20561,N_20696);
nor U20858 (N_20858,N_20662,N_20584);
xor U20859 (N_20859,N_20634,N_20505);
nor U20860 (N_20860,N_20585,N_20749);
or U20861 (N_20861,N_20691,N_20650);
xor U20862 (N_20862,N_20524,N_20615);
nand U20863 (N_20863,N_20517,N_20556);
nand U20864 (N_20864,N_20729,N_20646);
and U20865 (N_20865,N_20719,N_20699);
and U20866 (N_20866,N_20560,N_20508);
or U20867 (N_20867,N_20537,N_20682);
or U20868 (N_20868,N_20716,N_20511);
xnor U20869 (N_20869,N_20579,N_20673);
and U20870 (N_20870,N_20590,N_20510);
xnor U20871 (N_20871,N_20610,N_20667);
xor U20872 (N_20872,N_20701,N_20704);
xor U20873 (N_20873,N_20546,N_20692);
nand U20874 (N_20874,N_20668,N_20596);
nor U20875 (N_20875,N_20666,N_20591);
xnor U20876 (N_20876,N_20637,N_20744);
nand U20877 (N_20877,N_20633,N_20698);
nor U20878 (N_20878,N_20678,N_20615);
or U20879 (N_20879,N_20666,N_20712);
and U20880 (N_20880,N_20643,N_20578);
nand U20881 (N_20881,N_20567,N_20639);
or U20882 (N_20882,N_20535,N_20724);
xnor U20883 (N_20883,N_20679,N_20545);
nand U20884 (N_20884,N_20707,N_20601);
and U20885 (N_20885,N_20625,N_20669);
or U20886 (N_20886,N_20614,N_20671);
and U20887 (N_20887,N_20738,N_20704);
nand U20888 (N_20888,N_20628,N_20593);
xor U20889 (N_20889,N_20532,N_20667);
xor U20890 (N_20890,N_20668,N_20686);
xor U20891 (N_20891,N_20735,N_20749);
and U20892 (N_20892,N_20725,N_20598);
nor U20893 (N_20893,N_20530,N_20502);
or U20894 (N_20894,N_20614,N_20652);
or U20895 (N_20895,N_20607,N_20603);
nor U20896 (N_20896,N_20687,N_20660);
or U20897 (N_20897,N_20596,N_20601);
nand U20898 (N_20898,N_20552,N_20618);
nand U20899 (N_20899,N_20603,N_20737);
nor U20900 (N_20900,N_20654,N_20683);
nor U20901 (N_20901,N_20721,N_20578);
or U20902 (N_20902,N_20689,N_20539);
and U20903 (N_20903,N_20712,N_20694);
nor U20904 (N_20904,N_20509,N_20695);
xnor U20905 (N_20905,N_20729,N_20547);
nor U20906 (N_20906,N_20681,N_20510);
or U20907 (N_20907,N_20742,N_20732);
and U20908 (N_20908,N_20713,N_20691);
xor U20909 (N_20909,N_20702,N_20584);
nor U20910 (N_20910,N_20623,N_20642);
nand U20911 (N_20911,N_20643,N_20615);
and U20912 (N_20912,N_20716,N_20614);
xor U20913 (N_20913,N_20704,N_20533);
nand U20914 (N_20914,N_20542,N_20656);
xnor U20915 (N_20915,N_20664,N_20707);
xnor U20916 (N_20916,N_20580,N_20513);
and U20917 (N_20917,N_20680,N_20523);
nor U20918 (N_20918,N_20544,N_20574);
nor U20919 (N_20919,N_20684,N_20693);
xor U20920 (N_20920,N_20542,N_20593);
or U20921 (N_20921,N_20617,N_20596);
xor U20922 (N_20922,N_20657,N_20723);
or U20923 (N_20923,N_20553,N_20654);
nor U20924 (N_20924,N_20546,N_20571);
or U20925 (N_20925,N_20515,N_20727);
nor U20926 (N_20926,N_20612,N_20680);
xnor U20927 (N_20927,N_20580,N_20548);
nor U20928 (N_20928,N_20636,N_20628);
or U20929 (N_20929,N_20551,N_20657);
nand U20930 (N_20930,N_20673,N_20743);
nor U20931 (N_20931,N_20595,N_20588);
or U20932 (N_20932,N_20736,N_20641);
nand U20933 (N_20933,N_20553,N_20697);
or U20934 (N_20934,N_20646,N_20631);
or U20935 (N_20935,N_20536,N_20542);
or U20936 (N_20936,N_20581,N_20607);
or U20937 (N_20937,N_20590,N_20641);
xor U20938 (N_20938,N_20679,N_20649);
and U20939 (N_20939,N_20649,N_20732);
nand U20940 (N_20940,N_20588,N_20623);
nor U20941 (N_20941,N_20679,N_20591);
nor U20942 (N_20942,N_20711,N_20522);
nand U20943 (N_20943,N_20717,N_20594);
nand U20944 (N_20944,N_20522,N_20619);
nor U20945 (N_20945,N_20625,N_20605);
or U20946 (N_20946,N_20694,N_20744);
nand U20947 (N_20947,N_20561,N_20523);
xnor U20948 (N_20948,N_20536,N_20741);
xnor U20949 (N_20949,N_20563,N_20548);
nor U20950 (N_20950,N_20683,N_20696);
xnor U20951 (N_20951,N_20726,N_20679);
nand U20952 (N_20952,N_20541,N_20538);
nand U20953 (N_20953,N_20649,N_20654);
and U20954 (N_20954,N_20685,N_20576);
xnor U20955 (N_20955,N_20567,N_20525);
and U20956 (N_20956,N_20574,N_20672);
and U20957 (N_20957,N_20655,N_20585);
xnor U20958 (N_20958,N_20699,N_20623);
xor U20959 (N_20959,N_20674,N_20550);
nand U20960 (N_20960,N_20625,N_20536);
nor U20961 (N_20961,N_20607,N_20661);
nor U20962 (N_20962,N_20745,N_20598);
xor U20963 (N_20963,N_20558,N_20505);
and U20964 (N_20964,N_20590,N_20532);
xnor U20965 (N_20965,N_20570,N_20673);
xnor U20966 (N_20966,N_20699,N_20676);
xnor U20967 (N_20967,N_20506,N_20637);
or U20968 (N_20968,N_20556,N_20591);
nor U20969 (N_20969,N_20526,N_20682);
nand U20970 (N_20970,N_20596,N_20602);
nor U20971 (N_20971,N_20618,N_20566);
nand U20972 (N_20972,N_20693,N_20688);
xor U20973 (N_20973,N_20563,N_20544);
xor U20974 (N_20974,N_20659,N_20522);
nor U20975 (N_20975,N_20531,N_20585);
or U20976 (N_20976,N_20738,N_20739);
nor U20977 (N_20977,N_20659,N_20602);
nor U20978 (N_20978,N_20739,N_20704);
and U20979 (N_20979,N_20548,N_20656);
or U20980 (N_20980,N_20582,N_20554);
nand U20981 (N_20981,N_20719,N_20539);
nand U20982 (N_20982,N_20504,N_20716);
nor U20983 (N_20983,N_20552,N_20545);
nor U20984 (N_20984,N_20571,N_20552);
and U20985 (N_20985,N_20630,N_20710);
or U20986 (N_20986,N_20614,N_20690);
and U20987 (N_20987,N_20738,N_20725);
xor U20988 (N_20988,N_20732,N_20546);
nor U20989 (N_20989,N_20620,N_20593);
nand U20990 (N_20990,N_20632,N_20598);
and U20991 (N_20991,N_20667,N_20714);
and U20992 (N_20992,N_20696,N_20619);
nand U20993 (N_20993,N_20629,N_20657);
xnor U20994 (N_20994,N_20627,N_20666);
and U20995 (N_20995,N_20505,N_20612);
xor U20996 (N_20996,N_20736,N_20614);
and U20997 (N_20997,N_20702,N_20734);
xnor U20998 (N_20998,N_20681,N_20632);
or U20999 (N_20999,N_20670,N_20713);
and U21000 (N_21000,N_20800,N_20999);
xnor U21001 (N_21001,N_20859,N_20909);
nor U21002 (N_21002,N_20759,N_20823);
and U21003 (N_21003,N_20952,N_20946);
and U21004 (N_21004,N_20850,N_20878);
and U21005 (N_21005,N_20791,N_20920);
or U21006 (N_21006,N_20788,N_20911);
nand U21007 (N_21007,N_20940,N_20983);
nor U21008 (N_21008,N_20831,N_20921);
or U21009 (N_21009,N_20972,N_20836);
and U21010 (N_21010,N_20906,N_20846);
xnor U21011 (N_21011,N_20916,N_20973);
nor U21012 (N_21012,N_20755,N_20847);
nand U21013 (N_21013,N_20774,N_20996);
nor U21014 (N_21014,N_20821,N_20751);
nand U21015 (N_21015,N_20867,N_20876);
nor U21016 (N_21016,N_20785,N_20837);
or U21017 (N_21017,N_20956,N_20765);
and U21018 (N_21018,N_20967,N_20805);
nand U21019 (N_21019,N_20769,N_20919);
and U21020 (N_21020,N_20816,N_20969);
nand U21021 (N_21021,N_20994,N_20779);
nand U21022 (N_21022,N_20950,N_20943);
nand U21023 (N_21023,N_20976,N_20776);
or U21024 (N_21024,N_20792,N_20866);
and U21025 (N_21025,N_20913,N_20945);
and U21026 (N_21026,N_20966,N_20980);
xnor U21027 (N_21027,N_20822,N_20982);
or U21028 (N_21028,N_20926,N_20908);
or U21029 (N_21029,N_20931,N_20869);
or U21030 (N_21030,N_20885,N_20957);
and U21031 (N_21031,N_20937,N_20958);
nand U21032 (N_21032,N_20806,N_20812);
nor U21033 (N_21033,N_20933,N_20875);
nand U21034 (N_21034,N_20883,N_20796);
nand U21035 (N_21035,N_20891,N_20760);
and U21036 (N_21036,N_20750,N_20888);
and U21037 (N_21037,N_20862,N_20993);
nand U21038 (N_21038,N_20863,N_20855);
nand U21039 (N_21039,N_20762,N_20948);
nand U21040 (N_21040,N_20947,N_20842);
or U21041 (N_21041,N_20826,N_20808);
nor U21042 (N_21042,N_20813,N_20893);
and U21043 (N_21043,N_20934,N_20971);
or U21044 (N_21044,N_20927,N_20907);
nor U21045 (N_21045,N_20900,N_20984);
nor U21046 (N_21046,N_20845,N_20793);
and U21047 (N_21047,N_20865,N_20778);
nor U21048 (N_21048,N_20914,N_20897);
nand U21049 (N_21049,N_20757,N_20917);
and U21050 (N_21050,N_20942,N_20861);
and U21051 (N_21051,N_20856,N_20928);
or U21052 (N_21052,N_20879,N_20789);
nor U21053 (N_21053,N_20987,N_20781);
nor U21054 (N_21054,N_20756,N_20870);
and U21055 (N_21055,N_20777,N_20895);
or U21056 (N_21056,N_20827,N_20955);
xor U21057 (N_21057,N_20959,N_20949);
or U21058 (N_21058,N_20998,N_20767);
xor U21059 (N_21059,N_20995,N_20766);
and U21060 (N_21060,N_20975,N_20902);
xnor U21061 (N_21061,N_20835,N_20990);
nor U21062 (N_21062,N_20936,N_20992);
nor U21063 (N_21063,N_20832,N_20843);
and U21064 (N_21064,N_20773,N_20887);
or U21065 (N_21065,N_20828,N_20801);
xor U21066 (N_21066,N_20840,N_20841);
xnor U21067 (N_21067,N_20962,N_20978);
nand U21068 (N_21068,N_20951,N_20991);
nand U21069 (N_21069,N_20794,N_20886);
nand U21070 (N_21070,N_20881,N_20960);
nand U21071 (N_21071,N_20854,N_20811);
xor U21072 (N_21072,N_20804,N_20964);
nand U21073 (N_21073,N_20925,N_20938);
and U21074 (N_21074,N_20896,N_20814);
or U21075 (N_21075,N_20944,N_20981);
nand U21076 (N_21076,N_20953,N_20935);
xnor U21077 (N_21077,N_20884,N_20820);
nor U21078 (N_21078,N_20930,N_20817);
or U21079 (N_21079,N_20844,N_20795);
or U21080 (N_21080,N_20758,N_20890);
xor U21081 (N_21081,N_20918,N_20783);
nand U21082 (N_21082,N_20852,N_20797);
nand U21083 (N_21083,N_20877,N_20880);
and U21084 (N_21084,N_20974,N_20873);
xor U21085 (N_21085,N_20803,N_20868);
and U21086 (N_21086,N_20834,N_20899);
and U21087 (N_21087,N_20768,N_20772);
and U21088 (N_21088,N_20929,N_20864);
and U21089 (N_21089,N_20818,N_20860);
nor U21090 (N_21090,N_20924,N_20963);
xnor U21091 (N_21091,N_20824,N_20858);
nor U21092 (N_21092,N_20849,N_20753);
nand U21093 (N_21093,N_20882,N_20851);
and U21094 (N_21094,N_20985,N_20839);
nor U21095 (N_21095,N_20912,N_20871);
or U21096 (N_21096,N_20915,N_20810);
xnor U21097 (N_21097,N_20954,N_20905);
or U21098 (N_21098,N_20941,N_20986);
or U21099 (N_21099,N_20922,N_20819);
nand U21100 (N_21100,N_20979,N_20754);
nand U21101 (N_21101,N_20825,N_20904);
xor U21102 (N_21102,N_20988,N_20968);
or U21103 (N_21103,N_20807,N_20898);
and U21104 (N_21104,N_20784,N_20770);
nor U21105 (N_21105,N_20889,N_20802);
and U21106 (N_21106,N_20872,N_20894);
or U21107 (N_21107,N_20815,N_20961);
or U21108 (N_21108,N_20809,N_20977);
and U21109 (N_21109,N_20892,N_20782);
xnor U21110 (N_21110,N_20833,N_20853);
nor U21111 (N_21111,N_20857,N_20848);
nand U21112 (N_21112,N_20798,N_20780);
nor U21113 (N_21113,N_20874,N_20799);
xor U21114 (N_21114,N_20923,N_20932);
and U21115 (N_21115,N_20775,N_20752);
xor U21116 (N_21116,N_20901,N_20939);
or U21117 (N_21117,N_20787,N_20761);
nand U21118 (N_21118,N_20965,N_20764);
nor U21119 (N_21119,N_20910,N_20763);
or U21120 (N_21120,N_20790,N_20830);
or U21121 (N_21121,N_20829,N_20771);
xnor U21122 (N_21122,N_20786,N_20970);
xnor U21123 (N_21123,N_20997,N_20989);
or U21124 (N_21124,N_20903,N_20838);
nor U21125 (N_21125,N_20841,N_20995);
nor U21126 (N_21126,N_20861,N_20945);
and U21127 (N_21127,N_20818,N_20977);
or U21128 (N_21128,N_20932,N_20871);
and U21129 (N_21129,N_20769,N_20837);
nor U21130 (N_21130,N_20862,N_20874);
or U21131 (N_21131,N_20945,N_20852);
nand U21132 (N_21132,N_20755,N_20800);
xor U21133 (N_21133,N_20939,N_20864);
and U21134 (N_21134,N_20915,N_20907);
or U21135 (N_21135,N_20965,N_20952);
or U21136 (N_21136,N_20831,N_20889);
or U21137 (N_21137,N_20915,N_20938);
and U21138 (N_21138,N_20810,N_20790);
and U21139 (N_21139,N_20926,N_20803);
nand U21140 (N_21140,N_20986,N_20902);
xor U21141 (N_21141,N_20956,N_20906);
and U21142 (N_21142,N_20990,N_20788);
and U21143 (N_21143,N_20968,N_20867);
nand U21144 (N_21144,N_20948,N_20804);
nor U21145 (N_21145,N_20840,N_20870);
nand U21146 (N_21146,N_20824,N_20855);
nand U21147 (N_21147,N_20927,N_20781);
and U21148 (N_21148,N_20767,N_20872);
and U21149 (N_21149,N_20932,N_20839);
xor U21150 (N_21150,N_20843,N_20809);
or U21151 (N_21151,N_20945,N_20955);
nor U21152 (N_21152,N_20952,N_20889);
or U21153 (N_21153,N_20756,N_20968);
nand U21154 (N_21154,N_20942,N_20866);
nor U21155 (N_21155,N_20946,N_20934);
or U21156 (N_21156,N_20901,N_20753);
xor U21157 (N_21157,N_20877,N_20844);
and U21158 (N_21158,N_20784,N_20793);
or U21159 (N_21159,N_20855,N_20902);
or U21160 (N_21160,N_20856,N_20753);
xor U21161 (N_21161,N_20862,N_20920);
xor U21162 (N_21162,N_20895,N_20906);
nand U21163 (N_21163,N_20932,N_20938);
nor U21164 (N_21164,N_20809,N_20776);
and U21165 (N_21165,N_20888,N_20833);
xnor U21166 (N_21166,N_20882,N_20836);
nand U21167 (N_21167,N_20978,N_20798);
or U21168 (N_21168,N_20984,N_20964);
or U21169 (N_21169,N_20920,N_20919);
nor U21170 (N_21170,N_20867,N_20808);
xor U21171 (N_21171,N_20960,N_20860);
nand U21172 (N_21172,N_20984,N_20994);
and U21173 (N_21173,N_20777,N_20840);
nor U21174 (N_21174,N_20964,N_20997);
nand U21175 (N_21175,N_20835,N_20837);
xnor U21176 (N_21176,N_20882,N_20780);
xor U21177 (N_21177,N_20983,N_20907);
xnor U21178 (N_21178,N_20844,N_20980);
and U21179 (N_21179,N_20860,N_20914);
nand U21180 (N_21180,N_20827,N_20924);
nand U21181 (N_21181,N_20998,N_20756);
nand U21182 (N_21182,N_20893,N_20939);
nor U21183 (N_21183,N_20917,N_20853);
nor U21184 (N_21184,N_20879,N_20950);
nor U21185 (N_21185,N_20888,N_20950);
nor U21186 (N_21186,N_20826,N_20842);
xnor U21187 (N_21187,N_20784,N_20780);
xnor U21188 (N_21188,N_20945,N_20766);
or U21189 (N_21189,N_20896,N_20816);
nor U21190 (N_21190,N_20756,N_20825);
nand U21191 (N_21191,N_20921,N_20840);
and U21192 (N_21192,N_20843,N_20825);
or U21193 (N_21193,N_20770,N_20814);
nor U21194 (N_21194,N_20797,N_20789);
xor U21195 (N_21195,N_20844,N_20763);
xor U21196 (N_21196,N_20834,N_20896);
nand U21197 (N_21197,N_20807,N_20836);
xor U21198 (N_21198,N_20906,N_20858);
nand U21199 (N_21199,N_20846,N_20858);
xor U21200 (N_21200,N_20881,N_20906);
xor U21201 (N_21201,N_20799,N_20934);
and U21202 (N_21202,N_20837,N_20824);
and U21203 (N_21203,N_20969,N_20892);
or U21204 (N_21204,N_20757,N_20982);
xnor U21205 (N_21205,N_20894,N_20898);
and U21206 (N_21206,N_20888,N_20898);
and U21207 (N_21207,N_20809,N_20796);
nor U21208 (N_21208,N_20780,N_20981);
nor U21209 (N_21209,N_20928,N_20933);
and U21210 (N_21210,N_20919,N_20883);
nand U21211 (N_21211,N_20857,N_20927);
and U21212 (N_21212,N_20919,N_20854);
nor U21213 (N_21213,N_20764,N_20859);
xor U21214 (N_21214,N_20962,N_20905);
xnor U21215 (N_21215,N_20780,N_20973);
or U21216 (N_21216,N_20803,N_20992);
nor U21217 (N_21217,N_20864,N_20984);
and U21218 (N_21218,N_20835,N_20997);
or U21219 (N_21219,N_20908,N_20818);
and U21220 (N_21220,N_20834,N_20995);
or U21221 (N_21221,N_20774,N_20813);
nor U21222 (N_21222,N_20859,N_20756);
nand U21223 (N_21223,N_20807,N_20876);
nor U21224 (N_21224,N_20871,N_20929);
and U21225 (N_21225,N_20811,N_20885);
nand U21226 (N_21226,N_20915,N_20953);
and U21227 (N_21227,N_20826,N_20911);
and U21228 (N_21228,N_20913,N_20754);
or U21229 (N_21229,N_20763,N_20843);
nand U21230 (N_21230,N_20775,N_20956);
xnor U21231 (N_21231,N_20965,N_20761);
or U21232 (N_21232,N_20954,N_20993);
nor U21233 (N_21233,N_20923,N_20913);
nand U21234 (N_21234,N_20976,N_20859);
and U21235 (N_21235,N_20862,N_20995);
nand U21236 (N_21236,N_20896,N_20820);
xor U21237 (N_21237,N_20952,N_20831);
or U21238 (N_21238,N_20990,N_20903);
nor U21239 (N_21239,N_20762,N_20939);
or U21240 (N_21240,N_20827,N_20831);
and U21241 (N_21241,N_20823,N_20948);
nand U21242 (N_21242,N_20969,N_20885);
nand U21243 (N_21243,N_20928,N_20870);
xor U21244 (N_21244,N_20871,N_20888);
nand U21245 (N_21245,N_20823,N_20795);
or U21246 (N_21246,N_20905,N_20880);
xnor U21247 (N_21247,N_20947,N_20857);
or U21248 (N_21248,N_20859,N_20800);
nor U21249 (N_21249,N_20950,N_20804);
nor U21250 (N_21250,N_21181,N_21134);
nand U21251 (N_21251,N_21028,N_21137);
or U21252 (N_21252,N_21073,N_21245);
xnor U21253 (N_21253,N_21130,N_21023);
nor U21254 (N_21254,N_21176,N_21201);
nor U21255 (N_21255,N_21125,N_21162);
or U21256 (N_21256,N_21043,N_21032);
nand U21257 (N_21257,N_21042,N_21191);
or U21258 (N_21258,N_21107,N_21129);
or U21259 (N_21259,N_21058,N_21116);
or U21260 (N_21260,N_21157,N_21105);
xnor U21261 (N_21261,N_21206,N_21117);
nor U21262 (N_21262,N_21048,N_21173);
nand U21263 (N_21263,N_21193,N_21056);
nor U21264 (N_21264,N_21188,N_21054);
nand U21265 (N_21265,N_21099,N_21213);
nand U21266 (N_21266,N_21174,N_21161);
xor U21267 (N_21267,N_21217,N_21052);
and U21268 (N_21268,N_21121,N_21092);
or U21269 (N_21269,N_21140,N_21154);
and U21270 (N_21270,N_21138,N_21202);
nand U21271 (N_21271,N_21205,N_21064);
and U21272 (N_21272,N_21085,N_21050);
and U21273 (N_21273,N_21061,N_21172);
and U21274 (N_21274,N_21063,N_21007);
and U21275 (N_21275,N_21127,N_21024);
nor U21276 (N_21276,N_21170,N_21096);
xor U21277 (N_21277,N_21038,N_21102);
nand U21278 (N_21278,N_21242,N_21076);
or U21279 (N_21279,N_21097,N_21207);
xnor U21280 (N_21280,N_21104,N_21029);
nand U21281 (N_21281,N_21214,N_21017);
nand U21282 (N_21282,N_21068,N_21204);
nor U21283 (N_21283,N_21194,N_21031);
and U21284 (N_21284,N_21158,N_21036);
and U21285 (N_21285,N_21080,N_21163);
xor U21286 (N_21286,N_21062,N_21014);
and U21287 (N_21287,N_21227,N_21118);
nand U21288 (N_21288,N_21153,N_21071);
or U21289 (N_21289,N_21215,N_21113);
and U21290 (N_21290,N_21196,N_21133);
and U21291 (N_21291,N_21175,N_21115);
and U21292 (N_21292,N_21082,N_21072);
and U21293 (N_21293,N_21090,N_21112);
and U21294 (N_21294,N_21094,N_21209);
xnor U21295 (N_21295,N_21146,N_21233);
xor U21296 (N_21296,N_21084,N_21069);
and U21297 (N_21297,N_21100,N_21034);
nor U21298 (N_21298,N_21136,N_21103);
and U21299 (N_21299,N_21210,N_21177);
or U21300 (N_21300,N_21087,N_21211);
nor U21301 (N_21301,N_21051,N_21044);
nor U21302 (N_21302,N_21171,N_21225);
and U21303 (N_21303,N_21234,N_21132);
nor U21304 (N_21304,N_21220,N_21030);
and U21305 (N_21305,N_21070,N_21012);
xor U21306 (N_21306,N_21183,N_21186);
nor U21307 (N_21307,N_21095,N_21159);
nand U21308 (N_21308,N_21086,N_21238);
and U21309 (N_21309,N_21222,N_21179);
xor U21310 (N_21310,N_21144,N_21057);
nand U21311 (N_21311,N_21083,N_21147);
or U21312 (N_21312,N_21009,N_21109);
and U21313 (N_21313,N_21018,N_21025);
xor U21314 (N_21314,N_21003,N_21165);
xor U21315 (N_21315,N_21198,N_21046);
nor U21316 (N_21316,N_21218,N_21232);
nand U21317 (N_21317,N_21224,N_21008);
xnor U21318 (N_21318,N_21013,N_21026);
or U21319 (N_21319,N_21192,N_21166);
and U21320 (N_21320,N_21143,N_21216);
xnor U21321 (N_21321,N_21247,N_21195);
or U21322 (N_21322,N_21093,N_21119);
xnor U21323 (N_21323,N_21049,N_21156);
or U21324 (N_21324,N_21122,N_21239);
and U21325 (N_21325,N_21067,N_21244);
nor U21326 (N_21326,N_21190,N_21055);
xnor U21327 (N_21327,N_21019,N_21135);
and U21328 (N_21328,N_21223,N_21237);
xor U21329 (N_21329,N_21221,N_21015);
or U21330 (N_21330,N_21141,N_21005);
nor U21331 (N_21331,N_21088,N_21074);
nand U21332 (N_21332,N_21182,N_21240);
nor U21333 (N_21333,N_21006,N_21059);
nor U21334 (N_21334,N_21001,N_21108);
nand U21335 (N_21335,N_21145,N_21123);
xor U21336 (N_21336,N_21139,N_21155);
and U21337 (N_21337,N_21126,N_21168);
and U21338 (N_21338,N_21066,N_21065);
or U21339 (N_21339,N_21040,N_21151);
and U21340 (N_21340,N_21047,N_21004);
or U21341 (N_21341,N_21178,N_21053);
and U21342 (N_21342,N_21111,N_21000);
or U21343 (N_21343,N_21021,N_21212);
or U21344 (N_21344,N_21185,N_21039);
xor U21345 (N_21345,N_21081,N_21114);
nor U21346 (N_21346,N_21045,N_21219);
xor U21347 (N_21347,N_21152,N_21035);
nor U21348 (N_21348,N_21241,N_21128);
and U21349 (N_21349,N_21164,N_21022);
nor U21350 (N_21350,N_21189,N_21120);
and U21351 (N_21351,N_21101,N_21167);
or U21352 (N_21352,N_21110,N_21089);
or U21353 (N_21353,N_21160,N_21243);
or U21354 (N_21354,N_21020,N_21231);
nand U21355 (N_21355,N_21037,N_21077);
or U21356 (N_21356,N_21197,N_21184);
and U21357 (N_21357,N_21106,N_21149);
xnor U21358 (N_21358,N_21249,N_21248);
nand U21359 (N_21359,N_21228,N_21011);
xor U21360 (N_21360,N_21203,N_21229);
nor U21361 (N_21361,N_21027,N_21002);
nor U21362 (N_21362,N_21010,N_21236);
xor U21363 (N_21363,N_21226,N_21131);
xnor U21364 (N_21364,N_21033,N_21098);
nor U21365 (N_21365,N_21016,N_21079);
xor U21366 (N_21366,N_21150,N_21078);
or U21367 (N_21367,N_21075,N_21230);
and U21368 (N_21368,N_21200,N_21041);
or U21369 (N_21369,N_21124,N_21180);
xor U21370 (N_21370,N_21148,N_21208);
or U21371 (N_21371,N_21169,N_21142);
xnor U21372 (N_21372,N_21091,N_21060);
nor U21373 (N_21373,N_21199,N_21235);
nor U21374 (N_21374,N_21187,N_21246);
and U21375 (N_21375,N_21057,N_21116);
nand U21376 (N_21376,N_21128,N_21163);
nand U21377 (N_21377,N_21195,N_21049);
or U21378 (N_21378,N_21236,N_21247);
xnor U21379 (N_21379,N_21071,N_21058);
and U21380 (N_21380,N_21062,N_21215);
nand U21381 (N_21381,N_21181,N_21175);
or U21382 (N_21382,N_21105,N_21142);
nand U21383 (N_21383,N_21043,N_21053);
or U21384 (N_21384,N_21043,N_21027);
nor U21385 (N_21385,N_21041,N_21030);
xnor U21386 (N_21386,N_21031,N_21071);
and U21387 (N_21387,N_21057,N_21191);
xnor U21388 (N_21388,N_21249,N_21141);
nor U21389 (N_21389,N_21111,N_21153);
nor U21390 (N_21390,N_21022,N_21240);
nand U21391 (N_21391,N_21078,N_21185);
nand U21392 (N_21392,N_21116,N_21034);
xnor U21393 (N_21393,N_21102,N_21152);
xor U21394 (N_21394,N_21073,N_21042);
and U21395 (N_21395,N_21195,N_21189);
xnor U21396 (N_21396,N_21025,N_21108);
or U21397 (N_21397,N_21062,N_21221);
nand U21398 (N_21398,N_21176,N_21225);
and U21399 (N_21399,N_21217,N_21133);
nor U21400 (N_21400,N_21228,N_21133);
or U21401 (N_21401,N_21118,N_21183);
nand U21402 (N_21402,N_21162,N_21170);
or U21403 (N_21403,N_21137,N_21092);
xor U21404 (N_21404,N_21148,N_21036);
nand U21405 (N_21405,N_21013,N_21090);
xnor U21406 (N_21406,N_21007,N_21246);
nor U21407 (N_21407,N_21213,N_21203);
nand U21408 (N_21408,N_21153,N_21124);
or U21409 (N_21409,N_21042,N_21236);
nor U21410 (N_21410,N_21008,N_21240);
nor U21411 (N_21411,N_21083,N_21081);
xnor U21412 (N_21412,N_21226,N_21112);
and U21413 (N_21413,N_21062,N_21245);
nand U21414 (N_21414,N_21009,N_21187);
and U21415 (N_21415,N_21024,N_21093);
nand U21416 (N_21416,N_21223,N_21213);
or U21417 (N_21417,N_21220,N_21097);
nor U21418 (N_21418,N_21171,N_21158);
nor U21419 (N_21419,N_21103,N_21096);
nand U21420 (N_21420,N_21086,N_21180);
and U21421 (N_21421,N_21077,N_21127);
xnor U21422 (N_21422,N_21154,N_21022);
or U21423 (N_21423,N_21040,N_21093);
xnor U21424 (N_21424,N_21194,N_21076);
xor U21425 (N_21425,N_21234,N_21143);
xnor U21426 (N_21426,N_21204,N_21214);
xor U21427 (N_21427,N_21014,N_21004);
or U21428 (N_21428,N_21071,N_21026);
and U21429 (N_21429,N_21122,N_21022);
xor U21430 (N_21430,N_21198,N_21182);
or U21431 (N_21431,N_21117,N_21113);
or U21432 (N_21432,N_21004,N_21128);
xnor U21433 (N_21433,N_21246,N_21059);
and U21434 (N_21434,N_21169,N_21139);
or U21435 (N_21435,N_21026,N_21082);
and U21436 (N_21436,N_21204,N_21185);
nor U21437 (N_21437,N_21088,N_21030);
and U21438 (N_21438,N_21145,N_21125);
nor U21439 (N_21439,N_21054,N_21211);
and U21440 (N_21440,N_21144,N_21113);
nand U21441 (N_21441,N_21141,N_21093);
xnor U21442 (N_21442,N_21076,N_21202);
nand U21443 (N_21443,N_21075,N_21003);
xor U21444 (N_21444,N_21133,N_21158);
xnor U21445 (N_21445,N_21183,N_21088);
xnor U21446 (N_21446,N_21144,N_21051);
nand U21447 (N_21447,N_21170,N_21211);
or U21448 (N_21448,N_21052,N_21070);
or U21449 (N_21449,N_21165,N_21112);
and U21450 (N_21450,N_21221,N_21191);
nand U21451 (N_21451,N_21069,N_21075);
nor U21452 (N_21452,N_21231,N_21194);
and U21453 (N_21453,N_21224,N_21158);
nor U21454 (N_21454,N_21100,N_21031);
xnor U21455 (N_21455,N_21041,N_21149);
nor U21456 (N_21456,N_21094,N_21161);
xnor U21457 (N_21457,N_21068,N_21035);
xor U21458 (N_21458,N_21171,N_21004);
and U21459 (N_21459,N_21176,N_21010);
nor U21460 (N_21460,N_21032,N_21234);
nor U21461 (N_21461,N_21158,N_21240);
nor U21462 (N_21462,N_21046,N_21099);
nor U21463 (N_21463,N_21208,N_21222);
and U21464 (N_21464,N_21049,N_21200);
and U21465 (N_21465,N_21125,N_21161);
nand U21466 (N_21466,N_21237,N_21083);
or U21467 (N_21467,N_21180,N_21126);
nand U21468 (N_21468,N_21033,N_21011);
and U21469 (N_21469,N_21020,N_21071);
xor U21470 (N_21470,N_21124,N_21213);
and U21471 (N_21471,N_21155,N_21046);
nand U21472 (N_21472,N_21202,N_21046);
nand U21473 (N_21473,N_21226,N_21065);
xnor U21474 (N_21474,N_21142,N_21243);
or U21475 (N_21475,N_21009,N_21233);
nor U21476 (N_21476,N_21246,N_21228);
nand U21477 (N_21477,N_21243,N_21066);
xor U21478 (N_21478,N_21032,N_21156);
nand U21479 (N_21479,N_21197,N_21060);
xnor U21480 (N_21480,N_21241,N_21032);
nor U21481 (N_21481,N_21147,N_21112);
and U21482 (N_21482,N_21050,N_21055);
xor U21483 (N_21483,N_21188,N_21094);
or U21484 (N_21484,N_21156,N_21048);
nor U21485 (N_21485,N_21083,N_21158);
nor U21486 (N_21486,N_21089,N_21151);
xor U21487 (N_21487,N_21116,N_21223);
or U21488 (N_21488,N_21186,N_21064);
nor U21489 (N_21489,N_21019,N_21048);
nor U21490 (N_21490,N_21011,N_21078);
and U21491 (N_21491,N_21162,N_21063);
nand U21492 (N_21492,N_21108,N_21237);
and U21493 (N_21493,N_21047,N_21031);
nand U21494 (N_21494,N_21229,N_21018);
nor U21495 (N_21495,N_21133,N_21004);
or U21496 (N_21496,N_21000,N_21019);
or U21497 (N_21497,N_21157,N_21112);
nand U21498 (N_21498,N_21249,N_21116);
and U21499 (N_21499,N_21026,N_21102);
nand U21500 (N_21500,N_21403,N_21318);
nor U21501 (N_21501,N_21341,N_21386);
or U21502 (N_21502,N_21289,N_21335);
nand U21503 (N_21503,N_21405,N_21374);
xnor U21504 (N_21504,N_21266,N_21449);
xor U21505 (N_21505,N_21267,N_21452);
and U21506 (N_21506,N_21316,N_21338);
and U21507 (N_21507,N_21361,N_21344);
and U21508 (N_21508,N_21432,N_21474);
xnor U21509 (N_21509,N_21421,N_21417);
and U21510 (N_21510,N_21489,N_21402);
xor U21511 (N_21511,N_21310,N_21493);
or U21512 (N_21512,N_21290,N_21451);
xnor U21513 (N_21513,N_21298,N_21332);
or U21514 (N_21514,N_21391,N_21360);
nor U21515 (N_21515,N_21381,N_21424);
nand U21516 (N_21516,N_21484,N_21467);
or U21517 (N_21517,N_21321,N_21465);
xnor U21518 (N_21518,N_21477,N_21485);
nor U21519 (N_21519,N_21393,N_21460);
nor U21520 (N_21520,N_21254,N_21384);
or U21521 (N_21521,N_21470,N_21385);
or U21522 (N_21522,N_21416,N_21377);
nor U21523 (N_21523,N_21275,N_21345);
nor U21524 (N_21524,N_21276,N_21435);
and U21525 (N_21525,N_21271,N_21395);
nand U21526 (N_21526,N_21499,N_21328);
or U21527 (N_21527,N_21487,N_21354);
nor U21528 (N_21528,N_21407,N_21413);
xor U21529 (N_21529,N_21269,N_21394);
xnor U21530 (N_21530,N_21359,N_21280);
or U21531 (N_21531,N_21371,N_21346);
nand U21532 (N_21532,N_21491,N_21431);
or U21533 (N_21533,N_21387,N_21414);
nor U21534 (N_21534,N_21426,N_21274);
xnor U21535 (N_21535,N_21370,N_21258);
and U21536 (N_21536,N_21253,N_21320);
nor U21537 (N_21537,N_21392,N_21323);
or U21538 (N_21538,N_21389,N_21488);
xor U21539 (N_21539,N_21494,N_21436);
or U21540 (N_21540,N_21482,N_21270);
or U21541 (N_21541,N_21388,N_21446);
nor U21542 (N_21542,N_21268,N_21262);
nand U21543 (N_21543,N_21342,N_21364);
xor U21544 (N_21544,N_21429,N_21325);
or U21545 (N_21545,N_21376,N_21339);
and U21546 (N_21546,N_21461,N_21422);
nand U21547 (N_21547,N_21322,N_21352);
and U21548 (N_21548,N_21495,N_21336);
nand U21549 (N_21549,N_21383,N_21473);
or U21550 (N_21550,N_21442,N_21273);
xnor U21551 (N_21551,N_21366,N_21418);
nand U21552 (N_21552,N_21445,N_21420);
nand U21553 (N_21553,N_21285,N_21288);
nand U21554 (N_21554,N_21434,N_21411);
and U21555 (N_21555,N_21347,N_21257);
nor U21556 (N_21556,N_21311,N_21369);
or U21557 (N_21557,N_21343,N_21476);
and U21558 (N_21558,N_21443,N_21396);
nand U21559 (N_21559,N_21304,N_21287);
nand U21560 (N_21560,N_21256,N_21313);
xnor U21561 (N_21561,N_21469,N_21471);
nand U21562 (N_21562,N_21462,N_21472);
or U21563 (N_21563,N_21307,N_21357);
and U21564 (N_21564,N_21382,N_21334);
or U21565 (N_21565,N_21264,N_21277);
xnor U21566 (N_21566,N_21265,N_21312);
and U21567 (N_21567,N_21301,N_21375);
xnor U21568 (N_21568,N_21250,N_21358);
or U21569 (N_21569,N_21475,N_21379);
nor U21570 (N_21570,N_21299,N_21331);
xor U21571 (N_21571,N_21279,N_21373);
or U21572 (N_21572,N_21315,N_21433);
or U21573 (N_21573,N_21306,N_21294);
nand U21574 (N_21574,N_21278,N_21464);
nand U21575 (N_21575,N_21309,N_21297);
and U21576 (N_21576,N_21291,N_21439);
or U21577 (N_21577,N_21456,N_21365);
or U21578 (N_21578,N_21261,N_21490);
and U21579 (N_21579,N_21444,N_21355);
xor U21580 (N_21580,N_21367,N_21272);
nor U21581 (N_21581,N_21314,N_21438);
xor U21582 (N_21582,N_21259,N_21459);
or U21583 (N_21583,N_21319,N_21292);
nand U21584 (N_21584,N_21453,N_21255);
and U21585 (N_21585,N_21478,N_21480);
and U21586 (N_21586,N_21425,N_21326);
nor U21587 (N_21587,N_21496,N_21457);
or U21588 (N_21588,N_21455,N_21498);
xnor U21589 (N_21589,N_21308,N_21348);
xnor U21590 (N_21590,N_21430,N_21448);
and U21591 (N_21591,N_21428,N_21305);
or U21592 (N_21592,N_21351,N_21399);
nand U21593 (N_21593,N_21330,N_21380);
or U21594 (N_21594,N_21363,N_21327);
nor U21595 (N_21595,N_21468,N_21440);
nor U21596 (N_21596,N_21437,N_21410);
xnor U21597 (N_21597,N_21412,N_21390);
or U21598 (N_21598,N_21404,N_21295);
xnor U21599 (N_21599,N_21441,N_21362);
nand U21600 (N_21600,N_21281,N_21353);
xor U21601 (N_21601,N_21458,N_21378);
nand U21602 (N_21602,N_21333,N_21401);
xor U21603 (N_21603,N_21400,N_21368);
xor U21604 (N_21604,N_21324,N_21349);
or U21605 (N_21605,N_21481,N_21492);
or U21606 (N_21606,N_21293,N_21397);
or U21607 (N_21607,N_21252,N_21329);
nor U21608 (N_21608,N_21423,N_21447);
nor U21609 (N_21609,N_21409,N_21356);
or U21610 (N_21610,N_21260,N_21450);
xnor U21611 (N_21611,N_21406,N_21282);
and U21612 (N_21612,N_21415,N_21300);
nand U21613 (N_21613,N_21427,N_21263);
nor U21614 (N_21614,N_21283,N_21454);
nand U21615 (N_21615,N_21337,N_21251);
or U21616 (N_21616,N_21303,N_21302);
nand U21617 (N_21617,N_21408,N_21497);
or U21618 (N_21618,N_21479,N_21372);
nand U21619 (N_21619,N_21463,N_21317);
nor U21620 (N_21620,N_21398,N_21483);
nor U21621 (N_21621,N_21296,N_21340);
or U21622 (N_21622,N_21350,N_21419);
and U21623 (N_21623,N_21286,N_21466);
nand U21624 (N_21624,N_21486,N_21284);
or U21625 (N_21625,N_21480,N_21286);
nor U21626 (N_21626,N_21416,N_21307);
or U21627 (N_21627,N_21317,N_21414);
xor U21628 (N_21628,N_21296,N_21431);
and U21629 (N_21629,N_21456,N_21311);
and U21630 (N_21630,N_21346,N_21339);
nand U21631 (N_21631,N_21373,N_21364);
and U21632 (N_21632,N_21391,N_21287);
nor U21633 (N_21633,N_21488,N_21324);
and U21634 (N_21634,N_21377,N_21375);
or U21635 (N_21635,N_21486,N_21360);
nand U21636 (N_21636,N_21270,N_21384);
and U21637 (N_21637,N_21467,N_21497);
nor U21638 (N_21638,N_21260,N_21428);
nand U21639 (N_21639,N_21381,N_21337);
nor U21640 (N_21640,N_21450,N_21374);
and U21641 (N_21641,N_21261,N_21392);
nand U21642 (N_21642,N_21342,N_21430);
xnor U21643 (N_21643,N_21403,N_21324);
xnor U21644 (N_21644,N_21380,N_21378);
nand U21645 (N_21645,N_21433,N_21394);
xnor U21646 (N_21646,N_21402,N_21384);
and U21647 (N_21647,N_21286,N_21490);
nand U21648 (N_21648,N_21469,N_21299);
xor U21649 (N_21649,N_21272,N_21479);
nor U21650 (N_21650,N_21485,N_21424);
nand U21651 (N_21651,N_21420,N_21321);
or U21652 (N_21652,N_21378,N_21471);
xnor U21653 (N_21653,N_21361,N_21373);
or U21654 (N_21654,N_21303,N_21443);
nand U21655 (N_21655,N_21453,N_21311);
xor U21656 (N_21656,N_21350,N_21416);
xnor U21657 (N_21657,N_21376,N_21472);
and U21658 (N_21658,N_21387,N_21403);
and U21659 (N_21659,N_21418,N_21341);
or U21660 (N_21660,N_21296,N_21391);
or U21661 (N_21661,N_21269,N_21302);
nor U21662 (N_21662,N_21333,N_21251);
and U21663 (N_21663,N_21451,N_21487);
or U21664 (N_21664,N_21298,N_21318);
or U21665 (N_21665,N_21444,N_21460);
nand U21666 (N_21666,N_21470,N_21348);
nand U21667 (N_21667,N_21322,N_21448);
and U21668 (N_21668,N_21427,N_21360);
and U21669 (N_21669,N_21356,N_21325);
or U21670 (N_21670,N_21445,N_21261);
nand U21671 (N_21671,N_21489,N_21333);
and U21672 (N_21672,N_21259,N_21490);
nand U21673 (N_21673,N_21455,N_21339);
and U21674 (N_21674,N_21350,N_21391);
and U21675 (N_21675,N_21356,N_21498);
nand U21676 (N_21676,N_21348,N_21399);
and U21677 (N_21677,N_21434,N_21254);
nand U21678 (N_21678,N_21325,N_21444);
nand U21679 (N_21679,N_21396,N_21342);
nand U21680 (N_21680,N_21366,N_21391);
xor U21681 (N_21681,N_21394,N_21499);
or U21682 (N_21682,N_21387,N_21476);
and U21683 (N_21683,N_21466,N_21382);
and U21684 (N_21684,N_21283,N_21314);
and U21685 (N_21685,N_21299,N_21319);
nand U21686 (N_21686,N_21437,N_21462);
or U21687 (N_21687,N_21410,N_21258);
xnor U21688 (N_21688,N_21422,N_21411);
nand U21689 (N_21689,N_21332,N_21329);
xnor U21690 (N_21690,N_21413,N_21259);
or U21691 (N_21691,N_21359,N_21260);
xnor U21692 (N_21692,N_21386,N_21344);
nand U21693 (N_21693,N_21260,N_21342);
and U21694 (N_21694,N_21325,N_21395);
nor U21695 (N_21695,N_21372,N_21444);
or U21696 (N_21696,N_21290,N_21459);
and U21697 (N_21697,N_21381,N_21467);
nor U21698 (N_21698,N_21300,N_21289);
nor U21699 (N_21699,N_21401,N_21313);
nand U21700 (N_21700,N_21411,N_21322);
and U21701 (N_21701,N_21256,N_21263);
and U21702 (N_21702,N_21380,N_21352);
and U21703 (N_21703,N_21423,N_21412);
or U21704 (N_21704,N_21417,N_21389);
nor U21705 (N_21705,N_21285,N_21443);
and U21706 (N_21706,N_21482,N_21369);
and U21707 (N_21707,N_21333,N_21442);
nand U21708 (N_21708,N_21295,N_21496);
nor U21709 (N_21709,N_21346,N_21398);
nor U21710 (N_21710,N_21484,N_21384);
xnor U21711 (N_21711,N_21361,N_21471);
nand U21712 (N_21712,N_21268,N_21277);
nand U21713 (N_21713,N_21332,N_21379);
or U21714 (N_21714,N_21397,N_21491);
and U21715 (N_21715,N_21432,N_21435);
nor U21716 (N_21716,N_21303,N_21384);
nand U21717 (N_21717,N_21260,N_21475);
nor U21718 (N_21718,N_21309,N_21338);
xor U21719 (N_21719,N_21413,N_21460);
and U21720 (N_21720,N_21403,N_21255);
nand U21721 (N_21721,N_21260,N_21285);
nand U21722 (N_21722,N_21432,N_21381);
and U21723 (N_21723,N_21316,N_21435);
or U21724 (N_21724,N_21357,N_21387);
or U21725 (N_21725,N_21427,N_21303);
xnor U21726 (N_21726,N_21444,N_21418);
and U21727 (N_21727,N_21357,N_21282);
nor U21728 (N_21728,N_21257,N_21442);
xor U21729 (N_21729,N_21449,N_21436);
nor U21730 (N_21730,N_21449,N_21301);
or U21731 (N_21731,N_21285,N_21310);
nor U21732 (N_21732,N_21385,N_21456);
nor U21733 (N_21733,N_21311,N_21435);
nand U21734 (N_21734,N_21369,N_21376);
and U21735 (N_21735,N_21276,N_21311);
xnor U21736 (N_21736,N_21280,N_21483);
nand U21737 (N_21737,N_21499,N_21349);
nor U21738 (N_21738,N_21444,N_21485);
or U21739 (N_21739,N_21373,N_21374);
nor U21740 (N_21740,N_21299,N_21416);
and U21741 (N_21741,N_21440,N_21370);
nand U21742 (N_21742,N_21320,N_21312);
or U21743 (N_21743,N_21432,N_21386);
nor U21744 (N_21744,N_21488,N_21270);
or U21745 (N_21745,N_21446,N_21316);
nor U21746 (N_21746,N_21334,N_21289);
xor U21747 (N_21747,N_21454,N_21414);
and U21748 (N_21748,N_21296,N_21318);
and U21749 (N_21749,N_21300,N_21440);
and U21750 (N_21750,N_21580,N_21566);
and U21751 (N_21751,N_21738,N_21749);
or U21752 (N_21752,N_21651,N_21676);
xor U21753 (N_21753,N_21581,N_21590);
nand U21754 (N_21754,N_21511,N_21643);
xor U21755 (N_21755,N_21552,N_21509);
or U21756 (N_21756,N_21512,N_21744);
nand U21757 (N_21757,N_21565,N_21617);
or U21758 (N_21758,N_21538,N_21558);
nand U21759 (N_21759,N_21628,N_21630);
and U21760 (N_21760,N_21573,N_21678);
or U21761 (N_21761,N_21739,N_21632);
nand U21762 (N_21762,N_21626,N_21549);
nor U21763 (N_21763,N_21690,N_21747);
xor U21764 (N_21764,N_21714,N_21505);
and U21765 (N_21765,N_21681,N_21534);
xor U21766 (N_21766,N_21696,N_21555);
and U21767 (N_21767,N_21646,N_21662);
or U21768 (N_21768,N_21671,N_21680);
nand U21769 (N_21769,N_21720,N_21689);
nor U21770 (N_21770,N_21730,N_21703);
or U21771 (N_21771,N_21621,N_21612);
nand U21772 (N_21772,N_21688,N_21645);
xor U21773 (N_21773,N_21515,N_21652);
or U21774 (N_21774,N_21508,N_21530);
nor U21775 (N_21775,N_21639,N_21564);
and U21776 (N_21776,N_21597,N_21571);
nand U21777 (N_21777,N_21705,N_21546);
nand U21778 (N_21778,N_21584,N_21598);
or U21779 (N_21779,N_21582,N_21684);
xnor U21780 (N_21780,N_21721,N_21700);
xnor U21781 (N_21781,N_21735,N_21629);
nand U21782 (N_21782,N_21537,N_21596);
xnor U21783 (N_21783,N_21618,N_21669);
or U21784 (N_21784,N_21586,N_21579);
nor U21785 (N_21785,N_21545,N_21624);
xnor U21786 (N_21786,N_21610,N_21711);
or U21787 (N_21787,N_21550,N_21649);
nand U21788 (N_21788,N_21504,N_21506);
or U21789 (N_21789,N_21620,N_21611);
nor U21790 (N_21790,N_21616,N_21535);
nor U21791 (N_21791,N_21679,N_21575);
or U21792 (N_21792,N_21660,N_21603);
and U21793 (N_21793,N_21593,N_21619);
nor U21794 (N_21794,N_21698,N_21722);
nand U21795 (N_21795,N_21525,N_21729);
or U21796 (N_21796,N_21683,N_21501);
or U21797 (N_21797,N_21604,N_21523);
xor U21798 (N_21798,N_21583,N_21658);
or U21799 (N_21799,N_21595,N_21716);
nand U21800 (N_21800,N_21673,N_21708);
or U21801 (N_21801,N_21636,N_21740);
nand U21802 (N_21802,N_21528,N_21502);
nor U21803 (N_21803,N_21613,N_21702);
nor U21804 (N_21804,N_21541,N_21706);
and U21805 (N_21805,N_21576,N_21642);
nor U21806 (N_21806,N_21561,N_21633);
nand U21807 (N_21807,N_21631,N_21574);
nand U21808 (N_21808,N_21605,N_21713);
xnor U21809 (N_21809,N_21627,N_21514);
or U21810 (N_21810,N_21691,N_21724);
xor U21811 (N_21811,N_21727,N_21615);
xnor U21812 (N_21812,N_21663,N_21726);
nand U21813 (N_21813,N_21507,N_21520);
nor U21814 (N_21814,N_21570,N_21704);
xnor U21815 (N_21815,N_21719,N_21527);
nand U21816 (N_21816,N_21718,N_21622);
nand U21817 (N_21817,N_21606,N_21667);
or U21818 (N_21818,N_21653,N_21589);
nand U21819 (N_21819,N_21614,N_21664);
nor U21820 (N_21820,N_21510,N_21559);
or U21821 (N_21821,N_21602,N_21715);
and U21822 (N_21822,N_21743,N_21567);
nor U21823 (N_21823,N_21563,N_21732);
or U21824 (N_21824,N_21594,N_21682);
nor U21825 (N_21825,N_21547,N_21553);
or U21826 (N_21826,N_21588,N_21542);
nand U21827 (N_21827,N_21518,N_21725);
and U21828 (N_21828,N_21551,N_21522);
xor U21829 (N_21829,N_21585,N_21686);
or U21830 (N_21830,N_21742,N_21647);
xnor U21831 (N_21831,N_21699,N_21513);
xor U21832 (N_21832,N_21635,N_21560);
or U21833 (N_21833,N_21548,N_21674);
and U21834 (N_21834,N_21695,N_21637);
xnor U21835 (N_21835,N_21665,N_21657);
and U21836 (N_21836,N_21634,N_21737);
xnor U21837 (N_21837,N_21685,N_21609);
xor U21838 (N_21838,N_21692,N_21503);
and U21839 (N_21839,N_21531,N_21524);
and U21840 (N_21840,N_21648,N_21638);
nand U21841 (N_21841,N_21517,N_21557);
or U21842 (N_21842,N_21697,N_21672);
nor U21843 (N_21843,N_21693,N_21625);
xor U21844 (N_21844,N_21540,N_21599);
xnor U21845 (N_21845,N_21577,N_21532);
nand U21846 (N_21846,N_21707,N_21650);
xnor U21847 (N_21847,N_21569,N_21723);
or U21848 (N_21848,N_21568,N_21745);
xnor U21849 (N_21849,N_21601,N_21656);
nand U21850 (N_21850,N_21748,N_21500);
nand U21851 (N_21851,N_21668,N_21675);
nand U21852 (N_21852,N_21556,N_21519);
and U21853 (N_21853,N_21701,N_21709);
nor U21854 (N_21854,N_21736,N_21644);
nand U21855 (N_21855,N_21554,N_21572);
or U21856 (N_21856,N_21640,N_21741);
xnor U21857 (N_21857,N_21746,N_21654);
or U21858 (N_21858,N_21687,N_21623);
or U21859 (N_21859,N_21600,N_21731);
nand U21860 (N_21860,N_21670,N_21733);
and U21861 (N_21861,N_21607,N_21544);
nand U21862 (N_21862,N_21734,N_21694);
nand U21863 (N_21863,N_21608,N_21539);
and U21864 (N_21864,N_21728,N_21587);
nor U21865 (N_21865,N_21712,N_21516);
nor U21866 (N_21866,N_21591,N_21592);
nand U21867 (N_21867,N_21543,N_21521);
xnor U21868 (N_21868,N_21536,N_21529);
nor U21869 (N_21869,N_21641,N_21710);
xnor U21870 (N_21870,N_21717,N_21562);
nand U21871 (N_21871,N_21578,N_21533);
nand U21872 (N_21872,N_21661,N_21659);
nand U21873 (N_21873,N_21677,N_21655);
or U21874 (N_21874,N_21666,N_21526);
nor U21875 (N_21875,N_21704,N_21517);
nand U21876 (N_21876,N_21574,N_21626);
nand U21877 (N_21877,N_21603,N_21715);
nand U21878 (N_21878,N_21668,N_21521);
xor U21879 (N_21879,N_21670,N_21524);
and U21880 (N_21880,N_21502,N_21504);
xnor U21881 (N_21881,N_21502,N_21600);
and U21882 (N_21882,N_21667,N_21622);
nor U21883 (N_21883,N_21727,N_21698);
or U21884 (N_21884,N_21651,N_21525);
nor U21885 (N_21885,N_21694,N_21643);
nand U21886 (N_21886,N_21548,N_21646);
and U21887 (N_21887,N_21616,N_21580);
nor U21888 (N_21888,N_21579,N_21540);
nand U21889 (N_21889,N_21504,N_21620);
nor U21890 (N_21890,N_21605,N_21598);
or U21891 (N_21891,N_21609,N_21521);
and U21892 (N_21892,N_21699,N_21619);
xnor U21893 (N_21893,N_21732,N_21630);
or U21894 (N_21894,N_21663,N_21625);
or U21895 (N_21895,N_21698,N_21549);
nand U21896 (N_21896,N_21500,N_21629);
nand U21897 (N_21897,N_21641,N_21513);
and U21898 (N_21898,N_21623,N_21743);
nor U21899 (N_21899,N_21702,N_21739);
nor U21900 (N_21900,N_21613,N_21565);
nand U21901 (N_21901,N_21644,N_21547);
nand U21902 (N_21902,N_21684,N_21650);
nand U21903 (N_21903,N_21696,N_21620);
xnor U21904 (N_21904,N_21643,N_21603);
xor U21905 (N_21905,N_21596,N_21630);
xnor U21906 (N_21906,N_21645,N_21739);
and U21907 (N_21907,N_21535,N_21713);
nor U21908 (N_21908,N_21534,N_21663);
xor U21909 (N_21909,N_21533,N_21706);
nand U21910 (N_21910,N_21565,N_21555);
xor U21911 (N_21911,N_21723,N_21596);
nor U21912 (N_21912,N_21517,N_21620);
and U21913 (N_21913,N_21705,N_21535);
nor U21914 (N_21914,N_21585,N_21529);
xnor U21915 (N_21915,N_21518,N_21731);
nor U21916 (N_21916,N_21674,N_21524);
nor U21917 (N_21917,N_21724,N_21723);
and U21918 (N_21918,N_21555,N_21566);
nor U21919 (N_21919,N_21549,N_21577);
xnor U21920 (N_21920,N_21656,N_21599);
xnor U21921 (N_21921,N_21732,N_21536);
nor U21922 (N_21922,N_21621,N_21539);
nor U21923 (N_21923,N_21726,N_21646);
xor U21924 (N_21924,N_21649,N_21656);
and U21925 (N_21925,N_21716,N_21513);
nor U21926 (N_21926,N_21581,N_21644);
nand U21927 (N_21927,N_21655,N_21742);
and U21928 (N_21928,N_21581,N_21725);
nand U21929 (N_21929,N_21709,N_21534);
or U21930 (N_21930,N_21721,N_21695);
xor U21931 (N_21931,N_21586,N_21673);
nor U21932 (N_21932,N_21617,N_21566);
nor U21933 (N_21933,N_21588,N_21652);
or U21934 (N_21934,N_21721,N_21581);
and U21935 (N_21935,N_21649,N_21596);
or U21936 (N_21936,N_21599,N_21620);
and U21937 (N_21937,N_21658,N_21683);
nand U21938 (N_21938,N_21629,N_21634);
nor U21939 (N_21939,N_21664,N_21508);
and U21940 (N_21940,N_21536,N_21570);
or U21941 (N_21941,N_21706,N_21660);
nor U21942 (N_21942,N_21590,N_21555);
or U21943 (N_21943,N_21652,N_21684);
xor U21944 (N_21944,N_21510,N_21608);
and U21945 (N_21945,N_21619,N_21719);
and U21946 (N_21946,N_21673,N_21554);
xor U21947 (N_21947,N_21519,N_21668);
xor U21948 (N_21948,N_21500,N_21576);
nor U21949 (N_21949,N_21507,N_21640);
or U21950 (N_21950,N_21548,N_21621);
nand U21951 (N_21951,N_21556,N_21646);
and U21952 (N_21952,N_21551,N_21712);
nor U21953 (N_21953,N_21557,N_21704);
xor U21954 (N_21954,N_21672,N_21715);
or U21955 (N_21955,N_21636,N_21700);
xnor U21956 (N_21956,N_21732,N_21522);
xor U21957 (N_21957,N_21631,N_21617);
nand U21958 (N_21958,N_21731,N_21564);
or U21959 (N_21959,N_21554,N_21651);
xnor U21960 (N_21960,N_21743,N_21717);
and U21961 (N_21961,N_21538,N_21516);
nand U21962 (N_21962,N_21526,N_21587);
nand U21963 (N_21963,N_21573,N_21543);
and U21964 (N_21964,N_21560,N_21650);
or U21965 (N_21965,N_21518,N_21686);
nor U21966 (N_21966,N_21587,N_21708);
nor U21967 (N_21967,N_21609,N_21709);
nand U21968 (N_21968,N_21528,N_21556);
nand U21969 (N_21969,N_21509,N_21689);
nor U21970 (N_21970,N_21542,N_21705);
nand U21971 (N_21971,N_21702,N_21639);
nand U21972 (N_21972,N_21513,N_21695);
nor U21973 (N_21973,N_21670,N_21553);
and U21974 (N_21974,N_21521,N_21606);
nand U21975 (N_21975,N_21597,N_21689);
nor U21976 (N_21976,N_21512,N_21687);
nand U21977 (N_21977,N_21715,N_21584);
nand U21978 (N_21978,N_21675,N_21509);
nand U21979 (N_21979,N_21544,N_21519);
and U21980 (N_21980,N_21729,N_21748);
or U21981 (N_21981,N_21574,N_21632);
nor U21982 (N_21982,N_21682,N_21522);
nand U21983 (N_21983,N_21594,N_21726);
xor U21984 (N_21984,N_21676,N_21557);
and U21985 (N_21985,N_21731,N_21670);
xnor U21986 (N_21986,N_21576,N_21542);
and U21987 (N_21987,N_21726,N_21580);
and U21988 (N_21988,N_21648,N_21651);
xnor U21989 (N_21989,N_21749,N_21731);
nand U21990 (N_21990,N_21503,N_21633);
and U21991 (N_21991,N_21542,N_21515);
or U21992 (N_21992,N_21581,N_21660);
and U21993 (N_21993,N_21675,N_21564);
nor U21994 (N_21994,N_21551,N_21552);
xnor U21995 (N_21995,N_21627,N_21710);
nor U21996 (N_21996,N_21734,N_21612);
and U21997 (N_21997,N_21700,N_21681);
nor U21998 (N_21998,N_21624,N_21547);
and U21999 (N_21999,N_21635,N_21738);
and U22000 (N_22000,N_21758,N_21788);
or U22001 (N_22001,N_21874,N_21959);
nor U22002 (N_22002,N_21849,N_21885);
and U22003 (N_22003,N_21873,N_21985);
or U22004 (N_22004,N_21893,N_21976);
or U22005 (N_22005,N_21800,N_21752);
xor U22006 (N_22006,N_21787,N_21770);
nand U22007 (N_22007,N_21848,N_21950);
or U22008 (N_22008,N_21980,N_21986);
or U22009 (N_22009,N_21938,N_21844);
or U22010 (N_22010,N_21915,N_21979);
or U22011 (N_22011,N_21780,N_21819);
nand U22012 (N_22012,N_21762,N_21997);
xor U22013 (N_22013,N_21835,N_21771);
nand U22014 (N_22014,N_21984,N_21899);
and U22015 (N_22015,N_21811,N_21930);
and U22016 (N_22016,N_21908,N_21853);
nor U22017 (N_22017,N_21785,N_21756);
nand U22018 (N_22018,N_21881,N_21989);
nand U22019 (N_22019,N_21822,N_21939);
and U22020 (N_22020,N_21929,N_21907);
or U22021 (N_22021,N_21883,N_21827);
and U22022 (N_22022,N_21942,N_21951);
nand U22023 (N_22023,N_21875,N_21944);
xnor U22024 (N_22024,N_21920,N_21936);
and U22025 (N_22025,N_21775,N_21839);
nor U22026 (N_22026,N_21921,N_21791);
nand U22027 (N_22027,N_21948,N_21768);
nor U22028 (N_22028,N_21766,N_21841);
xor U22029 (N_22029,N_21851,N_21918);
and U22030 (N_22030,N_21896,N_21796);
xor U22031 (N_22031,N_21911,N_21926);
or U22032 (N_22032,N_21868,N_21957);
xor U22033 (N_22033,N_21812,N_21760);
xnor U22034 (N_22034,N_21751,N_21990);
xor U22035 (N_22035,N_21808,N_21803);
nor U22036 (N_22036,N_21809,N_21952);
nand U22037 (N_22037,N_21922,N_21772);
and U22038 (N_22038,N_21838,N_21993);
and U22039 (N_22039,N_21886,N_21904);
nand U22040 (N_22040,N_21978,N_21933);
nor U22041 (N_22041,N_21784,N_21935);
and U22042 (N_22042,N_21917,N_21887);
nor U22043 (N_22043,N_21974,N_21840);
or U22044 (N_22044,N_21842,N_21831);
nand U22045 (N_22045,N_21925,N_21971);
nand U22046 (N_22046,N_21913,N_21807);
or U22047 (N_22047,N_21818,N_21958);
nor U22048 (N_22048,N_21755,N_21916);
xor U22049 (N_22049,N_21854,N_21963);
and U22050 (N_22050,N_21850,N_21778);
nor U22051 (N_22051,N_21816,N_21995);
or U22052 (N_22052,N_21906,N_21824);
nor U22053 (N_22053,N_21802,N_21956);
nand U22054 (N_22054,N_21937,N_21829);
and U22055 (N_22055,N_21955,N_21817);
nand U22056 (N_22056,N_21799,N_21765);
nand U22057 (N_22057,N_21894,N_21863);
nor U22058 (N_22058,N_21970,N_21813);
or U22059 (N_22059,N_21864,N_21859);
xor U22060 (N_22060,N_21814,N_21776);
nor U22061 (N_22061,N_21972,N_21769);
nand U22062 (N_22062,N_21794,N_21783);
nor U22063 (N_22063,N_21833,N_21781);
nor U22064 (N_22064,N_21805,N_21876);
xor U22065 (N_22065,N_21763,N_21890);
xnor U22066 (N_22066,N_21919,N_21999);
or U22067 (N_22067,N_21882,N_21941);
nor U22068 (N_22068,N_21949,N_21815);
nor U22069 (N_22069,N_21973,N_21786);
and U22070 (N_22070,N_21947,N_21880);
or U22071 (N_22071,N_21836,N_21975);
xor U22072 (N_22072,N_21759,N_21982);
and U22073 (N_22073,N_21996,N_21845);
or U22074 (N_22074,N_21945,N_21891);
and U22075 (N_22075,N_21750,N_21968);
and U22076 (N_22076,N_21923,N_21782);
xor U22077 (N_22077,N_21792,N_21810);
nand U22078 (N_22078,N_21773,N_21825);
nor U22079 (N_22079,N_21869,N_21820);
and U22080 (N_22080,N_21753,N_21994);
nand U22081 (N_22081,N_21927,N_21924);
nor U22082 (N_22082,N_21892,N_21878);
nand U22083 (N_22083,N_21910,N_21761);
or U22084 (N_22084,N_21983,N_21914);
xor U22085 (N_22085,N_21867,N_21877);
or U22086 (N_22086,N_21879,N_21858);
and U22087 (N_22087,N_21795,N_21832);
xnor U22088 (N_22088,N_21789,N_21754);
and U22089 (N_22089,N_21898,N_21888);
xnor U22090 (N_22090,N_21856,N_21837);
xnor U22091 (N_22091,N_21900,N_21862);
or U22092 (N_22092,N_21987,N_21871);
nor U22093 (N_22093,N_21857,N_21866);
nor U22094 (N_22094,N_21932,N_21793);
nor U22095 (N_22095,N_21826,N_21909);
and U22096 (N_22096,N_21889,N_21798);
nor U22097 (N_22097,N_21774,N_21847);
and U22098 (N_22098,N_21855,N_21846);
xnor U22099 (N_22099,N_21884,N_21903);
or U22100 (N_22100,N_21860,N_21905);
or U22101 (N_22101,N_21821,N_21830);
nand U22102 (N_22102,N_21967,N_21895);
nand U22103 (N_22103,N_21801,N_21964);
nor U22104 (N_22104,N_21953,N_21764);
and U22105 (N_22105,N_21961,N_21954);
or U22106 (N_22106,N_21897,N_21998);
nand U22107 (N_22107,N_21931,N_21977);
nor U22108 (N_22108,N_21843,N_21872);
xor U22109 (N_22109,N_21861,N_21767);
or U22110 (N_22110,N_21902,N_21777);
and U22111 (N_22111,N_21828,N_21988);
and U22112 (N_22112,N_21934,N_21966);
xnor U22113 (N_22113,N_21823,N_21852);
nand U22114 (N_22114,N_21806,N_21946);
nand U22115 (N_22115,N_21940,N_21804);
and U22116 (N_22116,N_21870,N_21960);
xor U22117 (N_22117,N_21962,N_21969);
and U22118 (N_22118,N_21943,N_21757);
and U22119 (N_22119,N_21865,N_21797);
xnor U22120 (N_22120,N_21965,N_21790);
and U22121 (N_22121,N_21991,N_21912);
xor U22122 (N_22122,N_21981,N_21992);
or U22123 (N_22123,N_21901,N_21779);
nand U22124 (N_22124,N_21928,N_21834);
or U22125 (N_22125,N_21789,N_21825);
and U22126 (N_22126,N_21975,N_21995);
xor U22127 (N_22127,N_21918,N_21949);
or U22128 (N_22128,N_21923,N_21797);
and U22129 (N_22129,N_21963,N_21908);
and U22130 (N_22130,N_21761,N_21785);
xor U22131 (N_22131,N_21813,N_21783);
nand U22132 (N_22132,N_21840,N_21946);
nand U22133 (N_22133,N_21968,N_21905);
nand U22134 (N_22134,N_21844,N_21794);
nor U22135 (N_22135,N_21762,N_21974);
or U22136 (N_22136,N_21869,N_21823);
nor U22137 (N_22137,N_21850,N_21821);
nand U22138 (N_22138,N_21965,N_21919);
or U22139 (N_22139,N_21791,N_21889);
xor U22140 (N_22140,N_21769,N_21931);
or U22141 (N_22141,N_21895,N_21783);
or U22142 (N_22142,N_21754,N_21935);
xnor U22143 (N_22143,N_21987,N_21806);
xnor U22144 (N_22144,N_21907,N_21752);
or U22145 (N_22145,N_21752,N_21912);
nand U22146 (N_22146,N_21795,N_21972);
nand U22147 (N_22147,N_21810,N_21907);
xnor U22148 (N_22148,N_21798,N_21922);
nand U22149 (N_22149,N_21860,N_21974);
nor U22150 (N_22150,N_21782,N_21919);
nor U22151 (N_22151,N_21929,N_21834);
and U22152 (N_22152,N_21790,N_21787);
nor U22153 (N_22153,N_21883,N_21965);
and U22154 (N_22154,N_21786,N_21836);
xor U22155 (N_22155,N_21753,N_21953);
or U22156 (N_22156,N_21941,N_21808);
nor U22157 (N_22157,N_21890,N_21806);
nor U22158 (N_22158,N_21764,N_21924);
nor U22159 (N_22159,N_21958,N_21809);
or U22160 (N_22160,N_21902,N_21839);
xnor U22161 (N_22161,N_21974,N_21956);
or U22162 (N_22162,N_21820,N_21889);
or U22163 (N_22163,N_21881,N_21868);
xnor U22164 (N_22164,N_21914,N_21856);
or U22165 (N_22165,N_21877,N_21940);
xnor U22166 (N_22166,N_21841,N_21895);
and U22167 (N_22167,N_21800,N_21938);
nand U22168 (N_22168,N_21784,N_21754);
or U22169 (N_22169,N_21939,N_21955);
or U22170 (N_22170,N_21967,N_21909);
xnor U22171 (N_22171,N_21963,N_21965);
xor U22172 (N_22172,N_21842,N_21799);
or U22173 (N_22173,N_21892,N_21833);
nand U22174 (N_22174,N_21921,N_21974);
xnor U22175 (N_22175,N_21789,N_21782);
or U22176 (N_22176,N_21954,N_21861);
or U22177 (N_22177,N_21773,N_21765);
nand U22178 (N_22178,N_21759,N_21902);
nor U22179 (N_22179,N_21930,N_21766);
xor U22180 (N_22180,N_21864,N_21908);
xnor U22181 (N_22181,N_21785,N_21967);
or U22182 (N_22182,N_21978,N_21904);
xnor U22183 (N_22183,N_21977,N_21776);
nand U22184 (N_22184,N_21789,N_21978);
or U22185 (N_22185,N_21875,N_21809);
nor U22186 (N_22186,N_21759,N_21961);
nor U22187 (N_22187,N_21869,N_21871);
nand U22188 (N_22188,N_21816,N_21751);
or U22189 (N_22189,N_21946,N_21829);
nand U22190 (N_22190,N_21840,N_21950);
nand U22191 (N_22191,N_21783,N_21785);
nand U22192 (N_22192,N_21837,N_21840);
or U22193 (N_22193,N_21940,N_21821);
xnor U22194 (N_22194,N_21844,N_21887);
nor U22195 (N_22195,N_21798,N_21910);
xnor U22196 (N_22196,N_21950,N_21779);
nor U22197 (N_22197,N_21852,N_21993);
nor U22198 (N_22198,N_21880,N_21851);
nand U22199 (N_22199,N_21889,N_21990);
nor U22200 (N_22200,N_21756,N_21784);
and U22201 (N_22201,N_21976,N_21771);
xor U22202 (N_22202,N_21873,N_21815);
xor U22203 (N_22203,N_21922,N_21943);
xnor U22204 (N_22204,N_21872,N_21976);
or U22205 (N_22205,N_21888,N_21823);
or U22206 (N_22206,N_21870,N_21769);
xor U22207 (N_22207,N_21868,N_21942);
xnor U22208 (N_22208,N_21763,N_21804);
and U22209 (N_22209,N_21756,N_21820);
nor U22210 (N_22210,N_21879,N_21999);
nor U22211 (N_22211,N_21829,N_21870);
xor U22212 (N_22212,N_21964,N_21946);
nand U22213 (N_22213,N_21819,N_21905);
nand U22214 (N_22214,N_21874,N_21894);
and U22215 (N_22215,N_21929,N_21769);
nand U22216 (N_22216,N_21838,N_21981);
nor U22217 (N_22217,N_21880,N_21930);
and U22218 (N_22218,N_21997,N_21889);
or U22219 (N_22219,N_21917,N_21888);
or U22220 (N_22220,N_21853,N_21772);
xor U22221 (N_22221,N_21915,N_21989);
or U22222 (N_22222,N_21951,N_21750);
and U22223 (N_22223,N_21809,N_21997);
xnor U22224 (N_22224,N_21787,N_21779);
or U22225 (N_22225,N_21889,N_21831);
nand U22226 (N_22226,N_21889,N_21882);
or U22227 (N_22227,N_21871,N_21960);
nor U22228 (N_22228,N_21789,N_21955);
nand U22229 (N_22229,N_21798,N_21758);
or U22230 (N_22230,N_21780,N_21979);
or U22231 (N_22231,N_21971,N_21908);
or U22232 (N_22232,N_21950,N_21895);
nor U22233 (N_22233,N_21792,N_21801);
or U22234 (N_22234,N_21880,N_21835);
xor U22235 (N_22235,N_21897,N_21991);
xor U22236 (N_22236,N_21903,N_21986);
xor U22237 (N_22237,N_21917,N_21802);
nor U22238 (N_22238,N_21891,N_21973);
xnor U22239 (N_22239,N_21885,N_21990);
nor U22240 (N_22240,N_21931,N_21879);
or U22241 (N_22241,N_21775,N_21773);
and U22242 (N_22242,N_21792,N_21789);
nand U22243 (N_22243,N_21923,N_21750);
nand U22244 (N_22244,N_21839,N_21999);
and U22245 (N_22245,N_21760,N_21884);
xor U22246 (N_22246,N_21779,N_21977);
nor U22247 (N_22247,N_21978,N_21990);
and U22248 (N_22248,N_21973,N_21845);
xor U22249 (N_22249,N_21908,N_21992);
or U22250 (N_22250,N_22067,N_22064);
or U22251 (N_22251,N_22076,N_22068);
nand U22252 (N_22252,N_22165,N_22005);
xnor U22253 (N_22253,N_22231,N_22078);
or U22254 (N_22254,N_22109,N_22048);
nor U22255 (N_22255,N_22200,N_22233);
nand U22256 (N_22256,N_22188,N_22060);
and U22257 (N_22257,N_22139,N_22190);
or U22258 (N_22258,N_22083,N_22069);
nor U22259 (N_22259,N_22106,N_22239);
nor U22260 (N_22260,N_22079,N_22040);
nor U22261 (N_22261,N_22086,N_22147);
xor U22262 (N_22262,N_22043,N_22001);
or U22263 (N_22263,N_22010,N_22141);
nor U22264 (N_22264,N_22240,N_22159);
or U22265 (N_22265,N_22196,N_22038);
xnor U22266 (N_22266,N_22032,N_22114);
nor U22267 (N_22267,N_22130,N_22119);
xor U22268 (N_22268,N_22183,N_22166);
nor U22269 (N_22269,N_22126,N_22046);
and U22270 (N_22270,N_22207,N_22238);
nor U22271 (N_22271,N_22004,N_22047);
and U22272 (N_22272,N_22018,N_22158);
and U22273 (N_22273,N_22085,N_22042);
xnor U22274 (N_22274,N_22015,N_22181);
and U22275 (N_22275,N_22101,N_22153);
or U22276 (N_22276,N_22073,N_22011);
or U22277 (N_22277,N_22104,N_22054);
nand U22278 (N_22278,N_22112,N_22089);
nor U22279 (N_22279,N_22071,N_22057);
or U22280 (N_22280,N_22187,N_22221);
xnor U22281 (N_22281,N_22195,N_22063);
xnor U22282 (N_22282,N_22031,N_22092);
xor U22283 (N_22283,N_22102,N_22197);
nand U22284 (N_22284,N_22023,N_22125);
or U22285 (N_22285,N_22027,N_22097);
nand U22286 (N_22286,N_22241,N_22167);
or U22287 (N_22287,N_22058,N_22222);
nor U22288 (N_22288,N_22172,N_22148);
nand U22289 (N_22289,N_22155,N_22151);
xnor U22290 (N_22290,N_22045,N_22194);
xnor U22291 (N_22291,N_22229,N_22163);
or U22292 (N_22292,N_22029,N_22100);
xnor U22293 (N_22293,N_22162,N_22033);
xor U22294 (N_22294,N_22227,N_22072);
xor U22295 (N_22295,N_22140,N_22108);
and U22296 (N_22296,N_22247,N_22120);
and U22297 (N_22297,N_22050,N_22093);
nand U22298 (N_22298,N_22211,N_22127);
xnor U22299 (N_22299,N_22156,N_22087);
xnor U22300 (N_22300,N_22145,N_22210);
nand U22301 (N_22301,N_22180,N_22149);
or U22302 (N_22302,N_22124,N_22173);
nor U22303 (N_22303,N_22075,N_22061);
nor U22304 (N_22304,N_22003,N_22184);
or U22305 (N_22305,N_22041,N_22123);
nand U22306 (N_22306,N_22174,N_22036);
or U22307 (N_22307,N_22117,N_22094);
and U22308 (N_22308,N_22113,N_22204);
nor U22309 (N_22309,N_22170,N_22037);
nand U22310 (N_22310,N_22171,N_22202);
nor U22311 (N_22311,N_22066,N_22230);
nand U22312 (N_22312,N_22154,N_22129);
nand U22313 (N_22313,N_22177,N_22020);
and U22314 (N_22314,N_22216,N_22193);
nor U22315 (N_22315,N_22228,N_22199);
and U22316 (N_22316,N_22122,N_22215);
and U22317 (N_22317,N_22059,N_22235);
xnor U22318 (N_22318,N_22107,N_22098);
xor U22319 (N_22319,N_22135,N_22191);
xnor U22320 (N_22320,N_22164,N_22161);
or U22321 (N_22321,N_22056,N_22065);
nand U22322 (N_22322,N_22143,N_22179);
and U22323 (N_22323,N_22115,N_22116);
nand U22324 (N_22324,N_22030,N_22000);
nor U22325 (N_22325,N_22213,N_22133);
nor U22326 (N_22326,N_22185,N_22077);
or U22327 (N_22327,N_22160,N_22223);
xnor U22328 (N_22328,N_22219,N_22009);
nand U22329 (N_22329,N_22248,N_22225);
or U22330 (N_22330,N_22090,N_22017);
nor U22331 (N_22331,N_22246,N_22035);
nor U22332 (N_22332,N_22105,N_22039);
nand U22333 (N_22333,N_22111,N_22157);
or U22334 (N_22334,N_22176,N_22152);
nor U22335 (N_22335,N_22084,N_22236);
xnor U22336 (N_22336,N_22091,N_22007);
or U22337 (N_22337,N_22082,N_22245);
and U22338 (N_22338,N_22146,N_22062);
and U22339 (N_22339,N_22206,N_22074);
xor U22340 (N_22340,N_22209,N_22237);
nor U22341 (N_22341,N_22178,N_22019);
and U22342 (N_22342,N_22044,N_22096);
or U22343 (N_22343,N_22034,N_22186);
xnor U22344 (N_22344,N_22232,N_22220);
and U22345 (N_22345,N_22242,N_22224);
and U22346 (N_22346,N_22006,N_22203);
or U22347 (N_22347,N_22080,N_22137);
nand U22348 (N_22348,N_22051,N_22189);
or U22349 (N_22349,N_22144,N_22168);
and U22350 (N_22350,N_22055,N_22021);
and U22351 (N_22351,N_22169,N_22024);
nand U22352 (N_22352,N_22138,N_22192);
and U22353 (N_22353,N_22244,N_22198);
nor U22354 (N_22354,N_22088,N_22014);
nand U22355 (N_22355,N_22012,N_22110);
or U22356 (N_22356,N_22128,N_22212);
nand U22357 (N_22357,N_22226,N_22218);
and U22358 (N_22358,N_22201,N_22208);
xor U22359 (N_22359,N_22131,N_22026);
nand U22360 (N_22360,N_22142,N_22175);
and U22361 (N_22361,N_22070,N_22013);
nor U22362 (N_22362,N_22118,N_22234);
and U22363 (N_22363,N_22205,N_22099);
and U22364 (N_22364,N_22134,N_22121);
nand U22365 (N_22365,N_22103,N_22132);
nor U22366 (N_22366,N_22053,N_22217);
nor U22367 (N_22367,N_22081,N_22150);
nor U22368 (N_22368,N_22025,N_22052);
nor U22369 (N_22369,N_22028,N_22002);
or U22370 (N_22370,N_22016,N_22249);
and U22371 (N_22371,N_22095,N_22008);
nor U22372 (N_22372,N_22136,N_22049);
or U22373 (N_22373,N_22243,N_22182);
xor U22374 (N_22374,N_22214,N_22022);
nor U22375 (N_22375,N_22176,N_22122);
or U22376 (N_22376,N_22243,N_22044);
xor U22377 (N_22377,N_22178,N_22064);
xor U22378 (N_22378,N_22054,N_22130);
xor U22379 (N_22379,N_22232,N_22238);
xor U22380 (N_22380,N_22226,N_22141);
or U22381 (N_22381,N_22071,N_22011);
and U22382 (N_22382,N_22184,N_22084);
xnor U22383 (N_22383,N_22101,N_22155);
and U22384 (N_22384,N_22082,N_22040);
and U22385 (N_22385,N_22124,N_22109);
xor U22386 (N_22386,N_22238,N_22161);
nor U22387 (N_22387,N_22156,N_22021);
or U22388 (N_22388,N_22134,N_22169);
nand U22389 (N_22389,N_22149,N_22231);
and U22390 (N_22390,N_22053,N_22071);
xnor U22391 (N_22391,N_22021,N_22050);
xor U22392 (N_22392,N_22149,N_22119);
and U22393 (N_22393,N_22200,N_22095);
or U22394 (N_22394,N_22240,N_22085);
and U22395 (N_22395,N_22064,N_22145);
or U22396 (N_22396,N_22026,N_22159);
and U22397 (N_22397,N_22175,N_22188);
or U22398 (N_22398,N_22069,N_22062);
and U22399 (N_22399,N_22188,N_22215);
xor U22400 (N_22400,N_22219,N_22189);
nor U22401 (N_22401,N_22218,N_22112);
xor U22402 (N_22402,N_22248,N_22240);
nor U22403 (N_22403,N_22240,N_22220);
and U22404 (N_22404,N_22233,N_22171);
and U22405 (N_22405,N_22235,N_22157);
nand U22406 (N_22406,N_22106,N_22043);
nand U22407 (N_22407,N_22128,N_22160);
nor U22408 (N_22408,N_22236,N_22168);
or U22409 (N_22409,N_22122,N_22071);
or U22410 (N_22410,N_22246,N_22241);
or U22411 (N_22411,N_22123,N_22247);
nand U22412 (N_22412,N_22054,N_22155);
xnor U22413 (N_22413,N_22246,N_22195);
xor U22414 (N_22414,N_22147,N_22039);
or U22415 (N_22415,N_22176,N_22154);
xnor U22416 (N_22416,N_22225,N_22062);
nor U22417 (N_22417,N_22178,N_22197);
and U22418 (N_22418,N_22070,N_22211);
or U22419 (N_22419,N_22234,N_22159);
nand U22420 (N_22420,N_22157,N_22228);
nand U22421 (N_22421,N_22103,N_22163);
and U22422 (N_22422,N_22216,N_22016);
and U22423 (N_22423,N_22224,N_22219);
nand U22424 (N_22424,N_22126,N_22079);
nor U22425 (N_22425,N_22113,N_22065);
nor U22426 (N_22426,N_22001,N_22212);
nand U22427 (N_22427,N_22045,N_22086);
xnor U22428 (N_22428,N_22133,N_22115);
and U22429 (N_22429,N_22050,N_22026);
nand U22430 (N_22430,N_22057,N_22087);
or U22431 (N_22431,N_22003,N_22138);
nor U22432 (N_22432,N_22179,N_22224);
nor U22433 (N_22433,N_22094,N_22106);
nand U22434 (N_22434,N_22133,N_22055);
and U22435 (N_22435,N_22125,N_22117);
xnor U22436 (N_22436,N_22176,N_22173);
xnor U22437 (N_22437,N_22041,N_22177);
and U22438 (N_22438,N_22101,N_22112);
xnor U22439 (N_22439,N_22070,N_22223);
or U22440 (N_22440,N_22061,N_22066);
nor U22441 (N_22441,N_22244,N_22169);
nand U22442 (N_22442,N_22061,N_22039);
nand U22443 (N_22443,N_22099,N_22197);
or U22444 (N_22444,N_22144,N_22063);
nand U22445 (N_22445,N_22108,N_22109);
or U22446 (N_22446,N_22008,N_22110);
and U22447 (N_22447,N_22175,N_22065);
and U22448 (N_22448,N_22157,N_22205);
and U22449 (N_22449,N_22060,N_22231);
nand U22450 (N_22450,N_22245,N_22081);
and U22451 (N_22451,N_22005,N_22096);
nand U22452 (N_22452,N_22166,N_22067);
and U22453 (N_22453,N_22048,N_22030);
xor U22454 (N_22454,N_22124,N_22245);
xnor U22455 (N_22455,N_22175,N_22011);
or U22456 (N_22456,N_22155,N_22078);
or U22457 (N_22457,N_22064,N_22195);
xnor U22458 (N_22458,N_22172,N_22072);
and U22459 (N_22459,N_22107,N_22093);
and U22460 (N_22460,N_22160,N_22134);
and U22461 (N_22461,N_22111,N_22203);
and U22462 (N_22462,N_22234,N_22122);
and U22463 (N_22463,N_22232,N_22010);
nand U22464 (N_22464,N_22138,N_22077);
nand U22465 (N_22465,N_22230,N_22205);
nand U22466 (N_22466,N_22014,N_22094);
xnor U22467 (N_22467,N_22106,N_22219);
nand U22468 (N_22468,N_22121,N_22103);
nand U22469 (N_22469,N_22069,N_22052);
xnor U22470 (N_22470,N_22237,N_22086);
or U22471 (N_22471,N_22148,N_22185);
and U22472 (N_22472,N_22100,N_22136);
xor U22473 (N_22473,N_22045,N_22229);
xor U22474 (N_22474,N_22027,N_22180);
and U22475 (N_22475,N_22069,N_22110);
nor U22476 (N_22476,N_22112,N_22096);
xnor U22477 (N_22477,N_22168,N_22143);
nand U22478 (N_22478,N_22005,N_22012);
and U22479 (N_22479,N_22153,N_22181);
xor U22480 (N_22480,N_22032,N_22172);
nand U22481 (N_22481,N_22019,N_22240);
nand U22482 (N_22482,N_22123,N_22174);
xnor U22483 (N_22483,N_22138,N_22107);
xnor U22484 (N_22484,N_22037,N_22122);
nand U22485 (N_22485,N_22075,N_22214);
nand U22486 (N_22486,N_22227,N_22057);
nor U22487 (N_22487,N_22225,N_22246);
xnor U22488 (N_22488,N_22080,N_22174);
nor U22489 (N_22489,N_22154,N_22020);
xor U22490 (N_22490,N_22072,N_22104);
nand U22491 (N_22491,N_22093,N_22196);
or U22492 (N_22492,N_22176,N_22042);
nand U22493 (N_22493,N_22227,N_22130);
or U22494 (N_22494,N_22002,N_22238);
and U22495 (N_22495,N_22121,N_22139);
nor U22496 (N_22496,N_22188,N_22062);
or U22497 (N_22497,N_22029,N_22235);
and U22498 (N_22498,N_22000,N_22005);
xor U22499 (N_22499,N_22086,N_22124);
and U22500 (N_22500,N_22496,N_22495);
and U22501 (N_22501,N_22494,N_22308);
or U22502 (N_22502,N_22417,N_22284);
nor U22503 (N_22503,N_22302,N_22359);
and U22504 (N_22504,N_22362,N_22320);
nand U22505 (N_22505,N_22263,N_22366);
nor U22506 (N_22506,N_22381,N_22271);
and U22507 (N_22507,N_22399,N_22497);
and U22508 (N_22508,N_22352,N_22253);
nor U22509 (N_22509,N_22457,N_22478);
nand U22510 (N_22510,N_22305,N_22294);
nor U22511 (N_22511,N_22347,N_22374);
nor U22512 (N_22512,N_22467,N_22350);
nor U22513 (N_22513,N_22491,N_22436);
and U22514 (N_22514,N_22346,N_22461);
or U22515 (N_22515,N_22397,N_22490);
or U22516 (N_22516,N_22485,N_22469);
or U22517 (N_22517,N_22298,N_22369);
or U22518 (N_22518,N_22419,N_22272);
and U22519 (N_22519,N_22270,N_22325);
nor U22520 (N_22520,N_22439,N_22438);
nand U22521 (N_22521,N_22285,N_22288);
or U22522 (N_22522,N_22363,N_22408);
nand U22523 (N_22523,N_22473,N_22327);
nand U22524 (N_22524,N_22411,N_22306);
nor U22525 (N_22525,N_22442,N_22372);
nor U22526 (N_22526,N_22474,N_22416);
and U22527 (N_22527,N_22317,N_22268);
and U22528 (N_22528,N_22315,N_22480);
xnor U22529 (N_22529,N_22384,N_22475);
nand U22530 (N_22530,N_22289,N_22486);
or U22531 (N_22531,N_22477,N_22356);
or U22532 (N_22532,N_22336,N_22345);
nor U22533 (N_22533,N_22349,N_22394);
nand U22534 (N_22534,N_22286,N_22357);
or U22535 (N_22535,N_22387,N_22261);
nand U22536 (N_22536,N_22487,N_22358);
nand U22537 (N_22537,N_22407,N_22489);
nand U22538 (N_22538,N_22251,N_22333);
nor U22539 (N_22539,N_22360,N_22388);
xnor U22540 (N_22540,N_22367,N_22254);
nor U22541 (N_22541,N_22418,N_22390);
or U22542 (N_22542,N_22328,N_22392);
and U22543 (N_22543,N_22344,N_22331);
or U22544 (N_22544,N_22319,N_22312);
or U22545 (N_22545,N_22450,N_22282);
xnor U22546 (N_22546,N_22299,N_22444);
nand U22547 (N_22547,N_22403,N_22414);
or U22548 (N_22548,N_22383,N_22313);
or U22549 (N_22549,N_22323,N_22413);
nor U22550 (N_22550,N_22437,N_22452);
and U22551 (N_22551,N_22318,N_22409);
nand U22552 (N_22552,N_22269,N_22425);
nor U22553 (N_22553,N_22458,N_22273);
and U22554 (N_22554,N_22396,N_22440);
nor U22555 (N_22555,N_22295,N_22342);
nand U22556 (N_22556,N_22348,N_22443);
or U22557 (N_22557,N_22355,N_22258);
and U22558 (N_22558,N_22321,N_22470);
and U22559 (N_22559,N_22351,N_22262);
and U22560 (N_22560,N_22446,N_22279);
nand U22561 (N_22561,N_22329,N_22424);
nand U22562 (N_22562,N_22370,N_22364);
or U22563 (N_22563,N_22277,N_22304);
xor U22564 (N_22564,N_22296,N_22483);
nor U22565 (N_22565,N_22493,N_22426);
nand U22566 (N_22566,N_22307,N_22481);
or U22567 (N_22567,N_22423,N_22451);
xnor U22568 (N_22568,N_22265,N_22453);
xor U22569 (N_22569,N_22311,N_22400);
and U22570 (N_22570,N_22448,N_22391);
nor U22571 (N_22571,N_22267,N_22441);
nor U22572 (N_22572,N_22472,N_22338);
nand U22573 (N_22573,N_22429,N_22379);
xor U22574 (N_22574,N_22476,N_22492);
xnor U22575 (N_22575,N_22464,N_22385);
nand U22576 (N_22576,N_22433,N_22341);
xor U22577 (N_22577,N_22445,N_22332);
nor U22578 (N_22578,N_22449,N_22431);
and U22579 (N_22579,N_22398,N_22406);
or U22580 (N_22580,N_22498,N_22264);
xnor U22581 (N_22581,N_22463,N_22393);
nor U22582 (N_22582,N_22430,N_22488);
nand U22583 (N_22583,N_22455,N_22365);
or U22584 (N_22584,N_22276,N_22405);
xor U22585 (N_22585,N_22422,N_22326);
xor U22586 (N_22586,N_22468,N_22460);
nand U22587 (N_22587,N_22471,N_22266);
or U22588 (N_22588,N_22432,N_22256);
nor U22589 (N_22589,N_22324,N_22300);
and U22590 (N_22590,N_22421,N_22339);
or U22591 (N_22591,N_22259,N_22353);
xnor U22592 (N_22592,N_22466,N_22482);
xnor U22593 (N_22593,N_22410,N_22343);
and U22594 (N_22594,N_22375,N_22281);
or U22595 (N_22595,N_22462,N_22297);
or U22596 (N_22596,N_22465,N_22310);
nor U22597 (N_22597,N_22361,N_22404);
or U22598 (N_22598,N_22316,N_22287);
nand U22599 (N_22599,N_22257,N_22278);
xnor U22600 (N_22600,N_22314,N_22395);
and U22601 (N_22601,N_22283,N_22255);
nor U22602 (N_22602,N_22402,N_22415);
and U22603 (N_22603,N_22380,N_22435);
xnor U22604 (N_22604,N_22301,N_22292);
or U22605 (N_22605,N_22371,N_22401);
nand U22606 (N_22606,N_22454,N_22386);
nor U22607 (N_22607,N_22322,N_22274);
nand U22608 (N_22608,N_22428,N_22373);
nand U22609 (N_22609,N_22382,N_22293);
or U22610 (N_22610,N_22434,N_22303);
xnor U22611 (N_22611,N_22250,N_22335);
and U22612 (N_22612,N_22378,N_22427);
xor U22613 (N_22613,N_22420,N_22499);
nor U22614 (N_22614,N_22456,N_22340);
nand U22615 (N_22615,N_22260,N_22368);
nor U22616 (N_22616,N_22280,N_22291);
xor U22617 (N_22617,N_22389,N_22252);
and U22618 (N_22618,N_22377,N_22330);
and U22619 (N_22619,N_22290,N_22334);
or U22620 (N_22620,N_22484,N_22479);
nor U22621 (N_22621,N_22447,N_22376);
nand U22622 (N_22622,N_22275,N_22309);
nor U22623 (N_22623,N_22459,N_22412);
xnor U22624 (N_22624,N_22354,N_22337);
and U22625 (N_22625,N_22487,N_22435);
and U22626 (N_22626,N_22446,N_22415);
or U22627 (N_22627,N_22375,N_22490);
xnor U22628 (N_22628,N_22409,N_22422);
nor U22629 (N_22629,N_22433,N_22462);
or U22630 (N_22630,N_22438,N_22451);
xnor U22631 (N_22631,N_22489,N_22283);
xor U22632 (N_22632,N_22290,N_22307);
xor U22633 (N_22633,N_22261,N_22368);
xnor U22634 (N_22634,N_22338,N_22420);
nor U22635 (N_22635,N_22325,N_22397);
nand U22636 (N_22636,N_22307,N_22383);
nor U22637 (N_22637,N_22477,N_22440);
xnor U22638 (N_22638,N_22466,N_22442);
nand U22639 (N_22639,N_22394,N_22362);
or U22640 (N_22640,N_22344,N_22316);
nor U22641 (N_22641,N_22446,N_22433);
xor U22642 (N_22642,N_22343,N_22270);
or U22643 (N_22643,N_22277,N_22469);
and U22644 (N_22644,N_22456,N_22364);
nand U22645 (N_22645,N_22452,N_22312);
or U22646 (N_22646,N_22378,N_22434);
xor U22647 (N_22647,N_22499,N_22314);
and U22648 (N_22648,N_22379,N_22425);
nand U22649 (N_22649,N_22489,N_22271);
xnor U22650 (N_22650,N_22297,N_22257);
nor U22651 (N_22651,N_22415,N_22304);
and U22652 (N_22652,N_22344,N_22273);
or U22653 (N_22653,N_22259,N_22324);
and U22654 (N_22654,N_22466,N_22434);
nand U22655 (N_22655,N_22415,N_22488);
xnor U22656 (N_22656,N_22478,N_22357);
nor U22657 (N_22657,N_22465,N_22407);
and U22658 (N_22658,N_22467,N_22451);
nand U22659 (N_22659,N_22343,N_22498);
xor U22660 (N_22660,N_22397,N_22338);
or U22661 (N_22661,N_22275,N_22483);
or U22662 (N_22662,N_22287,N_22302);
nand U22663 (N_22663,N_22258,N_22315);
nor U22664 (N_22664,N_22425,N_22442);
nand U22665 (N_22665,N_22298,N_22478);
xnor U22666 (N_22666,N_22447,N_22347);
or U22667 (N_22667,N_22255,N_22270);
nor U22668 (N_22668,N_22275,N_22478);
nand U22669 (N_22669,N_22433,N_22412);
nor U22670 (N_22670,N_22428,N_22321);
and U22671 (N_22671,N_22332,N_22433);
nand U22672 (N_22672,N_22495,N_22392);
nor U22673 (N_22673,N_22453,N_22466);
or U22674 (N_22674,N_22303,N_22444);
or U22675 (N_22675,N_22358,N_22343);
xnor U22676 (N_22676,N_22416,N_22363);
nor U22677 (N_22677,N_22469,N_22407);
nor U22678 (N_22678,N_22470,N_22395);
xnor U22679 (N_22679,N_22344,N_22302);
xor U22680 (N_22680,N_22398,N_22283);
nand U22681 (N_22681,N_22326,N_22402);
xnor U22682 (N_22682,N_22487,N_22366);
xnor U22683 (N_22683,N_22415,N_22469);
nor U22684 (N_22684,N_22270,N_22268);
and U22685 (N_22685,N_22339,N_22444);
or U22686 (N_22686,N_22273,N_22314);
and U22687 (N_22687,N_22422,N_22284);
nor U22688 (N_22688,N_22358,N_22474);
nand U22689 (N_22689,N_22345,N_22389);
or U22690 (N_22690,N_22321,N_22349);
nand U22691 (N_22691,N_22344,N_22326);
and U22692 (N_22692,N_22305,N_22463);
and U22693 (N_22693,N_22439,N_22336);
or U22694 (N_22694,N_22427,N_22409);
xnor U22695 (N_22695,N_22494,N_22414);
or U22696 (N_22696,N_22439,N_22454);
xor U22697 (N_22697,N_22315,N_22473);
or U22698 (N_22698,N_22396,N_22446);
nand U22699 (N_22699,N_22437,N_22310);
and U22700 (N_22700,N_22285,N_22250);
nand U22701 (N_22701,N_22326,N_22490);
or U22702 (N_22702,N_22458,N_22331);
nand U22703 (N_22703,N_22375,N_22498);
nand U22704 (N_22704,N_22372,N_22371);
or U22705 (N_22705,N_22438,N_22419);
or U22706 (N_22706,N_22462,N_22400);
and U22707 (N_22707,N_22452,N_22406);
nand U22708 (N_22708,N_22351,N_22483);
nand U22709 (N_22709,N_22334,N_22466);
xnor U22710 (N_22710,N_22375,N_22367);
nand U22711 (N_22711,N_22414,N_22286);
and U22712 (N_22712,N_22250,N_22479);
and U22713 (N_22713,N_22344,N_22258);
and U22714 (N_22714,N_22294,N_22396);
xnor U22715 (N_22715,N_22382,N_22301);
xor U22716 (N_22716,N_22325,N_22362);
xor U22717 (N_22717,N_22445,N_22468);
or U22718 (N_22718,N_22428,N_22333);
nand U22719 (N_22719,N_22381,N_22378);
nor U22720 (N_22720,N_22306,N_22445);
and U22721 (N_22721,N_22436,N_22285);
or U22722 (N_22722,N_22351,N_22427);
and U22723 (N_22723,N_22365,N_22408);
or U22724 (N_22724,N_22365,N_22251);
or U22725 (N_22725,N_22354,N_22351);
nand U22726 (N_22726,N_22329,N_22288);
nand U22727 (N_22727,N_22350,N_22341);
nor U22728 (N_22728,N_22439,N_22253);
xor U22729 (N_22729,N_22387,N_22250);
nand U22730 (N_22730,N_22376,N_22499);
nand U22731 (N_22731,N_22366,N_22393);
or U22732 (N_22732,N_22424,N_22331);
nand U22733 (N_22733,N_22446,N_22321);
nand U22734 (N_22734,N_22353,N_22436);
nand U22735 (N_22735,N_22282,N_22357);
nor U22736 (N_22736,N_22463,N_22314);
nand U22737 (N_22737,N_22467,N_22416);
or U22738 (N_22738,N_22459,N_22435);
xnor U22739 (N_22739,N_22308,N_22323);
xnor U22740 (N_22740,N_22274,N_22319);
xor U22741 (N_22741,N_22328,N_22403);
nand U22742 (N_22742,N_22253,N_22285);
and U22743 (N_22743,N_22429,N_22409);
and U22744 (N_22744,N_22450,N_22423);
nor U22745 (N_22745,N_22472,N_22493);
xor U22746 (N_22746,N_22375,N_22269);
and U22747 (N_22747,N_22250,N_22450);
and U22748 (N_22748,N_22377,N_22453);
nor U22749 (N_22749,N_22475,N_22424);
xor U22750 (N_22750,N_22559,N_22505);
and U22751 (N_22751,N_22740,N_22736);
xor U22752 (N_22752,N_22697,N_22577);
nor U22753 (N_22753,N_22538,N_22598);
or U22754 (N_22754,N_22566,N_22550);
nand U22755 (N_22755,N_22721,N_22596);
and U22756 (N_22756,N_22664,N_22618);
nor U22757 (N_22757,N_22585,N_22643);
nor U22758 (N_22758,N_22680,N_22526);
and U22759 (N_22759,N_22708,N_22686);
nor U22760 (N_22760,N_22645,N_22517);
nor U22761 (N_22761,N_22616,N_22569);
or U22762 (N_22762,N_22570,N_22628);
and U22763 (N_22763,N_22738,N_22531);
xnor U22764 (N_22764,N_22611,N_22675);
nor U22765 (N_22765,N_22734,N_22743);
nor U22766 (N_22766,N_22695,N_22667);
nor U22767 (N_22767,N_22516,N_22520);
nor U22768 (N_22768,N_22701,N_22603);
nand U22769 (N_22769,N_22523,N_22732);
xor U22770 (N_22770,N_22625,N_22744);
and U22771 (N_22771,N_22678,N_22528);
or U22772 (N_22772,N_22606,N_22655);
nor U22773 (N_22773,N_22703,N_22692);
or U22774 (N_22774,N_22614,N_22612);
and U22775 (N_22775,N_22557,N_22620);
nor U22776 (N_22776,N_22709,N_22513);
and U22777 (N_22777,N_22601,N_22632);
nor U22778 (N_22778,N_22574,N_22619);
and U22779 (N_22779,N_22607,N_22699);
or U22780 (N_22780,N_22580,N_22737);
and U22781 (N_22781,N_22705,N_22503);
nor U22782 (N_22782,N_22656,N_22524);
and U22783 (N_22783,N_22545,N_22706);
and U22784 (N_22784,N_22514,N_22565);
or U22785 (N_22785,N_22593,N_22636);
nor U22786 (N_22786,N_22584,N_22689);
nand U22787 (N_22787,N_22543,N_22600);
xor U22788 (N_22788,N_22613,N_22717);
nand U22789 (N_22789,N_22561,N_22579);
nor U22790 (N_22790,N_22556,N_22749);
and U22791 (N_22791,N_22534,N_22564);
or U22792 (N_22792,N_22581,N_22509);
and U22793 (N_22793,N_22602,N_22535);
nor U22794 (N_22794,N_22525,N_22739);
xor U22795 (N_22795,N_22595,N_22672);
or U22796 (N_22796,N_22633,N_22508);
xnor U22797 (N_22797,N_22500,N_22702);
xor U22798 (N_22798,N_22591,N_22502);
and U22799 (N_22799,N_22587,N_22573);
and U22800 (N_22800,N_22677,N_22712);
xor U22801 (N_22801,N_22653,N_22527);
nor U22802 (N_22802,N_22647,N_22548);
nor U22803 (N_22803,N_22745,N_22644);
nor U22804 (N_22804,N_22637,N_22714);
xor U22805 (N_22805,N_22501,N_22729);
nor U22806 (N_22806,N_22670,N_22683);
or U22807 (N_22807,N_22666,N_22617);
and U22808 (N_22808,N_22693,N_22571);
xor U22809 (N_22809,N_22641,N_22624);
nor U22810 (N_22810,N_22568,N_22642);
and U22811 (N_22811,N_22506,N_22583);
nand U22812 (N_22812,N_22630,N_22631);
xnor U22813 (N_22813,N_22536,N_22687);
nor U22814 (N_22814,N_22518,N_22649);
nor U22815 (N_22815,N_22541,N_22588);
or U22816 (N_22816,N_22623,N_22594);
or U22817 (N_22817,N_22676,N_22662);
xnor U22818 (N_22818,N_22741,N_22589);
and U22819 (N_22819,N_22747,N_22519);
and U22820 (N_22820,N_22746,N_22731);
nor U22821 (N_22821,N_22562,N_22638);
or U22822 (N_22822,N_22651,N_22665);
and U22823 (N_22823,N_22515,N_22733);
and U22824 (N_22824,N_22544,N_22742);
xnor U22825 (N_22825,N_22671,N_22553);
and U22826 (N_22826,N_22660,N_22661);
xor U22827 (N_22827,N_22521,N_22627);
and U22828 (N_22828,N_22681,N_22720);
or U22829 (N_22829,N_22572,N_22694);
nand U22830 (N_22830,N_22552,N_22510);
xnor U22831 (N_22831,N_22567,N_22599);
and U22832 (N_22832,N_22540,N_22657);
nand U22833 (N_22833,N_22615,N_22622);
nor U22834 (N_22834,N_22608,N_22654);
and U22835 (N_22835,N_22533,N_22609);
nor U22836 (N_22836,N_22512,N_22711);
nor U22837 (N_22837,N_22719,N_22725);
and U22838 (N_22838,N_22529,N_22727);
nand U22839 (N_22839,N_22610,N_22646);
nand U22840 (N_22840,N_22707,N_22555);
nor U22841 (N_22841,N_22718,N_22626);
or U22842 (N_22842,N_22582,N_22507);
nand U22843 (N_22843,N_22648,N_22723);
nand U22844 (N_22844,N_22639,N_22704);
and U22845 (N_22845,N_22668,N_22669);
xnor U22846 (N_22846,N_22549,N_22578);
nor U22847 (N_22847,N_22592,N_22722);
nand U22848 (N_22848,N_22640,N_22537);
xnor U22849 (N_22849,N_22716,N_22728);
or U22850 (N_22850,N_22700,N_22522);
nor U22851 (N_22851,N_22635,N_22730);
or U22852 (N_22852,N_22575,N_22684);
nand U22853 (N_22853,N_22554,N_22547);
nand U22854 (N_22854,N_22688,N_22696);
or U22855 (N_22855,N_22576,N_22530);
xnor U22856 (N_22856,N_22673,N_22590);
or U22857 (N_22857,N_22663,N_22539);
and U22858 (N_22858,N_22605,N_22551);
or U22859 (N_22859,N_22679,N_22690);
nor U22860 (N_22860,N_22504,N_22604);
nand U22861 (N_22861,N_22629,N_22621);
or U22862 (N_22862,N_22659,N_22650);
or U22863 (N_22863,N_22735,N_22511);
or U22864 (N_22864,N_22713,N_22726);
and U22865 (N_22865,N_22685,N_22558);
and U22866 (N_22866,N_22532,N_22652);
nor U22867 (N_22867,N_22586,N_22698);
or U22868 (N_22868,N_22560,N_22682);
or U22869 (N_22869,N_22542,N_22715);
and U22870 (N_22870,N_22674,N_22597);
xnor U22871 (N_22871,N_22546,N_22710);
nand U22872 (N_22872,N_22691,N_22724);
nand U22873 (N_22873,N_22658,N_22563);
nand U22874 (N_22874,N_22748,N_22634);
xor U22875 (N_22875,N_22545,N_22600);
nor U22876 (N_22876,N_22514,N_22744);
nor U22877 (N_22877,N_22590,N_22716);
nand U22878 (N_22878,N_22667,N_22584);
nand U22879 (N_22879,N_22712,N_22662);
and U22880 (N_22880,N_22740,N_22723);
and U22881 (N_22881,N_22667,N_22697);
nand U22882 (N_22882,N_22720,N_22669);
or U22883 (N_22883,N_22715,N_22716);
nand U22884 (N_22884,N_22586,N_22566);
nand U22885 (N_22885,N_22729,N_22706);
xnor U22886 (N_22886,N_22570,N_22555);
nand U22887 (N_22887,N_22728,N_22696);
nand U22888 (N_22888,N_22645,N_22675);
nor U22889 (N_22889,N_22620,N_22611);
or U22890 (N_22890,N_22508,N_22747);
or U22891 (N_22891,N_22701,N_22728);
nor U22892 (N_22892,N_22580,N_22587);
xnor U22893 (N_22893,N_22552,N_22614);
nor U22894 (N_22894,N_22541,N_22597);
xnor U22895 (N_22895,N_22737,N_22687);
or U22896 (N_22896,N_22524,N_22727);
and U22897 (N_22897,N_22682,N_22641);
and U22898 (N_22898,N_22593,N_22619);
nor U22899 (N_22899,N_22521,N_22698);
xnor U22900 (N_22900,N_22512,N_22589);
and U22901 (N_22901,N_22541,N_22594);
and U22902 (N_22902,N_22686,N_22665);
nand U22903 (N_22903,N_22501,N_22571);
nor U22904 (N_22904,N_22505,N_22551);
or U22905 (N_22905,N_22660,N_22606);
and U22906 (N_22906,N_22512,N_22655);
nor U22907 (N_22907,N_22717,N_22731);
xor U22908 (N_22908,N_22698,N_22644);
nand U22909 (N_22909,N_22624,N_22609);
and U22910 (N_22910,N_22703,N_22688);
nor U22911 (N_22911,N_22535,N_22710);
and U22912 (N_22912,N_22695,N_22689);
or U22913 (N_22913,N_22680,N_22608);
xor U22914 (N_22914,N_22726,N_22595);
nand U22915 (N_22915,N_22711,N_22644);
and U22916 (N_22916,N_22614,N_22508);
xor U22917 (N_22917,N_22569,N_22658);
and U22918 (N_22918,N_22628,N_22695);
and U22919 (N_22919,N_22718,N_22520);
nand U22920 (N_22920,N_22542,N_22560);
nor U22921 (N_22921,N_22503,N_22667);
xor U22922 (N_22922,N_22552,N_22738);
nand U22923 (N_22923,N_22528,N_22721);
xnor U22924 (N_22924,N_22577,N_22641);
or U22925 (N_22925,N_22732,N_22662);
or U22926 (N_22926,N_22530,N_22591);
nor U22927 (N_22927,N_22554,N_22715);
nor U22928 (N_22928,N_22574,N_22685);
or U22929 (N_22929,N_22625,N_22710);
nor U22930 (N_22930,N_22693,N_22583);
and U22931 (N_22931,N_22631,N_22570);
nor U22932 (N_22932,N_22624,N_22678);
nor U22933 (N_22933,N_22720,N_22602);
nand U22934 (N_22934,N_22572,N_22638);
nand U22935 (N_22935,N_22543,N_22611);
or U22936 (N_22936,N_22528,N_22737);
xnor U22937 (N_22937,N_22674,N_22602);
nand U22938 (N_22938,N_22646,N_22628);
xor U22939 (N_22939,N_22545,N_22659);
xnor U22940 (N_22940,N_22557,N_22743);
nand U22941 (N_22941,N_22633,N_22698);
xnor U22942 (N_22942,N_22603,N_22593);
or U22943 (N_22943,N_22592,N_22682);
and U22944 (N_22944,N_22628,N_22523);
nand U22945 (N_22945,N_22512,N_22661);
nand U22946 (N_22946,N_22729,N_22570);
xor U22947 (N_22947,N_22678,N_22674);
nor U22948 (N_22948,N_22669,N_22535);
nor U22949 (N_22949,N_22702,N_22635);
nand U22950 (N_22950,N_22747,N_22554);
nand U22951 (N_22951,N_22667,N_22648);
nor U22952 (N_22952,N_22742,N_22643);
and U22953 (N_22953,N_22535,N_22734);
and U22954 (N_22954,N_22673,N_22675);
and U22955 (N_22955,N_22653,N_22716);
and U22956 (N_22956,N_22733,N_22728);
and U22957 (N_22957,N_22597,N_22515);
nor U22958 (N_22958,N_22526,N_22625);
xor U22959 (N_22959,N_22723,N_22510);
nor U22960 (N_22960,N_22554,N_22703);
xor U22961 (N_22961,N_22633,N_22614);
xor U22962 (N_22962,N_22503,N_22582);
nor U22963 (N_22963,N_22600,N_22522);
xor U22964 (N_22964,N_22632,N_22679);
or U22965 (N_22965,N_22515,N_22726);
nand U22966 (N_22966,N_22569,N_22731);
and U22967 (N_22967,N_22581,N_22695);
nor U22968 (N_22968,N_22660,N_22735);
nor U22969 (N_22969,N_22562,N_22697);
nor U22970 (N_22970,N_22606,N_22713);
nor U22971 (N_22971,N_22591,N_22508);
or U22972 (N_22972,N_22649,N_22580);
and U22973 (N_22973,N_22533,N_22598);
xor U22974 (N_22974,N_22524,N_22728);
and U22975 (N_22975,N_22534,N_22576);
xnor U22976 (N_22976,N_22568,N_22506);
nor U22977 (N_22977,N_22626,N_22610);
nand U22978 (N_22978,N_22708,N_22576);
and U22979 (N_22979,N_22632,N_22735);
or U22980 (N_22980,N_22697,N_22532);
xnor U22981 (N_22981,N_22676,N_22604);
or U22982 (N_22982,N_22586,N_22570);
xnor U22983 (N_22983,N_22673,N_22605);
or U22984 (N_22984,N_22542,N_22599);
nand U22985 (N_22985,N_22716,N_22602);
or U22986 (N_22986,N_22593,N_22564);
or U22987 (N_22987,N_22714,N_22675);
or U22988 (N_22988,N_22716,N_22652);
nand U22989 (N_22989,N_22580,N_22586);
nand U22990 (N_22990,N_22640,N_22689);
and U22991 (N_22991,N_22730,N_22584);
nand U22992 (N_22992,N_22560,N_22689);
and U22993 (N_22993,N_22566,N_22722);
or U22994 (N_22994,N_22625,N_22630);
nor U22995 (N_22995,N_22726,N_22551);
and U22996 (N_22996,N_22692,N_22709);
nor U22997 (N_22997,N_22719,N_22671);
nand U22998 (N_22998,N_22501,N_22677);
and U22999 (N_22999,N_22555,N_22713);
nor U23000 (N_23000,N_22819,N_22877);
nor U23001 (N_23001,N_22796,N_22751);
and U23002 (N_23002,N_22879,N_22957);
and U23003 (N_23003,N_22864,N_22804);
nor U23004 (N_23004,N_22894,N_22897);
nand U23005 (N_23005,N_22997,N_22985);
or U23006 (N_23006,N_22931,N_22867);
nand U23007 (N_23007,N_22945,N_22916);
nand U23008 (N_23008,N_22885,N_22801);
or U23009 (N_23009,N_22893,N_22798);
nand U23010 (N_23010,N_22881,N_22861);
and U23011 (N_23011,N_22770,N_22942);
xor U23012 (N_23012,N_22757,N_22859);
nand U23013 (N_23013,N_22763,N_22995);
or U23014 (N_23014,N_22788,N_22871);
and U23015 (N_23015,N_22803,N_22836);
nand U23016 (N_23016,N_22809,N_22907);
and U23017 (N_23017,N_22849,N_22996);
or U23018 (N_23018,N_22758,N_22903);
nand U23019 (N_23019,N_22845,N_22905);
and U23020 (N_23020,N_22834,N_22917);
and U23021 (N_23021,N_22781,N_22984);
nor U23022 (N_23022,N_22908,N_22896);
nand U23023 (N_23023,N_22844,N_22765);
nand U23024 (N_23024,N_22777,N_22938);
and U23025 (N_23025,N_22878,N_22780);
and U23026 (N_23026,N_22838,N_22767);
xor U23027 (N_23027,N_22817,N_22776);
xnor U23028 (N_23028,N_22883,N_22806);
nor U23029 (N_23029,N_22914,N_22768);
or U23030 (N_23030,N_22766,N_22888);
xnor U23031 (N_23031,N_22755,N_22863);
xnor U23032 (N_23032,N_22855,N_22784);
xnor U23033 (N_23033,N_22912,N_22818);
xor U23034 (N_23034,N_22927,N_22955);
nor U23035 (N_23035,N_22994,N_22899);
or U23036 (N_23036,N_22876,N_22968);
xnor U23037 (N_23037,N_22810,N_22828);
xor U23038 (N_23038,N_22975,N_22926);
and U23039 (N_23039,N_22753,N_22973);
nand U23040 (N_23040,N_22948,N_22872);
nor U23041 (N_23041,N_22841,N_22986);
or U23042 (N_23042,N_22779,N_22808);
nand U23043 (N_23043,N_22981,N_22873);
nor U23044 (N_23044,N_22869,N_22762);
and U23045 (N_23045,N_22936,N_22771);
or U23046 (N_23046,N_22971,N_22987);
xnor U23047 (N_23047,N_22998,N_22901);
and U23048 (N_23048,N_22812,N_22830);
nor U23049 (N_23049,N_22963,N_22786);
xor U23050 (N_23050,N_22949,N_22865);
or U23051 (N_23051,N_22946,N_22935);
xnor U23052 (N_23052,N_22813,N_22993);
nand U23053 (N_23053,N_22799,N_22842);
and U23054 (N_23054,N_22759,N_22937);
and U23055 (N_23055,N_22795,N_22892);
or U23056 (N_23056,N_22951,N_22891);
or U23057 (N_23057,N_22953,N_22923);
and U23058 (N_23058,N_22807,N_22852);
nor U23059 (N_23059,N_22827,N_22970);
or U23060 (N_23060,N_22843,N_22823);
and U23061 (N_23061,N_22911,N_22857);
and U23062 (N_23062,N_22778,N_22764);
nor U23063 (N_23063,N_22825,N_22824);
xnor U23064 (N_23064,N_22754,N_22954);
nand U23065 (N_23065,N_22805,N_22972);
or U23066 (N_23066,N_22976,N_22909);
nor U23067 (N_23067,N_22956,N_22884);
or U23068 (N_23068,N_22761,N_22882);
and U23069 (N_23069,N_22750,N_22904);
xor U23070 (N_23070,N_22832,N_22977);
xnor U23071 (N_23071,N_22835,N_22858);
and U23072 (N_23072,N_22958,N_22895);
xor U23073 (N_23073,N_22840,N_22846);
and U23074 (N_23074,N_22815,N_22769);
or U23075 (N_23075,N_22811,N_22792);
xor U23076 (N_23076,N_22928,N_22760);
nand U23077 (N_23077,N_22831,N_22790);
nor U23078 (N_23078,N_22874,N_22964);
xnor U23079 (N_23079,N_22921,N_22837);
nor U23080 (N_23080,N_22965,N_22829);
nand U23081 (N_23081,N_22851,N_22756);
and U23082 (N_23082,N_22772,N_22787);
or U23083 (N_23083,N_22919,N_22880);
and U23084 (N_23084,N_22794,N_22800);
nand U23085 (N_23085,N_22943,N_22952);
nand U23086 (N_23086,N_22922,N_22791);
and U23087 (N_23087,N_22939,N_22982);
nor U23088 (N_23088,N_22816,N_22814);
xor U23089 (N_23089,N_22782,N_22980);
and U23090 (N_23090,N_22925,N_22797);
xor U23091 (N_23091,N_22886,N_22868);
nor U23092 (N_23092,N_22913,N_22860);
and U23093 (N_23093,N_22822,N_22989);
nor U23094 (N_23094,N_22934,N_22802);
nand U23095 (N_23095,N_22785,N_22906);
xor U23096 (N_23096,N_22870,N_22889);
nor U23097 (N_23097,N_22950,N_22941);
nand U23098 (N_23098,N_22752,N_22966);
nor U23099 (N_23099,N_22862,N_22826);
nand U23100 (N_23100,N_22856,N_22990);
or U23101 (N_23101,N_22978,N_22932);
xnor U23102 (N_23102,N_22789,N_22967);
and U23103 (N_23103,N_22839,N_22960);
nand U23104 (N_23104,N_22773,N_22898);
and U23105 (N_23105,N_22979,N_22774);
nor U23106 (N_23106,N_22930,N_22961);
xnor U23107 (N_23107,N_22783,N_22820);
nor U23108 (N_23108,N_22902,N_22848);
or U23109 (N_23109,N_22833,N_22924);
or U23110 (N_23110,N_22821,N_22969);
nand U23111 (N_23111,N_22959,N_22983);
xnor U23112 (N_23112,N_22992,N_22962);
nor U23113 (N_23113,N_22910,N_22793);
xor U23114 (N_23114,N_22890,N_22887);
nand U23115 (N_23115,N_22918,N_22974);
xor U23116 (N_23116,N_22988,N_22875);
nor U23117 (N_23117,N_22991,N_22850);
nand U23118 (N_23118,N_22866,N_22775);
nand U23119 (N_23119,N_22940,N_22853);
or U23120 (N_23120,N_22929,N_22847);
xnor U23121 (N_23121,N_22915,N_22900);
nand U23122 (N_23122,N_22933,N_22944);
nand U23123 (N_23123,N_22999,N_22920);
xor U23124 (N_23124,N_22854,N_22947);
and U23125 (N_23125,N_22894,N_22953);
nor U23126 (N_23126,N_22936,N_22914);
or U23127 (N_23127,N_22787,N_22979);
and U23128 (N_23128,N_22964,N_22848);
xnor U23129 (N_23129,N_22763,N_22806);
and U23130 (N_23130,N_22785,N_22810);
xor U23131 (N_23131,N_22804,N_22839);
xnor U23132 (N_23132,N_22927,N_22795);
or U23133 (N_23133,N_22836,N_22752);
xor U23134 (N_23134,N_22994,N_22794);
or U23135 (N_23135,N_22896,N_22934);
nor U23136 (N_23136,N_22875,N_22909);
and U23137 (N_23137,N_22833,N_22886);
nand U23138 (N_23138,N_22999,N_22985);
or U23139 (N_23139,N_22938,N_22884);
and U23140 (N_23140,N_22795,N_22998);
nand U23141 (N_23141,N_22820,N_22905);
nor U23142 (N_23142,N_22789,N_22994);
xnor U23143 (N_23143,N_22804,N_22756);
nor U23144 (N_23144,N_22771,N_22777);
nand U23145 (N_23145,N_22791,N_22814);
or U23146 (N_23146,N_22764,N_22838);
xor U23147 (N_23147,N_22999,N_22800);
xor U23148 (N_23148,N_22854,N_22771);
nand U23149 (N_23149,N_22870,N_22900);
xor U23150 (N_23150,N_22843,N_22910);
xnor U23151 (N_23151,N_22873,N_22976);
and U23152 (N_23152,N_22761,N_22811);
and U23153 (N_23153,N_22842,N_22802);
or U23154 (N_23154,N_22849,N_22998);
xnor U23155 (N_23155,N_22979,N_22864);
or U23156 (N_23156,N_22750,N_22789);
xnor U23157 (N_23157,N_22969,N_22808);
and U23158 (N_23158,N_22851,N_22926);
xor U23159 (N_23159,N_22755,N_22952);
and U23160 (N_23160,N_22798,N_22888);
nor U23161 (N_23161,N_22918,N_22913);
nand U23162 (N_23162,N_22977,N_22986);
nor U23163 (N_23163,N_22879,N_22839);
nor U23164 (N_23164,N_22757,N_22877);
nand U23165 (N_23165,N_22789,N_22937);
nand U23166 (N_23166,N_22864,N_22823);
nor U23167 (N_23167,N_22761,N_22915);
and U23168 (N_23168,N_22840,N_22863);
nand U23169 (N_23169,N_22753,N_22967);
and U23170 (N_23170,N_22802,N_22977);
nand U23171 (N_23171,N_22810,N_22816);
xnor U23172 (N_23172,N_22940,N_22865);
or U23173 (N_23173,N_22755,N_22785);
nand U23174 (N_23174,N_22820,N_22823);
nor U23175 (N_23175,N_22787,N_22882);
or U23176 (N_23176,N_22763,N_22981);
or U23177 (N_23177,N_22831,N_22835);
xor U23178 (N_23178,N_22987,N_22862);
nand U23179 (N_23179,N_22905,N_22987);
nor U23180 (N_23180,N_22965,N_22855);
nor U23181 (N_23181,N_22932,N_22755);
nor U23182 (N_23182,N_22906,N_22870);
or U23183 (N_23183,N_22789,N_22849);
and U23184 (N_23184,N_22982,N_22755);
nand U23185 (N_23185,N_22833,N_22768);
xnor U23186 (N_23186,N_22768,N_22943);
xor U23187 (N_23187,N_22859,N_22823);
nor U23188 (N_23188,N_22960,N_22895);
or U23189 (N_23189,N_22792,N_22923);
or U23190 (N_23190,N_22813,N_22932);
or U23191 (N_23191,N_22889,N_22959);
xor U23192 (N_23192,N_22774,N_22770);
xnor U23193 (N_23193,N_22944,N_22927);
xor U23194 (N_23194,N_22805,N_22950);
nand U23195 (N_23195,N_22802,N_22912);
and U23196 (N_23196,N_22819,N_22906);
nor U23197 (N_23197,N_22893,N_22920);
or U23198 (N_23198,N_22788,N_22791);
nand U23199 (N_23199,N_22803,N_22855);
or U23200 (N_23200,N_22778,N_22790);
nor U23201 (N_23201,N_22790,N_22982);
or U23202 (N_23202,N_22883,N_22971);
and U23203 (N_23203,N_22920,N_22896);
or U23204 (N_23204,N_22840,N_22860);
or U23205 (N_23205,N_22908,N_22800);
or U23206 (N_23206,N_22839,N_22767);
nand U23207 (N_23207,N_22816,N_22819);
and U23208 (N_23208,N_22837,N_22779);
xnor U23209 (N_23209,N_22888,N_22930);
nand U23210 (N_23210,N_22952,N_22838);
nand U23211 (N_23211,N_22966,N_22886);
nor U23212 (N_23212,N_22787,N_22942);
nor U23213 (N_23213,N_22817,N_22952);
or U23214 (N_23214,N_22911,N_22785);
and U23215 (N_23215,N_22967,N_22765);
nand U23216 (N_23216,N_22783,N_22832);
nor U23217 (N_23217,N_22962,N_22784);
nand U23218 (N_23218,N_22891,N_22980);
and U23219 (N_23219,N_22790,N_22966);
xor U23220 (N_23220,N_22859,N_22940);
nand U23221 (N_23221,N_22877,N_22812);
nand U23222 (N_23222,N_22842,N_22833);
nand U23223 (N_23223,N_22852,N_22870);
or U23224 (N_23224,N_22883,N_22963);
nand U23225 (N_23225,N_22931,N_22757);
nor U23226 (N_23226,N_22860,N_22985);
nand U23227 (N_23227,N_22929,N_22920);
nor U23228 (N_23228,N_22884,N_22787);
and U23229 (N_23229,N_22835,N_22792);
nor U23230 (N_23230,N_22816,N_22964);
xor U23231 (N_23231,N_22971,N_22810);
nand U23232 (N_23232,N_22837,N_22763);
and U23233 (N_23233,N_22922,N_22982);
nand U23234 (N_23234,N_22918,N_22770);
xor U23235 (N_23235,N_22854,N_22790);
nand U23236 (N_23236,N_22761,N_22972);
xor U23237 (N_23237,N_22789,N_22766);
and U23238 (N_23238,N_22871,N_22924);
nor U23239 (N_23239,N_22815,N_22935);
and U23240 (N_23240,N_22900,N_22939);
or U23241 (N_23241,N_22823,N_22791);
xnor U23242 (N_23242,N_22884,N_22816);
nor U23243 (N_23243,N_22924,N_22912);
nor U23244 (N_23244,N_22857,N_22885);
nand U23245 (N_23245,N_22855,N_22755);
and U23246 (N_23246,N_22994,N_22812);
xor U23247 (N_23247,N_22819,N_22975);
xor U23248 (N_23248,N_22815,N_22751);
xnor U23249 (N_23249,N_22894,N_22780);
nand U23250 (N_23250,N_23139,N_23177);
nor U23251 (N_23251,N_23098,N_23220);
xnor U23252 (N_23252,N_23238,N_23173);
or U23253 (N_23253,N_23086,N_23130);
or U23254 (N_23254,N_23198,N_23137);
and U23255 (N_23255,N_23223,N_23176);
nand U23256 (N_23256,N_23032,N_23247);
and U23257 (N_23257,N_23231,N_23246);
nand U23258 (N_23258,N_23071,N_23197);
xnor U23259 (N_23259,N_23169,N_23070);
nand U23260 (N_23260,N_23044,N_23015);
nor U23261 (N_23261,N_23208,N_23064);
nand U23262 (N_23262,N_23055,N_23203);
nand U23263 (N_23263,N_23166,N_23230);
or U23264 (N_23264,N_23034,N_23110);
or U23265 (N_23265,N_23073,N_23028);
xor U23266 (N_23266,N_23219,N_23156);
nor U23267 (N_23267,N_23199,N_23026);
or U23268 (N_23268,N_23186,N_23193);
nand U23269 (N_23269,N_23222,N_23004);
or U23270 (N_23270,N_23120,N_23038);
and U23271 (N_23271,N_23128,N_23147);
xnor U23272 (N_23272,N_23067,N_23085);
and U23273 (N_23273,N_23168,N_23190);
nor U23274 (N_23274,N_23017,N_23171);
xnor U23275 (N_23275,N_23094,N_23194);
nand U23276 (N_23276,N_23043,N_23213);
xnor U23277 (N_23277,N_23083,N_23112);
and U23278 (N_23278,N_23207,N_23123);
nand U23279 (N_23279,N_23188,N_23196);
and U23280 (N_23280,N_23226,N_23144);
xor U23281 (N_23281,N_23142,N_23146);
nor U23282 (N_23282,N_23162,N_23093);
or U23283 (N_23283,N_23016,N_23159);
nor U23284 (N_23284,N_23012,N_23129);
nor U23285 (N_23285,N_23101,N_23145);
and U23286 (N_23286,N_23050,N_23007);
nand U23287 (N_23287,N_23239,N_23107);
and U23288 (N_23288,N_23102,N_23150);
or U23289 (N_23289,N_23087,N_23075);
and U23290 (N_23290,N_23136,N_23019);
and U23291 (N_23291,N_23108,N_23051);
xnor U23292 (N_23292,N_23245,N_23116);
nor U23293 (N_23293,N_23174,N_23240);
and U23294 (N_23294,N_23057,N_23224);
nand U23295 (N_23295,N_23131,N_23049);
or U23296 (N_23296,N_23235,N_23154);
nand U23297 (N_23297,N_23165,N_23185);
nand U23298 (N_23298,N_23233,N_23027);
or U23299 (N_23299,N_23031,N_23180);
nand U23300 (N_23300,N_23062,N_23088);
nor U23301 (N_23301,N_23029,N_23157);
and U23302 (N_23302,N_23042,N_23068);
nand U23303 (N_23303,N_23124,N_23151);
nor U23304 (N_23304,N_23234,N_23024);
nor U23305 (N_23305,N_23148,N_23065);
xnor U23306 (N_23306,N_23006,N_23109);
nand U23307 (N_23307,N_23210,N_23164);
xnor U23308 (N_23308,N_23091,N_23183);
or U23309 (N_23309,N_23018,N_23010);
and U23310 (N_23310,N_23077,N_23084);
xnor U23311 (N_23311,N_23160,N_23033);
nand U23312 (N_23312,N_23105,N_23097);
and U23313 (N_23313,N_23125,N_23022);
nand U23314 (N_23314,N_23149,N_23099);
xor U23315 (N_23315,N_23200,N_23003);
or U23316 (N_23316,N_23013,N_23106);
nor U23317 (N_23317,N_23104,N_23111);
nand U23318 (N_23318,N_23000,N_23229);
nand U23319 (N_23319,N_23076,N_23132);
nand U23320 (N_23320,N_23115,N_23216);
xor U23321 (N_23321,N_23113,N_23126);
or U23322 (N_23322,N_23072,N_23181);
xnor U23323 (N_23323,N_23054,N_23056);
nand U23324 (N_23324,N_23122,N_23047);
nor U23325 (N_23325,N_23211,N_23079);
and U23326 (N_23326,N_23119,N_23249);
nand U23327 (N_23327,N_23036,N_23189);
nor U23328 (N_23328,N_23178,N_23011);
and U23329 (N_23329,N_23035,N_23103);
nand U23330 (N_23330,N_23117,N_23138);
nand U23331 (N_23331,N_23041,N_23179);
nand U23332 (N_23332,N_23046,N_23040);
or U23333 (N_23333,N_23069,N_23228);
and U23334 (N_23334,N_23187,N_23161);
nand U23335 (N_23335,N_23172,N_23121);
xnor U23336 (N_23336,N_23167,N_23025);
or U23337 (N_23337,N_23158,N_23221);
and U23338 (N_23338,N_23143,N_23236);
xnor U23339 (N_23339,N_23175,N_23090);
or U23340 (N_23340,N_23045,N_23244);
or U23341 (N_23341,N_23048,N_23214);
xnor U23342 (N_23342,N_23118,N_23005);
nor U23343 (N_23343,N_23021,N_23227);
nor U23344 (N_23344,N_23081,N_23002);
or U23345 (N_23345,N_23243,N_23023);
and U23346 (N_23346,N_23060,N_23201);
xnor U23347 (N_23347,N_23061,N_23248);
nand U23348 (N_23348,N_23089,N_23078);
xor U23349 (N_23349,N_23192,N_23184);
nand U23350 (N_23350,N_23080,N_23066);
nor U23351 (N_23351,N_23153,N_23212);
nor U23352 (N_23352,N_23205,N_23030);
or U23353 (N_23353,N_23141,N_23058);
or U23354 (N_23354,N_23134,N_23074);
nand U23355 (N_23355,N_23092,N_23237);
xor U23356 (N_23356,N_23063,N_23008);
nand U23357 (N_23357,N_23242,N_23037);
nand U23358 (N_23358,N_23204,N_23096);
and U23359 (N_23359,N_23020,N_23114);
and U23360 (N_23360,N_23135,N_23059);
nor U23361 (N_23361,N_23163,N_23215);
and U23362 (N_23362,N_23140,N_23195);
nor U23363 (N_23363,N_23053,N_23052);
nor U23364 (N_23364,N_23152,N_23217);
or U23365 (N_23365,N_23232,N_23001);
and U23366 (N_23366,N_23082,N_23191);
nor U23367 (N_23367,N_23202,N_23095);
nor U23368 (N_23368,N_23206,N_23133);
nor U23369 (N_23369,N_23182,N_23039);
and U23370 (N_23370,N_23170,N_23225);
xor U23371 (N_23371,N_23127,N_23209);
xor U23372 (N_23372,N_23100,N_23155);
or U23373 (N_23373,N_23241,N_23014);
or U23374 (N_23374,N_23009,N_23218);
xnor U23375 (N_23375,N_23249,N_23118);
or U23376 (N_23376,N_23170,N_23139);
or U23377 (N_23377,N_23167,N_23208);
or U23378 (N_23378,N_23083,N_23231);
nor U23379 (N_23379,N_23022,N_23164);
xor U23380 (N_23380,N_23188,N_23118);
nor U23381 (N_23381,N_23169,N_23248);
and U23382 (N_23382,N_23087,N_23106);
nand U23383 (N_23383,N_23180,N_23168);
and U23384 (N_23384,N_23207,N_23206);
nand U23385 (N_23385,N_23245,N_23019);
and U23386 (N_23386,N_23003,N_23153);
nand U23387 (N_23387,N_23012,N_23044);
or U23388 (N_23388,N_23186,N_23032);
nor U23389 (N_23389,N_23151,N_23134);
and U23390 (N_23390,N_23092,N_23221);
xor U23391 (N_23391,N_23239,N_23047);
and U23392 (N_23392,N_23158,N_23125);
nand U23393 (N_23393,N_23217,N_23009);
and U23394 (N_23394,N_23044,N_23123);
and U23395 (N_23395,N_23103,N_23090);
nor U23396 (N_23396,N_23106,N_23029);
or U23397 (N_23397,N_23144,N_23048);
or U23398 (N_23398,N_23183,N_23094);
or U23399 (N_23399,N_23005,N_23102);
and U23400 (N_23400,N_23189,N_23091);
xnor U23401 (N_23401,N_23006,N_23100);
xnor U23402 (N_23402,N_23165,N_23060);
and U23403 (N_23403,N_23043,N_23244);
nand U23404 (N_23404,N_23016,N_23035);
nand U23405 (N_23405,N_23164,N_23104);
nand U23406 (N_23406,N_23047,N_23191);
and U23407 (N_23407,N_23109,N_23071);
and U23408 (N_23408,N_23175,N_23079);
xor U23409 (N_23409,N_23073,N_23236);
nor U23410 (N_23410,N_23148,N_23071);
and U23411 (N_23411,N_23020,N_23073);
xor U23412 (N_23412,N_23091,N_23199);
nand U23413 (N_23413,N_23190,N_23110);
nor U23414 (N_23414,N_23086,N_23109);
nand U23415 (N_23415,N_23006,N_23029);
or U23416 (N_23416,N_23166,N_23134);
and U23417 (N_23417,N_23125,N_23086);
xor U23418 (N_23418,N_23023,N_23240);
nand U23419 (N_23419,N_23160,N_23196);
nand U23420 (N_23420,N_23247,N_23227);
xor U23421 (N_23421,N_23196,N_23185);
and U23422 (N_23422,N_23150,N_23157);
nor U23423 (N_23423,N_23197,N_23157);
and U23424 (N_23424,N_23227,N_23143);
and U23425 (N_23425,N_23118,N_23121);
nor U23426 (N_23426,N_23247,N_23066);
nor U23427 (N_23427,N_23095,N_23217);
or U23428 (N_23428,N_23006,N_23224);
and U23429 (N_23429,N_23178,N_23099);
and U23430 (N_23430,N_23122,N_23182);
or U23431 (N_23431,N_23074,N_23087);
nand U23432 (N_23432,N_23082,N_23099);
or U23433 (N_23433,N_23121,N_23187);
and U23434 (N_23434,N_23140,N_23001);
xor U23435 (N_23435,N_23087,N_23080);
xor U23436 (N_23436,N_23235,N_23247);
nor U23437 (N_23437,N_23156,N_23062);
or U23438 (N_23438,N_23092,N_23134);
nand U23439 (N_23439,N_23045,N_23032);
and U23440 (N_23440,N_23193,N_23086);
or U23441 (N_23441,N_23226,N_23110);
xnor U23442 (N_23442,N_23180,N_23131);
or U23443 (N_23443,N_23163,N_23213);
nor U23444 (N_23444,N_23109,N_23079);
nor U23445 (N_23445,N_23040,N_23218);
and U23446 (N_23446,N_23244,N_23190);
nor U23447 (N_23447,N_23183,N_23138);
nand U23448 (N_23448,N_23023,N_23014);
or U23449 (N_23449,N_23016,N_23243);
or U23450 (N_23450,N_23001,N_23241);
or U23451 (N_23451,N_23235,N_23018);
nor U23452 (N_23452,N_23147,N_23173);
nand U23453 (N_23453,N_23211,N_23109);
or U23454 (N_23454,N_23207,N_23092);
and U23455 (N_23455,N_23059,N_23180);
nor U23456 (N_23456,N_23142,N_23199);
or U23457 (N_23457,N_23227,N_23092);
or U23458 (N_23458,N_23066,N_23004);
xnor U23459 (N_23459,N_23093,N_23211);
and U23460 (N_23460,N_23184,N_23062);
and U23461 (N_23461,N_23228,N_23081);
or U23462 (N_23462,N_23240,N_23002);
nor U23463 (N_23463,N_23133,N_23194);
nand U23464 (N_23464,N_23158,N_23121);
xor U23465 (N_23465,N_23052,N_23074);
nand U23466 (N_23466,N_23068,N_23177);
nand U23467 (N_23467,N_23193,N_23218);
and U23468 (N_23468,N_23106,N_23158);
or U23469 (N_23469,N_23043,N_23171);
xor U23470 (N_23470,N_23002,N_23175);
or U23471 (N_23471,N_23150,N_23061);
nor U23472 (N_23472,N_23068,N_23204);
or U23473 (N_23473,N_23222,N_23010);
and U23474 (N_23474,N_23056,N_23220);
and U23475 (N_23475,N_23004,N_23159);
or U23476 (N_23476,N_23091,N_23244);
nand U23477 (N_23477,N_23070,N_23049);
nor U23478 (N_23478,N_23168,N_23225);
and U23479 (N_23479,N_23144,N_23074);
xnor U23480 (N_23480,N_23195,N_23159);
nand U23481 (N_23481,N_23093,N_23080);
nand U23482 (N_23482,N_23239,N_23131);
nand U23483 (N_23483,N_23078,N_23074);
nor U23484 (N_23484,N_23064,N_23128);
or U23485 (N_23485,N_23210,N_23204);
nor U23486 (N_23486,N_23096,N_23121);
nand U23487 (N_23487,N_23164,N_23182);
or U23488 (N_23488,N_23128,N_23094);
and U23489 (N_23489,N_23116,N_23173);
or U23490 (N_23490,N_23100,N_23227);
nand U23491 (N_23491,N_23189,N_23095);
and U23492 (N_23492,N_23221,N_23064);
nand U23493 (N_23493,N_23083,N_23017);
nand U23494 (N_23494,N_23187,N_23194);
xor U23495 (N_23495,N_23197,N_23077);
nand U23496 (N_23496,N_23100,N_23080);
or U23497 (N_23497,N_23145,N_23095);
nand U23498 (N_23498,N_23144,N_23016);
nand U23499 (N_23499,N_23228,N_23019);
and U23500 (N_23500,N_23286,N_23371);
nand U23501 (N_23501,N_23261,N_23486);
or U23502 (N_23502,N_23414,N_23403);
nand U23503 (N_23503,N_23474,N_23341);
xor U23504 (N_23504,N_23287,N_23299);
and U23505 (N_23505,N_23460,N_23266);
or U23506 (N_23506,N_23492,N_23306);
nor U23507 (N_23507,N_23454,N_23320);
nor U23508 (N_23508,N_23356,N_23375);
nand U23509 (N_23509,N_23373,N_23305);
nand U23510 (N_23510,N_23459,N_23289);
nand U23511 (N_23511,N_23277,N_23465);
nand U23512 (N_23512,N_23444,N_23466);
nor U23513 (N_23513,N_23328,N_23340);
nor U23514 (N_23514,N_23360,N_23362);
nand U23515 (N_23515,N_23345,N_23260);
nor U23516 (N_23516,N_23411,N_23353);
and U23517 (N_23517,N_23409,N_23370);
nor U23518 (N_23518,N_23430,N_23386);
or U23519 (N_23519,N_23354,N_23379);
nand U23520 (N_23520,N_23359,N_23429);
nand U23521 (N_23521,N_23313,N_23272);
nand U23522 (N_23522,N_23480,N_23477);
nor U23523 (N_23523,N_23452,N_23327);
nor U23524 (N_23524,N_23269,N_23295);
nand U23525 (N_23525,N_23298,N_23268);
and U23526 (N_23526,N_23329,N_23488);
nand U23527 (N_23527,N_23445,N_23338);
nand U23528 (N_23528,N_23383,N_23424);
xor U23529 (N_23529,N_23257,N_23322);
nor U23530 (N_23530,N_23493,N_23254);
or U23531 (N_23531,N_23442,N_23302);
xor U23532 (N_23532,N_23263,N_23450);
nand U23533 (N_23533,N_23319,N_23363);
nand U23534 (N_23534,N_23326,N_23418);
xnor U23535 (N_23535,N_23361,N_23337);
and U23536 (N_23536,N_23250,N_23312);
and U23537 (N_23537,N_23355,N_23495);
and U23538 (N_23538,N_23453,N_23336);
or U23539 (N_23539,N_23273,N_23331);
nand U23540 (N_23540,N_23297,N_23404);
nor U23541 (N_23541,N_23315,N_23303);
xor U23542 (N_23542,N_23296,N_23292);
and U23543 (N_23543,N_23401,N_23334);
or U23544 (N_23544,N_23490,N_23389);
and U23545 (N_23545,N_23410,N_23441);
and U23546 (N_23546,N_23284,N_23256);
xnor U23547 (N_23547,N_23462,N_23432);
nand U23548 (N_23548,N_23300,N_23461);
or U23549 (N_23549,N_23397,N_23288);
and U23550 (N_23550,N_23449,N_23366);
or U23551 (N_23551,N_23275,N_23385);
xnor U23552 (N_23552,N_23267,N_23372);
xor U23553 (N_23553,N_23440,N_23309);
and U23554 (N_23554,N_23431,N_23482);
xor U23555 (N_23555,N_23475,N_23346);
xnor U23556 (N_23556,N_23464,N_23374);
and U23557 (N_23557,N_23252,N_23253);
nand U23558 (N_23558,N_23307,N_23467);
nor U23559 (N_23559,N_23378,N_23427);
or U23560 (N_23560,N_23262,N_23265);
or U23561 (N_23561,N_23343,N_23390);
nand U23562 (N_23562,N_23382,N_23405);
or U23563 (N_23563,N_23478,N_23434);
or U23564 (N_23564,N_23280,N_23476);
and U23565 (N_23565,N_23368,N_23443);
nor U23566 (N_23566,N_23412,N_23437);
or U23567 (N_23567,N_23487,N_23451);
or U23568 (N_23568,N_23350,N_23439);
nor U23569 (N_23569,N_23264,N_23285);
or U23570 (N_23570,N_23325,N_23447);
nor U23571 (N_23571,N_23351,N_23426);
nor U23572 (N_23572,N_23419,N_23310);
nand U23573 (N_23573,N_23259,N_23278);
or U23574 (N_23574,N_23271,N_23407);
nor U23575 (N_23575,N_23398,N_23408);
and U23576 (N_23576,N_23364,N_23330);
and U23577 (N_23577,N_23335,N_23416);
and U23578 (N_23578,N_23323,N_23406);
xor U23579 (N_23579,N_23294,N_23384);
nor U23580 (N_23580,N_23413,N_23469);
or U23581 (N_23581,N_23314,N_23352);
or U23582 (N_23582,N_23324,N_23396);
nor U23583 (N_23583,N_23470,N_23318);
or U23584 (N_23584,N_23483,N_23281);
and U23585 (N_23585,N_23436,N_23399);
or U23586 (N_23586,N_23494,N_23394);
nor U23587 (N_23587,N_23342,N_23463);
or U23588 (N_23588,N_23392,N_23433);
nor U23589 (N_23589,N_23317,N_23255);
nand U23590 (N_23590,N_23291,N_23428);
or U23591 (N_23591,N_23402,N_23489);
nand U23592 (N_23592,N_23311,N_23290);
nor U23593 (N_23593,N_23301,N_23455);
and U23594 (N_23594,N_23458,N_23283);
nand U23595 (N_23595,N_23400,N_23473);
nor U23596 (N_23596,N_23438,N_23456);
or U23597 (N_23597,N_23276,N_23472);
xnor U23598 (N_23598,N_23425,N_23274);
nand U23599 (N_23599,N_23422,N_23479);
xnor U23600 (N_23600,N_23393,N_23497);
nand U23601 (N_23601,N_23498,N_23258);
nand U23602 (N_23602,N_23332,N_23423);
nand U23603 (N_23603,N_23491,N_23421);
nand U23604 (N_23604,N_23484,N_23358);
nand U23605 (N_23605,N_23380,N_23446);
and U23606 (N_23606,N_23485,N_23499);
nor U23607 (N_23607,N_23282,N_23344);
nand U23608 (N_23608,N_23348,N_23349);
nor U23609 (N_23609,N_23308,N_23367);
and U23610 (N_23610,N_23365,N_23387);
xor U23611 (N_23611,N_23496,N_23381);
and U23612 (N_23612,N_23279,N_23377);
and U23613 (N_23613,N_23471,N_23468);
nand U23614 (N_23614,N_23251,N_23270);
nor U23615 (N_23615,N_23376,N_23391);
nor U23616 (N_23616,N_23357,N_23448);
or U23617 (N_23617,N_23457,N_23481);
nand U23618 (N_23618,N_23415,N_23369);
nor U23619 (N_23619,N_23339,N_23333);
nand U23620 (N_23620,N_23417,N_23321);
or U23621 (N_23621,N_23304,N_23293);
xnor U23622 (N_23622,N_23395,N_23388);
nor U23623 (N_23623,N_23435,N_23347);
or U23624 (N_23624,N_23420,N_23316);
xnor U23625 (N_23625,N_23314,N_23300);
xnor U23626 (N_23626,N_23294,N_23372);
and U23627 (N_23627,N_23383,N_23324);
xor U23628 (N_23628,N_23285,N_23353);
or U23629 (N_23629,N_23296,N_23315);
or U23630 (N_23630,N_23481,N_23468);
or U23631 (N_23631,N_23427,N_23254);
xnor U23632 (N_23632,N_23253,N_23496);
nand U23633 (N_23633,N_23403,N_23380);
and U23634 (N_23634,N_23412,N_23268);
nand U23635 (N_23635,N_23255,N_23493);
nor U23636 (N_23636,N_23406,N_23430);
xor U23637 (N_23637,N_23378,N_23471);
nor U23638 (N_23638,N_23412,N_23392);
nand U23639 (N_23639,N_23263,N_23466);
or U23640 (N_23640,N_23458,N_23464);
or U23641 (N_23641,N_23448,N_23287);
nand U23642 (N_23642,N_23401,N_23282);
nor U23643 (N_23643,N_23379,N_23416);
nand U23644 (N_23644,N_23338,N_23372);
nor U23645 (N_23645,N_23335,N_23472);
and U23646 (N_23646,N_23274,N_23340);
nand U23647 (N_23647,N_23314,N_23445);
nand U23648 (N_23648,N_23482,N_23383);
nor U23649 (N_23649,N_23256,N_23371);
nand U23650 (N_23650,N_23460,N_23371);
and U23651 (N_23651,N_23301,N_23335);
or U23652 (N_23652,N_23290,N_23364);
or U23653 (N_23653,N_23265,N_23485);
nor U23654 (N_23654,N_23368,N_23465);
nand U23655 (N_23655,N_23495,N_23332);
nand U23656 (N_23656,N_23498,N_23278);
nor U23657 (N_23657,N_23292,N_23454);
nor U23658 (N_23658,N_23354,N_23434);
and U23659 (N_23659,N_23432,N_23461);
xor U23660 (N_23660,N_23361,N_23289);
and U23661 (N_23661,N_23291,N_23298);
nor U23662 (N_23662,N_23483,N_23368);
and U23663 (N_23663,N_23437,N_23334);
xnor U23664 (N_23664,N_23439,N_23455);
and U23665 (N_23665,N_23365,N_23332);
nand U23666 (N_23666,N_23313,N_23284);
nand U23667 (N_23667,N_23467,N_23417);
and U23668 (N_23668,N_23421,N_23319);
and U23669 (N_23669,N_23464,N_23340);
and U23670 (N_23670,N_23287,N_23470);
xor U23671 (N_23671,N_23356,N_23317);
or U23672 (N_23672,N_23398,N_23285);
or U23673 (N_23673,N_23386,N_23428);
xor U23674 (N_23674,N_23338,N_23347);
nor U23675 (N_23675,N_23370,N_23284);
nor U23676 (N_23676,N_23313,N_23394);
or U23677 (N_23677,N_23459,N_23328);
nand U23678 (N_23678,N_23482,N_23441);
nor U23679 (N_23679,N_23402,N_23297);
and U23680 (N_23680,N_23255,N_23316);
xor U23681 (N_23681,N_23457,N_23262);
and U23682 (N_23682,N_23453,N_23340);
nand U23683 (N_23683,N_23318,N_23368);
xor U23684 (N_23684,N_23259,N_23370);
nor U23685 (N_23685,N_23440,N_23346);
nor U23686 (N_23686,N_23272,N_23277);
nor U23687 (N_23687,N_23438,N_23397);
or U23688 (N_23688,N_23357,N_23404);
or U23689 (N_23689,N_23320,N_23325);
and U23690 (N_23690,N_23254,N_23417);
and U23691 (N_23691,N_23461,N_23453);
or U23692 (N_23692,N_23324,N_23453);
and U23693 (N_23693,N_23396,N_23419);
and U23694 (N_23694,N_23443,N_23332);
nor U23695 (N_23695,N_23408,N_23291);
xor U23696 (N_23696,N_23348,N_23265);
nand U23697 (N_23697,N_23358,N_23370);
xnor U23698 (N_23698,N_23309,N_23471);
or U23699 (N_23699,N_23404,N_23294);
and U23700 (N_23700,N_23324,N_23290);
and U23701 (N_23701,N_23285,N_23346);
and U23702 (N_23702,N_23316,N_23484);
nor U23703 (N_23703,N_23344,N_23290);
nand U23704 (N_23704,N_23302,N_23292);
or U23705 (N_23705,N_23410,N_23316);
nand U23706 (N_23706,N_23408,N_23481);
or U23707 (N_23707,N_23352,N_23460);
or U23708 (N_23708,N_23352,N_23484);
xor U23709 (N_23709,N_23393,N_23433);
and U23710 (N_23710,N_23263,N_23463);
or U23711 (N_23711,N_23395,N_23260);
or U23712 (N_23712,N_23406,N_23401);
and U23713 (N_23713,N_23312,N_23360);
nand U23714 (N_23714,N_23463,N_23391);
and U23715 (N_23715,N_23391,N_23403);
nor U23716 (N_23716,N_23438,N_23320);
xor U23717 (N_23717,N_23285,N_23445);
and U23718 (N_23718,N_23326,N_23492);
xnor U23719 (N_23719,N_23449,N_23346);
nor U23720 (N_23720,N_23289,N_23323);
and U23721 (N_23721,N_23269,N_23474);
nand U23722 (N_23722,N_23397,N_23395);
or U23723 (N_23723,N_23441,N_23444);
xor U23724 (N_23724,N_23324,N_23404);
nor U23725 (N_23725,N_23446,N_23253);
and U23726 (N_23726,N_23460,N_23476);
nor U23727 (N_23727,N_23364,N_23433);
nand U23728 (N_23728,N_23279,N_23349);
nand U23729 (N_23729,N_23313,N_23385);
xor U23730 (N_23730,N_23267,N_23432);
or U23731 (N_23731,N_23463,N_23421);
xnor U23732 (N_23732,N_23452,N_23282);
nor U23733 (N_23733,N_23405,N_23270);
or U23734 (N_23734,N_23473,N_23494);
or U23735 (N_23735,N_23447,N_23379);
and U23736 (N_23736,N_23366,N_23265);
xor U23737 (N_23737,N_23355,N_23384);
or U23738 (N_23738,N_23491,N_23469);
nor U23739 (N_23739,N_23280,N_23335);
or U23740 (N_23740,N_23387,N_23260);
or U23741 (N_23741,N_23283,N_23480);
nor U23742 (N_23742,N_23292,N_23318);
or U23743 (N_23743,N_23376,N_23324);
nand U23744 (N_23744,N_23361,N_23314);
xor U23745 (N_23745,N_23401,N_23388);
or U23746 (N_23746,N_23433,N_23312);
or U23747 (N_23747,N_23477,N_23374);
xor U23748 (N_23748,N_23361,N_23325);
nand U23749 (N_23749,N_23312,N_23422);
or U23750 (N_23750,N_23615,N_23505);
nor U23751 (N_23751,N_23739,N_23700);
nor U23752 (N_23752,N_23648,N_23634);
xnor U23753 (N_23753,N_23629,N_23545);
nor U23754 (N_23754,N_23542,N_23692);
or U23755 (N_23755,N_23562,N_23567);
or U23756 (N_23756,N_23506,N_23660);
or U23757 (N_23757,N_23585,N_23541);
nor U23758 (N_23758,N_23680,N_23738);
or U23759 (N_23759,N_23544,N_23716);
nand U23760 (N_23760,N_23713,N_23695);
or U23761 (N_23761,N_23651,N_23569);
nand U23762 (N_23762,N_23656,N_23726);
and U23763 (N_23763,N_23743,N_23608);
nor U23764 (N_23764,N_23635,N_23500);
nand U23765 (N_23765,N_23637,N_23558);
and U23766 (N_23766,N_23714,N_23661);
nor U23767 (N_23767,N_23535,N_23578);
and U23768 (N_23768,N_23669,N_23598);
nor U23769 (N_23769,N_23691,N_23625);
or U23770 (N_23770,N_23742,N_23630);
xnor U23771 (N_23771,N_23554,N_23559);
and U23772 (N_23772,N_23626,N_23737);
nor U23773 (N_23773,N_23612,N_23747);
nor U23774 (N_23774,N_23540,N_23606);
nor U23775 (N_23775,N_23686,N_23592);
or U23776 (N_23776,N_23621,N_23677);
and U23777 (N_23777,N_23657,N_23574);
and U23778 (N_23778,N_23633,N_23572);
nor U23779 (N_23779,N_23610,N_23557);
nor U23780 (N_23780,N_23520,N_23519);
or U23781 (N_23781,N_23719,N_23591);
or U23782 (N_23782,N_23674,N_23539);
or U23783 (N_23783,N_23683,N_23525);
nand U23784 (N_23784,N_23576,N_23720);
and U23785 (N_23785,N_23673,N_23706);
or U23786 (N_23786,N_23516,N_23590);
and U23787 (N_23787,N_23746,N_23518);
xnor U23788 (N_23788,N_23509,N_23701);
xnor U23789 (N_23789,N_23676,N_23698);
nor U23790 (N_23790,N_23556,N_23528);
nor U23791 (N_23791,N_23687,N_23532);
nand U23792 (N_23792,N_23573,N_23584);
and U23793 (N_23793,N_23580,N_23718);
nor U23794 (N_23794,N_23607,N_23512);
xnor U23795 (N_23795,N_23546,N_23605);
or U23796 (N_23796,N_23594,N_23555);
xor U23797 (N_23797,N_23721,N_23667);
or U23798 (N_23798,N_23543,N_23589);
xor U23799 (N_23799,N_23632,N_23678);
or U23800 (N_23800,N_23704,N_23647);
and U23801 (N_23801,N_23568,N_23502);
nand U23802 (N_23802,N_23552,N_23577);
or U23803 (N_23803,N_23586,N_23507);
xor U23804 (N_23804,N_23534,N_23614);
and U23805 (N_23805,N_23732,N_23665);
or U23806 (N_23806,N_23530,N_23570);
and U23807 (N_23807,N_23553,N_23703);
nand U23808 (N_23808,N_23641,N_23616);
and U23809 (N_23809,N_23697,N_23638);
nand U23810 (N_23810,N_23510,N_23728);
and U23811 (N_23811,N_23644,N_23645);
nand U23812 (N_23812,N_23699,N_23508);
nand U23813 (N_23813,N_23531,N_23688);
or U23814 (N_23814,N_23653,N_23603);
or U23815 (N_23815,N_23550,N_23702);
xor U23816 (N_23816,N_23740,N_23731);
and U23817 (N_23817,N_23551,N_23654);
or U23818 (N_23818,N_23682,N_23547);
nand U23819 (N_23819,N_23566,N_23596);
and U23820 (N_23820,N_23636,N_23609);
nand U23821 (N_23821,N_23521,N_23602);
xor U23822 (N_23822,N_23622,N_23563);
nor U23823 (N_23823,N_23613,N_23748);
and U23824 (N_23824,N_23684,N_23696);
or U23825 (N_23825,N_23708,N_23565);
or U23826 (N_23826,N_23689,N_23575);
or U23827 (N_23827,N_23623,N_23735);
or U23828 (N_23828,N_23724,N_23593);
or U23829 (N_23829,N_23723,N_23522);
nand U23830 (N_23830,N_23620,N_23581);
xor U23831 (N_23831,N_23685,N_23549);
or U23832 (N_23832,N_23529,N_23655);
nor U23833 (N_23833,N_23643,N_23733);
nor U23834 (N_23834,N_23707,N_23631);
and U23835 (N_23835,N_23600,N_23741);
and U23836 (N_23836,N_23599,N_23517);
nor U23837 (N_23837,N_23611,N_23675);
or U23838 (N_23838,N_23712,N_23668);
nor U23839 (N_23839,N_23659,N_23514);
xor U23840 (N_23840,N_23734,N_23639);
and U23841 (N_23841,N_23670,N_23715);
and U23842 (N_23842,N_23717,N_23736);
xor U23843 (N_23843,N_23503,N_23548);
xnor U23844 (N_23844,N_23501,N_23564);
nand U23845 (N_23845,N_23640,N_23662);
nor U23846 (N_23846,N_23601,N_23694);
nand U23847 (N_23847,N_23536,N_23526);
nor U23848 (N_23848,N_23561,N_23730);
and U23849 (N_23849,N_23646,N_23666);
nand U23850 (N_23850,N_23711,N_23729);
xor U23851 (N_23851,N_23504,N_23537);
nand U23852 (N_23852,N_23523,N_23527);
nand U23853 (N_23853,N_23745,N_23727);
xnor U23854 (N_23854,N_23511,N_23587);
nor U23855 (N_23855,N_23652,N_23560);
or U23856 (N_23856,N_23690,N_23533);
and U23857 (N_23857,N_23588,N_23617);
xnor U23858 (N_23858,N_23604,N_23658);
xnor U23859 (N_23859,N_23725,N_23642);
or U23860 (N_23860,N_23664,N_23649);
nand U23861 (N_23861,N_23628,N_23710);
or U23862 (N_23862,N_23579,N_23650);
nor U23863 (N_23863,N_23513,N_23671);
and U23864 (N_23864,N_23571,N_23627);
nand U23865 (N_23865,N_23681,N_23582);
xor U23866 (N_23866,N_23595,N_23515);
or U23867 (N_23867,N_23679,N_23722);
xnor U23868 (N_23868,N_23619,N_23663);
and U23869 (N_23869,N_23583,N_23744);
nand U23870 (N_23870,N_23672,N_23597);
and U23871 (N_23871,N_23618,N_23624);
and U23872 (N_23872,N_23749,N_23524);
nand U23873 (N_23873,N_23709,N_23693);
xor U23874 (N_23874,N_23705,N_23538);
nor U23875 (N_23875,N_23528,N_23517);
or U23876 (N_23876,N_23652,N_23621);
xnor U23877 (N_23877,N_23542,N_23739);
nor U23878 (N_23878,N_23548,N_23516);
nor U23879 (N_23879,N_23522,N_23717);
nand U23880 (N_23880,N_23749,N_23616);
nor U23881 (N_23881,N_23742,N_23679);
or U23882 (N_23882,N_23606,N_23515);
nand U23883 (N_23883,N_23576,N_23673);
or U23884 (N_23884,N_23704,N_23501);
and U23885 (N_23885,N_23591,N_23741);
xnor U23886 (N_23886,N_23680,N_23555);
xor U23887 (N_23887,N_23504,N_23638);
nand U23888 (N_23888,N_23592,N_23594);
nand U23889 (N_23889,N_23643,N_23689);
and U23890 (N_23890,N_23618,N_23632);
nor U23891 (N_23891,N_23657,N_23581);
or U23892 (N_23892,N_23619,N_23735);
nand U23893 (N_23893,N_23613,N_23614);
or U23894 (N_23894,N_23520,N_23536);
or U23895 (N_23895,N_23557,N_23626);
nand U23896 (N_23896,N_23537,N_23510);
or U23897 (N_23897,N_23702,N_23732);
nand U23898 (N_23898,N_23580,N_23647);
or U23899 (N_23899,N_23651,N_23723);
nor U23900 (N_23900,N_23565,N_23681);
and U23901 (N_23901,N_23695,N_23557);
nand U23902 (N_23902,N_23524,N_23511);
xor U23903 (N_23903,N_23652,N_23581);
xor U23904 (N_23904,N_23684,N_23660);
or U23905 (N_23905,N_23505,N_23506);
and U23906 (N_23906,N_23685,N_23735);
and U23907 (N_23907,N_23562,N_23733);
nor U23908 (N_23908,N_23695,N_23618);
and U23909 (N_23909,N_23676,N_23671);
xor U23910 (N_23910,N_23700,N_23589);
or U23911 (N_23911,N_23528,N_23657);
or U23912 (N_23912,N_23697,N_23673);
xnor U23913 (N_23913,N_23561,N_23642);
and U23914 (N_23914,N_23686,N_23518);
and U23915 (N_23915,N_23555,N_23671);
and U23916 (N_23916,N_23728,N_23607);
and U23917 (N_23917,N_23523,N_23592);
and U23918 (N_23918,N_23543,N_23652);
and U23919 (N_23919,N_23657,N_23538);
nor U23920 (N_23920,N_23597,N_23511);
and U23921 (N_23921,N_23589,N_23533);
or U23922 (N_23922,N_23577,N_23649);
xor U23923 (N_23923,N_23630,N_23627);
and U23924 (N_23924,N_23525,N_23564);
nand U23925 (N_23925,N_23521,N_23520);
xor U23926 (N_23926,N_23695,N_23520);
nand U23927 (N_23927,N_23515,N_23508);
or U23928 (N_23928,N_23539,N_23658);
xnor U23929 (N_23929,N_23555,N_23740);
or U23930 (N_23930,N_23506,N_23653);
or U23931 (N_23931,N_23634,N_23687);
nor U23932 (N_23932,N_23709,N_23597);
xnor U23933 (N_23933,N_23520,N_23661);
nor U23934 (N_23934,N_23520,N_23606);
or U23935 (N_23935,N_23624,N_23659);
xor U23936 (N_23936,N_23633,N_23721);
or U23937 (N_23937,N_23589,N_23667);
or U23938 (N_23938,N_23634,N_23643);
nor U23939 (N_23939,N_23653,N_23607);
xnor U23940 (N_23940,N_23674,N_23601);
nand U23941 (N_23941,N_23748,N_23569);
and U23942 (N_23942,N_23686,N_23675);
nor U23943 (N_23943,N_23667,N_23585);
or U23944 (N_23944,N_23666,N_23509);
or U23945 (N_23945,N_23629,N_23736);
nor U23946 (N_23946,N_23671,N_23631);
and U23947 (N_23947,N_23561,N_23704);
nand U23948 (N_23948,N_23633,N_23682);
or U23949 (N_23949,N_23746,N_23526);
and U23950 (N_23950,N_23604,N_23719);
nand U23951 (N_23951,N_23713,N_23582);
nor U23952 (N_23952,N_23645,N_23656);
or U23953 (N_23953,N_23557,N_23600);
xor U23954 (N_23954,N_23575,N_23567);
xor U23955 (N_23955,N_23521,N_23685);
and U23956 (N_23956,N_23668,N_23591);
nand U23957 (N_23957,N_23501,N_23552);
nor U23958 (N_23958,N_23631,N_23501);
nor U23959 (N_23959,N_23627,N_23632);
nand U23960 (N_23960,N_23601,N_23608);
nor U23961 (N_23961,N_23692,N_23703);
xor U23962 (N_23962,N_23559,N_23652);
or U23963 (N_23963,N_23518,N_23564);
nand U23964 (N_23964,N_23553,N_23595);
xnor U23965 (N_23965,N_23569,N_23550);
or U23966 (N_23966,N_23714,N_23567);
nor U23967 (N_23967,N_23562,N_23594);
and U23968 (N_23968,N_23517,N_23593);
nand U23969 (N_23969,N_23590,N_23549);
or U23970 (N_23970,N_23538,N_23632);
nor U23971 (N_23971,N_23669,N_23667);
nand U23972 (N_23972,N_23671,N_23608);
xnor U23973 (N_23973,N_23702,N_23506);
nor U23974 (N_23974,N_23721,N_23583);
nand U23975 (N_23975,N_23666,N_23547);
nor U23976 (N_23976,N_23567,N_23512);
nand U23977 (N_23977,N_23665,N_23735);
or U23978 (N_23978,N_23678,N_23604);
xor U23979 (N_23979,N_23668,N_23715);
nor U23980 (N_23980,N_23610,N_23670);
and U23981 (N_23981,N_23692,N_23623);
xor U23982 (N_23982,N_23684,N_23605);
xor U23983 (N_23983,N_23582,N_23530);
xnor U23984 (N_23984,N_23612,N_23645);
nand U23985 (N_23985,N_23531,N_23683);
and U23986 (N_23986,N_23634,N_23613);
nor U23987 (N_23987,N_23579,N_23583);
and U23988 (N_23988,N_23688,N_23525);
nand U23989 (N_23989,N_23667,N_23743);
nor U23990 (N_23990,N_23543,N_23512);
and U23991 (N_23991,N_23713,N_23623);
xor U23992 (N_23992,N_23601,N_23580);
and U23993 (N_23993,N_23619,N_23726);
and U23994 (N_23994,N_23513,N_23635);
xnor U23995 (N_23995,N_23538,N_23607);
nor U23996 (N_23996,N_23583,N_23651);
nor U23997 (N_23997,N_23678,N_23713);
or U23998 (N_23998,N_23718,N_23732);
nand U23999 (N_23999,N_23571,N_23714);
nor U24000 (N_24000,N_23959,N_23781);
nor U24001 (N_24001,N_23810,N_23870);
nor U24002 (N_24002,N_23878,N_23981);
or U24003 (N_24003,N_23835,N_23825);
xnor U24004 (N_24004,N_23945,N_23924);
or U24005 (N_24005,N_23960,N_23951);
xor U24006 (N_24006,N_23844,N_23907);
nor U24007 (N_24007,N_23950,N_23982);
nand U24008 (N_24008,N_23956,N_23866);
or U24009 (N_24009,N_23886,N_23839);
nor U24010 (N_24010,N_23799,N_23890);
nand U24011 (N_24011,N_23805,N_23979);
nand U24012 (N_24012,N_23840,N_23916);
xor U24013 (N_24013,N_23988,N_23853);
or U24014 (N_24014,N_23824,N_23797);
nand U24015 (N_24015,N_23875,N_23763);
nand U24016 (N_24016,N_23789,N_23996);
and U24017 (N_24017,N_23784,N_23817);
and U24018 (N_24018,N_23782,N_23926);
or U24019 (N_24019,N_23814,N_23934);
nor U24020 (N_24020,N_23938,N_23813);
nand U24021 (N_24021,N_23929,N_23828);
nand U24022 (N_24022,N_23859,N_23874);
and U24023 (N_24023,N_23928,N_23761);
nand U24024 (N_24024,N_23837,N_23957);
nor U24025 (N_24025,N_23823,N_23937);
nand U24026 (N_24026,N_23752,N_23885);
xnor U24027 (N_24027,N_23983,N_23976);
or U24028 (N_24028,N_23990,N_23949);
nand U24029 (N_24029,N_23834,N_23992);
and U24030 (N_24030,N_23766,N_23922);
nor U24031 (N_24031,N_23857,N_23898);
nor U24032 (N_24032,N_23940,N_23863);
nor U24033 (N_24033,N_23794,N_23822);
xor U24034 (N_24034,N_23793,N_23917);
xor U24035 (N_24035,N_23830,N_23942);
xnor U24036 (N_24036,N_23903,N_23865);
or U24037 (N_24037,N_23787,N_23849);
nand U24038 (N_24038,N_23827,N_23754);
nand U24039 (N_24039,N_23927,N_23902);
nor U24040 (N_24040,N_23963,N_23759);
and U24041 (N_24041,N_23894,N_23993);
xor U24042 (N_24042,N_23967,N_23795);
or U24043 (N_24043,N_23977,N_23848);
nor U24044 (N_24044,N_23798,N_23913);
nor U24045 (N_24045,N_23932,N_23912);
or U24046 (N_24046,N_23832,N_23775);
xor U24047 (N_24047,N_23931,N_23770);
nand U24048 (N_24048,N_23884,N_23774);
xor U24049 (N_24049,N_23920,N_23887);
nor U24050 (N_24050,N_23838,N_23842);
xor U24051 (N_24051,N_23802,N_23829);
nand U24052 (N_24052,N_23820,N_23773);
and U24053 (N_24053,N_23964,N_23883);
nand U24054 (N_24054,N_23851,N_23779);
nand U24055 (N_24055,N_23955,N_23850);
xor U24056 (N_24056,N_23944,N_23783);
xor U24057 (N_24057,N_23984,N_23915);
and U24058 (N_24058,N_23987,N_23991);
xnor U24059 (N_24059,N_23941,N_23879);
xor U24060 (N_24060,N_23757,N_23873);
or U24061 (N_24061,N_23925,N_23896);
nand U24062 (N_24062,N_23943,N_23997);
nand U24063 (N_24063,N_23919,N_23900);
nor U24064 (N_24064,N_23998,N_23847);
nand U24065 (N_24065,N_23762,N_23792);
nand U24066 (N_24066,N_23891,N_23860);
and U24067 (N_24067,N_23804,N_23897);
nor U24068 (N_24068,N_23901,N_23858);
and U24069 (N_24069,N_23867,N_23816);
nand U24070 (N_24070,N_23953,N_23769);
nand U24071 (N_24071,N_23871,N_23936);
nand U24072 (N_24072,N_23765,N_23809);
or U24073 (N_24073,N_23961,N_23877);
and U24074 (N_24074,N_23994,N_23876);
or U24075 (N_24075,N_23948,N_23930);
and U24076 (N_24076,N_23845,N_23999);
or U24077 (N_24077,N_23826,N_23753);
nand U24078 (N_24078,N_23771,N_23911);
or U24079 (N_24079,N_23852,N_23946);
nor U24080 (N_24080,N_23975,N_23764);
nand U24081 (N_24081,N_23815,N_23755);
nand U24082 (N_24082,N_23855,N_23785);
and U24083 (N_24083,N_23864,N_23807);
and U24084 (N_24084,N_23846,N_23889);
or U24085 (N_24085,N_23880,N_23954);
or U24086 (N_24086,N_23767,N_23856);
nor U24087 (N_24087,N_23899,N_23972);
xor U24088 (N_24088,N_23918,N_23808);
nand U24089 (N_24089,N_23868,N_23908);
and U24090 (N_24090,N_23862,N_23966);
xnor U24091 (N_24091,N_23973,N_23935);
xnor U24092 (N_24092,N_23892,N_23818);
and U24093 (N_24093,N_23962,N_23843);
or U24094 (N_24094,N_23751,N_23872);
xnor U24095 (N_24095,N_23786,N_23811);
and U24096 (N_24096,N_23882,N_23906);
nor U24097 (N_24097,N_23970,N_23978);
xnor U24098 (N_24098,N_23939,N_23952);
xor U24099 (N_24099,N_23888,N_23947);
and U24100 (N_24100,N_23758,N_23772);
nand U24101 (N_24101,N_23923,N_23833);
or U24102 (N_24102,N_23760,N_23971);
nor U24103 (N_24103,N_23777,N_23780);
nand U24104 (N_24104,N_23895,N_23914);
nand U24105 (N_24105,N_23788,N_23841);
or U24106 (N_24106,N_23756,N_23995);
nand U24107 (N_24107,N_23831,N_23989);
nor U24108 (N_24108,N_23986,N_23909);
nor U24109 (N_24109,N_23958,N_23910);
nor U24110 (N_24110,N_23974,N_23980);
and U24111 (N_24111,N_23968,N_23933);
nor U24112 (N_24112,N_23803,N_23893);
and U24113 (N_24113,N_23791,N_23750);
and U24114 (N_24114,N_23790,N_23768);
xnor U24115 (N_24115,N_23796,N_23921);
nand U24116 (N_24116,N_23836,N_23778);
and U24117 (N_24117,N_23969,N_23861);
nand U24118 (N_24118,N_23819,N_23905);
nor U24119 (N_24119,N_23812,N_23965);
or U24120 (N_24120,N_23881,N_23800);
or U24121 (N_24121,N_23806,N_23904);
or U24122 (N_24122,N_23985,N_23869);
nor U24123 (N_24123,N_23821,N_23776);
and U24124 (N_24124,N_23801,N_23854);
xor U24125 (N_24125,N_23872,N_23834);
nand U24126 (N_24126,N_23850,N_23838);
and U24127 (N_24127,N_23801,N_23783);
xor U24128 (N_24128,N_23865,N_23863);
nand U24129 (N_24129,N_23878,N_23818);
nand U24130 (N_24130,N_23953,N_23753);
nor U24131 (N_24131,N_23955,N_23797);
nor U24132 (N_24132,N_23837,N_23778);
xor U24133 (N_24133,N_23954,N_23928);
xor U24134 (N_24134,N_23801,N_23786);
nor U24135 (N_24135,N_23998,N_23928);
or U24136 (N_24136,N_23847,N_23769);
xnor U24137 (N_24137,N_23996,N_23791);
or U24138 (N_24138,N_23794,N_23932);
nor U24139 (N_24139,N_23864,N_23911);
nor U24140 (N_24140,N_23978,N_23780);
nor U24141 (N_24141,N_23988,N_23776);
xor U24142 (N_24142,N_23973,N_23824);
xnor U24143 (N_24143,N_23944,N_23912);
xnor U24144 (N_24144,N_23821,N_23789);
or U24145 (N_24145,N_23853,N_23795);
nor U24146 (N_24146,N_23802,N_23918);
nor U24147 (N_24147,N_23867,N_23905);
nor U24148 (N_24148,N_23941,N_23974);
and U24149 (N_24149,N_23912,N_23780);
and U24150 (N_24150,N_23865,N_23765);
xor U24151 (N_24151,N_23974,N_23949);
or U24152 (N_24152,N_23926,N_23868);
and U24153 (N_24153,N_23880,N_23885);
xor U24154 (N_24154,N_23860,N_23915);
or U24155 (N_24155,N_23877,N_23946);
nand U24156 (N_24156,N_23888,N_23982);
nand U24157 (N_24157,N_23753,N_23767);
nand U24158 (N_24158,N_23988,N_23803);
nand U24159 (N_24159,N_23759,N_23865);
xnor U24160 (N_24160,N_23956,N_23787);
or U24161 (N_24161,N_23888,N_23977);
and U24162 (N_24162,N_23933,N_23863);
nand U24163 (N_24163,N_23791,N_23936);
nor U24164 (N_24164,N_23832,N_23985);
or U24165 (N_24165,N_23983,N_23918);
nand U24166 (N_24166,N_23949,N_23957);
nor U24167 (N_24167,N_23881,N_23815);
nor U24168 (N_24168,N_23841,N_23758);
nor U24169 (N_24169,N_23789,N_23933);
xnor U24170 (N_24170,N_23813,N_23951);
or U24171 (N_24171,N_23776,N_23970);
nor U24172 (N_24172,N_23869,N_23862);
nand U24173 (N_24173,N_23829,N_23855);
nand U24174 (N_24174,N_23989,N_23775);
and U24175 (N_24175,N_23960,N_23876);
or U24176 (N_24176,N_23789,N_23800);
and U24177 (N_24177,N_23816,N_23841);
or U24178 (N_24178,N_23993,N_23896);
and U24179 (N_24179,N_23758,N_23930);
xnor U24180 (N_24180,N_23899,N_23942);
xnor U24181 (N_24181,N_23777,N_23965);
nand U24182 (N_24182,N_23866,N_23881);
and U24183 (N_24183,N_23875,N_23780);
nand U24184 (N_24184,N_23785,N_23949);
nor U24185 (N_24185,N_23929,N_23877);
and U24186 (N_24186,N_23888,N_23859);
xnor U24187 (N_24187,N_23872,N_23832);
or U24188 (N_24188,N_23922,N_23772);
and U24189 (N_24189,N_23881,N_23963);
or U24190 (N_24190,N_23926,N_23989);
or U24191 (N_24191,N_23909,N_23833);
or U24192 (N_24192,N_23792,N_23773);
xor U24193 (N_24193,N_23867,N_23755);
nor U24194 (N_24194,N_23934,N_23819);
or U24195 (N_24195,N_23987,N_23951);
or U24196 (N_24196,N_23765,N_23855);
and U24197 (N_24197,N_23948,N_23945);
nor U24198 (N_24198,N_23875,N_23953);
nand U24199 (N_24199,N_23996,N_23796);
and U24200 (N_24200,N_23838,N_23919);
xor U24201 (N_24201,N_23832,N_23752);
or U24202 (N_24202,N_23781,N_23772);
and U24203 (N_24203,N_23794,N_23893);
and U24204 (N_24204,N_23765,N_23904);
nor U24205 (N_24205,N_23940,N_23859);
or U24206 (N_24206,N_23966,N_23995);
xor U24207 (N_24207,N_23985,N_23891);
nand U24208 (N_24208,N_23868,N_23756);
nand U24209 (N_24209,N_23859,N_23831);
nand U24210 (N_24210,N_23925,N_23879);
nor U24211 (N_24211,N_23766,N_23831);
xor U24212 (N_24212,N_23886,N_23797);
nor U24213 (N_24213,N_23752,N_23972);
nor U24214 (N_24214,N_23754,N_23800);
nand U24215 (N_24215,N_23945,N_23953);
or U24216 (N_24216,N_23870,N_23777);
nand U24217 (N_24217,N_23969,N_23808);
and U24218 (N_24218,N_23999,N_23775);
or U24219 (N_24219,N_23999,N_23793);
nand U24220 (N_24220,N_23921,N_23901);
nor U24221 (N_24221,N_23848,N_23967);
xnor U24222 (N_24222,N_23868,N_23915);
nor U24223 (N_24223,N_23846,N_23931);
and U24224 (N_24224,N_23847,N_23891);
and U24225 (N_24225,N_23984,N_23924);
nand U24226 (N_24226,N_23794,N_23964);
and U24227 (N_24227,N_23778,N_23843);
nor U24228 (N_24228,N_23801,N_23972);
or U24229 (N_24229,N_23820,N_23770);
and U24230 (N_24230,N_23779,N_23945);
or U24231 (N_24231,N_23885,N_23787);
nor U24232 (N_24232,N_23960,N_23821);
and U24233 (N_24233,N_23963,N_23791);
nand U24234 (N_24234,N_23756,N_23838);
and U24235 (N_24235,N_23887,N_23816);
and U24236 (N_24236,N_23915,N_23809);
or U24237 (N_24237,N_23786,N_23952);
or U24238 (N_24238,N_23820,N_23757);
nor U24239 (N_24239,N_23782,N_23834);
and U24240 (N_24240,N_23831,N_23968);
and U24241 (N_24241,N_23783,N_23787);
and U24242 (N_24242,N_23775,N_23835);
xnor U24243 (N_24243,N_23966,N_23894);
or U24244 (N_24244,N_23890,N_23993);
xnor U24245 (N_24245,N_23794,N_23779);
nor U24246 (N_24246,N_23878,N_23811);
nor U24247 (N_24247,N_23864,N_23890);
and U24248 (N_24248,N_23903,N_23831);
or U24249 (N_24249,N_23940,N_23882);
nor U24250 (N_24250,N_24200,N_24073);
nor U24251 (N_24251,N_24238,N_24030);
or U24252 (N_24252,N_24131,N_24235);
and U24253 (N_24253,N_24080,N_24094);
or U24254 (N_24254,N_24075,N_24015);
or U24255 (N_24255,N_24069,N_24142);
nor U24256 (N_24256,N_24156,N_24204);
or U24257 (N_24257,N_24019,N_24231);
xor U24258 (N_24258,N_24000,N_24010);
or U24259 (N_24259,N_24249,N_24039);
xor U24260 (N_24260,N_24117,N_24097);
nand U24261 (N_24261,N_24038,N_24008);
xor U24262 (N_24262,N_24182,N_24107);
and U24263 (N_24263,N_24222,N_24183);
nand U24264 (N_24264,N_24018,N_24140);
xor U24265 (N_24265,N_24060,N_24158);
or U24266 (N_24266,N_24221,N_24091);
or U24267 (N_24267,N_24164,N_24198);
or U24268 (N_24268,N_24079,N_24001);
nand U24269 (N_24269,N_24227,N_24224);
nor U24270 (N_24270,N_24064,N_24102);
xor U24271 (N_24271,N_24218,N_24003);
xnor U24272 (N_24272,N_24034,N_24111);
and U24273 (N_24273,N_24212,N_24004);
or U24274 (N_24274,N_24192,N_24247);
or U24275 (N_24275,N_24155,N_24240);
xnor U24276 (N_24276,N_24110,N_24220);
nor U24277 (N_24277,N_24052,N_24225);
nor U24278 (N_24278,N_24207,N_24245);
and U24279 (N_24279,N_24096,N_24209);
or U24280 (N_24280,N_24127,N_24202);
xnor U24281 (N_24281,N_24159,N_24049);
nor U24282 (N_24282,N_24063,N_24042);
or U24283 (N_24283,N_24172,N_24241);
or U24284 (N_24284,N_24006,N_24233);
nor U24285 (N_24285,N_24068,N_24154);
nand U24286 (N_24286,N_24028,N_24051);
xor U24287 (N_24287,N_24002,N_24187);
and U24288 (N_24288,N_24136,N_24208);
nor U24289 (N_24289,N_24074,N_24070);
or U24290 (N_24290,N_24134,N_24032);
and U24291 (N_24291,N_24114,N_24011);
xor U24292 (N_24292,N_24116,N_24168);
nand U24293 (N_24293,N_24223,N_24062);
or U24294 (N_24294,N_24082,N_24165);
or U24295 (N_24295,N_24184,N_24016);
nor U24296 (N_24296,N_24242,N_24054);
nor U24297 (N_24297,N_24099,N_24174);
or U24298 (N_24298,N_24029,N_24175);
or U24299 (N_24299,N_24194,N_24141);
and U24300 (N_24300,N_24146,N_24139);
and U24301 (N_24301,N_24193,N_24021);
and U24302 (N_24302,N_24213,N_24128);
nor U24303 (N_24303,N_24076,N_24186);
or U24304 (N_24304,N_24033,N_24169);
nand U24305 (N_24305,N_24157,N_24118);
nand U24306 (N_24306,N_24196,N_24173);
xor U24307 (N_24307,N_24210,N_24057);
xor U24308 (N_24308,N_24205,N_24066);
or U24309 (N_24309,N_24103,N_24031);
and U24310 (N_24310,N_24059,N_24126);
and U24311 (N_24311,N_24077,N_24053);
xnor U24312 (N_24312,N_24177,N_24124);
xor U24313 (N_24313,N_24211,N_24226);
xnor U24314 (N_24314,N_24190,N_24244);
xnor U24315 (N_24315,N_24214,N_24129);
nand U24316 (N_24316,N_24152,N_24151);
or U24317 (N_24317,N_24147,N_24228);
and U24318 (N_24318,N_24093,N_24012);
or U24319 (N_24319,N_24014,N_24009);
nor U24320 (N_24320,N_24206,N_24181);
and U24321 (N_24321,N_24007,N_24027);
xnor U24322 (N_24322,N_24170,N_24067);
or U24323 (N_24323,N_24125,N_24232);
and U24324 (N_24324,N_24098,N_24092);
and U24325 (N_24325,N_24148,N_24189);
and U24326 (N_24326,N_24041,N_24120);
nor U24327 (N_24327,N_24217,N_24132);
nand U24328 (N_24328,N_24239,N_24215);
or U24329 (N_24329,N_24121,N_24088);
xnor U24330 (N_24330,N_24043,N_24026);
nor U24331 (N_24331,N_24101,N_24203);
nand U24332 (N_24332,N_24237,N_24044);
nand U24333 (N_24333,N_24234,N_24106);
xor U24334 (N_24334,N_24023,N_24176);
xor U24335 (N_24335,N_24145,N_24149);
and U24336 (N_24336,N_24085,N_24071);
and U24337 (N_24337,N_24119,N_24188);
and U24338 (N_24338,N_24115,N_24072);
nor U24339 (N_24339,N_24166,N_24086);
nand U24340 (N_24340,N_24020,N_24078);
nor U24341 (N_24341,N_24100,N_24083);
xnor U24342 (N_24342,N_24179,N_24095);
and U24343 (N_24343,N_24195,N_24122);
nor U24344 (N_24344,N_24047,N_24138);
and U24345 (N_24345,N_24236,N_24229);
nor U24346 (N_24346,N_24037,N_24199);
or U24347 (N_24347,N_24036,N_24035);
and U24348 (N_24348,N_24058,N_24022);
nor U24349 (N_24349,N_24108,N_24017);
nor U24350 (N_24350,N_24065,N_24171);
xor U24351 (N_24351,N_24143,N_24081);
and U24352 (N_24352,N_24219,N_24090);
nor U24353 (N_24353,N_24178,N_24048);
xnor U24354 (N_24354,N_24153,N_24185);
xnor U24355 (N_24355,N_24113,N_24050);
nand U24356 (N_24356,N_24055,N_24061);
nand U24357 (N_24357,N_24230,N_24137);
and U24358 (N_24358,N_24084,N_24112);
xnor U24359 (N_24359,N_24180,N_24013);
xor U24360 (N_24360,N_24040,N_24087);
or U24361 (N_24361,N_24046,N_24150);
or U24362 (N_24362,N_24216,N_24167);
nand U24363 (N_24363,N_24246,N_24160);
nor U24364 (N_24364,N_24056,N_24123);
xnor U24365 (N_24365,N_24045,N_24105);
nor U24366 (N_24366,N_24248,N_24024);
nor U24367 (N_24367,N_24161,N_24025);
xnor U24368 (N_24368,N_24191,N_24243);
and U24369 (N_24369,N_24109,N_24005);
nand U24370 (N_24370,N_24163,N_24197);
or U24371 (N_24371,N_24130,N_24089);
nand U24372 (N_24372,N_24104,N_24162);
xor U24373 (N_24373,N_24133,N_24135);
nand U24374 (N_24374,N_24144,N_24201);
nand U24375 (N_24375,N_24240,N_24129);
and U24376 (N_24376,N_24006,N_24220);
nand U24377 (N_24377,N_24198,N_24186);
nand U24378 (N_24378,N_24074,N_24177);
and U24379 (N_24379,N_24030,N_24127);
nand U24380 (N_24380,N_24129,N_24231);
or U24381 (N_24381,N_24162,N_24054);
or U24382 (N_24382,N_24020,N_24093);
nand U24383 (N_24383,N_24202,N_24010);
nand U24384 (N_24384,N_24012,N_24109);
and U24385 (N_24385,N_24194,N_24099);
xnor U24386 (N_24386,N_24162,N_24119);
nor U24387 (N_24387,N_24078,N_24142);
nor U24388 (N_24388,N_24183,N_24198);
nand U24389 (N_24389,N_24009,N_24186);
and U24390 (N_24390,N_24020,N_24043);
nand U24391 (N_24391,N_24049,N_24247);
xor U24392 (N_24392,N_24133,N_24184);
xnor U24393 (N_24393,N_24164,N_24032);
and U24394 (N_24394,N_24239,N_24226);
nor U24395 (N_24395,N_24044,N_24219);
nand U24396 (N_24396,N_24148,N_24165);
nand U24397 (N_24397,N_24208,N_24072);
nand U24398 (N_24398,N_24102,N_24027);
nor U24399 (N_24399,N_24186,N_24221);
xor U24400 (N_24400,N_24155,N_24161);
nand U24401 (N_24401,N_24092,N_24221);
and U24402 (N_24402,N_24007,N_24155);
and U24403 (N_24403,N_24219,N_24236);
nor U24404 (N_24404,N_24000,N_24121);
nor U24405 (N_24405,N_24111,N_24194);
and U24406 (N_24406,N_24131,N_24186);
nor U24407 (N_24407,N_24140,N_24146);
nand U24408 (N_24408,N_24119,N_24226);
nor U24409 (N_24409,N_24178,N_24184);
and U24410 (N_24410,N_24057,N_24109);
nand U24411 (N_24411,N_24093,N_24228);
nor U24412 (N_24412,N_24116,N_24170);
nand U24413 (N_24413,N_24075,N_24243);
and U24414 (N_24414,N_24048,N_24233);
and U24415 (N_24415,N_24192,N_24207);
xor U24416 (N_24416,N_24021,N_24216);
and U24417 (N_24417,N_24076,N_24079);
xnor U24418 (N_24418,N_24119,N_24061);
nor U24419 (N_24419,N_24014,N_24248);
nand U24420 (N_24420,N_24151,N_24105);
and U24421 (N_24421,N_24014,N_24219);
nand U24422 (N_24422,N_24118,N_24100);
xor U24423 (N_24423,N_24109,N_24002);
xnor U24424 (N_24424,N_24153,N_24132);
nor U24425 (N_24425,N_24191,N_24195);
xor U24426 (N_24426,N_24227,N_24010);
nand U24427 (N_24427,N_24160,N_24243);
xnor U24428 (N_24428,N_24235,N_24044);
nor U24429 (N_24429,N_24163,N_24228);
nand U24430 (N_24430,N_24238,N_24192);
xnor U24431 (N_24431,N_24069,N_24241);
nand U24432 (N_24432,N_24019,N_24037);
and U24433 (N_24433,N_24112,N_24039);
xor U24434 (N_24434,N_24018,N_24173);
or U24435 (N_24435,N_24191,N_24228);
nor U24436 (N_24436,N_24072,N_24146);
xor U24437 (N_24437,N_24011,N_24032);
and U24438 (N_24438,N_24208,N_24020);
and U24439 (N_24439,N_24204,N_24180);
nor U24440 (N_24440,N_24016,N_24062);
nand U24441 (N_24441,N_24104,N_24112);
and U24442 (N_24442,N_24138,N_24039);
nor U24443 (N_24443,N_24094,N_24211);
or U24444 (N_24444,N_24003,N_24035);
or U24445 (N_24445,N_24223,N_24240);
nand U24446 (N_24446,N_24230,N_24101);
xor U24447 (N_24447,N_24217,N_24082);
or U24448 (N_24448,N_24161,N_24002);
nand U24449 (N_24449,N_24013,N_24140);
xnor U24450 (N_24450,N_24144,N_24005);
nand U24451 (N_24451,N_24108,N_24073);
and U24452 (N_24452,N_24106,N_24225);
xor U24453 (N_24453,N_24041,N_24217);
nor U24454 (N_24454,N_24086,N_24070);
or U24455 (N_24455,N_24049,N_24246);
nor U24456 (N_24456,N_24094,N_24224);
nor U24457 (N_24457,N_24021,N_24189);
nor U24458 (N_24458,N_24159,N_24095);
or U24459 (N_24459,N_24116,N_24032);
and U24460 (N_24460,N_24198,N_24224);
nor U24461 (N_24461,N_24020,N_24163);
or U24462 (N_24462,N_24169,N_24132);
nand U24463 (N_24463,N_24174,N_24118);
or U24464 (N_24464,N_24061,N_24040);
xor U24465 (N_24465,N_24177,N_24146);
and U24466 (N_24466,N_24034,N_24072);
nand U24467 (N_24467,N_24052,N_24156);
xor U24468 (N_24468,N_24086,N_24202);
nor U24469 (N_24469,N_24106,N_24179);
nor U24470 (N_24470,N_24027,N_24201);
xnor U24471 (N_24471,N_24168,N_24122);
and U24472 (N_24472,N_24086,N_24190);
nor U24473 (N_24473,N_24122,N_24139);
or U24474 (N_24474,N_24020,N_24190);
xor U24475 (N_24475,N_24043,N_24079);
nand U24476 (N_24476,N_24058,N_24166);
xor U24477 (N_24477,N_24082,N_24176);
or U24478 (N_24478,N_24203,N_24169);
xor U24479 (N_24479,N_24159,N_24188);
xor U24480 (N_24480,N_24005,N_24242);
and U24481 (N_24481,N_24180,N_24145);
and U24482 (N_24482,N_24043,N_24219);
nor U24483 (N_24483,N_24048,N_24005);
and U24484 (N_24484,N_24101,N_24084);
and U24485 (N_24485,N_24170,N_24107);
nor U24486 (N_24486,N_24153,N_24117);
or U24487 (N_24487,N_24220,N_24128);
xor U24488 (N_24488,N_24020,N_24229);
or U24489 (N_24489,N_24020,N_24196);
nor U24490 (N_24490,N_24010,N_24059);
xnor U24491 (N_24491,N_24077,N_24024);
nand U24492 (N_24492,N_24109,N_24214);
and U24493 (N_24493,N_24170,N_24152);
and U24494 (N_24494,N_24124,N_24144);
or U24495 (N_24495,N_24027,N_24227);
nor U24496 (N_24496,N_24027,N_24123);
nand U24497 (N_24497,N_24154,N_24065);
nor U24498 (N_24498,N_24017,N_24205);
xor U24499 (N_24499,N_24224,N_24190);
nand U24500 (N_24500,N_24392,N_24262);
nor U24501 (N_24501,N_24450,N_24364);
nor U24502 (N_24502,N_24478,N_24287);
nor U24503 (N_24503,N_24296,N_24292);
xor U24504 (N_24504,N_24488,N_24268);
nand U24505 (N_24505,N_24434,N_24383);
or U24506 (N_24506,N_24410,N_24324);
or U24507 (N_24507,N_24265,N_24336);
and U24508 (N_24508,N_24275,N_24283);
nand U24509 (N_24509,N_24301,N_24323);
or U24510 (N_24510,N_24338,N_24329);
nand U24511 (N_24511,N_24468,N_24489);
xnor U24512 (N_24512,N_24398,N_24496);
and U24513 (N_24513,N_24288,N_24310);
and U24514 (N_24514,N_24472,N_24443);
and U24515 (N_24515,N_24422,N_24269);
or U24516 (N_24516,N_24344,N_24290);
nand U24517 (N_24517,N_24424,N_24384);
nand U24518 (N_24518,N_24377,N_24388);
and U24519 (N_24519,N_24367,N_24448);
nor U24520 (N_24520,N_24390,N_24463);
nand U24521 (N_24521,N_24252,N_24475);
and U24522 (N_24522,N_24473,N_24445);
nand U24523 (N_24523,N_24335,N_24479);
nor U24524 (N_24524,N_24294,N_24406);
nand U24525 (N_24525,N_24404,N_24272);
nand U24526 (N_24526,N_24427,N_24351);
or U24527 (N_24527,N_24251,N_24300);
or U24528 (N_24528,N_24311,N_24391);
or U24529 (N_24529,N_24365,N_24372);
and U24530 (N_24530,N_24442,N_24495);
and U24531 (N_24531,N_24431,N_24277);
or U24532 (N_24532,N_24417,N_24413);
and U24533 (N_24533,N_24433,N_24358);
xnor U24534 (N_24534,N_24374,N_24444);
and U24535 (N_24535,N_24363,N_24407);
nor U24536 (N_24536,N_24451,N_24459);
xor U24537 (N_24537,N_24481,N_24425);
nor U24538 (N_24538,N_24462,N_24399);
nor U24539 (N_24539,N_24334,N_24486);
or U24540 (N_24540,N_24333,N_24313);
nor U24541 (N_24541,N_24352,N_24379);
nor U24542 (N_24542,N_24318,N_24293);
xor U24543 (N_24543,N_24456,N_24341);
or U24544 (N_24544,N_24331,N_24371);
xnor U24545 (N_24545,N_24273,N_24499);
and U24546 (N_24546,N_24426,N_24278);
nand U24547 (N_24547,N_24360,N_24285);
nand U24548 (N_24548,N_24259,N_24393);
or U24549 (N_24549,N_24299,N_24357);
nand U24550 (N_24550,N_24385,N_24423);
xnor U24551 (N_24551,N_24254,N_24416);
nand U24552 (N_24552,N_24271,N_24325);
nor U24553 (N_24553,N_24327,N_24411);
nand U24554 (N_24554,N_24315,N_24326);
xnor U24555 (N_24555,N_24439,N_24470);
or U24556 (N_24556,N_24447,N_24400);
nor U24557 (N_24557,N_24493,N_24304);
xnor U24558 (N_24558,N_24253,N_24342);
nor U24559 (N_24559,N_24343,N_24368);
xor U24560 (N_24560,N_24405,N_24266);
and U24561 (N_24561,N_24322,N_24464);
xnor U24562 (N_24562,N_24366,N_24485);
nor U24563 (N_24563,N_24467,N_24449);
or U24564 (N_24564,N_24440,N_24484);
nand U24565 (N_24565,N_24257,N_24471);
nand U24566 (N_24566,N_24381,N_24250);
and U24567 (N_24567,N_24345,N_24476);
and U24568 (N_24568,N_24282,N_24480);
and U24569 (N_24569,N_24328,N_24307);
nand U24570 (N_24570,N_24261,N_24286);
nor U24571 (N_24571,N_24332,N_24498);
nor U24572 (N_24572,N_24330,N_24319);
xor U24573 (N_24573,N_24289,N_24491);
xnor U24574 (N_24574,N_24403,N_24376);
xnor U24575 (N_24575,N_24477,N_24340);
nor U24576 (N_24576,N_24370,N_24362);
nand U24577 (N_24577,N_24432,N_24380);
xnor U24578 (N_24578,N_24302,N_24437);
and U24579 (N_24579,N_24492,N_24314);
nor U24580 (N_24580,N_24460,N_24429);
and U24581 (N_24581,N_24386,N_24487);
xnor U24582 (N_24582,N_24474,N_24375);
xor U24583 (N_24583,N_24312,N_24441);
nor U24584 (N_24584,N_24316,N_24321);
xor U24585 (N_24585,N_24466,N_24483);
and U24586 (N_24586,N_24276,N_24305);
or U24587 (N_24587,N_24256,N_24308);
and U24588 (N_24588,N_24255,N_24420);
nor U24589 (N_24589,N_24401,N_24309);
nor U24590 (N_24590,N_24455,N_24452);
xor U24591 (N_24591,N_24280,N_24414);
or U24592 (N_24592,N_24497,N_24458);
nor U24593 (N_24593,N_24260,N_24279);
nand U24594 (N_24594,N_24490,N_24430);
or U24595 (N_24595,N_24284,N_24387);
nand U24596 (N_24596,N_24461,N_24438);
nor U24597 (N_24597,N_24446,N_24291);
nand U24598 (N_24598,N_24270,N_24465);
or U24599 (N_24599,N_24274,N_24349);
nand U24600 (N_24600,N_24353,N_24418);
nand U24601 (N_24601,N_24373,N_24482);
nand U24602 (N_24602,N_24454,N_24457);
or U24603 (N_24603,N_24267,N_24298);
or U24604 (N_24604,N_24408,N_24494);
or U24605 (N_24605,N_24435,N_24354);
and U24606 (N_24606,N_24412,N_24264);
or U24607 (N_24607,N_24320,N_24306);
nand U24608 (N_24608,N_24337,N_24263);
nor U24609 (N_24609,N_24428,N_24346);
nor U24610 (N_24610,N_24395,N_24347);
xor U24611 (N_24611,N_24258,N_24297);
xnor U24612 (N_24612,N_24453,N_24382);
nand U24613 (N_24613,N_24369,N_24396);
and U24614 (N_24614,N_24317,N_24350);
xor U24615 (N_24615,N_24359,N_24402);
xor U24616 (N_24616,N_24415,N_24303);
and U24617 (N_24617,N_24421,N_24409);
nor U24618 (N_24618,N_24397,N_24355);
and U24619 (N_24619,N_24295,N_24469);
nor U24620 (N_24620,N_24394,N_24378);
nor U24621 (N_24621,N_24389,N_24348);
or U24622 (N_24622,N_24281,N_24356);
xor U24623 (N_24623,N_24436,N_24361);
and U24624 (N_24624,N_24339,N_24419);
xor U24625 (N_24625,N_24323,N_24417);
nand U24626 (N_24626,N_24276,N_24422);
xor U24627 (N_24627,N_24405,N_24372);
or U24628 (N_24628,N_24401,N_24258);
xnor U24629 (N_24629,N_24342,N_24345);
nor U24630 (N_24630,N_24393,N_24442);
or U24631 (N_24631,N_24318,N_24340);
and U24632 (N_24632,N_24270,N_24321);
and U24633 (N_24633,N_24303,N_24407);
xor U24634 (N_24634,N_24467,N_24394);
nor U24635 (N_24635,N_24395,N_24306);
xnor U24636 (N_24636,N_24285,N_24354);
or U24637 (N_24637,N_24289,N_24315);
nor U24638 (N_24638,N_24463,N_24456);
xnor U24639 (N_24639,N_24488,N_24374);
and U24640 (N_24640,N_24252,N_24344);
nand U24641 (N_24641,N_24328,N_24472);
xnor U24642 (N_24642,N_24350,N_24264);
nor U24643 (N_24643,N_24404,N_24348);
nor U24644 (N_24644,N_24365,N_24467);
and U24645 (N_24645,N_24412,N_24307);
nor U24646 (N_24646,N_24400,N_24449);
and U24647 (N_24647,N_24429,N_24406);
or U24648 (N_24648,N_24390,N_24296);
and U24649 (N_24649,N_24442,N_24386);
xor U24650 (N_24650,N_24254,N_24258);
or U24651 (N_24651,N_24296,N_24490);
nand U24652 (N_24652,N_24387,N_24385);
and U24653 (N_24653,N_24391,N_24272);
and U24654 (N_24654,N_24454,N_24491);
xor U24655 (N_24655,N_24405,N_24434);
and U24656 (N_24656,N_24429,N_24291);
xnor U24657 (N_24657,N_24463,N_24377);
and U24658 (N_24658,N_24486,N_24470);
nand U24659 (N_24659,N_24344,N_24437);
and U24660 (N_24660,N_24424,N_24293);
or U24661 (N_24661,N_24347,N_24343);
xor U24662 (N_24662,N_24368,N_24286);
or U24663 (N_24663,N_24295,N_24410);
xnor U24664 (N_24664,N_24440,N_24266);
xnor U24665 (N_24665,N_24452,N_24331);
or U24666 (N_24666,N_24325,N_24356);
or U24667 (N_24667,N_24253,N_24436);
and U24668 (N_24668,N_24436,N_24283);
and U24669 (N_24669,N_24455,N_24435);
nor U24670 (N_24670,N_24358,N_24351);
xnor U24671 (N_24671,N_24446,N_24250);
or U24672 (N_24672,N_24483,N_24290);
or U24673 (N_24673,N_24296,N_24265);
xnor U24674 (N_24674,N_24471,N_24270);
xor U24675 (N_24675,N_24263,N_24360);
nand U24676 (N_24676,N_24484,N_24448);
xnor U24677 (N_24677,N_24492,N_24354);
nor U24678 (N_24678,N_24499,N_24406);
nor U24679 (N_24679,N_24474,N_24451);
xnor U24680 (N_24680,N_24303,N_24270);
and U24681 (N_24681,N_24361,N_24334);
nor U24682 (N_24682,N_24320,N_24375);
nand U24683 (N_24683,N_24427,N_24366);
xor U24684 (N_24684,N_24380,N_24355);
and U24685 (N_24685,N_24462,N_24431);
xor U24686 (N_24686,N_24358,N_24279);
nor U24687 (N_24687,N_24405,N_24365);
nor U24688 (N_24688,N_24338,N_24461);
nand U24689 (N_24689,N_24314,N_24370);
xor U24690 (N_24690,N_24358,N_24459);
and U24691 (N_24691,N_24393,N_24441);
nor U24692 (N_24692,N_24345,N_24312);
xor U24693 (N_24693,N_24412,N_24493);
and U24694 (N_24694,N_24301,N_24333);
and U24695 (N_24695,N_24392,N_24450);
or U24696 (N_24696,N_24488,N_24257);
and U24697 (N_24697,N_24299,N_24399);
and U24698 (N_24698,N_24422,N_24351);
or U24699 (N_24699,N_24422,N_24279);
xnor U24700 (N_24700,N_24439,N_24438);
nor U24701 (N_24701,N_24296,N_24403);
nand U24702 (N_24702,N_24315,N_24312);
nor U24703 (N_24703,N_24463,N_24484);
or U24704 (N_24704,N_24320,N_24398);
and U24705 (N_24705,N_24322,N_24467);
nand U24706 (N_24706,N_24410,N_24312);
nand U24707 (N_24707,N_24305,N_24327);
and U24708 (N_24708,N_24366,N_24362);
nand U24709 (N_24709,N_24332,N_24408);
nor U24710 (N_24710,N_24278,N_24410);
and U24711 (N_24711,N_24399,N_24341);
xnor U24712 (N_24712,N_24466,N_24363);
nand U24713 (N_24713,N_24485,N_24438);
or U24714 (N_24714,N_24256,N_24494);
xnor U24715 (N_24715,N_24453,N_24358);
and U24716 (N_24716,N_24277,N_24327);
or U24717 (N_24717,N_24399,N_24270);
xnor U24718 (N_24718,N_24316,N_24282);
and U24719 (N_24719,N_24443,N_24323);
or U24720 (N_24720,N_24347,N_24375);
nor U24721 (N_24721,N_24413,N_24380);
nor U24722 (N_24722,N_24336,N_24451);
xnor U24723 (N_24723,N_24263,N_24331);
nand U24724 (N_24724,N_24289,N_24278);
nand U24725 (N_24725,N_24253,N_24275);
nor U24726 (N_24726,N_24406,N_24400);
nor U24727 (N_24727,N_24386,N_24355);
and U24728 (N_24728,N_24355,N_24302);
nor U24729 (N_24729,N_24308,N_24331);
and U24730 (N_24730,N_24330,N_24257);
nor U24731 (N_24731,N_24424,N_24446);
and U24732 (N_24732,N_24330,N_24464);
or U24733 (N_24733,N_24384,N_24391);
and U24734 (N_24734,N_24277,N_24361);
xnor U24735 (N_24735,N_24315,N_24467);
xor U24736 (N_24736,N_24462,N_24319);
or U24737 (N_24737,N_24297,N_24278);
and U24738 (N_24738,N_24469,N_24334);
and U24739 (N_24739,N_24341,N_24400);
xor U24740 (N_24740,N_24266,N_24275);
and U24741 (N_24741,N_24293,N_24259);
nand U24742 (N_24742,N_24378,N_24389);
or U24743 (N_24743,N_24465,N_24266);
nand U24744 (N_24744,N_24466,N_24498);
and U24745 (N_24745,N_24499,N_24419);
nor U24746 (N_24746,N_24439,N_24314);
and U24747 (N_24747,N_24493,N_24386);
or U24748 (N_24748,N_24359,N_24426);
or U24749 (N_24749,N_24338,N_24428);
nor U24750 (N_24750,N_24627,N_24571);
or U24751 (N_24751,N_24698,N_24618);
or U24752 (N_24752,N_24561,N_24688);
nand U24753 (N_24753,N_24702,N_24685);
nor U24754 (N_24754,N_24638,N_24542);
nand U24755 (N_24755,N_24531,N_24600);
nand U24756 (N_24756,N_24739,N_24729);
and U24757 (N_24757,N_24512,N_24631);
xor U24758 (N_24758,N_24540,N_24690);
nand U24759 (N_24759,N_24615,N_24641);
nor U24760 (N_24760,N_24606,N_24720);
or U24761 (N_24761,N_24582,N_24695);
xor U24762 (N_24762,N_24522,N_24673);
or U24763 (N_24763,N_24676,N_24506);
or U24764 (N_24764,N_24643,N_24577);
nor U24765 (N_24765,N_24722,N_24664);
nand U24766 (N_24766,N_24629,N_24634);
or U24767 (N_24767,N_24710,N_24593);
xor U24768 (N_24768,N_24516,N_24687);
nor U24769 (N_24769,N_24658,N_24548);
and U24770 (N_24770,N_24713,N_24611);
nor U24771 (N_24771,N_24630,N_24741);
or U24772 (N_24772,N_24632,N_24511);
or U24773 (N_24773,N_24502,N_24507);
nand U24774 (N_24774,N_24671,N_24662);
xor U24775 (N_24775,N_24591,N_24552);
nand U24776 (N_24776,N_24694,N_24547);
and U24777 (N_24777,N_24564,N_24563);
xnor U24778 (N_24778,N_24579,N_24723);
xnor U24779 (N_24779,N_24665,N_24738);
nand U24780 (N_24780,N_24706,N_24523);
nand U24781 (N_24781,N_24545,N_24728);
and U24782 (N_24782,N_24566,N_24602);
nor U24783 (N_24783,N_24649,N_24529);
xor U24784 (N_24784,N_24733,N_24576);
xor U24785 (N_24785,N_24518,N_24709);
xnor U24786 (N_24786,N_24644,N_24521);
nand U24787 (N_24787,N_24537,N_24660);
xor U24788 (N_24788,N_24684,N_24520);
xnor U24789 (N_24789,N_24726,N_24554);
or U24790 (N_24790,N_24693,N_24652);
xnor U24791 (N_24791,N_24683,N_24674);
nor U24792 (N_24792,N_24725,N_24501);
nor U24793 (N_24793,N_24642,N_24678);
nor U24794 (N_24794,N_24508,N_24704);
and U24795 (N_24795,N_24635,N_24603);
xnor U24796 (N_24796,N_24715,N_24543);
and U24797 (N_24797,N_24569,N_24595);
nor U24798 (N_24798,N_24609,N_24539);
or U24799 (N_24799,N_24639,N_24736);
or U24800 (N_24800,N_24650,N_24553);
nor U24801 (N_24801,N_24747,N_24617);
xnor U24802 (N_24802,N_24742,N_24515);
nand U24803 (N_24803,N_24653,N_24610);
or U24804 (N_24804,N_24580,N_24573);
or U24805 (N_24805,N_24605,N_24705);
nand U24806 (N_24806,N_24680,N_24614);
xnor U24807 (N_24807,N_24568,N_24712);
xor U24808 (N_24808,N_24556,N_24669);
nand U24809 (N_24809,N_24621,N_24596);
and U24810 (N_24810,N_24581,N_24717);
and U24811 (N_24811,N_24743,N_24656);
nor U24812 (N_24812,N_24585,N_24624);
nor U24813 (N_24813,N_24551,N_24558);
and U24814 (N_24814,N_24746,N_24696);
or U24815 (N_24815,N_24503,N_24536);
xnor U24816 (N_24816,N_24730,N_24748);
or U24817 (N_24817,N_24578,N_24549);
nand U24818 (N_24818,N_24519,N_24724);
xnor U24819 (N_24819,N_24535,N_24677);
nor U24820 (N_24820,N_24588,N_24657);
and U24821 (N_24821,N_24744,N_24703);
nand U24822 (N_24822,N_24533,N_24594);
and U24823 (N_24823,N_24625,N_24623);
nand U24824 (N_24824,N_24574,N_24646);
nand U24825 (N_24825,N_24682,N_24740);
nand U24826 (N_24826,N_24557,N_24708);
or U24827 (N_24827,N_24721,N_24679);
or U24828 (N_24828,N_24672,N_24616);
xor U24829 (N_24829,N_24716,N_24514);
xnor U24830 (N_24830,N_24636,N_24647);
or U24831 (N_24831,N_24598,N_24661);
nor U24832 (N_24832,N_24697,N_24538);
nor U24833 (N_24833,N_24604,N_24622);
nor U24834 (N_24834,N_24675,N_24544);
nor U24835 (N_24835,N_24525,N_24524);
and U24836 (N_24836,N_24648,N_24637);
nand U24837 (N_24837,N_24667,N_24587);
and U24838 (N_24838,N_24526,N_24668);
and U24839 (N_24839,N_24601,N_24654);
and U24840 (N_24840,N_24714,N_24541);
or U24841 (N_24841,N_24560,N_24612);
xnor U24842 (N_24842,N_24559,N_24719);
xnor U24843 (N_24843,N_24607,N_24555);
xor U24844 (N_24844,N_24626,N_24613);
nor U24845 (N_24845,N_24735,N_24711);
nand U24846 (N_24846,N_24586,N_24510);
nand U24847 (N_24847,N_24500,N_24590);
and U24848 (N_24848,N_24528,N_24749);
nor U24849 (N_24849,N_24663,N_24718);
nor U24850 (N_24850,N_24651,N_24567);
nor U24851 (N_24851,N_24686,N_24589);
and U24852 (N_24852,N_24659,N_24691);
or U24853 (N_24853,N_24534,N_24745);
or U24854 (N_24854,N_24546,N_24592);
nor U24855 (N_24855,N_24597,N_24628);
nand U24856 (N_24856,N_24737,N_24701);
or U24857 (N_24857,N_24599,N_24527);
or U24858 (N_24858,N_24530,N_24562);
and U24859 (N_24859,N_24509,N_24505);
xnor U24860 (N_24860,N_24700,N_24655);
nand U24861 (N_24861,N_24692,N_24565);
or U24862 (N_24862,N_24619,N_24645);
xnor U24863 (N_24863,N_24727,N_24734);
nor U24864 (N_24864,N_24513,N_24699);
xnor U24865 (N_24865,N_24608,N_24670);
xor U24866 (N_24866,N_24517,N_24504);
xor U24867 (N_24867,N_24532,N_24583);
nand U24868 (N_24868,N_24640,N_24620);
nor U24869 (N_24869,N_24689,N_24575);
nand U24870 (N_24870,N_24732,N_24633);
xor U24871 (N_24871,N_24681,N_24584);
nor U24872 (N_24872,N_24666,N_24550);
xor U24873 (N_24873,N_24707,N_24570);
nand U24874 (N_24874,N_24731,N_24572);
and U24875 (N_24875,N_24551,N_24506);
or U24876 (N_24876,N_24668,N_24587);
nand U24877 (N_24877,N_24542,N_24624);
nand U24878 (N_24878,N_24549,N_24687);
nor U24879 (N_24879,N_24644,N_24509);
or U24880 (N_24880,N_24719,N_24621);
or U24881 (N_24881,N_24681,N_24696);
nor U24882 (N_24882,N_24613,N_24734);
nand U24883 (N_24883,N_24601,N_24535);
xor U24884 (N_24884,N_24660,N_24652);
nand U24885 (N_24885,N_24592,N_24585);
or U24886 (N_24886,N_24510,N_24749);
xnor U24887 (N_24887,N_24597,N_24664);
nor U24888 (N_24888,N_24502,N_24682);
xor U24889 (N_24889,N_24533,N_24701);
xor U24890 (N_24890,N_24579,N_24655);
nor U24891 (N_24891,N_24660,N_24523);
and U24892 (N_24892,N_24677,N_24665);
and U24893 (N_24893,N_24709,N_24633);
xor U24894 (N_24894,N_24728,N_24596);
or U24895 (N_24895,N_24662,N_24519);
nor U24896 (N_24896,N_24661,N_24664);
nand U24897 (N_24897,N_24518,N_24748);
xnor U24898 (N_24898,N_24727,N_24645);
nor U24899 (N_24899,N_24737,N_24710);
and U24900 (N_24900,N_24725,N_24642);
nor U24901 (N_24901,N_24703,N_24585);
nor U24902 (N_24902,N_24686,N_24588);
and U24903 (N_24903,N_24543,N_24654);
nor U24904 (N_24904,N_24696,N_24665);
nand U24905 (N_24905,N_24589,N_24684);
xor U24906 (N_24906,N_24567,N_24617);
or U24907 (N_24907,N_24606,N_24504);
and U24908 (N_24908,N_24543,N_24501);
nand U24909 (N_24909,N_24632,N_24633);
and U24910 (N_24910,N_24649,N_24584);
nor U24911 (N_24911,N_24661,N_24654);
or U24912 (N_24912,N_24680,N_24523);
or U24913 (N_24913,N_24632,N_24515);
xor U24914 (N_24914,N_24622,N_24609);
and U24915 (N_24915,N_24519,N_24727);
or U24916 (N_24916,N_24642,N_24720);
xnor U24917 (N_24917,N_24520,N_24523);
xnor U24918 (N_24918,N_24588,N_24722);
and U24919 (N_24919,N_24580,N_24680);
nand U24920 (N_24920,N_24733,N_24558);
nand U24921 (N_24921,N_24612,N_24552);
and U24922 (N_24922,N_24660,N_24530);
nor U24923 (N_24923,N_24606,N_24659);
xor U24924 (N_24924,N_24599,N_24621);
nor U24925 (N_24925,N_24620,N_24578);
nor U24926 (N_24926,N_24733,N_24723);
xor U24927 (N_24927,N_24653,N_24618);
and U24928 (N_24928,N_24714,N_24628);
and U24929 (N_24929,N_24650,N_24511);
nand U24930 (N_24930,N_24644,N_24537);
nand U24931 (N_24931,N_24587,N_24674);
nor U24932 (N_24932,N_24706,N_24628);
nand U24933 (N_24933,N_24597,N_24739);
and U24934 (N_24934,N_24611,N_24527);
nor U24935 (N_24935,N_24600,N_24545);
nor U24936 (N_24936,N_24744,N_24557);
nor U24937 (N_24937,N_24671,N_24645);
and U24938 (N_24938,N_24662,N_24713);
xor U24939 (N_24939,N_24592,N_24596);
xor U24940 (N_24940,N_24581,N_24503);
or U24941 (N_24941,N_24740,N_24615);
or U24942 (N_24942,N_24599,N_24533);
or U24943 (N_24943,N_24543,N_24620);
and U24944 (N_24944,N_24647,N_24590);
xnor U24945 (N_24945,N_24701,N_24580);
or U24946 (N_24946,N_24630,N_24502);
nor U24947 (N_24947,N_24599,N_24689);
or U24948 (N_24948,N_24502,N_24555);
or U24949 (N_24949,N_24569,N_24744);
xor U24950 (N_24950,N_24743,N_24609);
and U24951 (N_24951,N_24665,N_24614);
and U24952 (N_24952,N_24688,N_24669);
nand U24953 (N_24953,N_24724,N_24563);
xor U24954 (N_24954,N_24617,N_24685);
and U24955 (N_24955,N_24618,N_24596);
or U24956 (N_24956,N_24611,N_24506);
xor U24957 (N_24957,N_24714,N_24614);
nand U24958 (N_24958,N_24577,N_24524);
and U24959 (N_24959,N_24629,N_24605);
nor U24960 (N_24960,N_24610,N_24726);
nand U24961 (N_24961,N_24692,N_24631);
xnor U24962 (N_24962,N_24562,N_24528);
xnor U24963 (N_24963,N_24727,N_24594);
or U24964 (N_24964,N_24599,N_24706);
or U24965 (N_24965,N_24526,N_24570);
or U24966 (N_24966,N_24506,N_24655);
or U24967 (N_24967,N_24592,N_24552);
xnor U24968 (N_24968,N_24699,N_24612);
or U24969 (N_24969,N_24564,N_24514);
or U24970 (N_24970,N_24679,N_24667);
nor U24971 (N_24971,N_24530,N_24563);
and U24972 (N_24972,N_24599,N_24691);
nand U24973 (N_24973,N_24697,N_24506);
nor U24974 (N_24974,N_24740,N_24656);
and U24975 (N_24975,N_24703,N_24627);
or U24976 (N_24976,N_24682,N_24621);
and U24977 (N_24977,N_24667,N_24663);
nor U24978 (N_24978,N_24720,N_24651);
xnor U24979 (N_24979,N_24657,N_24683);
and U24980 (N_24980,N_24669,N_24514);
and U24981 (N_24981,N_24672,N_24532);
and U24982 (N_24982,N_24703,N_24531);
nand U24983 (N_24983,N_24736,N_24747);
xnor U24984 (N_24984,N_24660,N_24712);
xnor U24985 (N_24985,N_24578,N_24611);
nor U24986 (N_24986,N_24512,N_24563);
or U24987 (N_24987,N_24524,N_24713);
nand U24988 (N_24988,N_24512,N_24721);
or U24989 (N_24989,N_24682,N_24681);
nand U24990 (N_24990,N_24658,N_24726);
and U24991 (N_24991,N_24748,N_24695);
or U24992 (N_24992,N_24515,N_24731);
nand U24993 (N_24993,N_24593,N_24584);
or U24994 (N_24994,N_24586,N_24610);
xor U24995 (N_24995,N_24550,N_24614);
nand U24996 (N_24996,N_24717,N_24720);
xor U24997 (N_24997,N_24679,N_24500);
and U24998 (N_24998,N_24720,N_24673);
xnor U24999 (N_24999,N_24727,N_24684);
nand U25000 (N_25000,N_24819,N_24908);
nand U25001 (N_25001,N_24821,N_24828);
or U25002 (N_25002,N_24831,N_24861);
xor U25003 (N_25003,N_24995,N_24941);
or U25004 (N_25004,N_24980,N_24790);
nor U25005 (N_25005,N_24862,N_24864);
or U25006 (N_25006,N_24834,N_24939);
nor U25007 (N_25007,N_24800,N_24762);
and U25008 (N_25008,N_24925,N_24898);
or U25009 (N_25009,N_24945,N_24927);
or U25010 (N_25010,N_24998,N_24962);
and U25011 (N_25011,N_24884,N_24996);
xor U25012 (N_25012,N_24863,N_24934);
nor U25013 (N_25013,N_24817,N_24794);
nor U25014 (N_25014,N_24988,N_24993);
nand U25015 (N_25015,N_24948,N_24901);
xor U25016 (N_25016,N_24932,N_24920);
nor U25017 (N_25017,N_24857,N_24913);
nor U25018 (N_25018,N_24965,N_24893);
xor U25019 (N_25019,N_24890,N_24809);
nand U25020 (N_25020,N_24795,N_24771);
xnor U25021 (N_25021,N_24798,N_24785);
and U25022 (N_25022,N_24974,N_24887);
nand U25023 (N_25023,N_24899,N_24838);
nor U25024 (N_25024,N_24982,N_24793);
nor U25025 (N_25025,N_24791,N_24815);
or U25026 (N_25026,N_24879,N_24903);
or U25027 (N_25027,N_24847,N_24865);
xnor U25028 (N_25028,N_24975,N_24813);
nand U25029 (N_25029,N_24990,N_24849);
nor U25030 (N_25030,N_24937,N_24875);
nand U25031 (N_25031,N_24753,N_24846);
xor U25032 (N_25032,N_24891,N_24818);
nand U25033 (N_25033,N_24970,N_24827);
nor U25034 (N_25034,N_24867,N_24919);
nand U25035 (N_25035,N_24967,N_24900);
nor U25036 (N_25036,N_24829,N_24772);
or U25037 (N_25037,N_24757,N_24873);
and U25038 (N_25038,N_24897,N_24957);
nor U25039 (N_25039,N_24839,N_24769);
nor U25040 (N_25040,N_24788,N_24853);
nand U25041 (N_25041,N_24959,N_24935);
and U25042 (N_25042,N_24947,N_24924);
nor U25043 (N_25043,N_24981,N_24997);
nor U25044 (N_25044,N_24953,N_24782);
or U25045 (N_25045,N_24816,N_24783);
xnor U25046 (N_25046,N_24910,N_24999);
xor U25047 (N_25047,N_24835,N_24911);
or U25048 (N_25048,N_24840,N_24807);
nand U25049 (N_25049,N_24752,N_24960);
xor U25050 (N_25050,N_24781,N_24869);
and U25051 (N_25051,N_24928,N_24804);
nor U25052 (N_25052,N_24767,N_24918);
or U25053 (N_25053,N_24758,N_24973);
nand U25054 (N_25054,N_24797,N_24796);
nand U25055 (N_25055,N_24933,N_24989);
or U25056 (N_25056,N_24986,N_24904);
and U25057 (N_25057,N_24824,N_24880);
xnor U25058 (N_25058,N_24885,N_24836);
or U25059 (N_25059,N_24860,N_24765);
and U25060 (N_25060,N_24801,N_24950);
or U25061 (N_25061,N_24978,N_24940);
nand U25062 (N_25062,N_24979,N_24876);
xnor U25063 (N_25063,N_24754,N_24912);
nor U25064 (N_25064,N_24915,N_24949);
nor U25065 (N_25065,N_24905,N_24942);
or U25066 (N_25066,N_24868,N_24907);
xnor U25067 (N_25067,N_24803,N_24766);
xnor U25068 (N_25068,N_24844,N_24751);
and U25069 (N_25069,N_24780,N_24787);
nand U25070 (N_25070,N_24922,N_24814);
xnor U25071 (N_25071,N_24851,N_24823);
nand U25072 (N_25072,N_24972,N_24943);
xor U25073 (N_25073,N_24810,N_24811);
and U25074 (N_25074,N_24837,N_24969);
xor U25075 (N_25075,N_24768,N_24878);
and U25076 (N_25076,N_24888,N_24841);
nand U25077 (N_25077,N_24854,N_24799);
xnor U25078 (N_25078,N_24786,N_24968);
nand U25079 (N_25079,N_24802,N_24761);
and U25080 (N_25080,N_24806,N_24850);
or U25081 (N_25081,N_24994,N_24833);
and U25082 (N_25082,N_24773,N_24936);
nor U25083 (N_25083,N_24984,N_24845);
xnor U25084 (N_25084,N_24874,N_24755);
nand U25085 (N_25085,N_24777,N_24848);
or U25086 (N_25086,N_24938,N_24930);
or U25087 (N_25087,N_24871,N_24764);
nand U25088 (N_25088,N_24923,N_24832);
nand U25089 (N_25089,N_24921,N_24991);
nand U25090 (N_25090,N_24842,N_24983);
nor U25091 (N_25091,N_24902,N_24843);
and U25092 (N_25092,N_24951,N_24866);
or U25093 (N_25093,N_24808,N_24852);
and U25094 (N_25094,N_24870,N_24770);
nor U25095 (N_25095,N_24856,N_24830);
nor U25096 (N_25096,N_24775,N_24763);
xor U25097 (N_25097,N_24859,N_24909);
or U25098 (N_25098,N_24776,N_24971);
nor U25099 (N_25099,N_24882,N_24877);
or U25100 (N_25100,N_24822,N_24976);
or U25101 (N_25101,N_24812,N_24826);
nor U25102 (N_25102,N_24805,N_24855);
or U25103 (N_25103,N_24759,N_24774);
or U25104 (N_25104,N_24987,N_24883);
nor U25105 (N_25105,N_24958,N_24944);
nand U25106 (N_25106,N_24964,N_24985);
nand U25107 (N_25107,N_24858,N_24926);
xor U25108 (N_25108,N_24886,N_24881);
nor U25109 (N_25109,N_24916,N_24929);
xor U25110 (N_25110,N_24914,N_24917);
nand U25111 (N_25111,N_24820,N_24954);
xor U25112 (N_25112,N_24756,N_24778);
nor U25113 (N_25113,N_24963,N_24895);
nand U25114 (N_25114,N_24789,N_24889);
and U25115 (N_25115,N_24779,N_24896);
nor U25116 (N_25116,N_24952,N_24992);
nor U25117 (N_25117,N_24750,N_24961);
xor U25118 (N_25118,N_24966,N_24784);
xnor U25119 (N_25119,N_24872,N_24906);
or U25120 (N_25120,N_24956,N_24825);
nor U25121 (N_25121,N_24792,N_24892);
nand U25122 (N_25122,N_24931,N_24894);
or U25123 (N_25123,N_24946,N_24955);
xor U25124 (N_25124,N_24760,N_24977);
and U25125 (N_25125,N_24819,N_24766);
nor U25126 (N_25126,N_24752,N_24892);
nor U25127 (N_25127,N_24774,N_24901);
nand U25128 (N_25128,N_24821,N_24910);
nor U25129 (N_25129,N_24852,N_24911);
xor U25130 (N_25130,N_24992,N_24862);
nor U25131 (N_25131,N_24797,N_24979);
or U25132 (N_25132,N_24770,N_24913);
and U25133 (N_25133,N_24868,N_24882);
and U25134 (N_25134,N_24920,N_24916);
or U25135 (N_25135,N_24980,N_24903);
or U25136 (N_25136,N_24912,N_24750);
nor U25137 (N_25137,N_24929,N_24990);
xnor U25138 (N_25138,N_24822,N_24997);
and U25139 (N_25139,N_24821,N_24806);
or U25140 (N_25140,N_24786,N_24902);
nor U25141 (N_25141,N_24760,N_24781);
xor U25142 (N_25142,N_24925,N_24754);
xnor U25143 (N_25143,N_24883,N_24775);
and U25144 (N_25144,N_24855,N_24942);
xor U25145 (N_25145,N_24782,N_24871);
xnor U25146 (N_25146,N_24850,N_24819);
nand U25147 (N_25147,N_24810,N_24759);
nand U25148 (N_25148,N_24775,N_24859);
xor U25149 (N_25149,N_24984,N_24953);
xnor U25150 (N_25150,N_24906,N_24999);
and U25151 (N_25151,N_24833,N_24998);
or U25152 (N_25152,N_24941,N_24866);
xor U25153 (N_25153,N_24778,N_24874);
or U25154 (N_25154,N_24845,N_24965);
nand U25155 (N_25155,N_24977,N_24922);
nand U25156 (N_25156,N_24951,N_24948);
or U25157 (N_25157,N_24848,N_24990);
or U25158 (N_25158,N_24841,N_24855);
xor U25159 (N_25159,N_24759,N_24932);
and U25160 (N_25160,N_24940,N_24873);
or U25161 (N_25161,N_24858,N_24997);
nand U25162 (N_25162,N_24815,N_24942);
nand U25163 (N_25163,N_24876,N_24892);
and U25164 (N_25164,N_24813,N_24873);
xnor U25165 (N_25165,N_24993,N_24839);
nand U25166 (N_25166,N_24915,N_24919);
and U25167 (N_25167,N_24753,N_24983);
or U25168 (N_25168,N_24866,N_24795);
nor U25169 (N_25169,N_24835,N_24891);
nand U25170 (N_25170,N_24826,N_24787);
xnor U25171 (N_25171,N_24772,N_24864);
or U25172 (N_25172,N_24865,N_24755);
nand U25173 (N_25173,N_24942,N_24793);
xor U25174 (N_25174,N_24888,N_24786);
nand U25175 (N_25175,N_24909,N_24755);
xnor U25176 (N_25176,N_24824,N_24935);
nand U25177 (N_25177,N_24804,N_24977);
or U25178 (N_25178,N_24853,N_24852);
xor U25179 (N_25179,N_24976,N_24982);
and U25180 (N_25180,N_24996,N_24757);
xor U25181 (N_25181,N_24753,N_24937);
xor U25182 (N_25182,N_24936,N_24844);
or U25183 (N_25183,N_24885,N_24853);
nand U25184 (N_25184,N_24927,N_24942);
nand U25185 (N_25185,N_24777,N_24942);
nand U25186 (N_25186,N_24754,N_24870);
nor U25187 (N_25187,N_24998,N_24906);
or U25188 (N_25188,N_24804,N_24948);
and U25189 (N_25189,N_24919,N_24950);
nor U25190 (N_25190,N_24839,N_24802);
nand U25191 (N_25191,N_24902,N_24911);
nor U25192 (N_25192,N_24755,N_24889);
nand U25193 (N_25193,N_24759,N_24829);
nand U25194 (N_25194,N_24894,N_24928);
or U25195 (N_25195,N_24932,N_24792);
and U25196 (N_25196,N_24778,N_24945);
and U25197 (N_25197,N_24952,N_24796);
nand U25198 (N_25198,N_24932,N_24853);
and U25199 (N_25199,N_24873,N_24797);
xnor U25200 (N_25200,N_24956,N_24921);
nand U25201 (N_25201,N_24850,N_24866);
nor U25202 (N_25202,N_24901,N_24899);
or U25203 (N_25203,N_24978,N_24889);
nor U25204 (N_25204,N_24974,N_24907);
nor U25205 (N_25205,N_24792,N_24767);
or U25206 (N_25206,N_24783,N_24874);
and U25207 (N_25207,N_24904,N_24878);
nor U25208 (N_25208,N_24774,N_24904);
nor U25209 (N_25209,N_24835,N_24958);
nor U25210 (N_25210,N_24829,N_24998);
xnor U25211 (N_25211,N_24870,N_24789);
nor U25212 (N_25212,N_24919,N_24990);
or U25213 (N_25213,N_24923,N_24887);
xor U25214 (N_25214,N_24967,N_24856);
and U25215 (N_25215,N_24816,N_24869);
nor U25216 (N_25216,N_24955,N_24876);
and U25217 (N_25217,N_24882,N_24874);
or U25218 (N_25218,N_24971,N_24952);
nor U25219 (N_25219,N_24798,N_24953);
xnor U25220 (N_25220,N_24840,N_24891);
xor U25221 (N_25221,N_24869,N_24755);
and U25222 (N_25222,N_24829,N_24880);
nand U25223 (N_25223,N_24947,N_24842);
xnor U25224 (N_25224,N_24942,N_24985);
nand U25225 (N_25225,N_24934,N_24948);
xor U25226 (N_25226,N_24809,N_24781);
nand U25227 (N_25227,N_24985,N_24773);
xor U25228 (N_25228,N_24793,N_24753);
nor U25229 (N_25229,N_24758,N_24895);
and U25230 (N_25230,N_24930,N_24959);
nand U25231 (N_25231,N_24888,N_24853);
or U25232 (N_25232,N_24800,N_24869);
nor U25233 (N_25233,N_24908,N_24792);
nand U25234 (N_25234,N_24894,N_24797);
and U25235 (N_25235,N_24881,N_24992);
nor U25236 (N_25236,N_24950,N_24880);
and U25237 (N_25237,N_24760,N_24946);
nor U25238 (N_25238,N_24796,N_24763);
nand U25239 (N_25239,N_24962,N_24995);
or U25240 (N_25240,N_24862,N_24801);
nand U25241 (N_25241,N_24923,N_24830);
nand U25242 (N_25242,N_24845,N_24776);
or U25243 (N_25243,N_24872,N_24893);
nand U25244 (N_25244,N_24954,N_24957);
xor U25245 (N_25245,N_24886,N_24772);
xnor U25246 (N_25246,N_24911,N_24901);
or U25247 (N_25247,N_24950,N_24861);
or U25248 (N_25248,N_24869,N_24853);
or U25249 (N_25249,N_24882,N_24841);
nor U25250 (N_25250,N_25066,N_25170);
xor U25251 (N_25251,N_25033,N_25050);
xor U25252 (N_25252,N_25076,N_25063);
or U25253 (N_25253,N_25117,N_25139);
or U25254 (N_25254,N_25042,N_25086);
and U25255 (N_25255,N_25005,N_25093);
and U25256 (N_25256,N_25031,N_25201);
nand U25257 (N_25257,N_25237,N_25132);
xnor U25258 (N_25258,N_25202,N_25136);
and U25259 (N_25259,N_25186,N_25133);
and U25260 (N_25260,N_25032,N_25011);
and U25261 (N_25261,N_25159,N_25147);
and U25262 (N_25262,N_25046,N_25069);
and U25263 (N_25263,N_25240,N_25087);
and U25264 (N_25264,N_25001,N_25099);
nor U25265 (N_25265,N_25016,N_25096);
or U25266 (N_25266,N_25241,N_25056);
nand U25267 (N_25267,N_25009,N_25165);
nor U25268 (N_25268,N_25143,N_25034);
and U25269 (N_25269,N_25052,N_25198);
or U25270 (N_25270,N_25141,N_25120);
xnor U25271 (N_25271,N_25224,N_25024);
xor U25272 (N_25272,N_25043,N_25223);
and U25273 (N_25273,N_25209,N_25000);
and U25274 (N_25274,N_25212,N_25184);
nand U25275 (N_25275,N_25064,N_25220);
nand U25276 (N_25276,N_25178,N_25015);
nor U25277 (N_25277,N_25007,N_25194);
and U25278 (N_25278,N_25127,N_25107);
and U25279 (N_25279,N_25183,N_25062);
xor U25280 (N_25280,N_25053,N_25082);
and U25281 (N_25281,N_25190,N_25094);
and U25282 (N_25282,N_25074,N_25123);
nor U25283 (N_25283,N_25036,N_25145);
nor U25284 (N_25284,N_25073,N_25051);
and U25285 (N_25285,N_25238,N_25142);
xnor U25286 (N_25286,N_25232,N_25246);
xor U25287 (N_25287,N_25089,N_25155);
and U25288 (N_25288,N_25029,N_25134);
nand U25289 (N_25289,N_25030,N_25037);
xnor U25290 (N_25290,N_25163,N_25226);
and U25291 (N_25291,N_25188,N_25185);
or U25292 (N_25292,N_25217,N_25167);
and U25293 (N_25293,N_25208,N_25017);
nor U25294 (N_25294,N_25152,N_25078);
nand U25295 (N_25295,N_25138,N_25164);
or U25296 (N_25296,N_25041,N_25021);
and U25297 (N_25297,N_25070,N_25199);
nand U25298 (N_25298,N_25072,N_25195);
or U25299 (N_25299,N_25023,N_25144);
nand U25300 (N_25300,N_25045,N_25088);
and U25301 (N_25301,N_25181,N_25026);
nor U25302 (N_25302,N_25112,N_25192);
xor U25303 (N_25303,N_25210,N_25101);
nor U25304 (N_25304,N_25214,N_25048);
and U25305 (N_25305,N_25137,N_25233);
or U25306 (N_25306,N_25110,N_25028);
xnor U25307 (N_25307,N_25105,N_25013);
or U25308 (N_25308,N_25124,N_25244);
nand U25309 (N_25309,N_25189,N_25049);
or U25310 (N_25310,N_25219,N_25229);
nor U25311 (N_25311,N_25039,N_25111);
nand U25312 (N_25312,N_25221,N_25079);
nand U25313 (N_25313,N_25077,N_25010);
or U25314 (N_25314,N_25040,N_25191);
or U25315 (N_25315,N_25003,N_25216);
xor U25316 (N_25316,N_25239,N_25154);
and U25317 (N_25317,N_25098,N_25203);
and U25318 (N_25318,N_25228,N_25100);
nor U25319 (N_25319,N_25204,N_25193);
and U25320 (N_25320,N_25174,N_25162);
nor U25321 (N_25321,N_25166,N_25230);
or U25322 (N_25322,N_25047,N_25084);
xnor U25323 (N_25323,N_25108,N_25083);
nand U25324 (N_25324,N_25057,N_25218);
nor U25325 (N_25325,N_25243,N_25182);
nor U25326 (N_25326,N_25151,N_25231);
nor U25327 (N_25327,N_25106,N_25177);
and U25328 (N_25328,N_25156,N_25027);
xnor U25329 (N_25329,N_25125,N_25002);
or U25330 (N_25330,N_25104,N_25058);
xnor U25331 (N_25331,N_25242,N_25012);
and U25332 (N_25332,N_25222,N_25158);
nor U25333 (N_25333,N_25160,N_25175);
and U25334 (N_25334,N_25196,N_25197);
xnor U25335 (N_25335,N_25187,N_25095);
and U25336 (N_25336,N_25071,N_25067);
nand U25337 (N_25337,N_25019,N_25014);
nand U25338 (N_25338,N_25103,N_25249);
nor U25339 (N_25339,N_25092,N_25206);
or U25340 (N_25340,N_25006,N_25004);
nor U25341 (N_25341,N_25200,N_25245);
nor U25342 (N_25342,N_25115,N_25128);
or U25343 (N_25343,N_25227,N_25131);
nor U25344 (N_25344,N_25234,N_25135);
nand U25345 (N_25345,N_25247,N_25207);
or U25346 (N_25346,N_25236,N_25179);
nor U25347 (N_25347,N_25122,N_25114);
and U25348 (N_25348,N_25161,N_25215);
nor U25349 (N_25349,N_25061,N_25038);
nand U25350 (N_25350,N_25109,N_25059);
nor U25351 (N_25351,N_25149,N_25169);
xnor U25352 (N_25352,N_25168,N_25211);
and U25353 (N_25353,N_25025,N_25081);
nor U25354 (N_25354,N_25055,N_25060);
or U25355 (N_25355,N_25126,N_25119);
or U25356 (N_25356,N_25044,N_25090);
nor U25357 (N_25357,N_25176,N_25150);
xor U25358 (N_25358,N_25097,N_25157);
nor U25359 (N_25359,N_25091,N_25129);
nand U25360 (N_25360,N_25180,N_25054);
nor U25361 (N_25361,N_25116,N_25022);
xnor U25362 (N_25362,N_25171,N_25068);
nand U25363 (N_25363,N_25146,N_25018);
or U25364 (N_25364,N_25080,N_25248);
or U25365 (N_25365,N_25173,N_25172);
nand U25366 (N_25366,N_25102,N_25121);
or U25367 (N_25367,N_25035,N_25235);
nor U25368 (N_25368,N_25065,N_25075);
xor U25369 (N_25369,N_25008,N_25148);
and U25370 (N_25370,N_25213,N_25118);
xor U25371 (N_25371,N_25130,N_25140);
or U25372 (N_25372,N_25020,N_25153);
nand U25373 (N_25373,N_25113,N_25205);
xnor U25374 (N_25374,N_25225,N_25085);
or U25375 (N_25375,N_25212,N_25084);
xor U25376 (N_25376,N_25161,N_25050);
and U25377 (N_25377,N_25234,N_25124);
nor U25378 (N_25378,N_25179,N_25129);
or U25379 (N_25379,N_25038,N_25003);
nor U25380 (N_25380,N_25231,N_25012);
or U25381 (N_25381,N_25059,N_25196);
and U25382 (N_25382,N_25085,N_25000);
and U25383 (N_25383,N_25147,N_25212);
nor U25384 (N_25384,N_25146,N_25025);
xnor U25385 (N_25385,N_25012,N_25094);
nand U25386 (N_25386,N_25063,N_25052);
or U25387 (N_25387,N_25007,N_25182);
and U25388 (N_25388,N_25182,N_25201);
xor U25389 (N_25389,N_25074,N_25234);
or U25390 (N_25390,N_25074,N_25162);
and U25391 (N_25391,N_25236,N_25227);
xor U25392 (N_25392,N_25037,N_25245);
nand U25393 (N_25393,N_25067,N_25185);
xor U25394 (N_25394,N_25210,N_25002);
and U25395 (N_25395,N_25202,N_25060);
xor U25396 (N_25396,N_25155,N_25035);
nand U25397 (N_25397,N_25130,N_25008);
or U25398 (N_25398,N_25187,N_25096);
nor U25399 (N_25399,N_25010,N_25047);
or U25400 (N_25400,N_25124,N_25176);
or U25401 (N_25401,N_25127,N_25208);
and U25402 (N_25402,N_25220,N_25155);
nor U25403 (N_25403,N_25074,N_25174);
nand U25404 (N_25404,N_25108,N_25186);
nor U25405 (N_25405,N_25044,N_25227);
nand U25406 (N_25406,N_25206,N_25001);
and U25407 (N_25407,N_25106,N_25222);
or U25408 (N_25408,N_25070,N_25187);
or U25409 (N_25409,N_25007,N_25132);
nand U25410 (N_25410,N_25055,N_25110);
nand U25411 (N_25411,N_25089,N_25106);
and U25412 (N_25412,N_25160,N_25053);
or U25413 (N_25413,N_25011,N_25138);
and U25414 (N_25414,N_25001,N_25244);
or U25415 (N_25415,N_25185,N_25068);
nand U25416 (N_25416,N_25013,N_25054);
or U25417 (N_25417,N_25113,N_25000);
nand U25418 (N_25418,N_25194,N_25201);
nand U25419 (N_25419,N_25109,N_25189);
and U25420 (N_25420,N_25156,N_25032);
xnor U25421 (N_25421,N_25221,N_25097);
or U25422 (N_25422,N_25079,N_25094);
nand U25423 (N_25423,N_25071,N_25241);
nand U25424 (N_25424,N_25047,N_25144);
nand U25425 (N_25425,N_25165,N_25090);
nand U25426 (N_25426,N_25145,N_25095);
nand U25427 (N_25427,N_25091,N_25209);
nor U25428 (N_25428,N_25036,N_25052);
and U25429 (N_25429,N_25151,N_25070);
nor U25430 (N_25430,N_25229,N_25091);
nor U25431 (N_25431,N_25098,N_25048);
xnor U25432 (N_25432,N_25199,N_25206);
nor U25433 (N_25433,N_25221,N_25163);
nand U25434 (N_25434,N_25243,N_25163);
nor U25435 (N_25435,N_25120,N_25169);
and U25436 (N_25436,N_25078,N_25167);
and U25437 (N_25437,N_25227,N_25000);
xor U25438 (N_25438,N_25087,N_25071);
nor U25439 (N_25439,N_25247,N_25219);
xnor U25440 (N_25440,N_25232,N_25172);
xnor U25441 (N_25441,N_25112,N_25011);
xnor U25442 (N_25442,N_25058,N_25170);
xnor U25443 (N_25443,N_25085,N_25087);
and U25444 (N_25444,N_25051,N_25197);
or U25445 (N_25445,N_25010,N_25206);
or U25446 (N_25446,N_25232,N_25202);
nand U25447 (N_25447,N_25145,N_25087);
nor U25448 (N_25448,N_25089,N_25198);
and U25449 (N_25449,N_25190,N_25216);
xor U25450 (N_25450,N_25204,N_25047);
xor U25451 (N_25451,N_25209,N_25007);
or U25452 (N_25452,N_25115,N_25242);
nand U25453 (N_25453,N_25017,N_25097);
and U25454 (N_25454,N_25109,N_25120);
nor U25455 (N_25455,N_25061,N_25159);
nand U25456 (N_25456,N_25095,N_25143);
and U25457 (N_25457,N_25131,N_25028);
and U25458 (N_25458,N_25150,N_25189);
nand U25459 (N_25459,N_25101,N_25077);
nor U25460 (N_25460,N_25101,N_25179);
xnor U25461 (N_25461,N_25157,N_25087);
xor U25462 (N_25462,N_25237,N_25067);
or U25463 (N_25463,N_25224,N_25191);
nor U25464 (N_25464,N_25083,N_25030);
and U25465 (N_25465,N_25174,N_25143);
or U25466 (N_25466,N_25122,N_25046);
nor U25467 (N_25467,N_25235,N_25075);
or U25468 (N_25468,N_25035,N_25044);
nor U25469 (N_25469,N_25077,N_25074);
xnor U25470 (N_25470,N_25023,N_25127);
xnor U25471 (N_25471,N_25196,N_25175);
nor U25472 (N_25472,N_25074,N_25242);
nand U25473 (N_25473,N_25049,N_25018);
xor U25474 (N_25474,N_25073,N_25015);
or U25475 (N_25475,N_25149,N_25207);
or U25476 (N_25476,N_25057,N_25113);
xnor U25477 (N_25477,N_25001,N_25152);
and U25478 (N_25478,N_25143,N_25004);
or U25479 (N_25479,N_25048,N_25093);
and U25480 (N_25480,N_25017,N_25085);
nand U25481 (N_25481,N_25124,N_25030);
nor U25482 (N_25482,N_25139,N_25072);
and U25483 (N_25483,N_25220,N_25165);
xor U25484 (N_25484,N_25043,N_25004);
and U25485 (N_25485,N_25058,N_25222);
nand U25486 (N_25486,N_25145,N_25158);
or U25487 (N_25487,N_25059,N_25053);
nand U25488 (N_25488,N_25084,N_25104);
nor U25489 (N_25489,N_25113,N_25008);
nand U25490 (N_25490,N_25116,N_25136);
nand U25491 (N_25491,N_25192,N_25082);
nor U25492 (N_25492,N_25183,N_25225);
nand U25493 (N_25493,N_25098,N_25191);
nand U25494 (N_25494,N_25186,N_25248);
and U25495 (N_25495,N_25041,N_25106);
or U25496 (N_25496,N_25087,N_25131);
and U25497 (N_25497,N_25022,N_25018);
and U25498 (N_25498,N_25199,N_25192);
and U25499 (N_25499,N_25170,N_25182);
or U25500 (N_25500,N_25283,N_25462);
nor U25501 (N_25501,N_25435,N_25334);
nand U25502 (N_25502,N_25261,N_25320);
and U25503 (N_25503,N_25287,N_25436);
and U25504 (N_25504,N_25359,N_25487);
nand U25505 (N_25505,N_25361,N_25256);
or U25506 (N_25506,N_25338,N_25410);
or U25507 (N_25507,N_25270,N_25304);
nand U25508 (N_25508,N_25281,N_25385);
xor U25509 (N_25509,N_25279,N_25407);
xor U25510 (N_25510,N_25355,N_25346);
and U25511 (N_25511,N_25401,N_25404);
and U25512 (N_25512,N_25459,N_25384);
nand U25513 (N_25513,N_25329,N_25455);
nand U25514 (N_25514,N_25262,N_25305);
or U25515 (N_25515,N_25485,N_25483);
xnor U25516 (N_25516,N_25366,N_25426);
and U25517 (N_25517,N_25336,N_25491);
and U25518 (N_25518,N_25365,N_25448);
or U25519 (N_25519,N_25339,N_25343);
nand U25520 (N_25520,N_25431,N_25374);
nand U25521 (N_25521,N_25382,N_25432);
nor U25522 (N_25522,N_25379,N_25423);
or U25523 (N_25523,N_25497,N_25333);
or U25524 (N_25524,N_25417,N_25328);
nor U25525 (N_25525,N_25392,N_25367);
or U25526 (N_25526,N_25461,N_25416);
or U25527 (N_25527,N_25429,N_25450);
or U25528 (N_25528,N_25311,N_25332);
and U25529 (N_25529,N_25330,N_25280);
or U25530 (N_25530,N_25388,N_25399);
xor U25531 (N_25531,N_25495,N_25402);
xor U25532 (N_25532,N_25335,N_25299);
xnor U25533 (N_25533,N_25319,N_25327);
xor U25534 (N_25534,N_25493,N_25375);
nor U25535 (N_25535,N_25363,N_25378);
nor U25536 (N_25536,N_25425,N_25482);
or U25537 (N_25537,N_25460,N_25456);
and U25538 (N_25538,N_25389,N_25468);
xnor U25539 (N_25539,N_25325,N_25344);
and U25540 (N_25540,N_25427,N_25413);
and U25541 (N_25541,N_25323,N_25411);
or U25542 (N_25542,N_25386,N_25342);
and U25543 (N_25543,N_25472,N_25463);
nand U25544 (N_25544,N_25263,N_25418);
and U25545 (N_25545,N_25309,N_25394);
nand U25546 (N_25546,N_25358,N_25451);
xor U25547 (N_25547,N_25449,N_25318);
and U25548 (N_25548,N_25391,N_25293);
and U25549 (N_25549,N_25266,N_25443);
nor U25550 (N_25550,N_25422,N_25282);
nand U25551 (N_25551,N_25314,N_25369);
xnor U25552 (N_25552,N_25258,N_25254);
xor U25553 (N_25553,N_25364,N_25313);
nand U25554 (N_25554,N_25454,N_25446);
nor U25555 (N_25555,N_25352,N_25420);
and U25556 (N_25556,N_25277,N_25298);
nor U25557 (N_25557,N_25408,N_25381);
nand U25558 (N_25558,N_25347,N_25310);
xor U25559 (N_25559,N_25350,N_25296);
nor U25560 (N_25560,N_25373,N_25372);
and U25561 (N_25561,N_25295,N_25269);
nand U25562 (N_25562,N_25357,N_25253);
or U25563 (N_25563,N_25292,N_25438);
nor U25564 (N_25564,N_25396,N_25440);
or U25565 (N_25565,N_25437,N_25312);
nand U25566 (N_25566,N_25291,N_25405);
xor U25567 (N_25567,N_25273,N_25457);
xor U25568 (N_25568,N_25301,N_25272);
nand U25569 (N_25569,N_25471,N_25268);
nor U25570 (N_25570,N_25478,N_25479);
nand U25571 (N_25571,N_25286,N_25331);
or U25572 (N_25572,N_25419,N_25349);
and U25573 (N_25573,N_25289,N_25315);
or U25574 (N_25574,N_25288,N_25445);
xnor U25575 (N_25575,N_25345,N_25383);
xnor U25576 (N_25576,N_25257,N_25476);
or U25577 (N_25577,N_25467,N_25284);
xnor U25578 (N_25578,N_25424,N_25496);
xnor U25579 (N_25579,N_25481,N_25442);
and U25580 (N_25580,N_25341,N_25351);
nand U25581 (N_25581,N_25356,N_25492);
xor U25582 (N_25582,N_25326,N_25348);
nor U25583 (N_25583,N_25395,N_25477);
and U25584 (N_25584,N_25490,N_25360);
nand U25585 (N_25585,N_25294,N_25264);
nor U25586 (N_25586,N_25499,N_25397);
nor U25587 (N_25587,N_25473,N_25303);
xor U25588 (N_25588,N_25412,N_25469);
xnor U25589 (N_25589,N_25317,N_25362);
nand U25590 (N_25590,N_25453,N_25260);
nor U25591 (N_25591,N_25489,N_25465);
and U25592 (N_25592,N_25377,N_25337);
nand U25593 (N_25593,N_25406,N_25390);
xnor U25594 (N_25594,N_25444,N_25458);
or U25595 (N_25595,N_25316,N_25371);
nor U25596 (N_25596,N_25433,N_25308);
and U25597 (N_25597,N_25480,N_25421);
or U25598 (N_25598,N_25276,N_25409);
or U25599 (N_25599,N_25475,N_25354);
nand U25600 (N_25600,N_25259,N_25285);
or U25601 (N_25601,N_25484,N_25265);
xnor U25602 (N_25602,N_25474,N_25380);
and U25603 (N_25603,N_25403,N_25250);
nor U25604 (N_25604,N_25321,N_25466);
xnor U25605 (N_25605,N_25400,N_25439);
xnor U25606 (N_25606,N_25393,N_25353);
and U25607 (N_25607,N_25290,N_25252);
nand U25608 (N_25608,N_25452,N_25488);
xor U25609 (N_25609,N_25376,N_25274);
and U25610 (N_25610,N_25398,N_25255);
or U25611 (N_25611,N_25370,N_25322);
nor U25612 (N_25612,N_25278,N_25300);
nand U25613 (N_25613,N_25340,N_25324);
nand U25614 (N_25614,N_25306,N_25430);
xnor U25615 (N_25615,N_25251,N_25486);
and U25616 (N_25616,N_25441,N_25271);
xor U25617 (N_25617,N_25297,N_25414);
nand U25618 (N_25618,N_25464,N_25387);
and U25619 (N_25619,N_25267,N_25470);
or U25620 (N_25620,N_25307,N_25275);
xor U25621 (N_25621,N_25302,N_25415);
nor U25622 (N_25622,N_25434,N_25498);
or U25623 (N_25623,N_25447,N_25428);
xor U25624 (N_25624,N_25494,N_25368);
nor U25625 (N_25625,N_25387,N_25339);
nand U25626 (N_25626,N_25470,N_25373);
nor U25627 (N_25627,N_25414,N_25484);
nand U25628 (N_25628,N_25475,N_25337);
or U25629 (N_25629,N_25345,N_25398);
and U25630 (N_25630,N_25261,N_25334);
nand U25631 (N_25631,N_25284,N_25408);
nor U25632 (N_25632,N_25405,N_25431);
xnor U25633 (N_25633,N_25394,N_25262);
xnor U25634 (N_25634,N_25351,N_25289);
and U25635 (N_25635,N_25449,N_25360);
and U25636 (N_25636,N_25468,N_25387);
nand U25637 (N_25637,N_25309,N_25307);
and U25638 (N_25638,N_25270,N_25320);
or U25639 (N_25639,N_25400,N_25322);
nor U25640 (N_25640,N_25461,N_25463);
or U25641 (N_25641,N_25257,N_25496);
nand U25642 (N_25642,N_25379,N_25314);
nor U25643 (N_25643,N_25465,N_25415);
xor U25644 (N_25644,N_25260,N_25379);
or U25645 (N_25645,N_25447,N_25474);
and U25646 (N_25646,N_25274,N_25251);
nand U25647 (N_25647,N_25295,N_25466);
nand U25648 (N_25648,N_25356,N_25423);
or U25649 (N_25649,N_25272,N_25466);
and U25650 (N_25650,N_25458,N_25467);
or U25651 (N_25651,N_25342,N_25446);
xnor U25652 (N_25652,N_25492,N_25431);
and U25653 (N_25653,N_25343,N_25321);
or U25654 (N_25654,N_25278,N_25282);
nand U25655 (N_25655,N_25291,N_25368);
nand U25656 (N_25656,N_25442,N_25344);
and U25657 (N_25657,N_25331,N_25366);
xor U25658 (N_25658,N_25494,N_25305);
nand U25659 (N_25659,N_25361,N_25370);
or U25660 (N_25660,N_25287,N_25384);
or U25661 (N_25661,N_25445,N_25456);
and U25662 (N_25662,N_25432,N_25417);
and U25663 (N_25663,N_25384,N_25300);
and U25664 (N_25664,N_25269,N_25357);
nor U25665 (N_25665,N_25391,N_25435);
nand U25666 (N_25666,N_25406,N_25435);
and U25667 (N_25667,N_25361,N_25487);
nor U25668 (N_25668,N_25315,N_25413);
nor U25669 (N_25669,N_25418,N_25260);
nand U25670 (N_25670,N_25331,N_25411);
and U25671 (N_25671,N_25411,N_25415);
nor U25672 (N_25672,N_25350,N_25308);
xor U25673 (N_25673,N_25458,N_25445);
or U25674 (N_25674,N_25268,N_25261);
nor U25675 (N_25675,N_25365,N_25312);
nor U25676 (N_25676,N_25413,N_25354);
nor U25677 (N_25677,N_25474,N_25382);
and U25678 (N_25678,N_25315,N_25492);
and U25679 (N_25679,N_25399,N_25449);
nor U25680 (N_25680,N_25258,N_25274);
nand U25681 (N_25681,N_25251,N_25371);
nor U25682 (N_25682,N_25313,N_25345);
xnor U25683 (N_25683,N_25256,N_25423);
xor U25684 (N_25684,N_25420,N_25461);
and U25685 (N_25685,N_25375,N_25252);
nand U25686 (N_25686,N_25470,N_25309);
or U25687 (N_25687,N_25389,N_25251);
nor U25688 (N_25688,N_25489,N_25417);
or U25689 (N_25689,N_25436,N_25309);
nor U25690 (N_25690,N_25276,N_25444);
nor U25691 (N_25691,N_25288,N_25436);
nand U25692 (N_25692,N_25318,N_25252);
nand U25693 (N_25693,N_25390,N_25467);
nand U25694 (N_25694,N_25283,N_25340);
or U25695 (N_25695,N_25348,N_25302);
and U25696 (N_25696,N_25367,N_25464);
nor U25697 (N_25697,N_25457,N_25309);
nand U25698 (N_25698,N_25496,N_25457);
and U25699 (N_25699,N_25287,N_25355);
or U25700 (N_25700,N_25454,N_25466);
and U25701 (N_25701,N_25405,N_25469);
xnor U25702 (N_25702,N_25345,N_25472);
or U25703 (N_25703,N_25349,N_25314);
nand U25704 (N_25704,N_25437,N_25459);
nor U25705 (N_25705,N_25361,N_25262);
nor U25706 (N_25706,N_25321,N_25273);
nor U25707 (N_25707,N_25331,N_25302);
or U25708 (N_25708,N_25410,N_25342);
xor U25709 (N_25709,N_25418,N_25296);
or U25710 (N_25710,N_25374,N_25402);
nand U25711 (N_25711,N_25266,N_25370);
nor U25712 (N_25712,N_25443,N_25344);
xor U25713 (N_25713,N_25474,N_25354);
and U25714 (N_25714,N_25392,N_25372);
nor U25715 (N_25715,N_25495,N_25477);
nor U25716 (N_25716,N_25486,N_25490);
or U25717 (N_25717,N_25413,N_25408);
or U25718 (N_25718,N_25450,N_25421);
nand U25719 (N_25719,N_25297,N_25308);
xnor U25720 (N_25720,N_25445,N_25477);
and U25721 (N_25721,N_25407,N_25447);
xor U25722 (N_25722,N_25262,N_25338);
xor U25723 (N_25723,N_25486,N_25431);
or U25724 (N_25724,N_25298,N_25423);
nand U25725 (N_25725,N_25403,N_25388);
xnor U25726 (N_25726,N_25491,N_25334);
nand U25727 (N_25727,N_25270,N_25479);
xor U25728 (N_25728,N_25474,N_25374);
xnor U25729 (N_25729,N_25344,N_25389);
nand U25730 (N_25730,N_25263,N_25443);
nand U25731 (N_25731,N_25473,N_25267);
nand U25732 (N_25732,N_25266,N_25430);
nand U25733 (N_25733,N_25309,N_25317);
xor U25734 (N_25734,N_25440,N_25392);
nor U25735 (N_25735,N_25414,N_25454);
and U25736 (N_25736,N_25316,N_25399);
nand U25737 (N_25737,N_25409,N_25410);
or U25738 (N_25738,N_25485,N_25455);
or U25739 (N_25739,N_25265,N_25398);
xnor U25740 (N_25740,N_25280,N_25407);
nand U25741 (N_25741,N_25276,N_25384);
nor U25742 (N_25742,N_25395,N_25345);
nor U25743 (N_25743,N_25472,N_25391);
and U25744 (N_25744,N_25268,N_25266);
nor U25745 (N_25745,N_25473,N_25465);
and U25746 (N_25746,N_25452,N_25282);
or U25747 (N_25747,N_25291,N_25392);
xnor U25748 (N_25748,N_25388,N_25476);
xnor U25749 (N_25749,N_25408,N_25335);
nand U25750 (N_25750,N_25684,N_25546);
and U25751 (N_25751,N_25730,N_25689);
or U25752 (N_25752,N_25603,N_25548);
nand U25753 (N_25753,N_25588,N_25747);
nor U25754 (N_25754,N_25593,N_25652);
or U25755 (N_25755,N_25714,N_25649);
nor U25756 (N_25756,N_25519,N_25557);
and U25757 (N_25757,N_25637,N_25562);
or U25758 (N_25758,N_25582,N_25626);
nor U25759 (N_25759,N_25567,N_25718);
or U25760 (N_25760,N_25648,N_25625);
nor U25761 (N_25761,N_25712,N_25583);
and U25762 (N_25762,N_25550,N_25722);
or U25763 (N_25763,N_25622,N_25672);
and U25764 (N_25764,N_25655,N_25696);
nor U25765 (N_25765,N_25660,N_25690);
and U25766 (N_25766,N_25725,N_25563);
and U25767 (N_25767,N_25678,N_25579);
nand U25768 (N_25768,N_25573,N_25598);
and U25769 (N_25769,N_25701,N_25601);
or U25770 (N_25770,N_25527,N_25568);
and U25771 (N_25771,N_25732,N_25556);
xnor U25772 (N_25772,N_25552,N_25742);
or U25773 (N_25773,N_25572,N_25731);
nor U25774 (N_25774,N_25607,N_25728);
nor U25775 (N_25775,N_25615,N_25681);
or U25776 (N_25776,N_25659,N_25530);
nor U25777 (N_25777,N_25560,N_25570);
nor U25778 (N_25778,N_25636,N_25537);
nor U25779 (N_25779,N_25576,N_25506);
nor U25780 (N_25780,N_25736,N_25633);
nor U25781 (N_25781,N_25578,N_25707);
or U25782 (N_25782,N_25565,N_25710);
or U25783 (N_25783,N_25679,N_25638);
or U25784 (N_25784,N_25551,N_25629);
xnor U25785 (N_25785,N_25674,N_25535);
nor U25786 (N_25786,N_25726,N_25504);
or U25787 (N_25787,N_25713,N_25525);
xnor U25788 (N_25788,N_25580,N_25602);
and U25789 (N_25789,N_25585,N_25564);
and U25790 (N_25790,N_25640,N_25539);
nand U25791 (N_25791,N_25569,N_25665);
xnor U25792 (N_25792,N_25651,N_25555);
or U25793 (N_25793,N_25639,N_25597);
nand U25794 (N_25794,N_25677,N_25612);
xnor U25795 (N_25795,N_25592,N_25693);
and U25796 (N_25796,N_25610,N_25683);
and U25797 (N_25797,N_25514,N_25587);
and U25798 (N_25798,N_25536,N_25724);
or U25799 (N_25799,N_25661,N_25694);
nor U25800 (N_25800,N_25508,N_25618);
nand U25801 (N_25801,N_25513,N_25676);
or U25802 (N_25802,N_25520,N_25675);
xor U25803 (N_25803,N_25624,N_25616);
and U25804 (N_25804,N_25507,N_25631);
or U25805 (N_25805,N_25595,N_25687);
and U25806 (N_25806,N_25735,N_25542);
nor U25807 (N_25807,N_25549,N_25680);
and U25808 (N_25808,N_25748,N_25695);
or U25809 (N_25809,N_25518,N_25666);
and U25810 (N_25810,N_25511,N_25739);
or U25811 (N_25811,N_25554,N_25606);
nand U25812 (N_25812,N_25500,N_25531);
nand U25813 (N_25813,N_25643,N_25599);
nor U25814 (N_25814,N_25517,N_25503);
or U25815 (N_25815,N_25559,N_25737);
nor U25816 (N_25816,N_25526,N_25734);
xor U25817 (N_25817,N_25620,N_25682);
nor U25818 (N_25818,N_25541,N_25654);
or U25819 (N_25819,N_25529,N_25604);
nor U25820 (N_25820,N_25581,N_25609);
and U25821 (N_25821,N_25706,N_25749);
xnor U25822 (N_25822,N_25717,N_25711);
or U25823 (N_25823,N_25553,N_25703);
nand U25824 (N_25824,N_25729,N_25558);
and U25825 (N_25825,N_25591,N_25608);
and U25826 (N_25826,N_25670,N_25534);
or U25827 (N_25827,N_25611,N_25702);
or U25828 (N_25828,N_25613,N_25516);
or U25829 (N_25829,N_25692,N_25658);
or U25830 (N_25830,N_25574,N_25653);
nand U25831 (N_25831,N_25532,N_25662);
and U25832 (N_25832,N_25528,N_25547);
nand U25833 (N_25833,N_25708,N_25650);
and U25834 (N_25834,N_25575,N_25745);
or U25835 (N_25835,N_25627,N_25746);
nor U25836 (N_25836,N_25663,N_25720);
xor U25837 (N_25837,N_25614,N_25645);
xnor U25838 (N_25838,N_25538,N_25540);
nor U25839 (N_25839,N_25644,N_25719);
nand U25840 (N_25840,N_25727,N_25512);
nand U25841 (N_25841,N_25669,N_25630);
nand U25842 (N_25842,N_25740,N_25671);
xnor U25843 (N_25843,N_25571,N_25691);
nor U25844 (N_25844,N_25590,N_25664);
or U25845 (N_25845,N_25744,N_25617);
nor U25846 (N_25846,N_25586,N_25686);
nand U25847 (N_25847,N_25673,N_25515);
nor U25848 (N_25848,N_25619,N_25589);
or U25849 (N_25849,N_25741,N_25733);
or U25850 (N_25850,N_25688,N_25699);
or U25851 (N_25851,N_25698,N_25715);
or U25852 (N_25852,N_25566,N_25561);
and U25853 (N_25853,N_25621,N_25668);
xnor U25854 (N_25854,N_25646,N_25594);
nand U25855 (N_25855,N_25685,N_25605);
xnor U25856 (N_25856,N_25647,N_25501);
nand U25857 (N_25857,N_25544,N_25700);
and U25858 (N_25858,N_25667,N_25704);
or U25859 (N_25859,N_25596,N_25709);
or U25860 (N_25860,N_25628,N_25743);
nor U25861 (N_25861,N_25716,N_25533);
xor U25862 (N_25862,N_25656,N_25521);
or U25863 (N_25863,N_25524,N_25523);
nor U25864 (N_25864,N_25522,N_25509);
nand U25865 (N_25865,N_25641,N_25721);
or U25866 (N_25866,N_25584,N_25705);
or U25867 (N_25867,N_25600,N_25642);
and U25868 (N_25868,N_25738,N_25632);
nand U25869 (N_25869,N_25657,N_25505);
and U25870 (N_25870,N_25510,N_25623);
and U25871 (N_25871,N_25697,N_25577);
and U25872 (N_25872,N_25634,N_25502);
xnor U25873 (N_25873,N_25545,N_25543);
nand U25874 (N_25874,N_25723,N_25635);
xor U25875 (N_25875,N_25665,N_25669);
and U25876 (N_25876,N_25719,N_25625);
xor U25877 (N_25877,N_25612,N_25602);
xor U25878 (N_25878,N_25622,N_25568);
nor U25879 (N_25879,N_25712,N_25688);
or U25880 (N_25880,N_25741,N_25728);
nand U25881 (N_25881,N_25607,N_25739);
nor U25882 (N_25882,N_25727,N_25506);
nand U25883 (N_25883,N_25663,N_25670);
nand U25884 (N_25884,N_25564,N_25501);
nor U25885 (N_25885,N_25715,N_25704);
xor U25886 (N_25886,N_25725,N_25673);
nor U25887 (N_25887,N_25612,N_25525);
or U25888 (N_25888,N_25676,N_25506);
or U25889 (N_25889,N_25594,N_25628);
and U25890 (N_25890,N_25749,N_25503);
nor U25891 (N_25891,N_25584,N_25579);
or U25892 (N_25892,N_25693,N_25526);
nand U25893 (N_25893,N_25500,N_25628);
nand U25894 (N_25894,N_25667,N_25582);
nand U25895 (N_25895,N_25726,N_25612);
nand U25896 (N_25896,N_25700,N_25726);
nand U25897 (N_25897,N_25690,N_25510);
xnor U25898 (N_25898,N_25527,N_25638);
nor U25899 (N_25899,N_25560,N_25655);
and U25900 (N_25900,N_25577,N_25705);
xor U25901 (N_25901,N_25648,N_25610);
nand U25902 (N_25902,N_25582,N_25686);
nand U25903 (N_25903,N_25644,N_25621);
nand U25904 (N_25904,N_25611,N_25586);
nand U25905 (N_25905,N_25732,N_25590);
or U25906 (N_25906,N_25711,N_25619);
nand U25907 (N_25907,N_25547,N_25607);
nor U25908 (N_25908,N_25525,N_25571);
nand U25909 (N_25909,N_25678,N_25548);
nor U25910 (N_25910,N_25502,N_25621);
or U25911 (N_25911,N_25727,N_25682);
xnor U25912 (N_25912,N_25621,N_25734);
and U25913 (N_25913,N_25521,N_25633);
nand U25914 (N_25914,N_25697,N_25536);
nand U25915 (N_25915,N_25516,N_25541);
nand U25916 (N_25916,N_25593,N_25654);
and U25917 (N_25917,N_25657,N_25593);
and U25918 (N_25918,N_25517,N_25624);
nand U25919 (N_25919,N_25649,N_25700);
nand U25920 (N_25920,N_25509,N_25524);
xnor U25921 (N_25921,N_25544,N_25559);
and U25922 (N_25922,N_25561,N_25702);
or U25923 (N_25923,N_25564,N_25722);
xnor U25924 (N_25924,N_25548,N_25511);
nand U25925 (N_25925,N_25683,N_25705);
and U25926 (N_25926,N_25612,N_25532);
nor U25927 (N_25927,N_25723,N_25506);
and U25928 (N_25928,N_25705,N_25512);
nor U25929 (N_25929,N_25743,N_25741);
xor U25930 (N_25930,N_25530,N_25634);
and U25931 (N_25931,N_25615,N_25505);
xor U25932 (N_25932,N_25519,N_25729);
or U25933 (N_25933,N_25706,N_25639);
or U25934 (N_25934,N_25690,N_25624);
nand U25935 (N_25935,N_25650,N_25516);
xor U25936 (N_25936,N_25705,N_25533);
xor U25937 (N_25937,N_25547,N_25514);
nor U25938 (N_25938,N_25725,N_25522);
and U25939 (N_25939,N_25512,N_25523);
or U25940 (N_25940,N_25586,N_25595);
xnor U25941 (N_25941,N_25585,N_25591);
nand U25942 (N_25942,N_25601,N_25691);
or U25943 (N_25943,N_25592,N_25503);
xor U25944 (N_25944,N_25722,N_25749);
or U25945 (N_25945,N_25535,N_25679);
nand U25946 (N_25946,N_25579,N_25659);
xnor U25947 (N_25947,N_25512,N_25571);
nand U25948 (N_25948,N_25733,N_25624);
or U25949 (N_25949,N_25683,N_25702);
nor U25950 (N_25950,N_25670,N_25624);
and U25951 (N_25951,N_25731,N_25506);
nand U25952 (N_25952,N_25733,N_25570);
nand U25953 (N_25953,N_25728,N_25589);
or U25954 (N_25954,N_25686,N_25563);
nor U25955 (N_25955,N_25601,N_25747);
nand U25956 (N_25956,N_25606,N_25561);
or U25957 (N_25957,N_25705,N_25549);
nor U25958 (N_25958,N_25708,N_25571);
or U25959 (N_25959,N_25616,N_25595);
xor U25960 (N_25960,N_25624,N_25743);
and U25961 (N_25961,N_25660,N_25725);
nor U25962 (N_25962,N_25609,N_25608);
and U25963 (N_25963,N_25736,N_25511);
and U25964 (N_25964,N_25666,N_25726);
xnor U25965 (N_25965,N_25542,N_25652);
nand U25966 (N_25966,N_25624,N_25596);
nand U25967 (N_25967,N_25541,N_25539);
xor U25968 (N_25968,N_25689,N_25591);
xor U25969 (N_25969,N_25691,N_25670);
nand U25970 (N_25970,N_25661,N_25565);
nor U25971 (N_25971,N_25610,N_25532);
nor U25972 (N_25972,N_25655,N_25635);
nand U25973 (N_25973,N_25739,N_25664);
or U25974 (N_25974,N_25738,N_25688);
and U25975 (N_25975,N_25723,N_25609);
xnor U25976 (N_25976,N_25646,N_25746);
and U25977 (N_25977,N_25581,N_25637);
nor U25978 (N_25978,N_25526,N_25609);
nor U25979 (N_25979,N_25594,N_25657);
nor U25980 (N_25980,N_25524,N_25584);
nand U25981 (N_25981,N_25740,N_25535);
and U25982 (N_25982,N_25660,N_25603);
nor U25983 (N_25983,N_25703,N_25713);
nor U25984 (N_25984,N_25638,N_25736);
nand U25985 (N_25985,N_25643,N_25720);
or U25986 (N_25986,N_25744,N_25630);
and U25987 (N_25987,N_25653,N_25576);
nor U25988 (N_25988,N_25700,N_25709);
and U25989 (N_25989,N_25502,N_25660);
xnor U25990 (N_25990,N_25669,N_25539);
nor U25991 (N_25991,N_25651,N_25578);
xnor U25992 (N_25992,N_25638,N_25568);
or U25993 (N_25993,N_25737,N_25538);
and U25994 (N_25994,N_25661,N_25710);
xor U25995 (N_25995,N_25733,N_25569);
nand U25996 (N_25996,N_25601,N_25528);
nand U25997 (N_25997,N_25704,N_25500);
xnor U25998 (N_25998,N_25726,N_25515);
nand U25999 (N_25999,N_25576,N_25574);
or U26000 (N_26000,N_25955,N_25802);
nor U26001 (N_26001,N_25757,N_25970);
and U26002 (N_26002,N_25929,N_25959);
xor U26003 (N_26003,N_25886,N_25811);
nand U26004 (N_26004,N_25977,N_25779);
nand U26005 (N_26005,N_25855,N_25760);
nand U26006 (N_26006,N_25922,N_25763);
nor U26007 (N_26007,N_25989,N_25917);
and U26008 (N_26008,N_25883,N_25775);
nor U26009 (N_26009,N_25828,N_25780);
xor U26010 (N_26010,N_25964,N_25909);
nor U26011 (N_26011,N_25818,N_25856);
or U26012 (N_26012,N_25822,N_25918);
and U26013 (N_26013,N_25840,N_25995);
or U26014 (N_26014,N_25801,N_25889);
nor U26015 (N_26015,N_25887,N_25876);
and U26016 (N_26016,N_25846,N_25994);
or U26017 (N_26017,N_25902,N_25864);
or U26018 (N_26018,N_25903,N_25753);
or U26019 (N_26019,N_25860,N_25789);
nor U26020 (N_26020,N_25915,N_25784);
xnor U26021 (N_26021,N_25971,N_25859);
nor U26022 (N_26022,N_25892,N_25940);
and U26023 (N_26023,N_25999,N_25987);
or U26024 (N_26024,N_25952,N_25793);
nand U26025 (N_26025,N_25881,N_25783);
nor U26026 (N_26026,N_25895,N_25978);
or U26027 (N_26027,N_25849,N_25824);
nor U26028 (N_26028,N_25821,N_25945);
nand U26029 (N_26029,N_25804,N_25782);
or U26030 (N_26030,N_25930,N_25815);
nor U26031 (N_26031,N_25936,N_25773);
or U26032 (N_26032,N_25799,N_25877);
or U26033 (N_26033,N_25816,N_25997);
and U26034 (N_26034,N_25831,N_25944);
or U26035 (N_26035,N_25866,N_25991);
nor U26036 (N_26036,N_25845,N_25833);
or U26037 (N_26037,N_25812,N_25869);
and U26038 (N_26038,N_25872,N_25847);
nor U26039 (N_26039,N_25981,N_25858);
xor U26040 (N_26040,N_25848,N_25838);
xor U26041 (N_26041,N_25751,N_25950);
and U26042 (N_26042,N_25862,N_25755);
nor U26043 (N_26043,N_25960,N_25853);
and U26044 (N_26044,N_25830,N_25919);
nor U26045 (N_26045,N_25974,N_25980);
and U26046 (N_26046,N_25770,N_25958);
or U26047 (N_26047,N_25946,N_25901);
and U26048 (N_26048,N_25907,N_25916);
xor U26049 (N_26049,N_25820,N_25905);
xor U26050 (N_26050,N_25809,N_25835);
nor U26051 (N_26051,N_25879,N_25867);
and U26052 (N_26052,N_25928,N_25827);
and U26053 (N_26053,N_25988,N_25888);
nand U26054 (N_26054,N_25943,N_25957);
nand U26055 (N_26055,N_25932,N_25985);
xnor U26056 (N_26056,N_25885,N_25948);
nor U26057 (N_26057,N_25826,N_25898);
nand U26058 (N_26058,N_25756,N_25842);
nand U26059 (N_26059,N_25899,N_25914);
and U26060 (N_26060,N_25857,N_25781);
nand U26061 (N_26061,N_25807,N_25976);
or U26062 (N_26062,N_25990,N_25806);
and U26063 (N_26063,N_25754,N_25800);
nand U26064 (N_26064,N_25777,N_25787);
and U26065 (N_26065,N_25832,N_25951);
nand U26066 (N_26066,N_25984,N_25791);
or U26067 (N_26067,N_25837,N_25967);
xnor U26068 (N_26068,N_25942,N_25759);
nor U26069 (N_26069,N_25794,N_25891);
nor U26070 (N_26070,N_25873,N_25844);
xor U26071 (N_26071,N_25774,N_25851);
nor U26072 (N_26072,N_25954,N_25772);
or U26073 (N_26073,N_25797,N_25813);
xnor U26074 (N_26074,N_25874,N_25910);
or U26075 (N_26075,N_25765,N_25850);
and U26076 (N_26076,N_25893,N_25785);
nor U26077 (N_26077,N_25920,N_25923);
nand U26078 (N_26078,N_25788,N_25803);
nor U26079 (N_26079,N_25966,N_25897);
nor U26080 (N_26080,N_25947,N_25817);
xor U26081 (N_26081,N_25894,N_25761);
xnor U26082 (N_26082,N_25839,N_25998);
and U26083 (N_26083,N_25776,N_25939);
xnor U26084 (N_26084,N_25805,N_25882);
xor U26085 (N_26085,N_25834,N_25829);
xnor U26086 (N_26086,N_25854,N_25852);
nand U26087 (N_26087,N_25863,N_25979);
or U26088 (N_26088,N_25778,N_25972);
or U26089 (N_26089,N_25975,N_25973);
nand U26090 (N_26090,N_25758,N_25880);
nand U26091 (N_26091,N_25961,N_25836);
nor U26092 (N_26092,N_25884,N_25769);
nand U26093 (N_26093,N_25871,N_25941);
nor U26094 (N_26094,N_25870,N_25968);
nand U26095 (N_26095,N_25878,N_25904);
and U26096 (N_26096,N_25982,N_25993);
or U26097 (N_26097,N_25906,N_25992);
and U26098 (N_26098,N_25790,N_25956);
or U26099 (N_26099,N_25931,N_25911);
nor U26100 (N_26100,N_25771,N_25814);
nor U26101 (N_26101,N_25927,N_25896);
nand U26102 (N_26102,N_25819,N_25768);
nand U26103 (N_26103,N_25865,N_25937);
and U26104 (N_26104,N_25933,N_25921);
xor U26105 (N_26105,N_25764,N_25949);
or U26106 (N_26106,N_25925,N_25752);
nor U26107 (N_26107,N_25963,N_25926);
nand U26108 (N_26108,N_25841,N_25934);
nor U26109 (N_26109,N_25935,N_25750);
xnor U26110 (N_26110,N_25969,N_25861);
or U26111 (N_26111,N_25983,N_25767);
and U26112 (N_26112,N_25938,N_25986);
nor U26113 (N_26113,N_25962,N_25965);
xor U26114 (N_26114,N_25766,N_25908);
or U26115 (N_26115,N_25868,N_25796);
and U26116 (N_26116,N_25762,N_25843);
xor U26117 (N_26117,N_25792,N_25924);
nor U26118 (N_26118,N_25808,N_25786);
nor U26119 (N_26119,N_25875,N_25810);
xnor U26120 (N_26120,N_25996,N_25912);
nor U26121 (N_26121,N_25798,N_25913);
nor U26122 (N_26122,N_25795,N_25900);
or U26123 (N_26123,N_25953,N_25823);
nand U26124 (N_26124,N_25890,N_25825);
nor U26125 (N_26125,N_25937,N_25838);
xnor U26126 (N_26126,N_25754,N_25768);
xnor U26127 (N_26127,N_25829,N_25984);
and U26128 (N_26128,N_25798,N_25926);
nand U26129 (N_26129,N_25779,N_25970);
nor U26130 (N_26130,N_25875,N_25936);
nand U26131 (N_26131,N_25914,N_25872);
xnor U26132 (N_26132,N_25853,N_25974);
nor U26133 (N_26133,N_25908,N_25994);
nor U26134 (N_26134,N_25827,N_25876);
nand U26135 (N_26135,N_25788,N_25945);
nand U26136 (N_26136,N_25884,N_25761);
and U26137 (N_26137,N_25846,N_25794);
nand U26138 (N_26138,N_25790,N_25876);
nor U26139 (N_26139,N_25816,N_25862);
and U26140 (N_26140,N_25949,N_25945);
and U26141 (N_26141,N_25918,N_25893);
xnor U26142 (N_26142,N_25845,N_25836);
nor U26143 (N_26143,N_25930,N_25911);
nor U26144 (N_26144,N_25826,N_25783);
nand U26145 (N_26145,N_25772,N_25935);
or U26146 (N_26146,N_25762,N_25771);
or U26147 (N_26147,N_25894,N_25990);
nor U26148 (N_26148,N_25878,N_25893);
nor U26149 (N_26149,N_25875,N_25768);
nand U26150 (N_26150,N_25775,N_25928);
and U26151 (N_26151,N_25870,N_25856);
nor U26152 (N_26152,N_25931,N_25800);
xor U26153 (N_26153,N_25847,N_25848);
or U26154 (N_26154,N_25813,N_25863);
xor U26155 (N_26155,N_25777,N_25845);
and U26156 (N_26156,N_25755,N_25925);
and U26157 (N_26157,N_25892,N_25792);
xor U26158 (N_26158,N_25942,N_25986);
xor U26159 (N_26159,N_25869,N_25923);
or U26160 (N_26160,N_25823,N_25861);
nand U26161 (N_26161,N_25843,N_25858);
xnor U26162 (N_26162,N_25750,N_25844);
or U26163 (N_26163,N_25825,N_25850);
nand U26164 (N_26164,N_25961,N_25925);
and U26165 (N_26165,N_25753,N_25867);
nor U26166 (N_26166,N_25750,N_25887);
nor U26167 (N_26167,N_25776,N_25847);
or U26168 (N_26168,N_25840,N_25991);
xnor U26169 (N_26169,N_25868,N_25911);
xnor U26170 (N_26170,N_25891,N_25970);
and U26171 (N_26171,N_25947,N_25815);
or U26172 (N_26172,N_25830,N_25761);
nor U26173 (N_26173,N_25907,N_25839);
xnor U26174 (N_26174,N_25932,N_25930);
xor U26175 (N_26175,N_25836,N_25969);
nor U26176 (N_26176,N_25799,N_25872);
or U26177 (N_26177,N_25757,N_25760);
xor U26178 (N_26178,N_25955,N_25755);
or U26179 (N_26179,N_25921,N_25758);
or U26180 (N_26180,N_25986,N_25903);
nand U26181 (N_26181,N_25764,N_25921);
xor U26182 (N_26182,N_25776,N_25827);
or U26183 (N_26183,N_25954,N_25909);
and U26184 (N_26184,N_25877,N_25763);
or U26185 (N_26185,N_25905,N_25947);
and U26186 (N_26186,N_25834,N_25896);
and U26187 (N_26187,N_25994,N_25785);
nand U26188 (N_26188,N_25957,N_25789);
and U26189 (N_26189,N_25970,N_25817);
and U26190 (N_26190,N_25969,N_25937);
nor U26191 (N_26191,N_25879,N_25844);
or U26192 (N_26192,N_25847,N_25972);
and U26193 (N_26193,N_25952,N_25873);
xnor U26194 (N_26194,N_25757,N_25873);
nand U26195 (N_26195,N_25951,N_25952);
or U26196 (N_26196,N_25947,N_25808);
nand U26197 (N_26197,N_25816,N_25773);
and U26198 (N_26198,N_25768,N_25841);
nor U26199 (N_26199,N_25956,N_25946);
and U26200 (N_26200,N_25942,N_25833);
and U26201 (N_26201,N_25822,N_25905);
and U26202 (N_26202,N_25861,N_25856);
and U26203 (N_26203,N_25798,N_25753);
and U26204 (N_26204,N_25905,N_25945);
nor U26205 (N_26205,N_25789,N_25759);
xor U26206 (N_26206,N_25872,N_25756);
and U26207 (N_26207,N_25871,N_25838);
and U26208 (N_26208,N_25806,N_25801);
nor U26209 (N_26209,N_25848,N_25978);
and U26210 (N_26210,N_25786,N_25963);
xor U26211 (N_26211,N_25898,N_25801);
nand U26212 (N_26212,N_25913,N_25997);
or U26213 (N_26213,N_25779,N_25751);
nand U26214 (N_26214,N_25878,N_25949);
xnor U26215 (N_26215,N_25843,N_25929);
nand U26216 (N_26216,N_25871,N_25844);
and U26217 (N_26217,N_25882,N_25756);
nor U26218 (N_26218,N_25758,N_25913);
or U26219 (N_26219,N_25976,N_25882);
or U26220 (N_26220,N_25895,N_25992);
nand U26221 (N_26221,N_25813,N_25895);
or U26222 (N_26222,N_25855,N_25823);
or U26223 (N_26223,N_25945,N_25924);
nand U26224 (N_26224,N_25850,N_25986);
or U26225 (N_26225,N_25779,N_25999);
xnor U26226 (N_26226,N_25884,N_25929);
and U26227 (N_26227,N_25932,N_25968);
nand U26228 (N_26228,N_25850,N_25766);
nand U26229 (N_26229,N_25775,N_25789);
xnor U26230 (N_26230,N_25928,N_25881);
and U26231 (N_26231,N_25985,N_25815);
nand U26232 (N_26232,N_25875,N_25970);
nor U26233 (N_26233,N_25922,N_25823);
or U26234 (N_26234,N_25819,N_25832);
xnor U26235 (N_26235,N_25803,N_25974);
nor U26236 (N_26236,N_25750,N_25775);
and U26237 (N_26237,N_25824,N_25868);
nor U26238 (N_26238,N_25833,N_25793);
nand U26239 (N_26239,N_25811,N_25788);
or U26240 (N_26240,N_25918,N_25764);
and U26241 (N_26241,N_25935,N_25955);
nand U26242 (N_26242,N_25963,N_25830);
nand U26243 (N_26243,N_25884,N_25791);
and U26244 (N_26244,N_25866,N_25796);
nand U26245 (N_26245,N_25911,N_25900);
xnor U26246 (N_26246,N_25964,N_25773);
xnor U26247 (N_26247,N_25807,N_25842);
nor U26248 (N_26248,N_25810,N_25893);
and U26249 (N_26249,N_25868,N_25872);
and U26250 (N_26250,N_26167,N_26054);
xor U26251 (N_26251,N_26012,N_26169);
or U26252 (N_26252,N_26162,N_26112);
or U26253 (N_26253,N_26065,N_26014);
nand U26254 (N_26254,N_26066,N_26021);
and U26255 (N_26255,N_26027,N_26038);
nor U26256 (N_26256,N_26024,N_26108);
xor U26257 (N_26257,N_26061,N_26222);
xnor U26258 (N_26258,N_26089,N_26033);
and U26259 (N_26259,N_26000,N_26225);
nor U26260 (N_26260,N_26107,N_26182);
xor U26261 (N_26261,N_26245,N_26010);
nand U26262 (N_26262,N_26045,N_26181);
nor U26263 (N_26263,N_26177,N_26067);
and U26264 (N_26264,N_26221,N_26140);
nand U26265 (N_26265,N_26151,N_26039);
xor U26266 (N_26266,N_26059,N_26204);
or U26267 (N_26267,N_26217,N_26088);
or U26268 (N_26268,N_26147,N_26022);
or U26269 (N_26269,N_26043,N_26034);
nor U26270 (N_26270,N_26133,N_26243);
and U26271 (N_26271,N_26226,N_26073);
xnor U26272 (N_26272,N_26083,N_26068);
or U26273 (N_26273,N_26080,N_26161);
xnor U26274 (N_26274,N_26192,N_26241);
nand U26275 (N_26275,N_26050,N_26053);
nand U26276 (N_26276,N_26145,N_26219);
and U26277 (N_26277,N_26238,N_26002);
nor U26278 (N_26278,N_26207,N_26017);
xor U26279 (N_26279,N_26004,N_26086);
and U26280 (N_26280,N_26110,N_26224);
nor U26281 (N_26281,N_26214,N_26117);
and U26282 (N_26282,N_26212,N_26157);
nand U26283 (N_26283,N_26101,N_26160);
nor U26284 (N_26284,N_26206,N_26098);
xnor U26285 (N_26285,N_26114,N_26006);
nor U26286 (N_26286,N_26023,N_26058);
or U26287 (N_26287,N_26173,N_26210);
xor U26288 (N_26288,N_26248,N_26148);
or U26289 (N_26289,N_26227,N_26247);
and U26290 (N_26290,N_26026,N_26116);
xnor U26291 (N_26291,N_26115,N_26146);
nor U26292 (N_26292,N_26163,N_26168);
or U26293 (N_26293,N_26049,N_26103);
or U26294 (N_26294,N_26082,N_26190);
nor U26295 (N_26295,N_26239,N_26183);
nand U26296 (N_26296,N_26121,N_26235);
and U26297 (N_26297,N_26104,N_26005);
or U26298 (N_26298,N_26109,N_26020);
nand U26299 (N_26299,N_26075,N_26209);
and U26300 (N_26300,N_26134,N_26159);
xnor U26301 (N_26301,N_26123,N_26124);
nand U26302 (N_26302,N_26019,N_26172);
xor U26303 (N_26303,N_26113,N_26102);
xor U26304 (N_26304,N_26051,N_26071);
nor U26305 (N_26305,N_26196,N_26249);
or U26306 (N_26306,N_26037,N_26072);
or U26307 (N_26307,N_26223,N_26186);
nor U26308 (N_26308,N_26074,N_26197);
xnor U26309 (N_26309,N_26236,N_26200);
and U26310 (N_26310,N_26127,N_26139);
nor U26311 (N_26311,N_26091,N_26016);
xnor U26312 (N_26312,N_26048,N_26090);
xor U26313 (N_26313,N_26057,N_26141);
and U26314 (N_26314,N_26211,N_26137);
and U26315 (N_26315,N_26240,N_26152);
xor U26316 (N_26316,N_26205,N_26085);
and U26317 (N_26317,N_26164,N_26009);
nor U26318 (N_26318,N_26001,N_26111);
or U26319 (N_26319,N_26078,N_26025);
nor U26320 (N_26320,N_26191,N_26178);
nand U26321 (N_26321,N_26097,N_26105);
and U26322 (N_26322,N_26220,N_26188);
or U26323 (N_26323,N_26120,N_26154);
xnor U26324 (N_26324,N_26150,N_26234);
or U26325 (N_26325,N_26063,N_26093);
xnor U26326 (N_26326,N_26047,N_26184);
nor U26327 (N_26327,N_26099,N_26155);
and U26328 (N_26328,N_26230,N_26062);
or U26329 (N_26329,N_26041,N_26171);
or U26330 (N_26330,N_26028,N_26128);
nor U26331 (N_26331,N_26144,N_26052);
or U26332 (N_26332,N_26189,N_26199);
and U26333 (N_26333,N_26198,N_26084);
nor U26334 (N_26334,N_26011,N_26203);
xnor U26335 (N_26335,N_26100,N_26081);
nand U26336 (N_26336,N_26046,N_26180);
or U26337 (N_26337,N_26237,N_26216);
nand U26338 (N_26338,N_26193,N_26179);
or U26339 (N_26339,N_26032,N_26044);
nor U26340 (N_26340,N_26218,N_26035);
and U26341 (N_26341,N_26158,N_26018);
nand U26342 (N_26342,N_26185,N_26246);
or U26343 (N_26343,N_26030,N_26132);
xnor U26344 (N_26344,N_26228,N_26142);
nand U26345 (N_26345,N_26095,N_26013);
or U26346 (N_26346,N_26231,N_26092);
xnor U26347 (N_26347,N_26215,N_26036);
nand U26348 (N_26348,N_26208,N_26143);
or U26349 (N_26349,N_26242,N_26055);
and U26350 (N_26350,N_26138,N_26126);
nor U26351 (N_26351,N_26229,N_26119);
and U26352 (N_26352,N_26056,N_26202);
nand U26353 (N_26353,N_26076,N_26176);
nand U26354 (N_26354,N_26125,N_26060);
xor U26355 (N_26355,N_26031,N_26118);
and U26356 (N_26356,N_26015,N_26106);
nand U26357 (N_26357,N_26070,N_26187);
and U26358 (N_26358,N_26003,N_26007);
nor U26359 (N_26359,N_26233,N_26165);
nand U26360 (N_26360,N_26213,N_26087);
nor U26361 (N_26361,N_26194,N_26131);
or U26362 (N_26362,N_26096,N_26029);
nor U26363 (N_26363,N_26153,N_26069);
or U26364 (N_26364,N_26201,N_26170);
and U26365 (N_26365,N_26232,N_26166);
and U26366 (N_26366,N_26042,N_26122);
nand U26367 (N_26367,N_26135,N_26077);
or U26368 (N_26368,N_26008,N_26136);
nand U26369 (N_26369,N_26094,N_26064);
and U26370 (N_26370,N_26195,N_26130);
nor U26371 (N_26371,N_26156,N_26244);
nand U26372 (N_26372,N_26175,N_26149);
or U26373 (N_26373,N_26129,N_26040);
or U26374 (N_26374,N_26174,N_26079);
nor U26375 (N_26375,N_26018,N_26019);
nand U26376 (N_26376,N_26190,N_26033);
xnor U26377 (N_26377,N_26094,N_26044);
and U26378 (N_26378,N_26036,N_26202);
or U26379 (N_26379,N_26110,N_26245);
xor U26380 (N_26380,N_26094,N_26003);
or U26381 (N_26381,N_26002,N_26152);
nand U26382 (N_26382,N_26210,N_26122);
nand U26383 (N_26383,N_26059,N_26183);
xnor U26384 (N_26384,N_26110,N_26175);
nand U26385 (N_26385,N_26071,N_26158);
and U26386 (N_26386,N_26114,N_26086);
and U26387 (N_26387,N_26071,N_26034);
and U26388 (N_26388,N_26074,N_26209);
and U26389 (N_26389,N_26153,N_26104);
xnor U26390 (N_26390,N_26113,N_26002);
nand U26391 (N_26391,N_26048,N_26118);
and U26392 (N_26392,N_26014,N_26172);
xnor U26393 (N_26393,N_26215,N_26073);
and U26394 (N_26394,N_26133,N_26226);
xnor U26395 (N_26395,N_26038,N_26182);
and U26396 (N_26396,N_26249,N_26244);
and U26397 (N_26397,N_26124,N_26015);
and U26398 (N_26398,N_26216,N_26242);
nor U26399 (N_26399,N_26043,N_26082);
or U26400 (N_26400,N_26046,N_26226);
xor U26401 (N_26401,N_26178,N_26108);
nor U26402 (N_26402,N_26127,N_26210);
nor U26403 (N_26403,N_26195,N_26064);
nand U26404 (N_26404,N_26176,N_26111);
nor U26405 (N_26405,N_26136,N_26170);
or U26406 (N_26406,N_26206,N_26144);
nor U26407 (N_26407,N_26160,N_26055);
nand U26408 (N_26408,N_26102,N_26120);
nand U26409 (N_26409,N_26041,N_26130);
nand U26410 (N_26410,N_26149,N_26044);
nor U26411 (N_26411,N_26066,N_26093);
nand U26412 (N_26412,N_26119,N_26051);
or U26413 (N_26413,N_26039,N_26193);
nor U26414 (N_26414,N_26041,N_26136);
nand U26415 (N_26415,N_26000,N_26159);
nor U26416 (N_26416,N_26123,N_26121);
or U26417 (N_26417,N_26133,N_26056);
xnor U26418 (N_26418,N_26185,N_26191);
nand U26419 (N_26419,N_26249,N_26226);
nor U26420 (N_26420,N_26074,N_26107);
nor U26421 (N_26421,N_26233,N_26167);
or U26422 (N_26422,N_26122,N_26023);
nor U26423 (N_26423,N_26195,N_26043);
nand U26424 (N_26424,N_26103,N_26215);
and U26425 (N_26425,N_26121,N_26051);
nand U26426 (N_26426,N_26086,N_26133);
xor U26427 (N_26427,N_26213,N_26012);
or U26428 (N_26428,N_26056,N_26222);
xnor U26429 (N_26429,N_26081,N_26058);
nor U26430 (N_26430,N_26063,N_26026);
xor U26431 (N_26431,N_26216,N_26227);
xnor U26432 (N_26432,N_26002,N_26151);
and U26433 (N_26433,N_26112,N_26048);
nand U26434 (N_26434,N_26095,N_26066);
or U26435 (N_26435,N_26050,N_26173);
and U26436 (N_26436,N_26111,N_26144);
or U26437 (N_26437,N_26001,N_26101);
or U26438 (N_26438,N_26167,N_26183);
or U26439 (N_26439,N_26005,N_26241);
nand U26440 (N_26440,N_26080,N_26157);
and U26441 (N_26441,N_26056,N_26163);
and U26442 (N_26442,N_26040,N_26063);
xnor U26443 (N_26443,N_26198,N_26110);
nand U26444 (N_26444,N_26240,N_26089);
nor U26445 (N_26445,N_26226,N_26115);
or U26446 (N_26446,N_26158,N_26195);
nand U26447 (N_26447,N_26196,N_26029);
nor U26448 (N_26448,N_26172,N_26017);
or U26449 (N_26449,N_26194,N_26226);
xnor U26450 (N_26450,N_26087,N_26187);
nand U26451 (N_26451,N_26110,N_26006);
and U26452 (N_26452,N_26032,N_26225);
nand U26453 (N_26453,N_26189,N_26031);
or U26454 (N_26454,N_26237,N_26166);
nor U26455 (N_26455,N_26025,N_26198);
and U26456 (N_26456,N_26067,N_26111);
nand U26457 (N_26457,N_26029,N_26184);
xnor U26458 (N_26458,N_26036,N_26102);
nand U26459 (N_26459,N_26163,N_26221);
xnor U26460 (N_26460,N_26102,N_26061);
xnor U26461 (N_26461,N_26216,N_26012);
or U26462 (N_26462,N_26228,N_26135);
xor U26463 (N_26463,N_26241,N_26184);
nand U26464 (N_26464,N_26061,N_26069);
nand U26465 (N_26465,N_26178,N_26182);
nand U26466 (N_26466,N_26078,N_26205);
and U26467 (N_26467,N_26227,N_26164);
xnor U26468 (N_26468,N_26087,N_26056);
or U26469 (N_26469,N_26009,N_26004);
and U26470 (N_26470,N_26024,N_26087);
nand U26471 (N_26471,N_26112,N_26050);
nand U26472 (N_26472,N_26105,N_26141);
nor U26473 (N_26473,N_26139,N_26237);
xor U26474 (N_26474,N_26189,N_26172);
and U26475 (N_26475,N_26236,N_26052);
or U26476 (N_26476,N_26110,N_26021);
nor U26477 (N_26477,N_26238,N_26092);
and U26478 (N_26478,N_26078,N_26150);
xor U26479 (N_26479,N_26197,N_26228);
or U26480 (N_26480,N_26000,N_26169);
nor U26481 (N_26481,N_26009,N_26012);
nor U26482 (N_26482,N_26063,N_26043);
xor U26483 (N_26483,N_26203,N_26070);
nor U26484 (N_26484,N_26104,N_26102);
and U26485 (N_26485,N_26210,N_26221);
nand U26486 (N_26486,N_26191,N_26094);
xnor U26487 (N_26487,N_26002,N_26170);
and U26488 (N_26488,N_26199,N_26238);
or U26489 (N_26489,N_26148,N_26129);
nand U26490 (N_26490,N_26139,N_26094);
nor U26491 (N_26491,N_26115,N_26070);
or U26492 (N_26492,N_26175,N_26171);
or U26493 (N_26493,N_26040,N_26182);
and U26494 (N_26494,N_26066,N_26185);
and U26495 (N_26495,N_26023,N_26094);
xnor U26496 (N_26496,N_26220,N_26180);
xnor U26497 (N_26497,N_26066,N_26068);
or U26498 (N_26498,N_26048,N_26050);
or U26499 (N_26499,N_26223,N_26233);
nor U26500 (N_26500,N_26366,N_26460);
nand U26501 (N_26501,N_26308,N_26318);
and U26502 (N_26502,N_26386,N_26383);
nand U26503 (N_26503,N_26401,N_26255);
and U26504 (N_26504,N_26341,N_26471);
xor U26505 (N_26505,N_26440,N_26320);
xnor U26506 (N_26506,N_26497,N_26419);
nor U26507 (N_26507,N_26448,N_26380);
and U26508 (N_26508,N_26256,N_26283);
xor U26509 (N_26509,N_26420,N_26319);
nand U26510 (N_26510,N_26357,N_26444);
nand U26511 (N_26511,N_26381,N_26262);
nand U26512 (N_26512,N_26391,N_26402);
nor U26513 (N_26513,N_26332,N_26297);
nand U26514 (N_26514,N_26446,N_26355);
and U26515 (N_26515,N_26483,N_26323);
or U26516 (N_26516,N_26315,N_26378);
and U26517 (N_26517,N_26447,N_26451);
and U26518 (N_26518,N_26266,N_26275);
and U26519 (N_26519,N_26480,N_26331);
nand U26520 (N_26520,N_26409,N_26470);
nor U26521 (N_26521,N_26410,N_26449);
xnor U26522 (N_26522,N_26426,N_26258);
and U26523 (N_26523,N_26389,N_26476);
or U26524 (N_26524,N_26488,N_26345);
or U26525 (N_26525,N_26379,N_26423);
nor U26526 (N_26526,N_26272,N_26414);
and U26527 (N_26527,N_26385,N_26435);
or U26528 (N_26528,N_26392,N_26282);
nand U26529 (N_26529,N_26362,N_26291);
xnor U26530 (N_26530,N_26454,N_26493);
and U26531 (N_26531,N_26344,N_26261);
nor U26532 (N_26532,N_26382,N_26350);
nor U26533 (N_26533,N_26431,N_26399);
nor U26534 (N_26534,N_26430,N_26356);
or U26535 (N_26535,N_26418,N_26474);
nand U26536 (N_26536,N_26374,N_26330);
and U26537 (N_26537,N_26364,N_26496);
and U26538 (N_26538,N_26398,N_26264);
nand U26539 (N_26539,N_26433,N_26333);
nor U26540 (N_26540,N_26478,N_26343);
nor U26541 (N_26541,N_26462,N_26427);
and U26542 (N_26542,N_26481,N_26295);
and U26543 (N_26543,N_26473,N_26280);
nand U26544 (N_26544,N_26487,N_26342);
nor U26545 (N_26545,N_26375,N_26347);
xor U26546 (N_26546,N_26491,N_26403);
nor U26547 (N_26547,N_26467,N_26259);
or U26548 (N_26548,N_26411,N_26421);
nor U26549 (N_26549,N_26325,N_26270);
or U26550 (N_26550,N_26466,N_26321);
or U26551 (N_26551,N_26336,N_26436);
nor U26552 (N_26552,N_26287,N_26456);
nor U26553 (N_26553,N_26316,N_26377);
or U26554 (N_26554,N_26251,N_26359);
nor U26555 (N_26555,N_26369,N_26458);
or U26556 (N_26556,N_26276,N_26368);
xor U26557 (N_26557,N_26387,N_26305);
and U26558 (N_26558,N_26438,N_26307);
or U26559 (N_26559,N_26455,N_26292);
and U26560 (N_26560,N_26425,N_26329);
nor U26561 (N_26561,N_26290,N_26468);
nor U26562 (N_26562,N_26335,N_26299);
xnor U26563 (N_26563,N_26490,N_26365);
nor U26564 (N_26564,N_26294,N_26396);
nand U26565 (N_26565,N_26390,N_26317);
or U26566 (N_26566,N_26465,N_26477);
or U26567 (N_26567,N_26252,N_26485);
nand U26568 (N_26568,N_26303,N_26313);
or U26569 (N_26569,N_26353,N_26253);
xor U26570 (N_26570,N_26263,N_26302);
or U26571 (N_26571,N_26416,N_26312);
xor U26572 (N_26572,N_26417,N_26482);
nor U26573 (N_26573,N_26254,N_26489);
nor U26574 (N_26574,N_26289,N_26388);
nand U26575 (N_26575,N_26346,N_26437);
and U26576 (N_26576,N_26337,N_26326);
or U26577 (N_26577,N_26439,N_26373);
xnor U26578 (N_26578,N_26372,N_26265);
xor U26579 (N_26579,N_26404,N_26306);
nand U26580 (N_26580,N_26351,N_26257);
and U26581 (N_26581,N_26370,N_26277);
and U26582 (N_26582,N_26459,N_26415);
xor U26583 (N_26583,N_26327,N_26405);
nor U26584 (N_26584,N_26457,N_26268);
or U26585 (N_26585,N_26429,N_26453);
and U26586 (N_26586,N_26492,N_26408);
nand U26587 (N_26587,N_26279,N_26352);
nor U26588 (N_26588,N_26428,N_26484);
xnor U26589 (N_26589,N_26413,N_26441);
or U26590 (N_26590,N_26494,N_26400);
nor U26591 (N_26591,N_26309,N_26393);
and U26592 (N_26592,N_26498,N_26475);
xor U26593 (N_26593,N_26432,N_26434);
or U26594 (N_26594,N_26450,N_26463);
and U26595 (N_26595,N_26314,N_26348);
nor U26596 (N_26596,N_26384,N_26472);
nor U26597 (N_26597,N_26499,N_26339);
or U26598 (N_26598,N_26461,N_26288);
nor U26599 (N_26599,N_26363,N_26495);
nand U26600 (N_26600,N_26443,N_26424);
and U26601 (N_26601,N_26361,N_26338);
xor U26602 (N_26602,N_26469,N_26397);
or U26603 (N_26603,N_26269,N_26334);
xnor U26604 (N_26604,N_26296,N_26394);
nand U26605 (N_26605,N_26322,N_26260);
nand U26606 (N_26606,N_26376,N_26274);
nand U26607 (N_26607,N_26293,N_26442);
nand U26608 (N_26608,N_26360,N_26354);
and U26609 (N_26609,N_26300,N_26349);
nand U26610 (N_26610,N_26452,N_26285);
nand U26611 (N_26611,N_26311,N_26395);
xor U26612 (N_26612,N_26304,N_26340);
or U26613 (N_26613,N_26407,N_26371);
or U26614 (N_26614,N_26486,N_26479);
or U26615 (N_26615,N_26412,N_26406);
nor U26616 (N_26616,N_26267,N_26310);
or U26617 (N_26617,N_26422,N_26328);
and U26618 (N_26618,N_26271,N_26281);
xnor U26619 (N_26619,N_26324,N_26273);
or U26620 (N_26620,N_26284,N_26367);
nand U26621 (N_26621,N_26301,N_26250);
xor U26622 (N_26622,N_26278,N_26286);
xnor U26623 (N_26623,N_26445,N_26358);
and U26624 (N_26624,N_26298,N_26464);
or U26625 (N_26625,N_26394,N_26315);
nand U26626 (N_26626,N_26441,N_26257);
nor U26627 (N_26627,N_26338,N_26496);
nand U26628 (N_26628,N_26417,N_26498);
xor U26629 (N_26629,N_26258,N_26435);
and U26630 (N_26630,N_26492,N_26304);
nor U26631 (N_26631,N_26429,N_26439);
xnor U26632 (N_26632,N_26291,N_26358);
nand U26633 (N_26633,N_26284,N_26494);
xor U26634 (N_26634,N_26254,N_26337);
and U26635 (N_26635,N_26329,N_26338);
or U26636 (N_26636,N_26289,N_26354);
nor U26637 (N_26637,N_26444,N_26382);
and U26638 (N_26638,N_26367,N_26446);
xor U26639 (N_26639,N_26335,N_26309);
nor U26640 (N_26640,N_26367,N_26314);
nand U26641 (N_26641,N_26366,N_26494);
xor U26642 (N_26642,N_26403,N_26348);
and U26643 (N_26643,N_26353,N_26286);
nor U26644 (N_26644,N_26482,N_26302);
xor U26645 (N_26645,N_26281,N_26288);
xor U26646 (N_26646,N_26495,N_26357);
nor U26647 (N_26647,N_26429,N_26434);
or U26648 (N_26648,N_26280,N_26345);
or U26649 (N_26649,N_26367,N_26363);
nor U26650 (N_26650,N_26444,N_26278);
nor U26651 (N_26651,N_26311,N_26289);
xor U26652 (N_26652,N_26437,N_26460);
and U26653 (N_26653,N_26453,N_26394);
xnor U26654 (N_26654,N_26351,N_26435);
or U26655 (N_26655,N_26414,N_26404);
and U26656 (N_26656,N_26416,N_26340);
and U26657 (N_26657,N_26451,N_26392);
xor U26658 (N_26658,N_26283,N_26470);
xnor U26659 (N_26659,N_26355,N_26308);
xor U26660 (N_26660,N_26470,N_26478);
and U26661 (N_26661,N_26313,N_26402);
or U26662 (N_26662,N_26465,N_26342);
nand U26663 (N_26663,N_26473,N_26376);
xnor U26664 (N_26664,N_26289,N_26446);
or U26665 (N_26665,N_26374,N_26261);
and U26666 (N_26666,N_26317,N_26340);
xnor U26667 (N_26667,N_26261,N_26288);
or U26668 (N_26668,N_26485,N_26415);
xnor U26669 (N_26669,N_26396,N_26351);
nor U26670 (N_26670,N_26396,N_26483);
xnor U26671 (N_26671,N_26458,N_26477);
nand U26672 (N_26672,N_26356,N_26366);
or U26673 (N_26673,N_26382,N_26397);
nor U26674 (N_26674,N_26440,N_26303);
nor U26675 (N_26675,N_26444,N_26460);
xor U26676 (N_26676,N_26293,N_26408);
xnor U26677 (N_26677,N_26432,N_26356);
and U26678 (N_26678,N_26484,N_26315);
xnor U26679 (N_26679,N_26473,N_26461);
nand U26680 (N_26680,N_26349,N_26429);
and U26681 (N_26681,N_26308,N_26329);
and U26682 (N_26682,N_26494,N_26402);
and U26683 (N_26683,N_26410,N_26454);
or U26684 (N_26684,N_26361,N_26325);
nor U26685 (N_26685,N_26467,N_26438);
and U26686 (N_26686,N_26299,N_26309);
or U26687 (N_26687,N_26375,N_26315);
or U26688 (N_26688,N_26423,N_26455);
or U26689 (N_26689,N_26468,N_26264);
or U26690 (N_26690,N_26436,N_26347);
nand U26691 (N_26691,N_26282,N_26465);
or U26692 (N_26692,N_26439,N_26378);
and U26693 (N_26693,N_26471,N_26322);
and U26694 (N_26694,N_26448,N_26367);
nand U26695 (N_26695,N_26380,N_26377);
nand U26696 (N_26696,N_26478,N_26340);
xnor U26697 (N_26697,N_26477,N_26286);
xnor U26698 (N_26698,N_26251,N_26354);
or U26699 (N_26699,N_26391,N_26306);
nand U26700 (N_26700,N_26443,N_26265);
nand U26701 (N_26701,N_26445,N_26338);
and U26702 (N_26702,N_26258,N_26259);
or U26703 (N_26703,N_26318,N_26253);
and U26704 (N_26704,N_26304,N_26450);
nand U26705 (N_26705,N_26432,N_26481);
xnor U26706 (N_26706,N_26446,N_26464);
nor U26707 (N_26707,N_26263,N_26425);
nand U26708 (N_26708,N_26334,N_26473);
xnor U26709 (N_26709,N_26337,N_26276);
nor U26710 (N_26710,N_26314,N_26330);
and U26711 (N_26711,N_26391,N_26467);
and U26712 (N_26712,N_26280,N_26315);
nor U26713 (N_26713,N_26354,N_26323);
and U26714 (N_26714,N_26344,N_26434);
nor U26715 (N_26715,N_26319,N_26353);
and U26716 (N_26716,N_26432,N_26467);
or U26717 (N_26717,N_26470,N_26466);
nor U26718 (N_26718,N_26436,N_26402);
nor U26719 (N_26719,N_26288,N_26302);
nor U26720 (N_26720,N_26309,N_26307);
and U26721 (N_26721,N_26384,N_26386);
and U26722 (N_26722,N_26349,N_26250);
and U26723 (N_26723,N_26436,N_26290);
and U26724 (N_26724,N_26431,N_26251);
xor U26725 (N_26725,N_26418,N_26365);
nor U26726 (N_26726,N_26367,N_26424);
or U26727 (N_26727,N_26361,N_26481);
or U26728 (N_26728,N_26489,N_26378);
and U26729 (N_26729,N_26337,N_26478);
and U26730 (N_26730,N_26257,N_26379);
nor U26731 (N_26731,N_26282,N_26407);
and U26732 (N_26732,N_26381,N_26438);
or U26733 (N_26733,N_26484,N_26328);
or U26734 (N_26734,N_26288,N_26385);
xnor U26735 (N_26735,N_26477,N_26490);
or U26736 (N_26736,N_26378,N_26318);
xor U26737 (N_26737,N_26337,N_26413);
nand U26738 (N_26738,N_26305,N_26306);
and U26739 (N_26739,N_26299,N_26377);
nand U26740 (N_26740,N_26257,N_26488);
xnor U26741 (N_26741,N_26460,N_26300);
nor U26742 (N_26742,N_26431,N_26444);
xnor U26743 (N_26743,N_26469,N_26301);
and U26744 (N_26744,N_26320,N_26379);
or U26745 (N_26745,N_26325,N_26385);
nor U26746 (N_26746,N_26266,N_26264);
and U26747 (N_26747,N_26383,N_26436);
and U26748 (N_26748,N_26439,N_26294);
and U26749 (N_26749,N_26288,N_26482);
xnor U26750 (N_26750,N_26521,N_26716);
nand U26751 (N_26751,N_26594,N_26573);
nand U26752 (N_26752,N_26605,N_26583);
nor U26753 (N_26753,N_26625,N_26679);
and U26754 (N_26754,N_26582,N_26658);
xor U26755 (N_26755,N_26733,N_26590);
nor U26756 (N_26756,N_26647,N_26681);
nand U26757 (N_26757,N_26559,N_26713);
nand U26758 (N_26758,N_26690,N_26640);
and U26759 (N_26759,N_26629,N_26689);
xor U26760 (N_26760,N_26637,N_26552);
nand U26761 (N_26761,N_26504,N_26705);
nor U26762 (N_26762,N_26725,N_26718);
or U26763 (N_26763,N_26668,N_26683);
and U26764 (N_26764,N_26588,N_26530);
or U26765 (N_26765,N_26643,N_26694);
or U26766 (N_26766,N_26632,N_26736);
xor U26767 (N_26767,N_26674,N_26641);
nand U26768 (N_26768,N_26607,N_26574);
nor U26769 (N_26769,N_26724,N_26548);
or U26770 (N_26770,N_26517,N_26747);
nor U26771 (N_26771,N_26741,N_26506);
nand U26772 (N_26772,N_26734,N_26737);
nor U26773 (N_26773,N_26650,N_26648);
xor U26774 (N_26774,N_26610,N_26619);
and U26775 (N_26775,N_26666,N_26722);
xnor U26776 (N_26776,N_26631,N_26720);
nor U26777 (N_26777,N_26685,N_26654);
and U26778 (N_26778,N_26719,N_26622);
or U26779 (N_26779,N_26721,N_26682);
or U26780 (N_26780,N_26592,N_26744);
or U26781 (N_26781,N_26554,N_26555);
and U26782 (N_26782,N_26696,N_26701);
nand U26783 (N_26783,N_26717,N_26616);
and U26784 (N_26784,N_26510,N_26728);
nand U26785 (N_26785,N_26630,N_26730);
xnor U26786 (N_26786,N_26620,N_26512);
or U26787 (N_26787,N_26529,N_26662);
and U26788 (N_26788,N_26556,N_26646);
and U26789 (N_26789,N_26535,N_26618);
and U26790 (N_26790,N_26591,N_26599);
xnor U26791 (N_26791,N_26514,N_26739);
or U26792 (N_26792,N_26714,N_26693);
and U26793 (N_26793,N_26667,N_26533);
nor U26794 (N_26794,N_26553,N_26505);
nand U26795 (N_26795,N_26670,N_26612);
xnor U26796 (N_26796,N_26746,N_26561);
and U26797 (N_26797,N_26522,N_26707);
and U26798 (N_26798,N_26710,N_26664);
nand U26799 (N_26799,N_26597,N_26604);
or U26800 (N_26800,N_26563,N_26738);
or U26801 (N_26801,N_26581,N_26532);
and U26802 (N_26802,N_26603,N_26577);
nand U26803 (N_26803,N_26623,N_26525);
or U26804 (N_26804,N_26572,N_26723);
nor U26805 (N_26805,N_26665,N_26671);
nand U26806 (N_26806,N_26749,N_26500);
nand U26807 (N_26807,N_26642,N_26542);
xor U26808 (N_26808,N_26684,N_26543);
and U26809 (N_26809,N_26614,N_26566);
and U26810 (N_26810,N_26729,N_26508);
nor U26811 (N_26811,N_26613,N_26633);
nand U26812 (N_26812,N_26695,N_26732);
and U26813 (N_26813,N_26691,N_26540);
nor U26814 (N_26814,N_26606,N_26698);
nand U26815 (N_26815,N_26546,N_26518);
or U26816 (N_26816,N_26537,N_26692);
xor U26817 (N_26817,N_26507,N_26528);
xnor U26818 (N_26818,N_26519,N_26651);
nor U26819 (N_26819,N_26520,N_26557);
nand U26820 (N_26820,N_26609,N_26558);
xor U26821 (N_26821,N_26731,N_26653);
nand U26822 (N_26822,N_26541,N_26656);
nor U26823 (N_26823,N_26536,N_26501);
xor U26824 (N_26824,N_26748,N_26702);
xor U26825 (N_26825,N_26727,N_26601);
xnor U26826 (N_26826,N_26587,N_26627);
and U26827 (N_26827,N_26657,N_26675);
and U26828 (N_26828,N_26634,N_26688);
nor U26829 (N_26829,N_26678,N_26743);
nor U26830 (N_26830,N_26663,N_26661);
or U26831 (N_26831,N_26595,N_26711);
nor U26832 (N_26832,N_26598,N_26515);
and U26833 (N_26833,N_26513,N_26545);
nand U26834 (N_26834,N_26579,N_26596);
or U26835 (N_26835,N_26709,N_26672);
or U26836 (N_26836,N_26669,N_26742);
or U26837 (N_26837,N_26602,N_26569);
xor U26838 (N_26838,N_26699,N_26740);
nor U26839 (N_26839,N_26659,N_26502);
and U26840 (N_26840,N_26551,N_26547);
nand U26841 (N_26841,N_26509,N_26715);
and U26842 (N_26842,N_26735,N_26611);
and U26843 (N_26843,N_26655,N_26534);
nand U26844 (N_26844,N_26538,N_26575);
xor U26845 (N_26845,N_26503,N_26704);
and U26846 (N_26846,N_26628,N_26639);
or U26847 (N_26847,N_26624,N_26652);
nor U26848 (N_26848,N_26539,N_26589);
or U26849 (N_26849,N_26660,N_26712);
or U26850 (N_26850,N_26527,N_26580);
nand U26851 (N_26851,N_26524,N_26549);
nand U26852 (N_26852,N_26544,N_26578);
or U26853 (N_26853,N_26531,N_26697);
and U26854 (N_26854,N_26560,N_26644);
xnor U26855 (N_26855,N_26645,N_26550);
xnor U26856 (N_26856,N_26565,N_26617);
or U26857 (N_26857,N_26673,N_26621);
and U26858 (N_26858,N_26680,N_26568);
nand U26859 (N_26859,N_26706,N_26608);
nand U26860 (N_26860,N_26726,N_26570);
or U26861 (N_26861,N_26636,N_26562);
nand U26862 (N_26862,N_26576,N_26567);
and U26863 (N_26863,N_26511,N_26626);
or U26864 (N_26864,N_26677,N_26615);
nand U26865 (N_26865,N_26516,N_26593);
and U26866 (N_26866,N_26676,N_26686);
and U26867 (N_26867,N_26638,N_26687);
nand U26868 (N_26868,N_26523,N_26526);
nand U26869 (N_26869,N_26708,N_26700);
or U26870 (N_26870,N_26600,N_26584);
or U26871 (N_26871,N_26635,N_26564);
nand U26872 (N_26872,N_26745,N_26649);
nor U26873 (N_26873,N_26586,N_26571);
or U26874 (N_26874,N_26703,N_26585);
xnor U26875 (N_26875,N_26523,N_26641);
nor U26876 (N_26876,N_26725,N_26716);
and U26877 (N_26877,N_26612,N_26547);
nor U26878 (N_26878,N_26581,N_26662);
nand U26879 (N_26879,N_26576,N_26575);
and U26880 (N_26880,N_26517,N_26645);
nor U26881 (N_26881,N_26707,N_26702);
nand U26882 (N_26882,N_26619,N_26570);
and U26883 (N_26883,N_26562,N_26724);
or U26884 (N_26884,N_26658,N_26666);
nor U26885 (N_26885,N_26638,N_26731);
and U26886 (N_26886,N_26608,N_26533);
or U26887 (N_26887,N_26516,N_26548);
or U26888 (N_26888,N_26682,N_26563);
nand U26889 (N_26889,N_26541,N_26739);
and U26890 (N_26890,N_26518,N_26604);
xor U26891 (N_26891,N_26646,N_26730);
and U26892 (N_26892,N_26601,N_26703);
nor U26893 (N_26893,N_26711,N_26503);
nor U26894 (N_26894,N_26570,N_26560);
and U26895 (N_26895,N_26640,N_26607);
nand U26896 (N_26896,N_26542,N_26523);
nand U26897 (N_26897,N_26608,N_26503);
xor U26898 (N_26898,N_26693,N_26595);
and U26899 (N_26899,N_26528,N_26669);
and U26900 (N_26900,N_26541,N_26702);
xnor U26901 (N_26901,N_26709,N_26680);
nand U26902 (N_26902,N_26721,N_26556);
nand U26903 (N_26903,N_26606,N_26584);
or U26904 (N_26904,N_26598,N_26540);
nor U26905 (N_26905,N_26513,N_26587);
nor U26906 (N_26906,N_26728,N_26627);
and U26907 (N_26907,N_26528,N_26749);
xor U26908 (N_26908,N_26694,N_26677);
nor U26909 (N_26909,N_26575,N_26652);
nand U26910 (N_26910,N_26705,N_26599);
nand U26911 (N_26911,N_26721,N_26731);
or U26912 (N_26912,N_26710,N_26600);
or U26913 (N_26913,N_26554,N_26708);
nand U26914 (N_26914,N_26690,N_26615);
or U26915 (N_26915,N_26740,N_26747);
or U26916 (N_26916,N_26563,N_26559);
nand U26917 (N_26917,N_26573,N_26581);
xor U26918 (N_26918,N_26528,N_26523);
xnor U26919 (N_26919,N_26589,N_26609);
nand U26920 (N_26920,N_26687,N_26505);
xnor U26921 (N_26921,N_26532,N_26589);
and U26922 (N_26922,N_26682,N_26747);
and U26923 (N_26923,N_26658,N_26553);
nand U26924 (N_26924,N_26645,N_26745);
or U26925 (N_26925,N_26611,N_26637);
nand U26926 (N_26926,N_26593,N_26733);
xnor U26927 (N_26927,N_26683,N_26580);
and U26928 (N_26928,N_26622,N_26669);
and U26929 (N_26929,N_26560,N_26608);
xor U26930 (N_26930,N_26583,N_26639);
nand U26931 (N_26931,N_26505,N_26668);
or U26932 (N_26932,N_26658,N_26520);
nor U26933 (N_26933,N_26717,N_26534);
nand U26934 (N_26934,N_26615,N_26612);
nor U26935 (N_26935,N_26532,N_26735);
or U26936 (N_26936,N_26688,N_26500);
nand U26937 (N_26937,N_26689,N_26550);
and U26938 (N_26938,N_26626,N_26607);
nor U26939 (N_26939,N_26657,N_26694);
and U26940 (N_26940,N_26583,N_26662);
and U26941 (N_26941,N_26650,N_26550);
nand U26942 (N_26942,N_26666,N_26555);
or U26943 (N_26943,N_26621,N_26558);
and U26944 (N_26944,N_26542,N_26736);
or U26945 (N_26945,N_26651,N_26644);
and U26946 (N_26946,N_26606,N_26738);
nor U26947 (N_26947,N_26502,N_26507);
or U26948 (N_26948,N_26533,N_26732);
nor U26949 (N_26949,N_26685,N_26620);
and U26950 (N_26950,N_26531,N_26631);
nor U26951 (N_26951,N_26660,N_26642);
nand U26952 (N_26952,N_26723,N_26713);
or U26953 (N_26953,N_26590,N_26731);
and U26954 (N_26954,N_26535,N_26680);
nor U26955 (N_26955,N_26727,N_26504);
xor U26956 (N_26956,N_26585,N_26601);
nand U26957 (N_26957,N_26700,N_26549);
nand U26958 (N_26958,N_26707,N_26587);
xor U26959 (N_26959,N_26703,N_26501);
or U26960 (N_26960,N_26580,N_26632);
nand U26961 (N_26961,N_26705,N_26510);
nor U26962 (N_26962,N_26665,N_26609);
and U26963 (N_26963,N_26720,N_26665);
or U26964 (N_26964,N_26602,N_26599);
xnor U26965 (N_26965,N_26634,N_26629);
nor U26966 (N_26966,N_26640,N_26728);
nor U26967 (N_26967,N_26689,N_26735);
or U26968 (N_26968,N_26535,N_26575);
nand U26969 (N_26969,N_26564,N_26681);
or U26970 (N_26970,N_26614,N_26724);
nor U26971 (N_26971,N_26586,N_26565);
or U26972 (N_26972,N_26713,N_26546);
and U26973 (N_26973,N_26647,N_26695);
nand U26974 (N_26974,N_26504,N_26543);
nand U26975 (N_26975,N_26538,N_26643);
or U26976 (N_26976,N_26666,N_26588);
and U26977 (N_26977,N_26599,N_26513);
nand U26978 (N_26978,N_26717,N_26628);
xor U26979 (N_26979,N_26679,N_26670);
nand U26980 (N_26980,N_26581,N_26519);
xnor U26981 (N_26981,N_26504,N_26582);
nor U26982 (N_26982,N_26699,N_26673);
and U26983 (N_26983,N_26736,N_26714);
nand U26984 (N_26984,N_26674,N_26651);
xnor U26985 (N_26985,N_26623,N_26683);
nand U26986 (N_26986,N_26666,N_26650);
nor U26987 (N_26987,N_26589,N_26624);
nand U26988 (N_26988,N_26709,N_26742);
and U26989 (N_26989,N_26709,N_26718);
and U26990 (N_26990,N_26623,N_26622);
nor U26991 (N_26991,N_26641,N_26586);
nand U26992 (N_26992,N_26553,N_26511);
nor U26993 (N_26993,N_26673,N_26552);
nand U26994 (N_26994,N_26695,N_26712);
and U26995 (N_26995,N_26692,N_26656);
nor U26996 (N_26996,N_26618,N_26667);
nor U26997 (N_26997,N_26680,N_26504);
nor U26998 (N_26998,N_26659,N_26719);
or U26999 (N_26999,N_26687,N_26506);
and U27000 (N_27000,N_26843,N_26777);
nand U27001 (N_27001,N_26992,N_26836);
nor U27002 (N_27002,N_26819,N_26960);
xnor U27003 (N_27003,N_26753,N_26780);
or U27004 (N_27004,N_26834,N_26799);
nand U27005 (N_27005,N_26824,N_26872);
nand U27006 (N_27006,N_26976,N_26791);
or U27007 (N_27007,N_26883,N_26981);
xor U27008 (N_27008,N_26811,N_26830);
and U27009 (N_27009,N_26877,N_26949);
and U27010 (N_27010,N_26876,N_26886);
nor U27011 (N_27011,N_26764,N_26855);
nand U27012 (N_27012,N_26888,N_26947);
or U27013 (N_27013,N_26793,N_26972);
nor U27014 (N_27014,N_26999,N_26952);
or U27015 (N_27015,N_26977,N_26930);
nand U27016 (N_27016,N_26990,N_26916);
and U27017 (N_27017,N_26773,N_26871);
nor U27018 (N_27018,N_26827,N_26920);
xor U27019 (N_27019,N_26912,N_26779);
and U27020 (N_27020,N_26806,N_26860);
nand U27021 (N_27021,N_26818,N_26863);
and U27022 (N_27022,N_26924,N_26852);
or U27023 (N_27023,N_26911,N_26885);
xnor U27024 (N_27024,N_26787,N_26758);
nor U27025 (N_27025,N_26807,N_26932);
xnor U27026 (N_27026,N_26896,N_26866);
nor U27027 (N_27027,N_26998,N_26835);
nor U27028 (N_27028,N_26781,N_26897);
xnor U27029 (N_27029,N_26881,N_26765);
and U27030 (N_27030,N_26805,N_26769);
nor U27031 (N_27031,N_26803,N_26870);
or U27032 (N_27032,N_26917,N_26776);
nand U27033 (N_27033,N_26857,N_26783);
and U27034 (N_27034,N_26821,N_26891);
nor U27035 (N_27035,N_26950,N_26809);
or U27036 (N_27036,N_26802,N_26941);
or U27037 (N_27037,N_26768,N_26894);
or U27038 (N_27038,N_26808,N_26944);
xnor U27039 (N_27039,N_26804,N_26928);
nand U27040 (N_27040,N_26859,N_26760);
nor U27041 (N_27041,N_26794,N_26974);
nor U27042 (N_27042,N_26962,N_26767);
and U27043 (N_27043,N_26850,N_26994);
and U27044 (N_27044,N_26782,N_26832);
nand U27045 (N_27045,N_26795,N_26820);
nor U27046 (N_27046,N_26889,N_26757);
nand U27047 (N_27047,N_26923,N_26786);
nand U27048 (N_27048,N_26961,N_26948);
nand U27049 (N_27049,N_26801,N_26945);
nand U27050 (N_27050,N_26858,N_26996);
nand U27051 (N_27051,N_26997,N_26775);
nand U27052 (N_27052,N_26926,N_26831);
nor U27053 (N_27053,N_26893,N_26868);
and U27054 (N_27054,N_26839,N_26865);
nand U27055 (N_27055,N_26861,N_26762);
or U27056 (N_27056,N_26914,N_26937);
and U27057 (N_27057,N_26841,N_26823);
xnor U27058 (N_27058,N_26970,N_26918);
nand U27059 (N_27059,N_26789,N_26822);
and U27060 (N_27060,N_26958,N_26954);
xor U27061 (N_27061,N_26902,N_26921);
xnor U27062 (N_27062,N_26939,N_26880);
nor U27063 (N_27063,N_26750,N_26908);
nor U27064 (N_27064,N_26873,N_26965);
nor U27065 (N_27065,N_26752,N_26982);
and U27066 (N_27066,N_26854,N_26826);
or U27067 (N_27067,N_26771,N_26979);
nand U27068 (N_27068,N_26864,N_26878);
and U27069 (N_27069,N_26959,N_26851);
or U27070 (N_27070,N_26985,N_26910);
nand U27071 (N_27071,N_26975,N_26967);
nor U27072 (N_27072,N_26848,N_26840);
or U27073 (N_27073,N_26798,N_26838);
nor U27074 (N_27074,N_26963,N_26813);
nand U27075 (N_27075,N_26906,N_26966);
nor U27076 (N_27076,N_26988,N_26774);
xor U27077 (N_27077,N_26943,N_26971);
nand U27078 (N_27078,N_26935,N_26882);
or U27079 (N_27079,N_26956,N_26862);
nor U27080 (N_27080,N_26833,N_26927);
xor U27081 (N_27081,N_26812,N_26788);
or U27082 (N_27082,N_26761,N_26915);
and U27083 (N_27083,N_26968,N_26991);
nor U27084 (N_27084,N_26770,N_26973);
nand U27085 (N_27085,N_26987,N_26796);
and U27086 (N_27086,N_26931,N_26800);
or U27087 (N_27087,N_26817,N_26810);
nor U27088 (N_27088,N_26828,N_26995);
nand U27089 (N_27089,N_26792,N_26898);
nor U27090 (N_27090,N_26867,N_26933);
xor U27091 (N_27091,N_26955,N_26900);
or U27092 (N_27092,N_26847,N_26778);
and U27093 (N_27093,N_26907,N_26909);
nand U27094 (N_27094,N_26755,N_26797);
nand U27095 (N_27095,N_26856,N_26892);
xor U27096 (N_27096,N_26829,N_26989);
nor U27097 (N_27097,N_26751,N_26986);
and U27098 (N_27098,N_26969,N_26845);
xnor U27099 (N_27099,N_26853,N_26938);
nand U27100 (N_27100,N_26895,N_26919);
nand U27101 (N_27101,N_26887,N_26837);
nor U27102 (N_27102,N_26846,N_26904);
and U27103 (N_27103,N_26874,N_26925);
nand U27104 (N_27104,N_26814,N_26825);
xor U27105 (N_27105,N_26763,N_26844);
and U27106 (N_27106,N_26754,N_26784);
nand U27107 (N_27107,N_26980,N_26929);
and U27108 (N_27108,N_26934,N_26884);
xor U27109 (N_27109,N_26905,N_26913);
or U27110 (N_27110,N_26766,N_26946);
and U27111 (N_27111,N_26869,N_26993);
or U27112 (N_27112,N_26951,N_26983);
nand U27113 (N_27113,N_26759,N_26901);
xor U27114 (N_27114,N_26756,N_26953);
xor U27115 (N_27115,N_26984,N_26815);
and U27116 (N_27116,N_26957,N_26940);
and U27117 (N_27117,N_26899,N_26875);
and U27118 (N_27118,N_26964,N_26842);
and U27119 (N_27119,N_26890,N_26978);
nand U27120 (N_27120,N_26790,N_26942);
nor U27121 (N_27121,N_26785,N_26936);
xor U27122 (N_27122,N_26903,N_26772);
nand U27123 (N_27123,N_26849,N_26816);
or U27124 (N_27124,N_26922,N_26879);
xnor U27125 (N_27125,N_26910,N_26907);
or U27126 (N_27126,N_26841,N_26883);
xor U27127 (N_27127,N_26886,N_26833);
and U27128 (N_27128,N_26862,N_26899);
xnor U27129 (N_27129,N_26880,N_26957);
or U27130 (N_27130,N_26876,N_26951);
xor U27131 (N_27131,N_26771,N_26827);
nand U27132 (N_27132,N_26851,N_26777);
xnor U27133 (N_27133,N_26891,N_26767);
and U27134 (N_27134,N_26759,N_26865);
and U27135 (N_27135,N_26979,N_26952);
xor U27136 (N_27136,N_26820,N_26823);
xor U27137 (N_27137,N_26853,N_26955);
and U27138 (N_27138,N_26768,N_26956);
nand U27139 (N_27139,N_26932,N_26827);
nor U27140 (N_27140,N_26754,N_26895);
nand U27141 (N_27141,N_26944,N_26885);
or U27142 (N_27142,N_26819,N_26982);
nor U27143 (N_27143,N_26944,N_26978);
nor U27144 (N_27144,N_26836,N_26910);
or U27145 (N_27145,N_26890,N_26833);
nand U27146 (N_27146,N_26915,N_26840);
or U27147 (N_27147,N_26766,N_26901);
and U27148 (N_27148,N_26908,N_26876);
and U27149 (N_27149,N_26988,N_26902);
nor U27150 (N_27150,N_26909,N_26953);
nor U27151 (N_27151,N_26983,N_26898);
nor U27152 (N_27152,N_26810,N_26818);
and U27153 (N_27153,N_26935,N_26948);
or U27154 (N_27154,N_26920,N_26982);
nor U27155 (N_27155,N_26936,N_26812);
and U27156 (N_27156,N_26886,N_26998);
nand U27157 (N_27157,N_26937,N_26843);
and U27158 (N_27158,N_26906,N_26947);
nor U27159 (N_27159,N_26961,N_26978);
nor U27160 (N_27160,N_26758,N_26859);
and U27161 (N_27161,N_26853,N_26789);
nand U27162 (N_27162,N_26994,N_26918);
or U27163 (N_27163,N_26862,N_26967);
and U27164 (N_27164,N_26947,N_26875);
nor U27165 (N_27165,N_26789,N_26957);
nand U27166 (N_27166,N_26872,N_26951);
or U27167 (N_27167,N_26971,N_26908);
xnor U27168 (N_27168,N_26847,N_26935);
or U27169 (N_27169,N_26930,N_26799);
nor U27170 (N_27170,N_26803,N_26919);
nor U27171 (N_27171,N_26999,N_26881);
and U27172 (N_27172,N_26949,N_26977);
and U27173 (N_27173,N_26835,N_26983);
and U27174 (N_27174,N_26810,N_26925);
nor U27175 (N_27175,N_26751,N_26778);
xor U27176 (N_27176,N_26835,N_26878);
nand U27177 (N_27177,N_26801,N_26763);
xnor U27178 (N_27178,N_26963,N_26774);
nand U27179 (N_27179,N_26784,N_26805);
xnor U27180 (N_27180,N_26809,N_26804);
nand U27181 (N_27181,N_26786,N_26925);
or U27182 (N_27182,N_26891,N_26887);
xnor U27183 (N_27183,N_26754,N_26973);
and U27184 (N_27184,N_26935,N_26776);
or U27185 (N_27185,N_26753,N_26972);
nand U27186 (N_27186,N_26951,N_26948);
nand U27187 (N_27187,N_26938,N_26757);
xor U27188 (N_27188,N_26882,N_26796);
and U27189 (N_27189,N_26767,N_26853);
nor U27190 (N_27190,N_26798,N_26959);
or U27191 (N_27191,N_26977,N_26797);
and U27192 (N_27192,N_26824,N_26992);
or U27193 (N_27193,N_26970,N_26932);
nor U27194 (N_27194,N_26939,N_26835);
xor U27195 (N_27195,N_26880,N_26998);
nor U27196 (N_27196,N_26886,N_26961);
xnor U27197 (N_27197,N_26861,N_26821);
nand U27198 (N_27198,N_26878,N_26828);
nor U27199 (N_27199,N_26778,N_26823);
nor U27200 (N_27200,N_26766,N_26926);
and U27201 (N_27201,N_26810,N_26802);
nor U27202 (N_27202,N_26821,N_26754);
nor U27203 (N_27203,N_26922,N_26887);
nand U27204 (N_27204,N_26943,N_26990);
nor U27205 (N_27205,N_26848,N_26967);
or U27206 (N_27206,N_26846,N_26984);
or U27207 (N_27207,N_26775,N_26758);
xor U27208 (N_27208,N_26755,N_26953);
or U27209 (N_27209,N_26955,N_26790);
xor U27210 (N_27210,N_26904,N_26985);
nand U27211 (N_27211,N_26778,N_26866);
and U27212 (N_27212,N_26955,N_26934);
xnor U27213 (N_27213,N_26756,N_26981);
xnor U27214 (N_27214,N_26896,N_26755);
nor U27215 (N_27215,N_26919,N_26819);
nor U27216 (N_27216,N_26968,N_26939);
xnor U27217 (N_27217,N_26959,N_26807);
nand U27218 (N_27218,N_26802,N_26951);
nor U27219 (N_27219,N_26779,N_26777);
nor U27220 (N_27220,N_26959,N_26871);
nor U27221 (N_27221,N_26936,N_26860);
and U27222 (N_27222,N_26918,N_26986);
or U27223 (N_27223,N_26976,N_26990);
nand U27224 (N_27224,N_26933,N_26860);
nor U27225 (N_27225,N_26775,N_26869);
nand U27226 (N_27226,N_26936,N_26813);
and U27227 (N_27227,N_26899,N_26868);
nor U27228 (N_27228,N_26793,N_26771);
nand U27229 (N_27229,N_26932,N_26985);
xor U27230 (N_27230,N_26760,N_26872);
xor U27231 (N_27231,N_26818,N_26958);
nor U27232 (N_27232,N_26974,N_26835);
or U27233 (N_27233,N_26835,N_26850);
nor U27234 (N_27234,N_26845,N_26881);
nand U27235 (N_27235,N_26964,N_26845);
or U27236 (N_27236,N_26841,N_26875);
xnor U27237 (N_27237,N_26816,N_26853);
xor U27238 (N_27238,N_26750,N_26955);
or U27239 (N_27239,N_26977,N_26896);
and U27240 (N_27240,N_26913,N_26967);
xor U27241 (N_27241,N_26771,N_26879);
nand U27242 (N_27242,N_26876,N_26762);
and U27243 (N_27243,N_26787,N_26796);
or U27244 (N_27244,N_26954,N_26755);
nor U27245 (N_27245,N_26998,N_26891);
nand U27246 (N_27246,N_26997,N_26899);
nor U27247 (N_27247,N_26765,N_26853);
xor U27248 (N_27248,N_26881,N_26823);
or U27249 (N_27249,N_26807,N_26850);
nand U27250 (N_27250,N_27023,N_27014);
and U27251 (N_27251,N_27036,N_27146);
nor U27252 (N_27252,N_27041,N_27069);
and U27253 (N_27253,N_27020,N_27142);
nand U27254 (N_27254,N_27159,N_27178);
xor U27255 (N_27255,N_27131,N_27109);
nor U27256 (N_27256,N_27003,N_27090);
nand U27257 (N_27257,N_27065,N_27057);
nand U27258 (N_27258,N_27165,N_27234);
xnor U27259 (N_27259,N_27096,N_27229);
nand U27260 (N_27260,N_27058,N_27009);
nor U27261 (N_27261,N_27201,N_27237);
and U27262 (N_27262,N_27227,N_27174);
or U27263 (N_27263,N_27054,N_27028);
xnor U27264 (N_27264,N_27018,N_27015);
and U27265 (N_27265,N_27120,N_27195);
nand U27266 (N_27266,N_27166,N_27162);
and U27267 (N_27267,N_27158,N_27102);
or U27268 (N_27268,N_27156,N_27243);
xor U27269 (N_27269,N_27068,N_27145);
nor U27270 (N_27270,N_27236,N_27128);
and U27271 (N_27271,N_27000,N_27043);
or U27272 (N_27272,N_27124,N_27141);
nand U27273 (N_27273,N_27080,N_27033);
nor U27274 (N_27274,N_27218,N_27170);
xor U27275 (N_27275,N_27172,N_27113);
nor U27276 (N_27276,N_27040,N_27211);
and U27277 (N_27277,N_27193,N_27077);
nor U27278 (N_27278,N_27032,N_27107);
nor U27279 (N_27279,N_27073,N_27002);
nand U27280 (N_27280,N_27074,N_27210);
and U27281 (N_27281,N_27121,N_27209);
xor U27282 (N_27282,N_27007,N_27030);
nor U27283 (N_27283,N_27075,N_27085);
and U27284 (N_27284,N_27034,N_27104);
xor U27285 (N_27285,N_27059,N_27238);
nor U27286 (N_27286,N_27199,N_27192);
or U27287 (N_27287,N_27125,N_27150);
nand U27288 (N_27288,N_27176,N_27200);
xor U27289 (N_27289,N_27010,N_27087);
xor U27290 (N_27290,N_27097,N_27179);
or U27291 (N_27291,N_27070,N_27207);
or U27292 (N_27292,N_27230,N_27233);
nand U27293 (N_27293,N_27086,N_27039);
or U27294 (N_27294,N_27016,N_27212);
or U27295 (N_27295,N_27194,N_27042);
or U27296 (N_27296,N_27248,N_27114);
or U27297 (N_27297,N_27130,N_27183);
nor U27298 (N_27298,N_27082,N_27066);
or U27299 (N_27299,N_27220,N_27117);
and U27300 (N_27300,N_27242,N_27094);
xor U27301 (N_27301,N_27045,N_27231);
nand U27302 (N_27302,N_27052,N_27129);
and U27303 (N_27303,N_27160,N_27126);
xor U27304 (N_27304,N_27013,N_27191);
xnor U27305 (N_27305,N_27245,N_27076);
or U27306 (N_27306,N_27098,N_27008);
nor U27307 (N_27307,N_27055,N_27224);
or U27308 (N_27308,N_27180,N_27019);
xnor U27309 (N_27309,N_27168,N_27006);
or U27310 (N_27310,N_27153,N_27217);
nor U27311 (N_27311,N_27155,N_27175);
or U27312 (N_27312,N_27228,N_27127);
or U27313 (N_27313,N_27048,N_27169);
nor U27314 (N_27314,N_27110,N_27148);
nor U27315 (N_27315,N_27101,N_27044);
and U27316 (N_27316,N_27163,N_27235);
nand U27317 (N_27317,N_27105,N_27037);
nor U27318 (N_27318,N_27249,N_27241);
or U27319 (N_27319,N_27134,N_27111);
xnor U27320 (N_27320,N_27140,N_27035);
nor U27321 (N_27321,N_27181,N_27112);
nand U27322 (N_27322,N_27203,N_27092);
nand U27323 (N_27323,N_27029,N_27022);
nand U27324 (N_27324,N_27205,N_27161);
nand U27325 (N_27325,N_27106,N_27061);
nor U27326 (N_27326,N_27053,N_27143);
xnor U27327 (N_27327,N_27026,N_27064);
xor U27328 (N_27328,N_27063,N_27206);
and U27329 (N_27329,N_27147,N_27246);
nand U27330 (N_27330,N_27116,N_27185);
nand U27331 (N_27331,N_27021,N_27232);
xor U27332 (N_27332,N_27001,N_27099);
nand U27333 (N_27333,N_27100,N_27177);
or U27334 (N_27334,N_27089,N_27216);
xor U27335 (N_27335,N_27024,N_27157);
and U27336 (N_27336,N_27190,N_27078);
nor U27337 (N_27337,N_27144,N_27164);
nand U27338 (N_27338,N_27071,N_27154);
and U27339 (N_27339,N_27221,N_27051);
or U27340 (N_27340,N_27152,N_27208);
nand U27341 (N_27341,N_27088,N_27196);
or U27342 (N_27342,N_27115,N_27017);
or U27343 (N_27343,N_27188,N_27138);
xor U27344 (N_27344,N_27198,N_27202);
nor U27345 (N_27345,N_27011,N_27214);
and U27346 (N_27346,N_27137,N_27122);
nand U27347 (N_27347,N_27244,N_27123);
nand U27348 (N_27348,N_27136,N_27132);
and U27349 (N_27349,N_27213,N_27046);
or U27350 (N_27350,N_27038,N_27167);
xor U27351 (N_27351,N_27239,N_27186);
xnor U27352 (N_27352,N_27083,N_27060);
and U27353 (N_27353,N_27067,N_27204);
nor U27354 (N_27354,N_27095,N_27050);
or U27355 (N_27355,N_27103,N_27215);
nor U27356 (N_27356,N_27119,N_27072);
nand U27357 (N_27357,N_27219,N_27133);
and U27358 (N_27358,N_27247,N_27173);
nand U27359 (N_27359,N_27223,N_27184);
xor U27360 (N_27360,N_27093,N_27240);
nand U27361 (N_27361,N_27197,N_27135);
and U27362 (N_27362,N_27047,N_27182);
xor U27363 (N_27363,N_27062,N_27226);
and U27364 (N_27364,N_27084,N_27118);
nor U27365 (N_27365,N_27151,N_27056);
nor U27366 (N_27366,N_27108,N_27091);
nand U27367 (N_27367,N_27149,N_27079);
xor U27368 (N_27368,N_27004,N_27187);
xor U27369 (N_27369,N_27049,N_27025);
nor U27370 (N_27370,N_27005,N_27225);
nor U27371 (N_27371,N_27081,N_27189);
nand U27372 (N_27372,N_27171,N_27222);
xor U27373 (N_27373,N_27031,N_27139);
xnor U27374 (N_27374,N_27012,N_27027);
nand U27375 (N_27375,N_27091,N_27101);
or U27376 (N_27376,N_27051,N_27097);
xnor U27377 (N_27377,N_27076,N_27017);
nand U27378 (N_27378,N_27031,N_27003);
nor U27379 (N_27379,N_27012,N_27235);
and U27380 (N_27380,N_27057,N_27204);
nor U27381 (N_27381,N_27121,N_27232);
nand U27382 (N_27382,N_27050,N_27013);
nor U27383 (N_27383,N_27114,N_27244);
nand U27384 (N_27384,N_27029,N_27102);
and U27385 (N_27385,N_27239,N_27180);
nand U27386 (N_27386,N_27173,N_27137);
nand U27387 (N_27387,N_27215,N_27235);
nand U27388 (N_27388,N_27145,N_27073);
nand U27389 (N_27389,N_27006,N_27076);
xor U27390 (N_27390,N_27196,N_27162);
nor U27391 (N_27391,N_27063,N_27101);
nand U27392 (N_27392,N_27081,N_27125);
xor U27393 (N_27393,N_27189,N_27033);
and U27394 (N_27394,N_27217,N_27134);
nand U27395 (N_27395,N_27028,N_27233);
or U27396 (N_27396,N_27248,N_27097);
or U27397 (N_27397,N_27232,N_27130);
nor U27398 (N_27398,N_27011,N_27202);
and U27399 (N_27399,N_27247,N_27159);
nand U27400 (N_27400,N_27070,N_27090);
nand U27401 (N_27401,N_27035,N_27204);
nor U27402 (N_27402,N_27178,N_27223);
nand U27403 (N_27403,N_27041,N_27154);
xor U27404 (N_27404,N_27086,N_27103);
xnor U27405 (N_27405,N_27001,N_27018);
or U27406 (N_27406,N_27054,N_27092);
xor U27407 (N_27407,N_27191,N_27094);
nand U27408 (N_27408,N_27168,N_27193);
or U27409 (N_27409,N_27003,N_27231);
nand U27410 (N_27410,N_27097,N_27164);
xor U27411 (N_27411,N_27208,N_27080);
and U27412 (N_27412,N_27091,N_27202);
or U27413 (N_27413,N_27122,N_27195);
xor U27414 (N_27414,N_27119,N_27062);
or U27415 (N_27415,N_27235,N_27196);
xor U27416 (N_27416,N_27188,N_27243);
or U27417 (N_27417,N_27161,N_27045);
xor U27418 (N_27418,N_27179,N_27174);
nand U27419 (N_27419,N_27248,N_27195);
nand U27420 (N_27420,N_27028,N_27197);
nand U27421 (N_27421,N_27163,N_27158);
xor U27422 (N_27422,N_27056,N_27023);
nor U27423 (N_27423,N_27238,N_27031);
or U27424 (N_27424,N_27145,N_27036);
or U27425 (N_27425,N_27014,N_27067);
and U27426 (N_27426,N_27145,N_27085);
or U27427 (N_27427,N_27086,N_27138);
nor U27428 (N_27428,N_27245,N_27027);
nand U27429 (N_27429,N_27152,N_27063);
xnor U27430 (N_27430,N_27045,N_27190);
xnor U27431 (N_27431,N_27133,N_27001);
and U27432 (N_27432,N_27150,N_27049);
and U27433 (N_27433,N_27006,N_27073);
and U27434 (N_27434,N_27176,N_27121);
xnor U27435 (N_27435,N_27134,N_27133);
xor U27436 (N_27436,N_27018,N_27083);
and U27437 (N_27437,N_27228,N_27073);
or U27438 (N_27438,N_27154,N_27231);
nor U27439 (N_27439,N_27145,N_27195);
xnor U27440 (N_27440,N_27039,N_27030);
xor U27441 (N_27441,N_27228,N_27083);
nand U27442 (N_27442,N_27076,N_27114);
nor U27443 (N_27443,N_27025,N_27004);
nor U27444 (N_27444,N_27072,N_27106);
xnor U27445 (N_27445,N_27110,N_27238);
or U27446 (N_27446,N_27171,N_27172);
nand U27447 (N_27447,N_27104,N_27046);
and U27448 (N_27448,N_27161,N_27144);
nor U27449 (N_27449,N_27094,N_27057);
xor U27450 (N_27450,N_27198,N_27034);
nand U27451 (N_27451,N_27046,N_27225);
or U27452 (N_27452,N_27048,N_27201);
and U27453 (N_27453,N_27169,N_27215);
nand U27454 (N_27454,N_27217,N_27214);
or U27455 (N_27455,N_27034,N_27073);
nand U27456 (N_27456,N_27111,N_27048);
nand U27457 (N_27457,N_27003,N_27162);
nor U27458 (N_27458,N_27229,N_27130);
nand U27459 (N_27459,N_27111,N_27186);
or U27460 (N_27460,N_27013,N_27194);
and U27461 (N_27461,N_27087,N_27152);
xnor U27462 (N_27462,N_27066,N_27000);
xnor U27463 (N_27463,N_27213,N_27220);
nand U27464 (N_27464,N_27177,N_27155);
and U27465 (N_27465,N_27229,N_27127);
xnor U27466 (N_27466,N_27172,N_27006);
nor U27467 (N_27467,N_27119,N_27150);
nand U27468 (N_27468,N_27105,N_27079);
nand U27469 (N_27469,N_27190,N_27181);
xnor U27470 (N_27470,N_27139,N_27170);
and U27471 (N_27471,N_27091,N_27126);
nor U27472 (N_27472,N_27224,N_27045);
nand U27473 (N_27473,N_27247,N_27187);
nand U27474 (N_27474,N_27000,N_27168);
nand U27475 (N_27475,N_27086,N_27051);
nor U27476 (N_27476,N_27095,N_27145);
nand U27477 (N_27477,N_27033,N_27224);
or U27478 (N_27478,N_27234,N_27225);
xor U27479 (N_27479,N_27047,N_27025);
nor U27480 (N_27480,N_27053,N_27068);
nand U27481 (N_27481,N_27054,N_27217);
or U27482 (N_27482,N_27020,N_27222);
nor U27483 (N_27483,N_27140,N_27070);
nand U27484 (N_27484,N_27230,N_27122);
nand U27485 (N_27485,N_27188,N_27060);
and U27486 (N_27486,N_27239,N_27147);
and U27487 (N_27487,N_27197,N_27164);
nor U27488 (N_27488,N_27034,N_27006);
xor U27489 (N_27489,N_27132,N_27003);
xnor U27490 (N_27490,N_27042,N_27199);
or U27491 (N_27491,N_27144,N_27218);
and U27492 (N_27492,N_27223,N_27091);
and U27493 (N_27493,N_27010,N_27064);
or U27494 (N_27494,N_27029,N_27198);
or U27495 (N_27495,N_27129,N_27081);
nand U27496 (N_27496,N_27049,N_27127);
and U27497 (N_27497,N_27233,N_27015);
or U27498 (N_27498,N_27207,N_27089);
nand U27499 (N_27499,N_27221,N_27021);
nor U27500 (N_27500,N_27481,N_27485);
or U27501 (N_27501,N_27309,N_27370);
or U27502 (N_27502,N_27276,N_27388);
and U27503 (N_27503,N_27442,N_27338);
xor U27504 (N_27504,N_27415,N_27319);
or U27505 (N_27505,N_27264,N_27283);
or U27506 (N_27506,N_27457,N_27460);
and U27507 (N_27507,N_27324,N_27286);
nand U27508 (N_27508,N_27311,N_27459);
nor U27509 (N_27509,N_27348,N_27463);
or U27510 (N_27510,N_27380,N_27429);
nand U27511 (N_27511,N_27312,N_27361);
nand U27512 (N_27512,N_27328,N_27474);
xnor U27513 (N_27513,N_27495,N_27341);
nand U27514 (N_27514,N_27456,N_27322);
and U27515 (N_27515,N_27398,N_27473);
and U27516 (N_27516,N_27377,N_27381);
nor U27517 (N_27517,N_27360,N_27493);
xor U27518 (N_27518,N_27339,N_27342);
nor U27519 (N_27519,N_27395,N_27372);
and U27520 (N_27520,N_27303,N_27336);
or U27521 (N_27521,N_27394,N_27428);
nor U27522 (N_27522,N_27424,N_27335);
or U27523 (N_27523,N_27347,N_27332);
xnor U27524 (N_27524,N_27273,N_27318);
nor U27525 (N_27525,N_27354,N_27468);
or U27526 (N_27526,N_27497,N_27301);
or U27527 (N_27527,N_27490,N_27453);
nor U27528 (N_27528,N_27365,N_27475);
nor U27529 (N_27529,N_27469,N_27467);
and U27530 (N_27530,N_27254,N_27447);
nor U27531 (N_27531,N_27480,N_27340);
nor U27532 (N_27532,N_27320,N_27408);
nor U27533 (N_27533,N_27329,N_27326);
or U27534 (N_27534,N_27257,N_27421);
and U27535 (N_27535,N_27357,N_27393);
nor U27536 (N_27536,N_27337,N_27484);
xnor U27537 (N_27537,N_27269,N_27378);
nand U27538 (N_27538,N_27419,N_27349);
nand U27539 (N_27539,N_27278,N_27439);
xnor U27540 (N_27540,N_27478,N_27376);
nand U27541 (N_27541,N_27280,N_27367);
nand U27542 (N_27542,N_27444,N_27288);
or U27543 (N_27543,N_27374,N_27253);
and U27544 (N_27544,N_27445,N_27434);
nor U27545 (N_27545,N_27363,N_27386);
xnor U27546 (N_27546,N_27477,N_27255);
and U27547 (N_27547,N_27413,N_27427);
nor U27548 (N_27548,N_27300,N_27330);
and U27549 (N_27549,N_27496,N_27275);
and U27550 (N_27550,N_27268,N_27359);
nor U27551 (N_27551,N_27316,N_27383);
nor U27552 (N_27552,N_27299,N_27295);
and U27553 (N_27553,N_27410,N_27289);
or U27554 (N_27554,N_27290,N_27498);
and U27555 (N_27555,N_27431,N_27317);
and U27556 (N_27556,N_27375,N_27479);
nand U27557 (N_27557,N_27440,N_27250);
or U27558 (N_27558,N_27455,N_27256);
xor U27559 (N_27559,N_27401,N_27302);
xnor U27560 (N_27560,N_27272,N_27356);
and U27561 (N_27561,N_27279,N_27389);
or U27562 (N_27562,N_27314,N_27449);
xnor U27563 (N_27563,N_27409,N_27282);
nor U27564 (N_27564,N_27266,N_27271);
and U27565 (N_27565,N_27373,N_27443);
nor U27566 (N_27566,N_27458,N_27452);
or U27567 (N_27567,N_27284,N_27426);
nand U27568 (N_27568,N_27472,N_27450);
and U27569 (N_27569,N_27306,N_27392);
xnor U27570 (N_27570,N_27406,N_27464);
or U27571 (N_27571,N_27400,N_27397);
xor U27572 (N_27572,N_27323,N_27446);
nor U27573 (N_27573,N_27385,N_27267);
and U27574 (N_27574,N_27499,N_27277);
nor U27575 (N_27575,N_27313,N_27344);
nand U27576 (N_27576,N_27294,N_27404);
xnor U27577 (N_27577,N_27403,N_27334);
xor U27578 (N_27578,N_27263,N_27258);
xnor U27579 (N_27579,N_27327,N_27345);
xor U27580 (N_27580,N_27382,N_27451);
nand U27581 (N_27581,N_27414,N_27270);
or U27582 (N_27582,N_27425,N_27492);
or U27583 (N_27583,N_27417,N_27430);
nor U27584 (N_27584,N_27416,N_27364);
nand U27585 (N_27585,N_27287,N_27402);
or U27586 (N_27586,N_27351,N_27261);
or U27587 (N_27587,N_27387,N_27259);
xor U27588 (N_27588,N_27297,N_27494);
and U27589 (N_27589,N_27448,N_27412);
nor U27590 (N_27590,N_27350,N_27441);
xnor U27591 (N_27591,N_27384,N_27321);
nor U27592 (N_27592,N_27399,N_27281);
xor U27593 (N_27593,N_27438,N_27353);
nor U27594 (N_27594,N_27422,N_27298);
xnor U27595 (N_27595,N_27487,N_27405);
nor U27596 (N_27596,N_27292,N_27423);
or U27597 (N_27597,N_27489,N_27462);
xnor U27598 (N_27598,N_27418,N_27331);
nand U27599 (N_27599,N_27396,N_27465);
or U27600 (N_27600,N_27432,N_27461);
or U27601 (N_27601,N_27491,N_27407);
xnor U27602 (N_27602,N_27358,N_27291);
xor U27603 (N_27603,N_27437,N_27488);
nand U27604 (N_27604,N_27483,N_27471);
or U27605 (N_27605,N_27379,N_27466);
nand U27606 (N_27606,N_27293,N_27476);
or U27607 (N_27607,N_27436,N_27343);
and U27608 (N_27608,N_27352,N_27482);
nor U27609 (N_27609,N_27260,N_27308);
and U27610 (N_27610,N_27285,N_27251);
xor U27611 (N_27611,N_27420,N_27391);
or U27612 (N_27612,N_27433,N_27355);
and U27613 (N_27613,N_27333,N_27307);
nor U27614 (N_27614,N_27265,N_27362);
xnor U27615 (N_27615,N_27366,N_27310);
nor U27616 (N_27616,N_27252,N_27435);
nor U27617 (N_27617,N_27411,N_27274);
and U27618 (N_27618,N_27262,N_27304);
nand U27619 (N_27619,N_27325,N_27368);
nor U27620 (N_27620,N_27346,N_27315);
nor U27621 (N_27621,N_27454,N_27296);
nand U27622 (N_27622,N_27486,N_27371);
xnor U27623 (N_27623,N_27470,N_27369);
or U27624 (N_27624,N_27305,N_27390);
nand U27625 (N_27625,N_27311,N_27444);
nand U27626 (N_27626,N_27267,N_27490);
and U27627 (N_27627,N_27333,N_27258);
nand U27628 (N_27628,N_27395,N_27277);
xor U27629 (N_27629,N_27399,N_27305);
or U27630 (N_27630,N_27461,N_27329);
and U27631 (N_27631,N_27298,N_27437);
nand U27632 (N_27632,N_27264,N_27418);
nand U27633 (N_27633,N_27252,N_27390);
and U27634 (N_27634,N_27257,N_27303);
xor U27635 (N_27635,N_27395,N_27285);
nor U27636 (N_27636,N_27369,N_27429);
nand U27637 (N_27637,N_27453,N_27316);
nand U27638 (N_27638,N_27307,N_27399);
or U27639 (N_27639,N_27318,N_27372);
or U27640 (N_27640,N_27453,N_27472);
xnor U27641 (N_27641,N_27342,N_27465);
xnor U27642 (N_27642,N_27320,N_27350);
and U27643 (N_27643,N_27462,N_27271);
xor U27644 (N_27644,N_27315,N_27430);
nand U27645 (N_27645,N_27305,N_27414);
nor U27646 (N_27646,N_27413,N_27265);
nor U27647 (N_27647,N_27299,N_27337);
and U27648 (N_27648,N_27432,N_27407);
xor U27649 (N_27649,N_27319,N_27422);
and U27650 (N_27650,N_27251,N_27274);
nand U27651 (N_27651,N_27426,N_27481);
xnor U27652 (N_27652,N_27413,N_27465);
xor U27653 (N_27653,N_27418,N_27442);
nand U27654 (N_27654,N_27392,N_27334);
and U27655 (N_27655,N_27472,N_27433);
nor U27656 (N_27656,N_27353,N_27313);
or U27657 (N_27657,N_27334,N_27369);
nand U27658 (N_27658,N_27419,N_27335);
nand U27659 (N_27659,N_27356,N_27485);
xor U27660 (N_27660,N_27405,N_27474);
xor U27661 (N_27661,N_27319,N_27431);
and U27662 (N_27662,N_27390,N_27436);
xor U27663 (N_27663,N_27451,N_27419);
nand U27664 (N_27664,N_27270,N_27421);
xnor U27665 (N_27665,N_27379,N_27319);
nor U27666 (N_27666,N_27271,N_27453);
xor U27667 (N_27667,N_27373,N_27452);
or U27668 (N_27668,N_27460,N_27492);
nand U27669 (N_27669,N_27258,N_27341);
nor U27670 (N_27670,N_27304,N_27389);
xnor U27671 (N_27671,N_27399,N_27442);
nand U27672 (N_27672,N_27378,N_27309);
xor U27673 (N_27673,N_27351,N_27386);
and U27674 (N_27674,N_27293,N_27414);
or U27675 (N_27675,N_27330,N_27426);
xor U27676 (N_27676,N_27433,N_27346);
nor U27677 (N_27677,N_27441,N_27484);
nor U27678 (N_27678,N_27344,N_27400);
and U27679 (N_27679,N_27427,N_27383);
nand U27680 (N_27680,N_27338,N_27274);
and U27681 (N_27681,N_27280,N_27381);
or U27682 (N_27682,N_27317,N_27335);
nand U27683 (N_27683,N_27381,N_27266);
or U27684 (N_27684,N_27318,N_27423);
nor U27685 (N_27685,N_27277,N_27476);
xnor U27686 (N_27686,N_27479,N_27354);
or U27687 (N_27687,N_27353,N_27493);
and U27688 (N_27688,N_27396,N_27386);
nand U27689 (N_27689,N_27366,N_27300);
or U27690 (N_27690,N_27421,N_27274);
nor U27691 (N_27691,N_27324,N_27262);
xor U27692 (N_27692,N_27345,N_27391);
and U27693 (N_27693,N_27317,N_27387);
nand U27694 (N_27694,N_27333,N_27476);
xnor U27695 (N_27695,N_27495,N_27315);
and U27696 (N_27696,N_27287,N_27316);
nor U27697 (N_27697,N_27467,N_27281);
xnor U27698 (N_27698,N_27257,N_27331);
nand U27699 (N_27699,N_27334,N_27373);
nand U27700 (N_27700,N_27373,N_27375);
and U27701 (N_27701,N_27456,N_27457);
and U27702 (N_27702,N_27328,N_27272);
or U27703 (N_27703,N_27374,N_27482);
xnor U27704 (N_27704,N_27333,N_27337);
or U27705 (N_27705,N_27487,N_27253);
nand U27706 (N_27706,N_27411,N_27406);
and U27707 (N_27707,N_27479,N_27457);
nand U27708 (N_27708,N_27305,N_27252);
nor U27709 (N_27709,N_27409,N_27427);
nor U27710 (N_27710,N_27433,N_27417);
xnor U27711 (N_27711,N_27371,N_27469);
nor U27712 (N_27712,N_27287,N_27386);
nor U27713 (N_27713,N_27493,N_27329);
xor U27714 (N_27714,N_27429,N_27326);
nor U27715 (N_27715,N_27428,N_27402);
nor U27716 (N_27716,N_27272,N_27373);
and U27717 (N_27717,N_27322,N_27265);
nand U27718 (N_27718,N_27472,N_27458);
or U27719 (N_27719,N_27250,N_27432);
xnor U27720 (N_27720,N_27478,N_27443);
nand U27721 (N_27721,N_27462,N_27485);
or U27722 (N_27722,N_27314,N_27444);
and U27723 (N_27723,N_27389,N_27366);
nor U27724 (N_27724,N_27346,N_27497);
xnor U27725 (N_27725,N_27380,N_27489);
xor U27726 (N_27726,N_27408,N_27411);
and U27727 (N_27727,N_27456,N_27401);
nand U27728 (N_27728,N_27346,N_27429);
or U27729 (N_27729,N_27393,N_27492);
xor U27730 (N_27730,N_27321,N_27411);
nor U27731 (N_27731,N_27347,N_27488);
or U27732 (N_27732,N_27415,N_27370);
nand U27733 (N_27733,N_27251,N_27284);
or U27734 (N_27734,N_27479,N_27488);
and U27735 (N_27735,N_27468,N_27463);
or U27736 (N_27736,N_27327,N_27496);
or U27737 (N_27737,N_27483,N_27274);
xor U27738 (N_27738,N_27463,N_27293);
and U27739 (N_27739,N_27437,N_27431);
nor U27740 (N_27740,N_27312,N_27315);
xnor U27741 (N_27741,N_27265,N_27467);
nor U27742 (N_27742,N_27269,N_27275);
or U27743 (N_27743,N_27295,N_27296);
or U27744 (N_27744,N_27429,N_27381);
nand U27745 (N_27745,N_27374,N_27258);
nor U27746 (N_27746,N_27285,N_27427);
nand U27747 (N_27747,N_27407,N_27339);
and U27748 (N_27748,N_27280,N_27483);
and U27749 (N_27749,N_27497,N_27433);
nor U27750 (N_27750,N_27654,N_27506);
nand U27751 (N_27751,N_27698,N_27634);
or U27752 (N_27752,N_27500,N_27726);
xnor U27753 (N_27753,N_27731,N_27734);
or U27754 (N_27754,N_27741,N_27701);
xor U27755 (N_27755,N_27720,N_27614);
xnor U27756 (N_27756,N_27704,N_27607);
nor U27757 (N_27757,N_27583,N_27718);
nand U27758 (N_27758,N_27655,N_27564);
nor U27759 (N_27759,N_27590,N_27642);
xnor U27760 (N_27760,N_27603,N_27586);
xnor U27761 (N_27761,N_27703,N_27572);
nor U27762 (N_27762,N_27580,N_27695);
and U27763 (N_27763,N_27576,N_27524);
xnor U27764 (N_27764,N_27566,N_27595);
nand U27765 (N_27765,N_27507,N_27615);
or U27766 (N_27766,N_27693,N_27717);
or U27767 (N_27767,N_27543,N_27570);
nand U27768 (N_27768,N_27582,N_27640);
nor U27769 (N_27769,N_27697,N_27567);
xnor U27770 (N_27770,N_27732,N_27530);
nand U27771 (N_27771,N_27633,N_27581);
and U27772 (N_27772,N_27645,N_27558);
or U27773 (N_27773,N_27600,N_27554);
and U27774 (N_27774,N_27544,N_27516);
or U27775 (N_27775,N_27647,N_27626);
or U27776 (N_27776,N_27523,N_27534);
nor U27777 (N_27777,N_27522,N_27670);
and U27778 (N_27778,N_27539,N_27521);
nor U27779 (N_27779,N_27632,N_27520);
xor U27780 (N_27780,N_27676,N_27688);
and U27781 (N_27781,N_27672,N_27605);
or U27782 (N_27782,N_27628,N_27702);
xnor U27783 (N_27783,N_27608,N_27706);
or U27784 (N_27784,N_27743,N_27664);
nor U27785 (N_27785,N_27638,N_27501);
nand U27786 (N_27786,N_27598,N_27659);
nand U27787 (N_27787,N_27735,N_27678);
or U27788 (N_27788,N_27518,N_27677);
or U27789 (N_27789,N_27675,N_27641);
and U27790 (N_27790,N_27574,N_27616);
and U27791 (N_27791,N_27680,N_27740);
or U27792 (N_27792,N_27656,N_27591);
nor U27793 (N_27793,N_27571,N_27728);
nor U27794 (N_27794,N_27660,N_27681);
nor U27795 (N_27795,N_27588,N_27708);
nor U27796 (N_27796,N_27705,N_27631);
xor U27797 (N_27797,N_27589,N_27696);
and U27798 (N_27798,N_27744,N_27739);
nand U27799 (N_27799,N_27613,N_27716);
nand U27800 (N_27800,N_27714,N_27537);
xor U27801 (N_27801,N_27617,N_27612);
or U27802 (N_27802,N_27721,N_27709);
nor U27803 (N_27803,N_27729,N_27687);
nor U27804 (N_27804,N_27668,N_27649);
nor U27805 (N_27805,N_27563,N_27749);
xor U27806 (N_27806,N_27587,N_27609);
nand U27807 (N_27807,N_27604,N_27528);
nand U27808 (N_27808,N_27690,N_27723);
nand U27809 (N_27809,N_27556,N_27549);
and U27810 (N_27810,N_27514,N_27541);
nor U27811 (N_27811,N_27618,N_27665);
or U27812 (N_27812,N_27531,N_27747);
nor U27813 (N_27813,N_27686,N_27635);
and U27814 (N_27814,N_27636,N_27673);
and U27815 (N_27815,N_27551,N_27658);
and U27816 (N_27816,N_27577,N_27637);
and U27817 (N_27817,N_27646,N_27684);
nand U27818 (N_27818,N_27727,N_27713);
xor U27819 (N_27819,N_27512,N_27578);
and U27820 (N_27820,N_27509,N_27525);
and U27821 (N_27821,N_27532,N_27517);
xor U27822 (N_27822,N_27685,N_27553);
nand U27823 (N_27823,N_27663,N_27742);
xnor U27824 (N_27824,N_27527,N_27529);
xnor U27825 (N_27825,N_27503,N_27573);
xor U27826 (N_27826,N_27643,N_27594);
and U27827 (N_27827,N_27624,N_27565);
nor U27828 (N_27828,N_27515,N_27505);
nor U27829 (N_27829,N_27657,N_27715);
xor U27830 (N_27830,N_27644,N_27599);
and U27831 (N_27831,N_27682,N_27519);
and U27832 (N_27832,N_27546,N_27666);
xor U27833 (N_27833,N_27569,N_27535);
and U27834 (N_27834,N_27653,N_27691);
nor U27835 (N_27835,N_27737,N_27540);
nor U27836 (N_27836,N_27504,N_27526);
and U27837 (N_27837,N_27597,N_27555);
nand U27838 (N_27838,N_27700,N_27662);
xor U27839 (N_27839,N_27538,N_27606);
or U27840 (N_27840,N_27585,N_27560);
xnor U27841 (N_27841,N_27508,N_27510);
or U27842 (N_27842,N_27710,N_27610);
xor U27843 (N_27843,N_27619,N_27650);
xnor U27844 (N_27844,N_27502,N_27559);
or U27845 (N_27845,N_27561,N_27557);
xnor U27846 (N_27846,N_27547,N_27542);
or U27847 (N_27847,N_27674,N_27620);
xor U27848 (N_27848,N_27629,N_27648);
and U27849 (N_27849,N_27745,N_27623);
and U27850 (N_27850,N_27711,N_27621);
and U27851 (N_27851,N_27722,N_27513);
nor U27852 (N_27852,N_27736,N_27592);
or U27853 (N_27853,N_27712,N_27730);
xnor U27854 (N_27854,N_27601,N_27545);
xnor U27855 (N_27855,N_27746,N_27667);
xor U27856 (N_27856,N_27550,N_27602);
nor U27857 (N_27857,N_27627,N_27683);
nand U27858 (N_27858,N_27719,N_27679);
nor U27859 (N_27859,N_27625,N_27511);
nor U27860 (N_27860,N_27724,N_27692);
nand U27861 (N_27861,N_27748,N_27671);
xor U27862 (N_27862,N_27548,N_27738);
and U27863 (N_27863,N_27536,N_27651);
nand U27864 (N_27864,N_27533,N_27669);
nand U27865 (N_27865,N_27593,N_27575);
and U27866 (N_27866,N_27689,N_27630);
and U27867 (N_27867,N_27699,N_27733);
and U27868 (N_27868,N_27584,N_27622);
nor U27869 (N_27869,N_27694,N_27707);
nand U27870 (N_27870,N_27611,N_27562);
nand U27871 (N_27871,N_27552,N_27639);
and U27872 (N_27872,N_27725,N_27568);
nor U27873 (N_27873,N_27579,N_27661);
or U27874 (N_27874,N_27652,N_27596);
or U27875 (N_27875,N_27551,N_27608);
or U27876 (N_27876,N_27713,N_27503);
or U27877 (N_27877,N_27736,N_27628);
nand U27878 (N_27878,N_27642,N_27729);
nand U27879 (N_27879,N_27611,N_27661);
xnor U27880 (N_27880,N_27562,N_27552);
nand U27881 (N_27881,N_27567,N_27719);
xor U27882 (N_27882,N_27500,N_27585);
or U27883 (N_27883,N_27708,N_27703);
and U27884 (N_27884,N_27747,N_27603);
xor U27885 (N_27885,N_27565,N_27576);
nor U27886 (N_27886,N_27660,N_27588);
nor U27887 (N_27887,N_27624,N_27549);
xnor U27888 (N_27888,N_27646,N_27694);
nand U27889 (N_27889,N_27715,N_27699);
xor U27890 (N_27890,N_27527,N_27717);
nor U27891 (N_27891,N_27634,N_27600);
nor U27892 (N_27892,N_27549,N_27518);
nor U27893 (N_27893,N_27713,N_27685);
nand U27894 (N_27894,N_27662,N_27678);
xnor U27895 (N_27895,N_27698,N_27572);
nand U27896 (N_27896,N_27527,N_27681);
nor U27897 (N_27897,N_27692,N_27502);
nand U27898 (N_27898,N_27516,N_27629);
nand U27899 (N_27899,N_27513,N_27609);
xnor U27900 (N_27900,N_27685,N_27602);
xnor U27901 (N_27901,N_27529,N_27608);
and U27902 (N_27902,N_27594,N_27689);
and U27903 (N_27903,N_27629,N_27665);
and U27904 (N_27904,N_27683,N_27599);
and U27905 (N_27905,N_27662,N_27631);
and U27906 (N_27906,N_27745,N_27566);
nand U27907 (N_27907,N_27600,N_27509);
nor U27908 (N_27908,N_27536,N_27590);
nor U27909 (N_27909,N_27694,N_27738);
xor U27910 (N_27910,N_27705,N_27643);
nand U27911 (N_27911,N_27588,N_27536);
nor U27912 (N_27912,N_27545,N_27550);
xor U27913 (N_27913,N_27608,N_27652);
or U27914 (N_27914,N_27635,N_27621);
or U27915 (N_27915,N_27549,N_27676);
and U27916 (N_27916,N_27710,N_27711);
and U27917 (N_27917,N_27645,N_27635);
and U27918 (N_27918,N_27602,N_27656);
or U27919 (N_27919,N_27585,N_27594);
xor U27920 (N_27920,N_27691,N_27733);
or U27921 (N_27921,N_27556,N_27731);
nand U27922 (N_27922,N_27550,N_27701);
xnor U27923 (N_27923,N_27644,N_27585);
nand U27924 (N_27924,N_27647,N_27694);
xor U27925 (N_27925,N_27699,N_27616);
or U27926 (N_27926,N_27612,N_27560);
nor U27927 (N_27927,N_27504,N_27672);
or U27928 (N_27928,N_27519,N_27580);
nor U27929 (N_27929,N_27668,N_27581);
or U27930 (N_27930,N_27534,N_27689);
nand U27931 (N_27931,N_27729,N_27535);
nor U27932 (N_27932,N_27628,N_27554);
and U27933 (N_27933,N_27663,N_27550);
nand U27934 (N_27934,N_27617,N_27632);
or U27935 (N_27935,N_27696,N_27508);
xor U27936 (N_27936,N_27519,N_27641);
or U27937 (N_27937,N_27732,N_27673);
or U27938 (N_27938,N_27623,N_27537);
and U27939 (N_27939,N_27572,N_27548);
and U27940 (N_27940,N_27618,N_27538);
and U27941 (N_27941,N_27622,N_27720);
nand U27942 (N_27942,N_27501,N_27522);
nand U27943 (N_27943,N_27643,N_27575);
nor U27944 (N_27944,N_27649,N_27575);
nor U27945 (N_27945,N_27601,N_27541);
or U27946 (N_27946,N_27562,N_27695);
nor U27947 (N_27947,N_27520,N_27723);
nor U27948 (N_27948,N_27563,N_27723);
and U27949 (N_27949,N_27607,N_27629);
nor U27950 (N_27950,N_27522,N_27526);
nand U27951 (N_27951,N_27739,N_27643);
xor U27952 (N_27952,N_27743,N_27668);
or U27953 (N_27953,N_27519,N_27535);
or U27954 (N_27954,N_27531,N_27569);
and U27955 (N_27955,N_27653,N_27639);
and U27956 (N_27956,N_27500,N_27707);
nand U27957 (N_27957,N_27671,N_27514);
nor U27958 (N_27958,N_27599,N_27530);
nand U27959 (N_27959,N_27747,N_27703);
nand U27960 (N_27960,N_27695,N_27652);
xor U27961 (N_27961,N_27578,N_27535);
xnor U27962 (N_27962,N_27656,N_27731);
nand U27963 (N_27963,N_27697,N_27644);
or U27964 (N_27964,N_27550,N_27574);
or U27965 (N_27965,N_27691,N_27680);
nand U27966 (N_27966,N_27695,N_27712);
nor U27967 (N_27967,N_27644,N_27584);
nand U27968 (N_27968,N_27652,N_27581);
or U27969 (N_27969,N_27714,N_27622);
xor U27970 (N_27970,N_27612,N_27749);
nand U27971 (N_27971,N_27653,N_27733);
nand U27972 (N_27972,N_27738,N_27664);
or U27973 (N_27973,N_27561,N_27576);
xor U27974 (N_27974,N_27645,N_27596);
nand U27975 (N_27975,N_27611,N_27543);
xnor U27976 (N_27976,N_27586,N_27693);
nor U27977 (N_27977,N_27529,N_27683);
and U27978 (N_27978,N_27504,N_27534);
nand U27979 (N_27979,N_27631,N_27651);
xor U27980 (N_27980,N_27729,N_27656);
and U27981 (N_27981,N_27682,N_27518);
nor U27982 (N_27982,N_27690,N_27676);
or U27983 (N_27983,N_27675,N_27661);
xor U27984 (N_27984,N_27608,N_27705);
nand U27985 (N_27985,N_27504,N_27656);
or U27986 (N_27986,N_27535,N_27512);
xor U27987 (N_27987,N_27711,N_27593);
nor U27988 (N_27988,N_27516,N_27520);
nor U27989 (N_27989,N_27625,N_27527);
xnor U27990 (N_27990,N_27679,N_27676);
nor U27991 (N_27991,N_27551,N_27639);
xor U27992 (N_27992,N_27563,N_27617);
or U27993 (N_27993,N_27690,N_27711);
and U27994 (N_27994,N_27596,N_27555);
nor U27995 (N_27995,N_27681,N_27532);
and U27996 (N_27996,N_27714,N_27725);
and U27997 (N_27997,N_27515,N_27689);
xor U27998 (N_27998,N_27657,N_27705);
nand U27999 (N_27999,N_27698,N_27507);
nand U28000 (N_28000,N_27773,N_27875);
xnor U28001 (N_28001,N_27766,N_27783);
xnor U28002 (N_28002,N_27996,N_27913);
or U28003 (N_28003,N_27842,N_27889);
nand U28004 (N_28004,N_27919,N_27801);
nor U28005 (N_28005,N_27781,N_27943);
nor U28006 (N_28006,N_27771,N_27776);
and U28007 (N_28007,N_27917,N_27948);
xnor U28008 (N_28008,N_27908,N_27753);
nand U28009 (N_28009,N_27969,N_27861);
and U28010 (N_28010,N_27965,N_27864);
or U28011 (N_28011,N_27795,N_27854);
or U28012 (N_28012,N_27871,N_27934);
or U28013 (N_28013,N_27903,N_27900);
nor U28014 (N_28014,N_27761,N_27987);
nor U28015 (N_28015,N_27835,N_27961);
and U28016 (N_28016,N_27811,N_27905);
nor U28017 (N_28017,N_27865,N_27812);
nor U28018 (N_28018,N_27976,N_27981);
and U28019 (N_28019,N_27759,N_27847);
xor U28020 (N_28020,N_27798,N_27879);
xor U28021 (N_28021,N_27760,N_27848);
nand U28022 (N_28022,N_27912,N_27858);
nor U28023 (N_28023,N_27991,N_27866);
xnor U28024 (N_28024,N_27957,N_27886);
nor U28025 (N_28025,N_27916,N_27769);
and U28026 (N_28026,N_27821,N_27804);
nand U28027 (N_28027,N_27953,N_27809);
xor U28028 (N_28028,N_27844,N_27873);
xnor U28029 (N_28029,N_27883,N_27885);
xnor U28030 (N_28030,N_27929,N_27754);
and U28031 (N_28031,N_27995,N_27777);
xor U28032 (N_28032,N_27963,N_27926);
nand U28033 (N_28033,N_27980,N_27815);
nor U28034 (N_28034,N_27951,N_27837);
nand U28035 (N_28035,N_27925,N_27895);
and U28036 (N_28036,N_27849,N_27911);
nor U28037 (N_28037,N_27938,N_27958);
xor U28038 (N_28038,N_27756,N_27985);
nor U28039 (N_28039,N_27792,N_27762);
nand U28040 (N_28040,N_27874,N_27990);
or U28041 (N_28041,N_27878,N_27841);
nand U28042 (N_28042,N_27805,N_27971);
or U28043 (N_28043,N_27922,N_27876);
or U28044 (N_28044,N_27782,N_27898);
or U28045 (N_28045,N_27860,N_27877);
or U28046 (N_28046,N_27832,N_27954);
and U28047 (N_28047,N_27799,N_27850);
nor U28048 (N_28048,N_27775,N_27869);
or U28049 (N_28049,N_27863,N_27793);
and U28050 (N_28050,N_27867,N_27992);
or U28051 (N_28051,N_27808,N_27767);
xor U28052 (N_28052,N_27785,N_27755);
or U28053 (N_28053,N_27906,N_27824);
nand U28054 (N_28054,N_27882,N_27920);
or U28055 (N_28055,N_27802,N_27820);
and U28056 (N_28056,N_27946,N_27839);
nand U28057 (N_28057,N_27778,N_27870);
nor U28058 (N_28058,N_27803,N_27894);
and U28059 (N_28059,N_27765,N_27868);
nand U28060 (N_28060,N_27904,N_27955);
or U28061 (N_28061,N_27838,N_27977);
and U28062 (N_28062,N_27986,N_27822);
and U28063 (N_28063,N_27968,N_27831);
or U28064 (N_28064,N_27931,N_27952);
xnor U28065 (N_28065,N_27764,N_27887);
xnor U28066 (N_28066,N_27827,N_27978);
nor U28067 (N_28067,N_27779,N_27941);
and U28068 (N_28068,N_27774,N_27787);
nor U28069 (N_28069,N_27918,N_27915);
or U28070 (N_28070,N_27780,N_27997);
nand U28071 (N_28071,N_27829,N_27947);
or U28072 (N_28072,N_27999,N_27810);
and U28073 (N_28073,N_27914,N_27921);
nor U28074 (N_28074,N_27930,N_27944);
xnor U28075 (N_28075,N_27935,N_27843);
nand U28076 (N_28076,N_27826,N_27806);
and U28077 (N_28077,N_27979,N_27907);
nand U28078 (N_28078,N_27825,N_27789);
and U28079 (N_28079,N_27751,N_27855);
nand U28080 (N_28080,N_27828,N_27901);
nand U28081 (N_28081,N_27757,N_27891);
xnor U28082 (N_28082,N_27923,N_27772);
xnor U28083 (N_28083,N_27862,N_27924);
nor U28084 (N_28084,N_27819,N_27752);
nand U28085 (N_28085,N_27884,N_27989);
or U28086 (N_28086,N_27909,N_27942);
nand U28087 (N_28087,N_27956,N_27790);
nand U28088 (N_28088,N_27770,N_27786);
or U28089 (N_28089,N_27872,N_27836);
nand U28090 (N_28090,N_27998,N_27857);
nor U28091 (N_28091,N_27984,N_27856);
nor U28092 (N_28092,N_27945,N_27800);
or U28093 (N_28093,N_27818,N_27892);
or U28094 (N_28094,N_27845,N_27959);
nor U28095 (N_28095,N_27814,N_27796);
and U28096 (N_28096,N_27880,N_27928);
nand U28097 (N_28097,N_27983,N_27937);
or U28098 (N_28098,N_27970,N_27893);
nor U28099 (N_28099,N_27910,N_27960);
nor U28100 (N_28100,N_27830,N_27962);
and U28101 (N_28101,N_27966,N_27933);
nand U28102 (N_28102,N_27949,N_27853);
and U28103 (N_28103,N_27899,N_27807);
and U28104 (N_28104,N_27994,N_27974);
xor U28105 (N_28105,N_27816,N_27794);
xor U28106 (N_28106,N_27768,N_27927);
xnor U28107 (N_28107,N_27851,N_27936);
xnor U28108 (N_28108,N_27964,N_27896);
nor U28109 (N_28109,N_27852,N_27791);
nand U28110 (N_28110,N_27993,N_27846);
nand U28111 (N_28111,N_27967,N_27932);
nand U28112 (N_28112,N_27750,N_27817);
xnor U28113 (N_28113,N_27950,N_27902);
and U28114 (N_28114,N_27784,N_27973);
nand U28115 (N_28115,N_27982,N_27881);
nand U28116 (N_28116,N_27897,N_27890);
or U28117 (N_28117,N_27840,N_27939);
nand U28118 (N_28118,N_27972,N_27988);
nand U28119 (N_28119,N_27834,N_27797);
nand U28120 (N_28120,N_27833,N_27859);
nor U28121 (N_28121,N_27888,N_27758);
nor U28122 (N_28122,N_27940,N_27975);
or U28123 (N_28123,N_27813,N_27763);
or U28124 (N_28124,N_27823,N_27788);
xnor U28125 (N_28125,N_27876,N_27863);
xnor U28126 (N_28126,N_27835,N_27765);
nand U28127 (N_28127,N_27963,N_27847);
or U28128 (N_28128,N_27977,N_27755);
xor U28129 (N_28129,N_27750,N_27940);
xor U28130 (N_28130,N_27957,N_27806);
xor U28131 (N_28131,N_27866,N_27966);
xor U28132 (N_28132,N_27907,N_27798);
xor U28133 (N_28133,N_27985,N_27954);
and U28134 (N_28134,N_27992,N_27807);
nand U28135 (N_28135,N_27877,N_27871);
nor U28136 (N_28136,N_27807,N_27876);
xor U28137 (N_28137,N_27754,N_27991);
nand U28138 (N_28138,N_27766,N_27830);
nor U28139 (N_28139,N_27894,N_27873);
nand U28140 (N_28140,N_27946,N_27848);
xnor U28141 (N_28141,N_27768,N_27846);
xor U28142 (N_28142,N_27995,N_27846);
xnor U28143 (N_28143,N_27926,N_27833);
or U28144 (N_28144,N_27870,N_27949);
and U28145 (N_28145,N_27959,N_27905);
or U28146 (N_28146,N_27882,N_27931);
nor U28147 (N_28147,N_27982,N_27779);
xnor U28148 (N_28148,N_27800,N_27805);
or U28149 (N_28149,N_27802,N_27852);
or U28150 (N_28150,N_27977,N_27807);
nor U28151 (N_28151,N_27881,N_27802);
nand U28152 (N_28152,N_27888,N_27919);
nand U28153 (N_28153,N_27960,N_27928);
xnor U28154 (N_28154,N_27841,N_27852);
or U28155 (N_28155,N_27840,N_27999);
xor U28156 (N_28156,N_27991,N_27802);
and U28157 (N_28157,N_27804,N_27993);
or U28158 (N_28158,N_27798,N_27772);
xnor U28159 (N_28159,N_27913,N_27910);
nor U28160 (N_28160,N_27760,N_27948);
nand U28161 (N_28161,N_27940,N_27878);
nand U28162 (N_28162,N_27891,N_27814);
nor U28163 (N_28163,N_27872,N_27775);
or U28164 (N_28164,N_27772,N_27941);
nor U28165 (N_28165,N_27847,N_27762);
and U28166 (N_28166,N_27838,N_27775);
xnor U28167 (N_28167,N_27750,N_27834);
nor U28168 (N_28168,N_27995,N_27919);
and U28169 (N_28169,N_27899,N_27772);
nor U28170 (N_28170,N_27808,N_27951);
and U28171 (N_28171,N_27995,N_27900);
nor U28172 (N_28172,N_27891,N_27878);
xor U28173 (N_28173,N_27831,N_27902);
nand U28174 (N_28174,N_27807,N_27820);
nor U28175 (N_28175,N_27883,N_27777);
nand U28176 (N_28176,N_27855,N_27838);
xor U28177 (N_28177,N_27998,N_27929);
and U28178 (N_28178,N_27927,N_27929);
nand U28179 (N_28179,N_27783,N_27946);
and U28180 (N_28180,N_27820,N_27979);
xnor U28181 (N_28181,N_27853,N_27977);
nand U28182 (N_28182,N_27844,N_27966);
xnor U28183 (N_28183,N_27919,N_27952);
and U28184 (N_28184,N_27979,N_27879);
nor U28185 (N_28185,N_27964,N_27961);
nor U28186 (N_28186,N_27895,N_27833);
and U28187 (N_28187,N_27976,N_27808);
or U28188 (N_28188,N_27994,N_27864);
and U28189 (N_28189,N_27788,N_27751);
xor U28190 (N_28190,N_27751,N_27818);
nand U28191 (N_28191,N_27761,N_27846);
and U28192 (N_28192,N_27982,N_27937);
or U28193 (N_28193,N_27776,N_27854);
or U28194 (N_28194,N_27901,N_27802);
nand U28195 (N_28195,N_27906,N_27954);
xnor U28196 (N_28196,N_27862,N_27975);
nor U28197 (N_28197,N_27839,N_27760);
nand U28198 (N_28198,N_27862,N_27928);
nor U28199 (N_28199,N_27922,N_27777);
or U28200 (N_28200,N_27818,N_27788);
nor U28201 (N_28201,N_27792,N_27906);
nor U28202 (N_28202,N_27786,N_27829);
nor U28203 (N_28203,N_27929,N_27883);
and U28204 (N_28204,N_27768,N_27849);
nor U28205 (N_28205,N_27959,N_27807);
and U28206 (N_28206,N_27958,N_27837);
xor U28207 (N_28207,N_27879,N_27850);
and U28208 (N_28208,N_27914,N_27845);
and U28209 (N_28209,N_27815,N_27857);
xor U28210 (N_28210,N_27854,N_27761);
nand U28211 (N_28211,N_27827,N_27800);
xor U28212 (N_28212,N_27801,N_27907);
xnor U28213 (N_28213,N_27770,N_27972);
xor U28214 (N_28214,N_27999,N_27969);
and U28215 (N_28215,N_27994,N_27913);
nor U28216 (N_28216,N_27894,N_27751);
nor U28217 (N_28217,N_27883,N_27795);
nor U28218 (N_28218,N_27775,N_27777);
and U28219 (N_28219,N_27998,N_27997);
and U28220 (N_28220,N_27936,N_27811);
nand U28221 (N_28221,N_27940,N_27876);
xnor U28222 (N_28222,N_27752,N_27942);
nor U28223 (N_28223,N_27947,N_27923);
xnor U28224 (N_28224,N_27981,N_27991);
nand U28225 (N_28225,N_27777,N_27991);
xor U28226 (N_28226,N_27871,N_27777);
and U28227 (N_28227,N_27938,N_27882);
nor U28228 (N_28228,N_27830,N_27814);
and U28229 (N_28229,N_27772,N_27992);
nand U28230 (N_28230,N_27756,N_27978);
and U28231 (N_28231,N_27885,N_27839);
nor U28232 (N_28232,N_27872,N_27924);
xor U28233 (N_28233,N_27811,N_27837);
nand U28234 (N_28234,N_27962,N_27908);
nand U28235 (N_28235,N_27825,N_27978);
and U28236 (N_28236,N_27779,N_27957);
xnor U28237 (N_28237,N_27786,N_27934);
nor U28238 (N_28238,N_27891,N_27822);
xnor U28239 (N_28239,N_27838,N_27985);
nor U28240 (N_28240,N_27864,N_27981);
and U28241 (N_28241,N_27888,N_27764);
or U28242 (N_28242,N_27899,N_27808);
and U28243 (N_28243,N_27845,N_27968);
and U28244 (N_28244,N_27782,N_27891);
or U28245 (N_28245,N_27881,N_27823);
nand U28246 (N_28246,N_27855,N_27933);
or U28247 (N_28247,N_27955,N_27820);
nand U28248 (N_28248,N_27944,N_27910);
and U28249 (N_28249,N_27850,N_27836);
or U28250 (N_28250,N_28071,N_28088);
xor U28251 (N_28251,N_28093,N_28214);
nand U28252 (N_28252,N_28042,N_28145);
nand U28253 (N_28253,N_28232,N_28035);
nand U28254 (N_28254,N_28245,N_28208);
or U28255 (N_28255,N_28036,N_28159);
nand U28256 (N_28256,N_28120,N_28113);
or U28257 (N_28257,N_28015,N_28069);
and U28258 (N_28258,N_28164,N_28112);
xnor U28259 (N_28259,N_28106,N_28174);
xor U28260 (N_28260,N_28024,N_28139);
and U28261 (N_28261,N_28092,N_28194);
and U28262 (N_28262,N_28163,N_28017);
nand U28263 (N_28263,N_28222,N_28175);
nand U28264 (N_28264,N_28100,N_28207);
nand U28265 (N_28265,N_28212,N_28215);
or U28266 (N_28266,N_28022,N_28138);
nand U28267 (N_28267,N_28012,N_28249);
xnor U28268 (N_28268,N_28157,N_28204);
xnor U28269 (N_28269,N_28156,N_28028);
and U28270 (N_28270,N_28160,N_28054);
xnor U28271 (N_28271,N_28005,N_28130);
xnor U28272 (N_28272,N_28090,N_28030);
and U28273 (N_28273,N_28121,N_28099);
xor U28274 (N_28274,N_28228,N_28189);
nand U28275 (N_28275,N_28116,N_28230);
nor U28276 (N_28276,N_28183,N_28074);
or U28277 (N_28277,N_28011,N_28129);
xor U28278 (N_28278,N_28198,N_28199);
or U28279 (N_28279,N_28006,N_28033);
nor U28280 (N_28280,N_28000,N_28131);
nand U28281 (N_28281,N_28067,N_28010);
xor U28282 (N_28282,N_28196,N_28191);
nor U28283 (N_28283,N_28007,N_28047);
xor U28284 (N_28284,N_28097,N_28150);
xnor U28285 (N_28285,N_28085,N_28234);
or U28286 (N_28286,N_28083,N_28173);
or U28287 (N_28287,N_28117,N_28142);
nor U28288 (N_28288,N_28152,N_28066);
and U28289 (N_28289,N_28029,N_28125);
xor U28290 (N_28290,N_28225,N_28124);
and U28291 (N_28291,N_28154,N_28013);
and U28292 (N_28292,N_28072,N_28107);
or U28293 (N_28293,N_28170,N_28110);
and U28294 (N_28294,N_28244,N_28200);
or U28295 (N_28295,N_28240,N_28084);
nor U28296 (N_28296,N_28119,N_28050);
nand U28297 (N_28297,N_28102,N_28052);
nor U28298 (N_28298,N_28178,N_28239);
nand U28299 (N_28299,N_28027,N_28082);
nor U28300 (N_28300,N_28111,N_28123);
nor U28301 (N_28301,N_28053,N_28096);
xnor U28302 (N_28302,N_28179,N_28197);
and U28303 (N_28303,N_28018,N_28076);
nand U28304 (N_28304,N_28115,N_28192);
nor U28305 (N_28305,N_28026,N_28143);
nor U28306 (N_28306,N_28235,N_28188);
xnor U28307 (N_28307,N_28118,N_28002);
xor U28308 (N_28308,N_28168,N_28187);
or U28309 (N_28309,N_28141,N_28056);
and U28310 (N_28310,N_28216,N_28146);
nor U28311 (N_28311,N_28081,N_28248);
nand U28312 (N_28312,N_28064,N_28004);
or U28313 (N_28313,N_28247,N_28209);
or U28314 (N_28314,N_28223,N_28122);
nor U28315 (N_28315,N_28098,N_28180);
and U28316 (N_28316,N_28014,N_28190);
and U28317 (N_28317,N_28137,N_28077);
nand U28318 (N_28318,N_28109,N_28016);
or U28319 (N_28319,N_28233,N_28186);
nor U28320 (N_28320,N_28038,N_28044);
nor U28321 (N_28321,N_28039,N_28057);
and U28322 (N_28322,N_28095,N_28201);
xnor U28323 (N_28323,N_28217,N_28060);
or U28324 (N_28324,N_28227,N_28151);
nand U28325 (N_28325,N_28242,N_28003);
or U28326 (N_28326,N_28158,N_28087);
and U28327 (N_28327,N_28032,N_28127);
nand U28328 (N_28328,N_28231,N_28086);
and U28329 (N_28329,N_28103,N_28134);
nor U28330 (N_28330,N_28051,N_28034);
or U28331 (N_28331,N_28246,N_28148);
nand U28332 (N_28332,N_28155,N_28021);
nand U28333 (N_28333,N_28105,N_28220);
nand U28334 (N_28334,N_28009,N_28226);
xor U28335 (N_28335,N_28031,N_28205);
nand U28336 (N_28336,N_28065,N_28055);
and U28337 (N_28337,N_28177,N_28101);
or U28338 (N_28338,N_28075,N_28020);
xor U28339 (N_28339,N_28073,N_28237);
and U28340 (N_28340,N_28147,N_28079);
and U28341 (N_28341,N_28135,N_28162);
xnor U28342 (N_28342,N_28062,N_28008);
or U28343 (N_28343,N_28238,N_28213);
nand U28344 (N_28344,N_28241,N_28211);
nand U28345 (N_28345,N_28144,N_28126);
nand U28346 (N_28346,N_28149,N_28059);
and U28347 (N_28347,N_28061,N_28019);
nand U28348 (N_28348,N_28172,N_28063);
xor U28349 (N_28349,N_28219,N_28182);
nand U28350 (N_28350,N_28045,N_28195);
nand U28351 (N_28351,N_28133,N_28136);
and U28352 (N_28352,N_28025,N_28202);
and U28353 (N_28353,N_28167,N_28001);
nand U28354 (N_28354,N_28132,N_28037);
xor U28355 (N_28355,N_28108,N_28140);
and U28356 (N_28356,N_28070,N_28193);
and U28357 (N_28357,N_28184,N_28224);
nand U28358 (N_28358,N_28210,N_28041);
and U28359 (N_28359,N_28040,N_28229);
nand U28360 (N_28360,N_28068,N_28218);
and U28361 (N_28361,N_28048,N_28089);
xor U28362 (N_28362,N_28080,N_28058);
nand U28363 (N_28363,N_28161,N_28114);
xor U28364 (N_28364,N_28078,N_28049);
and U28365 (N_28365,N_28091,N_28243);
nor U28366 (N_28366,N_28236,N_28169);
and U28367 (N_28367,N_28104,N_28043);
or U28368 (N_28368,N_28185,N_28181);
nor U28369 (N_28369,N_28203,N_28046);
nand U28370 (N_28370,N_28171,N_28166);
xor U28371 (N_28371,N_28221,N_28176);
nand U28372 (N_28372,N_28153,N_28128);
or U28373 (N_28373,N_28023,N_28206);
and U28374 (N_28374,N_28094,N_28165);
or U28375 (N_28375,N_28128,N_28046);
nor U28376 (N_28376,N_28040,N_28177);
or U28377 (N_28377,N_28175,N_28141);
nor U28378 (N_28378,N_28034,N_28018);
nor U28379 (N_28379,N_28002,N_28069);
or U28380 (N_28380,N_28164,N_28075);
xor U28381 (N_28381,N_28140,N_28127);
xor U28382 (N_28382,N_28042,N_28196);
or U28383 (N_28383,N_28178,N_28154);
nand U28384 (N_28384,N_28098,N_28038);
and U28385 (N_28385,N_28016,N_28183);
nor U28386 (N_28386,N_28114,N_28019);
nor U28387 (N_28387,N_28070,N_28191);
and U28388 (N_28388,N_28102,N_28065);
xnor U28389 (N_28389,N_28218,N_28129);
xnor U28390 (N_28390,N_28142,N_28226);
nand U28391 (N_28391,N_28203,N_28134);
nor U28392 (N_28392,N_28128,N_28129);
or U28393 (N_28393,N_28102,N_28186);
and U28394 (N_28394,N_28138,N_28037);
xor U28395 (N_28395,N_28162,N_28140);
nand U28396 (N_28396,N_28166,N_28229);
or U28397 (N_28397,N_28169,N_28011);
nand U28398 (N_28398,N_28134,N_28008);
and U28399 (N_28399,N_28200,N_28224);
nor U28400 (N_28400,N_28107,N_28148);
and U28401 (N_28401,N_28029,N_28247);
and U28402 (N_28402,N_28077,N_28060);
nand U28403 (N_28403,N_28202,N_28094);
or U28404 (N_28404,N_28012,N_28076);
xnor U28405 (N_28405,N_28215,N_28099);
and U28406 (N_28406,N_28177,N_28082);
nor U28407 (N_28407,N_28014,N_28049);
and U28408 (N_28408,N_28218,N_28111);
nand U28409 (N_28409,N_28020,N_28077);
nor U28410 (N_28410,N_28041,N_28185);
and U28411 (N_28411,N_28182,N_28102);
xnor U28412 (N_28412,N_28034,N_28160);
or U28413 (N_28413,N_28004,N_28180);
and U28414 (N_28414,N_28201,N_28081);
and U28415 (N_28415,N_28154,N_28242);
xor U28416 (N_28416,N_28059,N_28196);
nor U28417 (N_28417,N_28171,N_28056);
nand U28418 (N_28418,N_28059,N_28028);
and U28419 (N_28419,N_28099,N_28069);
nor U28420 (N_28420,N_28162,N_28239);
xor U28421 (N_28421,N_28020,N_28013);
or U28422 (N_28422,N_28006,N_28009);
xor U28423 (N_28423,N_28118,N_28235);
nor U28424 (N_28424,N_28245,N_28235);
and U28425 (N_28425,N_28169,N_28141);
xor U28426 (N_28426,N_28121,N_28192);
nor U28427 (N_28427,N_28219,N_28068);
or U28428 (N_28428,N_28211,N_28145);
xor U28429 (N_28429,N_28017,N_28050);
or U28430 (N_28430,N_28079,N_28140);
nand U28431 (N_28431,N_28117,N_28141);
nor U28432 (N_28432,N_28212,N_28018);
or U28433 (N_28433,N_28019,N_28085);
nand U28434 (N_28434,N_28208,N_28114);
nor U28435 (N_28435,N_28126,N_28111);
xor U28436 (N_28436,N_28128,N_28214);
nor U28437 (N_28437,N_28239,N_28047);
nand U28438 (N_28438,N_28000,N_28087);
and U28439 (N_28439,N_28231,N_28112);
and U28440 (N_28440,N_28129,N_28050);
or U28441 (N_28441,N_28189,N_28191);
and U28442 (N_28442,N_28158,N_28137);
and U28443 (N_28443,N_28199,N_28057);
xnor U28444 (N_28444,N_28027,N_28050);
and U28445 (N_28445,N_28150,N_28109);
xnor U28446 (N_28446,N_28114,N_28180);
xnor U28447 (N_28447,N_28050,N_28137);
xor U28448 (N_28448,N_28161,N_28179);
and U28449 (N_28449,N_28106,N_28217);
or U28450 (N_28450,N_28240,N_28038);
xor U28451 (N_28451,N_28146,N_28075);
nand U28452 (N_28452,N_28185,N_28053);
and U28453 (N_28453,N_28023,N_28027);
nor U28454 (N_28454,N_28060,N_28071);
or U28455 (N_28455,N_28213,N_28247);
xor U28456 (N_28456,N_28243,N_28174);
nor U28457 (N_28457,N_28230,N_28104);
nor U28458 (N_28458,N_28041,N_28119);
nand U28459 (N_28459,N_28199,N_28077);
and U28460 (N_28460,N_28147,N_28135);
nand U28461 (N_28461,N_28192,N_28097);
nand U28462 (N_28462,N_28189,N_28186);
nor U28463 (N_28463,N_28017,N_28208);
nor U28464 (N_28464,N_28206,N_28123);
xnor U28465 (N_28465,N_28234,N_28018);
nor U28466 (N_28466,N_28141,N_28150);
xnor U28467 (N_28467,N_28108,N_28066);
nand U28468 (N_28468,N_28131,N_28033);
or U28469 (N_28469,N_28244,N_28080);
xnor U28470 (N_28470,N_28217,N_28130);
nor U28471 (N_28471,N_28245,N_28108);
or U28472 (N_28472,N_28190,N_28057);
nor U28473 (N_28473,N_28134,N_28080);
xnor U28474 (N_28474,N_28208,N_28053);
or U28475 (N_28475,N_28210,N_28181);
and U28476 (N_28476,N_28075,N_28002);
and U28477 (N_28477,N_28002,N_28207);
and U28478 (N_28478,N_28129,N_28235);
and U28479 (N_28479,N_28062,N_28073);
or U28480 (N_28480,N_28213,N_28242);
and U28481 (N_28481,N_28164,N_28152);
xor U28482 (N_28482,N_28194,N_28085);
xnor U28483 (N_28483,N_28206,N_28139);
and U28484 (N_28484,N_28139,N_28052);
or U28485 (N_28485,N_28162,N_28213);
or U28486 (N_28486,N_28007,N_28068);
and U28487 (N_28487,N_28182,N_28065);
or U28488 (N_28488,N_28239,N_28130);
xor U28489 (N_28489,N_28059,N_28092);
xor U28490 (N_28490,N_28141,N_28116);
xor U28491 (N_28491,N_28016,N_28205);
xnor U28492 (N_28492,N_28187,N_28238);
xor U28493 (N_28493,N_28003,N_28109);
or U28494 (N_28494,N_28215,N_28114);
or U28495 (N_28495,N_28216,N_28125);
xnor U28496 (N_28496,N_28191,N_28037);
nand U28497 (N_28497,N_28004,N_28143);
nor U28498 (N_28498,N_28166,N_28055);
and U28499 (N_28499,N_28170,N_28126);
nand U28500 (N_28500,N_28455,N_28283);
nor U28501 (N_28501,N_28297,N_28382);
and U28502 (N_28502,N_28419,N_28452);
and U28503 (N_28503,N_28262,N_28369);
nand U28504 (N_28504,N_28290,N_28460);
nand U28505 (N_28505,N_28451,N_28476);
nand U28506 (N_28506,N_28380,N_28309);
nor U28507 (N_28507,N_28305,N_28315);
or U28508 (N_28508,N_28449,N_28335);
and U28509 (N_28509,N_28362,N_28420);
nor U28510 (N_28510,N_28474,N_28396);
or U28511 (N_28511,N_28450,N_28466);
xnor U28512 (N_28512,N_28308,N_28354);
and U28513 (N_28513,N_28388,N_28433);
nand U28514 (N_28514,N_28348,N_28372);
or U28515 (N_28515,N_28491,N_28307);
or U28516 (N_28516,N_28263,N_28379);
nand U28517 (N_28517,N_28469,N_28467);
nand U28518 (N_28518,N_28434,N_28255);
nor U28519 (N_28519,N_28316,N_28492);
nand U28520 (N_28520,N_28443,N_28355);
or U28521 (N_28521,N_28393,N_28327);
or U28522 (N_28522,N_28456,N_28293);
xnor U28523 (N_28523,N_28320,N_28282);
or U28524 (N_28524,N_28352,N_28321);
nand U28525 (N_28525,N_28442,N_28444);
and U28526 (N_28526,N_28257,N_28252);
nand U28527 (N_28527,N_28383,N_28483);
nor U28528 (N_28528,N_28295,N_28394);
nor U28529 (N_28529,N_28421,N_28468);
nor U28530 (N_28530,N_28366,N_28266);
nor U28531 (N_28531,N_28415,N_28399);
xnor U28532 (N_28532,N_28303,N_28325);
nand U28533 (N_28533,N_28448,N_28342);
nand U28534 (N_28534,N_28404,N_28428);
or U28535 (N_28535,N_28438,N_28497);
xor U28536 (N_28536,N_28277,N_28322);
nand U28537 (N_28537,N_28403,N_28299);
and U28538 (N_28538,N_28312,N_28251);
nor U28539 (N_28539,N_28405,N_28333);
nor U28540 (N_28540,N_28271,N_28464);
nor U28541 (N_28541,N_28408,N_28311);
or U28542 (N_28542,N_28427,N_28317);
or U28543 (N_28543,N_28367,N_28445);
xnor U28544 (N_28544,N_28389,N_28259);
nor U28545 (N_28545,N_28281,N_28381);
or U28546 (N_28546,N_28306,N_28331);
xnor U28547 (N_28547,N_28414,N_28267);
nor U28548 (N_28548,N_28323,N_28345);
nor U28549 (N_28549,N_28296,N_28356);
xor U28550 (N_28550,N_28498,N_28338);
and U28551 (N_28551,N_28470,N_28370);
or U28552 (N_28552,N_28477,N_28481);
nor U28553 (N_28553,N_28463,N_28276);
xnor U28554 (N_28554,N_28446,N_28407);
or U28555 (N_28555,N_28471,N_28482);
and U28556 (N_28556,N_28301,N_28360);
or U28557 (N_28557,N_28373,N_28353);
nor U28558 (N_28558,N_28254,N_28411);
or U28559 (N_28559,N_28268,N_28346);
and U28560 (N_28560,N_28472,N_28364);
xor U28561 (N_28561,N_28391,N_28269);
or U28562 (N_28562,N_28319,N_28258);
nor U28563 (N_28563,N_28478,N_28330);
nor U28564 (N_28564,N_28435,N_28494);
nand U28565 (N_28565,N_28358,N_28359);
nor U28566 (N_28566,N_28377,N_28289);
or U28567 (N_28567,N_28326,N_28270);
nand U28568 (N_28568,N_28375,N_28337);
nor U28569 (N_28569,N_28458,N_28264);
and U28570 (N_28570,N_28417,N_28291);
nand U28571 (N_28571,N_28300,N_28447);
or U28572 (N_28572,N_28298,N_28390);
nand U28573 (N_28573,N_28288,N_28284);
and U28574 (N_28574,N_28285,N_28378);
or U28575 (N_28575,N_28313,N_28437);
nand U28576 (N_28576,N_28343,N_28499);
nor U28577 (N_28577,N_28473,N_28441);
nand U28578 (N_28578,N_28336,N_28406);
or U28579 (N_28579,N_28328,N_28430);
or U28580 (N_28580,N_28489,N_28371);
nand U28581 (N_28581,N_28385,N_28416);
xor U28582 (N_28582,N_28485,N_28410);
nand U28583 (N_28583,N_28357,N_28459);
or U28584 (N_28584,N_28304,N_28397);
nor U28585 (N_28585,N_28302,N_28495);
or U28586 (N_28586,N_28487,N_28368);
nand U28587 (N_28587,N_28454,N_28344);
xor U28588 (N_28588,N_28387,N_28429);
nor U28589 (N_28589,N_28436,N_28425);
and U28590 (N_28590,N_28440,N_28350);
nor U28591 (N_28591,N_28386,N_28310);
and U28592 (N_28592,N_28324,N_28423);
or U28593 (N_28593,N_28361,N_28363);
xor U28594 (N_28594,N_28457,N_28418);
or U28595 (N_28595,N_28401,N_28493);
and U28596 (N_28596,N_28465,N_28490);
nor U28597 (N_28597,N_28484,N_28480);
nor U28598 (N_28598,N_28365,N_28496);
or U28599 (N_28599,N_28272,N_28265);
nor U28600 (N_28600,N_28432,N_28398);
nor U28601 (N_28601,N_28349,N_28256);
nor U28602 (N_28602,N_28341,N_28400);
and U28603 (N_28603,N_28424,N_28392);
nand U28604 (N_28604,N_28250,N_28253);
xnor U28605 (N_28605,N_28279,N_28332);
or U28606 (N_28606,N_28488,N_28340);
nand U28607 (N_28607,N_28413,N_28273);
nand U28608 (N_28608,N_28351,N_28347);
nor U28609 (N_28609,N_28461,N_28314);
or U28610 (N_28610,N_28339,N_28286);
and U28611 (N_28611,N_28395,N_28462);
nor U28612 (N_28612,N_28479,N_28261);
or U28613 (N_28613,N_28260,N_28334);
xor U28614 (N_28614,N_28475,N_28274);
and U28615 (N_28615,N_28278,N_28426);
or U28616 (N_28616,N_28384,N_28422);
nand U28617 (N_28617,N_28280,N_28294);
nor U28618 (N_28618,N_28287,N_28275);
or U28619 (N_28619,N_28409,N_28329);
nor U28620 (N_28620,N_28453,N_28439);
or U28621 (N_28621,N_28318,N_28376);
or U28622 (N_28622,N_28486,N_28402);
nor U28623 (N_28623,N_28374,N_28292);
or U28624 (N_28624,N_28431,N_28412);
nor U28625 (N_28625,N_28279,N_28408);
xor U28626 (N_28626,N_28408,N_28297);
xnor U28627 (N_28627,N_28276,N_28472);
nor U28628 (N_28628,N_28342,N_28389);
or U28629 (N_28629,N_28345,N_28258);
nand U28630 (N_28630,N_28450,N_28371);
or U28631 (N_28631,N_28436,N_28290);
xnor U28632 (N_28632,N_28260,N_28257);
and U28633 (N_28633,N_28403,N_28392);
or U28634 (N_28634,N_28405,N_28421);
nand U28635 (N_28635,N_28324,N_28357);
xor U28636 (N_28636,N_28285,N_28267);
nand U28637 (N_28637,N_28264,N_28251);
nand U28638 (N_28638,N_28331,N_28340);
or U28639 (N_28639,N_28313,N_28395);
and U28640 (N_28640,N_28386,N_28406);
nand U28641 (N_28641,N_28367,N_28355);
or U28642 (N_28642,N_28480,N_28387);
and U28643 (N_28643,N_28255,N_28327);
and U28644 (N_28644,N_28301,N_28424);
xnor U28645 (N_28645,N_28391,N_28366);
nor U28646 (N_28646,N_28337,N_28392);
xnor U28647 (N_28647,N_28490,N_28253);
nor U28648 (N_28648,N_28347,N_28405);
xnor U28649 (N_28649,N_28405,N_28263);
nand U28650 (N_28650,N_28281,N_28319);
and U28651 (N_28651,N_28255,N_28307);
nor U28652 (N_28652,N_28483,N_28449);
or U28653 (N_28653,N_28341,N_28312);
or U28654 (N_28654,N_28265,N_28315);
xnor U28655 (N_28655,N_28491,N_28313);
and U28656 (N_28656,N_28347,N_28337);
nor U28657 (N_28657,N_28375,N_28420);
nor U28658 (N_28658,N_28332,N_28436);
and U28659 (N_28659,N_28346,N_28392);
nor U28660 (N_28660,N_28438,N_28498);
xnor U28661 (N_28661,N_28261,N_28391);
or U28662 (N_28662,N_28428,N_28310);
xnor U28663 (N_28663,N_28302,N_28403);
and U28664 (N_28664,N_28397,N_28407);
nor U28665 (N_28665,N_28291,N_28468);
nor U28666 (N_28666,N_28271,N_28318);
nor U28667 (N_28667,N_28452,N_28322);
nor U28668 (N_28668,N_28336,N_28363);
and U28669 (N_28669,N_28300,N_28305);
xor U28670 (N_28670,N_28434,N_28410);
xor U28671 (N_28671,N_28330,N_28348);
nand U28672 (N_28672,N_28361,N_28473);
nand U28673 (N_28673,N_28362,N_28281);
or U28674 (N_28674,N_28340,N_28316);
or U28675 (N_28675,N_28427,N_28458);
and U28676 (N_28676,N_28499,N_28257);
nor U28677 (N_28677,N_28473,N_28391);
or U28678 (N_28678,N_28296,N_28417);
xor U28679 (N_28679,N_28340,N_28314);
or U28680 (N_28680,N_28382,N_28318);
nand U28681 (N_28681,N_28442,N_28443);
nand U28682 (N_28682,N_28395,N_28282);
xnor U28683 (N_28683,N_28404,N_28338);
xnor U28684 (N_28684,N_28427,N_28390);
or U28685 (N_28685,N_28414,N_28429);
or U28686 (N_28686,N_28331,N_28479);
or U28687 (N_28687,N_28427,N_28271);
or U28688 (N_28688,N_28445,N_28497);
or U28689 (N_28689,N_28344,N_28324);
nor U28690 (N_28690,N_28384,N_28255);
nor U28691 (N_28691,N_28262,N_28499);
xor U28692 (N_28692,N_28438,N_28266);
xnor U28693 (N_28693,N_28355,N_28470);
or U28694 (N_28694,N_28467,N_28350);
and U28695 (N_28695,N_28496,N_28297);
nand U28696 (N_28696,N_28499,N_28270);
and U28697 (N_28697,N_28284,N_28488);
and U28698 (N_28698,N_28423,N_28391);
xnor U28699 (N_28699,N_28308,N_28374);
and U28700 (N_28700,N_28440,N_28496);
and U28701 (N_28701,N_28463,N_28486);
or U28702 (N_28702,N_28339,N_28322);
nand U28703 (N_28703,N_28406,N_28333);
xor U28704 (N_28704,N_28461,N_28275);
and U28705 (N_28705,N_28253,N_28466);
and U28706 (N_28706,N_28362,N_28406);
and U28707 (N_28707,N_28448,N_28450);
nand U28708 (N_28708,N_28262,N_28272);
nand U28709 (N_28709,N_28413,N_28312);
or U28710 (N_28710,N_28289,N_28485);
nand U28711 (N_28711,N_28410,N_28404);
nand U28712 (N_28712,N_28391,N_28444);
nand U28713 (N_28713,N_28306,N_28404);
and U28714 (N_28714,N_28456,N_28323);
nor U28715 (N_28715,N_28463,N_28488);
and U28716 (N_28716,N_28470,N_28375);
or U28717 (N_28717,N_28499,N_28404);
or U28718 (N_28718,N_28300,N_28392);
xnor U28719 (N_28719,N_28251,N_28324);
and U28720 (N_28720,N_28351,N_28465);
nor U28721 (N_28721,N_28439,N_28403);
nor U28722 (N_28722,N_28484,N_28382);
and U28723 (N_28723,N_28383,N_28469);
or U28724 (N_28724,N_28353,N_28305);
and U28725 (N_28725,N_28334,N_28429);
nand U28726 (N_28726,N_28483,N_28277);
xnor U28727 (N_28727,N_28424,N_28450);
xnor U28728 (N_28728,N_28395,N_28487);
xor U28729 (N_28729,N_28285,N_28467);
or U28730 (N_28730,N_28484,N_28283);
nor U28731 (N_28731,N_28335,N_28478);
nand U28732 (N_28732,N_28312,N_28350);
xor U28733 (N_28733,N_28367,N_28276);
nor U28734 (N_28734,N_28368,N_28252);
and U28735 (N_28735,N_28459,N_28383);
and U28736 (N_28736,N_28374,N_28321);
nand U28737 (N_28737,N_28303,N_28496);
and U28738 (N_28738,N_28310,N_28455);
nor U28739 (N_28739,N_28412,N_28293);
and U28740 (N_28740,N_28444,N_28318);
nor U28741 (N_28741,N_28475,N_28303);
nor U28742 (N_28742,N_28340,N_28420);
nand U28743 (N_28743,N_28399,N_28312);
nor U28744 (N_28744,N_28290,N_28386);
or U28745 (N_28745,N_28296,N_28476);
nand U28746 (N_28746,N_28432,N_28385);
and U28747 (N_28747,N_28336,N_28347);
nor U28748 (N_28748,N_28279,N_28280);
or U28749 (N_28749,N_28320,N_28354);
xor U28750 (N_28750,N_28611,N_28747);
xor U28751 (N_28751,N_28679,N_28659);
xnor U28752 (N_28752,N_28690,N_28535);
nor U28753 (N_28753,N_28614,N_28503);
and U28754 (N_28754,N_28525,N_28632);
and U28755 (N_28755,N_28568,N_28579);
xnor U28756 (N_28756,N_28674,N_28662);
and U28757 (N_28757,N_28732,N_28695);
or U28758 (N_28758,N_28528,N_28671);
and U28759 (N_28759,N_28650,N_28652);
or U28760 (N_28760,N_28546,N_28653);
xnor U28761 (N_28761,N_28642,N_28615);
and U28762 (N_28762,N_28543,N_28541);
nand U28763 (N_28763,N_28501,N_28622);
nor U28764 (N_28764,N_28573,N_28569);
or U28765 (N_28765,N_28624,N_28700);
and U28766 (N_28766,N_28547,N_28713);
nand U28767 (N_28767,N_28514,N_28635);
and U28768 (N_28768,N_28585,N_28716);
xor U28769 (N_28769,N_28548,N_28656);
nor U28770 (N_28770,N_28647,N_28651);
xnor U28771 (N_28771,N_28540,N_28565);
nor U28772 (N_28772,N_28698,N_28749);
and U28773 (N_28773,N_28575,N_28502);
and U28774 (N_28774,N_28578,N_28684);
or U28775 (N_28775,N_28744,N_28726);
nor U28776 (N_28776,N_28699,N_28688);
nor U28777 (N_28777,N_28741,N_28572);
and U28778 (N_28778,N_28566,N_28554);
nand U28779 (N_28779,N_28739,N_28550);
or U28780 (N_28780,N_28517,N_28666);
xor U28781 (N_28781,N_28717,N_28734);
and U28782 (N_28782,N_28567,N_28587);
and U28783 (N_28783,N_28733,N_28509);
nand U28784 (N_28784,N_28508,N_28602);
nor U28785 (N_28785,N_28746,N_28522);
and U28786 (N_28786,N_28560,N_28696);
or U28787 (N_28787,N_28603,N_28743);
nor U28788 (N_28788,N_28715,N_28636);
xnor U28789 (N_28789,N_28702,N_28516);
nor U28790 (N_28790,N_28559,N_28592);
xnor U28791 (N_28791,N_28580,N_28604);
and U28792 (N_28792,N_28708,N_28504);
xor U28793 (N_28793,N_28675,N_28710);
nand U28794 (N_28794,N_28551,N_28505);
and U28795 (N_28795,N_28660,N_28655);
or U28796 (N_28796,N_28731,N_28694);
and U28797 (N_28797,N_28558,N_28544);
or U28798 (N_28798,N_28513,N_28676);
nor U28799 (N_28799,N_28685,N_28610);
nand U28800 (N_28800,N_28521,N_28707);
nand U28801 (N_28801,N_28595,N_28616);
nand U28802 (N_28802,N_28657,N_28553);
and U28803 (N_28803,N_28582,N_28623);
nor U28804 (N_28804,N_28654,N_28518);
nand U28805 (N_28805,N_28649,N_28721);
or U28806 (N_28806,N_28570,N_28748);
or U28807 (N_28807,N_28594,N_28539);
nor U28808 (N_28808,N_28545,N_28712);
nor U28809 (N_28809,N_28735,N_28637);
xor U28810 (N_28810,N_28745,N_28533);
nand U28811 (N_28811,N_28672,N_28641);
and U28812 (N_28812,N_28630,N_28658);
nor U28813 (N_28813,N_28725,N_28620);
nand U28814 (N_28814,N_28597,N_28683);
or U28815 (N_28815,N_28571,N_28625);
or U28816 (N_28816,N_28538,N_28738);
and U28817 (N_28817,N_28621,N_28507);
xnor U28818 (N_28818,N_28520,N_28556);
or U28819 (N_28819,N_28686,N_28629);
and U28820 (N_28820,N_28704,N_28612);
xnor U28821 (N_28821,N_28606,N_28718);
or U28822 (N_28822,N_28697,N_28643);
xnor U28823 (N_28823,N_28607,N_28574);
or U28824 (N_28824,N_28729,N_28730);
or U28825 (N_28825,N_28628,N_28723);
nor U28826 (N_28826,N_28561,N_28682);
and U28827 (N_28827,N_28542,N_28705);
xor U28828 (N_28828,N_28589,N_28737);
xor U28829 (N_28829,N_28681,N_28633);
nand U28830 (N_28830,N_28691,N_28687);
xor U28831 (N_28831,N_28709,N_28706);
xnor U28832 (N_28832,N_28524,N_28663);
or U28833 (N_28833,N_28583,N_28667);
nand U28834 (N_28834,N_28586,N_28605);
nor U28835 (N_28835,N_28669,N_28665);
or U28836 (N_28836,N_28711,N_28529);
nor U28837 (N_28837,N_28512,N_28719);
xor U28838 (N_28838,N_28626,N_28506);
and U28839 (N_28839,N_28673,N_28500);
xor U28840 (N_28840,N_28639,N_28515);
nand U28841 (N_28841,N_28564,N_28678);
nor U28842 (N_28842,N_28530,N_28645);
nor U28843 (N_28843,N_28634,N_28536);
and U28844 (N_28844,N_28692,N_28549);
xnor U28845 (N_28845,N_28596,N_28562);
xor U28846 (N_28846,N_28617,N_28511);
and U28847 (N_28847,N_28740,N_28640);
or U28848 (N_28848,N_28555,N_28584);
or U28849 (N_28849,N_28526,N_28689);
or U28850 (N_28850,N_28576,N_28661);
and U28851 (N_28851,N_28598,N_28720);
nand U28852 (N_28852,N_28613,N_28618);
nand U28853 (N_28853,N_28519,N_28646);
nor U28854 (N_28854,N_28631,N_28527);
and U28855 (N_28855,N_28677,N_28644);
and U28856 (N_28856,N_28563,N_28608);
and U28857 (N_28857,N_28670,N_28742);
or U28858 (N_28858,N_28600,N_28588);
and U28859 (N_28859,N_28590,N_28664);
xor U28860 (N_28860,N_28693,N_28627);
and U28861 (N_28861,N_28680,N_28727);
and U28862 (N_28862,N_28619,N_28534);
nand U28863 (N_28863,N_28532,N_28736);
and U28864 (N_28864,N_28510,N_28728);
or U28865 (N_28865,N_28591,N_28609);
xnor U28866 (N_28866,N_28701,N_28577);
xnor U28867 (N_28867,N_28714,N_28557);
nand U28868 (N_28868,N_28648,N_28668);
xor U28869 (N_28869,N_28537,N_28581);
nand U28870 (N_28870,N_28724,N_28703);
xnor U28871 (N_28871,N_28552,N_28523);
nor U28872 (N_28872,N_28593,N_28531);
and U28873 (N_28873,N_28722,N_28601);
nand U28874 (N_28874,N_28599,N_28638);
nand U28875 (N_28875,N_28743,N_28529);
xnor U28876 (N_28876,N_28635,N_28563);
xnor U28877 (N_28877,N_28512,N_28657);
nand U28878 (N_28878,N_28621,N_28672);
xnor U28879 (N_28879,N_28656,N_28593);
or U28880 (N_28880,N_28727,N_28632);
and U28881 (N_28881,N_28746,N_28564);
and U28882 (N_28882,N_28697,N_28626);
nor U28883 (N_28883,N_28739,N_28573);
and U28884 (N_28884,N_28744,N_28749);
nor U28885 (N_28885,N_28612,N_28665);
xor U28886 (N_28886,N_28551,N_28523);
or U28887 (N_28887,N_28566,N_28532);
xor U28888 (N_28888,N_28692,N_28749);
xor U28889 (N_28889,N_28695,N_28548);
or U28890 (N_28890,N_28701,N_28632);
nand U28891 (N_28891,N_28723,N_28726);
nor U28892 (N_28892,N_28523,N_28605);
and U28893 (N_28893,N_28726,N_28646);
and U28894 (N_28894,N_28656,N_28644);
and U28895 (N_28895,N_28747,N_28635);
nand U28896 (N_28896,N_28696,N_28622);
and U28897 (N_28897,N_28541,N_28655);
and U28898 (N_28898,N_28501,N_28713);
or U28899 (N_28899,N_28678,N_28616);
and U28900 (N_28900,N_28626,N_28551);
and U28901 (N_28901,N_28728,N_28651);
or U28902 (N_28902,N_28617,N_28720);
or U28903 (N_28903,N_28540,N_28544);
nor U28904 (N_28904,N_28599,N_28701);
nand U28905 (N_28905,N_28599,N_28580);
nor U28906 (N_28906,N_28676,N_28560);
or U28907 (N_28907,N_28721,N_28586);
nand U28908 (N_28908,N_28643,N_28738);
or U28909 (N_28909,N_28729,N_28601);
xor U28910 (N_28910,N_28500,N_28708);
xnor U28911 (N_28911,N_28622,N_28565);
nand U28912 (N_28912,N_28627,N_28520);
and U28913 (N_28913,N_28550,N_28729);
and U28914 (N_28914,N_28543,N_28700);
xnor U28915 (N_28915,N_28558,N_28679);
or U28916 (N_28916,N_28734,N_28703);
nand U28917 (N_28917,N_28647,N_28583);
and U28918 (N_28918,N_28741,N_28679);
xnor U28919 (N_28919,N_28523,N_28596);
nor U28920 (N_28920,N_28726,N_28684);
xor U28921 (N_28921,N_28526,N_28648);
xnor U28922 (N_28922,N_28631,N_28660);
nand U28923 (N_28923,N_28514,N_28734);
and U28924 (N_28924,N_28727,N_28732);
or U28925 (N_28925,N_28540,N_28555);
nand U28926 (N_28926,N_28710,N_28708);
and U28927 (N_28927,N_28602,N_28655);
or U28928 (N_28928,N_28603,N_28654);
nand U28929 (N_28929,N_28728,N_28598);
and U28930 (N_28930,N_28583,N_28694);
and U28931 (N_28931,N_28726,N_28683);
and U28932 (N_28932,N_28524,N_28604);
or U28933 (N_28933,N_28749,N_28515);
and U28934 (N_28934,N_28743,N_28730);
nor U28935 (N_28935,N_28593,N_28740);
nand U28936 (N_28936,N_28663,N_28727);
xnor U28937 (N_28937,N_28584,N_28683);
or U28938 (N_28938,N_28636,N_28669);
or U28939 (N_28939,N_28518,N_28715);
or U28940 (N_28940,N_28710,N_28539);
nor U28941 (N_28941,N_28502,N_28699);
nand U28942 (N_28942,N_28668,N_28540);
and U28943 (N_28943,N_28610,N_28518);
and U28944 (N_28944,N_28508,N_28693);
nor U28945 (N_28945,N_28720,N_28632);
xor U28946 (N_28946,N_28733,N_28648);
xnor U28947 (N_28947,N_28542,N_28543);
xnor U28948 (N_28948,N_28694,N_28579);
and U28949 (N_28949,N_28676,N_28688);
and U28950 (N_28950,N_28710,N_28526);
nor U28951 (N_28951,N_28734,N_28674);
nand U28952 (N_28952,N_28596,N_28675);
or U28953 (N_28953,N_28617,N_28614);
xor U28954 (N_28954,N_28565,N_28730);
or U28955 (N_28955,N_28502,N_28516);
xor U28956 (N_28956,N_28567,N_28628);
and U28957 (N_28957,N_28601,N_28709);
or U28958 (N_28958,N_28535,N_28744);
or U28959 (N_28959,N_28695,N_28685);
and U28960 (N_28960,N_28501,N_28553);
and U28961 (N_28961,N_28574,N_28558);
xnor U28962 (N_28962,N_28593,N_28566);
xor U28963 (N_28963,N_28551,N_28620);
nor U28964 (N_28964,N_28691,N_28690);
nor U28965 (N_28965,N_28646,N_28745);
nand U28966 (N_28966,N_28667,N_28664);
xor U28967 (N_28967,N_28509,N_28653);
or U28968 (N_28968,N_28555,N_28628);
and U28969 (N_28969,N_28730,N_28594);
and U28970 (N_28970,N_28575,N_28580);
nand U28971 (N_28971,N_28542,N_28540);
and U28972 (N_28972,N_28734,N_28679);
nand U28973 (N_28973,N_28569,N_28547);
and U28974 (N_28974,N_28540,N_28593);
and U28975 (N_28975,N_28705,N_28515);
xnor U28976 (N_28976,N_28622,N_28720);
and U28977 (N_28977,N_28573,N_28678);
xor U28978 (N_28978,N_28742,N_28647);
or U28979 (N_28979,N_28694,N_28588);
nand U28980 (N_28980,N_28541,N_28698);
nand U28981 (N_28981,N_28612,N_28726);
and U28982 (N_28982,N_28717,N_28602);
and U28983 (N_28983,N_28543,N_28597);
xor U28984 (N_28984,N_28614,N_28622);
or U28985 (N_28985,N_28692,N_28545);
xor U28986 (N_28986,N_28685,N_28676);
nand U28987 (N_28987,N_28727,N_28533);
nand U28988 (N_28988,N_28695,N_28534);
or U28989 (N_28989,N_28504,N_28696);
nand U28990 (N_28990,N_28664,N_28678);
xnor U28991 (N_28991,N_28517,N_28552);
nand U28992 (N_28992,N_28690,N_28515);
and U28993 (N_28993,N_28610,N_28575);
nand U28994 (N_28994,N_28673,N_28619);
nand U28995 (N_28995,N_28631,N_28673);
nand U28996 (N_28996,N_28698,N_28613);
nand U28997 (N_28997,N_28548,N_28715);
and U28998 (N_28998,N_28718,N_28615);
nand U28999 (N_28999,N_28730,N_28745);
nand U29000 (N_29000,N_28936,N_28833);
or U29001 (N_29001,N_28951,N_28809);
and U29002 (N_29002,N_28861,N_28911);
nor U29003 (N_29003,N_28767,N_28890);
nand U29004 (N_29004,N_28779,N_28819);
or U29005 (N_29005,N_28942,N_28825);
nor U29006 (N_29006,N_28993,N_28888);
and U29007 (N_29007,N_28766,N_28863);
nand U29008 (N_29008,N_28789,N_28772);
and U29009 (N_29009,N_28816,N_28995);
xnor U29010 (N_29010,N_28929,N_28878);
nor U29011 (N_29011,N_28792,N_28797);
xor U29012 (N_29012,N_28967,N_28981);
or U29013 (N_29013,N_28832,N_28831);
nand U29014 (N_29014,N_28872,N_28877);
or U29015 (N_29015,N_28869,N_28912);
and U29016 (N_29016,N_28873,N_28791);
nand U29017 (N_29017,N_28774,N_28934);
or U29018 (N_29018,N_28979,N_28938);
nor U29019 (N_29019,N_28836,N_28773);
nor U29020 (N_29020,N_28879,N_28810);
or U29021 (N_29021,N_28870,N_28847);
nand U29022 (N_29022,N_28943,N_28959);
xnor U29023 (N_29023,N_28834,N_28788);
or U29024 (N_29024,N_28914,N_28953);
nor U29025 (N_29025,N_28957,N_28760);
or U29026 (N_29026,N_28970,N_28992);
nor U29027 (N_29027,N_28891,N_28762);
and U29028 (N_29028,N_28759,N_28867);
nand U29029 (N_29029,N_28826,N_28801);
nor U29030 (N_29030,N_28971,N_28996);
or U29031 (N_29031,N_28854,N_28848);
nor U29032 (N_29032,N_28906,N_28922);
nor U29033 (N_29033,N_28851,N_28786);
or U29034 (N_29034,N_28802,N_28865);
and U29035 (N_29035,N_28820,N_28884);
nand U29036 (N_29036,N_28923,N_28990);
or U29037 (N_29037,N_28883,N_28987);
nor U29038 (N_29038,N_28985,N_28780);
nand U29039 (N_29039,N_28966,N_28909);
nand U29040 (N_29040,N_28823,N_28986);
and U29041 (N_29041,N_28916,N_28806);
xor U29042 (N_29042,N_28905,N_28757);
or U29043 (N_29043,N_28962,N_28903);
nand U29044 (N_29044,N_28949,N_28900);
nand U29045 (N_29045,N_28928,N_28843);
and U29046 (N_29046,N_28895,N_28858);
nand U29047 (N_29047,N_28771,N_28965);
xnor U29048 (N_29048,N_28814,N_28755);
and U29049 (N_29049,N_28924,N_28796);
and U29050 (N_29050,N_28855,N_28963);
and U29051 (N_29051,N_28817,N_28874);
and U29052 (N_29052,N_28893,N_28940);
nand U29053 (N_29053,N_28783,N_28917);
nor U29054 (N_29054,N_28821,N_28840);
nand U29055 (N_29055,N_28787,N_28756);
and U29056 (N_29056,N_28980,N_28887);
xor U29057 (N_29057,N_28808,N_28844);
and U29058 (N_29058,N_28918,N_28952);
or U29059 (N_29059,N_28849,N_28857);
or U29060 (N_29060,N_28886,N_28902);
xnor U29061 (N_29061,N_28982,N_28950);
and U29062 (N_29062,N_28829,N_28919);
nor U29063 (N_29063,N_28750,N_28991);
and U29064 (N_29064,N_28958,N_28930);
or U29065 (N_29065,N_28835,N_28812);
nand U29066 (N_29066,N_28793,N_28860);
xor U29067 (N_29067,N_28856,N_28968);
and U29068 (N_29068,N_28811,N_28866);
and U29069 (N_29069,N_28846,N_28948);
nor U29070 (N_29070,N_28868,N_28853);
nor U29071 (N_29071,N_28818,N_28827);
xor U29072 (N_29072,N_28975,N_28815);
nand U29073 (N_29073,N_28947,N_28941);
nand U29074 (N_29074,N_28813,N_28778);
and U29075 (N_29075,N_28784,N_28897);
nand U29076 (N_29076,N_28775,N_28973);
or U29077 (N_29077,N_28910,N_28799);
nor U29078 (N_29078,N_28768,N_28794);
or U29079 (N_29079,N_28763,N_28998);
or U29080 (N_29080,N_28798,N_28881);
and U29081 (N_29081,N_28770,N_28978);
or U29082 (N_29082,N_28969,N_28976);
or U29083 (N_29083,N_28927,N_28790);
and U29084 (N_29084,N_28932,N_28901);
nand U29085 (N_29085,N_28805,N_28753);
xnor U29086 (N_29086,N_28871,N_28955);
or U29087 (N_29087,N_28935,N_28882);
nor U29088 (N_29088,N_28937,N_28830);
nand U29089 (N_29089,N_28841,N_28974);
and U29090 (N_29090,N_28837,N_28915);
nand U29091 (N_29091,N_28859,N_28754);
and U29092 (N_29092,N_28999,N_28781);
nor U29093 (N_29093,N_28988,N_28795);
xor U29094 (N_29094,N_28994,N_28758);
nand U29095 (N_29095,N_28752,N_28972);
or U29096 (N_29096,N_28907,N_28944);
xor U29097 (N_29097,N_28862,N_28761);
and U29098 (N_29098,N_28964,N_28769);
nand U29099 (N_29099,N_28997,N_28852);
nand U29100 (N_29100,N_28875,N_28961);
and U29101 (N_29101,N_28989,N_28984);
or U29102 (N_29102,N_28913,N_28785);
nand U29103 (N_29103,N_28977,N_28939);
or U29104 (N_29104,N_28800,N_28925);
nand U29105 (N_29105,N_28889,N_28926);
xor U29106 (N_29106,N_28822,N_28892);
or U29107 (N_29107,N_28945,N_28804);
xor U29108 (N_29108,N_28921,N_28885);
nand U29109 (N_29109,N_28896,N_28839);
and U29110 (N_29110,N_28845,N_28838);
nand U29111 (N_29111,N_28842,N_28956);
nor U29112 (N_29112,N_28876,N_28894);
and U29113 (N_29113,N_28920,N_28828);
xnor U29114 (N_29114,N_28777,N_28908);
xor U29115 (N_29115,N_28803,N_28904);
nand U29116 (N_29116,N_28983,N_28898);
xor U29117 (N_29117,N_28782,N_28751);
nor U29118 (N_29118,N_28899,N_28807);
nand U29119 (N_29119,N_28946,N_28880);
nand U29120 (N_29120,N_28931,N_28764);
nor U29121 (N_29121,N_28954,N_28824);
or U29122 (N_29122,N_28765,N_28864);
nand U29123 (N_29123,N_28850,N_28933);
or U29124 (N_29124,N_28776,N_28960);
nor U29125 (N_29125,N_28811,N_28790);
nand U29126 (N_29126,N_28901,N_28809);
and U29127 (N_29127,N_28887,N_28924);
or U29128 (N_29128,N_28786,N_28847);
nand U29129 (N_29129,N_28979,N_28870);
and U29130 (N_29130,N_28929,N_28923);
or U29131 (N_29131,N_28923,N_28985);
xor U29132 (N_29132,N_28887,N_28931);
xnor U29133 (N_29133,N_28925,N_28894);
nand U29134 (N_29134,N_28850,N_28771);
xnor U29135 (N_29135,N_28865,N_28979);
and U29136 (N_29136,N_28922,N_28814);
and U29137 (N_29137,N_28970,N_28784);
nor U29138 (N_29138,N_28806,N_28819);
and U29139 (N_29139,N_28930,N_28824);
nor U29140 (N_29140,N_28831,N_28825);
and U29141 (N_29141,N_28802,N_28886);
nor U29142 (N_29142,N_28822,N_28783);
nor U29143 (N_29143,N_28886,N_28872);
and U29144 (N_29144,N_28827,N_28828);
nor U29145 (N_29145,N_28995,N_28790);
nor U29146 (N_29146,N_28908,N_28914);
xor U29147 (N_29147,N_28809,N_28920);
xor U29148 (N_29148,N_28906,N_28958);
xnor U29149 (N_29149,N_28829,N_28867);
nand U29150 (N_29150,N_28824,N_28976);
nor U29151 (N_29151,N_28756,N_28984);
nor U29152 (N_29152,N_28820,N_28862);
and U29153 (N_29153,N_28953,N_28885);
and U29154 (N_29154,N_28758,N_28953);
and U29155 (N_29155,N_28866,N_28873);
and U29156 (N_29156,N_28782,N_28879);
or U29157 (N_29157,N_28981,N_28771);
xor U29158 (N_29158,N_28789,N_28945);
or U29159 (N_29159,N_28786,N_28759);
and U29160 (N_29160,N_28912,N_28787);
nand U29161 (N_29161,N_28811,N_28831);
xnor U29162 (N_29162,N_28915,N_28797);
nor U29163 (N_29163,N_28929,N_28832);
nand U29164 (N_29164,N_28767,N_28951);
nor U29165 (N_29165,N_28975,N_28987);
xor U29166 (N_29166,N_28887,N_28903);
and U29167 (N_29167,N_28974,N_28936);
nor U29168 (N_29168,N_28999,N_28944);
and U29169 (N_29169,N_28822,N_28974);
nor U29170 (N_29170,N_28955,N_28948);
xnor U29171 (N_29171,N_28930,N_28886);
nand U29172 (N_29172,N_28969,N_28967);
nor U29173 (N_29173,N_28764,N_28795);
xnor U29174 (N_29174,N_28931,N_28970);
xnor U29175 (N_29175,N_28853,N_28768);
nand U29176 (N_29176,N_28863,N_28936);
and U29177 (N_29177,N_28831,N_28993);
xnor U29178 (N_29178,N_28809,N_28797);
nor U29179 (N_29179,N_28927,N_28960);
xor U29180 (N_29180,N_28751,N_28846);
and U29181 (N_29181,N_28921,N_28864);
and U29182 (N_29182,N_28859,N_28993);
nor U29183 (N_29183,N_28850,N_28965);
xnor U29184 (N_29184,N_28913,N_28926);
and U29185 (N_29185,N_28930,N_28762);
nor U29186 (N_29186,N_28981,N_28774);
or U29187 (N_29187,N_28825,N_28971);
or U29188 (N_29188,N_28788,N_28881);
nand U29189 (N_29189,N_28772,N_28880);
nor U29190 (N_29190,N_28772,N_28754);
nor U29191 (N_29191,N_28950,N_28891);
nand U29192 (N_29192,N_28804,N_28881);
and U29193 (N_29193,N_28797,N_28834);
nor U29194 (N_29194,N_28777,N_28987);
and U29195 (N_29195,N_28848,N_28947);
and U29196 (N_29196,N_28973,N_28761);
or U29197 (N_29197,N_28814,N_28888);
and U29198 (N_29198,N_28779,N_28876);
or U29199 (N_29199,N_28797,N_28920);
nand U29200 (N_29200,N_28966,N_28778);
and U29201 (N_29201,N_28959,N_28900);
or U29202 (N_29202,N_28936,N_28757);
or U29203 (N_29203,N_28815,N_28982);
nor U29204 (N_29204,N_28838,N_28929);
and U29205 (N_29205,N_28796,N_28963);
or U29206 (N_29206,N_28849,N_28882);
nor U29207 (N_29207,N_28760,N_28968);
nor U29208 (N_29208,N_28825,N_28834);
nand U29209 (N_29209,N_28937,N_28764);
or U29210 (N_29210,N_28881,N_28962);
xor U29211 (N_29211,N_28802,N_28861);
xor U29212 (N_29212,N_28996,N_28776);
xnor U29213 (N_29213,N_28927,N_28903);
and U29214 (N_29214,N_28981,N_28795);
xnor U29215 (N_29215,N_28828,N_28959);
and U29216 (N_29216,N_28759,N_28843);
nand U29217 (N_29217,N_28890,N_28796);
xor U29218 (N_29218,N_28987,N_28925);
xor U29219 (N_29219,N_28839,N_28873);
nand U29220 (N_29220,N_28790,N_28922);
nand U29221 (N_29221,N_28996,N_28992);
nor U29222 (N_29222,N_28876,N_28758);
nor U29223 (N_29223,N_28772,N_28867);
or U29224 (N_29224,N_28915,N_28941);
and U29225 (N_29225,N_28806,N_28868);
nand U29226 (N_29226,N_28830,N_28857);
xor U29227 (N_29227,N_28882,N_28952);
xor U29228 (N_29228,N_28940,N_28997);
or U29229 (N_29229,N_28807,N_28849);
and U29230 (N_29230,N_28877,N_28750);
and U29231 (N_29231,N_28767,N_28786);
nand U29232 (N_29232,N_28954,N_28880);
or U29233 (N_29233,N_28942,N_28969);
or U29234 (N_29234,N_28846,N_28939);
nor U29235 (N_29235,N_28760,N_28846);
nand U29236 (N_29236,N_28768,N_28854);
nor U29237 (N_29237,N_28861,N_28858);
or U29238 (N_29238,N_28764,N_28842);
xnor U29239 (N_29239,N_28808,N_28942);
xnor U29240 (N_29240,N_28892,N_28799);
xor U29241 (N_29241,N_28774,N_28773);
xnor U29242 (N_29242,N_28958,N_28793);
xnor U29243 (N_29243,N_28863,N_28835);
nand U29244 (N_29244,N_28988,N_28888);
nand U29245 (N_29245,N_28862,N_28962);
xor U29246 (N_29246,N_28932,N_28853);
nor U29247 (N_29247,N_28896,N_28972);
and U29248 (N_29248,N_28757,N_28812);
xnor U29249 (N_29249,N_28776,N_28840);
nor U29250 (N_29250,N_29168,N_29163);
xnor U29251 (N_29251,N_29121,N_29106);
and U29252 (N_29252,N_29234,N_29068);
xor U29253 (N_29253,N_29178,N_29043);
nand U29254 (N_29254,N_29119,N_29045);
nor U29255 (N_29255,N_29114,N_29172);
xor U29256 (N_29256,N_29102,N_29115);
and U29257 (N_29257,N_29012,N_29143);
or U29258 (N_29258,N_29123,N_29064);
xor U29259 (N_29259,N_29004,N_29118);
xor U29260 (N_29260,N_29108,N_29061);
xnor U29261 (N_29261,N_29097,N_29036);
and U29262 (N_29262,N_29050,N_29190);
nand U29263 (N_29263,N_29194,N_29048);
xnor U29264 (N_29264,N_29035,N_29238);
nand U29265 (N_29265,N_29140,N_29040);
nand U29266 (N_29266,N_29037,N_29113);
nand U29267 (N_29267,N_29204,N_29104);
and U29268 (N_29268,N_29007,N_29155);
and U29269 (N_29269,N_29205,N_29221);
xnor U29270 (N_29270,N_29105,N_29165);
or U29271 (N_29271,N_29162,N_29028);
nor U29272 (N_29272,N_29066,N_29233);
nand U29273 (N_29273,N_29084,N_29089);
or U29274 (N_29274,N_29224,N_29207);
nand U29275 (N_29275,N_29131,N_29135);
nand U29276 (N_29276,N_29167,N_29175);
and U29277 (N_29277,N_29060,N_29023);
or U29278 (N_29278,N_29055,N_29197);
or U29279 (N_29279,N_29242,N_29147);
nand U29280 (N_29280,N_29183,N_29006);
nand U29281 (N_29281,N_29169,N_29141);
xor U29282 (N_29282,N_29085,N_29029);
nor U29283 (N_29283,N_29201,N_29015);
and U29284 (N_29284,N_29019,N_29039);
and U29285 (N_29285,N_29216,N_29005);
xnor U29286 (N_29286,N_29145,N_29239);
nand U29287 (N_29287,N_29200,N_29189);
or U29288 (N_29288,N_29003,N_29100);
xor U29289 (N_29289,N_29014,N_29179);
or U29290 (N_29290,N_29110,N_29170);
xnor U29291 (N_29291,N_29134,N_29126);
or U29292 (N_29292,N_29191,N_29228);
nand U29293 (N_29293,N_29151,N_29054);
nor U29294 (N_29294,N_29246,N_29127);
nor U29295 (N_29295,N_29001,N_29120);
nand U29296 (N_29296,N_29022,N_29219);
and U29297 (N_29297,N_29171,N_29111);
or U29298 (N_29298,N_29230,N_29236);
or U29299 (N_29299,N_29034,N_29229);
nor U29300 (N_29300,N_29020,N_29152);
xnor U29301 (N_29301,N_29052,N_29027);
nand U29302 (N_29302,N_29166,N_29033);
or U29303 (N_29303,N_29182,N_29099);
nor U29304 (N_29304,N_29016,N_29018);
and U29305 (N_29305,N_29196,N_29009);
xnor U29306 (N_29306,N_29227,N_29109);
nor U29307 (N_29307,N_29214,N_29133);
xnor U29308 (N_29308,N_29128,N_29241);
nand U29309 (N_29309,N_29209,N_29180);
or U29310 (N_29310,N_29138,N_29103);
xor U29311 (N_29311,N_29144,N_29074);
nand U29312 (N_29312,N_29210,N_29011);
xnor U29313 (N_29313,N_29116,N_29218);
nor U29314 (N_29314,N_29146,N_29161);
nand U29315 (N_29315,N_29038,N_29096);
xor U29316 (N_29316,N_29046,N_29002);
or U29317 (N_29317,N_29042,N_29093);
xnor U29318 (N_29318,N_29053,N_29211);
nor U29319 (N_29319,N_29206,N_29160);
nand U29320 (N_29320,N_29184,N_29159);
xor U29321 (N_29321,N_29245,N_29157);
xnor U29322 (N_29322,N_29030,N_29031);
xor U29323 (N_29323,N_29149,N_29235);
nand U29324 (N_29324,N_29112,N_29044);
nand U29325 (N_29325,N_29008,N_29076);
or U29326 (N_29326,N_29185,N_29208);
nor U29327 (N_29327,N_29021,N_29177);
nand U29328 (N_29328,N_29153,N_29173);
or U29329 (N_29329,N_29198,N_29081);
nor U29330 (N_29330,N_29243,N_29083);
nor U29331 (N_29331,N_29174,N_29058);
nand U29332 (N_29332,N_29130,N_29215);
nor U29333 (N_29333,N_29193,N_29057);
or U29334 (N_29334,N_29148,N_29080);
or U29335 (N_29335,N_29079,N_29176);
or U29336 (N_29336,N_29217,N_29063);
or U29337 (N_29337,N_29158,N_29122);
xnor U29338 (N_29338,N_29186,N_29013);
and U29339 (N_29339,N_29137,N_29240);
and U29340 (N_29340,N_29117,N_29095);
xnor U29341 (N_29341,N_29222,N_29010);
nor U29342 (N_29342,N_29077,N_29107);
nand U29343 (N_29343,N_29067,N_29248);
and U29344 (N_29344,N_29032,N_29212);
and U29345 (N_29345,N_29087,N_29164);
xnor U29346 (N_29346,N_29059,N_29192);
and U29347 (N_29347,N_29203,N_29223);
nand U29348 (N_29348,N_29195,N_29139);
nor U29349 (N_29349,N_29000,N_29199);
xnor U29350 (N_29350,N_29136,N_29069);
nand U29351 (N_29351,N_29082,N_29125);
and U29352 (N_29352,N_29231,N_29098);
xor U29353 (N_29353,N_29244,N_29075);
and U29354 (N_29354,N_29226,N_29154);
nor U29355 (N_29355,N_29220,N_29142);
or U29356 (N_29356,N_29086,N_29078);
nand U29357 (N_29357,N_29049,N_29051);
or U29358 (N_29358,N_29041,N_29088);
nor U29359 (N_29359,N_29017,N_29094);
or U29360 (N_29360,N_29092,N_29090);
nand U29361 (N_29361,N_29156,N_29124);
or U29362 (N_29362,N_29072,N_29101);
and U29363 (N_29363,N_29225,N_29073);
and U29364 (N_29364,N_29213,N_29232);
or U29365 (N_29365,N_29249,N_29202);
xnor U29366 (N_29366,N_29056,N_29026);
and U29367 (N_29367,N_29091,N_29132);
xor U29368 (N_29368,N_29047,N_29065);
nand U29369 (N_29369,N_29071,N_29129);
nor U29370 (N_29370,N_29025,N_29187);
nor U29371 (N_29371,N_29237,N_29181);
nand U29372 (N_29372,N_29024,N_29070);
xnor U29373 (N_29373,N_29188,N_29247);
or U29374 (N_29374,N_29150,N_29062);
and U29375 (N_29375,N_29035,N_29082);
and U29376 (N_29376,N_29167,N_29154);
nand U29377 (N_29377,N_29024,N_29135);
nand U29378 (N_29378,N_29221,N_29224);
and U29379 (N_29379,N_29142,N_29096);
nand U29380 (N_29380,N_29156,N_29032);
nand U29381 (N_29381,N_29130,N_29148);
nand U29382 (N_29382,N_29024,N_29111);
nand U29383 (N_29383,N_29240,N_29174);
and U29384 (N_29384,N_29001,N_29050);
or U29385 (N_29385,N_29024,N_29066);
or U29386 (N_29386,N_29039,N_29220);
nor U29387 (N_29387,N_29121,N_29228);
and U29388 (N_29388,N_29176,N_29131);
xnor U29389 (N_29389,N_29114,N_29027);
nor U29390 (N_29390,N_29110,N_29076);
and U29391 (N_29391,N_29041,N_29125);
nor U29392 (N_29392,N_29044,N_29131);
xnor U29393 (N_29393,N_29225,N_29066);
nand U29394 (N_29394,N_29107,N_29201);
nand U29395 (N_29395,N_29230,N_29164);
and U29396 (N_29396,N_29206,N_29021);
or U29397 (N_29397,N_29091,N_29218);
and U29398 (N_29398,N_29034,N_29046);
nor U29399 (N_29399,N_29181,N_29147);
and U29400 (N_29400,N_29134,N_29130);
xor U29401 (N_29401,N_29020,N_29099);
nand U29402 (N_29402,N_29145,N_29036);
or U29403 (N_29403,N_29199,N_29221);
and U29404 (N_29404,N_29192,N_29230);
xor U29405 (N_29405,N_29111,N_29210);
nor U29406 (N_29406,N_29132,N_29006);
xor U29407 (N_29407,N_29075,N_29243);
nor U29408 (N_29408,N_29150,N_29013);
xnor U29409 (N_29409,N_29233,N_29026);
and U29410 (N_29410,N_29064,N_29012);
nand U29411 (N_29411,N_29025,N_29136);
or U29412 (N_29412,N_29044,N_29226);
nor U29413 (N_29413,N_29118,N_29171);
nand U29414 (N_29414,N_29154,N_29076);
nor U29415 (N_29415,N_29081,N_29075);
nor U29416 (N_29416,N_29168,N_29199);
or U29417 (N_29417,N_29129,N_29167);
or U29418 (N_29418,N_29107,N_29168);
nor U29419 (N_29419,N_29057,N_29154);
or U29420 (N_29420,N_29215,N_29157);
or U29421 (N_29421,N_29178,N_29155);
nor U29422 (N_29422,N_29059,N_29248);
or U29423 (N_29423,N_29006,N_29046);
and U29424 (N_29424,N_29100,N_29238);
nand U29425 (N_29425,N_29053,N_29206);
nand U29426 (N_29426,N_29192,N_29238);
nand U29427 (N_29427,N_29055,N_29110);
nor U29428 (N_29428,N_29164,N_29040);
nor U29429 (N_29429,N_29126,N_29082);
xnor U29430 (N_29430,N_29087,N_29066);
nor U29431 (N_29431,N_29207,N_29092);
nor U29432 (N_29432,N_29215,N_29005);
nor U29433 (N_29433,N_29227,N_29176);
and U29434 (N_29434,N_29199,N_29137);
or U29435 (N_29435,N_29062,N_29064);
and U29436 (N_29436,N_29102,N_29118);
and U29437 (N_29437,N_29174,N_29092);
and U29438 (N_29438,N_29018,N_29128);
nand U29439 (N_29439,N_29122,N_29095);
nor U29440 (N_29440,N_29138,N_29160);
and U29441 (N_29441,N_29046,N_29172);
xnor U29442 (N_29442,N_29162,N_29084);
and U29443 (N_29443,N_29230,N_29146);
xor U29444 (N_29444,N_29216,N_29142);
nand U29445 (N_29445,N_29230,N_29017);
or U29446 (N_29446,N_29105,N_29152);
nor U29447 (N_29447,N_29113,N_29041);
and U29448 (N_29448,N_29138,N_29099);
or U29449 (N_29449,N_29139,N_29248);
and U29450 (N_29450,N_29174,N_29126);
nor U29451 (N_29451,N_29152,N_29045);
nor U29452 (N_29452,N_29048,N_29180);
and U29453 (N_29453,N_29005,N_29130);
xor U29454 (N_29454,N_29043,N_29018);
and U29455 (N_29455,N_29210,N_29096);
and U29456 (N_29456,N_29205,N_29170);
xor U29457 (N_29457,N_29065,N_29036);
nand U29458 (N_29458,N_29150,N_29163);
xor U29459 (N_29459,N_29019,N_29103);
or U29460 (N_29460,N_29035,N_29040);
nor U29461 (N_29461,N_29040,N_29001);
or U29462 (N_29462,N_29054,N_29217);
xor U29463 (N_29463,N_29014,N_29018);
and U29464 (N_29464,N_29228,N_29053);
nand U29465 (N_29465,N_29082,N_29132);
xnor U29466 (N_29466,N_29165,N_29210);
xor U29467 (N_29467,N_29076,N_29200);
xor U29468 (N_29468,N_29130,N_29049);
xor U29469 (N_29469,N_29000,N_29172);
or U29470 (N_29470,N_29197,N_29224);
and U29471 (N_29471,N_29226,N_29061);
and U29472 (N_29472,N_29128,N_29088);
and U29473 (N_29473,N_29000,N_29130);
nand U29474 (N_29474,N_29200,N_29213);
and U29475 (N_29475,N_29232,N_29119);
xor U29476 (N_29476,N_29038,N_29046);
and U29477 (N_29477,N_29159,N_29026);
and U29478 (N_29478,N_29168,N_29122);
or U29479 (N_29479,N_29075,N_29112);
xor U29480 (N_29480,N_29075,N_29018);
nand U29481 (N_29481,N_29170,N_29203);
xor U29482 (N_29482,N_29010,N_29089);
and U29483 (N_29483,N_29044,N_29096);
nor U29484 (N_29484,N_29201,N_29085);
and U29485 (N_29485,N_29170,N_29149);
and U29486 (N_29486,N_29099,N_29130);
or U29487 (N_29487,N_29185,N_29228);
and U29488 (N_29488,N_29180,N_29021);
and U29489 (N_29489,N_29112,N_29002);
and U29490 (N_29490,N_29003,N_29198);
xnor U29491 (N_29491,N_29124,N_29135);
and U29492 (N_29492,N_29002,N_29227);
xnor U29493 (N_29493,N_29038,N_29125);
nand U29494 (N_29494,N_29158,N_29231);
or U29495 (N_29495,N_29063,N_29213);
and U29496 (N_29496,N_29205,N_29115);
xor U29497 (N_29497,N_29100,N_29207);
nand U29498 (N_29498,N_29205,N_29088);
nand U29499 (N_29499,N_29025,N_29057);
or U29500 (N_29500,N_29372,N_29326);
xnor U29501 (N_29501,N_29388,N_29269);
nand U29502 (N_29502,N_29268,N_29395);
nor U29503 (N_29503,N_29391,N_29282);
nand U29504 (N_29504,N_29411,N_29433);
or U29505 (N_29505,N_29412,N_29496);
nand U29506 (N_29506,N_29470,N_29347);
and U29507 (N_29507,N_29351,N_29416);
nand U29508 (N_29508,N_29295,N_29324);
nor U29509 (N_29509,N_29485,N_29283);
and U29510 (N_29510,N_29493,N_29498);
nor U29511 (N_29511,N_29370,N_29253);
xnor U29512 (N_29512,N_29284,N_29374);
nor U29513 (N_29513,N_29309,N_29438);
or U29514 (N_29514,N_29273,N_29301);
or U29515 (N_29515,N_29319,N_29421);
or U29516 (N_29516,N_29341,N_29442);
and U29517 (N_29517,N_29257,N_29336);
nand U29518 (N_29518,N_29311,N_29436);
nand U29519 (N_29519,N_29457,N_29304);
and U29520 (N_29520,N_29437,N_29486);
and U29521 (N_29521,N_29356,N_29400);
nor U29522 (N_29522,N_29499,N_29300);
nand U29523 (N_29523,N_29463,N_29358);
and U29524 (N_29524,N_29320,N_29318);
or U29525 (N_29525,N_29366,N_29260);
or U29526 (N_29526,N_29277,N_29445);
nor U29527 (N_29527,N_29443,N_29387);
xor U29528 (N_29528,N_29354,N_29275);
xnor U29529 (N_29529,N_29394,N_29346);
nand U29530 (N_29530,N_29325,N_29480);
and U29531 (N_29531,N_29410,N_29430);
nor U29532 (N_29532,N_29270,N_29469);
xnor U29533 (N_29533,N_29456,N_29413);
nor U29534 (N_29534,N_29397,N_29392);
nand U29535 (N_29535,N_29314,N_29407);
xnor U29536 (N_29536,N_29434,N_29353);
and U29537 (N_29537,N_29479,N_29481);
nor U29538 (N_29538,N_29322,N_29348);
nor U29539 (N_29539,N_29290,N_29276);
xnor U29540 (N_29540,N_29255,N_29382);
nand U29541 (N_29541,N_29333,N_29425);
or U29542 (N_29542,N_29450,N_29254);
nand U29543 (N_29543,N_29334,N_29383);
nor U29544 (N_29544,N_29451,N_29471);
and U29545 (N_29545,N_29298,N_29377);
nor U29546 (N_29546,N_29250,N_29251);
nor U29547 (N_29547,N_29332,N_29310);
or U29548 (N_29548,N_29490,N_29261);
xnor U29549 (N_29549,N_29449,N_29452);
or U29550 (N_29550,N_29288,N_29335);
or U29551 (N_29551,N_29426,N_29466);
nor U29552 (N_29552,N_29308,N_29287);
and U29553 (N_29553,N_29475,N_29403);
nand U29554 (N_29554,N_29398,N_29262);
nor U29555 (N_29555,N_29307,N_29313);
nand U29556 (N_29556,N_29345,N_29404);
nand U29557 (N_29557,N_29331,N_29483);
xnor U29558 (N_29558,N_29381,N_29352);
nor U29559 (N_29559,N_29409,N_29289);
nor U29560 (N_29560,N_29462,N_29267);
or U29561 (N_29561,N_29266,N_29464);
nor U29562 (N_29562,N_29292,N_29484);
xor U29563 (N_29563,N_29459,N_29495);
xnor U29564 (N_29564,N_29274,N_29359);
nand U29565 (N_29565,N_29460,N_29367);
nand U29566 (N_29566,N_29256,N_29265);
and U29567 (N_29567,N_29429,N_29427);
or U29568 (N_29568,N_29378,N_29379);
and U29569 (N_29569,N_29355,N_29375);
or U29570 (N_29570,N_29406,N_29448);
xor U29571 (N_29571,N_29357,N_29362);
nand U29572 (N_29572,N_29390,N_29419);
nor U29573 (N_29573,N_29339,N_29306);
or U29574 (N_29574,N_29293,N_29491);
xnor U29575 (N_29575,N_29323,N_29414);
nand U29576 (N_29576,N_29384,N_29302);
xnor U29577 (N_29577,N_29278,N_29472);
and U29578 (N_29578,N_29312,N_29369);
nor U29579 (N_29579,N_29476,N_29497);
nor U29580 (N_29580,N_29477,N_29363);
nand U29581 (N_29581,N_29316,N_29371);
nand U29582 (N_29582,N_29350,N_29368);
and U29583 (N_29583,N_29386,N_29465);
nor U29584 (N_29584,N_29330,N_29263);
or U29585 (N_29585,N_29281,N_29399);
or U29586 (N_29586,N_29294,N_29482);
and U29587 (N_29587,N_29286,N_29373);
or U29588 (N_29588,N_29328,N_29258);
or U29589 (N_29589,N_29280,N_29279);
xnor U29590 (N_29590,N_29401,N_29297);
xnor U29591 (N_29591,N_29252,N_29299);
xnor U29592 (N_29592,N_29271,N_29343);
and U29593 (N_29593,N_29360,N_29380);
and U29594 (N_29594,N_29361,N_29424);
nand U29595 (N_29595,N_29285,N_29487);
or U29596 (N_29596,N_29444,N_29420);
and U29597 (N_29597,N_29473,N_29303);
nand U29598 (N_29598,N_29454,N_29364);
nand U29599 (N_29599,N_29440,N_29337);
xor U29600 (N_29600,N_29467,N_29264);
and U29601 (N_29601,N_29494,N_29422);
xor U29602 (N_29602,N_29340,N_29455);
xor U29603 (N_29603,N_29291,N_29458);
xor U29604 (N_29604,N_29329,N_29305);
xor U29605 (N_29605,N_29492,N_29418);
nor U29606 (N_29606,N_29342,N_29478);
nor U29607 (N_29607,N_29393,N_29272);
nor U29608 (N_29608,N_29327,N_29435);
and U29609 (N_29609,N_29408,N_29441);
and U29610 (N_29610,N_29344,N_29461);
and U29611 (N_29611,N_29317,N_29417);
or U29612 (N_29612,N_29338,N_29489);
nor U29613 (N_29613,N_29385,N_29321);
xnor U29614 (N_29614,N_29428,N_29453);
nand U29615 (N_29615,N_29296,N_29468);
nor U29616 (N_29616,N_29259,N_29405);
and U29617 (N_29617,N_29415,N_29376);
nand U29618 (N_29618,N_29474,N_29389);
nand U29619 (N_29619,N_29365,N_29488);
nand U29620 (N_29620,N_29315,N_29431);
nor U29621 (N_29621,N_29439,N_29396);
or U29622 (N_29622,N_29423,N_29349);
and U29623 (N_29623,N_29447,N_29402);
xnor U29624 (N_29624,N_29432,N_29446);
nand U29625 (N_29625,N_29491,N_29276);
xnor U29626 (N_29626,N_29384,N_29486);
nand U29627 (N_29627,N_29335,N_29266);
xnor U29628 (N_29628,N_29443,N_29406);
and U29629 (N_29629,N_29323,N_29437);
or U29630 (N_29630,N_29281,N_29278);
nand U29631 (N_29631,N_29426,N_29355);
nand U29632 (N_29632,N_29495,N_29485);
xor U29633 (N_29633,N_29267,N_29429);
and U29634 (N_29634,N_29487,N_29420);
nand U29635 (N_29635,N_29405,N_29338);
and U29636 (N_29636,N_29496,N_29484);
and U29637 (N_29637,N_29484,N_29267);
or U29638 (N_29638,N_29333,N_29378);
nand U29639 (N_29639,N_29401,N_29284);
or U29640 (N_29640,N_29362,N_29382);
and U29641 (N_29641,N_29279,N_29393);
xor U29642 (N_29642,N_29435,N_29388);
nor U29643 (N_29643,N_29312,N_29318);
and U29644 (N_29644,N_29279,N_29281);
and U29645 (N_29645,N_29259,N_29396);
xor U29646 (N_29646,N_29271,N_29432);
xnor U29647 (N_29647,N_29271,N_29348);
and U29648 (N_29648,N_29437,N_29412);
or U29649 (N_29649,N_29496,N_29293);
and U29650 (N_29650,N_29364,N_29398);
and U29651 (N_29651,N_29332,N_29383);
or U29652 (N_29652,N_29417,N_29286);
xnor U29653 (N_29653,N_29423,N_29497);
nand U29654 (N_29654,N_29339,N_29397);
xor U29655 (N_29655,N_29373,N_29337);
xnor U29656 (N_29656,N_29497,N_29458);
nand U29657 (N_29657,N_29478,N_29395);
nor U29658 (N_29658,N_29290,N_29423);
or U29659 (N_29659,N_29387,N_29408);
nor U29660 (N_29660,N_29433,N_29446);
and U29661 (N_29661,N_29388,N_29461);
xor U29662 (N_29662,N_29346,N_29481);
or U29663 (N_29663,N_29356,N_29428);
xnor U29664 (N_29664,N_29358,N_29260);
xnor U29665 (N_29665,N_29398,N_29425);
nand U29666 (N_29666,N_29381,N_29445);
and U29667 (N_29667,N_29402,N_29314);
or U29668 (N_29668,N_29262,N_29386);
or U29669 (N_29669,N_29370,N_29279);
nor U29670 (N_29670,N_29462,N_29456);
and U29671 (N_29671,N_29352,N_29436);
or U29672 (N_29672,N_29360,N_29268);
nor U29673 (N_29673,N_29271,N_29382);
xor U29674 (N_29674,N_29315,N_29497);
nor U29675 (N_29675,N_29275,N_29434);
nand U29676 (N_29676,N_29487,N_29466);
or U29677 (N_29677,N_29465,N_29298);
and U29678 (N_29678,N_29359,N_29431);
nor U29679 (N_29679,N_29286,N_29301);
or U29680 (N_29680,N_29343,N_29413);
xnor U29681 (N_29681,N_29450,N_29323);
xor U29682 (N_29682,N_29485,N_29432);
or U29683 (N_29683,N_29274,N_29357);
nor U29684 (N_29684,N_29266,N_29403);
xnor U29685 (N_29685,N_29411,N_29449);
and U29686 (N_29686,N_29478,N_29494);
nand U29687 (N_29687,N_29413,N_29416);
and U29688 (N_29688,N_29382,N_29354);
nand U29689 (N_29689,N_29446,N_29337);
and U29690 (N_29690,N_29402,N_29303);
or U29691 (N_29691,N_29490,N_29260);
or U29692 (N_29692,N_29482,N_29287);
and U29693 (N_29693,N_29378,N_29395);
nor U29694 (N_29694,N_29283,N_29404);
nor U29695 (N_29695,N_29403,N_29306);
nand U29696 (N_29696,N_29393,N_29291);
or U29697 (N_29697,N_29259,N_29323);
nor U29698 (N_29698,N_29384,N_29476);
and U29699 (N_29699,N_29414,N_29399);
or U29700 (N_29700,N_29340,N_29496);
xor U29701 (N_29701,N_29460,N_29492);
xnor U29702 (N_29702,N_29375,N_29282);
or U29703 (N_29703,N_29316,N_29324);
and U29704 (N_29704,N_29374,N_29393);
xnor U29705 (N_29705,N_29498,N_29352);
and U29706 (N_29706,N_29268,N_29404);
and U29707 (N_29707,N_29353,N_29391);
nor U29708 (N_29708,N_29482,N_29276);
nand U29709 (N_29709,N_29446,N_29470);
and U29710 (N_29710,N_29303,N_29462);
or U29711 (N_29711,N_29338,N_29378);
nor U29712 (N_29712,N_29433,N_29304);
or U29713 (N_29713,N_29455,N_29462);
nor U29714 (N_29714,N_29293,N_29453);
or U29715 (N_29715,N_29492,N_29270);
nor U29716 (N_29716,N_29290,N_29373);
nor U29717 (N_29717,N_29279,N_29350);
nand U29718 (N_29718,N_29264,N_29409);
nor U29719 (N_29719,N_29303,N_29371);
or U29720 (N_29720,N_29432,N_29471);
nand U29721 (N_29721,N_29283,N_29465);
and U29722 (N_29722,N_29473,N_29284);
xnor U29723 (N_29723,N_29343,N_29323);
xnor U29724 (N_29724,N_29456,N_29328);
nand U29725 (N_29725,N_29420,N_29465);
nor U29726 (N_29726,N_29418,N_29448);
or U29727 (N_29727,N_29277,N_29373);
xnor U29728 (N_29728,N_29349,N_29282);
or U29729 (N_29729,N_29426,N_29492);
xor U29730 (N_29730,N_29405,N_29473);
nor U29731 (N_29731,N_29481,N_29429);
or U29732 (N_29732,N_29452,N_29455);
nand U29733 (N_29733,N_29427,N_29370);
nand U29734 (N_29734,N_29370,N_29388);
xor U29735 (N_29735,N_29272,N_29285);
nor U29736 (N_29736,N_29360,N_29379);
xnor U29737 (N_29737,N_29285,N_29388);
nand U29738 (N_29738,N_29395,N_29458);
nor U29739 (N_29739,N_29362,N_29322);
xor U29740 (N_29740,N_29441,N_29286);
nor U29741 (N_29741,N_29333,N_29464);
xor U29742 (N_29742,N_29490,N_29349);
nor U29743 (N_29743,N_29484,N_29251);
or U29744 (N_29744,N_29315,N_29328);
nor U29745 (N_29745,N_29273,N_29379);
xor U29746 (N_29746,N_29333,N_29434);
xor U29747 (N_29747,N_29340,N_29336);
and U29748 (N_29748,N_29274,N_29367);
nand U29749 (N_29749,N_29417,N_29250);
nand U29750 (N_29750,N_29638,N_29709);
nand U29751 (N_29751,N_29726,N_29548);
and U29752 (N_29752,N_29596,N_29713);
xor U29753 (N_29753,N_29604,N_29724);
xnor U29754 (N_29754,N_29582,N_29579);
nand U29755 (N_29755,N_29568,N_29518);
nor U29756 (N_29756,N_29689,N_29619);
xor U29757 (N_29757,N_29748,N_29667);
nor U29758 (N_29758,N_29678,N_29676);
and U29759 (N_29759,N_29672,N_29690);
nand U29760 (N_29760,N_29613,N_29730);
or U29761 (N_29761,N_29505,N_29686);
xor U29762 (N_29762,N_29661,N_29520);
xor U29763 (N_29763,N_29610,N_29653);
nand U29764 (N_29764,N_29578,N_29607);
nor U29765 (N_29765,N_29515,N_29500);
xor U29766 (N_29766,N_29595,N_29727);
nand U29767 (N_29767,N_29647,N_29564);
nand U29768 (N_29768,N_29587,N_29631);
xor U29769 (N_29769,N_29592,N_29719);
nand U29770 (N_29770,N_29616,N_29572);
xnor U29771 (N_29771,N_29696,N_29585);
xor U29772 (N_29772,N_29669,N_29606);
or U29773 (N_29773,N_29714,N_29560);
nor U29774 (N_29774,N_29544,N_29557);
nor U29775 (N_29775,N_29654,N_29567);
nor U29776 (N_29776,N_29575,N_29543);
or U29777 (N_29777,N_29675,N_29723);
or U29778 (N_29778,N_29683,N_29721);
or U29779 (N_29779,N_29644,N_29687);
nand U29780 (N_29780,N_29706,N_29549);
xor U29781 (N_29781,N_29627,N_29536);
and U29782 (N_29782,N_29577,N_29569);
or U29783 (N_29783,N_29747,N_29733);
nand U29784 (N_29784,N_29666,N_29522);
nand U29785 (N_29785,N_29664,N_29720);
nor U29786 (N_29786,N_29708,N_29673);
xnor U29787 (N_29787,N_29540,N_29697);
xnor U29788 (N_29788,N_29502,N_29710);
or U29789 (N_29789,N_29609,N_29651);
nand U29790 (N_29790,N_29597,N_29702);
xnor U29791 (N_29791,N_29642,N_29660);
nor U29792 (N_29792,N_29692,N_29605);
and U29793 (N_29793,N_29739,N_29711);
and U29794 (N_29794,N_29657,N_29700);
xor U29795 (N_29795,N_29506,N_29599);
nand U29796 (N_29796,N_29684,N_29538);
and U29797 (N_29797,N_29519,N_29583);
nand U29798 (N_29798,N_29531,N_29523);
and U29799 (N_29799,N_29593,N_29509);
and U29800 (N_29800,N_29704,N_29510);
xnor U29801 (N_29801,N_29680,N_29581);
nand U29802 (N_29802,N_29632,N_29628);
xor U29803 (N_29803,N_29741,N_29646);
or U29804 (N_29804,N_29580,N_29655);
nor U29805 (N_29805,N_29508,N_29542);
nor U29806 (N_29806,N_29641,N_29617);
or U29807 (N_29807,N_29624,N_29643);
xnor U29808 (N_29808,N_29551,N_29566);
nor U29809 (N_29809,N_29640,N_29698);
xnor U29810 (N_29810,N_29731,N_29591);
xor U29811 (N_29811,N_29512,N_29504);
xor U29812 (N_29812,N_29717,N_29728);
xnor U29813 (N_29813,N_29695,N_29746);
or U29814 (N_29814,N_29535,N_29740);
or U29815 (N_29815,N_29659,N_29744);
or U29816 (N_29816,N_29552,N_29511);
and U29817 (N_29817,N_29586,N_29537);
nand U29818 (N_29818,N_29663,N_29550);
and U29819 (N_29819,N_29681,N_29693);
and U29820 (N_29820,N_29594,N_29530);
xor U29821 (N_29821,N_29611,N_29735);
xor U29822 (N_29822,N_29742,N_29658);
nor U29823 (N_29823,N_29598,N_29691);
nand U29824 (N_29824,N_29612,N_29555);
nand U29825 (N_29825,N_29534,N_29745);
xnor U29826 (N_29826,N_29722,N_29629);
nor U29827 (N_29827,N_29635,N_29526);
and U29828 (N_29828,N_29529,N_29625);
and U29829 (N_29829,N_29749,N_29737);
or U29830 (N_29830,N_29561,N_29620);
or U29831 (N_29831,N_29662,N_29715);
xor U29832 (N_29832,N_29725,N_29553);
and U29833 (N_29833,N_29712,N_29630);
and U29834 (N_29834,N_29614,N_29716);
xor U29835 (N_29835,N_29685,N_29615);
xnor U29836 (N_29836,N_29584,N_29602);
xnor U29837 (N_29837,N_29718,N_29688);
and U29838 (N_29838,N_29736,N_29626);
and U29839 (N_29839,N_29528,N_29565);
nand U29840 (N_29840,N_29645,N_29514);
and U29841 (N_29841,N_29590,N_29633);
nor U29842 (N_29842,N_29573,N_29541);
nor U29843 (N_29843,N_29732,N_29603);
or U29844 (N_29844,N_29707,N_29558);
nand U29845 (N_29845,N_29694,N_29743);
and U29846 (N_29846,N_29554,N_29637);
or U29847 (N_29847,N_29588,N_29532);
and U29848 (N_29848,N_29559,N_29513);
or U29849 (N_29849,N_29527,N_29668);
nor U29850 (N_29850,N_29623,N_29556);
nand U29851 (N_29851,N_29671,N_29703);
xnor U29852 (N_29852,N_29665,N_29563);
nor U29853 (N_29853,N_29547,N_29699);
or U29854 (N_29854,N_29533,N_29639);
and U29855 (N_29855,N_29516,N_29682);
nor U29856 (N_29856,N_29601,N_29618);
nand U29857 (N_29857,N_29525,N_29608);
and U29858 (N_29858,N_29705,N_29656);
xor U29859 (N_29859,N_29652,N_29574);
and U29860 (N_29860,N_29734,N_29634);
nand U29861 (N_29861,N_29521,N_29576);
xor U29862 (N_29862,N_29729,N_29524);
xor U29863 (N_29863,N_29738,N_29501);
and U29864 (N_29864,N_29600,N_29589);
nor U29865 (N_29865,N_29677,N_29545);
and U29866 (N_29866,N_29701,N_29649);
or U29867 (N_29867,N_29539,N_29674);
and U29868 (N_29868,N_29562,N_29571);
and U29869 (N_29869,N_29648,N_29507);
nor U29870 (N_29870,N_29570,N_29670);
nand U29871 (N_29871,N_29622,N_29636);
or U29872 (N_29872,N_29621,N_29503);
xnor U29873 (N_29873,N_29517,N_29679);
nand U29874 (N_29874,N_29650,N_29546);
or U29875 (N_29875,N_29593,N_29581);
nor U29876 (N_29876,N_29586,N_29695);
nand U29877 (N_29877,N_29669,N_29577);
nand U29878 (N_29878,N_29626,N_29559);
nor U29879 (N_29879,N_29544,N_29570);
and U29880 (N_29880,N_29510,N_29722);
nor U29881 (N_29881,N_29718,N_29644);
and U29882 (N_29882,N_29598,N_29683);
nand U29883 (N_29883,N_29725,N_29582);
nor U29884 (N_29884,N_29696,N_29666);
and U29885 (N_29885,N_29717,N_29731);
nor U29886 (N_29886,N_29565,N_29695);
or U29887 (N_29887,N_29594,N_29710);
and U29888 (N_29888,N_29721,N_29607);
or U29889 (N_29889,N_29586,N_29611);
xnor U29890 (N_29890,N_29737,N_29645);
nand U29891 (N_29891,N_29741,N_29723);
xor U29892 (N_29892,N_29695,N_29510);
xor U29893 (N_29893,N_29696,N_29700);
or U29894 (N_29894,N_29553,N_29534);
xnor U29895 (N_29895,N_29744,N_29730);
xor U29896 (N_29896,N_29692,N_29667);
nor U29897 (N_29897,N_29509,N_29577);
and U29898 (N_29898,N_29701,N_29529);
or U29899 (N_29899,N_29735,N_29567);
nand U29900 (N_29900,N_29570,N_29648);
nor U29901 (N_29901,N_29602,N_29623);
nor U29902 (N_29902,N_29571,N_29667);
nand U29903 (N_29903,N_29547,N_29570);
nand U29904 (N_29904,N_29728,N_29531);
and U29905 (N_29905,N_29553,N_29516);
nor U29906 (N_29906,N_29576,N_29670);
or U29907 (N_29907,N_29744,N_29500);
and U29908 (N_29908,N_29735,N_29501);
and U29909 (N_29909,N_29558,N_29522);
nor U29910 (N_29910,N_29740,N_29648);
nand U29911 (N_29911,N_29667,N_29651);
xor U29912 (N_29912,N_29682,N_29692);
or U29913 (N_29913,N_29739,N_29554);
xor U29914 (N_29914,N_29595,N_29744);
or U29915 (N_29915,N_29516,N_29600);
or U29916 (N_29916,N_29652,N_29692);
nand U29917 (N_29917,N_29578,N_29613);
nand U29918 (N_29918,N_29731,N_29679);
nor U29919 (N_29919,N_29706,N_29530);
xor U29920 (N_29920,N_29709,N_29565);
or U29921 (N_29921,N_29596,N_29505);
and U29922 (N_29922,N_29743,N_29548);
nor U29923 (N_29923,N_29728,N_29656);
xor U29924 (N_29924,N_29608,N_29614);
xor U29925 (N_29925,N_29589,N_29593);
nand U29926 (N_29926,N_29721,N_29636);
and U29927 (N_29927,N_29540,N_29693);
nand U29928 (N_29928,N_29716,N_29593);
xor U29929 (N_29929,N_29608,N_29543);
nor U29930 (N_29930,N_29560,N_29686);
and U29931 (N_29931,N_29706,N_29522);
nand U29932 (N_29932,N_29689,N_29665);
or U29933 (N_29933,N_29572,N_29727);
or U29934 (N_29934,N_29635,N_29512);
nor U29935 (N_29935,N_29517,N_29592);
or U29936 (N_29936,N_29717,N_29649);
and U29937 (N_29937,N_29561,N_29562);
and U29938 (N_29938,N_29675,N_29691);
nor U29939 (N_29939,N_29636,N_29537);
or U29940 (N_29940,N_29626,N_29748);
or U29941 (N_29941,N_29602,N_29552);
nor U29942 (N_29942,N_29736,N_29713);
nor U29943 (N_29943,N_29674,N_29528);
nand U29944 (N_29944,N_29710,N_29651);
nor U29945 (N_29945,N_29568,N_29679);
or U29946 (N_29946,N_29620,N_29591);
or U29947 (N_29947,N_29548,N_29731);
nor U29948 (N_29948,N_29650,N_29542);
xor U29949 (N_29949,N_29691,N_29744);
nand U29950 (N_29950,N_29719,N_29502);
nor U29951 (N_29951,N_29547,N_29606);
or U29952 (N_29952,N_29539,N_29630);
and U29953 (N_29953,N_29519,N_29617);
xor U29954 (N_29954,N_29668,N_29727);
nand U29955 (N_29955,N_29625,N_29534);
nand U29956 (N_29956,N_29586,N_29744);
xnor U29957 (N_29957,N_29619,N_29585);
xor U29958 (N_29958,N_29519,N_29717);
or U29959 (N_29959,N_29625,N_29702);
nand U29960 (N_29960,N_29606,N_29665);
nor U29961 (N_29961,N_29743,N_29710);
and U29962 (N_29962,N_29508,N_29604);
and U29963 (N_29963,N_29633,N_29610);
nand U29964 (N_29964,N_29507,N_29654);
xnor U29965 (N_29965,N_29700,N_29633);
xor U29966 (N_29966,N_29626,N_29591);
or U29967 (N_29967,N_29727,N_29693);
nor U29968 (N_29968,N_29619,N_29582);
nor U29969 (N_29969,N_29605,N_29719);
or U29970 (N_29970,N_29683,N_29734);
xnor U29971 (N_29971,N_29572,N_29744);
or U29972 (N_29972,N_29581,N_29739);
nor U29973 (N_29973,N_29742,N_29681);
or U29974 (N_29974,N_29640,N_29654);
and U29975 (N_29975,N_29512,N_29667);
or U29976 (N_29976,N_29547,N_29627);
xor U29977 (N_29977,N_29722,N_29702);
xnor U29978 (N_29978,N_29679,N_29570);
and U29979 (N_29979,N_29562,N_29523);
nand U29980 (N_29980,N_29587,N_29666);
nor U29981 (N_29981,N_29552,N_29699);
or U29982 (N_29982,N_29677,N_29744);
nand U29983 (N_29983,N_29533,N_29600);
or U29984 (N_29984,N_29719,N_29558);
and U29985 (N_29985,N_29652,N_29603);
nor U29986 (N_29986,N_29697,N_29521);
and U29987 (N_29987,N_29507,N_29619);
nand U29988 (N_29988,N_29736,N_29541);
or U29989 (N_29989,N_29675,N_29612);
or U29990 (N_29990,N_29675,N_29683);
and U29991 (N_29991,N_29712,N_29578);
or U29992 (N_29992,N_29503,N_29545);
and U29993 (N_29993,N_29606,N_29679);
xnor U29994 (N_29994,N_29652,N_29591);
and U29995 (N_29995,N_29623,N_29680);
or U29996 (N_29996,N_29573,N_29521);
or U29997 (N_29997,N_29540,N_29554);
nand U29998 (N_29998,N_29703,N_29599);
xnor U29999 (N_29999,N_29748,N_29723);
or U30000 (N_30000,N_29844,N_29826);
or U30001 (N_30001,N_29927,N_29765);
nand U30002 (N_30002,N_29892,N_29984);
nor U30003 (N_30003,N_29950,N_29801);
nor U30004 (N_30004,N_29852,N_29949);
nand U30005 (N_30005,N_29754,N_29922);
nand U30006 (N_30006,N_29763,N_29916);
and U30007 (N_30007,N_29943,N_29799);
or U30008 (N_30008,N_29838,N_29815);
or U30009 (N_30009,N_29993,N_29920);
nand U30010 (N_30010,N_29829,N_29964);
or U30011 (N_30011,N_29785,N_29997);
or U30012 (N_30012,N_29759,N_29875);
and U30013 (N_30013,N_29860,N_29847);
nor U30014 (N_30014,N_29868,N_29986);
nor U30015 (N_30015,N_29784,N_29791);
or U30016 (N_30016,N_29930,N_29814);
or U30017 (N_30017,N_29774,N_29899);
or U30018 (N_30018,N_29770,N_29985);
nand U30019 (N_30019,N_29808,N_29960);
or U30020 (N_30020,N_29767,N_29775);
nand U30021 (N_30021,N_29809,N_29793);
and U30022 (N_30022,N_29863,N_29753);
or U30023 (N_30023,N_29810,N_29924);
or U30024 (N_30024,N_29836,N_29812);
and U30025 (N_30025,N_29976,N_29970);
and U30026 (N_30026,N_29796,N_29982);
nand U30027 (N_30027,N_29828,N_29777);
nor U30028 (N_30028,N_29848,N_29833);
and U30029 (N_30029,N_29932,N_29913);
nor U30030 (N_30030,N_29845,N_29968);
xor U30031 (N_30031,N_29764,N_29898);
nor U30032 (N_30032,N_29813,N_29840);
xnor U30033 (N_30033,N_29803,N_29837);
xor U30034 (N_30034,N_29937,N_29851);
nand U30035 (N_30035,N_29900,N_29945);
or U30036 (N_30036,N_29980,N_29965);
nor U30037 (N_30037,N_29839,N_29963);
nand U30038 (N_30038,N_29865,N_29832);
xnor U30039 (N_30039,N_29977,N_29905);
xor U30040 (N_30040,N_29907,N_29991);
or U30041 (N_30041,N_29972,N_29956);
and U30042 (N_30042,N_29842,N_29856);
xnor U30043 (N_30043,N_29923,N_29870);
nor U30044 (N_30044,N_29961,N_29798);
nand U30045 (N_30045,N_29885,N_29919);
or U30046 (N_30046,N_29896,N_29938);
nand U30047 (N_30047,N_29978,N_29953);
nand U30048 (N_30048,N_29756,N_29891);
nor U30049 (N_30049,N_29929,N_29989);
or U30050 (N_30050,N_29786,N_29918);
xnor U30051 (N_30051,N_29955,N_29797);
or U30052 (N_30052,N_29939,N_29926);
nand U30053 (N_30053,N_29792,N_29872);
nor U30054 (N_30054,N_29757,N_29768);
xor U30055 (N_30055,N_29951,N_29902);
or U30056 (N_30056,N_29879,N_29954);
and U30057 (N_30057,N_29794,N_29790);
nor U30058 (N_30058,N_29788,N_29958);
and U30059 (N_30059,N_29992,N_29800);
and U30060 (N_30060,N_29861,N_29822);
nor U30061 (N_30061,N_29874,N_29878);
nor U30062 (N_30062,N_29909,N_29987);
xor U30063 (N_30063,N_29967,N_29886);
nor U30064 (N_30064,N_29890,N_29947);
nor U30065 (N_30065,N_29928,N_29871);
xor U30066 (N_30066,N_29783,N_29787);
nor U30067 (N_30067,N_29771,N_29818);
and U30068 (N_30068,N_29883,N_29750);
and U30069 (N_30069,N_29975,N_29841);
nand U30070 (N_30070,N_29802,N_29855);
or U30071 (N_30071,N_29998,N_29912);
xor U30072 (N_30072,N_29867,N_29766);
nor U30073 (N_30073,N_29773,N_29859);
nor U30074 (N_30074,N_29897,N_29819);
nor U30075 (N_30075,N_29887,N_29911);
nor U30076 (N_30076,N_29877,N_29761);
xor U30077 (N_30077,N_29846,N_29880);
nor U30078 (N_30078,N_29906,N_29971);
nand U30079 (N_30079,N_29843,N_29864);
nor U30080 (N_30080,N_29959,N_29936);
or U30081 (N_30081,N_29853,N_29934);
nor U30082 (N_30082,N_29979,N_29941);
xor U30083 (N_30083,N_29769,N_29994);
nor U30084 (N_30084,N_29948,N_29857);
and U30085 (N_30085,N_29910,N_29895);
nor U30086 (N_30086,N_29944,N_29834);
or U30087 (N_30087,N_29805,N_29914);
xnor U30088 (N_30088,N_29946,N_29827);
xnor U30089 (N_30089,N_29940,N_29850);
nor U30090 (N_30090,N_29973,N_29917);
nand U30091 (N_30091,N_29760,N_29789);
xnor U30092 (N_30092,N_29933,N_29866);
or U30093 (N_30093,N_29882,N_29830);
or U30094 (N_30094,N_29888,N_29969);
xor U30095 (N_30095,N_29804,N_29903);
xor U30096 (N_30096,N_29981,N_29881);
nor U30097 (N_30097,N_29925,N_29901);
nor U30098 (N_30098,N_29893,N_29849);
and U30099 (N_30099,N_29889,N_29762);
xor U30100 (N_30100,N_29876,N_29996);
and U30101 (N_30101,N_29990,N_29780);
nor U30102 (N_30102,N_29781,N_29858);
or U30103 (N_30103,N_29904,N_29966);
or U30104 (N_30104,N_29962,N_29835);
xnor U30105 (N_30105,N_29999,N_29894);
nand U30106 (N_30106,N_29957,N_29807);
xor U30107 (N_30107,N_29873,N_29825);
and U30108 (N_30108,N_29824,N_29811);
nand U30109 (N_30109,N_29942,N_29816);
and U30110 (N_30110,N_29795,N_29823);
nor U30111 (N_30111,N_29806,N_29772);
nand U30112 (N_30112,N_29758,N_29782);
and U30113 (N_30113,N_29752,N_29778);
xor U30114 (N_30114,N_29751,N_29983);
xnor U30115 (N_30115,N_29935,N_29755);
nor U30116 (N_30116,N_29988,N_29908);
xor U30117 (N_30117,N_29884,N_29952);
and U30118 (N_30118,N_29974,N_29862);
and U30119 (N_30119,N_29820,N_29869);
and U30120 (N_30120,N_29995,N_29831);
or U30121 (N_30121,N_29931,N_29817);
nor U30122 (N_30122,N_29821,N_29921);
nor U30123 (N_30123,N_29854,N_29776);
nand U30124 (N_30124,N_29779,N_29915);
nor U30125 (N_30125,N_29898,N_29821);
and U30126 (N_30126,N_29987,N_29863);
or U30127 (N_30127,N_29828,N_29978);
or U30128 (N_30128,N_29834,N_29954);
and U30129 (N_30129,N_29994,N_29886);
nor U30130 (N_30130,N_29762,N_29791);
or U30131 (N_30131,N_29928,N_29791);
or U30132 (N_30132,N_29866,N_29816);
xor U30133 (N_30133,N_29899,N_29800);
and U30134 (N_30134,N_29963,N_29798);
nand U30135 (N_30135,N_29885,N_29947);
or U30136 (N_30136,N_29798,N_29777);
nor U30137 (N_30137,N_29803,N_29767);
and U30138 (N_30138,N_29998,N_29768);
nand U30139 (N_30139,N_29833,N_29812);
and U30140 (N_30140,N_29999,N_29992);
xnor U30141 (N_30141,N_29976,N_29952);
nand U30142 (N_30142,N_29946,N_29772);
nor U30143 (N_30143,N_29943,N_29782);
and U30144 (N_30144,N_29865,N_29765);
xnor U30145 (N_30145,N_29757,N_29894);
nor U30146 (N_30146,N_29791,N_29772);
or U30147 (N_30147,N_29800,N_29914);
nor U30148 (N_30148,N_29779,N_29970);
or U30149 (N_30149,N_29926,N_29963);
nand U30150 (N_30150,N_29900,N_29835);
xnor U30151 (N_30151,N_29928,N_29790);
nor U30152 (N_30152,N_29773,N_29861);
and U30153 (N_30153,N_29799,N_29852);
xor U30154 (N_30154,N_29751,N_29772);
nor U30155 (N_30155,N_29787,N_29898);
or U30156 (N_30156,N_29818,N_29900);
or U30157 (N_30157,N_29916,N_29780);
and U30158 (N_30158,N_29820,N_29997);
nor U30159 (N_30159,N_29802,N_29838);
nor U30160 (N_30160,N_29977,N_29849);
nand U30161 (N_30161,N_29970,N_29773);
or U30162 (N_30162,N_29944,N_29954);
and U30163 (N_30163,N_29824,N_29966);
and U30164 (N_30164,N_29939,N_29943);
nor U30165 (N_30165,N_29998,N_29930);
nor U30166 (N_30166,N_29811,N_29801);
xor U30167 (N_30167,N_29907,N_29955);
and U30168 (N_30168,N_29818,N_29940);
and U30169 (N_30169,N_29833,N_29805);
and U30170 (N_30170,N_29855,N_29878);
xnor U30171 (N_30171,N_29814,N_29967);
xnor U30172 (N_30172,N_29852,N_29803);
xnor U30173 (N_30173,N_29963,N_29962);
nand U30174 (N_30174,N_29907,N_29949);
and U30175 (N_30175,N_29954,N_29899);
and U30176 (N_30176,N_29860,N_29903);
nand U30177 (N_30177,N_29942,N_29925);
xor U30178 (N_30178,N_29798,N_29874);
and U30179 (N_30179,N_29762,N_29792);
and U30180 (N_30180,N_29875,N_29957);
nor U30181 (N_30181,N_29783,N_29865);
or U30182 (N_30182,N_29897,N_29803);
nor U30183 (N_30183,N_29929,N_29768);
or U30184 (N_30184,N_29843,N_29882);
xor U30185 (N_30185,N_29821,N_29864);
or U30186 (N_30186,N_29898,N_29852);
nand U30187 (N_30187,N_29969,N_29854);
and U30188 (N_30188,N_29857,N_29980);
or U30189 (N_30189,N_29909,N_29780);
xnor U30190 (N_30190,N_29812,N_29874);
or U30191 (N_30191,N_29876,N_29960);
and U30192 (N_30192,N_29914,N_29873);
nor U30193 (N_30193,N_29907,N_29954);
xnor U30194 (N_30194,N_29988,N_29880);
nor U30195 (N_30195,N_29884,N_29910);
and U30196 (N_30196,N_29881,N_29782);
nand U30197 (N_30197,N_29962,N_29862);
xnor U30198 (N_30198,N_29761,N_29845);
and U30199 (N_30199,N_29988,N_29992);
or U30200 (N_30200,N_29796,N_29996);
and U30201 (N_30201,N_29790,N_29939);
nor U30202 (N_30202,N_29869,N_29864);
or U30203 (N_30203,N_29984,N_29897);
xnor U30204 (N_30204,N_29946,N_29859);
nand U30205 (N_30205,N_29787,N_29779);
nand U30206 (N_30206,N_29983,N_29914);
or U30207 (N_30207,N_29982,N_29826);
xor U30208 (N_30208,N_29928,N_29864);
and U30209 (N_30209,N_29989,N_29774);
or U30210 (N_30210,N_29911,N_29783);
nor U30211 (N_30211,N_29892,N_29757);
nand U30212 (N_30212,N_29871,N_29832);
nand U30213 (N_30213,N_29950,N_29963);
or U30214 (N_30214,N_29807,N_29934);
and U30215 (N_30215,N_29833,N_29802);
xor U30216 (N_30216,N_29830,N_29877);
xnor U30217 (N_30217,N_29886,N_29906);
nor U30218 (N_30218,N_29845,N_29753);
nand U30219 (N_30219,N_29956,N_29925);
nor U30220 (N_30220,N_29986,N_29909);
and U30221 (N_30221,N_29769,N_29765);
nand U30222 (N_30222,N_29922,N_29936);
and U30223 (N_30223,N_29804,N_29814);
or U30224 (N_30224,N_29847,N_29922);
xnor U30225 (N_30225,N_29904,N_29796);
xor U30226 (N_30226,N_29817,N_29853);
or U30227 (N_30227,N_29844,N_29779);
nor U30228 (N_30228,N_29766,N_29993);
nor U30229 (N_30229,N_29819,N_29779);
or U30230 (N_30230,N_29899,N_29808);
xor U30231 (N_30231,N_29769,N_29954);
or U30232 (N_30232,N_29960,N_29980);
nand U30233 (N_30233,N_29964,N_29792);
and U30234 (N_30234,N_29900,N_29962);
and U30235 (N_30235,N_29962,N_29953);
and U30236 (N_30236,N_29901,N_29822);
nand U30237 (N_30237,N_29911,N_29920);
nand U30238 (N_30238,N_29929,N_29963);
and U30239 (N_30239,N_29778,N_29887);
and U30240 (N_30240,N_29766,N_29857);
nand U30241 (N_30241,N_29910,N_29913);
nand U30242 (N_30242,N_29933,N_29991);
xor U30243 (N_30243,N_29958,N_29963);
xnor U30244 (N_30244,N_29868,N_29978);
nand U30245 (N_30245,N_29925,N_29985);
nand U30246 (N_30246,N_29968,N_29870);
and U30247 (N_30247,N_29959,N_29853);
nand U30248 (N_30248,N_29775,N_29893);
nor U30249 (N_30249,N_29957,N_29867);
and U30250 (N_30250,N_30055,N_30119);
xnor U30251 (N_30251,N_30188,N_30133);
or U30252 (N_30252,N_30045,N_30073);
xnor U30253 (N_30253,N_30093,N_30123);
nand U30254 (N_30254,N_30075,N_30230);
or U30255 (N_30255,N_30134,N_30053);
and U30256 (N_30256,N_30097,N_30237);
and U30257 (N_30257,N_30038,N_30063);
xnor U30258 (N_30258,N_30044,N_30142);
or U30259 (N_30259,N_30013,N_30124);
xnor U30260 (N_30260,N_30215,N_30248);
nor U30261 (N_30261,N_30099,N_30004);
nor U30262 (N_30262,N_30014,N_30036);
nor U30263 (N_30263,N_30076,N_30191);
nor U30264 (N_30264,N_30209,N_30033);
or U30265 (N_30265,N_30087,N_30246);
or U30266 (N_30266,N_30072,N_30108);
nand U30267 (N_30267,N_30236,N_30005);
nand U30268 (N_30268,N_30154,N_30098);
xnor U30269 (N_30269,N_30159,N_30096);
nand U30270 (N_30270,N_30168,N_30051);
nor U30271 (N_30271,N_30083,N_30224);
nand U30272 (N_30272,N_30126,N_30177);
nor U30273 (N_30273,N_30143,N_30040);
and U30274 (N_30274,N_30222,N_30042);
and U30275 (N_30275,N_30104,N_30064);
and U30276 (N_30276,N_30232,N_30118);
nor U30277 (N_30277,N_30068,N_30181);
nor U30278 (N_30278,N_30012,N_30107);
and U30279 (N_30279,N_30060,N_30247);
xnor U30280 (N_30280,N_30028,N_30027);
nand U30281 (N_30281,N_30086,N_30009);
nor U30282 (N_30282,N_30214,N_30220);
or U30283 (N_30283,N_30217,N_30058);
or U30284 (N_30284,N_30178,N_30234);
nand U30285 (N_30285,N_30201,N_30231);
nand U30286 (N_30286,N_30106,N_30114);
or U30287 (N_30287,N_30113,N_30031);
or U30288 (N_30288,N_30037,N_30008);
xnor U30289 (N_30289,N_30092,N_30243);
xor U30290 (N_30290,N_30077,N_30155);
nor U30291 (N_30291,N_30228,N_30029);
and U30292 (N_30292,N_30039,N_30233);
or U30293 (N_30293,N_30199,N_30144);
xnor U30294 (N_30294,N_30015,N_30043);
xor U30295 (N_30295,N_30157,N_30059);
or U30296 (N_30296,N_30057,N_30111);
and U30297 (N_30297,N_30105,N_30207);
nor U30298 (N_30298,N_30078,N_30184);
nor U30299 (N_30299,N_30117,N_30235);
nor U30300 (N_30300,N_30206,N_30130);
nand U30301 (N_30301,N_30032,N_30100);
or U30302 (N_30302,N_30022,N_30164);
nor U30303 (N_30303,N_30035,N_30094);
nor U30304 (N_30304,N_30103,N_30085);
and U30305 (N_30305,N_30193,N_30244);
nand U30306 (N_30306,N_30054,N_30225);
nand U30307 (N_30307,N_30109,N_30186);
or U30308 (N_30308,N_30131,N_30041);
nor U30309 (N_30309,N_30125,N_30223);
nand U30310 (N_30310,N_30030,N_30192);
nor U30311 (N_30311,N_30166,N_30066);
nand U30312 (N_30312,N_30150,N_30172);
or U30313 (N_30313,N_30001,N_30180);
nand U30314 (N_30314,N_30091,N_30216);
and U30315 (N_30315,N_30148,N_30121);
nand U30316 (N_30316,N_30242,N_30149);
and U30317 (N_30317,N_30240,N_30046);
xnor U30318 (N_30318,N_30171,N_30019);
xnor U30319 (N_30319,N_30136,N_30218);
nor U30320 (N_30320,N_30175,N_30211);
xnor U30321 (N_30321,N_30081,N_30203);
or U30322 (N_30322,N_30056,N_30173);
and U30323 (N_30323,N_30003,N_30227);
and U30324 (N_30324,N_30146,N_30007);
nand U30325 (N_30325,N_30020,N_30048);
or U30326 (N_30326,N_30002,N_30205);
and U30327 (N_30327,N_30070,N_30151);
xor U30328 (N_30328,N_30069,N_30065);
nand U30329 (N_30329,N_30170,N_30132);
xor U30330 (N_30330,N_30129,N_30208);
nor U30331 (N_30331,N_30152,N_30116);
nand U30332 (N_30332,N_30017,N_30212);
xnor U30333 (N_30333,N_30011,N_30249);
xnor U30334 (N_30334,N_30153,N_30120);
or U30335 (N_30335,N_30052,N_30163);
and U30336 (N_30336,N_30145,N_30169);
xor U30337 (N_30337,N_30190,N_30101);
nor U30338 (N_30338,N_30139,N_30062);
xnor U30339 (N_30339,N_30161,N_30229);
nor U30340 (N_30340,N_30195,N_30194);
nor U30341 (N_30341,N_30082,N_30089);
and U30342 (N_30342,N_30174,N_30016);
or U30343 (N_30343,N_30219,N_30090);
and U30344 (N_30344,N_30115,N_30198);
and U30345 (N_30345,N_30200,N_30147);
and U30346 (N_30346,N_30138,N_30088);
nand U30347 (N_30347,N_30204,N_30182);
xor U30348 (N_30348,N_30238,N_30140);
and U30349 (N_30349,N_30245,N_30156);
nand U30350 (N_30350,N_30079,N_30025);
and U30351 (N_30351,N_30158,N_30102);
and U30352 (N_30352,N_30127,N_30095);
or U30353 (N_30353,N_30239,N_30135);
xor U30354 (N_30354,N_30185,N_30061);
nand U30355 (N_30355,N_30226,N_30084);
nand U30356 (N_30356,N_30024,N_30110);
or U30357 (N_30357,N_30034,N_30128);
xor U30358 (N_30358,N_30241,N_30197);
nor U30359 (N_30359,N_30141,N_30165);
nor U30360 (N_30360,N_30112,N_30049);
nor U30361 (N_30361,N_30196,N_30213);
nor U30362 (N_30362,N_30162,N_30026);
or U30363 (N_30363,N_30074,N_30176);
xnor U30364 (N_30364,N_30210,N_30080);
nor U30365 (N_30365,N_30122,N_30183);
nand U30366 (N_30366,N_30000,N_30023);
or U30367 (N_30367,N_30010,N_30202);
nor U30368 (N_30368,N_30067,N_30221);
nor U30369 (N_30369,N_30071,N_30189);
and U30370 (N_30370,N_30167,N_30018);
nor U30371 (N_30371,N_30021,N_30050);
and U30372 (N_30372,N_30187,N_30047);
nand U30373 (N_30373,N_30179,N_30160);
nand U30374 (N_30374,N_30137,N_30006);
nor U30375 (N_30375,N_30035,N_30058);
and U30376 (N_30376,N_30026,N_30245);
xor U30377 (N_30377,N_30003,N_30120);
and U30378 (N_30378,N_30195,N_30186);
nand U30379 (N_30379,N_30111,N_30086);
and U30380 (N_30380,N_30231,N_30090);
or U30381 (N_30381,N_30114,N_30217);
xnor U30382 (N_30382,N_30211,N_30185);
or U30383 (N_30383,N_30220,N_30168);
nor U30384 (N_30384,N_30147,N_30233);
or U30385 (N_30385,N_30026,N_30169);
nand U30386 (N_30386,N_30077,N_30167);
nor U30387 (N_30387,N_30201,N_30219);
nor U30388 (N_30388,N_30019,N_30055);
xor U30389 (N_30389,N_30152,N_30147);
xnor U30390 (N_30390,N_30059,N_30035);
nor U30391 (N_30391,N_30187,N_30144);
and U30392 (N_30392,N_30153,N_30236);
and U30393 (N_30393,N_30056,N_30206);
xnor U30394 (N_30394,N_30051,N_30034);
nor U30395 (N_30395,N_30080,N_30096);
xnor U30396 (N_30396,N_30049,N_30222);
nor U30397 (N_30397,N_30249,N_30036);
nor U30398 (N_30398,N_30230,N_30027);
or U30399 (N_30399,N_30015,N_30084);
and U30400 (N_30400,N_30062,N_30098);
and U30401 (N_30401,N_30023,N_30047);
nor U30402 (N_30402,N_30070,N_30226);
and U30403 (N_30403,N_30116,N_30008);
and U30404 (N_30404,N_30035,N_30233);
nand U30405 (N_30405,N_30148,N_30042);
nand U30406 (N_30406,N_30185,N_30159);
nand U30407 (N_30407,N_30019,N_30213);
nand U30408 (N_30408,N_30175,N_30130);
nand U30409 (N_30409,N_30183,N_30228);
or U30410 (N_30410,N_30227,N_30159);
or U30411 (N_30411,N_30128,N_30093);
xor U30412 (N_30412,N_30082,N_30196);
or U30413 (N_30413,N_30134,N_30157);
nor U30414 (N_30414,N_30002,N_30091);
nand U30415 (N_30415,N_30237,N_30229);
or U30416 (N_30416,N_30216,N_30008);
or U30417 (N_30417,N_30016,N_30136);
nor U30418 (N_30418,N_30136,N_30217);
xor U30419 (N_30419,N_30140,N_30177);
or U30420 (N_30420,N_30203,N_30037);
and U30421 (N_30421,N_30102,N_30055);
or U30422 (N_30422,N_30136,N_30073);
nor U30423 (N_30423,N_30200,N_30072);
and U30424 (N_30424,N_30241,N_30025);
nand U30425 (N_30425,N_30176,N_30106);
xnor U30426 (N_30426,N_30224,N_30030);
and U30427 (N_30427,N_30027,N_30133);
nor U30428 (N_30428,N_30026,N_30164);
nand U30429 (N_30429,N_30023,N_30073);
xnor U30430 (N_30430,N_30050,N_30154);
or U30431 (N_30431,N_30180,N_30039);
xor U30432 (N_30432,N_30013,N_30162);
xor U30433 (N_30433,N_30179,N_30223);
nand U30434 (N_30434,N_30055,N_30068);
xor U30435 (N_30435,N_30196,N_30057);
xor U30436 (N_30436,N_30020,N_30174);
and U30437 (N_30437,N_30033,N_30115);
nand U30438 (N_30438,N_30172,N_30030);
and U30439 (N_30439,N_30159,N_30089);
xnor U30440 (N_30440,N_30123,N_30101);
and U30441 (N_30441,N_30156,N_30036);
or U30442 (N_30442,N_30224,N_30168);
nand U30443 (N_30443,N_30121,N_30009);
xor U30444 (N_30444,N_30087,N_30155);
nand U30445 (N_30445,N_30180,N_30048);
xnor U30446 (N_30446,N_30097,N_30116);
nand U30447 (N_30447,N_30083,N_30129);
nor U30448 (N_30448,N_30174,N_30243);
xor U30449 (N_30449,N_30049,N_30233);
nor U30450 (N_30450,N_30145,N_30107);
and U30451 (N_30451,N_30236,N_30116);
nand U30452 (N_30452,N_30233,N_30074);
nor U30453 (N_30453,N_30058,N_30020);
nand U30454 (N_30454,N_30071,N_30098);
xor U30455 (N_30455,N_30090,N_30199);
and U30456 (N_30456,N_30231,N_30176);
xor U30457 (N_30457,N_30148,N_30109);
nor U30458 (N_30458,N_30055,N_30028);
nor U30459 (N_30459,N_30194,N_30081);
xnor U30460 (N_30460,N_30147,N_30109);
and U30461 (N_30461,N_30100,N_30191);
nand U30462 (N_30462,N_30032,N_30229);
nand U30463 (N_30463,N_30175,N_30074);
xor U30464 (N_30464,N_30039,N_30131);
nor U30465 (N_30465,N_30021,N_30034);
xor U30466 (N_30466,N_30035,N_30049);
and U30467 (N_30467,N_30189,N_30232);
and U30468 (N_30468,N_30167,N_30205);
nor U30469 (N_30469,N_30173,N_30091);
xor U30470 (N_30470,N_30132,N_30108);
nand U30471 (N_30471,N_30071,N_30138);
nor U30472 (N_30472,N_30001,N_30167);
xnor U30473 (N_30473,N_30062,N_30054);
and U30474 (N_30474,N_30009,N_30162);
and U30475 (N_30475,N_30164,N_30109);
nor U30476 (N_30476,N_30137,N_30184);
and U30477 (N_30477,N_30015,N_30111);
xnor U30478 (N_30478,N_30116,N_30223);
xnor U30479 (N_30479,N_30201,N_30095);
and U30480 (N_30480,N_30065,N_30014);
and U30481 (N_30481,N_30019,N_30130);
or U30482 (N_30482,N_30227,N_30083);
and U30483 (N_30483,N_30121,N_30161);
nand U30484 (N_30484,N_30126,N_30062);
nand U30485 (N_30485,N_30080,N_30170);
xnor U30486 (N_30486,N_30182,N_30078);
nand U30487 (N_30487,N_30159,N_30048);
nand U30488 (N_30488,N_30138,N_30244);
nand U30489 (N_30489,N_30133,N_30240);
xor U30490 (N_30490,N_30133,N_30083);
nand U30491 (N_30491,N_30206,N_30249);
nor U30492 (N_30492,N_30237,N_30061);
nor U30493 (N_30493,N_30240,N_30062);
and U30494 (N_30494,N_30230,N_30079);
and U30495 (N_30495,N_30225,N_30071);
nand U30496 (N_30496,N_30225,N_30101);
nor U30497 (N_30497,N_30180,N_30000);
xnor U30498 (N_30498,N_30105,N_30188);
nor U30499 (N_30499,N_30156,N_30243);
or U30500 (N_30500,N_30363,N_30351);
nor U30501 (N_30501,N_30388,N_30486);
nand U30502 (N_30502,N_30459,N_30410);
xor U30503 (N_30503,N_30330,N_30406);
and U30504 (N_30504,N_30342,N_30457);
and U30505 (N_30505,N_30321,N_30362);
and U30506 (N_30506,N_30372,N_30254);
and U30507 (N_30507,N_30313,N_30401);
xnor U30508 (N_30508,N_30380,N_30439);
xnor U30509 (N_30509,N_30304,N_30455);
nor U30510 (N_30510,N_30374,N_30443);
or U30511 (N_30511,N_30437,N_30408);
xor U30512 (N_30512,N_30349,N_30373);
xnor U30513 (N_30513,N_30463,N_30471);
nor U30514 (N_30514,N_30376,N_30293);
and U30515 (N_30515,N_30390,N_30440);
xnor U30516 (N_30516,N_30338,N_30283);
xor U30517 (N_30517,N_30354,N_30479);
or U30518 (N_30518,N_30447,N_30418);
nor U30519 (N_30519,N_30345,N_30493);
or U30520 (N_30520,N_30339,N_30287);
nand U30521 (N_30521,N_30465,N_30333);
and U30522 (N_30522,N_30475,N_30472);
and U30523 (N_30523,N_30485,N_30441);
and U30524 (N_30524,N_30424,N_30446);
or U30525 (N_30525,N_30312,N_30385);
nor U30526 (N_30526,N_30409,N_30488);
nand U30527 (N_30527,N_30365,N_30481);
nor U30528 (N_30528,N_30251,N_30497);
or U30529 (N_30529,N_30375,N_30477);
nand U30530 (N_30530,N_30297,N_30395);
or U30531 (N_30531,N_30429,N_30482);
nand U30532 (N_30532,N_30478,N_30270);
nand U30533 (N_30533,N_30266,N_30379);
nand U30534 (N_30534,N_30402,N_30296);
and U30535 (N_30535,N_30428,N_30267);
and U30536 (N_30536,N_30412,N_30259);
and U30537 (N_30537,N_30360,N_30343);
nand U30538 (N_30538,N_30417,N_30291);
nor U30539 (N_30539,N_30445,N_30290);
xnor U30540 (N_30540,N_30314,N_30265);
nand U30541 (N_30541,N_30277,N_30332);
and U30542 (N_30542,N_30299,N_30381);
xor U30543 (N_30543,N_30327,N_30444);
or U30544 (N_30544,N_30268,N_30498);
nand U30545 (N_30545,N_30423,N_30255);
and U30546 (N_30546,N_30377,N_30416);
xor U30547 (N_30547,N_30448,N_30495);
xor U30548 (N_30548,N_30367,N_30250);
and U30549 (N_30549,N_30334,N_30260);
nor U30550 (N_30550,N_30364,N_30425);
xnor U30551 (N_30551,N_30421,N_30355);
nand U30552 (N_30552,N_30326,N_30331);
or U30553 (N_30553,N_30308,N_30430);
xor U30554 (N_30554,N_30384,N_30294);
xor U30555 (N_30555,N_30269,N_30361);
xnor U30556 (N_30556,N_30352,N_30336);
and U30557 (N_30557,N_30398,N_30318);
nor U30558 (N_30558,N_30261,N_30278);
or U30559 (N_30559,N_30470,N_30257);
xnor U30560 (N_30560,N_30275,N_30407);
or U30561 (N_30561,N_30347,N_30289);
and U30562 (N_30562,N_30378,N_30382);
and U30563 (N_30563,N_30458,N_30391);
nor U30564 (N_30564,N_30434,N_30264);
or U30565 (N_30565,N_30285,N_30311);
or U30566 (N_30566,N_30274,N_30263);
xor U30567 (N_30567,N_30344,N_30483);
nand U30568 (N_30568,N_30328,N_30348);
nor U30569 (N_30569,N_30282,N_30325);
or U30570 (N_30570,N_30281,N_30252);
nand U30571 (N_30571,N_30442,N_30403);
and U30572 (N_30572,N_30435,N_30492);
and U30573 (N_30573,N_30438,N_30490);
and U30574 (N_30574,N_30366,N_30394);
nand U30575 (N_30575,N_30419,N_30451);
or U30576 (N_30576,N_30272,N_30397);
nand U30577 (N_30577,N_30337,N_30454);
or U30578 (N_30578,N_30487,N_30316);
or U30579 (N_30579,N_30273,N_30309);
xnor U30580 (N_30580,N_30306,N_30358);
nor U30581 (N_30581,N_30370,N_30473);
and U30582 (N_30582,N_30399,N_30340);
or U30583 (N_30583,N_30307,N_30284);
or U30584 (N_30584,N_30460,N_30357);
nand U30585 (N_30585,N_30292,N_30324);
xor U30586 (N_30586,N_30303,N_30420);
or U30587 (N_30587,N_30298,N_30484);
or U30588 (N_30588,N_30393,N_30315);
xor U30589 (N_30589,N_30405,N_30280);
xor U30590 (N_30590,N_30414,N_30301);
nand U30591 (N_30591,N_30392,N_30422);
nand U30592 (N_30592,N_30258,N_30323);
xnor U30593 (N_30593,N_30279,N_30288);
and U30594 (N_30594,N_30300,N_30496);
nand U30595 (N_30595,N_30453,N_30413);
and U30596 (N_30596,N_30415,N_30353);
xnor U30597 (N_30597,N_30461,N_30356);
and U30598 (N_30598,N_30489,N_30368);
or U30599 (N_30599,N_30383,N_30295);
or U30600 (N_30600,N_30286,N_30427);
or U30601 (N_30601,N_30411,N_30494);
nor U30602 (N_30602,N_30386,N_30404);
nor U30603 (N_30603,N_30320,N_30400);
nor U30604 (N_30604,N_30253,N_30317);
xor U30605 (N_30605,N_30359,N_30469);
or U30606 (N_30606,N_30346,N_30462);
xnor U30607 (N_30607,N_30256,N_30450);
xnor U30608 (N_30608,N_30431,N_30369);
nor U30609 (N_30609,N_30341,N_30466);
or U30610 (N_30610,N_30319,N_30262);
nand U30611 (N_30611,N_30452,N_30449);
xnor U30612 (N_30612,N_30456,N_30436);
or U30613 (N_30613,N_30387,N_30467);
or U30614 (N_30614,N_30480,N_30305);
or U30615 (N_30615,N_30389,N_30371);
nor U30616 (N_30616,N_30350,N_30271);
and U30617 (N_30617,N_30322,N_30302);
xnor U30618 (N_30618,N_30432,N_30433);
nand U30619 (N_30619,N_30276,N_30491);
or U30620 (N_30620,N_30329,N_30499);
xor U30621 (N_30621,N_30474,N_30310);
nand U30622 (N_30622,N_30426,N_30396);
nor U30623 (N_30623,N_30464,N_30476);
nand U30624 (N_30624,N_30468,N_30335);
and U30625 (N_30625,N_30482,N_30353);
nand U30626 (N_30626,N_30264,N_30454);
and U30627 (N_30627,N_30384,N_30394);
or U30628 (N_30628,N_30388,N_30386);
and U30629 (N_30629,N_30267,N_30430);
nand U30630 (N_30630,N_30448,N_30485);
or U30631 (N_30631,N_30368,N_30435);
xor U30632 (N_30632,N_30397,N_30451);
and U30633 (N_30633,N_30357,N_30326);
or U30634 (N_30634,N_30311,N_30251);
xnor U30635 (N_30635,N_30454,N_30427);
or U30636 (N_30636,N_30352,N_30366);
xnor U30637 (N_30637,N_30451,N_30320);
nor U30638 (N_30638,N_30342,N_30448);
and U30639 (N_30639,N_30353,N_30335);
or U30640 (N_30640,N_30328,N_30353);
xor U30641 (N_30641,N_30332,N_30286);
nand U30642 (N_30642,N_30427,N_30364);
or U30643 (N_30643,N_30412,N_30422);
or U30644 (N_30644,N_30463,N_30309);
nor U30645 (N_30645,N_30372,N_30255);
and U30646 (N_30646,N_30349,N_30413);
nor U30647 (N_30647,N_30370,N_30319);
nand U30648 (N_30648,N_30469,N_30277);
nor U30649 (N_30649,N_30321,N_30496);
xnor U30650 (N_30650,N_30250,N_30290);
xor U30651 (N_30651,N_30458,N_30250);
xor U30652 (N_30652,N_30396,N_30428);
nand U30653 (N_30653,N_30424,N_30358);
nor U30654 (N_30654,N_30250,N_30311);
xor U30655 (N_30655,N_30499,N_30363);
and U30656 (N_30656,N_30464,N_30288);
or U30657 (N_30657,N_30445,N_30465);
and U30658 (N_30658,N_30491,N_30449);
or U30659 (N_30659,N_30451,N_30363);
and U30660 (N_30660,N_30254,N_30303);
and U30661 (N_30661,N_30322,N_30329);
or U30662 (N_30662,N_30341,N_30292);
and U30663 (N_30663,N_30413,N_30455);
nor U30664 (N_30664,N_30294,N_30462);
and U30665 (N_30665,N_30282,N_30347);
and U30666 (N_30666,N_30404,N_30494);
xnor U30667 (N_30667,N_30289,N_30358);
xnor U30668 (N_30668,N_30313,N_30431);
or U30669 (N_30669,N_30391,N_30362);
nand U30670 (N_30670,N_30319,N_30488);
and U30671 (N_30671,N_30360,N_30298);
and U30672 (N_30672,N_30444,N_30268);
xor U30673 (N_30673,N_30270,N_30269);
or U30674 (N_30674,N_30426,N_30436);
xnor U30675 (N_30675,N_30314,N_30491);
and U30676 (N_30676,N_30343,N_30318);
and U30677 (N_30677,N_30464,N_30336);
or U30678 (N_30678,N_30281,N_30259);
and U30679 (N_30679,N_30390,N_30417);
and U30680 (N_30680,N_30329,N_30380);
nand U30681 (N_30681,N_30270,N_30277);
and U30682 (N_30682,N_30333,N_30399);
xnor U30683 (N_30683,N_30298,N_30261);
xor U30684 (N_30684,N_30278,N_30469);
nand U30685 (N_30685,N_30397,N_30333);
or U30686 (N_30686,N_30290,N_30378);
nand U30687 (N_30687,N_30402,N_30483);
or U30688 (N_30688,N_30284,N_30493);
xnor U30689 (N_30689,N_30370,N_30285);
and U30690 (N_30690,N_30331,N_30402);
nor U30691 (N_30691,N_30264,N_30301);
nor U30692 (N_30692,N_30447,N_30305);
or U30693 (N_30693,N_30455,N_30316);
or U30694 (N_30694,N_30251,N_30483);
xor U30695 (N_30695,N_30492,N_30463);
nor U30696 (N_30696,N_30420,N_30314);
nor U30697 (N_30697,N_30328,N_30367);
or U30698 (N_30698,N_30447,N_30457);
or U30699 (N_30699,N_30458,N_30494);
nand U30700 (N_30700,N_30449,N_30461);
nor U30701 (N_30701,N_30253,N_30376);
or U30702 (N_30702,N_30264,N_30490);
or U30703 (N_30703,N_30450,N_30266);
and U30704 (N_30704,N_30329,N_30303);
xnor U30705 (N_30705,N_30331,N_30364);
xor U30706 (N_30706,N_30426,N_30295);
or U30707 (N_30707,N_30287,N_30448);
and U30708 (N_30708,N_30261,N_30459);
nor U30709 (N_30709,N_30321,N_30438);
nor U30710 (N_30710,N_30362,N_30312);
nor U30711 (N_30711,N_30359,N_30308);
nand U30712 (N_30712,N_30492,N_30260);
nor U30713 (N_30713,N_30278,N_30479);
xor U30714 (N_30714,N_30323,N_30273);
and U30715 (N_30715,N_30409,N_30259);
nand U30716 (N_30716,N_30343,N_30471);
nor U30717 (N_30717,N_30484,N_30416);
and U30718 (N_30718,N_30337,N_30348);
nor U30719 (N_30719,N_30250,N_30409);
nand U30720 (N_30720,N_30283,N_30332);
xor U30721 (N_30721,N_30309,N_30460);
and U30722 (N_30722,N_30327,N_30362);
and U30723 (N_30723,N_30470,N_30288);
xnor U30724 (N_30724,N_30347,N_30388);
or U30725 (N_30725,N_30285,N_30317);
or U30726 (N_30726,N_30415,N_30453);
nand U30727 (N_30727,N_30463,N_30268);
and U30728 (N_30728,N_30457,N_30391);
nand U30729 (N_30729,N_30387,N_30255);
nand U30730 (N_30730,N_30368,N_30338);
nor U30731 (N_30731,N_30334,N_30375);
nor U30732 (N_30732,N_30280,N_30474);
xor U30733 (N_30733,N_30417,N_30490);
and U30734 (N_30734,N_30492,N_30346);
nor U30735 (N_30735,N_30379,N_30390);
nand U30736 (N_30736,N_30304,N_30463);
xor U30737 (N_30737,N_30334,N_30451);
nand U30738 (N_30738,N_30285,N_30310);
and U30739 (N_30739,N_30363,N_30276);
nor U30740 (N_30740,N_30297,N_30380);
nand U30741 (N_30741,N_30313,N_30367);
or U30742 (N_30742,N_30285,N_30298);
nor U30743 (N_30743,N_30341,N_30445);
or U30744 (N_30744,N_30285,N_30441);
nand U30745 (N_30745,N_30402,N_30263);
nand U30746 (N_30746,N_30454,N_30281);
and U30747 (N_30747,N_30451,N_30367);
or U30748 (N_30748,N_30392,N_30430);
or U30749 (N_30749,N_30301,N_30483);
nor U30750 (N_30750,N_30740,N_30557);
and U30751 (N_30751,N_30595,N_30569);
xor U30752 (N_30752,N_30673,N_30598);
nand U30753 (N_30753,N_30702,N_30577);
nor U30754 (N_30754,N_30642,N_30564);
and U30755 (N_30755,N_30527,N_30678);
nor U30756 (N_30756,N_30713,N_30668);
nor U30757 (N_30757,N_30709,N_30622);
or U30758 (N_30758,N_30742,N_30609);
nand U30759 (N_30759,N_30525,N_30655);
and U30760 (N_30760,N_30591,N_30541);
nor U30761 (N_30761,N_30672,N_30546);
nor U30762 (N_30762,N_30719,N_30718);
and U30763 (N_30763,N_30539,N_30634);
or U30764 (N_30764,N_30679,N_30640);
nand U30765 (N_30765,N_30682,N_30728);
and U30766 (N_30766,N_30532,N_30657);
and U30767 (N_30767,N_30638,N_30608);
xor U30768 (N_30768,N_30524,N_30544);
or U30769 (N_30769,N_30739,N_30665);
nor U30770 (N_30770,N_30641,N_30732);
and U30771 (N_30771,N_30573,N_30664);
and U30772 (N_30772,N_30612,N_30552);
nand U30773 (N_30773,N_30645,N_30670);
and U30774 (N_30774,N_30725,N_30520);
nor U30775 (N_30775,N_30736,N_30734);
xor U30776 (N_30776,N_30536,N_30695);
nand U30777 (N_30777,N_30688,N_30528);
nor U30778 (N_30778,N_30721,N_30523);
or U30779 (N_30779,N_30731,N_30511);
and U30780 (N_30780,N_30667,N_30508);
and U30781 (N_30781,N_30716,N_30547);
nand U30782 (N_30782,N_30626,N_30749);
or U30783 (N_30783,N_30677,N_30554);
nand U30784 (N_30784,N_30733,N_30606);
xnor U30785 (N_30785,N_30637,N_30601);
and U30786 (N_30786,N_30644,N_30654);
nand U30787 (N_30787,N_30616,N_30540);
xnor U30788 (N_30788,N_30694,N_30555);
nor U30789 (N_30789,N_30636,N_30561);
nor U30790 (N_30790,N_30572,N_30615);
nand U30791 (N_30791,N_30576,N_30501);
nand U30792 (N_30792,N_30617,N_30559);
and U30793 (N_30793,N_30549,N_30747);
nand U30794 (N_30794,N_30723,N_30610);
xnor U30795 (N_30795,N_30521,N_30744);
xnor U30796 (N_30796,N_30538,N_30701);
and U30797 (N_30797,N_30628,N_30659);
and U30798 (N_30798,N_30669,N_30696);
xnor U30799 (N_30799,N_30568,N_30565);
xor U30800 (N_30800,N_30737,N_30588);
xor U30801 (N_30801,N_30652,N_30602);
or U30802 (N_30802,N_30711,N_30522);
and U30803 (N_30803,N_30727,N_30579);
nor U30804 (N_30804,N_30666,N_30560);
or U30805 (N_30805,N_30745,N_30593);
xnor U30806 (N_30806,N_30624,N_30629);
nor U30807 (N_30807,N_30648,N_30699);
and U30808 (N_30808,N_30684,N_30708);
and U30809 (N_30809,N_30597,N_30563);
nor U30810 (N_30810,N_30605,N_30510);
or U30811 (N_30811,N_30720,N_30726);
or U30812 (N_30812,N_30551,N_30611);
and U30813 (N_30813,N_30643,N_30505);
nor U30814 (N_30814,N_30681,N_30604);
nor U30815 (N_30815,N_30574,N_30542);
or U30816 (N_30816,N_30633,N_30550);
xnor U30817 (N_30817,N_30509,N_30500);
and U30818 (N_30818,N_30582,N_30571);
nand U30819 (N_30819,N_30594,N_30515);
xnor U30820 (N_30820,N_30558,N_30548);
or U30821 (N_30821,N_30712,N_30599);
or U30822 (N_30822,N_30502,N_30683);
nand U30823 (N_30823,N_30623,N_30537);
and U30824 (N_30824,N_30639,N_30738);
or U30825 (N_30825,N_30556,N_30661);
xnor U30826 (N_30826,N_30580,N_30647);
nand U30827 (N_30827,N_30578,N_30715);
xnor U30828 (N_30828,N_30656,N_30596);
nor U30829 (N_30829,N_30735,N_30586);
nand U30830 (N_30830,N_30675,N_30706);
nand U30831 (N_30831,N_30503,N_30660);
or U30832 (N_30832,N_30512,N_30704);
nand U30833 (N_30833,N_30632,N_30685);
nor U30834 (N_30834,N_30693,N_30590);
nand U30835 (N_30835,N_30692,N_30553);
xnor U30836 (N_30836,N_30630,N_30651);
nand U30837 (N_30837,N_30627,N_30662);
and U30838 (N_30838,N_30585,N_30671);
xor U30839 (N_30839,N_30631,N_30589);
or U30840 (N_30840,N_30545,N_30587);
nand U30841 (N_30841,N_30575,N_30618);
or U30842 (N_30842,N_30698,N_30543);
or U30843 (N_30843,N_30741,N_30570);
xor U30844 (N_30844,N_30613,N_30748);
xnor U30845 (N_30845,N_30707,N_30583);
or U30846 (N_30846,N_30506,N_30746);
nand U30847 (N_30847,N_30680,N_30689);
nor U30848 (N_30848,N_30619,N_30722);
nand U30849 (N_30849,N_30530,N_30729);
nor U30850 (N_30850,N_30690,N_30566);
nand U30851 (N_30851,N_30691,N_30603);
or U30852 (N_30852,N_30517,N_30653);
xnor U30853 (N_30853,N_30534,N_30529);
and U30854 (N_30854,N_30650,N_30533);
or U30855 (N_30855,N_30562,N_30676);
nand U30856 (N_30856,N_30620,N_30687);
nand U30857 (N_30857,N_30700,N_30514);
or U30858 (N_30858,N_30710,N_30519);
and U30859 (N_30859,N_30625,N_30614);
xor U30860 (N_30860,N_30516,N_30658);
and U30861 (N_30861,N_30663,N_30581);
xor U30862 (N_30862,N_30607,N_30535);
and U30863 (N_30863,N_30724,N_30526);
xor U30864 (N_30864,N_30567,N_30686);
nor U30865 (N_30865,N_30518,N_30705);
xor U30866 (N_30866,N_30674,N_30513);
nand U30867 (N_30867,N_30649,N_30714);
xor U30868 (N_30868,N_30743,N_30504);
or U30869 (N_30869,N_30531,N_30584);
or U30870 (N_30870,N_30592,N_30621);
or U30871 (N_30871,N_30507,N_30697);
nor U30872 (N_30872,N_30730,N_30717);
nand U30873 (N_30873,N_30646,N_30600);
xnor U30874 (N_30874,N_30703,N_30635);
and U30875 (N_30875,N_30748,N_30539);
xor U30876 (N_30876,N_30697,N_30593);
or U30877 (N_30877,N_30571,N_30718);
or U30878 (N_30878,N_30525,N_30569);
nor U30879 (N_30879,N_30604,N_30689);
nand U30880 (N_30880,N_30631,N_30500);
nor U30881 (N_30881,N_30717,N_30687);
xnor U30882 (N_30882,N_30709,N_30507);
nor U30883 (N_30883,N_30637,N_30558);
and U30884 (N_30884,N_30607,N_30614);
or U30885 (N_30885,N_30575,N_30673);
xor U30886 (N_30886,N_30635,N_30624);
and U30887 (N_30887,N_30636,N_30525);
nor U30888 (N_30888,N_30637,N_30740);
nor U30889 (N_30889,N_30603,N_30682);
xnor U30890 (N_30890,N_30710,N_30676);
or U30891 (N_30891,N_30605,N_30598);
nor U30892 (N_30892,N_30689,N_30561);
xor U30893 (N_30893,N_30726,N_30575);
or U30894 (N_30894,N_30744,N_30651);
or U30895 (N_30895,N_30551,N_30563);
xnor U30896 (N_30896,N_30734,N_30567);
or U30897 (N_30897,N_30501,N_30675);
or U30898 (N_30898,N_30673,N_30736);
nand U30899 (N_30899,N_30505,N_30601);
and U30900 (N_30900,N_30701,N_30501);
or U30901 (N_30901,N_30564,N_30541);
and U30902 (N_30902,N_30605,N_30726);
nand U30903 (N_30903,N_30676,N_30711);
nor U30904 (N_30904,N_30574,N_30537);
nand U30905 (N_30905,N_30644,N_30690);
or U30906 (N_30906,N_30549,N_30648);
nor U30907 (N_30907,N_30642,N_30638);
and U30908 (N_30908,N_30516,N_30644);
nor U30909 (N_30909,N_30681,N_30579);
and U30910 (N_30910,N_30662,N_30544);
nor U30911 (N_30911,N_30655,N_30717);
or U30912 (N_30912,N_30592,N_30509);
or U30913 (N_30913,N_30699,N_30511);
or U30914 (N_30914,N_30533,N_30679);
nand U30915 (N_30915,N_30747,N_30743);
nand U30916 (N_30916,N_30745,N_30626);
xor U30917 (N_30917,N_30686,N_30556);
or U30918 (N_30918,N_30710,N_30540);
or U30919 (N_30919,N_30539,N_30680);
xor U30920 (N_30920,N_30748,N_30746);
nand U30921 (N_30921,N_30545,N_30678);
or U30922 (N_30922,N_30694,N_30614);
nor U30923 (N_30923,N_30698,N_30736);
or U30924 (N_30924,N_30620,N_30542);
nand U30925 (N_30925,N_30572,N_30566);
xnor U30926 (N_30926,N_30684,N_30552);
and U30927 (N_30927,N_30513,N_30509);
xor U30928 (N_30928,N_30612,N_30722);
or U30929 (N_30929,N_30677,N_30512);
nand U30930 (N_30930,N_30517,N_30616);
or U30931 (N_30931,N_30527,N_30547);
nand U30932 (N_30932,N_30677,N_30580);
and U30933 (N_30933,N_30574,N_30573);
nor U30934 (N_30934,N_30611,N_30702);
xor U30935 (N_30935,N_30630,N_30644);
xnor U30936 (N_30936,N_30732,N_30519);
xnor U30937 (N_30937,N_30536,N_30676);
xor U30938 (N_30938,N_30633,N_30697);
nand U30939 (N_30939,N_30568,N_30564);
nand U30940 (N_30940,N_30506,N_30641);
or U30941 (N_30941,N_30667,N_30649);
nand U30942 (N_30942,N_30726,N_30610);
nor U30943 (N_30943,N_30513,N_30632);
nor U30944 (N_30944,N_30687,N_30661);
xnor U30945 (N_30945,N_30639,N_30645);
nor U30946 (N_30946,N_30599,N_30668);
nor U30947 (N_30947,N_30621,N_30526);
or U30948 (N_30948,N_30576,N_30654);
and U30949 (N_30949,N_30690,N_30570);
nand U30950 (N_30950,N_30704,N_30501);
nor U30951 (N_30951,N_30545,N_30675);
nor U30952 (N_30952,N_30599,N_30553);
nand U30953 (N_30953,N_30556,N_30544);
and U30954 (N_30954,N_30503,N_30564);
nand U30955 (N_30955,N_30580,N_30663);
nand U30956 (N_30956,N_30579,N_30653);
nor U30957 (N_30957,N_30676,N_30677);
or U30958 (N_30958,N_30626,N_30580);
or U30959 (N_30959,N_30748,N_30710);
and U30960 (N_30960,N_30708,N_30623);
nand U30961 (N_30961,N_30725,N_30655);
or U30962 (N_30962,N_30678,N_30532);
nor U30963 (N_30963,N_30740,N_30512);
nand U30964 (N_30964,N_30622,N_30676);
and U30965 (N_30965,N_30560,N_30640);
or U30966 (N_30966,N_30631,N_30529);
nor U30967 (N_30967,N_30503,N_30727);
and U30968 (N_30968,N_30749,N_30624);
nor U30969 (N_30969,N_30743,N_30528);
or U30970 (N_30970,N_30695,N_30603);
xor U30971 (N_30971,N_30625,N_30510);
or U30972 (N_30972,N_30690,N_30605);
xor U30973 (N_30973,N_30725,N_30524);
or U30974 (N_30974,N_30520,N_30584);
nor U30975 (N_30975,N_30636,N_30646);
xor U30976 (N_30976,N_30565,N_30666);
xor U30977 (N_30977,N_30576,N_30626);
nand U30978 (N_30978,N_30655,N_30646);
and U30979 (N_30979,N_30728,N_30649);
and U30980 (N_30980,N_30526,N_30660);
xnor U30981 (N_30981,N_30601,N_30580);
xnor U30982 (N_30982,N_30672,N_30670);
nand U30983 (N_30983,N_30684,N_30541);
and U30984 (N_30984,N_30526,N_30744);
xnor U30985 (N_30985,N_30731,N_30659);
or U30986 (N_30986,N_30578,N_30699);
and U30987 (N_30987,N_30738,N_30503);
or U30988 (N_30988,N_30657,N_30649);
nand U30989 (N_30989,N_30592,N_30692);
or U30990 (N_30990,N_30731,N_30502);
or U30991 (N_30991,N_30500,N_30722);
nand U30992 (N_30992,N_30714,N_30644);
nand U30993 (N_30993,N_30612,N_30745);
and U30994 (N_30994,N_30515,N_30707);
xnor U30995 (N_30995,N_30574,N_30673);
or U30996 (N_30996,N_30535,N_30576);
and U30997 (N_30997,N_30591,N_30738);
nor U30998 (N_30998,N_30621,N_30693);
xor U30999 (N_30999,N_30559,N_30732);
xnor U31000 (N_31000,N_30820,N_30953);
and U31001 (N_31001,N_30802,N_30851);
or U31002 (N_31002,N_30833,N_30893);
nand U31003 (N_31003,N_30843,N_30780);
nor U31004 (N_31004,N_30970,N_30862);
and U31005 (N_31005,N_30788,N_30899);
nand U31006 (N_31006,N_30954,N_30785);
nand U31007 (N_31007,N_30762,N_30921);
nor U31008 (N_31008,N_30922,N_30907);
or U31009 (N_31009,N_30823,N_30783);
nor U31010 (N_31010,N_30885,N_30772);
or U31011 (N_31011,N_30806,N_30997);
and U31012 (N_31012,N_30863,N_30972);
xor U31013 (N_31013,N_30965,N_30886);
or U31014 (N_31014,N_30926,N_30935);
and U31015 (N_31015,N_30878,N_30958);
nor U31016 (N_31016,N_30937,N_30829);
nor U31017 (N_31017,N_30795,N_30966);
or U31018 (N_31018,N_30944,N_30846);
xor U31019 (N_31019,N_30969,N_30912);
or U31020 (N_31020,N_30776,N_30987);
nand U31021 (N_31021,N_30955,N_30765);
and U31022 (N_31022,N_30978,N_30766);
and U31023 (N_31023,N_30801,N_30930);
nor U31024 (N_31024,N_30750,N_30857);
xnor U31025 (N_31025,N_30946,N_30814);
and U31026 (N_31026,N_30928,N_30852);
and U31027 (N_31027,N_30960,N_30841);
nor U31028 (N_31028,N_30971,N_30764);
nor U31029 (N_31029,N_30993,N_30781);
nand U31030 (N_31030,N_30932,N_30901);
or U31031 (N_31031,N_30821,N_30844);
and U31032 (N_31032,N_30879,N_30964);
nor U31033 (N_31033,N_30904,N_30819);
and U31034 (N_31034,N_30995,N_30824);
xnor U31035 (N_31035,N_30837,N_30870);
nor U31036 (N_31036,N_30810,N_30991);
and U31037 (N_31037,N_30790,N_30822);
or U31038 (N_31038,N_30897,N_30865);
and U31039 (N_31039,N_30962,N_30916);
nor U31040 (N_31040,N_30871,N_30873);
and U31041 (N_31041,N_30992,N_30891);
nand U31042 (N_31042,N_30920,N_30890);
xnor U31043 (N_31043,N_30805,N_30753);
nand U31044 (N_31044,N_30976,N_30797);
or U31045 (N_31045,N_30763,N_30784);
xnor U31046 (N_31046,N_30791,N_30812);
xor U31047 (N_31047,N_30798,N_30842);
nor U31048 (N_31048,N_30799,N_30792);
xor U31049 (N_31049,N_30939,N_30840);
nand U31050 (N_31050,N_30982,N_30758);
or U31051 (N_31051,N_30867,N_30881);
and U31052 (N_31052,N_30945,N_30773);
or U31053 (N_31053,N_30918,N_30914);
or U31054 (N_31054,N_30817,N_30884);
xnor U31055 (N_31055,N_30796,N_30818);
and U31056 (N_31056,N_30975,N_30850);
xnor U31057 (N_31057,N_30900,N_30999);
xnor U31058 (N_31058,N_30883,N_30950);
and U31059 (N_31059,N_30775,N_30808);
and U31060 (N_31060,N_30895,N_30880);
nor U31061 (N_31061,N_30752,N_30756);
xor U31062 (N_31062,N_30830,N_30777);
nor U31063 (N_31063,N_30967,N_30787);
or U31064 (N_31064,N_30770,N_30809);
and U31065 (N_31065,N_30915,N_30835);
nand U31066 (N_31066,N_30754,N_30858);
or U31067 (N_31067,N_30898,N_30888);
nor U31068 (N_31068,N_30959,N_30917);
and U31069 (N_31069,N_30941,N_30910);
or U31070 (N_31070,N_30866,N_30998);
xnor U31071 (N_31071,N_30903,N_30927);
and U31072 (N_31072,N_30789,N_30760);
xnor U31073 (N_31073,N_30925,N_30936);
xnor U31074 (N_31074,N_30848,N_30834);
xnor U31075 (N_31075,N_30948,N_30909);
or U31076 (N_31076,N_30827,N_30767);
xor U31077 (N_31077,N_30905,N_30815);
or U31078 (N_31078,N_30892,N_30940);
nand U31079 (N_31079,N_30952,N_30751);
or U31080 (N_31080,N_30874,N_30919);
nand U31081 (N_31081,N_30807,N_30872);
xor U31082 (N_31082,N_30831,N_30942);
or U31083 (N_31083,N_30911,N_30856);
nor U31084 (N_31084,N_30906,N_30968);
and U31085 (N_31085,N_30839,N_30804);
nand U31086 (N_31086,N_30786,N_30803);
or U31087 (N_31087,N_30813,N_30882);
nor U31088 (N_31088,N_30794,N_30951);
or U31089 (N_31089,N_30961,N_30908);
xor U31090 (N_31090,N_30868,N_30949);
nor U31091 (N_31091,N_30769,N_30887);
nand U31092 (N_31092,N_30986,N_30826);
xor U31093 (N_31093,N_30838,N_30990);
xnor U31094 (N_31094,N_30923,N_30913);
nand U31095 (N_31095,N_30793,N_30861);
and U31096 (N_31096,N_30979,N_30779);
and U31097 (N_31097,N_30934,N_30931);
or U31098 (N_31098,N_30855,N_30778);
and U31099 (N_31099,N_30980,N_30973);
nand U31100 (N_31100,N_30825,N_30875);
nor U31101 (N_31101,N_30994,N_30877);
and U31102 (N_31102,N_30947,N_30759);
or U31103 (N_31103,N_30782,N_30860);
xor U31104 (N_31104,N_30984,N_30774);
or U31105 (N_31105,N_30956,N_30963);
xnor U31106 (N_31106,N_30853,N_30988);
or U31107 (N_31107,N_30983,N_30889);
nor U31108 (N_31108,N_30876,N_30989);
or U31109 (N_31109,N_30938,N_30996);
nand U31110 (N_31110,N_30832,N_30836);
and U31111 (N_31111,N_30757,N_30864);
nand U31112 (N_31112,N_30985,N_30771);
or U31113 (N_31113,N_30847,N_30924);
and U31114 (N_31114,N_30929,N_30800);
and U31115 (N_31115,N_30977,N_30894);
nor U31116 (N_31116,N_30761,N_30974);
nor U31117 (N_31117,N_30849,N_30768);
and U31118 (N_31118,N_30859,N_30811);
xor U31119 (N_31119,N_30755,N_30854);
or U31120 (N_31120,N_30943,N_30869);
and U31121 (N_31121,N_30957,N_30896);
nand U31122 (N_31122,N_30981,N_30845);
nand U31123 (N_31123,N_30816,N_30828);
nor U31124 (N_31124,N_30933,N_30902);
xor U31125 (N_31125,N_30852,N_30794);
and U31126 (N_31126,N_30884,N_30972);
nand U31127 (N_31127,N_30782,N_30904);
xor U31128 (N_31128,N_30854,N_30959);
nand U31129 (N_31129,N_30820,N_30829);
xnor U31130 (N_31130,N_30757,N_30948);
nor U31131 (N_31131,N_30798,N_30795);
and U31132 (N_31132,N_30904,N_30914);
and U31133 (N_31133,N_30804,N_30866);
and U31134 (N_31134,N_30904,N_30753);
xor U31135 (N_31135,N_30935,N_30853);
nand U31136 (N_31136,N_30764,N_30936);
nand U31137 (N_31137,N_30878,N_30830);
and U31138 (N_31138,N_30885,N_30752);
or U31139 (N_31139,N_30936,N_30905);
and U31140 (N_31140,N_30822,N_30794);
nor U31141 (N_31141,N_30848,N_30785);
xor U31142 (N_31142,N_30838,N_30893);
xor U31143 (N_31143,N_30953,N_30853);
xnor U31144 (N_31144,N_30926,N_30755);
and U31145 (N_31145,N_30806,N_30804);
and U31146 (N_31146,N_30891,N_30914);
xor U31147 (N_31147,N_30902,N_30806);
nand U31148 (N_31148,N_30957,N_30792);
and U31149 (N_31149,N_30803,N_30758);
nand U31150 (N_31150,N_30832,N_30854);
nand U31151 (N_31151,N_30880,N_30869);
xnor U31152 (N_31152,N_30903,N_30891);
or U31153 (N_31153,N_30887,N_30913);
nand U31154 (N_31154,N_30866,N_30870);
or U31155 (N_31155,N_30843,N_30872);
nor U31156 (N_31156,N_30873,N_30996);
nand U31157 (N_31157,N_30860,N_30922);
and U31158 (N_31158,N_30875,N_30944);
or U31159 (N_31159,N_30891,N_30947);
nand U31160 (N_31160,N_30869,N_30841);
or U31161 (N_31161,N_30869,N_30975);
xnor U31162 (N_31162,N_30781,N_30979);
and U31163 (N_31163,N_30840,N_30767);
nor U31164 (N_31164,N_30854,N_30915);
nor U31165 (N_31165,N_30840,N_30771);
nand U31166 (N_31166,N_30923,N_30928);
nand U31167 (N_31167,N_30871,N_30828);
xnor U31168 (N_31168,N_30931,N_30985);
and U31169 (N_31169,N_30871,N_30865);
and U31170 (N_31170,N_30925,N_30891);
nand U31171 (N_31171,N_30988,N_30886);
or U31172 (N_31172,N_30951,N_30941);
nand U31173 (N_31173,N_30757,N_30997);
nand U31174 (N_31174,N_30774,N_30935);
nor U31175 (N_31175,N_30772,N_30989);
nor U31176 (N_31176,N_30761,N_30890);
nand U31177 (N_31177,N_30933,N_30827);
xnor U31178 (N_31178,N_30947,N_30927);
nand U31179 (N_31179,N_30871,N_30901);
and U31180 (N_31180,N_30752,N_30806);
or U31181 (N_31181,N_30905,N_30779);
and U31182 (N_31182,N_30768,N_30874);
or U31183 (N_31183,N_30808,N_30787);
and U31184 (N_31184,N_30872,N_30958);
or U31185 (N_31185,N_30923,N_30760);
nor U31186 (N_31186,N_30800,N_30873);
nor U31187 (N_31187,N_30827,N_30876);
xnor U31188 (N_31188,N_30929,N_30878);
nor U31189 (N_31189,N_30937,N_30960);
xor U31190 (N_31190,N_30753,N_30876);
or U31191 (N_31191,N_30892,N_30778);
or U31192 (N_31192,N_30987,N_30919);
and U31193 (N_31193,N_30977,N_30909);
xnor U31194 (N_31194,N_30765,N_30804);
or U31195 (N_31195,N_30878,N_30758);
nor U31196 (N_31196,N_30952,N_30859);
xor U31197 (N_31197,N_30771,N_30831);
or U31198 (N_31198,N_30996,N_30941);
xnor U31199 (N_31199,N_30828,N_30788);
and U31200 (N_31200,N_30842,N_30843);
nand U31201 (N_31201,N_30850,N_30925);
xor U31202 (N_31202,N_30981,N_30893);
and U31203 (N_31203,N_30927,N_30807);
nand U31204 (N_31204,N_30883,N_30781);
or U31205 (N_31205,N_30842,N_30964);
xnor U31206 (N_31206,N_30846,N_30861);
or U31207 (N_31207,N_30862,N_30793);
and U31208 (N_31208,N_30951,N_30893);
nand U31209 (N_31209,N_30829,N_30858);
nand U31210 (N_31210,N_30862,N_30757);
nand U31211 (N_31211,N_30896,N_30909);
or U31212 (N_31212,N_30920,N_30915);
nor U31213 (N_31213,N_30946,N_30915);
nand U31214 (N_31214,N_30940,N_30947);
and U31215 (N_31215,N_30963,N_30825);
nand U31216 (N_31216,N_30798,N_30953);
nand U31217 (N_31217,N_30900,N_30962);
nand U31218 (N_31218,N_30767,N_30934);
nor U31219 (N_31219,N_30904,N_30906);
or U31220 (N_31220,N_30971,N_30952);
nand U31221 (N_31221,N_30807,N_30770);
and U31222 (N_31222,N_30983,N_30860);
xnor U31223 (N_31223,N_30881,N_30953);
nand U31224 (N_31224,N_30957,N_30764);
and U31225 (N_31225,N_30896,N_30979);
xnor U31226 (N_31226,N_30792,N_30906);
and U31227 (N_31227,N_30793,N_30870);
xor U31228 (N_31228,N_30949,N_30967);
and U31229 (N_31229,N_30920,N_30866);
xor U31230 (N_31230,N_30892,N_30784);
xnor U31231 (N_31231,N_30958,N_30896);
or U31232 (N_31232,N_30778,N_30843);
nand U31233 (N_31233,N_30934,N_30756);
nand U31234 (N_31234,N_30798,N_30977);
and U31235 (N_31235,N_30980,N_30789);
and U31236 (N_31236,N_30936,N_30894);
or U31237 (N_31237,N_30963,N_30950);
xnor U31238 (N_31238,N_30912,N_30766);
xor U31239 (N_31239,N_30972,N_30780);
or U31240 (N_31240,N_30950,N_30943);
or U31241 (N_31241,N_30926,N_30994);
nor U31242 (N_31242,N_30829,N_30753);
nor U31243 (N_31243,N_30826,N_30998);
and U31244 (N_31244,N_30838,N_30885);
nor U31245 (N_31245,N_30988,N_30972);
and U31246 (N_31246,N_30831,N_30852);
and U31247 (N_31247,N_30762,N_30842);
xnor U31248 (N_31248,N_30928,N_30871);
or U31249 (N_31249,N_30959,N_30897);
and U31250 (N_31250,N_31181,N_31168);
nor U31251 (N_31251,N_31224,N_31107);
and U31252 (N_31252,N_31030,N_31118);
xnor U31253 (N_31253,N_31177,N_31040);
or U31254 (N_31254,N_31072,N_31152);
xor U31255 (N_31255,N_31154,N_31005);
nor U31256 (N_31256,N_31027,N_31101);
or U31257 (N_31257,N_31230,N_31212);
xor U31258 (N_31258,N_31075,N_31169);
xnor U31259 (N_31259,N_31007,N_31063);
nand U31260 (N_31260,N_31162,N_31034);
and U31261 (N_31261,N_31217,N_31013);
xor U31262 (N_31262,N_31202,N_31210);
nor U31263 (N_31263,N_31099,N_31110);
and U31264 (N_31264,N_31023,N_31014);
or U31265 (N_31265,N_31116,N_31026);
nand U31266 (N_31266,N_31125,N_31122);
nor U31267 (N_31267,N_31047,N_31247);
xnor U31268 (N_31268,N_31103,N_31143);
and U31269 (N_31269,N_31225,N_31223);
nand U31270 (N_31270,N_31094,N_31200);
xor U31271 (N_31271,N_31061,N_31095);
nand U31272 (N_31272,N_31245,N_31066);
nor U31273 (N_31273,N_31050,N_31201);
and U31274 (N_31274,N_31175,N_31028);
nor U31275 (N_31275,N_31093,N_31097);
nand U31276 (N_31276,N_31165,N_31008);
or U31277 (N_31277,N_31146,N_31074);
nand U31278 (N_31278,N_31071,N_31220);
nand U31279 (N_31279,N_31062,N_31046);
or U31280 (N_31280,N_31068,N_31057);
nor U31281 (N_31281,N_31158,N_31060);
or U31282 (N_31282,N_31003,N_31238);
nand U31283 (N_31283,N_31001,N_31240);
and U31284 (N_31284,N_31100,N_31229);
or U31285 (N_31285,N_31166,N_31002);
and U31286 (N_31286,N_31218,N_31183);
or U31287 (N_31287,N_31082,N_31138);
or U31288 (N_31288,N_31096,N_31032);
or U31289 (N_31289,N_31226,N_31073);
nand U31290 (N_31290,N_31248,N_31233);
xor U31291 (N_31291,N_31176,N_31130);
xor U31292 (N_31292,N_31174,N_31239);
and U31293 (N_31293,N_31024,N_31006);
nor U31294 (N_31294,N_31084,N_31052);
nor U31295 (N_31295,N_31081,N_31119);
or U31296 (N_31296,N_31187,N_31236);
nand U31297 (N_31297,N_31170,N_31235);
or U31298 (N_31298,N_31196,N_31038);
nand U31299 (N_31299,N_31194,N_31077);
xnor U31300 (N_31300,N_31197,N_31133);
nor U31301 (N_31301,N_31092,N_31115);
nand U31302 (N_31302,N_31159,N_31242);
or U31303 (N_31303,N_31051,N_31222);
nand U31304 (N_31304,N_31205,N_31244);
nor U31305 (N_31305,N_31121,N_31190);
and U31306 (N_31306,N_31114,N_31188);
nor U31307 (N_31307,N_31106,N_31018);
xor U31308 (N_31308,N_31022,N_31111);
and U31309 (N_31309,N_31144,N_31137);
or U31310 (N_31310,N_31173,N_31105);
nor U31311 (N_31311,N_31227,N_31070);
nand U31312 (N_31312,N_31069,N_31016);
nand U31313 (N_31313,N_31167,N_31098);
xnor U31314 (N_31314,N_31042,N_31059);
nand U31315 (N_31315,N_31141,N_31199);
and U31316 (N_31316,N_31109,N_31091);
nand U31317 (N_31317,N_31054,N_31151);
or U31318 (N_31318,N_31135,N_31039);
or U31319 (N_31319,N_31153,N_31085);
xnor U31320 (N_31320,N_31193,N_31241);
and U31321 (N_31321,N_31228,N_31161);
nor U31322 (N_31322,N_31056,N_31045);
xnor U31323 (N_31323,N_31029,N_31088);
xor U31324 (N_31324,N_31246,N_31086);
or U31325 (N_31325,N_31108,N_31120);
nor U31326 (N_31326,N_31185,N_31083);
nand U31327 (N_31327,N_31102,N_31172);
xor U31328 (N_31328,N_31204,N_31123);
and U31329 (N_31329,N_31243,N_31010);
nor U31330 (N_31330,N_31127,N_31134);
xor U31331 (N_31331,N_31148,N_31112);
or U31332 (N_31332,N_31163,N_31012);
or U31333 (N_31333,N_31155,N_31017);
xor U31334 (N_31334,N_31147,N_31019);
or U31335 (N_31335,N_31191,N_31139);
nand U31336 (N_31336,N_31221,N_31021);
nor U31337 (N_31337,N_31080,N_31213);
nor U31338 (N_31338,N_31171,N_31126);
nor U31339 (N_31339,N_31214,N_31044);
nand U31340 (N_31340,N_31009,N_31184);
nor U31341 (N_31341,N_31113,N_31164);
or U31342 (N_31342,N_31206,N_31058);
xor U31343 (N_31343,N_31182,N_31142);
nand U31344 (N_31344,N_31160,N_31195);
nor U31345 (N_31345,N_31079,N_31208);
or U31346 (N_31346,N_31249,N_31015);
nand U31347 (N_31347,N_31037,N_31136);
xnor U31348 (N_31348,N_31067,N_31041);
xnor U31349 (N_31349,N_31216,N_31237);
and U31350 (N_31350,N_31065,N_31000);
nor U31351 (N_31351,N_31104,N_31035);
nand U31352 (N_31352,N_31055,N_31231);
nor U31353 (N_31353,N_31215,N_31145);
or U31354 (N_31354,N_31129,N_31124);
and U31355 (N_31355,N_31128,N_31198);
or U31356 (N_31356,N_31132,N_31090);
xor U31357 (N_31357,N_31157,N_31180);
nor U31358 (N_31358,N_31011,N_31036);
or U31359 (N_31359,N_31043,N_31207);
nand U31360 (N_31360,N_31156,N_31031);
or U31361 (N_31361,N_31020,N_31149);
nor U31362 (N_31362,N_31048,N_31078);
xnor U31363 (N_31363,N_31064,N_31211);
or U31364 (N_31364,N_31203,N_31049);
or U31365 (N_31365,N_31025,N_31033);
xor U31366 (N_31366,N_31209,N_31186);
nor U31367 (N_31367,N_31089,N_31192);
xnor U31368 (N_31368,N_31131,N_31178);
nand U31369 (N_31369,N_31004,N_31232);
or U31370 (N_31370,N_31179,N_31117);
nand U31371 (N_31371,N_31076,N_31087);
nor U31372 (N_31372,N_31219,N_31189);
or U31373 (N_31373,N_31150,N_31140);
nand U31374 (N_31374,N_31053,N_31234);
nor U31375 (N_31375,N_31068,N_31045);
and U31376 (N_31376,N_31092,N_31025);
or U31377 (N_31377,N_31209,N_31056);
or U31378 (N_31378,N_31079,N_31158);
xor U31379 (N_31379,N_31211,N_31046);
xnor U31380 (N_31380,N_31171,N_31238);
nor U31381 (N_31381,N_31095,N_31055);
and U31382 (N_31382,N_31002,N_31213);
xnor U31383 (N_31383,N_31031,N_31195);
nand U31384 (N_31384,N_31195,N_31230);
and U31385 (N_31385,N_31246,N_31122);
nor U31386 (N_31386,N_31246,N_31188);
and U31387 (N_31387,N_31238,N_31136);
or U31388 (N_31388,N_31218,N_31099);
nand U31389 (N_31389,N_31170,N_31248);
xnor U31390 (N_31390,N_31129,N_31194);
nor U31391 (N_31391,N_31120,N_31160);
nand U31392 (N_31392,N_31228,N_31157);
nor U31393 (N_31393,N_31168,N_31017);
nand U31394 (N_31394,N_31213,N_31249);
xnor U31395 (N_31395,N_31225,N_31185);
nor U31396 (N_31396,N_31049,N_31196);
and U31397 (N_31397,N_31164,N_31189);
nand U31398 (N_31398,N_31230,N_31185);
and U31399 (N_31399,N_31033,N_31111);
xor U31400 (N_31400,N_31110,N_31176);
or U31401 (N_31401,N_31213,N_31097);
nand U31402 (N_31402,N_31234,N_31172);
nand U31403 (N_31403,N_31091,N_31072);
or U31404 (N_31404,N_31205,N_31224);
xnor U31405 (N_31405,N_31084,N_31086);
or U31406 (N_31406,N_31234,N_31069);
xor U31407 (N_31407,N_31224,N_31156);
or U31408 (N_31408,N_31091,N_31112);
xor U31409 (N_31409,N_31111,N_31119);
or U31410 (N_31410,N_31215,N_31225);
and U31411 (N_31411,N_31167,N_31066);
xor U31412 (N_31412,N_31038,N_31052);
nand U31413 (N_31413,N_31088,N_31212);
or U31414 (N_31414,N_31147,N_31207);
or U31415 (N_31415,N_31110,N_31036);
or U31416 (N_31416,N_31130,N_31060);
and U31417 (N_31417,N_31028,N_31198);
nand U31418 (N_31418,N_31142,N_31163);
nand U31419 (N_31419,N_31048,N_31202);
xnor U31420 (N_31420,N_31082,N_31156);
and U31421 (N_31421,N_31017,N_31074);
nor U31422 (N_31422,N_31103,N_31189);
nor U31423 (N_31423,N_31104,N_31093);
xor U31424 (N_31424,N_31016,N_31125);
nand U31425 (N_31425,N_31181,N_31200);
or U31426 (N_31426,N_31201,N_31208);
nand U31427 (N_31427,N_31069,N_31066);
or U31428 (N_31428,N_31158,N_31076);
or U31429 (N_31429,N_31222,N_31165);
nand U31430 (N_31430,N_31205,N_31141);
nand U31431 (N_31431,N_31081,N_31241);
nand U31432 (N_31432,N_31049,N_31073);
and U31433 (N_31433,N_31137,N_31203);
nor U31434 (N_31434,N_31232,N_31217);
nand U31435 (N_31435,N_31223,N_31159);
nor U31436 (N_31436,N_31244,N_31066);
xnor U31437 (N_31437,N_31133,N_31222);
nor U31438 (N_31438,N_31128,N_31227);
and U31439 (N_31439,N_31011,N_31243);
xnor U31440 (N_31440,N_31194,N_31215);
nor U31441 (N_31441,N_31228,N_31099);
and U31442 (N_31442,N_31102,N_31004);
xnor U31443 (N_31443,N_31000,N_31223);
nor U31444 (N_31444,N_31142,N_31201);
or U31445 (N_31445,N_31241,N_31111);
xor U31446 (N_31446,N_31008,N_31122);
and U31447 (N_31447,N_31029,N_31145);
xor U31448 (N_31448,N_31061,N_31160);
xor U31449 (N_31449,N_31135,N_31163);
nor U31450 (N_31450,N_31146,N_31228);
nand U31451 (N_31451,N_31192,N_31203);
nand U31452 (N_31452,N_31164,N_31106);
nand U31453 (N_31453,N_31140,N_31090);
nor U31454 (N_31454,N_31196,N_31057);
and U31455 (N_31455,N_31157,N_31076);
nor U31456 (N_31456,N_31003,N_31192);
and U31457 (N_31457,N_31102,N_31041);
xnor U31458 (N_31458,N_31076,N_31208);
or U31459 (N_31459,N_31203,N_31237);
or U31460 (N_31460,N_31246,N_31062);
nor U31461 (N_31461,N_31088,N_31150);
and U31462 (N_31462,N_31045,N_31080);
nand U31463 (N_31463,N_31217,N_31052);
or U31464 (N_31464,N_31097,N_31216);
or U31465 (N_31465,N_31103,N_31190);
nor U31466 (N_31466,N_31213,N_31134);
or U31467 (N_31467,N_31224,N_31076);
and U31468 (N_31468,N_31123,N_31114);
nor U31469 (N_31469,N_31113,N_31105);
and U31470 (N_31470,N_31034,N_31138);
xor U31471 (N_31471,N_31219,N_31041);
nor U31472 (N_31472,N_31149,N_31175);
nand U31473 (N_31473,N_31009,N_31206);
nand U31474 (N_31474,N_31005,N_31173);
nand U31475 (N_31475,N_31149,N_31024);
nand U31476 (N_31476,N_31192,N_31067);
xnor U31477 (N_31477,N_31167,N_31025);
xor U31478 (N_31478,N_31238,N_31219);
and U31479 (N_31479,N_31064,N_31072);
and U31480 (N_31480,N_31095,N_31080);
xor U31481 (N_31481,N_31017,N_31145);
and U31482 (N_31482,N_31248,N_31049);
or U31483 (N_31483,N_31133,N_31115);
xor U31484 (N_31484,N_31142,N_31148);
nor U31485 (N_31485,N_31013,N_31032);
nand U31486 (N_31486,N_31042,N_31192);
xnor U31487 (N_31487,N_31124,N_31100);
and U31488 (N_31488,N_31245,N_31131);
nor U31489 (N_31489,N_31186,N_31138);
nor U31490 (N_31490,N_31008,N_31057);
nor U31491 (N_31491,N_31040,N_31057);
xnor U31492 (N_31492,N_31204,N_31010);
or U31493 (N_31493,N_31215,N_31184);
nor U31494 (N_31494,N_31188,N_31053);
or U31495 (N_31495,N_31167,N_31214);
nor U31496 (N_31496,N_31094,N_31206);
nor U31497 (N_31497,N_31143,N_31017);
xnor U31498 (N_31498,N_31248,N_31078);
nand U31499 (N_31499,N_31091,N_31235);
nand U31500 (N_31500,N_31481,N_31309);
nor U31501 (N_31501,N_31458,N_31349);
and U31502 (N_31502,N_31332,N_31381);
xor U31503 (N_31503,N_31352,N_31343);
xor U31504 (N_31504,N_31346,N_31294);
nor U31505 (N_31505,N_31493,N_31266);
and U31506 (N_31506,N_31492,N_31400);
nor U31507 (N_31507,N_31288,N_31329);
nand U31508 (N_31508,N_31433,N_31369);
and U31509 (N_31509,N_31425,N_31334);
and U31510 (N_31510,N_31406,N_31322);
xor U31511 (N_31511,N_31363,N_31468);
nor U31512 (N_31512,N_31386,N_31415);
and U31513 (N_31513,N_31469,N_31438);
xnor U31514 (N_31514,N_31398,N_31310);
nand U31515 (N_31515,N_31348,N_31441);
nand U31516 (N_31516,N_31337,N_31353);
nor U31517 (N_31517,N_31282,N_31414);
and U31518 (N_31518,N_31361,N_31295);
or U31519 (N_31519,N_31411,N_31264);
and U31520 (N_31520,N_31396,N_31485);
nor U31521 (N_31521,N_31432,N_31491);
and U31522 (N_31522,N_31311,N_31304);
and U31523 (N_31523,N_31312,N_31466);
xor U31524 (N_31524,N_31255,N_31268);
nor U31525 (N_31525,N_31498,N_31300);
nor U31526 (N_31526,N_31475,N_31316);
xnor U31527 (N_31527,N_31461,N_31404);
nand U31528 (N_31528,N_31465,N_31424);
nand U31529 (N_31529,N_31420,N_31428);
and U31530 (N_31530,N_31449,N_31275);
xnor U31531 (N_31531,N_31431,N_31342);
xnor U31532 (N_31532,N_31375,N_31462);
xnor U31533 (N_31533,N_31486,N_31401);
or U31534 (N_31534,N_31259,N_31366);
or U31535 (N_31535,N_31326,N_31345);
nor U31536 (N_31536,N_31418,N_31410);
or U31537 (N_31537,N_31379,N_31490);
nor U31538 (N_31538,N_31339,N_31362);
nor U31539 (N_31539,N_31499,N_31471);
and U31540 (N_31540,N_31280,N_31318);
xor U31541 (N_31541,N_31459,N_31327);
or U31542 (N_31542,N_31358,N_31292);
and U31543 (N_31543,N_31365,N_31442);
xor U31544 (N_31544,N_31279,N_31390);
nand U31545 (N_31545,N_31262,N_31370);
nor U31546 (N_31546,N_31479,N_31416);
nand U31547 (N_31547,N_31271,N_31447);
or U31548 (N_31548,N_31388,N_31454);
or U31549 (N_31549,N_31409,N_31403);
nor U31550 (N_31550,N_31395,N_31333);
xor U31551 (N_31551,N_31357,N_31489);
nand U31552 (N_31552,N_31437,N_31487);
and U31553 (N_31553,N_31281,N_31315);
xor U31554 (N_31554,N_31445,N_31399);
nor U31555 (N_31555,N_31383,N_31374);
xor U31556 (N_31556,N_31338,N_31480);
nor U31557 (N_31557,N_31354,N_31260);
and U31558 (N_31558,N_31474,N_31376);
xnor U31559 (N_31559,N_31278,N_31405);
or U31560 (N_31560,N_31336,N_31269);
nand U31561 (N_31561,N_31495,N_31270);
and U31562 (N_31562,N_31297,N_31367);
nand U31563 (N_31563,N_31306,N_31301);
nand U31564 (N_31564,N_31303,N_31263);
nand U31565 (N_31565,N_31328,N_31472);
xnor U31566 (N_31566,N_31276,N_31456);
nand U31567 (N_31567,N_31307,N_31277);
nand U31568 (N_31568,N_31261,N_31319);
nor U31569 (N_31569,N_31457,N_31308);
nand U31570 (N_31570,N_31360,N_31453);
nor U31571 (N_31571,N_31347,N_31325);
or U31572 (N_31572,N_31330,N_31478);
nand U31573 (N_31573,N_31384,N_31422);
and U31574 (N_31574,N_31427,N_31446);
and U31575 (N_31575,N_31382,N_31443);
xor U31576 (N_31576,N_31448,N_31440);
and U31577 (N_31577,N_31385,N_31430);
or U31578 (N_31578,N_31299,N_31484);
nand U31579 (N_31579,N_31378,N_31253);
nor U31580 (N_31580,N_31402,N_31284);
and U31581 (N_31581,N_31256,N_31265);
nand U31582 (N_31582,N_31436,N_31283);
and U31583 (N_31583,N_31341,N_31377);
nand U31584 (N_31584,N_31391,N_31408);
and U31585 (N_31585,N_31317,N_31380);
nand U31586 (N_31586,N_31389,N_31397);
xnor U31587 (N_31587,N_31393,N_31464);
or U31588 (N_31588,N_31298,N_31272);
nand U31589 (N_31589,N_31289,N_31452);
xor U31590 (N_31590,N_31323,N_31413);
nor U31591 (N_31591,N_31476,N_31372);
nor U31592 (N_31592,N_31435,N_31313);
nand U31593 (N_31593,N_31296,N_31417);
nor U31594 (N_31594,N_31387,N_31302);
or U31595 (N_31595,N_31460,N_31254);
or U31596 (N_31596,N_31496,N_31305);
and U31597 (N_31597,N_31290,N_31273);
xnor U31598 (N_31598,N_31473,N_31455);
or U31599 (N_31599,N_31373,N_31286);
nand U31600 (N_31600,N_31451,N_31250);
or U31601 (N_31601,N_31291,N_31285);
or U31602 (N_31602,N_31321,N_31324);
xor U31603 (N_31603,N_31467,N_31482);
and U31604 (N_31604,N_31252,N_31421);
nand U31605 (N_31605,N_31320,N_31267);
nand U31606 (N_31606,N_31331,N_31274);
and U31607 (N_31607,N_31251,N_31426);
nand U31608 (N_31608,N_31477,N_31258);
or U31609 (N_31609,N_31371,N_31392);
nand U31610 (N_31610,N_31351,N_31419);
nand U31611 (N_31611,N_31463,N_31257);
or U31612 (N_31612,N_31494,N_31429);
nand U31613 (N_31613,N_31350,N_31364);
nand U31614 (N_31614,N_31293,N_31340);
nor U31615 (N_31615,N_31444,N_31355);
or U31616 (N_31616,N_31359,N_31450);
or U31617 (N_31617,N_31335,N_31287);
nand U31618 (N_31618,N_31488,N_31423);
or U31619 (N_31619,N_31439,N_31407);
and U31620 (N_31620,N_31470,N_31344);
nor U31621 (N_31621,N_31434,N_31497);
or U31622 (N_31622,N_31368,N_31394);
or U31623 (N_31623,N_31314,N_31483);
nand U31624 (N_31624,N_31412,N_31356);
nor U31625 (N_31625,N_31436,N_31364);
nor U31626 (N_31626,N_31259,N_31419);
xor U31627 (N_31627,N_31287,N_31397);
nand U31628 (N_31628,N_31445,N_31426);
and U31629 (N_31629,N_31478,N_31361);
nand U31630 (N_31630,N_31312,N_31347);
and U31631 (N_31631,N_31375,N_31381);
and U31632 (N_31632,N_31428,N_31459);
and U31633 (N_31633,N_31263,N_31298);
and U31634 (N_31634,N_31251,N_31289);
or U31635 (N_31635,N_31409,N_31452);
or U31636 (N_31636,N_31397,N_31254);
nor U31637 (N_31637,N_31354,N_31261);
or U31638 (N_31638,N_31371,N_31416);
and U31639 (N_31639,N_31415,N_31261);
nand U31640 (N_31640,N_31262,N_31271);
nor U31641 (N_31641,N_31356,N_31498);
and U31642 (N_31642,N_31470,N_31369);
nor U31643 (N_31643,N_31482,N_31307);
or U31644 (N_31644,N_31316,N_31343);
xnor U31645 (N_31645,N_31270,N_31379);
nand U31646 (N_31646,N_31294,N_31293);
nor U31647 (N_31647,N_31350,N_31271);
nand U31648 (N_31648,N_31435,N_31389);
and U31649 (N_31649,N_31440,N_31306);
nor U31650 (N_31650,N_31460,N_31368);
and U31651 (N_31651,N_31449,N_31297);
nor U31652 (N_31652,N_31415,N_31287);
and U31653 (N_31653,N_31348,N_31272);
xor U31654 (N_31654,N_31498,N_31309);
nor U31655 (N_31655,N_31292,N_31458);
or U31656 (N_31656,N_31374,N_31484);
xor U31657 (N_31657,N_31308,N_31335);
xor U31658 (N_31658,N_31439,N_31284);
nand U31659 (N_31659,N_31381,N_31431);
nand U31660 (N_31660,N_31401,N_31351);
or U31661 (N_31661,N_31254,N_31405);
and U31662 (N_31662,N_31380,N_31351);
or U31663 (N_31663,N_31320,N_31354);
or U31664 (N_31664,N_31332,N_31271);
or U31665 (N_31665,N_31271,N_31252);
or U31666 (N_31666,N_31306,N_31379);
or U31667 (N_31667,N_31363,N_31276);
xor U31668 (N_31668,N_31317,N_31374);
and U31669 (N_31669,N_31490,N_31403);
or U31670 (N_31670,N_31353,N_31305);
or U31671 (N_31671,N_31257,N_31254);
or U31672 (N_31672,N_31359,N_31330);
nor U31673 (N_31673,N_31436,N_31298);
and U31674 (N_31674,N_31361,N_31310);
or U31675 (N_31675,N_31257,N_31372);
and U31676 (N_31676,N_31327,N_31265);
xnor U31677 (N_31677,N_31344,N_31422);
and U31678 (N_31678,N_31386,N_31446);
nand U31679 (N_31679,N_31453,N_31442);
and U31680 (N_31680,N_31477,N_31435);
nor U31681 (N_31681,N_31384,N_31372);
xor U31682 (N_31682,N_31359,N_31441);
nand U31683 (N_31683,N_31261,N_31332);
or U31684 (N_31684,N_31477,N_31283);
and U31685 (N_31685,N_31391,N_31442);
xor U31686 (N_31686,N_31443,N_31463);
or U31687 (N_31687,N_31343,N_31305);
xnor U31688 (N_31688,N_31468,N_31319);
and U31689 (N_31689,N_31399,N_31306);
nor U31690 (N_31690,N_31250,N_31368);
or U31691 (N_31691,N_31454,N_31314);
xnor U31692 (N_31692,N_31343,N_31450);
xor U31693 (N_31693,N_31278,N_31431);
nand U31694 (N_31694,N_31400,N_31306);
nor U31695 (N_31695,N_31488,N_31296);
or U31696 (N_31696,N_31475,N_31461);
nand U31697 (N_31697,N_31297,N_31409);
and U31698 (N_31698,N_31413,N_31326);
and U31699 (N_31699,N_31365,N_31450);
and U31700 (N_31700,N_31385,N_31254);
nand U31701 (N_31701,N_31436,N_31280);
nand U31702 (N_31702,N_31409,N_31258);
xor U31703 (N_31703,N_31335,N_31278);
nor U31704 (N_31704,N_31252,N_31297);
and U31705 (N_31705,N_31480,N_31393);
nand U31706 (N_31706,N_31320,N_31290);
nand U31707 (N_31707,N_31398,N_31331);
xor U31708 (N_31708,N_31297,N_31339);
and U31709 (N_31709,N_31373,N_31274);
nand U31710 (N_31710,N_31495,N_31301);
xnor U31711 (N_31711,N_31412,N_31304);
and U31712 (N_31712,N_31288,N_31492);
nand U31713 (N_31713,N_31287,N_31474);
and U31714 (N_31714,N_31489,N_31285);
xor U31715 (N_31715,N_31302,N_31449);
nor U31716 (N_31716,N_31298,N_31447);
nand U31717 (N_31717,N_31309,N_31449);
nand U31718 (N_31718,N_31267,N_31287);
nand U31719 (N_31719,N_31311,N_31444);
or U31720 (N_31720,N_31308,N_31448);
nand U31721 (N_31721,N_31336,N_31272);
nand U31722 (N_31722,N_31351,N_31413);
xor U31723 (N_31723,N_31343,N_31300);
nand U31724 (N_31724,N_31450,N_31457);
or U31725 (N_31725,N_31453,N_31380);
xor U31726 (N_31726,N_31257,N_31262);
or U31727 (N_31727,N_31407,N_31466);
or U31728 (N_31728,N_31420,N_31333);
or U31729 (N_31729,N_31410,N_31444);
or U31730 (N_31730,N_31275,N_31267);
nor U31731 (N_31731,N_31472,N_31257);
or U31732 (N_31732,N_31258,N_31334);
nor U31733 (N_31733,N_31293,N_31353);
nor U31734 (N_31734,N_31361,N_31381);
nor U31735 (N_31735,N_31289,N_31406);
nor U31736 (N_31736,N_31309,N_31264);
nand U31737 (N_31737,N_31496,N_31339);
or U31738 (N_31738,N_31476,N_31348);
and U31739 (N_31739,N_31256,N_31446);
and U31740 (N_31740,N_31276,N_31313);
and U31741 (N_31741,N_31318,N_31443);
and U31742 (N_31742,N_31334,N_31388);
and U31743 (N_31743,N_31366,N_31465);
nor U31744 (N_31744,N_31434,N_31410);
and U31745 (N_31745,N_31258,N_31368);
or U31746 (N_31746,N_31429,N_31466);
nand U31747 (N_31747,N_31339,N_31288);
nor U31748 (N_31748,N_31277,N_31346);
nand U31749 (N_31749,N_31348,N_31321);
xor U31750 (N_31750,N_31725,N_31604);
xor U31751 (N_31751,N_31749,N_31587);
nand U31752 (N_31752,N_31686,N_31727);
or U31753 (N_31753,N_31730,N_31616);
nand U31754 (N_31754,N_31683,N_31501);
xor U31755 (N_31755,N_31573,N_31503);
nor U31756 (N_31756,N_31666,N_31559);
or U31757 (N_31757,N_31513,N_31557);
or U31758 (N_31758,N_31648,N_31505);
and U31759 (N_31759,N_31564,N_31664);
or U31760 (N_31760,N_31590,N_31650);
xor U31761 (N_31761,N_31563,N_31541);
or U31762 (N_31762,N_31553,N_31504);
nand U31763 (N_31763,N_31609,N_31698);
and U31764 (N_31764,N_31517,N_31585);
nand U31765 (N_31765,N_31610,N_31595);
or U31766 (N_31766,N_31511,N_31636);
nor U31767 (N_31767,N_31569,N_31623);
and U31768 (N_31768,N_31535,N_31586);
and U31769 (N_31769,N_31619,N_31746);
and U31770 (N_31770,N_31735,N_31672);
nand U31771 (N_31771,N_31649,N_31695);
xnor U31772 (N_31772,N_31721,N_31708);
and U31773 (N_31773,N_31567,N_31733);
and U31774 (N_31774,N_31568,N_31703);
xnor U31775 (N_31775,N_31651,N_31713);
or U31776 (N_31776,N_31618,N_31509);
or U31777 (N_31777,N_31642,N_31628);
nand U31778 (N_31778,N_31645,N_31533);
xor U31779 (N_31779,N_31722,N_31675);
nor U31780 (N_31780,N_31633,N_31680);
and U31781 (N_31781,N_31682,N_31589);
nand U31782 (N_31782,N_31524,N_31684);
or U31783 (N_31783,N_31669,N_31523);
nand U31784 (N_31784,N_31693,N_31577);
xor U31785 (N_31785,N_31705,N_31699);
and U31786 (N_31786,N_31744,N_31643);
nor U31787 (N_31787,N_31615,N_31570);
and U31788 (N_31788,N_31508,N_31606);
xor U31789 (N_31789,N_31690,N_31736);
or U31790 (N_31790,N_31528,N_31743);
nand U31791 (N_31791,N_31560,N_31627);
or U31792 (N_31792,N_31572,N_31670);
nor U31793 (N_31793,N_31625,N_31621);
xor U31794 (N_31794,N_31525,N_31565);
nand U31795 (N_31795,N_31566,N_31694);
and U31796 (N_31796,N_31696,N_31550);
or U31797 (N_31797,N_31520,N_31653);
and U31798 (N_31798,N_31608,N_31706);
or U31799 (N_31799,N_31717,N_31554);
nand U31800 (N_31800,N_31542,N_31647);
nor U31801 (N_31801,N_31540,N_31510);
xnor U31802 (N_31802,N_31659,N_31506);
xnor U31803 (N_31803,N_31552,N_31638);
nand U31804 (N_31804,N_31515,N_31747);
or U31805 (N_31805,N_31549,N_31734);
nand U31806 (N_31806,N_31597,N_31613);
and U31807 (N_31807,N_31514,N_31555);
nand U31808 (N_31808,N_31521,N_31728);
and U31809 (N_31809,N_31584,N_31729);
or U31810 (N_31810,N_31679,N_31726);
nand U31811 (N_31811,N_31671,N_31507);
and U31812 (N_31812,N_31576,N_31526);
or U31813 (N_31813,N_31716,N_31529);
xor U31814 (N_31814,N_31532,N_31723);
nand U31815 (N_31815,N_31662,N_31689);
or U31816 (N_31816,N_31538,N_31715);
or U31817 (N_31817,N_31592,N_31678);
xnor U31818 (N_31818,N_31711,N_31668);
and U31819 (N_31819,N_31620,N_31632);
and U31820 (N_31820,N_31740,N_31537);
xor U31821 (N_31821,N_31534,N_31677);
xnor U31822 (N_31822,N_31531,N_31667);
nand U31823 (N_31823,N_31704,N_31545);
xnor U31824 (N_31824,N_31731,N_31718);
and U31825 (N_31825,N_31579,N_31634);
xnor U31826 (N_31826,N_31539,N_31547);
nor U31827 (N_31827,N_31596,N_31732);
or U31828 (N_31828,N_31544,N_31548);
xnor U31829 (N_31829,N_31631,N_31603);
xor U31830 (N_31830,N_31700,N_31739);
xnor U31831 (N_31831,N_31712,N_31676);
and U31832 (N_31832,N_31530,N_31661);
nor U31833 (N_31833,N_31518,N_31702);
nor U31834 (N_31834,N_31607,N_31574);
xor U31835 (N_31835,N_31720,N_31561);
nand U31836 (N_31836,N_31630,N_31629);
nor U31837 (N_31837,N_31652,N_31685);
and U31838 (N_31838,N_31654,N_31737);
and U31839 (N_31839,N_31724,N_31626);
and U31840 (N_31840,N_31502,N_31637);
xor U31841 (N_31841,N_31692,N_31512);
xnor U31842 (N_31842,N_31543,N_31598);
nand U31843 (N_31843,N_31742,N_31583);
and U31844 (N_31844,N_31738,N_31655);
or U31845 (N_31845,N_31660,N_31635);
nand U31846 (N_31846,N_31710,N_31681);
and U31847 (N_31847,N_31593,N_31556);
nand U31848 (N_31848,N_31578,N_31500);
or U31849 (N_31849,N_31562,N_31599);
xor U31850 (N_31850,N_31674,N_31546);
or U31851 (N_31851,N_31656,N_31605);
nand U31852 (N_31852,N_31582,N_31575);
and U31853 (N_31853,N_31558,N_31571);
and U31854 (N_31854,N_31617,N_31591);
nand U31855 (N_31855,N_31657,N_31611);
nand U31856 (N_31856,N_31536,N_31741);
or U31857 (N_31857,N_31663,N_31519);
xor U31858 (N_31858,N_31640,N_31687);
xor U31859 (N_31859,N_31646,N_31691);
nand U31860 (N_31860,N_31665,N_31709);
and U31861 (N_31861,N_31719,N_31624);
xnor U31862 (N_31862,N_31644,N_31658);
and U31863 (N_31863,N_31639,N_31748);
and U31864 (N_31864,N_31522,N_31612);
or U31865 (N_31865,N_31622,N_31580);
or U31866 (N_31866,N_31641,N_31601);
nor U31867 (N_31867,N_31714,N_31594);
nand U31868 (N_31868,N_31551,N_31745);
nor U31869 (N_31869,N_31673,N_31581);
xor U31870 (N_31870,N_31701,N_31707);
xor U31871 (N_31871,N_31697,N_31527);
nor U31872 (N_31872,N_31588,N_31688);
nand U31873 (N_31873,N_31602,N_31516);
nor U31874 (N_31874,N_31600,N_31614);
nand U31875 (N_31875,N_31650,N_31721);
nand U31876 (N_31876,N_31620,N_31659);
xnor U31877 (N_31877,N_31501,N_31583);
or U31878 (N_31878,N_31745,N_31669);
and U31879 (N_31879,N_31510,N_31722);
and U31880 (N_31880,N_31526,N_31609);
or U31881 (N_31881,N_31743,N_31717);
xnor U31882 (N_31882,N_31581,N_31742);
xnor U31883 (N_31883,N_31613,N_31594);
and U31884 (N_31884,N_31554,N_31570);
nand U31885 (N_31885,N_31532,N_31742);
xor U31886 (N_31886,N_31615,N_31639);
nor U31887 (N_31887,N_31657,N_31534);
nand U31888 (N_31888,N_31636,N_31712);
or U31889 (N_31889,N_31632,N_31561);
xnor U31890 (N_31890,N_31596,N_31652);
nand U31891 (N_31891,N_31668,N_31718);
nor U31892 (N_31892,N_31551,N_31585);
or U31893 (N_31893,N_31519,N_31660);
nor U31894 (N_31894,N_31696,N_31577);
and U31895 (N_31895,N_31714,N_31685);
xor U31896 (N_31896,N_31526,N_31701);
nand U31897 (N_31897,N_31560,N_31575);
and U31898 (N_31898,N_31512,N_31510);
xnor U31899 (N_31899,N_31673,N_31701);
nor U31900 (N_31900,N_31506,N_31700);
and U31901 (N_31901,N_31661,N_31553);
nor U31902 (N_31902,N_31749,N_31586);
xnor U31903 (N_31903,N_31574,N_31625);
or U31904 (N_31904,N_31631,N_31684);
or U31905 (N_31905,N_31667,N_31612);
nand U31906 (N_31906,N_31657,N_31725);
nand U31907 (N_31907,N_31533,N_31514);
nand U31908 (N_31908,N_31693,N_31618);
xor U31909 (N_31909,N_31677,N_31745);
nor U31910 (N_31910,N_31505,N_31645);
nand U31911 (N_31911,N_31665,N_31580);
nand U31912 (N_31912,N_31604,N_31593);
and U31913 (N_31913,N_31618,N_31746);
or U31914 (N_31914,N_31548,N_31699);
or U31915 (N_31915,N_31573,N_31700);
and U31916 (N_31916,N_31585,N_31695);
xor U31917 (N_31917,N_31677,N_31575);
nand U31918 (N_31918,N_31550,N_31578);
or U31919 (N_31919,N_31698,N_31716);
xor U31920 (N_31920,N_31543,N_31576);
nand U31921 (N_31921,N_31660,N_31616);
and U31922 (N_31922,N_31561,N_31709);
nand U31923 (N_31923,N_31580,N_31723);
nand U31924 (N_31924,N_31519,N_31506);
xnor U31925 (N_31925,N_31628,N_31586);
nor U31926 (N_31926,N_31512,N_31593);
and U31927 (N_31927,N_31660,N_31553);
or U31928 (N_31928,N_31606,N_31533);
nor U31929 (N_31929,N_31671,N_31564);
xor U31930 (N_31930,N_31549,N_31641);
nor U31931 (N_31931,N_31698,N_31704);
nand U31932 (N_31932,N_31731,N_31538);
xnor U31933 (N_31933,N_31611,N_31641);
nor U31934 (N_31934,N_31513,N_31729);
and U31935 (N_31935,N_31590,N_31512);
nor U31936 (N_31936,N_31666,N_31603);
xor U31937 (N_31937,N_31578,N_31693);
or U31938 (N_31938,N_31523,N_31615);
nand U31939 (N_31939,N_31745,N_31577);
and U31940 (N_31940,N_31694,N_31510);
or U31941 (N_31941,N_31577,N_31623);
xnor U31942 (N_31942,N_31643,N_31622);
xnor U31943 (N_31943,N_31694,N_31627);
nor U31944 (N_31944,N_31651,N_31686);
nor U31945 (N_31945,N_31620,N_31713);
nand U31946 (N_31946,N_31680,N_31641);
nand U31947 (N_31947,N_31671,N_31733);
xnor U31948 (N_31948,N_31522,N_31689);
nor U31949 (N_31949,N_31508,N_31733);
nand U31950 (N_31950,N_31690,N_31517);
nand U31951 (N_31951,N_31586,N_31593);
and U31952 (N_31952,N_31539,N_31638);
xor U31953 (N_31953,N_31649,N_31590);
and U31954 (N_31954,N_31544,N_31516);
xor U31955 (N_31955,N_31710,N_31554);
xnor U31956 (N_31956,N_31586,N_31746);
and U31957 (N_31957,N_31671,N_31504);
nand U31958 (N_31958,N_31637,N_31716);
and U31959 (N_31959,N_31657,N_31510);
or U31960 (N_31960,N_31646,N_31543);
or U31961 (N_31961,N_31608,N_31599);
and U31962 (N_31962,N_31706,N_31749);
xor U31963 (N_31963,N_31605,N_31623);
xor U31964 (N_31964,N_31571,N_31529);
and U31965 (N_31965,N_31683,N_31575);
or U31966 (N_31966,N_31529,N_31736);
xor U31967 (N_31967,N_31679,N_31633);
xnor U31968 (N_31968,N_31728,N_31668);
and U31969 (N_31969,N_31610,N_31543);
nor U31970 (N_31970,N_31699,N_31611);
xor U31971 (N_31971,N_31597,N_31632);
or U31972 (N_31972,N_31542,N_31607);
nand U31973 (N_31973,N_31524,N_31626);
nor U31974 (N_31974,N_31510,N_31597);
or U31975 (N_31975,N_31531,N_31609);
and U31976 (N_31976,N_31709,N_31547);
or U31977 (N_31977,N_31745,N_31612);
or U31978 (N_31978,N_31509,N_31674);
or U31979 (N_31979,N_31657,N_31664);
or U31980 (N_31980,N_31606,N_31510);
nor U31981 (N_31981,N_31522,N_31567);
nand U31982 (N_31982,N_31593,N_31675);
nor U31983 (N_31983,N_31562,N_31629);
xor U31984 (N_31984,N_31578,N_31566);
and U31985 (N_31985,N_31679,N_31656);
xnor U31986 (N_31986,N_31748,N_31697);
and U31987 (N_31987,N_31567,N_31523);
or U31988 (N_31988,N_31688,N_31724);
xor U31989 (N_31989,N_31666,N_31695);
nor U31990 (N_31990,N_31615,N_31691);
nand U31991 (N_31991,N_31570,N_31714);
nor U31992 (N_31992,N_31510,N_31617);
nand U31993 (N_31993,N_31567,N_31730);
and U31994 (N_31994,N_31602,N_31702);
or U31995 (N_31995,N_31509,N_31619);
or U31996 (N_31996,N_31577,N_31649);
or U31997 (N_31997,N_31735,N_31557);
xor U31998 (N_31998,N_31612,N_31641);
nor U31999 (N_31999,N_31550,N_31584);
nand U32000 (N_32000,N_31805,N_31916);
and U32001 (N_32001,N_31991,N_31984);
or U32002 (N_32002,N_31933,N_31924);
or U32003 (N_32003,N_31918,N_31820);
nand U32004 (N_32004,N_31883,N_31829);
or U32005 (N_32005,N_31894,N_31761);
and U32006 (N_32006,N_31774,N_31983);
nor U32007 (N_32007,N_31967,N_31995);
and U32008 (N_32008,N_31977,N_31852);
and U32009 (N_32009,N_31886,N_31903);
xnor U32010 (N_32010,N_31838,N_31930);
xnor U32011 (N_32011,N_31937,N_31942);
nor U32012 (N_32012,N_31986,N_31970);
nor U32013 (N_32013,N_31853,N_31925);
nand U32014 (N_32014,N_31907,N_31823);
xor U32015 (N_32015,N_31885,N_31893);
and U32016 (N_32016,N_31815,N_31781);
and U32017 (N_32017,N_31811,N_31947);
nor U32018 (N_32018,N_31783,N_31888);
xnor U32019 (N_32019,N_31817,N_31834);
nand U32020 (N_32020,N_31826,N_31806);
nand U32021 (N_32021,N_31803,N_31813);
and U32022 (N_32022,N_31818,N_31985);
nand U32023 (N_32023,N_31982,N_31875);
or U32024 (N_32024,N_31862,N_31775);
nand U32025 (N_32025,N_31992,N_31821);
nor U32026 (N_32026,N_31996,N_31868);
xnor U32027 (N_32027,N_31994,N_31767);
or U32028 (N_32028,N_31856,N_31915);
xor U32029 (N_32029,N_31962,N_31766);
nand U32030 (N_32030,N_31851,N_31921);
or U32031 (N_32031,N_31861,N_31895);
or U32032 (N_32032,N_31989,N_31972);
and U32033 (N_32033,N_31874,N_31891);
nor U32034 (N_32034,N_31754,N_31906);
or U32035 (N_32035,N_31797,N_31863);
xor U32036 (N_32036,N_31917,N_31884);
xor U32037 (N_32037,N_31940,N_31946);
xor U32038 (N_32038,N_31948,N_31959);
or U32039 (N_32039,N_31901,N_31978);
nor U32040 (N_32040,N_31997,N_31810);
and U32041 (N_32041,N_31931,N_31908);
xor U32042 (N_32042,N_31787,N_31859);
and U32043 (N_32043,N_31943,N_31912);
nand U32044 (N_32044,N_31825,N_31858);
and U32045 (N_32045,N_31763,N_31794);
xnor U32046 (N_32046,N_31831,N_31929);
nand U32047 (N_32047,N_31869,N_31864);
xnor U32048 (N_32048,N_31846,N_31876);
nor U32049 (N_32049,N_31923,N_31824);
nand U32050 (N_32050,N_31758,N_31988);
or U32051 (N_32051,N_31779,N_31934);
nand U32052 (N_32052,N_31958,N_31936);
nor U32053 (N_32053,N_31975,N_31833);
nand U32054 (N_32054,N_31878,N_31960);
nand U32055 (N_32055,N_31932,N_31927);
nand U32056 (N_32056,N_31848,N_31777);
nand U32057 (N_32057,N_31966,N_31772);
and U32058 (N_32058,N_31780,N_31782);
or U32059 (N_32059,N_31757,N_31939);
and U32060 (N_32060,N_31765,N_31922);
xnor U32061 (N_32061,N_31755,N_31814);
nand U32062 (N_32062,N_31796,N_31870);
or U32063 (N_32063,N_31800,N_31841);
or U32064 (N_32064,N_31752,N_31961);
nand U32065 (N_32065,N_31809,N_31771);
and U32066 (N_32066,N_31873,N_31865);
or U32067 (N_32067,N_31785,N_31872);
or U32068 (N_32068,N_31920,N_31956);
xnor U32069 (N_32069,N_31999,N_31788);
or U32070 (N_32070,N_31849,N_31963);
or U32071 (N_32071,N_31981,N_31879);
or U32072 (N_32072,N_31974,N_31953);
and U32073 (N_32073,N_31786,N_31949);
nand U32074 (N_32074,N_31843,N_31902);
nor U32075 (N_32075,N_31990,N_31760);
or U32076 (N_32076,N_31898,N_31778);
or U32077 (N_32077,N_31768,N_31845);
and U32078 (N_32078,N_31890,N_31950);
or U32079 (N_32079,N_31877,N_31836);
or U32080 (N_32080,N_31957,N_31993);
nor U32081 (N_32081,N_31971,N_31881);
nand U32082 (N_32082,N_31954,N_31802);
nand U32083 (N_32083,N_31987,N_31832);
and U32084 (N_32084,N_31784,N_31790);
and U32085 (N_32085,N_31792,N_31855);
or U32086 (N_32086,N_31847,N_31854);
and U32087 (N_32087,N_31909,N_31835);
nand U32088 (N_32088,N_31762,N_31905);
and U32089 (N_32089,N_31795,N_31756);
or U32090 (N_32090,N_31839,N_31899);
nand U32091 (N_32091,N_31827,N_31976);
xor U32092 (N_32092,N_31871,N_31764);
xor U32093 (N_32093,N_31773,N_31919);
nor U32094 (N_32094,N_31945,N_31789);
nor U32095 (N_32095,N_31892,N_31882);
or U32096 (N_32096,N_31889,N_31842);
and U32097 (N_32097,N_31804,N_31840);
nand U32098 (N_32098,N_31822,N_31860);
nand U32099 (N_32099,N_31944,N_31955);
nand U32100 (N_32100,N_31769,N_31793);
xnor U32101 (N_32101,N_31968,N_31911);
or U32102 (N_32102,N_31951,N_31844);
nand U32103 (N_32103,N_31857,N_31807);
and U32104 (N_32104,N_31866,N_31799);
xnor U32105 (N_32105,N_31751,N_31897);
nor U32106 (N_32106,N_31850,N_31750);
xnor U32107 (N_32107,N_31798,N_31776);
nor U32108 (N_32108,N_31914,N_31808);
xor U32109 (N_32109,N_31770,N_31941);
nand U32110 (N_32110,N_31973,N_31969);
xor U32111 (N_32111,N_31791,N_31965);
nor U32112 (N_32112,N_31900,N_31828);
nor U32113 (N_32113,N_31980,N_31935);
and U32114 (N_32114,N_31928,N_31952);
nor U32115 (N_32115,N_31926,N_31896);
or U32116 (N_32116,N_31812,N_31998);
and U32117 (N_32117,N_31801,N_31867);
nor U32118 (N_32118,N_31837,N_31938);
nand U32119 (N_32119,N_31964,N_31816);
nor U32120 (N_32120,N_31830,N_31753);
or U32121 (N_32121,N_31910,N_31913);
or U32122 (N_32122,N_31887,N_31979);
or U32123 (N_32123,N_31819,N_31759);
or U32124 (N_32124,N_31904,N_31880);
xor U32125 (N_32125,N_31950,N_31854);
nand U32126 (N_32126,N_31777,N_31896);
or U32127 (N_32127,N_31959,N_31848);
xor U32128 (N_32128,N_31803,N_31794);
and U32129 (N_32129,N_31750,N_31810);
xor U32130 (N_32130,N_31827,N_31865);
or U32131 (N_32131,N_31998,N_31954);
nor U32132 (N_32132,N_31932,N_31815);
or U32133 (N_32133,N_31872,N_31943);
and U32134 (N_32134,N_31895,N_31867);
xor U32135 (N_32135,N_31846,N_31834);
nor U32136 (N_32136,N_31944,N_31761);
nor U32137 (N_32137,N_31962,N_31857);
xnor U32138 (N_32138,N_31910,N_31757);
xnor U32139 (N_32139,N_31873,N_31855);
nor U32140 (N_32140,N_31809,N_31995);
nand U32141 (N_32141,N_31794,N_31754);
nand U32142 (N_32142,N_31786,N_31798);
nor U32143 (N_32143,N_31810,N_31864);
nand U32144 (N_32144,N_31962,N_31966);
xnor U32145 (N_32145,N_31903,N_31781);
nand U32146 (N_32146,N_31985,N_31973);
xnor U32147 (N_32147,N_31773,N_31969);
or U32148 (N_32148,N_31975,N_31949);
and U32149 (N_32149,N_31973,N_31913);
and U32150 (N_32150,N_31947,N_31789);
and U32151 (N_32151,N_31760,N_31827);
or U32152 (N_32152,N_31830,N_31944);
nand U32153 (N_32153,N_31952,N_31844);
and U32154 (N_32154,N_31835,N_31978);
nand U32155 (N_32155,N_31823,N_31814);
and U32156 (N_32156,N_31966,N_31892);
or U32157 (N_32157,N_31786,N_31847);
xor U32158 (N_32158,N_31837,N_31762);
nor U32159 (N_32159,N_31812,N_31993);
and U32160 (N_32160,N_31995,N_31971);
xnor U32161 (N_32161,N_31820,N_31764);
or U32162 (N_32162,N_31962,N_31830);
nand U32163 (N_32163,N_31845,N_31916);
nand U32164 (N_32164,N_31993,N_31982);
nand U32165 (N_32165,N_31884,N_31939);
or U32166 (N_32166,N_31779,N_31849);
nor U32167 (N_32167,N_31941,N_31777);
nand U32168 (N_32168,N_31939,N_31797);
nand U32169 (N_32169,N_31909,N_31974);
nor U32170 (N_32170,N_31928,N_31876);
or U32171 (N_32171,N_31788,N_31961);
nor U32172 (N_32172,N_31989,N_31852);
xnor U32173 (N_32173,N_31971,N_31955);
or U32174 (N_32174,N_31861,N_31924);
xor U32175 (N_32175,N_31750,N_31769);
xor U32176 (N_32176,N_31809,N_31979);
nand U32177 (N_32177,N_31902,N_31802);
nor U32178 (N_32178,N_31846,N_31899);
xor U32179 (N_32179,N_31776,N_31981);
or U32180 (N_32180,N_31751,N_31870);
nand U32181 (N_32181,N_31933,N_31867);
nor U32182 (N_32182,N_31960,N_31795);
xor U32183 (N_32183,N_31921,N_31784);
xor U32184 (N_32184,N_31850,N_31958);
or U32185 (N_32185,N_31916,N_31818);
and U32186 (N_32186,N_31839,N_31833);
xor U32187 (N_32187,N_31991,N_31875);
nor U32188 (N_32188,N_31788,N_31802);
nand U32189 (N_32189,N_31764,N_31817);
and U32190 (N_32190,N_31999,N_31916);
nor U32191 (N_32191,N_31964,N_31835);
nor U32192 (N_32192,N_31810,N_31803);
xnor U32193 (N_32193,N_31891,N_31942);
or U32194 (N_32194,N_31837,N_31831);
and U32195 (N_32195,N_31752,N_31804);
nand U32196 (N_32196,N_31973,N_31752);
and U32197 (N_32197,N_31820,N_31962);
and U32198 (N_32198,N_31877,N_31799);
or U32199 (N_32199,N_31890,N_31990);
and U32200 (N_32200,N_31805,N_31863);
or U32201 (N_32201,N_31989,N_31824);
xor U32202 (N_32202,N_31867,N_31922);
or U32203 (N_32203,N_31859,N_31896);
nand U32204 (N_32204,N_31941,N_31781);
or U32205 (N_32205,N_31846,N_31875);
nand U32206 (N_32206,N_31913,N_31767);
nor U32207 (N_32207,N_31834,N_31919);
nand U32208 (N_32208,N_31782,N_31984);
nor U32209 (N_32209,N_31974,N_31906);
and U32210 (N_32210,N_31813,N_31783);
xnor U32211 (N_32211,N_31940,N_31933);
and U32212 (N_32212,N_31985,N_31810);
nand U32213 (N_32213,N_31851,N_31772);
or U32214 (N_32214,N_31947,N_31871);
or U32215 (N_32215,N_31860,N_31785);
xor U32216 (N_32216,N_31932,N_31898);
and U32217 (N_32217,N_31826,N_31864);
and U32218 (N_32218,N_31852,N_31785);
or U32219 (N_32219,N_31891,N_31844);
nand U32220 (N_32220,N_31999,N_31901);
xor U32221 (N_32221,N_31765,N_31889);
or U32222 (N_32222,N_31890,N_31852);
and U32223 (N_32223,N_31775,N_31995);
xnor U32224 (N_32224,N_31948,N_31775);
xnor U32225 (N_32225,N_31811,N_31988);
nor U32226 (N_32226,N_31964,N_31803);
xnor U32227 (N_32227,N_31786,N_31784);
nand U32228 (N_32228,N_31885,N_31970);
nand U32229 (N_32229,N_31892,N_31963);
nor U32230 (N_32230,N_31956,N_31978);
nand U32231 (N_32231,N_31980,N_31879);
xnor U32232 (N_32232,N_31822,N_31943);
nand U32233 (N_32233,N_31885,N_31866);
xor U32234 (N_32234,N_31968,N_31875);
nor U32235 (N_32235,N_31764,N_31770);
xor U32236 (N_32236,N_31781,N_31901);
and U32237 (N_32237,N_31967,N_31890);
xnor U32238 (N_32238,N_31844,N_31814);
nor U32239 (N_32239,N_31872,N_31902);
xor U32240 (N_32240,N_31877,N_31932);
nand U32241 (N_32241,N_31928,N_31752);
nand U32242 (N_32242,N_31864,N_31916);
and U32243 (N_32243,N_31954,N_31863);
nor U32244 (N_32244,N_31767,N_31894);
xor U32245 (N_32245,N_31766,N_31889);
xnor U32246 (N_32246,N_31979,N_31966);
nor U32247 (N_32247,N_31844,N_31768);
and U32248 (N_32248,N_31952,N_31764);
xnor U32249 (N_32249,N_31852,N_31751);
nand U32250 (N_32250,N_32063,N_32071);
xnor U32251 (N_32251,N_32148,N_32070);
xor U32252 (N_32252,N_32079,N_32019);
xnor U32253 (N_32253,N_32084,N_32180);
xor U32254 (N_32254,N_32026,N_32030);
and U32255 (N_32255,N_32229,N_32249);
xnor U32256 (N_32256,N_32198,N_32002);
and U32257 (N_32257,N_32149,N_32034);
nor U32258 (N_32258,N_32130,N_32075);
or U32259 (N_32259,N_32235,N_32200);
xnor U32260 (N_32260,N_32028,N_32111);
nand U32261 (N_32261,N_32205,N_32154);
xor U32262 (N_32262,N_32232,N_32006);
nor U32263 (N_32263,N_32013,N_32134);
nand U32264 (N_32264,N_32153,N_32039);
and U32265 (N_32265,N_32032,N_32053);
and U32266 (N_32266,N_32164,N_32201);
and U32267 (N_32267,N_32095,N_32114);
nor U32268 (N_32268,N_32021,N_32191);
and U32269 (N_32269,N_32179,N_32060);
xor U32270 (N_32270,N_32104,N_32231);
and U32271 (N_32271,N_32023,N_32196);
or U32272 (N_32272,N_32245,N_32100);
nor U32273 (N_32273,N_32062,N_32136);
nand U32274 (N_32274,N_32151,N_32049);
nor U32275 (N_32275,N_32225,N_32112);
nand U32276 (N_32276,N_32146,N_32190);
xor U32277 (N_32277,N_32212,N_32064);
xor U32278 (N_32278,N_32247,N_32208);
xnor U32279 (N_32279,N_32162,N_32078);
and U32280 (N_32280,N_32222,N_32025);
nor U32281 (N_32281,N_32044,N_32206);
nand U32282 (N_32282,N_32214,N_32096);
nand U32283 (N_32283,N_32169,N_32128);
xnor U32284 (N_32284,N_32077,N_32157);
nand U32285 (N_32285,N_32000,N_32193);
nor U32286 (N_32286,N_32132,N_32203);
nor U32287 (N_32287,N_32016,N_32102);
or U32288 (N_32288,N_32171,N_32218);
nand U32289 (N_32289,N_32195,N_32244);
nor U32290 (N_32290,N_32183,N_32216);
or U32291 (N_32291,N_32065,N_32088);
and U32292 (N_32292,N_32147,N_32210);
and U32293 (N_32293,N_32003,N_32174);
and U32294 (N_32294,N_32024,N_32159);
xor U32295 (N_32295,N_32061,N_32048);
nand U32296 (N_32296,N_32110,N_32005);
nand U32297 (N_32297,N_32068,N_32168);
or U32298 (N_32298,N_32054,N_32184);
nor U32299 (N_32299,N_32221,N_32083);
and U32300 (N_32300,N_32090,N_32046);
or U32301 (N_32301,N_32108,N_32226);
xnor U32302 (N_32302,N_32192,N_32129);
nor U32303 (N_32303,N_32033,N_32029);
nor U32304 (N_32304,N_32055,N_32194);
xnor U32305 (N_32305,N_32139,N_32144);
nor U32306 (N_32306,N_32118,N_32161);
xor U32307 (N_32307,N_32127,N_32175);
or U32308 (N_32308,N_32236,N_32176);
nor U32309 (N_32309,N_32215,N_32056);
nor U32310 (N_32310,N_32117,N_32242);
and U32311 (N_32311,N_32125,N_32240);
nor U32312 (N_32312,N_32042,N_32015);
nor U32313 (N_32313,N_32007,N_32124);
nor U32314 (N_32314,N_32241,N_32213);
nand U32315 (N_32315,N_32223,N_32099);
nor U32316 (N_32316,N_32069,N_32220);
nor U32317 (N_32317,N_32145,N_32237);
nand U32318 (N_32318,N_32089,N_32173);
or U32319 (N_32319,N_32121,N_32143);
and U32320 (N_32320,N_32008,N_32131);
and U32321 (N_32321,N_32073,N_32017);
nand U32322 (N_32322,N_32037,N_32076);
and U32323 (N_32323,N_32197,N_32094);
or U32324 (N_32324,N_32074,N_32209);
nand U32325 (N_32325,N_32160,N_32188);
and U32326 (N_32326,N_32067,N_32009);
or U32327 (N_32327,N_32057,N_32150);
and U32328 (N_32328,N_32081,N_32243);
nand U32329 (N_32329,N_32091,N_32022);
and U32330 (N_32330,N_32058,N_32041);
nand U32331 (N_32331,N_32217,N_32199);
and U32332 (N_32332,N_32186,N_32027);
xor U32333 (N_32333,N_32051,N_32172);
nand U32334 (N_32334,N_32142,N_32167);
and U32335 (N_32335,N_32155,N_32202);
or U32336 (N_32336,N_32211,N_32047);
xnor U32337 (N_32337,N_32101,N_32001);
or U32338 (N_32338,N_32248,N_32163);
and U32339 (N_32339,N_32072,N_32233);
or U32340 (N_32340,N_32170,N_32123);
and U32341 (N_32341,N_32105,N_32119);
nor U32342 (N_32342,N_32238,N_32230);
or U32343 (N_32343,N_32133,N_32219);
or U32344 (N_32344,N_32187,N_32038);
or U32345 (N_32345,N_32116,N_32126);
nor U32346 (N_32346,N_32020,N_32177);
or U32347 (N_32347,N_32097,N_32087);
and U32348 (N_32348,N_32107,N_32004);
nor U32349 (N_32349,N_32246,N_32012);
and U32350 (N_32350,N_32166,N_32045);
or U32351 (N_32351,N_32109,N_32137);
nand U32352 (N_32352,N_32189,N_32182);
and U32353 (N_32353,N_32010,N_32135);
and U32354 (N_32354,N_32085,N_32165);
and U32355 (N_32355,N_32122,N_32098);
or U32356 (N_32356,N_32185,N_32228);
xnor U32357 (N_32357,N_32086,N_32052);
or U32358 (N_32358,N_32093,N_32115);
and U32359 (N_32359,N_32040,N_32158);
nor U32360 (N_32360,N_32152,N_32059);
and U32361 (N_32361,N_32156,N_32043);
and U32362 (N_32362,N_32181,N_32120);
nor U32363 (N_32363,N_32011,N_32092);
nor U32364 (N_32364,N_32140,N_32080);
and U32365 (N_32365,N_32113,N_32066);
and U32366 (N_32366,N_32224,N_32106);
or U32367 (N_32367,N_32103,N_32138);
or U32368 (N_32368,N_32014,N_32239);
or U32369 (N_32369,N_32082,N_32050);
nand U32370 (N_32370,N_32018,N_32234);
or U32371 (N_32371,N_32204,N_32031);
and U32372 (N_32372,N_32141,N_32227);
nor U32373 (N_32373,N_32178,N_32036);
nand U32374 (N_32374,N_32035,N_32207);
or U32375 (N_32375,N_32192,N_32190);
or U32376 (N_32376,N_32201,N_32069);
and U32377 (N_32377,N_32061,N_32217);
xnor U32378 (N_32378,N_32163,N_32038);
nor U32379 (N_32379,N_32069,N_32113);
xnor U32380 (N_32380,N_32142,N_32184);
or U32381 (N_32381,N_32035,N_32031);
nor U32382 (N_32382,N_32106,N_32159);
nand U32383 (N_32383,N_32044,N_32107);
xnor U32384 (N_32384,N_32001,N_32092);
nor U32385 (N_32385,N_32015,N_32138);
and U32386 (N_32386,N_32028,N_32208);
nand U32387 (N_32387,N_32232,N_32166);
or U32388 (N_32388,N_32141,N_32007);
nor U32389 (N_32389,N_32170,N_32010);
nor U32390 (N_32390,N_32094,N_32114);
or U32391 (N_32391,N_32041,N_32049);
or U32392 (N_32392,N_32191,N_32249);
and U32393 (N_32393,N_32010,N_32069);
or U32394 (N_32394,N_32096,N_32161);
and U32395 (N_32395,N_32188,N_32022);
or U32396 (N_32396,N_32044,N_32045);
and U32397 (N_32397,N_32203,N_32218);
nor U32398 (N_32398,N_32027,N_32026);
xnor U32399 (N_32399,N_32074,N_32175);
and U32400 (N_32400,N_32092,N_32177);
xor U32401 (N_32401,N_32158,N_32199);
or U32402 (N_32402,N_32027,N_32246);
nor U32403 (N_32403,N_32223,N_32170);
or U32404 (N_32404,N_32175,N_32108);
xnor U32405 (N_32405,N_32012,N_32076);
xnor U32406 (N_32406,N_32014,N_32236);
xnor U32407 (N_32407,N_32219,N_32109);
or U32408 (N_32408,N_32026,N_32036);
xor U32409 (N_32409,N_32211,N_32091);
nor U32410 (N_32410,N_32138,N_32131);
or U32411 (N_32411,N_32052,N_32183);
nor U32412 (N_32412,N_32135,N_32243);
or U32413 (N_32413,N_32012,N_32036);
nand U32414 (N_32414,N_32020,N_32243);
nand U32415 (N_32415,N_32106,N_32032);
or U32416 (N_32416,N_32034,N_32245);
nand U32417 (N_32417,N_32109,N_32058);
nor U32418 (N_32418,N_32169,N_32118);
nor U32419 (N_32419,N_32201,N_32243);
nor U32420 (N_32420,N_32173,N_32175);
nand U32421 (N_32421,N_32074,N_32073);
and U32422 (N_32422,N_32221,N_32012);
xnor U32423 (N_32423,N_32241,N_32141);
and U32424 (N_32424,N_32103,N_32009);
nand U32425 (N_32425,N_32095,N_32093);
xor U32426 (N_32426,N_32235,N_32078);
nor U32427 (N_32427,N_32157,N_32079);
xor U32428 (N_32428,N_32100,N_32178);
xnor U32429 (N_32429,N_32044,N_32228);
or U32430 (N_32430,N_32141,N_32188);
nand U32431 (N_32431,N_32204,N_32016);
or U32432 (N_32432,N_32083,N_32070);
and U32433 (N_32433,N_32249,N_32217);
nand U32434 (N_32434,N_32229,N_32248);
xnor U32435 (N_32435,N_32009,N_32060);
nor U32436 (N_32436,N_32002,N_32096);
xnor U32437 (N_32437,N_32163,N_32091);
nor U32438 (N_32438,N_32155,N_32239);
xnor U32439 (N_32439,N_32244,N_32013);
xnor U32440 (N_32440,N_32189,N_32238);
xnor U32441 (N_32441,N_32000,N_32036);
and U32442 (N_32442,N_32010,N_32072);
and U32443 (N_32443,N_32168,N_32036);
xor U32444 (N_32444,N_32027,N_32033);
nand U32445 (N_32445,N_32094,N_32125);
and U32446 (N_32446,N_32193,N_32239);
and U32447 (N_32447,N_32061,N_32011);
nand U32448 (N_32448,N_32028,N_32141);
nand U32449 (N_32449,N_32216,N_32171);
and U32450 (N_32450,N_32228,N_32223);
or U32451 (N_32451,N_32226,N_32147);
and U32452 (N_32452,N_32213,N_32199);
nor U32453 (N_32453,N_32132,N_32192);
nor U32454 (N_32454,N_32095,N_32019);
and U32455 (N_32455,N_32086,N_32239);
or U32456 (N_32456,N_32073,N_32186);
nand U32457 (N_32457,N_32074,N_32094);
and U32458 (N_32458,N_32046,N_32207);
xnor U32459 (N_32459,N_32035,N_32046);
nor U32460 (N_32460,N_32229,N_32104);
xnor U32461 (N_32461,N_32206,N_32019);
or U32462 (N_32462,N_32080,N_32097);
nand U32463 (N_32463,N_32045,N_32224);
xor U32464 (N_32464,N_32058,N_32019);
nand U32465 (N_32465,N_32001,N_32188);
nand U32466 (N_32466,N_32013,N_32100);
and U32467 (N_32467,N_32221,N_32048);
nor U32468 (N_32468,N_32072,N_32186);
nor U32469 (N_32469,N_32075,N_32212);
or U32470 (N_32470,N_32064,N_32010);
and U32471 (N_32471,N_32133,N_32087);
and U32472 (N_32472,N_32152,N_32115);
nor U32473 (N_32473,N_32189,N_32043);
nand U32474 (N_32474,N_32244,N_32157);
nor U32475 (N_32475,N_32154,N_32133);
xnor U32476 (N_32476,N_32000,N_32186);
and U32477 (N_32477,N_32243,N_32078);
xnor U32478 (N_32478,N_32131,N_32006);
or U32479 (N_32479,N_32099,N_32162);
nand U32480 (N_32480,N_32228,N_32052);
and U32481 (N_32481,N_32230,N_32234);
or U32482 (N_32482,N_32076,N_32217);
and U32483 (N_32483,N_32079,N_32211);
nor U32484 (N_32484,N_32048,N_32052);
and U32485 (N_32485,N_32215,N_32182);
nand U32486 (N_32486,N_32200,N_32226);
nand U32487 (N_32487,N_32117,N_32193);
nand U32488 (N_32488,N_32129,N_32050);
and U32489 (N_32489,N_32088,N_32028);
nor U32490 (N_32490,N_32015,N_32136);
nor U32491 (N_32491,N_32207,N_32041);
xnor U32492 (N_32492,N_32207,N_32151);
xnor U32493 (N_32493,N_32024,N_32230);
nor U32494 (N_32494,N_32060,N_32164);
and U32495 (N_32495,N_32177,N_32001);
and U32496 (N_32496,N_32172,N_32214);
and U32497 (N_32497,N_32152,N_32047);
and U32498 (N_32498,N_32100,N_32195);
xnor U32499 (N_32499,N_32054,N_32140);
or U32500 (N_32500,N_32257,N_32286);
nand U32501 (N_32501,N_32341,N_32450);
xor U32502 (N_32502,N_32329,N_32491);
or U32503 (N_32503,N_32297,N_32356);
xor U32504 (N_32504,N_32413,N_32302);
or U32505 (N_32505,N_32360,N_32467);
xor U32506 (N_32506,N_32315,N_32466);
nor U32507 (N_32507,N_32392,N_32265);
nor U32508 (N_32508,N_32287,N_32310);
xor U32509 (N_32509,N_32277,N_32481);
nand U32510 (N_32510,N_32320,N_32379);
or U32511 (N_32511,N_32390,N_32458);
or U32512 (N_32512,N_32416,N_32407);
or U32513 (N_32513,N_32373,N_32300);
nor U32514 (N_32514,N_32281,N_32253);
nand U32515 (N_32515,N_32473,N_32478);
and U32516 (N_32516,N_32385,N_32486);
or U32517 (N_32517,N_32419,N_32279);
or U32518 (N_32518,N_32483,N_32410);
or U32519 (N_32519,N_32479,N_32293);
nor U32520 (N_32520,N_32388,N_32386);
or U32521 (N_32521,N_32381,N_32441);
and U32522 (N_32522,N_32397,N_32308);
xnor U32523 (N_32523,N_32280,N_32429);
or U32524 (N_32524,N_32463,N_32468);
or U32525 (N_32525,N_32430,N_32439);
xnor U32526 (N_32526,N_32278,N_32438);
nand U32527 (N_32527,N_32348,N_32260);
nand U32528 (N_32528,N_32372,N_32314);
and U32529 (N_32529,N_32275,N_32344);
or U32530 (N_32530,N_32459,N_32465);
nand U32531 (N_32531,N_32336,N_32366);
nor U32532 (N_32532,N_32284,N_32427);
nand U32533 (N_32533,N_32436,N_32487);
or U32534 (N_32534,N_32387,N_32290);
and U32535 (N_32535,N_32301,N_32259);
xor U32536 (N_32536,N_32461,N_32365);
or U32537 (N_32537,N_32440,N_32267);
nand U32538 (N_32538,N_32389,N_32402);
nor U32539 (N_32539,N_32250,N_32383);
xnor U32540 (N_32540,N_32269,N_32431);
or U32541 (N_32541,N_32362,N_32447);
nor U32542 (N_32542,N_32401,N_32499);
nand U32543 (N_32543,N_32420,N_32405);
and U32544 (N_32544,N_32444,N_32282);
xnor U32545 (N_32545,N_32437,N_32255);
and U32546 (N_32546,N_32477,N_32380);
nand U32547 (N_32547,N_32475,N_32361);
nand U32548 (N_32548,N_32271,N_32368);
and U32549 (N_32549,N_32324,N_32488);
and U32550 (N_32550,N_32307,N_32409);
xnor U32551 (N_32551,N_32332,N_32292);
xor U32552 (N_32552,N_32424,N_32495);
nor U32553 (N_32553,N_32350,N_32299);
or U32554 (N_32554,N_32484,N_32485);
and U32555 (N_32555,N_32305,N_32251);
and U32556 (N_32556,N_32496,N_32460);
and U32557 (N_32557,N_32262,N_32358);
xnor U32558 (N_32558,N_32489,N_32261);
and U32559 (N_32559,N_32454,N_32359);
xnor U32560 (N_32560,N_32342,N_32346);
or U32561 (N_32561,N_32377,N_32443);
and U32562 (N_32562,N_32474,N_32258);
and U32563 (N_32563,N_32497,N_32471);
xnor U32564 (N_32564,N_32462,N_32311);
and U32565 (N_32565,N_32325,N_32298);
nor U32566 (N_32566,N_32421,N_32445);
nor U32567 (N_32567,N_32422,N_32321);
nor U32568 (N_32568,N_32395,N_32349);
nand U32569 (N_32569,N_32352,N_32347);
or U32570 (N_32570,N_32351,N_32323);
and U32571 (N_32571,N_32370,N_32494);
nor U32572 (N_32572,N_32333,N_32452);
nor U32573 (N_32573,N_32406,N_32453);
nor U32574 (N_32574,N_32289,N_32451);
and U32575 (N_32575,N_32304,N_32476);
and U32576 (N_32576,N_32364,N_32328);
nor U32577 (N_32577,N_32403,N_32353);
nor U32578 (N_32578,N_32399,N_32480);
nand U32579 (N_32579,N_32291,N_32322);
xnor U32580 (N_32580,N_32283,N_32470);
and U32581 (N_32581,N_32382,N_32428);
xor U32582 (N_32582,N_32378,N_32433);
and U32583 (N_32583,N_32252,N_32254);
nor U32584 (N_32584,N_32331,N_32412);
nand U32585 (N_32585,N_32264,N_32270);
xor U32586 (N_32586,N_32337,N_32455);
nand U32587 (N_32587,N_32309,N_32376);
and U32588 (N_32588,N_32442,N_32273);
nand U32589 (N_32589,N_32394,N_32313);
nand U32590 (N_32590,N_32415,N_32374);
nor U32591 (N_32591,N_32369,N_32391);
xnor U32592 (N_32592,N_32256,N_32469);
xnor U32593 (N_32593,N_32426,N_32306);
xnor U32594 (N_32594,N_32285,N_32296);
or U32595 (N_32595,N_32456,N_32464);
nand U32596 (N_32596,N_32295,N_32411);
nor U32597 (N_32597,N_32448,N_32357);
xor U32598 (N_32598,N_32303,N_32363);
nor U32599 (N_32599,N_32418,N_32472);
nand U32600 (N_32600,N_32393,N_32354);
and U32601 (N_32601,N_32355,N_32498);
or U32602 (N_32602,N_32404,N_32457);
or U32603 (N_32603,N_32316,N_32340);
nand U32604 (N_32604,N_32330,N_32263);
or U32605 (N_32605,N_32425,N_32335);
nand U32606 (N_32606,N_32490,N_32414);
xor U32607 (N_32607,N_32446,N_32274);
nand U32608 (N_32608,N_32371,N_32449);
or U32609 (N_32609,N_32339,N_32268);
nor U32610 (N_32610,N_32326,N_32400);
or U32611 (N_32611,N_32435,N_32367);
and U32612 (N_32612,N_32276,N_32343);
nor U32613 (N_32613,N_32482,N_32434);
nor U32614 (N_32614,N_32334,N_32423);
and U32615 (N_32615,N_32398,N_32345);
and U32616 (N_32616,N_32492,N_32375);
or U32617 (N_32617,N_32432,N_32266);
or U32618 (N_32618,N_32317,N_32493);
xnor U32619 (N_32619,N_32327,N_32288);
nand U32620 (N_32620,N_32384,N_32338);
nor U32621 (N_32621,N_32318,N_32312);
nand U32622 (N_32622,N_32408,N_32396);
xor U32623 (N_32623,N_32294,N_32319);
or U32624 (N_32624,N_32417,N_32272);
xnor U32625 (N_32625,N_32448,N_32399);
and U32626 (N_32626,N_32491,N_32400);
nor U32627 (N_32627,N_32482,N_32311);
nand U32628 (N_32628,N_32480,N_32271);
nand U32629 (N_32629,N_32317,N_32262);
nor U32630 (N_32630,N_32289,N_32359);
xnor U32631 (N_32631,N_32325,N_32396);
nand U32632 (N_32632,N_32479,N_32374);
xnor U32633 (N_32633,N_32357,N_32356);
xnor U32634 (N_32634,N_32292,N_32378);
nor U32635 (N_32635,N_32394,N_32378);
nand U32636 (N_32636,N_32484,N_32372);
xor U32637 (N_32637,N_32391,N_32386);
nor U32638 (N_32638,N_32327,N_32276);
and U32639 (N_32639,N_32378,N_32311);
and U32640 (N_32640,N_32250,N_32387);
nand U32641 (N_32641,N_32341,N_32257);
xor U32642 (N_32642,N_32452,N_32423);
xnor U32643 (N_32643,N_32305,N_32351);
or U32644 (N_32644,N_32350,N_32494);
nor U32645 (N_32645,N_32293,N_32442);
xnor U32646 (N_32646,N_32374,N_32493);
or U32647 (N_32647,N_32477,N_32306);
and U32648 (N_32648,N_32411,N_32265);
xor U32649 (N_32649,N_32407,N_32290);
and U32650 (N_32650,N_32408,N_32494);
nand U32651 (N_32651,N_32296,N_32471);
and U32652 (N_32652,N_32305,N_32372);
or U32653 (N_32653,N_32313,N_32456);
or U32654 (N_32654,N_32278,N_32457);
nor U32655 (N_32655,N_32410,N_32281);
xor U32656 (N_32656,N_32295,N_32320);
nor U32657 (N_32657,N_32455,N_32447);
and U32658 (N_32658,N_32400,N_32455);
nor U32659 (N_32659,N_32361,N_32433);
nor U32660 (N_32660,N_32422,N_32375);
or U32661 (N_32661,N_32462,N_32450);
or U32662 (N_32662,N_32403,N_32474);
or U32663 (N_32663,N_32314,N_32287);
nand U32664 (N_32664,N_32271,N_32320);
xnor U32665 (N_32665,N_32385,N_32342);
or U32666 (N_32666,N_32482,N_32459);
nand U32667 (N_32667,N_32358,N_32390);
nand U32668 (N_32668,N_32442,N_32441);
and U32669 (N_32669,N_32476,N_32287);
nor U32670 (N_32670,N_32418,N_32405);
or U32671 (N_32671,N_32475,N_32266);
or U32672 (N_32672,N_32264,N_32398);
nand U32673 (N_32673,N_32251,N_32302);
xor U32674 (N_32674,N_32435,N_32388);
nor U32675 (N_32675,N_32342,N_32460);
xor U32676 (N_32676,N_32350,N_32309);
and U32677 (N_32677,N_32254,N_32492);
or U32678 (N_32678,N_32447,N_32351);
or U32679 (N_32679,N_32448,N_32421);
nand U32680 (N_32680,N_32462,N_32488);
and U32681 (N_32681,N_32493,N_32498);
and U32682 (N_32682,N_32342,N_32386);
or U32683 (N_32683,N_32287,N_32311);
nand U32684 (N_32684,N_32318,N_32354);
nor U32685 (N_32685,N_32319,N_32404);
nand U32686 (N_32686,N_32286,N_32326);
and U32687 (N_32687,N_32492,N_32449);
xnor U32688 (N_32688,N_32389,N_32436);
xnor U32689 (N_32689,N_32446,N_32319);
nand U32690 (N_32690,N_32372,N_32388);
and U32691 (N_32691,N_32290,N_32396);
nor U32692 (N_32692,N_32253,N_32430);
and U32693 (N_32693,N_32278,N_32450);
or U32694 (N_32694,N_32460,N_32251);
nand U32695 (N_32695,N_32450,N_32378);
or U32696 (N_32696,N_32331,N_32446);
or U32697 (N_32697,N_32410,N_32254);
xnor U32698 (N_32698,N_32355,N_32368);
nor U32699 (N_32699,N_32310,N_32353);
and U32700 (N_32700,N_32418,N_32441);
or U32701 (N_32701,N_32286,N_32276);
and U32702 (N_32702,N_32296,N_32340);
nor U32703 (N_32703,N_32397,N_32443);
xor U32704 (N_32704,N_32304,N_32418);
and U32705 (N_32705,N_32424,N_32478);
xor U32706 (N_32706,N_32401,N_32376);
and U32707 (N_32707,N_32290,N_32450);
xnor U32708 (N_32708,N_32294,N_32456);
nand U32709 (N_32709,N_32279,N_32356);
nor U32710 (N_32710,N_32313,N_32451);
or U32711 (N_32711,N_32435,N_32373);
xor U32712 (N_32712,N_32322,N_32429);
nor U32713 (N_32713,N_32251,N_32458);
and U32714 (N_32714,N_32305,N_32361);
xor U32715 (N_32715,N_32285,N_32250);
nor U32716 (N_32716,N_32344,N_32288);
nor U32717 (N_32717,N_32280,N_32309);
nand U32718 (N_32718,N_32378,N_32333);
or U32719 (N_32719,N_32344,N_32422);
xor U32720 (N_32720,N_32400,N_32446);
and U32721 (N_32721,N_32404,N_32251);
nor U32722 (N_32722,N_32356,N_32490);
or U32723 (N_32723,N_32347,N_32404);
and U32724 (N_32724,N_32251,N_32327);
xnor U32725 (N_32725,N_32443,N_32262);
nand U32726 (N_32726,N_32299,N_32374);
or U32727 (N_32727,N_32481,N_32368);
nor U32728 (N_32728,N_32278,N_32268);
or U32729 (N_32729,N_32340,N_32410);
nand U32730 (N_32730,N_32475,N_32385);
xor U32731 (N_32731,N_32285,N_32377);
xor U32732 (N_32732,N_32429,N_32289);
xor U32733 (N_32733,N_32388,N_32361);
nand U32734 (N_32734,N_32416,N_32427);
nor U32735 (N_32735,N_32483,N_32320);
xnor U32736 (N_32736,N_32273,N_32360);
xor U32737 (N_32737,N_32385,N_32270);
or U32738 (N_32738,N_32451,N_32358);
nand U32739 (N_32739,N_32429,N_32269);
and U32740 (N_32740,N_32483,N_32415);
nand U32741 (N_32741,N_32476,N_32389);
and U32742 (N_32742,N_32331,N_32478);
nor U32743 (N_32743,N_32420,N_32429);
nand U32744 (N_32744,N_32430,N_32324);
xnor U32745 (N_32745,N_32408,N_32424);
nand U32746 (N_32746,N_32436,N_32291);
nand U32747 (N_32747,N_32270,N_32267);
nand U32748 (N_32748,N_32367,N_32409);
or U32749 (N_32749,N_32452,N_32395);
or U32750 (N_32750,N_32551,N_32735);
xor U32751 (N_32751,N_32567,N_32722);
and U32752 (N_32752,N_32636,N_32583);
and U32753 (N_32753,N_32748,N_32515);
or U32754 (N_32754,N_32531,N_32621);
and U32755 (N_32755,N_32539,N_32705);
or U32756 (N_32756,N_32655,N_32598);
or U32757 (N_32757,N_32548,N_32549);
nand U32758 (N_32758,N_32668,N_32525);
xnor U32759 (N_32759,N_32633,N_32501);
or U32760 (N_32760,N_32686,N_32717);
nand U32761 (N_32761,N_32514,N_32546);
and U32762 (N_32762,N_32563,N_32641);
nor U32763 (N_32763,N_32529,N_32609);
and U32764 (N_32764,N_32683,N_32687);
or U32765 (N_32765,N_32580,N_32533);
or U32766 (N_32766,N_32632,N_32586);
nor U32767 (N_32767,N_32582,N_32726);
xor U32768 (N_32768,N_32638,N_32555);
and U32769 (N_32769,N_32723,N_32584);
xor U32770 (N_32770,N_32709,N_32509);
or U32771 (N_32771,N_32644,N_32725);
xor U32772 (N_32772,N_32696,N_32743);
nor U32773 (N_32773,N_32517,N_32716);
nor U32774 (N_32774,N_32659,N_32624);
or U32775 (N_32775,N_32541,N_32561);
nor U32776 (N_32776,N_32623,N_32628);
or U32777 (N_32777,N_32594,N_32610);
or U32778 (N_32778,N_32565,N_32654);
and U32779 (N_32779,N_32694,N_32554);
and U32780 (N_32780,N_32669,N_32570);
nor U32781 (N_32781,N_32714,N_32523);
and U32782 (N_32782,N_32685,N_32545);
xnor U32783 (N_32783,N_32608,N_32647);
and U32784 (N_32784,N_32699,N_32503);
or U32785 (N_32785,N_32592,N_32607);
nand U32786 (N_32786,N_32520,N_32662);
or U32787 (N_32787,N_32708,N_32663);
or U32788 (N_32788,N_32661,N_32508);
or U32789 (N_32789,N_32746,N_32579);
nand U32790 (N_32790,N_32619,N_32616);
nor U32791 (N_32791,N_32537,N_32587);
and U32792 (N_32792,N_32688,N_32728);
and U32793 (N_32793,N_32605,N_32600);
xnor U32794 (N_32794,N_32697,N_32693);
nand U32795 (N_32795,N_32741,N_32692);
and U32796 (N_32796,N_32742,N_32729);
or U32797 (N_32797,N_32684,N_32575);
and U32798 (N_32798,N_32682,N_32502);
xor U32799 (N_32799,N_32719,N_32552);
or U32800 (N_32800,N_32625,N_32569);
or U32801 (N_32801,N_32524,N_32639);
nor U32802 (N_32802,N_32657,N_32612);
nand U32803 (N_32803,N_32535,N_32680);
xnor U32804 (N_32804,N_32505,N_32576);
or U32805 (N_32805,N_32724,N_32574);
nand U32806 (N_32806,N_32626,N_32707);
or U32807 (N_32807,N_32677,N_32718);
and U32808 (N_32808,N_32635,N_32650);
xnor U32809 (N_32809,N_32681,N_32544);
nor U32810 (N_32810,N_32690,N_32643);
or U32811 (N_32811,N_32652,N_32599);
and U32812 (N_32812,N_32500,N_32711);
nand U32813 (N_32813,N_32634,N_32504);
and U32814 (N_32814,N_32511,N_32730);
nand U32815 (N_32815,N_32532,N_32671);
nor U32816 (N_32816,N_32595,N_32560);
or U32817 (N_32817,N_32648,N_32738);
and U32818 (N_32818,N_32704,N_32526);
and U32819 (N_32819,N_32720,N_32712);
and U32820 (N_32820,N_32557,N_32745);
xnor U32821 (N_32821,N_32553,N_32577);
nor U32822 (N_32822,N_32739,N_32572);
or U32823 (N_32823,N_32614,N_32613);
xnor U32824 (N_32824,N_32606,N_32627);
xnor U32825 (N_32825,N_32543,N_32540);
nor U32826 (N_32826,N_32665,N_32733);
or U32827 (N_32827,N_32744,N_32588);
xor U32828 (N_32828,N_32631,N_32597);
xnor U32829 (N_32829,N_32666,N_32528);
xnor U32830 (N_32830,N_32732,N_32603);
nor U32831 (N_32831,N_32700,N_32721);
nor U32832 (N_32832,N_32571,N_32566);
nand U32833 (N_32833,N_32506,N_32578);
or U32834 (N_32834,N_32637,N_32585);
xor U32835 (N_32835,N_32737,N_32695);
xor U32836 (N_32836,N_32670,N_32698);
nand U32837 (N_32837,N_32589,N_32736);
and U32838 (N_32838,N_32673,N_32701);
and U32839 (N_32839,N_32615,N_32556);
nand U32840 (N_32840,N_32510,N_32703);
nand U32841 (N_32841,N_32516,N_32596);
and U32842 (N_32842,N_32573,N_32689);
nand U32843 (N_32843,N_32660,N_32611);
nor U32844 (N_32844,N_32562,N_32581);
or U32845 (N_32845,N_32747,N_32713);
nand U32846 (N_32846,N_32678,N_32749);
nor U32847 (N_32847,N_32530,N_32564);
and U32848 (N_32848,N_32522,N_32674);
nand U32849 (N_32849,N_32653,N_32706);
xor U32850 (N_32850,N_32518,N_32675);
xnor U32851 (N_32851,N_32656,N_32536);
nand U32852 (N_32852,N_32538,N_32691);
xor U32853 (N_32853,N_32593,N_32649);
xor U32854 (N_32854,N_32629,N_32667);
nor U32855 (N_32855,N_32559,N_32601);
xor U32856 (N_32856,N_32527,N_32558);
or U32857 (N_32857,N_32715,N_32734);
nand U32858 (N_32858,N_32604,N_32513);
xnor U32859 (N_32859,N_32591,N_32550);
nand U32860 (N_32860,N_32640,N_32521);
xnor U32861 (N_32861,N_32590,N_32651);
xnor U32862 (N_32862,N_32602,N_32658);
or U32863 (N_32863,N_32664,N_32676);
nand U32864 (N_32864,N_32620,N_32512);
and U32865 (N_32865,N_32702,N_32618);
nand U32866 (N_32866,N_32740,N_32622);
or U32867 (N_32867,N_32534,N_32642);
and U32868 (N_32868,N_32727,N_32672);
or U32869 (N_32869,N_32646,N_32547);
xor U32870 (N_32870,N_32507,N_32617);
nor U32871 (N_32871,N_32519,N_32645);
nand U32872 (N_32872,N_32630,N_32568);
nand U32873 (N_32873,N_32731,N_32679);
nor U32874 (N_32874,N_32710,N_32542);
nand U32875 (N_32875,N_32721,N_32715);
or U32876 (N_32876,N_32718,N_32631);
or U32877 (N_32877,N_32698,N_32558);
and U32878 (N_32878,N_32590,N_32545);
xor U32879 (N_32879,N_32572,N_32542);
nand U32880 (N_32880,N_32689,N_32550);
and U32881 (N_32881,N_32566,N_32705);
xor U32882 (N_32882,N_32682,N_32534);
nor U32883 (N_32883,N_32610,N_32747);
nand U32884 (N_32884,N_32739,N_32540);
and U32885 (N_32885,N_32683,N_32524);
nor U32886 (N_32886,N_32604,N_32503);
nand U32887 (N_32887,N_32734,N_32563);
or U32888 (N_32888,N_32570,N_32742);
or U32889 (N_32889,N_32666,N_32745);
nor U32890 (N_32890,N_32570,N_32682);
nor U32891 (N_32891,N_32675,N_32588);
nor U32892 (N_32892,N_32523,N_32508);
and U32893 (N_32893,N_32692,N_32599);
or U32894 (N_32894,N_32636,N_32678);
xor U32895 (N_32895,N_32660,N_32515);
nor U32896 (N_32896,N_32640,N_32535);
xor U32897 (N_32897,N_32579,N_32521);
xnor U32898 (N_32898,N_32722,N_32718);
or U32899 (N_32899,N_32677,N_32641);
xor U32900 (N_32900,N_32651,N_32710);
and U32901 (N_32901,N_32574,N_32746);
or U32902 (N_32902,N_32718,N_32593);
nand U32903 (N_32903,N_32509,N_32699);
and U32904 (N_32904,N_32717,N_32705);
xor U32905 (N_32905,N_32664,N_32616);
and U32906 (N_32906,N_32628,N_32689);
xor U32907 (N_32907,N_32649,N_32646);
or U32908 (N_32908,N_32590,N_32684);
nor U32909 (N_32909,N_32663,N_32526);
or U32910 (N_32910,N_32537,N_32741);
or U32911 (N_32911,N_32534,N_32688);
and U32912 (N_32912,N_32558,N_32576);
nand U32913 (N_32913,N_32703,N_32623);
xnor U32914 (N_32914,N_32511,N_32616);
or U32915 (N_32915,N_32744,N_32645);
or U32916 (N_32916,N_32630,N_32644);
or U32917 (N_32917,N_32711,N_32617);
or U32918 (N_32918,N_32622,N_32684);
and U32919 (N_32919,N_32720,N_32703);
xor U32920 (N_32920,N_32732,N_32539);
and U32921 (N_32921,N_32561,N_32741);
and U32922 (N_32922,N_32528,N_32664);
xnor U32923 (N_32923,N_32514,N_32532);
nand U32924 (N_32924,N_32625,N_32539);
nand U32925 (N_32925,N_32535,N_32684);
or U32926 (N_32926,N_32673,N_32528);
nor U32927 (N_32927,N_32509,N_32745);
nor U32928 (N_32928,N_32676,N_32602);
xnor U32929 (N_32929,N_32552,N_32646);
nand U32930 (N_32930,N_32726,N_32746);
or U32931 (N_32931,N_32566,N_32713);
or U32932 (N_32932,N_32590,N_32567);
nor U32933 (N_32933,N_32746,N_32553);
or U32934 (N_32934,N_32546,N_32594);
or U32935 (N_32935,N_32537,N_32639);
xnor U32936 (N_32936,N_32513,N_32677);
and U32937 (N_32937,N_32624,N_32675);
or U32938 (N_32938,N_32636,N_32562);
and U32939 (N_32939,N_32715,N_32741);
and U32940 (N_32940,N_32613,N_32601);
xnor U32941 (N_32941,N_32689,N_32721);
xnor U32942 (N_32942,N_32603,N_32600);
xnor U32943 (N_32943,N_32605,N_32705);
nand U32944 (N_32944,N_32681,N_32643);
nand U32945 (N_32945,N_32724,N_32501);
or U32946 (N_32946,N_32669,N_32537);
nand U32947 (N_32947,N_32520,N_32655);
and U32948 (N_32948,N_32628,N_32742);
xnor U32949 (N_32949,N_32524,N_32711);
nor U32950 (N_32950,N_32554,N_32504);
nand U32951 (N_32951,N_32709,N_32547);
xor U32952 (N_32952,N_32649,N_32511);
xnor U32953 (N_32953,N_32535,N_32677);
nand U32954 (N_32954,N_32598,N_32621);
nand U32955 (N_32955,N_32573,N_32749);
xnor U32956 (N_32956,N_32675,N_32634);
and U32957 (N_32957,N_32671,N_32591);
or U32958 (N_32958,N_32729,N_32663);
nand U32959 (N_32959,N_32729,N_32685);
or U32960 (N_32960,N_32691,N_32600);
or U32961 (N_32961,N_32619,N_32679);
nor U32962 (N_32962,N_32563,N_32685);
nor U32963 (N_32963,N_32720,N_32534);
or U32964 (N_32964,N_32538,N_32650);
and U32965 (N_32965,N_32602,N_32633);
nor U32966 (N_32966,N_32514,N_32659);
or U32967 (N_32967,N_32610,N_32658);
xnor U32968 (N_32968,N_32610,N_32585);
xnor U32969 (N_32969,N_32627,N_32600);
and U32970 (N_32970,N_32676,N_32719);
and U32971 (N_32971,N_32743,N_32517);
nor U32972 (N_32972,N_32555,N_32526);
nor U32973 (N_32973,N_32501,N_32671);
and U32974 (N_32974,N_32579,N_32728);
and U32975 (N_32975,N_32636,N_32545);
or U32976 (N_32976,N_32732,N_32567);
nor U32977 (N_32977,N_32590,N_32621);
or U32978 (N_32978,N_32561,N_32681);
nor U32979 (N_32979,N_32571,N_32500);
and U32980 (N_32980,N_32544,N_32742);
nor U32981 (N_32981,N_32539,N_32556);
and U32982 (N_32982,N_32604,N_32512);
nand U32983 (N_32983,N_32616,N_32600);
and U32984 (N_32984,N_32603,N_32661);
nand U32985 (N_32985,N_32646,N_32559);
and U32986 (N_32986,N_32708,N_32607);
or U32987 (N_32987,N_32690,N_32639);
xnor U32988 (N_32988,N_32711,N_32561);
nor U32989 (N_32989,N_32733,N_32590);
and U32990 (N_32990,N_32577,N_32611);
nand U32991 (N_32991,N_32630,N_32745);
nand U32992 (N_32992,N_32685,N_32597);
or U32993 (N_32993,N_32523,N_32677);
nand U32994 (N_32994,N_32636,N_32605);
and U32995 (N_32995,N_32510,N_32597);
or U32996 (N_32996,N_32563,N_32639);
nand U32997 (N_32997,N_32725,N_32743);
and U32998 (N_32998,N_32694,N_32599);
and U32999 (N_32999,N_32697,N_32554);
xor U33000 (N_33000,N_32831,N_32897);
nor U33001 (N_33001,N_32952,N_32944);
xnor U33002 (N_33002,N_32966,N_32950);
nand U33003 (N_33003,N_32829,N_32888);
nor U33004 (N_33004,N_32968,N_32800);
nand U33005 (N_33005,N_32982,N_32791);
nor U33006 (N_33006,N_32814,N_32846);
and U33007 (N_33007,N_32927,N_32844);
xnor U33008 (N_33008,N_32917,N_32894);
nor U33009 (N_33009,N_32896,N_32793);
and U33010 (N_33010,N_32990,N_32902);
and U33011 (N_33011,N_32822,N_32879);
or U33012 (N_33012,N_32840,N_32853);
xor U33013 (N_33013,N_32889,N_32936);
or U33014 (N_33014,N_32898,N_32880);
and U33015 (N_33015,N_32816,N_32807);
or U33016 (N_33016,N_32905,N_32869);
or U33017 (N_33017,N_32995,N_32901);
or U33018 (N_33018,N_32969,N_32983);
or U33019 (N_33019,N_32752,N_32811);
xnor U33020 (N_33020,N_32953,N_32942);
and U33021 (N_33021,N_32970,N_32866);
nand U33022 (N_33022,N_32997,N_32923);
and U33023 (N_33023,N_32890,N_32813);
nand U33024 (N_33024,N_32922,N_32792);
and U33025 (N_33025,N_32833,N_32946);
and U33026 (N_33026,N_32921,N_32838);
nand U33027 (N_33027,N_32938,N_32918);
and U33028 (N_33028,N_32994,N_32940);
xor U33029 (N_33029,N_32836,N_32868);
and U33030 (N_33030,N_32786,N_32843);
and U33031 (N_33031,N_32911,N_32785);
nand U33032 (N_33032,N_32993,N_32788);
or U33033 (N_33033,N_32783,N_32850);
xor U33034 (N_33034,N_32998,N_32847);
or U33035 (N_33035,N_32766,N_32954);
xor U33036 (N_33036,N_32956,N_32958);
or U33037 (N_33037,N_32988,N_32774);
or U33038 (N_33038,N_32755,N_32949);
or U33039 (N_33039,N_32903,N_32961);
and U33040 (N_33040,N_32820,N_32775);
xor U33041 (N_33041,N_32893,N_32874);
xnor U33042 (N_33042,N_32830,N_32773);
nor U33043 (N_33043,N_32935,N_32803);
and U33044 (N_33044,N_32873,N_32828);
nand U33045 (N_33045,N_32857,N_32981);
xor U33046 (N_33046,N_32959,N_32799);
or U33047 (N_33047,N_32900,N_32978);
and U33048 (N_33048,N_32787,N_32794);
nor U33049 (N_33049,N_32849,N_32863);
nand U33050 (N_33050,N_32985,N_32928);
nor U33051 (N_33051,N_32835,N_32852);
xnor U33052 (N_33052,N_32907,N_32915);
xnor U33053 (N_33053,N_32974,N_32967);
xor U33054 (N_33054,N_32996,N_32804);
and U33055 (N_33055,N_32842,N_32817);
and U33056 (N_33056,N_32832,N_32826);
xor U33057 (N_33057,N_32945,N_32904);
nand U33058 (N_33058,N_32808,N_32761);
and U33059 (N_33059,N_32939,N_32845);
xor U33060 (N_33060,N_32906,N_32875);
xor U33061 (N_33061,N_32823,N_32815);
xor U33062 (N_33062,N_32963,N_32976);
xor U33063 (N_33063,N_32914,N_32769);
nor U33064 (N_33064,N_32760,N_32979);
or U33065 (N_33065,N_32870,N_32877);
nor U33066 (N_33066,N_32934,N_32884);
nand U33067 (N_33067,N_32802,N_32876);
or U33068 (N_33068,N_32933,N_32790);
and U33069 (N_33069,N_32782,N_32991);
or U33070 (N_33070,N_32768,N_32951);
nor U33071 (N_33071,N_32763,N_32930);
xor U33072 (N_33072,N_32926,N_32882);
nand U33073 (N_33073,N_32809,N_32765);
and U33074 (N_33074,N_32859,N_32973);
and U33075 (N_33075,N_32806,N_32908);
nand U33076 (N_33076,N_32778,N_32964);
or U33077 (N_33077,N_32771,N_32781);
and U33078 (N_33078,N_32941,N_32955);
nor U33079 (N_33079,N_32916,N_32795);
nand U33080 (N_33080,N_32762,N_32758);
xor U33081 (N_33081,N_32909,N_32932);
xor U33082 (N_33082,N_32891,N_32839);
and U33083 (N_33083,N_32848,N_32892);
xor U33084 (N_33084,N_32784,N_32984);
nor U33085 (N_33085,N_32919,N_32797);
nand U33086 (N_33086,N_32925,N_32818);
and U33087 (N_33087,N_32885,N_32862);
nand U33088 (N_33088,N_32929,N_32948);
nor U33089 (N_33089,N_32812,N_32810);
xor U33090 (N_33090,N_32759,N_32780);
or U33091 (N_33091,N_32871,N_32867);
nand U33092 (N_33092,N_32856,N_32855);
nand U33093 (N_33093,N_32750,N_32858);
xnor U33094 (N_33094,N_32872,N_32878);
nor U33095 (N_33095,N_32931,N_32913);
and U33096 (N_33096,N_32824,N_32851);
nor U33097 (N_33097,N_32825,N_32779);
and U33098 (N_33098,N_32819,N_32960);
or U33099 (N_33099,N_32772,N_32798);
xnor U33100 (N_33100,N_32764,N_32756);
and U33101 (N_33101,N_32860,N_32751);
nor U33102 (N_33102,N_32789,N_32883);
nor U33103 (N_33103,N_32767,N_32947);
and U33104 (N_33104,N_32972,N_32886);
and U33105 (N_33105,N_32992,N_32753);
and U33106 (N_33106,N_32912,N_32841);
nor U33107 (N_33107,N_32754,N_32899);
or U33108 (N_33108,N_32777,N_32943);
and U33109 (N_33109,N_32971,N_32920);
and U33110 (N_33110,N_32975,N_32910);
and U33111 (N_33111,N_32821,N_32757);
nand U33112 (N_33112,N_32801,N_32861);
or U33113 (N_33113,N_32881,N_32796);
nand U33114 (N_33114,N_32980,N_32776);
nand U33115 (N_33115,N_32962,N_32834);
and U33116 (N_33116,N_32865,N_32987);
xor U33117 (N_33117,N_32864,N_32937);
or U33118 (N_33118,N_32827,N_32957);
and U33119 (N_33119,N_32989,N_32770);
nand U33120 (N_33120,N_32837,N_32924);
and U33121 (N_33121,N_32999,N_32977);
nor U33122 (N_33122,N_32895,N_32965);
nand U33123 (N_33123,N_32887,N_32986);
and U33124 (N_33124,N_32854,N_32805);
or U33125 (N_33125,N_32903,N_32814);
and U33126 (N_33126,N_32867,N_32900);
nor U33127 (N_33127,N_32854,N_32979);
and U33128 (N_33128,N_32857,N_32990);
and U33129 (N_33129,N_32957,N_32792);
xor U33130 (N_33130,N_32769,N_32759);
nand U33131 (N_33131,N_32857,N_32849);
and U33132 (N_33132,N_32763,N_32832);
nand U33133 (N_33133,N_32876,N_32939);
xnor U33134 (N_33134,N_32977,N_32932);
xnor U33135 (N_33135,N_32933,N_32980);
or U33136 (N_33136,N_32975,N_32822);
or U33137 (N_33137,N_32961,N_32901);
nand U33138 (N_33138,N_32778,N_32936);
or U33139 (N_33139,N_32750,N_32953);
nor U33140 (N_33140,N_32932,N_32970);
nand U33141 (N_33141,N_32775,N_32756);
or U33142 (N_33142,N_32767,N_32847);
or U33143 (N_33143,N_32784,N_32965);
nor U33144 (N_33144,N_32916,N_32875);
xnor U33145 (N_33145,N_32958,N_32995);
and U33146 (N_33146,N_32881,N_32921);
nor U33147 (N_33147,N_32803,N_32994);
and U33148 (N_33148,N_32995,N_32951);
nand U33149 (N_33149,N_32812,N_32934);
or U33150 (N_33150,N_32966,N_32817);
and U33151 (N_33151,N_32994,N_32795);
or U33152 (N_33152,N_32900,N_32928);
or U33153 (N_33153,N_32914,N_32889);
nor U33154 (N_33154,N_32798,N_32845);
and U33155 (N_33155,N_32785,N_32864);
nand U33156 (N_33156,N_32914,N_32991);
xor U33157 (N_33157,N_32959,N_32956);
or U33158 (N_33158,N_32972,N_32917);
nand U33159 (N_33159,N_32812,N_32992);
xor U33160 (N_33160,N_32891,N_32772);
nor U33161 (N_33161,N_32783,N_32928);
nand U33162 (N_33162,N_32905,N_32906);
nor U33163 (N_33163,N_32871,N_32837);
nor U33164 (N_33164,N_32982,N_32766);
nand U33165 (N_33165,N_32888,N_32849);
nor U33166 (N_33166,N_32847,N_32759);
xnor U33167 (N_33167,N_32780,N_32754);
xor U33168 (N_33168,N_32958,N_32915);
or U33169 (N_33169,N_32915,N_32976);
and U33170 (N_33170,N_32830,N_32931);
nand U33171 (N_33171,N_32760,N_32978);
nand U33172 (N_33172,N_32793,N_32829);
nand U33173 (N_33173,N_32894,N_32789);
and U33174 (N_33174,N_32762,N_32993);
xnor U33175 (N_33175,N_32838,N_32770);
or U33176 (N_33176,N_32870,N_32780);
and U33177 (N_33177,N_32997,N_32761);
nor U33178 (N_33178,N_32894,N_32783);
nor U33179 (N_33179,N_32776,N_32903);
nand U33180 (N_33180,N_32927,N_32911);
or U33181 (N_33181,N_32896,N_32954);
xor U33182 (N_33182,N_32915,N_32889);
nand U33183 (N_33183,N_32814,N_32966);
nand U33184 (N_33184,N_32785,N_32959);
and U33185 (N_33185,N_32874,N_32834);
xor U33186 (N_33186,N_32780,N_32787);
and U33187 (N_33187,N_32840,N_32944);
xnor U33188 (N_33188,N_32798,N_32806);
nand U33189 (N_33189,N_32757,N_32781);
nor U33190 (N_33190,N_32935,N_32757);
nor U33191 (N_33191,N_32875,N_32808);
and U33192 (N_33192,N_32944,N_32760);
nor U33193 (N_33193,N_32873,N_32896);
nand U33194 (N_33194,N_32832,N_32872);
or U33195 (N_33195,N_32971,N_32821);
xnor U33196 (N_33196,N_32969,N_32943);
nor U33197 (N_33197,N_32974,N_32917);
nor U33198 (N_33198,N_32786,N_32988);
nand U33199 (N_33199,N_32862,N_32999);
or U33200 (N_33200,N_32881,N_32943);
nor U33201 (N_33201,N_32995,N_32917);
or U33202 (N_33202,N_32780,N_32792);
or U33203 (N_33203,N_32907,N_32956);
nor U33204 (N_33204,N_32911,N_32930);
and U33205 (N_33205,N_32905,N_32789);
and U33206 (N_33206,N_32842,N_32929);
or U33207 (N_33207,N_32751,N_32822);
xor U33208 (N_33208,N_32876,N_32962);
nand U33209 (N_33209,N_32850,N_32810);
or U33210 (N_33210,N_32920,N_32974);
xnor U33211 (N_33211,N_32887,N_32768);
xnor U33212 (N_33212,N_32980,N_32773);
and U33213 (N_33213,N_32965,N_32966);
xor U33214 (N_33214,N_32973,N_32926);
xor U33215 (N_33215,N_32923,N_32932);
nor U33216 (N_33216,N_32855,N_32835);
nand U33217 (N_33217,N_32914,N_32906);
xnor U33218 (N_33218,N_32867,N_32786);
or U33219 (N_33219,N_32901,N_32952);
or U33220 (N_33220,N_32844,N_32848);
or U33221 (N_33221,N_32819,N_32942);
nand U33222 (N_33222,N_32758,N_32812);
nand U33223 (N_33223,N_32965,N_32887);
xor U33224 (N_33224,N_32758,N_32991);
or U33225 (N_33225,N_32940,N_32793);
or U33226 (N_33226,N_32763,N_32865);
nand U33227 (N_33227,N_32898,N_32823);
xnor U33228 (N_33228,N_32796,N_32874);
nor U33229 (N_33229,N_32808,N_32787);
nand U33230 (N_33230,N_32840,N_32755);
or U33231 (N_33231,N_32903,N_32857);
nand U33232 (N_33232,N_32793,N_32920);
nand U33233 (N_33233,N_32872,N_32866);
nor U33234 (N_33234,N_32831,N_32989);
or U33235 (N_33235,N_32937,N_32911);
and U33236 (N_33236,N_32781,N_32922);
nor U33237 (N_33237,N_32964,N_32848);
nand U33238 (N_33238,N_32874,N_32933);
nor U33239 (N_33239,N_32910,N_32926);
and U33240 (N_33240,N_32812,N_32853);
nand U33241 (N_33241,N_32960,N_32846);
and U33242 (N_33242,N_32985,N_32983);
or U33243 (N_33243,N_32969,N_32809);
or U33244 (N_33244,N_32911,N_32845);
or U33245 (N_33245,N_32844,N_32879);
or U33246 (N_33246,N_32877,N_32827);
and U33247 (N_33247,N_32775,N_32815);
and U33248 (N_33248,N_32913,N_32861);
nor U33249 (N_33249,N_32757,N_32770);
xor U33250 (N_33250,N_33147,N_33130);
or U33251 (N_33251,N_33207,N_33110);
nor U33252 (N_33252,N_33043,N_33173);
nand U33253 (N_33253,N_33119,N_33148);
and U33254 (N_33254,N_33180,N_33052);
nor U33255 (N_33255,N_33181,N_33131);
nand U33256 (N_33256,N_33249,N_33112);
xor U33257 (N_33257,N_33023,N_33103);
nand U33258 (N_33258,N_33127,N_33111);
nand U33259 (N_33259,N_33172,N_33101);
and U33260 (N_33260,N_33033,N_33085);
nand U33261 (N_33261,N_33053,N_33109);
or U33262 (N_33262,N_33229,N_33062);
xnor U33263 (N_33263,N_33107,N_33201);
or U33264 (N_33264,N_33209,N_33047);
and U33265 (N_33265,N_33214,N_33219);
nor U33266 (N_33266,N_33097,N_33169);
and U33267 (N_33267,N_33026,N_33046);
and U33268 (N_33268,N_33223,N_33149);
nor U33269 (N_33269,N_33012,N_33082);
and U33270 (N_33270,N_33091,N_33065);
xnor U33271 (N_33271,N_33210,N_33032);
and U33272 (N_33272,N_33151,N_33071);
nand U33273 (N_33273,N_33126,N_33038);
nand U33274 (N_33274,N_33141,N_33197);
nand U33275 (N_33275,N_33029,N_33213);
or U33276 (N_33276,N_33000,N_33017);
nand U33277 (N_33277,N_33129,N_33054);
or U33278 (N_33278,N_33005,N_33189);
or U33279 (N_33279,N_33024,N_33123);
nand U33280 (N_33280,N_33102,N_33184);
xnor U33281 (N_33281,N_33079,N_33217);
nand U33282 (N_33282,N_33113,N_33146);
xnor U33283 (N_33283,N_33188,N_33004);
nor U33284 (N_33284,N_33028,N_33218);
nand U33285 (N_33285,N_33124,N_33185);
nor U33286 (N_33286,N_33084,N_33204);
or U33287 (N_33287,N_33042,N_33118);
nor U33288 (N_33288,N_33211,N_33049);
and U33289 (N_33289,N_33137,N_33060);
nor U33290 (N_33290,N_33171,N_33178);
nor U33291 (N_33291,N_33067,N_33075);
nand U33292 (N_33292,N_33036,N_33238);
or U33293 (N_33293,N_33064,N_33006);
or U33294 (N_33294,N_33048,N_33095);
nor U33295 (N_33295,N_33206,N_33233);
or U33296 (N_33296,N_33231,N_33163);
or U33297 (N_33297,N_33096,N_33212);
xor U33298 (N_33298,N_33037,N_33244);
and U33299 (N_33299,N_33132,N_33059);
nand U33300 (N_33300,N_33224,N_33108);
nor U33301 (N_33301,N_33166,N_33045);
nor U33302 (N_33302,N_33168,N_33125);
nand U33303 (N_33303,N_33240,N_33236);
nor U33304 (N_33304,N_33035,N_33155);
nor U33305 (N_33305,N_33070,N_33083);
nor U33306 (N_33306,N_33200,N_33235);
xor U33307 (N_33307,N_33039,N_33220);
nand U33308 (N_33308,N_33199,N_33022);
or U33309 (N_33309,N_33202,N_33056);
nor U33310 (N_33310,N_33159,N_33139);
or U33311 (N_33311,N_33226,N_33078);
xnor U33312 (N_33312,N_33007,N_33228);
nand U33313 (N_33313,N_33088,N_33100);
and U33314 (N_33314,N_33192,N_33058);
nand U33315 (N_33315,N_33241,N_33165);
nor U33316 (N_33316,N_33034,N_33183);
nand U33317 (N_33317,N_33208,N_33066);
and U33318 (N_33318,N_33089,N_33117);
and U33319 (N_33319,N_33162,N_33156);
xor U33320 (N_33320,N_33086,N_33080);
nor U33321 (N_33321,N_33248,N_33010);
or U33322 (N_33322,N_33073,N_33121);
nor U33323 (N_33323,N_33152,N_33051);
and U33324 (N_33324,N_33044,N_33225);
xnor U33325 (N_33325,N_33069,N_33143);
xor U33326 (N_33326,N_33128,N_33177);
xor U33327 (N_33327,N_33215,N_33187);
nand U33328 (N_33328,N_33190,N_33134);
nand U33329 (N_33329,N_33003,N_33205);
nor U33330 (N_33330,N_33114,N_33041);
nor U33331 (N_33331,N_33232,N_33013);
xnor U33332 (N_33332,N_33120,N_33179);
nand U33333 (N_33333,N_33090,N_33182);
and U33334 (N_33334,N_33170,N_33196);
xor U33335 (N_33335,N_33167,N_33105);
xnor U33336 (N_33336,N_33245,N_33175);
or U33337 (N_33337,N_33216,N_33153);
and U33338 (N_33338,N_33222,N_33040);
or U33339 (N_33339,N_33161,N_33001);
nor U33340 (N_33340,N_33239,N_33016);
xor U33341 (N_33341,N_33057,N_33027);
xnor U33342 (N_33342,N_33186,N_33176);
and U33343 (N_33343,N_33242,N_33191);
nand U33344 (N_33344,N_33099,N_33140);
nor U33345 (N_33345,N_33092,N_33025);
and U33346 (N_33346,N_33104,N_33020);
or U33347 (N_33347,N_33063,N_33227);
nor U33348 (N_33348,N_33009,N_33158);
nor U33349 (N_33349,N_33154,N_33106);
nand U33350 (N_33350,N_33122,N_33087);
and U33351 (N_33351,N_33098,N_33174);
xor U33352 (N_33352,N_33061,N_33203);
and U33353 (N_33353,N_33142,N_33195);
nor U33354 (N_33354,N_33150,N_33074);
nor U33355 (N_33355,N_33076,N_33077);
nor U33356 (N_33356,N_33014,N_33237);
and U33357 (N_33357,N_33050,N_33008);
nor U33358 (N_33358,N_33030,N_33138);
nand U33359 (N_33359,N_33068,N_33157);
nand U33360 (N_33360,N_33135,N_33116);
and U33361 (N_33361,N_33221,N_33194);
nand U33362 (N_33362,N_33031,N_33072);
or U33363 (N_33363,N_33015,N_33011);
and U33364 (N_33364,N_33164,N_33094);
nor U33365 (N_33365,N_33133,N_33115);
nor U33366 (N_33366,N_33093,N_33144);
xnor U33367 (N_33367,N_33230,N_33246);
nor U33368 (N_33368,N_33002,N_33243);
or U33369 (N_33369,N_33018,N_33247);
xnor U33370 (N_33370,N_33081,N_33019);
xnor U33371 (N_33371,N_33021,N_33145);
and U33372 (N_33372,N_33234,N_33193);
nor U33373 (N_33373,N_33055,N_33136);
nor U33374 (N_33374,N_33198,N_33160);
and U33375 (N_33375,N_33158,N_33083);
xor U33376 (N_33376,N_33130,N_33003);
and U33377 (N_33377,N_33023,N_33127);
nor U33378 (N_33378,N_33014,N_33090);
nand U33379 (N_33379,N_33087,N_33187);
xor U33380 (N_33380,N_33057,N_33210);
nand U33381 (N_33381,N_33236,N_33216);
or U33382 (N_33382,N_33242,N_33225);
nand U33383 (N_33383,N_33100,N_33183);
and U33384 (N_33384,N_33204,N_33217);
xor U33385 (N_33385,N_33197,N_33051);
or U33386 (N_33386,N_33068,N_33161);
and U33387 (N_33387,N_33025,N_33087);
nor U33388 (N_33388,N_33139,N_33249);
and U33389 (N_33389,N_33225,N_33017);
nand U33390 (N_33390,N_33142,N_33082);
nor U33391 (N_33391,N_33127,N_33128);
or U33392 (N_33392,N_33075,N_33219);
nor U33393 (N_33393,N_33011,N_33164);
xor U33394 (N_33394,N_33114,N_33050);
or U33395 (N_33395,N_33195,N_33113);
or U33396 (N_33396,N_33107,N_33106);
nor U33397 (N_33397,N_33017,N_33147);
nor U33398 (N_33398,N_33011,N_33052);
xnor U33399 (N_33399,N_33217,N_33036);
and U33400 (N_33400,N_33196,N_33243);
nand U33401 (N_33401,N_33070,N_33043);
and U33402 (N_33402,N_33221,N_33019);
and U33403 (N_33403,N_33218,N_33247);
or U33404 (N_33404,N_33170,N_33239);
nand U33405 (N_33405,N_33007,N_33095);
or U33406 (N_33406,N_33100,N_33102);
and U33407 (N_33407,N_33032,N_33163);
nor U33408 (N_33408,N_33054,N_33128);
xnor U33409 (N_33409,N_33023,N_33172);
nand U33410 (N_33410,N_33183,N_33028);
or U33411 (N_33411,N_33236,N_33031);
xor U33412 (N_33412,N_33049,N_33230);
xor U33413 (N_33413,N_33153,N_33018);
and U33414 (N_33414,N_33249,N_33230);
nand U33415 (N_33415,N_33182,N_33132);
nor U33416 (N_33416,N_33157,N_33083);
nand U33417 (N_33417,N_33101,N_33163);
and U33418 (N_33418,N_33132,N_33108);
nor U33419 (N_33419,N_33147,N_33165);
xor U33420 (N_33420,N_33061,N_33207);
nor U33421 (N_33421,N_33132,N_33214);
or U33422 (N_33422,N_33190,N_33233);
or U33423 (N_33423,N_33040,N_33198);
nor U33424 (N_33424,N_33096,N_33058);
and U33425 (N_33425,N_33137,N_33157);
xnor U33426 (N_33426,N_33067,N_33193);
nor U33427 (N_33427,N_33236,N_33156);
and U33428 (N_33428,N_33079,N_33121);
nand U33429 (N_33429,N_33033,N_33090);
or U33430 (N_33430,N_33103,N_33128);
nor U33431 (N_33431,N_33084,N_33156);
nor U33432 (N_33432,N_33010,N_33247);
and U33433 (N_33433,N_33170,N_33191);
and U33434 (N_33434,N_33184,N_33131);
nand U33435 (N_33435,N_33228,N_33243);
nand U33436 (N_33436,N_33224,N_33188);
nor U33437 (N_33437,N_33084,N_33001);
xnor U33438 (N_33438,N_33155,N_33090);
or U33439 (N_33439,N_33117,N_33001);
nor U33440 (N_33440,N_33148,N_33111);
xor U33441 (N_33441,N_33168,N_33025);
xnor U33442 (N_33442,N_33201,N_33128);
or U33443 (N_33443,N_33117,N_33044);
and U33444 (N_33444,N_33155,N_33076);
nor U33445 (N_33445,N_33018,N_33173);
nand U33446 (N_33446,N_33185,N_33143);
nor U33447 (N_33447,N_33232,N_33008);
and U33448 (N_33448,N_33217,N_33059);
and U33449 (N_33449,N_33231,N_33239);
xor U33450 (N_33450,N_33218,N_33147);
nor U33451 (N_33451,N_33225,N_33223);
nand U33452 (N_33452,N_33104,N_33095);
and U33453 (N_33453,N_33195,N_33151);
and U33454 (N_33454,N_33107,N_33076);
nand U33455 (N_33455,N_33105,N_33149);
or U33456 (N_33456,N_33116,N_33176);
nor U33457 (N_33457,N_33099,N_33063);
nor U33458 (N_33458,N_33064,N_33140);
xor U33459 (N_33459,N_33204,N_33047);
or U33460 (N_33460,N_33028,N_33076);
nand U33461 (N_33461,N_33216,N_33008);
nor U33462 (N_33462,N_33174,N_33100);
and U33463 (N_33463,N_33205,N_33096);
nand U33464 (N_33464,N_33086,N_33206);
or U33465 (N_33465,N_33239,N_33228);
and U33466 (N_33466,N_33117,N_33015);
xnor U33467 (N_33467,N_33086,N_33051);
or U33468 (N_33468,N_33023,N_33217);
nand U33469 (N_33469,N_33151,N_33154);
or U33470 (N_33470,N_33131,N_33202);
xnor U33471 (N_33471,N_33000,N_33043);
nand U33472 (N_33472,N_33129,N_33103);
nand U33473 (N_33473,N_33098,N_33166);
or U33474 (N_33474,N_33125,N_33181);
and U33475 (N_33475,N_33088,N_33040);
and U33476 (N_33476,N_33104,N_33155);
or U33477 (N_33477,N_33244,N_33231);
nand U33478 (N_33478,N_33024,N_33015);
or U33479 (N_33479,N_33092,N_33056);
and U33480 (N_33480,N_33171,N_33247);
nor U33481 (N_33481,N_33123,N_33246);
xnor U33482 (N_33482,N_33088,N_33208);
xnor U33483 (N_33483,N_33144,N_33024);
xnor U33484 (N_33484,N_33218,N_33222);
nor U33485 (N_33485,N_33025,N_33216);
and U33486 (N_33486,N_33224,N_33150);
xnor U33487 (N_33487,N_33086,N_33237);
and U33488 (N_33488,N_33207,N_33006);
nand U33489 (N_33489,N_33150,N_33111);
xnor U33490 (N_33490,N_33104,N_33013);
or U33491 (N_33491,N_33103,N_33082);
or U33492 (N_33492,N_33023,N_33234);
nor U33493 (N_33493,N_33075,N_33178);
xnor U33494 (N_33494,N_33045,N_33138);
and U33495 (N_33495,N_33014,N_33081);
or U33496 (N_33496,N_33196,N_33030);
and U33497 (N_33497,N_33077,N_33075);
nand U33498 (N_33498,N_33088,N_33113);
nand U33499 (N_33499,N_33182,N_33183);
and U33500 (N_33500,N_33436,N_33319);
or U33501 (N_33501,N_33454,N_33252);
nor U33502 (N_33502,N_33293,N_33484);
or U33503 (N_33503,N_33401,N_33276);
or U33504 (N_33504,N_33299,N_33289);
and U33505 (N_33505,N_33439,N_33441);
or U33506 (N_33506,N_33256,N_33492);
nand U33507 (N_33507,N_33445,N_33434);
nand U33508 (N_33508,N_33327,N_33368);
nor U33509 (N_33509,N_33452,N_33392);
and U33510 (N_33510,N_33433,N_33424);
nor U33511 (N_33511,N_33385,N_33339);
nand U33512 (N_33512,N_33334,N_33440);
xor U33513 (N_33513,N_33271,N_33371);
nand U33514 (N_33514,N_33481,N_33331);
nand U33515 (N_33515,N_33325,N_33322);
xnor U33516 (N_33516,N_33329,N_33386);
nor U33517 (N_33517,N_33423,N_33266);
nand U33518 (N_33518,N_33475,N_33474);
nor U33519 (N_33519,N_33328,N_33302);
and U33520 (N_33520,N_33451,N_33402);
xnor U33521 (N_33521,N_33430,N_33410);
and U33522 (N_33522,N_33312,N_33347);
nor U33523 (N_33523,N_33477,N_33485);
xor U33524 (N_33524,N_33429,N_33437);
xnor U33525 (N_33525,N_33333,N_33294);
and U33526 (N_33526,N_33316,N_33487);
nand U33527 (N_33527,N_33438,N_33335);
nand U33528 (N_33528,N_33281,N_33343);
xor U33529 (N_33529,N_33342,N_33444);
xor U33530 (N_33530,N_33262,N_33403);
nor U33531 (N_33531,N_33303,N_33382);
and U33532 (N_33532,N_33310,N_33283);
and U33533 (N_33533,N_33432,N_33446);
nand U33534 (N_33534,N_33355,N_33388);
nor U33535 (N_33535,N_33469,N_33273);
and U33536 (N_33536,N_33390,N_33336);
xnor U33537 (N_33537,N_33408,N_33473);
or U33538 (N_33538,N_33398,N_33391);
or U33539 (N_33539,N_33380,N_33397);
and U33540 (N_33540,N_33447,N_33365);
nor U33541 (N_33541,N_33460,N_33407);
nand U33542 (N_33542,N_33313,N_33478);
xnor U33543 (N_33543,N_33340,N_33346);
nor U33544 (N_33544,N_33349,N_33415);
or U33545 (N_33545,N_33458,N_33428);
and U33546 (N_33546,N_33277,N_33288);
nor U33547 (N_33547,N_33358,N_33264);
or U33548 (N_33548,N_33418,N_33462);
and U33549 (N_33549,N_33321,N_33364);
nor U33550 (N_33550,N_33389,N_33298);
xnor U33551 (N_33551,N_33274,N_33268);
xnor U33552 (N_33552,N_33459,N_33400);
or U33553 (N_33553,N_33307,N_33466);
and U33554 (N_33554,N_33431,N_33409);
and U33555 (N_33555,N_33304,N_33383);
nand U33556 (N_33556,N_33381,N_33270);
and U33557 (N_33557,N_33330,N_33300);
nand U33558 (N_33558,N_33396,N_33356);
nor U33559 (N_33559,N_33311,N_33297);
xnor U33560 (N_33560,N_33292,N_33414);
and U33561 (N_33561,N_33348,N_33287);
nor U33562 (N_33562,N_33326,N_33366);
or U33563 (N_33563,N_33282,N_33419);
xnor U33564 (N_33564,N_33370,N_33426);
or U33565 (N_33565,N_33305,N_33332);
xnor U33566 (N_33566,N_33253,N_33279);
nor U33567 (N_33567,N_33306,N_33496);
and U33568 (N_33568,N_33375,N_33448);
xor U33569 (N_33569,N_33280,N_33412);
nor U33570 (N_33570,N_33353,N_33317);
or U33571 (N_33571,N_33269,N_33422);
or U33572 (N_33572,N_33463,N_33362);
nand U33573 (N_33573,N_33373,N_33449);
or U33574 (N_33574,N_33479,N_33495);
nor U33575 (N_33575,N_33296,N_33338);
or U33576 (N_33576,N_33251,N_33351);
nor U33577 (N_33577,N_33341,N_33387);
and U33578 (N_33578,N_33378,N_33499);
xnor U33579 (N_33579,N_33494,N_33405);
xnor U33580 (N_33580,N_33361,N_33411);
nor U33581 (N_33581,N_33257,N_33465);
and U33582 (N_33582,N_33421,N_33435);
xor U33583 (N_33583,N_33472,N_33301);
xor U33584 (N_33584,N_33272,N_33291);
or U33585 (N_33585,N_33467,N_33489);
or U33586 (N_33586,N_33377,N_33374);
xor U33587 (N_33587,N_33324,N_33425);
nand U33588 (N_33588,N_33278,N_33265);
or U33589 (N_33589,N_33309,N_33285);
xor U33590 (N_33590,N_33320,N_33345);
or U33591 (N_33591,N_33295,N_33394);
nand U33592 (N_33592,N_33443,N_33267);
or U33593 (N_33593,N_33399,N_33357);
nand U33594 (N_33594,N_33486,N_33350);
and U33595 (N_33595,N_33490,N_33369);
nor U33596 (N_33596,N_33470,N_33286);
and U33597 (N_33597,N_33261,N_33488);
nand U33598 (N_33598,N_33354,N_33404);
nand U33599 (N_33599,N_33498,N_33254);
and U33600 (N_33600,N_33427,N_33315);
nor U33601 (N_33601,N_33420,N_33406);
nand U33602 (N_33602,N_33360,N_33260);
or U33603 (N_33603,N_33482,N_33417);
and U33604 (N_33604,N_33461,N_33367);
and U33605 (N_33605,N_33259,N_33250);
xnor U33606 (N_33606,N_33455,N_33290);
and U33607 (N_33607,N_33258,N_33363);
or U33608 (N_33608,N_33413,N_33464);
or U33609 (N_33609,N_33497,N_33491);
or U33610 (N_33610,N_33359,N_33255);
nor U33611 (N_33611,N_33352,N_33476);
nand U33612 (N_33612,N_33323,N_33480);
nor U33613 (N_33613,N_33376,N_33395);
xnor U33614 (N_33614,N_33275,N_33263);
nand U33615 (N_33615,N_33393,N_33372);
and U33616 (N_33616,N_33416,N_33284);
nand U33617 (N_33617,N_33471,N_33450);
xnor U33618 (N_33618,N_33493,N_33379);
nor U33619 (N_33619,N_33384,N_33457);
nand U33620 (N_33620,N_33453,N_33318);
or U33621 (N_33621,N_33337,N_33308);
xor U33622 (N_33622,N_33344,N_33314);
nand U33623 (N_33623,N_33483,N_33456);
xor U33624 (N_33624,N_33468,N_33442);
nor U33625 (N_33625,N_33481,N_33407);
nand U33626 (N_33626,N_33452,N_33490);
nand U33627 (N_33627,N_33438,N_33303);
or U33628 (N_33628,N_33283,N_33404);
or U33629 (N_33629,N_33450,N_33273);
nor U33630 (N_33630,N_33272,N_33304);
xor U33631 (N_33631,N_33307,N_33439);
and U33632 (N_33632,N_33250,N_33283);
and U33633 (N_33633,N_33332,N_33361);
or U33634 (N_33634,N_33311,N_33439);
nand U33635 (N_33635,N_33291,N_33298);
and U33636 (N_33636,N_33396,N_33486);
or U33637 (N_33637,N_33337,N_33398);
and U33638 (N_33638,N_33265,N_33274);
nor U33639 (N_33639,N_33283,N_33290);
and U33640 (N_33640,N_33395,N_33436);
or U33641 (N_33641,N_33349,N_33275);
and U33642 (N_33642,N_33480,N_33254);
or U33643 (N_33643,N_33456,N_33494);
xnor U33644 (N_33644,N_33432,N_33360);
nand U33645 (N_33645,N_33326,N_33406);
or U33646 (N_33646,N_33466,N_33330);
nor U33647 (N_33647,N_33334,N_33253);
and U33648 (N_33648,N_33265,N_33289);
and U33649 (N_33649,N_33360,N_33435);
nor U33650 (N_33650,N_33465,N_33363);
or U33651 (N_33651,N_33305,N_33462);
or U33652 (N_33652,N_33499,N_33387);
and U33653 (N_33653,N_33409,N_33392);
xor U33654 (N_33654,N_33283,N_33370);
and U33655 (N_33655,N_33452,N_33338);
and U33656 (N_33656,N_33413,N_33486);
nor U33657 (N_33657,N_33253,N_33296);
and U33658 (N_33658,N_33447,N_33384);
nor U33659 (N_33659,N_33339,N_33331);
nor U33660 (N_33660,N_33283,N_33418);
nor U33661 (N_33661,N_33393,N_33317);
xnor U33662 (N_33662,N_33464,N_33475);
nor U33663 (N_33663,N_33306,N_33488);
nand U33664 (N_33664,N_33399,N_33466);
or U33665 (N_33665,N_33406,N_33444);
or U33666 (N_33666,N_33300,N_33340);
xnor U33667 (N_33667,N_33432,N_33261);
nand U33668 (N_33668,N_33420,N_33347);
nor U33669 (N_33669,N_33462,N_33304);
and U33670 (N_33670,N_33325,N_33273);
or U33671 (N_33671,N_33420,N_33375);
and U33672 (N_33672,N_33343,N_33319);
nor U33673 (N_33673,N_33451,N_33490);
and U33674 (N_33674,N_33379,N_33320);
nor U33675 (N_33675,N_33360,N_33330);
and U33676 (N_33676,N_33398,N_33330);
xor U33677 (N_33677,N_33308,N_33456);
nand U33678 (N_33678,N_33278,N_33389);
xor U33679 (N_33679,N_33382,N_33337);
xnor U33680 (N_33680,N_33416,N_33340);
nand U33681 (N_33681,N_33375,N_33259);
and U33682 (N_33682,N_33293,N_33424);
and U33683 (N_33683,N_33289,N_33490);
or U33684 (N_33684,N_33273,N_33471);
xnor U33685 (N_33685,N_33251,N_33384);
nor U33686 (N_33686,N_33274,N_33311);
xor U33687 (N_33687,N_33334,N_33279);
xnor U33688 (N_33688,N_33399,N_33322);
xnor U33689 (N_33689,N_33331,N_33463);
and U33690 (N_33690,N_33370,N_33305);
nor U33691 (N_33691,N_33399,N_33278);
nor U33692 (N_33692,N_33470,N_33360);
and U33693 (N_33693,N_33335,N_33473);
nor U33694 (N_33694,N_33435,N_33433);
nand U33695 (N_33695,N_33373,N_33374);
nand U33696 (N_33696,N_33489,N_33408);
or U33697 (N_33697,N_33420,N_33413);
nand U33698 (N_33698,N_33389,N_33363);
xnor U33699 (N_33699,N_33358,N_33412);
or U33700 (N_33700,N_33287,N_33273);
and U33701 (N_33701,N_33464,N_33288);
nor U33702 (N_33702,N_33364,N_33322);
nand U33703 (N_33703,N_33284,N_33333);
xor U33704 (N_33704,N_33423,N_33252);
nor U33705 (N_33705,N_33441,N_33376);
xor U33706 (N_33706,N_33287,N_33340);
and U33707 (N_33707,N_33410,N_33443);
or U33708 (N_33708,N_33479,N_33294);
nor U33709 (N_33709,N_33446,N_33477);
and U33710 (N_33710,N_33396,N_33460);
or U33711 (N_33711,N_33271,N_33452);
nand U33712 (N_33712,N_33382,N_33400);
xnor U33713 (N_33713,N_33435,N_33480);
nor U33714 (N_33714,N_33255,N_33260);
nand U33715 (N_33715,N_33427,N_33400);
nor U33716 (N_33716,N_33466,N_33254);
or U33717 (N_33717,N_33484,N_33449);
or U33718 (N_33718,N_33319,N_33295);
nor U33719 (N_33719,N_33307,N_33392);
or U33720 (N_33720,N_33309,N_33297);
nand U33721 (N_33721,N_33466,N_33491);
nor U33722 (N_33722,N_33416,N_33321);
nand U33723 (N_33723,N_33381,N_33485);
nand U33724 (N_33724,N_33458,N_33375);
xor U33725 (N_33725,N_33307,N_33412);
and U33726 (N_33726,N_33488,N_33397);
nand U33727 (N_33727,N_33486,N_33292);
nand U33728 (N_33728,N_33257,N_33452);
and U33729 (N_33729,N_33339,N_33327);
nor U33730 (N_33730,N_33344,N_33443);
xnor U33731 (N_33731,N_33288,N_33478);
nand U33732 (N_33732,N_33465,N_33323);
and U33733 (N_33733,N_33399,N_33365);
or U33734 (N_33734,N_33253,N_33264);
and U33735 (N_33735,N_33352,N_33431);
nand U33736 (N_33736,N_33476,N_33397);
or U33737 (N_33737,N_33333,N_33382);
nand U33738 (N_33738,N_33251,N_33482);
nand U33739 (N_33739,N_33272,N_33462);
and U33740 (N_33740,N_33461,N_33293);
or U33741 (N_33741,N_33390,N_33466);
nand U33742 (N_33742,N_33391,N_33326);
nor U33743 (N_33743,N_33351,N_33382);
nor U33744 (N_33744,N_33479,N_33276);
xor U33745 (N_33745,N_33266,N_33380);
and U33746 (N_33746,N_33474,N_33393);
nor U33747 (N_33747,N_33486,N_33379);
nand U33748 (N_33748,N_33445,N_33451);
or U33749 (N_33749,N_33473,N_33455);
or U33750 (N_33750,N_33642,N_33649);
xor U33751 (N_33751,N_33568,N_33559);
nand U33752 (N_33752,N_33575,N_33555);
or U33753 (N_33753,N_33610,N_33669);
nor U33754 (N_33754,N_33604,N_33699);
and U33755 (N_33755,N_33519,N_33724);
and U33756 (N_33756,N_33566,N_33662);
xor U33757 (N_33757,N_33596,N_33525);
and U33758 (N_33758,N_33579,N_33515);
nor U33759 (N_33759,N_33520,N_33599);
xnor U33760 (N_33760,N_33589,N_33622);
nand U33761 (N_33761,N_33574,N_33506);
xor U33762 (N_33762,N_33693,N_33673);
xor U33763 (N_33763,N_33545,N_33625);
nor U33764 (N_33764,N_33563,N_33680);
or U33765 (N_33765,N_33618,N_33517);
or U33766 (N_33766,N_33558,N_33700);
xor U33767 (N_33767,N_33740,N_33733);
nor U33768 (N_33768,N_33727,N_33542);
xnor U33769 (N_33769,N_33514,N_33644);
nor U33770 (N_33770,N_33601,N_33527);
nor U33771 (N_33771,N_33677,N_33573);
nor U33772 (N_33772,N_33634,N_33584);
nand U33773 (N_33773,N_33675,N_33696);
nand U33774 (N_33774,N_33705,N_33684);
nand U33775 (N_33775,N_33683,N_33734);
nor U33776 (N_33776,N_33743,N_33549);
or U33777 (N_33777,N_33729,N_33586);
nand U33778 (N_33778,N_33690,N_33742);
xnor U33779 (N_33779,N_33714,N_33540);
and U33780 (N_33780,N_33702,N_33580);
or U33781 (N_33781,N_33524,N_33614);
nand U33782 (N_33782,N_33713,N_33624);
xor U33783 (N_33783,N_33666,N_33523);
nand U33784 (N_33784,N_33535,N_33674);
or U33785 (N_33785,N_33626,N_33630);
nor U33786 (N_33786,N_33716,N_33651);
or U33787 (N_33787,N_33647,N_33689);
or U33788 (N_33788,N_33537,N_33717);
nand U33789 (N_33789,N_33539,N_33657);
nand U33790 (N_33790,N_33688,N_33613);
and U33791 (N_33791,N_33725,N_33738);
xnor U33792 (N_33792,N_33681,N_33667);
or U33793 (N_33793,N_33578,N_33704);
nand U33794 (N_33794,N_33735,N_33562);
or U33795 (N_33795,N_33569,N_33526);
or U33796 (N_33796,N_33711,N_33576);
or U33797 (N_33797,N_33668,N_33646);
and U33798 (N_33798,N_33736,N_33544);
xor U33799 (N_33799,N_33612,N_33686);
nand U33800 (N_33800,N_33557,N_33664);
xnor U33801 (N_33801,N_33629,N_33739);
nand U33802 (N_33802,N_33726,N_33663);
xor U33803 (N_33803,N_33676,N_33691);
nand U33804 (N_33804,N_33516,N_33749);
nor U33805 (N_33805,N_33590,N_33528);
nor U33806 (N_33806,N_33581,N_33567);
xnor U33807 (N_33807,N_33511,N_33658);
or U33808 (N_33808,N_33744,N_33617);
or U33809 (N_33809,N_33593,N_33572);
and U33810 (N_33810,N_33672,N_33721);
nor U33811 (N_33811,N_33541,N_33747);
and U33812 (N_33812,N_33620,N_33670);
nor U33813 (N_33813,N_33595,N_33678);
and U33814 (N_33814,N_33638,N_33534);
or U33815 (N_33815,N_33718,N_33571);
nor U33816 (N_33816,N_33650,N_33521);
xnor U33817 (N_33817,N_33565,N_33655);
nand U33818 (N_33818,N_33619,N_33654);
or U33819 (N_33819,N_33548,N_33616);
nor U33820 (N_33820,N_33710,N_33732);
nand U33821 (N_33821,N_33697,N_33731);
xor U33822 (N_33822,N_33695,N_33577);
and U33823 (N_33823,N_33640,N_33536);
xnor U33824 (N_33824,N_33635,N_33741);
nor U33825 (N_33825,N_33633,N_33737);
xnor U33826 (N_33826,N_33600,N_33564);
nor U33827 (N_33827,N_33653,N_33685);
nand U33828 (N_33828,N_33728,N_33608);
or U33829 (N_33829,N_33543,N_33546);
and U33830 (N_33830,N_33636,N_33706);
xnor U33831 (N_33831,N_33628,N_33694);
and U33832 (N_33832,N_33708,N_33529);
xor U33833 (N_33833,N_33621,N_33682);
xnor U33834 (N_33834,N_33692,N_33532);
and U33835 (N_33835,N_33585,N_33631);
and U33836 (N_33836,N_33554,N_33550);
or U33837 (N_33837,N_33505,N_33748);
or U33838 (N_33838,N_33551,N_33538);
xnor U33839 (N_33839,N_33518,N_33501);
xor U33840 (N_33840,N_33587,N_33679);
or U33841 (N_33841,N_33513,N_33592);
nand U33842 (N_33842,N_33522,N_33583);
xor U33843 (N_33843,N_33627,N_33507);
and U33844 (N_33844,N_33660,N_33745);
nand U33845 (N_33845,N_33652,N_33656);
and U33846 (N_33846,N_33500,N_33643);
nor U33847 (N_33847,N_33637,N_33645);
and U33848 (N_33848,N_33605,N_33606);
nor U33849 (N_33849,N_33722,N_33530);
nor U33850 (N_33850,N_33598,N_33665);
or U33851 (N_33851,N_33591,N_33509);
and U33852 (N_33852,N_33639,N_33611);
and U33853 (N_33853,N_33531,N_33603);
or U33854 (N_33854,N_33648,N_33671);
nor U33855 (N_33855,N_33632,N_33746);
or U33856 (N_33856,N_33712,N_33730);
and U33857 (N_33857,N_33709,N_33597);
or U33858 (N_33858,N_33607,N_33659);
nand U33859 (N_33859,N_33615,N_33561);
nor U33860 (N_33860,N_33641,N_33552);
nor U33861 (N_33861,N_33687,N_33553);
and U33862 (N_33862,N_33533,N_33547);
and U33863 (N_33863,N_33560,N_33703);
xnor U33864 (N_33864,N_33582,N_33720);
nand U33865 (N_33865,N_33556,N_33661);
nor U33866 (N_33866,N_33508,N_33701);
and U33867 (N_33867,N_33707,N_33715);
or U33868 (N_33868,N_33502,N_33719);
nor U33869 (N_33869,N_33512,N_33623);
nand U33870 (N_33870,N_33588,N_33570);
or U33871 (N_33871,N_33594,N_33602);
nand U33872 (N_33872,N_33609,N_33723);
or U33873 (N_33873,N_33698,N_33510);
xnor U33874 (N_33874,N_33503,N_33504);
nor U33875 (N_33875,N_33567,N_33715);
or U33876 (N_33876,N_33613,N_33737);
and U33877 (N_33877,N_33505,N_33614);
nand U33878 (N_33878,N_33573,N_33601);
nand U33879 (N_33879,N_33628,N_33548);
xor U33880 (N_33880,N_33717,N_33529);
nand U33881 (N_33881,N_33664,N_33680);
nand U33882 (N_33882,N_33743,N_33709);
nor U33883 (N_33883,N_33568,N_33657);
xor U33884 (N_33884,N_33611,N_33593);
nand U33885 (N_33885,N_33635,N_33531);
and U33886 (N_33886,N_33592,N_33593);
nor U33887 (N_33887,N_33693,N_33668);
nand U33888 (N_33888,N_33604,N_33586);
or U33889 (N_33889,N_33688,N_33650);
and U33890 (N_33890,N_33666,N_33531);
and U33891 (N_33891,N_33650,N_33609);
nand U33892 (N_33892,N_33684,N_33503);
and U33893 (N_33893,N_33743,N_33566);
nand U33894 (N_33894,N_33557,N_33564);
nand U33895 (N_33895,N_33561,N_33693);
and U33896 (N_33896,N_33572,N_33630);
xor U33897 (N_33897,N_33663,N_33566);
and U33898 (N_33898,N_33744,N_33588);
nor U33899 (N_33899,N_33664,N_33579);
nor U33900 (N_33900,N_33654,N_33555);
nor U33901 (N_33901,N_33510,N_33719);
and U33902 (N_33902,N_33624,N_33649);
nand U33903 (N_33903,N_33667,N_33622);
or U33904 (N_33904,N_33660,N_33580);
nand U33905 (N_33905,N_33651,N_33745);
nand U33906 (N_33906,N_33576,N_33518);
or U33907 (N_33907,N_33661,N_33571);
and U33908 (N_33908,N_33561,N_33588);
nor U33909 (N_33909,N_33529,N_33605);
or U33910 (N_33910,N_33664,N_33601);
and U33911 (N_33911,N_33714,N_33748);
and U33912 (N_33912,N_33533,N_33501);
or U33913 (N_33913,N_33634,N_33608);
nand U33914 (N_33914,N_33659,N_33616);
nor U33915 (N_33915,N_33598,N_33628);
xnor U33916 (N_33916,N_33678,N_33718);
xor U33917 (N_33917,N_33687,N_33592);
nand U33918 (N_33918,N_33567,N_33632);
xor U33919 (N_33919,N_33674,N_33617);
nand U33920 (N_33920,N_33730,N_33605);
and U33921 (N_33921,N_33628,N_33567);
nor U33922 (N_33922,N_33716,N_33536);
or U33923 (N_33923,N_33545,N_33606);
or U33924 (N_33924,N_33742,N_33668);
and U33925 (N_33925,N_33584,N_33534);
xnor U33926 (N_33926,N_33603,N_33552);
nand U33927 (N_33927,N_33620,N_33739);
and U33928 (N_33928,N_33644,N_33672);
xor U33929 (N_33929,N_33636,N_33569);
xnor U33930 (N_33930,N_33642,N_33519);
nand U33931 (N_33931,N_33704,N_33725);
nand U33932 (N_33932,N_33707,N_33655);
nand U33933 (N_33933,N_33503,N_33702);
or U33934 (N_33934,N_33741,N_33632);
nor U33935 (N_33935,N_33580,N_33697);
xnor U33936 (N_33936,N_33680,N_33671);
or U33937 (N_33937,N_33682,N_33547);
nor U33938 (N_33938,N_33553,N_33613);
nand U33939 (N_33939,N_33729,N_33647);
xnor U33940 (N_33940,N_33671,N_33733);
and U33941 (N_33941,N_33535,N_33582);
nand U33942 (N_33942,N_33715,N_33584);
xnor U33943 (N_33943,N_33619,N_33737);
or U33944 (N_33944,N_33721,N_33565);
xor U33945 (N_33945,N_33594,N_33683);
and U33946 (N_33946,N_33708,N_33550);
or U33947 (N_33947,N_33517,N_33698);
or U33948 (N_33948,N_33620,N_33544);
and U33949 (N_33949,N_33679,N_33747);
xor U33950 (N_33950,N_33695,N_33551);
nor U33951 (N_33951,N_33671,N_33703);
nor U33952 (N_33952,N_33509,N_33741);
or U33953 (N_33953,N_33616,N_33534);
nand U33954 (N_33954,N_33512,N_33589);
nor U33955 (N_33955,N_33660,N_33554);
and U33956 (N_33956,N_33689,N_33626);
or U33957 (N_33957,N_33610,N_33710);
nand U33958 (N_33958,N_33547,N_33516);
xnor U33959 (N_33959,N_33553,N_33653);
or U33960 (N_33960,N_33591,N_33594);
or U33961 (N_33961,N_33525,N_33504);
and U33962 (N_33962,N_33587,N_33602);
and U33963 (N_33963,N_33664,N_33556);
nor U33964 (N_33964,N_33517,N_33659);
nand U33965 (N_33965,N_33745,N_33601);
or U33966 (N_33966,N_33615,N_33600);
and U33967 (N_33967,N_33530,N_33589);
nor U33968 (N_33968,N_33545,N_33568);
xor U33969 (N_33969,N_33544,N_33670);
nor U33970 (N_33970,N_33642,N_33617);
nand U33971 (N_33971,N_33654,N_33536);
xnor U33972 (N_33972,N_33535,N_33745);
nand U33973 (N_33973,N_33584,N_33576);
or U33974 (N_33974,N_33613,N_33708);
nand U33975 (N_33975,N_33657,N_33747);
nand U33976 (N_33976,N_33678,N_33585);
xnor U33977 (N_33977,N_33608,N_33642);
nor U33978 (N_33978,N_33545,N_33711);
xnor U33979 (N_33979,N_33707,N_33641);
and U33980 (N_33980,N_33690,N_33584);
and U33981 (N_33981,N_33684,N_33638);
nand U33982 (N_33982,N_33627,N_33551);
nand U33983 (N_33983,N_33740,N_33588);
nor U33984 (N_33984,N_33653,N_33626);
nor U33985 (N_33985,N_33747,N_33656);
nor U33986 (N_33986,N_33745,N_33652);
nand U33987 (N_33987,N_33569,N_33556);
and U33988 (N_33988,N_33732,N_33626);
nand U33989 (N_33989,N_33600,N_33526);
xor U33990 (N_33990,N_33590,N_33710);
nor U33991 (N_33991,N_33543,N_33623);
and U33992 (N_33992,N_33686,N_33665);
xor U33993 (N_33993,N_33682,N_33560);
and U33994 (N_33994,N_33698,N_33531);
and U33995 (N_33995,N_33613,N_33518);
nor U33996 (N_33996,N_33594,N_33532);
xnor U33997 (N_33997,N_33697,N_33539);
nor U33998 (N_33998,N_33711,N_33522);
xnor U33999 (N_33999,N_33537,N_33550);
nand U34000 (N_34000,N_33885,N_33947);
and U34001 (N_34001,N_33793,N_33910);
nor U34002 (N_34002,N_33905,N_33961);
and U34003 (N_34003,N_33950,N_33851);
nor U34004 (N_34004,N_33797,N_33893);
and U34005 (N_34005,N_33872,N_33941);
or U34006 (N_34006,N_33946,N_33993);
and U34007 (N_34007,N_33903,N_33952);
nor U34008 (N_34008,N_33915,N_33976);
nor U34009 (N_34009,N_33897,N_33871);
nand U34010 (N_34010,N_33768,N_33996);
xnor U34011 (N_34011,N_33972,N_33942);
or U34012 (N_34012,N_33756,N_33933);
xnor U34013 (N_34013,N_33896,N_33758);
nor U34014 (N_34014,N_33939,N_33775);
nand U34015 (N_34015,N_33778,N_33819);
or U34016 (N_34016,N_33795,N_33762);
nand U34017 (N_34017,N_33830,N_33837);
nand U34018 (N_34018,N_33811,N_33997);
or U34019 (N_34019,N_33981,N_33964);
or U34020 (N_34020,N_33813,N_33943);
and U34021 (N_34021,N_33859,N_33959);
and U34022 (N_34022,N_33889,N_33789);
nor U34023 (N_34023,N_33869,N_33876);
or U34024 (N_34024,N_33785,N_33990);
xor U34025 (N_34025,N_33757,N_33936);
or U34026 (N_34026,N_33867,N_33951);
nor U34027 (N_34027,N_33878,N_33751);
nor U34028 (N_34028,N_33884,N_33843);
and U34029 (N_34029,N_33865,N_33886);
and U34030 (N_34030,N_33948,N_33974);
nor U34031 (N_34031,N_33928,N_33938);
nand U34032 (N_34032,N_33994,N_33894);
nand U34033 (N_34033,N_33999,N_33787);
xnor U34034 (N_34034,N_33855,N_33783);
nor U34035 (N_34035,N_33983,N_33820);
xor U34036 (N_34036,N_33909,N_33927);
nor U34037 (N_34037,N_33779,N_33965);
nand U34038 (N_34038,N_33922,N_33888);
xnor U34039 (N_34039,N_33831,N_33823);
xnor U34040 (N_34040,N_33991,N_33968);
xnor U34041 (N_34041,N_33854,N_33873);
and U34042 (N_34042,N_33984,N_33931);
and U34043 (N_34043,N_33792,N_33791);
nor U34044 (N_34044,N_33826,N_33962);
or U34045 (N_34045,N_33861,N_33875);
nor U34046 (N_34046,N_33838,N_33835);
and U34047 (N_34047,N_33966,N_33963);
and U34048 (N_34048,N_33945,N_33995);
nor U34049 (N_34049,N_33887,N_33839);
and U34050 (N_34050,N_33816,N_33781);
nand U34051 (N_34051,N_33923,N_33800);
nand U34052 (N_34052,N_33862,N_33752);
or U34053 (N_34053,N_33847,N_33761);
nand U34054 (N_34054,N_33763,N_33920);
xor U34055 (N_34055,N_33892,N_33804);
xnor U34056 (N_34056,N_33801,N_33987);
and U34057 (N_34057,N_33770,N_33949);
xor U34058 (N_34058,N_33908,N_33891);
or U34059 (N_34059,N_33796,N_33930);
nor U34060 (N_34060,N_33784,N_33880);
nand U34061 (N_34061,N_33988,N_33754);
nor U34062 (N_34062,N_33954,N_33812);
and U34063 (N_34063,N_33918,N_33940);
or U34064 (N_34064,N_33841,N_33767);
nand U34065 (N_34065,N_33913,N_33921);
xnor U34066 (N_34066,N_33848,N_33924);
nor U34067 (N_34067,N_33973,N_33832);
nand U34068 (N_34068,N_33919,N_33794);
or U34069 (N_34069,N_33982,N_33771);
nor U34070 (N_34070,N_33776,N_33882);
xor U34071 (N_34071,N_33824,N_33822);
or U34072 (N_34072,N_33844,N_33975);
and U34073 (N_34073,N_33805,N_33850);
or U34074 (N_34074,N_33895,N_33955);
and U34075 (N_34075,N_33842,N_33817);
and U34076 (N_34076,N_33814,N_33807);
xnor U34077 (N_34077,N_33916,N_33753);
xor U34078 (N_34078,N_33937,N_33866);
and U34079 (N_34079,N_33772,N_33932);
and U34080 (N_34080,N_33960,N_33766);
and U34081 (N_34081,N_33845,N_33840);
xnor U34082 (N_34082,N_33985,N_33857);
and U34083 (N_34083,N_33836,N_33989);
nor U34084 (N_34084,N_33904,N_33774);
and U34085 (N_34085,N_33899,N_33864);
and U34086 (N_34086,N_33907,N_33925);
and U34087 (N_34087,N_33852,N_33788);
and U34088 (N_34088,N_33992,N_33890);
and U34089 (N_34089,N_33944,N_33956);
and U34090 (N_34090,N_33760,N_33929);
xnor U34091 (N_34091,N_33858,N_33828);
or U34092 (N_34092,N_33877,N_33773);
nor U34093 (N_34093,N_33912,N_33777);
and U34094 (N_34094,N_33998,N_33970);
nand U34095 (N_34095,N_33815,N_33803);
or U34096 (N_34096,N_33802,N_33986);
nand U34097 (N_34097,N_33846,N_33977);
nor U34098 (N_34098,N_33834,N_33901);
nand U34099 (N_34099,N_33786,N_33881);
nor U34100 (N_34100,N_33825,N_33809);
or U34101 (N_34101,N_33829,N_33902);
nor U34102 (N_34102,N_33868,N_33780);
nor U34103 (N_34103,N_33958,N_33874);
nand U34104 (N_34104,N_33755,N_33906);
nor U34105 (N_34105,N_33917,N_33860);
or U34106 (N_34106,N_33863,N_33759);
and U34107 (N_34107,N_33856,N_33980);
or U34108 (N_34108,N_33782,N_33914);
xnor U34109 (N_34109,N_33979,N_33827);
and U34110 (N_34110,N_33808,N_33934);
and U34111 (N_34111,N_33799,N_33926);
xnor U34112 (N_34112,N_33969,N_33911);
nand U34113 (N_34113,N_33790,N_33870);
nand U34114 (N_34114,N_33810,N_33900);
xor U34115 (N_34115,N_33953,N_33853);
xor U34116 (N_34116,N_33764,N_33750);
nor U34117 (N_34117,N_33935,N_33765);
nor U34118 (N_34118,N_33821,N_33769);
and U34119 (N_34119,N_33818,N_33849);
and U34120 (N_34120,N_33833,N_33957);
or U34121 (N_34121,N_33978,N_33798);
or U34122 (N_34122,N_33971,N_33806);
and U34123 (N_34123,N_33967,N_33898);
nand U34124 (N_34124,N_33883,N_33879);
nor U34125 (N_34125,N_33963,N_33762);
or U34126 (N_34126,N_33871,N_33843);
nand U34127 (N_34127,N_33887,N_33992);
or U34128 (N_34128,N_33924,N_33953);
or U34129 (N_34129,N_33988,N_33869);
nor U34130 (N_34130,N_33925,N_33819);
or U34131 (N_34131,N_33829,N_33837);
or U34132 (N_34132,N_33815,N_33911);
and U34133 (N_34133,N_33933,N_33919);
nand U34134 (N_34134,N_33889,N_33974);
nand U34135 (N_34135,N_33811,N_33913);
or U34136 (N_34136,N_33924,N_33945);
or U34137 (N_34137,N_33972,N_33783);
nor U34138 (N_34138,N_33831,N_33878);
nand U34139 (N_34139,N_33760,N_33840);
or U34140 (N_34140,N_33936,N_33871);
nand U34141 (N_34141,N_33934,N_33839);
nand U34142 (N_34142,N_33932,N_33783);
and U34143 (N_34143,N_33847,N_33966);
nor U34144 (N_34144,N_33885,N_33991);
nor U34145 (N_34145,N_33785,N_33927);
nor U34146 (N_34146,N_33881,N_33771);
or U34147 (N_34147,N_33871,N_33977);
nor U34148 (N_34148,N_33904,N_33933);
or U34149 (N_34149,N_33885,N_33846);
and U34150 (N_34150,N_33765,N_33973);
nand U34151 (N_34151,N_33918,N_33770);
nor U34152 (N_34152,N_33909,N_33853);
or U34153 (N_34153,N_33843,N_33918);
nand U34154 (N_34154,N_33909,N_33922);
or U34155 (N_34155,N_33986,N_33966);
xnor U34156 (N_34156,N_33902,N_33919);
nor U34157 (N_34157,N_33995,N_33928);
or U34158 (N_34158,N_33837,N_33788);
nor U34159 (N_34159,N_33893,N_33771);
nor U34160 (N_34160,N_33757,N_33999);
or U34161 (N_34161,N_33817,N_33865);
nor U34162 (N_34162,N_33761,N_33902);
and U34163 (N_34163,N_33928,N_33994);
nand U34164 (N_34164,N_33954,N_33998);
or U34165 (N_34165,N_33904,N_33994);
nor U34166 (N_34166,N_33813,N_33918);
nor U34167 (N_34167,N_33831,N_33848);
nor U34168 (N_34168,N_33808,N_33855);
nand U34169 (N_34169,N_33981,N_33854);
or U34170 (N_34170,N_33919,N_33766);
and U34171 (N_34171,N_33833,N_33927);
xor U34172 (N_34172,N_33795,N_33806);
nor U34173 (N_34173,N_33914,N_33993);
nand U34174 (N_34174,N_33823,N_33784);
nand U34175 (N_34175,N_33930,N_33851);
or U34176 (N_34176,N_33833,N_33939);
nand U34177 (N_34177,N_33755,N_33976);
nand U34178 (N_34178,N_33970,N_33758);
xnor U34179 (N_34179,N_33909,N_33946);
or U34180 (N_34180,N_33865,N_33896);
nand U34181 (N_34181,N_33971,N_33761);
nand U34182 (N_34182,N_33836,N_33863);
xor U34183 (N_34183,N_33976,N_33767);
nor U34184 (N_34184,N_33911,N_33856);
and U34185 (N_34185,N_33909,N_33876);
or U34186 (N_34186,N_33911,N_33878);
xor U34187 (N_34187,N_33929,N_33815);
and U34188 (N_34188,N_33862,N_33813);
and U34189 (N_34189,N_33986,N_33839);
nor U34190 (N_34190,N_33993,N_33911);
or U34191 (N_34191,N_33787,N_33778);
nand U34192 (N_34192,N_33770,N_33962);
or U34193 (N_34193,N_33900,N_33990);
nand U34194 (N_34194,N_33812,N_33950);
or U34195 (N_34195,N_33811,N_33855);
nand U34196 (N_34196,N_33979,N_33869);
or U34197 (N_34197,N_33809,N_33771);
xnor U34198 (N_34198,N_33776,N_33807);
nor U34199 (N_34199,N_33927,N_33796);
nor U34200 (N_34200,N_33845,N_33991);
nor U34201 (N_34201,N_33882,N_33891);
or U34202 (N_34202,N_33751,N_33859);
or U34203 (N_34203,N_33962,N_33845);
nand U34204 (N_34204,N_33914,N_33977);
xor U34205 (N_34205,N_33920,N_33796);
xnor U34206 (N_34206,N_33888,N_33975);
nor U34207 (N_34207,N_33762,N_33950);
and U34208 (N_34208,N_33780,N_33764);
nand U34209 (N_34209,N_33779,N_33881);
nor U34210 (N_34210,N_33992,N_33826);
nand U34211 (N_34211,N_33943,N_33878);
xnor U34212 (N_34212,N_33844,N_33864);
nand U34213 (N_34213,N_33965,N_33934);
or U34214 (N_34214,N_33763,N_33765);
nor U34215 (N_34215,N_33768,N_33904);
or U34216 (N_34216,N_33904,N_33839);
nand U34217 (N_34217,N_33804,N_33988);
nor U34218 (N_34218,N_33887,N_33924);
or U34219 (N_34219,N_33888,N_33914);
and U34220 (N_34220,N_33837,N_33859);
xnor U34221 (N_34221,N_33903,N_33752);
nor U34222 (N_34222,N_33756,N_33856);
nand U34223 (N_34223,N_33819,N_33971);
xnor U34224 (N_34224,N_33850,N_33969);
or U34225 (N_34225,N_33792,N_33947);
nand U34226 (N_34226,N_33802,N_33893);
nor U34227 (N_34227,N_33814,N_33946);
or U34228 (N_34228,N_33996,N_33867);
nor U34229 (N_34229,N_33861,N_33920);
nand U34230 (N_34230,N_33856,N_33951);
nand U34231 (N_34231,N_33951,N_33754);
xnor U34232 (N_34232,N_33906,N_33878);
or U34233 (N_34233,N_33789,N_33953);
or U34234 (N_34234,N_33750,N_33755);
nand U34235 (N_34235,N_33983,N_33811);
nor U34236 (N_34236,N_33787,N_33803);
nor U34237 (N_34237,N_33814,N_33779);
xnor U34238 (N_34238,N_33930,N_33951);
xor U34239 (N_34239,N_33794,N_33895);
or U34240 (N_34240,N_33819,N_33986);
nand U34241 (N_34241,N_33807,N_33996);
and U34242 (N_34242,N_33848,N_33965);
xor U34243 (N_34243,N_33888,N_33986);
or U34244 (N_34244,N_33972,N_33820);
and U34245 (N_34245,N_33900,N_33966);
xnor U34246 (N_34246,N_33911,N_33895);
xor U34247 (N_34247,N_33995,N_33895);
or U34248 (N_34248,N_33835,N_33849);
nor U34249 (N_34249,N_33795,N_33791);
and U34250 (N_34250,N_34010,N_34008);
nor U34251 (N_34251,N_34240,N_34223);
xnor U34252 (N_34252,N_34235,N_34085);
nor U34253 (N_34253,N_34215,N_34179);
nor U34254 (N_34254,N_34197,N_34149);
xnor U34255 (N_34255,N_34170,N_34156);
and U34256 (N_34256,N_34023,N_34222);
nor U34257 (N_34257,N_34234,N_34244);
and U34258 (N_34258,N_34020,N_34238);
and U34259 (N_34259,N_34060,N_34136);
or U34260 (N_34260,N_34206,N_34157);
nor U34261 (N_34261,N_34131,N_34117);
or U34262 (N_34262,N_34114,N_34226);
or U34263 (N_34263,N_34013,N_34087);
or U34264 (N_34264,N_34014,N_34181);
nand U34265 (N_34265,N_34221,N_34064);
nand U34266 (N_34266,N_34196,N_34052);
xor U34267 (N_34267,N_34134,N_34062);
or U34268 (N_34268,N_34152,N_34193);
nand U34269 (N_34269,N_34092,N_34048);
or U34270 (N_34270,N_34161,N_34009);
nor U34271 (N_34271,N_34146,N_34081);
or U34272 (N_34272,N_34204,N_34115);
and U34273 (N_34273,N_34214,N_34249);
or U34274 (N_34274,N_34162,N_34203);
xor U34275 (N_34275,N_34164,N_34248);
nor U34276 (N_34276,N_34137,N_34056);
xnor U34277 (N_34277,N_34088,N_34151);
nor U34278 (N_34278,N_34100,N_34180);
nand U34279 (N_34279,N_34074,N_34175);
nor U34280 (N_34280,N_34024,N_34033);
and U34281 (N_34281,N_34150,N_34201);
and U34282 (N_34282,N_34055,N_34118);
xor U34283 (N_34283,N_34194,N_34192);
and U34284 (N_34284,N_34028,N_34002);
xnor U34285 (N_34285,N_34163,N_34091);
nor U34286 (N_34286,N_34111,N_34158);
nand U34287 (N_34287,N_34126,N_34046);
nand U34288 (N_34288,N_34065,N_34069);
nor U34289 (N_34289,N_34217,N_34070);
nand U34290 (N_34290,N_34123,N_34075);
xnor U34291 (N_34291,N_34246,N_34095);
nor U34292 (N_34292,N_34236,N_34188);
nand U34293 (N_34293,N_34026,N_34172);
nor U34294 (N_34294,N_34237,N_34077);
and U34295 (N_34295,N_34232,N_34102);
and U34296 (N_34296,N_34053,N_34001);
nand U34297 (N_34297,N_34079,N_34177);
nand U34298 (N_34298,N_34015,N_34144);
nand U34299 (N_34299,N_34208,N_34145);
nor U34300 (N_34300,N_34120,N_34159);
xor U34301 (N_34301,N_34034,N_34030);
nand U34302 (N_34302,N_34209,N_34242);
xor U34303 (N_34303,N_34017,N_34216);
or U34304 (N_34304,N_34182,N_34012);
and U34305 (N_34305,N_34160,N_34220);
and U34306 (N_34306,N_34132,N_34143);
and U34307 (N_34307,N_34076,N_34141);
nand U34308 (N_34308,N_34099,N_34186);
and U34309 (N_34309,N_34029,N_34166);
and U34310 (N_34310,N_34059,N_34154);
nand U34311 (N_34311,N_34039,N_34219);
and U34312 (N_34312,N_34178,N_34116);
nand U34313 (N_34313,N_34190,N_34218);
or U34314 (N_34314,N_34006,N_34243);
nand U34315 (N_34315,N_34082,N_34142);
and U34316 (N_34316,N_34155,N_34121);
and U34317 (N_34317,N_34038,N_34113);
nor U34318 (N_34318,N_34035,N_34213);
or U34319 (N_34319,N_34231,N_34239);
or U34320 (N_34320,N_34057,N_34071);
xor U34321 (N_34321,N_34090,N_34225);
and U34322 (N_34322,N_34040,N_34054);
nor U34323 (N_34323,N_34000,N_34176);
or U34324 (N_34324,N_34049,N_34110);
nor U34325 (N_34325,N_34067,N_34138);
nand U34326 (N_34326,N_34021,N_34096);
or U34327 (N_34327,N_34078,N_34011);
nor U34328 (N_34328,N_34227,N_34198);
and U34329 (N_34329,N_34127,N_34068);
nand U34330 (N_34330,N_34041,N_34018);
xor U34331 (N_34331,N_34016,N_34129);
and U34332 (N_34332,N_34037,N_34004);
xnor U34333 (N_34333,N_34022,N_34247);
xor U34334 (N_34334,N_34089,N_34173);
nand U34335 (N_34335,N_34169,N_34093);
nand U34336 (N_34336,N_34147,N_34139);
nor U34337 (N_34337,N_34027,N_34171);
nand U34338 (N_34338,N_34105,N_34047);
and U34339 (N_34339,N_34122,N_34094);
nand U34340 (N_34340,N_34135,N_34224);
nor U34341 (N_34341,N_34083,N_34212);
nand U34342 (N_34342,N_34107,N_34073);
nor U34343 (N_34343,N_34195,N_34205);
nor U34344 (N_34344,N_34211,N_34032);
nor U34345 (N_34345,N_34167,N_34112);
and U34346 (N_34346,N_34228,N_34125);
nand U34347 (N_34347,N_34187,N_34168);
xnor U34348 (N_34348,N_34066,N_34080);
nand U34349 (N_34349,N_34229,N_34063);
nand U34350 (N_34350,N_34050,N_34005);
or U34351 (N_34351,N_34109,N_34084);
xnor U34352 (N_34352,N_34153,N_34140);
nor U34353 (N_34353,N_34148,N_34207);
nand U34354 (N_34354,N_34210,N_34106);
nor U34355 (N_34355,N_34174,N_34241);
or U34356 (N_34356,N_34101,N_34184);
nor U34357 (N_34357,N_34199,N_34007);
and U34358 (N_34358,N_34031,N_34130);
or U34359 (N_34359,N_34097,N_34108);
nand U34360 (N_34360,N_34124,N_34104);
and U34361 (N_34361,N_34183,N_34043);
nand U34362 (N_34362,N_34128,N_34191);
nand U34363 (N_34363,N_34098,N_34086);
or U34364 (N_34364,N_34072,N_34185);
xor U34365 (N_34365,N_34103,N_34045);
or U34366 (N_34366,N_34061,N_34230);
or U34367 (N_34367,N_34119,N_34133);
nand U34368 (N_34368,N_34025,N_34044);
xor U34369 (N_34369,N_34058,N_34042);
nand U34370 (N_34370,N_34189,N_34051);
or U34371 (N_34371,N_34202,N_34003);
nor U34372 (N_34372,N_34019,N_34245);
nor U34373 (N_34373,N_34200,N_34233);
and U34374 (N_34374,N_34036,N_34165);
xor U34375 (N_34375,N_34074,N_34037);
and U34376 (N_34376,N_34078,N_34244);
nor U34377 (N_34377,N_34128,N_34190);
xnor U34378 (N_34378,N_34225,N_34146);
and U34379 (N_34379,N_34132,N_34202);
and U34380 (N_34380,N_34076,N_34085);
xor U34381 (N_34381,N_34147,N_34176);
and U34382 (N_34382,N_34003,N_34151);
nand U34383 (N_34383,N_34157,N_34118);
or U34384 (N_34384,N_34238,N_34099);
or U34385 (N_34385,N_34093,N_34020);
and U34386 (N_34386,N_34187,N_34174);
and U34387 (N_34387,N_34191,N_34029);
or U34388 (N_34388,N_34145,N_34027);
and U34389 (N_34389,N_34151,N_34039);
nor U34390 (N_34390,N_34033,N_34175);
nor U34391 (N_34391,N_34220,N_34129);
xnor U34392 (N_34392,N_34055,N_34029);
nand U34393 (N_34393,N_34168,N_34058);
xor U34394 (N_34394,N_34161,N_34003);
and U34395 (N_34395,N_34081,N_34214);
nand U34396 (N_34396,N_34035,N_34079);
xnor U34397 (N_34397,N_34091,N_34189);
xnor U34398 (N_34398,N_34191,N_34200);
and U34399 (N_34399,N_34093,N_34146);
or U34400 (N_34400,N_34050,N_34169);
nor U34401 (N_34401,N_34066,N_34174);
xor U34402 (N_34402,N_34124,N_34037);
nand U34403 (N_34403,N_34211,N_34241);
nor U34404 (N_34404,N_34009,N_34038);
and U34405 (N_34405,N_34136,N_34096);
and U34406 (N_34406,N_34225,N_34205);
xnor U34407 (N_34407,N_34078,N_34115);
or U34408 (N_34408,N_34223,N_34169);
nor U34409 (N_34409,N_34039,N_34150);
or U34410 (N_34410,N_34087,N_34232);
nand U34411 (N_34411,N_34245,N_34054);
nor U34412 (N_34412,N_34203,N_34220);
nor U34413 (N_34413,N_34219,N_34087);
and U34414 (N_34414,N_34067,N_34109);
and U34415 (N_34415,N_34085,N_34079);
nor U34416 (N_34416,N_34069,N_34117);
xnor U34417 (N_34417,N_34099,N_34219);
xor U34418 (N_34418,N_34054,N_34194);
and U34419 (N_34419,N_34064,N_34020);
nor U34420 (N_34420,N_34143,N_34016);
xor U34421 (N_34421,N_34009,N_34116);
and U34422 (N_34422,N_34050,N_34012);
or U34423 (N_34423,N_34121,N_34244);
nor U34424 (N_34424,N_34110,N_34018);
or U34425 (N_34425,N_34227,N_34142);
nand U34426 (N_34426,N_34024,N_34018);
or U34427 (N_34427,N_34218,N_34242);
or U34428 (N_34428,N_34216,N_34038);
or U34429 (N_34429,N_34087,N_34032);
nand U34430 (N_34430,N_34166,N_34184);
or U34431 (N_34431,N_34067,N_34205);
and U34432 (N_34432,N_34120,N_34246);
xor U34433 (N_34433,N_34225,N_34101);
nand U34434 (N_34434,N_34231,N_34086);
xnor U34435 (N_34435,N_34239,N_34176);
or U34436 (N_34436,N_34218,N_34163);
xor U34437 (N_34437,N_34121,N_34011);
and U34438 (N_34438,N_34203,N_34085);
nand U34439 (N_34439,N_34106,N_34176);
xnor U34440 (N_34440,N_34067,N_34092);
xnor U34441 (N_34441,N_34187,N_34061);
xnor U34442 (N_34442,N_34195,N_34210);
nor U34443 (N_34443,N_34170,N_34063);
nor U34444 (N_34444,N_34094,N_34035);
and U34445 (N_34445,N_34076,N_34075);
nand U34446 (N_34446,N_34240,N_34145);
xnor U34447 (N_34447,N_34093,N_34085);
or U34448 (N_34448,N_34110,N_34094);
xor U34449 (N_34449,N_34110,N_34115);
nor U34450 (N_34450,N_34183,N_34062);
and U34451 (N_34451,N_34248,N_34065);
xnor U34452 (N_34452,N_34208,N_34081);
nor U34453 (N_34453,N_34149,N_34218);
nor U34454 (N_34454,N_34116,N_34099);
and U34455 (N_34455,N_34020,N_34128);
nor U34456 (N_34456,N_34155,N_34097);
and U34457 (N_34457,N_34107,N_34134);
or U34458 (N_34458,N_34198,N_34079);
and U34459 (N_34459,N_34034,N_34193);
nand U34460 (N_34460,N_34131,N_34228);
or U34461 (N_34461,N_34115,N_34215);
or U34462 (N_34462,N_34103,N_34204);
or U34463 (N_34463,N_34121,N_34031);
xor U34464 (N_34464,N_34123,N_34222);
and U34465 (N_34465,N_34120,N_34183);
nand U34466 (N_34466,N_34020,N_34108);
and U34467 (N_34467,N_34035,N_34117);
and U34468 (N_34468,N_34185,N_34008);
or U34469 (N_34469,N_34240,N_34135);
or U34470 (N_34470,N_34204,N_34022);
or U34471 (N_34471,N_34143,N_34207);
and U34472 (N_34472,N_34188,N_34084);
nand U34473 (N_34473,N_34177,N_34018);
nor U34474 (N_34474,N_34170,N_34167);
and U34475 (N_34475,N_34036,N_34199);
xnor U34476 (N_34476,N_34176,N_34083);
xor U34477 (N_34477,N_34115,N_34131);
nand U34478 (N_34478,N_34187,N_34190);
xor U34479 (N_34479,N_34173,N_34032);
nor U34480 (N_34480,N_34068,N_34197);
xnor U34481 (N_34481,N_34238,N_34211);
xnor U34482 (N_34482,N_34135,N_34033);
xnor U34483 (N_34483,N_34208,N_34200);
xor U34484 (N_34484,N_34086,N_34090);
or U34485 (N_34485,N_34040,N_34065);
xnor U34486 (N_34486,N_34043,N_34106);
nand U34487 (N_34487,N_34152,N_34065);
nor U34488 (N_34488,N_34065,N_34014);
xnor U34489 (N_34489,N_34122,N_34172);
or U34490 (N_34490,N_34086,N_34004);
nor U34491 (N_34491,N_34233,N_34145);
xnor U34492 (N_34492,N_34230,N_34129);
or U34493 (N_34493,N_34197,N_34235);
nor U34494 (N_34494,N_34196,N_34096);
xnor U34495 (N_34495,N_34153,N_34016);
xnor U34496 (N_34496,N_34219,N_34092);
or U34497 (N_34497,N_34013,N_34171);
xor U34498 (N_34498,N_34198,N_34056);
xnor U34499 (N_34499,N_34189,N_34231);
xnor U34500 (N_34500,N_34323,N_34493);
or U34501 (N_34501,N_34440,N_34257);
nand U34502 (N_34502,N_34260,N_34492);
or U34503 (N_34503,N_34471,N_34488);
or U34504 (N_34504,N_34322,N_34464);
xor U34505 (N_34505,N_34457,N_34458);
nor U34506 (N_34506,N_34359,N_34268);
nand U34507 (N_34507,N_34409,N_34309);
nand U34508 (N_34508,N_34274,N_34305);
or U34509 (N_34509,N_34265,N_34293);
nor U34510 (N_34510,N_34276,N_34413);
nor U34511 (N_34511,N_34315,N_34391);
and U34512 (N_34512,N_34427,N_34474);
nand U34513 (N_34513,N_34347,N_34373);
nand U34514 (N_34514,N_34299,N_34314);
and U34515 (N_34515,N_34449,N_34330);
and U34516 (N_34516,N_34366,N_34402);
and U34517 (N_34517,N_34415,N_34496);
or U34518 (N_34518,N_34311,N_34335);
xor U34519 (N_34519,N_34331,N_34460);
or U34520 (N_34520,N_34376,N_34439);
and U34521 (N_34521,N_34490,N_34332);
or U34522 (N_34522,N_34364,N_34499);
xnor U34523 (N_34523,N_34404,N_34400);
or U34524 (N_34524,N_34381,N_34319);
nor U34525 (N_34525,N_34423,N_34281);
nand U34526 (N_34526,N_34301,N_34452);
xnor U34527 (N_34527,N_34431,N_34422);
and U34528 (N_34528,N_34416,N_34395);
nand U34529 (N_34529,N_34481,N_34307);
xnor U34530 (N_34530,N_34258,N_34454);
nand U34531 (N_34531,N_34434,N_34362);
nand U34532 (N_34532,N_34387,N_34450);
xnor U34533 (N_34533,N_34393,N_34351);
nor U34534 (N_34534,N_34370,N_34252);
and U34535 (N_34535,N_34345,N_34382);
or U34536 (N_34536,N_34304,N_34285);
nor U34537 (N_34537,N_34491,N_34321);
and U34538 (N_34538,N_34463,N_34336);
nor U34539 (N_34539,N_34384,N_34302);
xnor U34540 (N_34540,N_34346,N_34455);
and U34541 (N_34541,N_34385,N_34442);
nand U34542 (N_34542,N_34446,N_34377);
and U34543 (N_34543,N_34353,N_34424);
xnor U34544 (N_34544,N_34448,N_34406);
xnor U34545 (N_34545,N_34361,N_34340);
xor U34546 (N_34546,N_34255,N_34467);
or U34547 (N_34547,N_34479,N_34392);
or U34548 (N_34548,N_34296,N_34365);
or U34549 (N_34549,N_34256,N_34269);
or U34550 (N_34550,N_34349,N_34473);
nand U34551 (N_34551,N_34444,N_34478);
nor U34552 (N_34552,N_34254,N_34287);
and U34553 (N_34553,N_34432,N_34277);
xor U34554 (N_34554,N_34379,N_34356);
xnor U34555 (N_34555,N_34263,N_34344);
and U34556 (N_34556,N_34380,N_34426);
or U34557 (N_34557,N_34408,N_34435);
nand U34558 (N_34558,N_34411,N_34262);
nor U34559 (N_34559,N_34494,N_34280);
nor U34560 (N_34560,N_34447,N_34477);
nand U34561 (N_34561,N_34306,N_34297);
nand U34562 (N_34562,N_34367,N_34484);
xnor U34563 (N_34563,N_34325,N_34355);
xor U34564 (N_34564,N_34456,N_34267);
or U34565 (N_34565,N_34453,N_34389);
or U34566 (N_34566,N_34418,N_34261);
xnor U34567 (N_34567,N_34390,N_34412);
xnor U34568 (N_34568,N_34295,N_34253);
nand U34569 (N_34569,N_34480,N_34405);
xor U34570 (N_34570,N_34337,N_34282);
nand U34571 (N_34571,N_34470,N_34300);
or U34572 (N_34572,N_34468,N_34371);
and U34573 (N_34573,N_34425,N_34388);
xnor U34574 (N_34574,N_34270,N_34279);
and U34575 (N_34575,N_34328,N_34310);
or U34576 (N_34576,N_34386,N_34437);
nor U34577 (N_34577,N_34461,N_34273);
nor U34578 (N_34578,N_34383,N_34317);
nor U34579 (N_34579,N_34368,N_34286);
and U34580 (N_34580,N_34363,N_34443);
or U34581 (N_34581,N_34329,N_34324);
and U34582 (N_34582,N_34466,N_34436);
or U34583 (N_34583,N_34401,N_34275);
and U34584 (N_34584,N_34266,N_34469);
nor U34585 (N_34585,N_34414,N_34482);
nand U34586 (N_34586,N_34360,N_34459);
or U34587 (N_34587,N_34420,N_34397);
nand U34588 (N_34588,N_34294,N_34292);
and U34589 (N_34589,N_34271,N_34372);
nand U34590 (N_34590,N_34326,N_34399);
nor U34591 (N_34591,N_34486,N_34250);
or U34592 (N_34592,N_34462,N_34378);
and U34593 (N_34593,N_34288,N_34289);
and U34594 (N_34594,N_34465,N_34433);
or U34595 (N_34595,N_34375,N_34483);
xnor U34596 (N_34596,N_34369,N_34316);
and U34597 (N_34597,N_34357,N_34343);
xor U34598 (N_34598,N_34290,N_34298);
and U34599 (N_34599,N_34394,N_34497);
nand U34600 (N_34600,N_34251,N_34445);
or U34601 (N_34601,N_34358,N_34374);
xnor U34602 (N_34602,N_34348,N_34264);
nor U34603 (N_34603,N_34352,N_34350);
xnor U34604 (N_34604,N_34398,N_34312);
and U34605 (N_34605,N_34313,N_34338);
xor U34606 (N_34606,N_34354,N_34272);
and U34607 (N_34607,N_34334,N_34421);
xor U34608 (N_34608,N_34438,N_34489);
or U34609 (N_34609,N_34333,N_34419);
xor U34610 (N_34610,N_34320,N_34339);
or U34611 (N_34611,N_34428,N_34430);
nor U34612 (N_34612,N_34417,N_34476);
nor U34613 (N_34613,N_34303,N_34403);
and U34614 (N_34614,N_34407,N_34410);
or U34615 (N_34615,N_34308,N_34485);
nor U34616 (N_34616,N_34429,N_34318);
nand U34617 (N_34617,N_34284,N_34472);
or U34618 (N_34618,N_34259,N_34475);
and U34619 (N_34619,N_34342,N_34451);
or U34620 (N_34620,N_34396,N_34341);
and U34621 (N_34621,N_34498,N_34327);
nand U34622 (N_34622,N_34283,N_34278);
and U34623 (N_34623,N_34441,N_34487);
nor U34624 (N_34624,N_34291,N_34495);
xor U34625 (N_34625,N_34432,N_34460);
nand U34626 (N_34626,N_34283,N_34382);
nor U34627 (N_34627,N_34323,N_34385);
nand U34628 (N_34628,N_34306,N_34290);
xor U34629 (N_34629,N_34403,N_34390);
and U34630 (N_34630,N_34313,N_34296);
xnor U34631 (N_34631,N_34301,N_34328);
nand U34632 (N_34632,N_34344,N_34341);
nand U34633 (N_34633,N_34389,N_34464);
nor U34634 (N_34634,N_34422,N_34457);
or U34635 (N_34635,N_34404,N_34331);
xor U34636 (N_34636,N_34422,N_34479);
or U34637 (N_34637,N_34318,N_34464);
nand U34638 (N_34638,N_34499,N_34405);
or U34639 (N_34639,N_34401,N_34288);
nor U34640 (N_34640,N_34273,N_34351);
nand U34641 (N_34641,N_34258,N_34307);
nor U34642 (N_34642,N_34375,N_34379);
and U34643 (N_34643,N_34408,N_34386);
and U34644 (N_34644,N_34355,N_34466);
and U34645 (N_34645,N_34288,N_34430);
nand U34646 (N_34646,N_34442,N_34286);
xor U34647 (N_34647,N_34490,N_34322);
xor U34648 (N_34648,N_34395,N_34373);
xor U34649 (N_34649,N_34461,N_34276);
xnor U34650 (N_34650,N_34483,N_34303);
nor U34651 (N_34651,N_34421,N_34332);
and U34652 (N_34652,N_34313,N_34280);
or U34653 (N_34653,N_34297,N_34337);
and U34654 (N_34654,N_34340,N_34278);
nand U34655 (N_34655,N_34499,N_34472);
nor U34656 (N_34656,N_34365,N_34418);
nor U34657 (N_34657,N_34425,N_34407);
or U34658 (N_34658,N_34476,N_34390);
xnor U34659 (N_34659,N_34298,N_34338);
xnor U34660 (N_34660,N_34366,N_34293);
nor U34661 (N_34661,N_34350,N_34292);
nor U34662 (N_34662,N_34312,N_34373);
nor U34663 (N_34663,N_34299,N_34440);
nor U34664 (N_34664,N_34256,N_34359);
xor U34665 (N_34665,N_34494,N_34435);
nand U34666 (N_34666,N_34296,N_34487);
xnor U34667 (N_34667,N_34457,N_34328);
nor U34668 (N_34668,N_34383,N_34453);
xnor U34669 (N_34669,N_34328,N_34492);
or U34670 (N_34670,N_34284,N_34298);
nand U34671 (N_34671,N_34319,N_34320);
and U34672 (N_34672,N_34388,N_34343);
nor U34673 (N_34673,N_34411,N_34474);
or U34674 (N_34674,N_34485,N_34379);
nand U34675 (N_34675,N_34255,N_34471);
xnor U34676 (N_34676,N_34361,N_34419);
nand U34677 (N_34677,N_34301,N_34499);
or U34678 (N_34678,N_34358,N_34407);
nor U34679 (N_34679,N_34459,N_34478);
and U34680 (N_34680,N_34295,N_34301);
xor U34681 (N_34681,N_34262,N_34320);
nor U34682 (N_34682,N_34295,N_34370);
and U34683 (N_34683,N_34300,N_34285);
nand U34684 (N_34684,N_34428,N_34443);
nor U34685 (N_34685,N_34351,N_34319);
xnor U34686 (N_34686,N_34410,N_34326);
nor U34687 (N_34687,N_34364,N_34383);
nor U34688 (N_34688,N_34293,N_34469);
nand U34689 (N_34689,N_34316,N_34364);
and U34690 (N_34690,N_34458,N_34290);
and U34691 (N_34691,N_34259,N_34402);
nor U34692 (N_34692,N_34258,N_34373);
or U34693 (N_34693,N_34433,N_34325);
nor U34694 (N_34694,N_34260,N_34494);
nor U34695 (N_34695,N_34408,N_34402);
or U34696 (N_34696,N_34366,N_34438);
nor U34697 (N_34697,N_34302,N_34343);
and U34698 (N_34698,N_34400,N_34475);
nor U34699 (N_34699,N_34471,N_34271);
xor U34700 (N_34700,N_34402,N_34367);
or U34701 (N_34701,N_34492,N_34372);
xor U34702 (N_34702,N_34386,N_34379);
and U34703 (N_34703,N_34481,N_34418);
and U34704 (N_34704,N_34437,N_34435);
xor U34705 (N_34705,N_34297,N_34296);
or U34706 (N_34706,N_34443,N_34468);
and U34707 (N_34707,N_34380,N_34444);
or U34708 (N_34708,N_34373,N_34396);
nand U34709 (N_34709,N_34282,N_34490);
or U34710 (N_34710,N_34307,N_34253);
xor U34711 (N_34711,N_34337,N_34338);
and U34712 (N_34712,N_34465,N_34261);
nand U34713 (N_34713,N_34326,N_34408);
nor U34714 (N_34714,N_34491,N_34389);
and U34715 (N_34715,N_34481,N_34431);
nor U34716 (N_34716,N_34475,N_34495);
or U34717 (N_34717,N_34321,N_34419);
nand U34718 (N_34718,N_34382,N_34449);
nand U34719 (N_34719,N_34341,N_34285);
nor U34720 (N_34720,N_34447,N_34320);
nor U34721 (N_34721,N_34371,N_34288);
or U34722 (N_34722,N_34373,N_34394);
xor U34723 (N_34723,N_34400,N_34280);
nand U34724 (N_34724,N_34494,N_34281);
xnor U34725 (N_34725,N_34366,N_34364);
and U34726 (N_34726,N_34378,N_34465);
or U34727 (N_34727,N_34378,N_34289);
nand U34728 (N_34728,N_34392,N_34494);
xor U34729 (N_34729,N_34298,N_34273);
or U34730 (N_34730,N_34253,N_34268);
nor U34731 (N_34731,N_34376,N_34313);
nor U34732 (N_34732,N_34296,N_34489);
xor U34733 (N_34733,N_34266,N_34335);
and U34734 (N_34734,N_34435,N_34483);
nor U34735 (N_34735,N_34431,N_34425);
nor U34736 (N_34736,N_34471,N_34328);
or U34737 (N_34737,N_34288,N_34343);
nand U34738 (N_34738,N_34373,N_34433);
and U34739 (N_34739,N_34471,N_34406);
and U34740 (N_34740,N_34268,N_34412);
nor U34741 (N_34741,N_34484,N_34473);
xnor U34742 (N_34742,N_34296,N_34295);
nand U34743 (N_34743,N_34290,N_34487);
nand U34744 (N_34744,N_34339,N_34261);
nand U34745 (N_34745,N_34441,N_34417);
xor U34746 (N_34746,N_34455,N_34369);
or U34747 (N_34747,N_34315,N_34380);
nor U34748 (N_34748,N_34284,N_34461);
nor U34749 (N_34749,N_34453,N_34385);
or U34750 (N_34750,N_34619,N_34520);
or U34751 (N_34751,N_34576,N_34706);
nor U34752 (N_34752,N_34655,N_34545);
nand U34753 (N_34753,N_34530,N_34737);
nor U34754 (N_34754,N_34584,N_34531);
and U34755 (N_34755,N_34620,N_34721);
or U34756 (N_34756,N_34521,N_34507);
or U34757 (N_34757,N_34656,N_34672);
and U34758 (N_34758,N_34708,N_34549);
nor U34759 (N_34759,N_34550,N_34733);
or U34760 (N_34760,N_34742,N_34730);
nor U34761 (N_34761,N_34664,N_34609);
nand U34762 (N_34762,N_34562,N_34718);
xor U34763 (N_34763,N_34692,N_34564);
and U34764 (N_34764,N_34675,N_34616);
nor U34765 (N_34765,N_34647,N_34663);
and U34766 (N_34766,N_34502,N_34665);
and U34767 (N_34767,N_34657,N_34695);
nor U34768 (N_34768,N_34691,N_34652);
or U34769 (N_34769,N_34518,N_34589);
xor U34770 (N_34770,N_34610,N_34709);
nor U34771 (N_34771,N_34746,N_34575);
and U34772 (N_34772,N_34683,N_34707);
or U34773 (N_34773,N_34661,N_34579);
nand U34774 (N_34774,N_34682,N_34563);
nand U34775 (N_34775,N_34537,N_34541);
nand U34776 (N_34776,N_34642,N_34741);
and U34777 (N_34777,N_34714,N_34535);
and U34778 (N_34778,N_34527,N_34641);
or U34779 (N_34779,N_34681,N_34582);
nand U34780 (N_34780,N_34660,N_34572);
nor U34781 (N_34781,N_34595,N_34585);
or U34782 (N_34782,N_34633,N_34534);
xor U34783 (N_34783,N_34732,N_34643);
or U34784 (N_34784,N_34587,N_34583);
nand U34785 (N_34785,N_34649,N_34634);
xnor U34786 (N_34786,N_34560,N_34561);
nand U34787 (N_34787,N_34710,N_34543);
nand U34788 (N_34788,N_34739,N_34601);
xor U34789 (N_34789,N_34577,N_34745);
nand U34790 (N_34790,N_34627,N_34640);
xor U34791 (N_34791,N_34626,N_34608);
and U34792 (N_34792,N_34523,N_34712);
nor U34793 (N_34793,N_34611,N_34635);
and U34794 (N_34794,N_34567,N_34510);
or U34795 (N_34795,N_34592,N_34728);
and U34796 (N_34796,N_34598,N_34696);
nand U34797 (N_34797,N_34738,N_34632);
or U34798 (N_34798,N_34704,N_34559);
and U34799 (N_34799,N_34613,N_34514);
nand U34800 (N_34800,N_34676,N_34720);
or U34801 (N_34801,N_34740,N_34658);
nor U34802 (N_34802,N_34662,N_34565);
xor U34803 (N_34803,N_34574,N_34668);
xnor U34804 (N_34804,N_34586,N_34693);
and U34805 (N_34805,N_34505,N_34606);
or U34806 (N_34806,N_34501,N_34529);
and U34807 (N_34807,N_34503,N_34686);
nor U34808 (N_34808,N_34628,N_34729);
and U34809 (N_34809,N_34605,N_34622);
xor U34810 (N_34810,N_34717,N_34525);
or U34811 (N_34811,N_34556,N_34536);
or U34812 (N_34812,N_34636,N_34517);
nand U34813 (N_34813,N_34684,N_34645);
xnor U34814 (N_34814,N_34734,N_34558);
xnor U34815 (N_34815,N_34749,N_34604);
nor U34816 (N_34816,N_34674,N_34509);
nor U34817 (N_34817,N_34702,N_34697);
xor U34818 (N_34818,N_34571,N_34594);
xnor U34819 (N_34819,N_34719,N_34698);
nor U34820 (N_34820,N_34731,N_34651);
nand U34821 (N_34821,N_34617,N_34666);
xnor U34822 (N_34822,N_34580,N_34516);
nand U34823 (N_34823,N_34679,N_34726);
or U34824 (N_34824,N_34654,N_34519);
and U34825 (N_34825,N_34639,N_34504);
or U34826 (N_34826,N_34694,N_34716);
xnor U34827 (N_34827,N_34670,N_34569);
xor U34828 (N_34828,N_34555,N_34687);
or U34829 (N_34829,N_34568,N_34690);
and U34830 (N_34830,N_34588,N_34596);
and U34831 (N_34831,N_34538,N_34593);
nor U34832 (N_34832,N_34603,N_34500);
or U34833 (N_34833,N_34624,N_34623);
or U34834 (N_34834,N_34557,N_34607);
nand U34835 (N_34835,N_34680,N_34621);
or U34836 (N_34836,N_34602,N_34650);
nand U34837 (N_34837,N_34638,N_34630);
and U34838 (N_34838,N_34700,N_34506);
nor U34839 (N_34839,N_34548,N_34673);
or U34840 (N_34840,N_34713,N_34533);
nor U34841 (N_34841,N_34615,N_34573);
nor U34842 (N_34842,N_34748,N_34532);
xnor U34843 (N_34843,N_34711,N_34590);
and U34844 (N_34844,N_34612,N_34540);
and U34845 (N_34845,N_34625,N_34512);
xor U34846 (N_34846,N_34648,N_34667);
xnor U34847 (N_34847,N_34554,N_34581);
nand U34848 (N_34848,N_34566,N_34547);
and U34849 (N_34849,N_34677,N_34699);
or U34850 (N_34850,N_34522,N_34618);
xor U34851 (N_34851,N_34544,N_34553);
nor U34852 (N_34852,N_34744,N_34526);
or U34853 (N_34853,N_34600,N_34685);
or U34854 (N_34854,N_34552,N_34546);
nor U34855 (N_34855,N_34715,N_34542);
or U34856 (N_34856,N_34644,N_34743);
nand U34857 (N_34857,N_34727,N_34678);
or U34858 (N_34858,N_34513,N_34578);
nor U34859 (N_34859,N_34637,N_34591);
and U34860 (N_34860,N_34597,N_34671);
nand U34861 (N_34861,N_34599,N_34669);
and U34862 (N_34862,N_34735,N_34508);
nor U34863 (N_34863,N_34689,N_34570);
xor U34864 (N_34864,N_34722,N_34703);
nor U34865 (N_34865,N_34701,N_34515);
xnor U34866 (N_34866,N_34551,N_34688);
nor U34867 (N_34867,N_34736,N_34725);
nor U34868 (N_34868,N_34511,N_34528);
and U34869 (N_34869,N_34653,N_34659);
xor U34870 (N_34870,N_34524,N_34631);
or U34871 (N_34871,N_34723,N_34629);
nor U34872 (N_34872,N_34705,N_34646);
nand U34873 (N_34873,N_34539,N_34614);
xnor U34874 (N_34874,N_34747,N_34724);
or U34875 (N_34875,N_34596,N_34720);
nand U34876 (N_34876,N_34504,N_34701);
and U34877 (N_34877,N_34692,N_34684);
nor U34878 (N_34878,N_34644,N_34583);
or U34879 (N_34879,N_34559,N_34650);
and U34880 (N_34880,N_34610,N_34663);
xnor U34881 (N_34881,N_34707,N_34571);
and U34882 (N_34882,N_34650,N_34510);
nand U34883 (N_34883,N_34576,N_34680);
xor U34884 (N_34884,N_34719,N_34654);
xor U34885 (N_34885,N_34714,N_34626);
nor U34886 (N_34886,N_34571,N_34744);
nor U34887 (N_34887,N_34509,N_34691);
or U34888 (N_34888,N_34712,N_34681);
xnor U34889 (N_34889,N_34747,N_34516);
nor U34890 (N_34890,N_34630,N_34610);
nand U34891 (N_34891,N_34717,N_34673);
xor U34892 (N_34892,N_34562,N_34535);
and U34893 (N_34893,N_34730,N_34523);
nor U34894 (N_34894,N_34592,N_34642);
or U34895 (N_34895,N_34579,N_34616);
xnor U34896 (N_34896,N_34665,N_34707);
or U34897 (N_34897,N_34548,N_34647);
or U34898 (N_34898,N_34549,N_34704);
and U34899 (N_34899,N_34663,N_34565);
and U34900 (N_34900,N_34659,N_34740);
nor U34901 (N_34901,N_34540,N_34614);
nor U34902 (N_34902,N_34677,N_34604);
nor U34903 (N_34903,N_34604,N_34603);
nand U34904 (N_34904,N_34641,N_34739);
and U34905 (N_34905,N_34718,N_34694);
nand U34906 (N_34906,N_34581,N_34602);
xor U34907 (N_34907,N_34660,N_34671);
nor U34908 (N_34908,N_34598,N_34596);
or U34909 (N_34909,N_34598,N_34538);
or U34910 (N_34910,N_34505,N_34624);
or U34911 (N_34911,N_34668,N_34702);
nand U34912 (N_34912,N_34566,N_34643);
nand U34913 (N_34913,N_34680,N_34568);
nor U34914 (N_34914,N_34509,N_34661);
nand U34915 (N_34915,N_34738,N_34667);
or U34916 (N_34916,N_34507,N_34721);
nand U34917 (N_34917,N_34617,N_34660);
xor U34918 (N_34918,N_34528,N_34699);
and U34919 (N_34919,N_34725,N_34539);
nor U34920 (N_34920,N_34632,N_34658);
and U34921 (N_34921,N_34612,N_34629);
nor U34922 (N_34922,N_34549,N_34723);
nand U34923 (N_34923,N_34669,N_34588);
and U34924 (N_34924,N_34648,N_34634);
xnor U34925 (N_34925,N_34725,N_34574);
nor U34926 (N_34926,N_34616,N_34614);
or U34927 (N_34927,N_34734,N_34601);
or U34928 (N_34928,N_34608,N_34684);
or U34929 (N_34929,N_34558,N_34621);
and U34930 (N_34930,N_34706,N_34716);
and U34931 (N_34931,N_34531,N_34726);
nand U34932 (N_34932,N_34530,N_34677);
nand U34933 (N_34933,N_34507,N_34640);
or U34934 (N_34934,N_34707,N_34572);
nand U34935 (N_34935,N_34665,N_34582);
xnor U34936 (N_34936,N_34502,N_34514);
or U34937 (N_34937,N_34622,N_34697);
or U34938 (N_34938,N_34530,N_34682);
or U34939 (N_34939,N_34565,N_34560);
and U34940 (N_34940,N_34730,N_34666);
nand U34941 (N_34941,N_34626,N_34576);
or U34942 (N_34942,N_34705,N_34647);
and U34943 (N_34943,N_34540,N_34627);
or U34944 (N_34944,N_34703,N_34566);
nor U34945 (N_34945,N_34696,N_34601);
or U34946 (N_34946,N_34726,N_34580);
xnor U34947 (N_34947,N_34582,N_34520);
nor U34948 (N_34948,N_34644,N_34564);
and U34949 (N_34949,N_34517,N_34661);
nand U34950 (N_34950,N_34713,N_34691);
nor U34951 (N_34951,N_34658,N_34690);
xor U34952 (N_34952,N_34567,N_34654);
nand U34953 (N_34953,N_34699,N_34672);
or U34954 (N_34954,N_34693,N_34606);
nor U34955 (N_34955,N_34573,N_34699);
and U34956 (N_34956,N_34685,N_34539);
or U34957 (N_34957,N_34548,N_34627);
xnor U34958 (N_34958,N_34742,N_34518);
nand U34959 (N_34959,N_34691,N_34580);
xor U34960 (N_34960,N_34624,N_34684);
xor U34961 (N_34961,N_34516,N_34682);
and U34962 (N_34962,N_34545,N_34634);
and U34963 (N_34963,N_34713,N_34675);
and U34964 (N_34964,N_34584,N_34576);
and U34965 (N_34965,N_34699,N_34708);
xor U34966 (N_34966,N_34694,N_34691);
nor U34967 (N_34967,N_34622,N_34681);
xor U34968 (N_34968,N_34600,N_34563);
nor U34969 (N_34969,N_34679,N_34738);
xor U34970 (N_34970,N_34566,N_34714);
xnor U34971 (N_34971,N_34572,N_34701);
xnor U34972 (N_34972,N_34714,N_34733);
nand U34973 (N_34973,N_34748,N_34609);
nand U34974 (N_34974,N_34701,N_34626);
xnor U34975 (N_34975,N_34591,N_34535);
nor U34976 (N_34976,N_34561,N_34642);
or U34977 (N_34977,N_34527,N_34702);
nand U34978 (N_34978,N_34667,N_34744);
or U34979 (N_34979,N_34745,N_34641);
nand U34980 (N_34980,N_34633,N_34740);
and U34981 (N_34981,N_34741,N_34577);
and U34982 (N_34982,N_34615,N_34524);
nand U34983 (N_34983,N_34521,N_34624);
or U34984 (N_34984,N_34551,N_34556);
and U34985 (N_34985,N_34739,N_34665);
nor U34986 (N_34986,N_34630,N_34518);
nand U34987 (N_34987,N_34501,N_34706);
and U34988 (N_34988,N_34543,N_34678);
nor U34989 (N_34989,N_34683,N_34649);
nor U34990 (N_34990,N_34671,N_34540);
nand U34991 (N_34991,N_34548,N_34516);
or U34992 (N_34992,N_34723,N_34527);
and U34993 (N_34993,N_34730,N_34694);
or U34994 (N_34994,N_34744,N_34604);
nand U34995 (N_34995,N_34509,N_34503);
and U34996 (N_34996,N_34593,N_34640);
xor U34997 (N_34997,N_34566,N_34545);
or U34998 (N_34998,N_34687,N_34576);
and U34999 (N_34999,N_34504,N_34655);
or U35000 (N_35000,N_34990,N_34847);
or U35001 (N_35001,N_34996,N_34916);
and U35002 (N_35002,N_34928,N_34865);
nor U35003 (N_35003,N_34827,N_34887);
or U35004 (N_35004,N_34919,N_34877);
nor U35005 (N_35005,N_34795,N_34857);
or U35006 (N_35006,N_34810,N_34771);
and U35007 (N_35007,N_34960,N_34943);
or U35008 (N_35008,N_34930,N_34811);
xnor U35009 (N_35009,N_34945,N_34859);
or U35010 (N_35010,N_34905,N_34954);
or U35011 (N_35011,N_34777,N_34867);
or U35012 (N_35012,N_34819,N_34883);
and U35013 (N_35013,N_34803,N_34765);
or U35014 (N_35014,N_34763,N_34999);
xnor U35015 (N_35015,N_34947,N_34951);
or U35016 (N_35016,N_34915,N_34938);
nor U35017 (N_35017,N_34845,N_34989);
or U35018 (N_35018,N_34844,N_34910);
xor U35019 (N_35019,N_34935,N_34758);
or U35020 (N_35020,N_34871,N_34812);
nand U35021 (N_35021,N_34965,N_34931);
xor U35022 (N_35022,N_34991,N_34902);
nand U35023 (N_35023,N_34879,N_34782);
xnor U35024 (N_35024,N_34881,N_34799);
xor U35025 (N_35025,N_34833,N_34878);
or U35026 (N_35026,N_34853,N_34988);
nand U35027 (N_35027,N_34775,N_34923);
and U35028 (N_35028,N_34882,N_34900);
nand U35029 (N_35029,N_34884,N_34912);
or U35030 (N_35030,N_34899,N_34970);
nand U35031 (N_35031,N_34851,N_34786);
xor U35032 (N_35032,N_34817,N_34816);
or U35033 (N_35033,N_34903,N_34908);
or U35034 (N_35034,N_34873,N_34805);
and U35035 (N_35035,N_34866,N_34776);
nand U35036 (N_35036,N_34956,N_34751);
or U35037 (N_35037,N_34784,N_34944);
nor U35038 (N_35038,N_34942,N_34924);
or U35039 (N_35039,N_34840,N_34860);
xnor U35040 (N_35040,N_34914,N_34972);
nor U35041 (N_35041,N_34848,N_34750);
and U35042 (N_35042,N_34918,N_34870);
nand U35043 (N_35043,N_34756,N_34774);
nand U35044 (N_35044,N_34779,N_34863);
and U35045 (N_35045,N_34843,N_34966);
or U35046 (N_35046,N_34981,N_34788);
nand U35047 (N_35047,N_34759,N_34936);
nor U35048 (N_35048,N_34933,N_34808);
xnor U35049 (N_35049,N_34909,N_34946);
nand U35050 (N_35050,N_34896,N_34815);
xor U35051 (N_35051,N_34926,N_34868);
and U35052 (N_35052,N_34953,N_34934);
and U35053 (N_35053,N_34984,N_34964);
and U35054 (N_35054,N_34921,N_34772);
nand U35055 (N_35055,N_34838,N_34793);
and U35056 (N_35056,N_34854,N_34801);
nand U35057 (N_35057,N_34757,N_34796);
nor U35058 (N_35058,N_34913,N_34929);
and U35059 (N_35059,N_34969,N_34980);
or U35060 (N_35060,N_34957,N_34783);
nor U35061 (N_35061,N_34925,N_34807);
or U35062 (N_35062,N_34927,N_34895);
and U35063 (N_35063,N_34952,N_34809);
or U35064 (N_35064,N_34804,N_34962);
and U35065 (N_35065,N_34993,N_34897);
and U35066 (N_35066,N_34979,N_34932);
xor U35067 (N_35067,N_34830,N_34820);
and U35068 (N_35068,N_34869,N_34955);
and U35069 (N_35069,N_34985,N_34973);
xnor U35070 (N_35070,N_34861,N_34898);
xor U35071 (N_35071,N_34814,N_34917);
nand U35072 (N_35072,N_34856,N_34849);
nor U35073 (N_35073,N_34813,N_34949);
xnor U35074 (N_35074,N_34904,N_34998);
or U35075 (N_35075,N_34920,N_34858);
or U35076 (N_35076,N_34986,N_34755);
or U35077 (N_35077,N_34790,N_34841);
nor U35078 (N_35078,N_34983,N_34907);
xnor U35079 (N_35079,N_34941,N_34958);
or U35080 (N_35080,N_34778,N_34967);
xor U35081 (N_35081,N_34880,N_34761);
and U35082 (N_35082,N_34976,N_34874);
xor U35083 (N_35083,N_34754,N_34995);
and U35084 (N_35084,N_34842,N_34764);
nor U35085 (N_35085,N_34886,N_34826);
and U35086 (N_35086,N_34906,N_34800);
or U35087 (N_35087,N_34876,N_34922);
and U35088 (N_35088,N_34789,N_34959);
nor U35089 (N_35089,N_34832,N_34974);
and U35090 (N_35090,N_34894,N_34785);
nand U35091 (N_35091,N_34982,N_34791);
and U35092 (N_35092,N_34862,N_34825);
and U35093 (N_35093,N_34839,N_34855);
xor U35094 (N_35094,N_34822,N_34852);
nor U35095 (N_35095,N_34948,N_34836);
nor U35096 (N_35096,N_34864,N_34994);
nor U35097 (N_35097,N_34823,N_34975);
and U35098 (N_35098,N_34939,N_34767);
or U35099 (N_35099,N_34806,N_34831);
and U35100 (N_35100,N_34872,N_34940);
xnor U35101 (N_35101,N_34987,N_34769);
or U35102 (N_35102,N_34950,N_34752);
nor U35103 (N_35103,N_34753,N_34961);
nand U35104 (N_35104,N_34911,N_34766);
or U35105 (N_35105,N_34968,N_34893);
xor U35106 (N_35106,N_34835,N_34792);
or U35107 (N_35107,N_34885,N_34997);
xor U35108 (N_35108,N_34888,N_34797);
and U35109 (N_35109,N_34787,N_34768);
nor U35110 (N_35110,N_34837,N_34828);
xnor U35111 (N_35111,N_34798,N_34992);
and U35112 (N_35112,N_34977,N_34794);
or U35113 (N_35113,N_34937,N_34781);
and U35114 (N_35114,N_34971,N_34890);
and U35115 (N_35115,N_34891,N_34963);
nor U35116 (N_35116,N_34762,N_34829);
and U35117 (N_35117,N_34780,N_34773);
nor U35118 (N_35118,N_34818,N_34892);
or U35119 (N_35119,N_34802,N_34850);
or U35120 (N_35120,N_34978,N_34889);
nand U35121 (N_35121,N_34901,N_34824);
and U35122 (N_35122,N_34760,N_34846);
nor U35123 (N_35123,N_34875,N_34770);
xor U35124 (N_35124,N_34834,N_34821);
or U35125 (N_35125,N_34871,N_34923);
and U35126 (N_35126,N_34787,N_34871);
xnor U35127 (N_35127,N_34957,N_34807);
and U35128 (N_35128,N_34865,N_34993);
nand U35129 (N_35129,N_34911,N_34893);
xnor U35130 (N_35130,N_34860,N_34890);
xnor U35131 (N_35131,N_34776,N_34897);
and U35132 (N_35132,N_34789,N_34820);
and U35133 (N_35133,N_34999,N_34982);
or U35134 (N_35134,N_34953,N_34947);
nor U35135 (N_35135,N_34845,N_34786);
xor U35136 (N_35136,N_34853,N_34976);
and U35137 (N_35137,N_34843,N_34775);
and U35138 (N_35138,N_34874,N_34814);
nand U35139 (N_35139,N_34786,N_34967);
nand U35140 (N_35140,N_34936,N_34951);
or U35141 (N_35141,N_34819,N_34896);
xnor U35142 (N_35142,N_34782,N_34759);
or U35143 (N_35143,N_34913,N_34962);
nor U35144 (N_35144,N_34833,N_34967);
or U35145 (N_35145,N_34801,N_34830);
and U35146 (N_35146,N_34956,N_34986);
xnor U35147 (N_35147,N_34909,N_34826);
nor U35148 (N_35148,N_34991,N_34767);
nor U35149 (N_35149,N_34985,N_34976);
nand U35150 (N_35150,N_34966,N_34958);
or U35151 (N_35151,N_34775,N_34759);
or U35152 (N_35152,N_34969,N_34758);
nor U35153 (N_35153,N_34867,N_34900);
nand U35154 (N_35154,N_34770,N_34972);
or U35155 (N_35155,N_34759,N_34803);
or U35156 (N_35156,N_34991,N_34898);
or U35157 (N_35157,N_34773,N_34864);
nor U35158 (N_35158,N_34789,N_34845);
nor U35159 (N_35159,N_34948,N_34779);
nand U35160 (N_35160,N_34880,N_34796);
or U35161 (N_35161,N_34943,N_34949);
nand U35162 (N_35162,N_34936,N_34958);
xnor U35163 (N_35163,N_34872,N_34881);
or U35164 (N_35164,N_34945,N_34900);
nand U35165 (N_35165,N_34934,N_34949);
and U35166 (N_35166,N_34864,N_34781);
or U35167 (N_35167,N_34882,N_34820);
or U35168 (N_35168,N_34955,N_34865);
nor U35169 (N_35169,N_34829,N_34896);
nor U35170 (N_35170,N_34825,N_34959);
or U35171 (N_35171,N_34775,N_34991);
xnor U35172 (N_35172,N_34958,N_34942);
xor U35173 (N_35173,N_34768,N_34760);
and U35174 (N_35174,N_34866,N_34794);
or U35175 (N_35175,N_34947,N_34857);
and U35176 (N_35176,N_34805,N_34926);
and U35177 (N_35177,N_34924,N_34932);
or U35178 (N_35178,N_34874,N_34838);
nor U35179 (N_35179,N_34913,N_34762);
and U35180 (N_35180,N_34909,N_34850);
xor U35181 (N_35181,N_34903,N_34832);
or U35182 (N_35182,N_34972,N_34924);
xor U35183 (N_35183,N_34856,N_34964);
or U35184 (N_35184,N_34836,N_34804);
nand U35185 (N_35185,N_34964,N_34824);
xor U35186 (N_35186,N_34875,N_34895);
nand U35187 (N_35187,N_34851,N_34982);
or U35188 (N_35188,N_34837,N_34759);
nand U35189 (N_35189,N_34765,N_34981);
nor U35190 (N_35190,N_34793,N_34837);
xnor U35191 (N_35191,N_34792,N_34883);
nor U35192 (N_35192,N_34919,N_34879);
nand U35193 (N_35193,N_34886,N_34871);
nor U35194 (N_35194,N_34768,N_34921);
and U35195 (N_35195,N_34995,N_34962);
or U35196 (N_35196,N_34768,N_34970);
nor U35197 (N_35197,N_34865,N_34788);
or U35198 (N_35198,N_34898,N_34885);
and U35199 (N_35199,N_34916,N_34806);
nand U35200 (N_35200,N_34815,N_34761);
or U35201 (N_35201,N_34990,N_34949);
xor U35202 (N_35202,N_34935,N_34927);
and U35203 (N_35203,N_34887,N_34872);
and U35204 (N_35204,N_34807,N_34846);
or U35205 (N_35205,N_34908,N_34844);
nor U35206 (N_35206,N_34841,N_34865);
and U35207 (N_35207,N_34762,N_34937);
nor U35208 (N_35208,N_34937,N_34907);
and U35209 (N_35209,N_34753,N_34830);
nor U35210 (N_35210,N_34862,N_34954);
and U35211 (N_35211,N_34815,N_34753);
nor U35212 (N_35212,N_34825,N_34931);
xor U35213 (N_35213,N_34932,N_34848);
xor U35214 (N_35214,N_34972,N_34998);
and U35215 (N_35215,N_34971,N_34940);
nor U35216 (N_35216,N_34989,N_34826);
nand U35217 (N_35217,N_34995,N_34758);
xor U35218 (N_35218,N_34975,N_34872);
xor U35219 (N_35219,N_34847,N_34872);
and U35220 (N_35220,N_34800,N_34943);
xnor U35221 (N_35221,N_34899,N_34896);
and U35222 (N_35222,N_34885,N_34909);
nor U35223 (N_35223,N_34813,N_34768);
xnor U35224 (N_35224,N_34778,N_34842);
or U35225 (N_35225,N_34843,N_34949);
or U35226 (N_35226,N_34885,N_34842);
and U35227 (N_35227,N_34844,N_34798);
and U35228 (N_35228,N_34846,N_34912);
and U35229 (N_35229,N_34914,N_34849);
xnor U35230 (N_35230,N_34769,N_34925);
nand U35231 (N_35231,N_34885,N_34762);
and U35232 (N_35232,N_34834,N_34863);
nand U35233 (N_35233,N_34804,N_34875);
and U35234 (N_35234,N_34938,N_34768);
nor U35235 (N_35235,N_34800,N_34903);
nand U35236 (N_35236,N_34812,N_34920);
xnor U35237 (N_35237,N_34842,N_34880);
or U35238 (N_35238,N_34915,N_34876);
nand U35239 (N_35239,N_34802,N_34813);
or U35240 (N_35240,N_34753,N_34997);
or U35241 (N_35241,N_34794,N_34958);
nor U35242 (N_35242,N_34976,N_34979);
and U35243 (N_35243,N_34938,N_34914);
and U35244 (N_35244,N_34773,N_34879);
and U35245 (N_35245,N_34848,N_34852);
or U35246 (N_35246,N_34790,N_34901);
nand U35247 (N_35247,N_34991,N_34882);
nor U35248 (N_35248,N_34774,N_34972);
and U35249 (N_35249,N_34828,N_34761);
or U35250 (N_35250,N_35145,N_35199);
or U35251 (N_35251,N_35006,N_35238);
and U35252 (N_35252,N_35112,N_35063);
nand U35253 (N_35253,N_35229,N_35144);
nor U35254 (N_35254,N_35027,N_35220);
or U35255 (N_35255,N_35175,N_35030);
nand U35256 (N_35256,N_35154,N_35079);
nand U35257 (N_35257,N_35209,N_35182);
and U35258 (N_35258,N_35146,N_35222);
and U35259 (N_35259,N_35106,N_35047);
or U35260 (N_35260,N_35200,N_35014);
and U35261 (N_35261,N_35223,N_35023);
nand U35262 (N_35262,N_35029,N_35031);
xnor U35263 (N_35263,N_35166,N_35129);
or U35264 (N_35264,N_35226,N_35032);
nand U35265 (N_35265,N_35093,N_35102);
or U35266 (N_35266,N_35241,N_35160);
nand U35267 (N_35267,N_35158,N_35099);
nand U35268 (N_35268,N_35138,N_35197);
or U35269 (N_35269,N_35073,N_35140);
or U35270 (N_35270,N_35089,N_35062);
or U35271 (N_35271,N_35204,N_35083);
nand U35272 (N_35272,N_35141,N_35022);
nor U35273 (N_35273,N_35069,N_35207);
and U35274 (N_35274,N_35159,N_35096);
nand U35275 (N_35275,N_35219,N_35080);
and U35276 (N_35276,N_35072,N_35143);
nand U35277 (N_35277,N_35076,N_35009);
nor U35278 (N_35278,N_35167,N_35218);
nand U35279 (N_35279,N_35206,N_35205);
xnor U35280 (N_35280,N_35150,N_35211);
nor U35281 (N_35281,N_35187,N_35246);
nor U35282 (N_35282,N_35021,N_35078);
and U35283 (N_35283,N_35111,N_35248);
and U35284 (N_35284,N_35126,N_35119);
nand U35285 (N_35285,N_35151,N_35245);
xor U35286 (N_35286,N_35217,N_35086);
nand U35287 (N_35287,N_35124,N_35048);
and U35288 (N_35288,N_35004,N_35042);
and U35289 (N_35289,N_35163,N_35149);
or U35290 (N_35290,N_35172,N_35176);
nand U35291 (N_35291,N_35017,N_35095);
or U35292 (N_35292,N_35186,N_35208);
xnor U35293 (N_35293,N_35034,N_35237);
and U35294 (N_35294,N_35087,N_35193);
xnor U35295 (N_35295,N_35066,N_35132);
nor U35296 (N_35296,N_35082,N_35227);
nand U35297 (N_35297,N_35003,N_35170);
xnor U35298 (N_35298,N_35068,N_35008);
or U35299 (N_35299,N_35100,N_35155);
nor U35300 (N_35300,N_35056,N_35188);
and U35301 (N_35301,N_35215,N_35232);
nor U35302 (N_35302,N_35233,N_35247);
and U35303 (N_35303,N_35128,N_35157);
or U35304 (N_35304,N_35152,N_35071);
or U35305 (N_35305,N_35104,N_35016);
nor U35306 (N_35306,N_35212,N_35005);
xnor U35307 (N_35307,N_35050,N_35213);
nor U35308 (N_35308,N_35053,N_35051);
or U35309 (N_35309,N_35044,N_35148);
and U35310 (N_35310,N_35239,N_35007);
and U35311 (N_35311,N_35242,N_35015);
and U35312 (N_35312,N_35130,N_35161);
xor U35313 (N_35313,N_35123,N_35125);
and U35314 (N_35314,N_35025,N_35164);
xnor U35315 (N_35315,N_35088,N_35061);
nand U35316 (N_35316,N_35228,N_35214);
or U35317 (N_35317,N_35018,N_35121);
xnor U35318 (N_35318,N_35216,N_35192);
and U35319 (N_35319,N_35178,N_35235);
nor U35320 (N_35320,N_35179,N_35052);
xor U35321 (N_35321,N_35243,N_35156);
and U35322 (N_35322,N_35024,N_35236);
and U35323 (N_35323,N_35039,N_35105);
xnor U35324 (N_35324,N_35026,N_35181);
nor U35325 (N_35325,N_35040,N_35142);
nor U35326 (N_35326,N_35116,N_35189);
nor U35327 (N_35327,N_35036,N_35169);
or U35328 (N_35328,N_35201,N_35133);
or U35329 (N_35329,N_35127,N_35225);
nor U35330 (N_35330,N_35221,N_35210);
and U35331 (N_35331,N_35075,N_35058);
xnor U35332 (N_35332,N_35117,N_35195);
nor U35333 (N_35333,N_35059,N_35180);
nand U35334 (N_35334,N_35184,N_35135);
nand U35335 (N_35335,N_35131,N_35054);
xnor U35336 (N_35336,N_35173,N_35097);
or U35337 (N_35337,N_35001,N_35012);
or U35338 (N_35338,N_35067,N_35183);
or U35339 (N_35339,N_35098,N_35077);
xnor U35340 (N_35340,N_35139,N_35074);
nand U35341 (N_35341,N_35168,N_35234);
and U35342 (N_35342,N_35120,N_35174);
xor U35343 (N_35343,N_35092,N_35055);
and U35344 (N_35344,N_35060,N_35231);
or U35345 (N_35345,N_35171,N_35064);
or U35346 (N_35346,N_35038,N_35118);
xor U35347 (N_35347,N_35081,N_35103);
and U35348 (N_35348,N_35091,N_35202);
or U35349 (N_35349,N_35043,N_35249);
nand U35350 (N_35350,N_35035,N_35085);
xor U35351 (N_35351,N_35090,N_35203);
xor U35352 (N_35352,N_35194,N_35198);
xor U35353 (N_35353,N_35153,N_35114);
and U35354 (N_35354,N_35190,N_35046);
or U35355 (N_35355,N_35101,N_35177);
or U35356 (N_35356,N_35084,N_35115);
nor U35357 (N_35357,N_35191,N_35049);
and U35358 (N_35358,N_35094,N_35224);
nor U35359 (N_35359,N_35011,N_35147);
nor U35360 (N_35360,N_35041,N_35045);
xnor U35361 (N_35361,N_35037,N_35057);
xor U35362 (N_35362,N_35122,N_35028);
xnor U35363 (N_35363,N_35002,N_35108);
or U35364 (N_35364,N_35196,N_35165);
and U35365 (N_35365,N_35110,N_35240);
nor U35366 (N_35366,N_35137,N_35033);
nor U35367 (N_35367,N_35162,N_35134);
nor U35368 (N_35368,N_35244,N_35013);
nand U35369 (N_35369,N_35113,N_35070);
or U35370 (N_35370,N_35019,N_35107);
nor U35371 (N_35371,N_35020,N_35000);
and U35372 (N_35372,N_35185,N_35065);
and U35373 (N_35373,N_35230,N_35010);
nor U35374 (N_35374,N_35109,N_35136);
nand U35375 (N_35375,N_35145,N_35151);
or U35376 (N_35376,N_35158,N_35215);
or U35377 (N_35377,N_35057,N_35084);
and U35378 (N_35378,N_35038,N_35011);
xor U35379 (N_35379,N_35229,N_35122);
nand U35380 (N_35380,N_35174,N_35043);
and U35381 (N_35381,N_35029,N_35102);
nor U35382 (N_35382,N_35088,N_35056);
nand U35383 (N_35383,N_35219,N_35099);
xnor U35384 (N_35384,N_35056,N_35133);
and U35385 (N_35385,N_35022,N_35019);
and U35386 (N_35386,N_35100,N_35075);
xnor U35387 (N_35387,N_35063,N_35151);
and U35388 (N_35388,N_35013,N_35161);
xnor U35389 (N_35389,N_35105,N_35084);
nand U35390 (N_35390,N_35172,N_35173);
nor U35391 (N_35391,N_35130,N_35198);
nand U35392 (N_35392,N_35226,N_35179);
or U35393 (N_35393,N_35165,N_35174);
xnor U35394 (N_35394,N_35040,N_35158);
nand U35395 (N_35395,N_35183,N_35040);
xor U35396 (N_35396,N_35043,N_35089);
and U35397 (N_35397,N_35151,N_35136);
nand U35398 (N_35398,N_35246,N_35217);
nand U35399 (N_35399,N_35107,N_35138);
or U35400 (N_35400,N_35085,N_35120);
and U35401 (N_35401,N_35034,N_35075);
or U35402 (N_35402,N_35213,N_35102);
nand U35403 (N_35403,N_35043,N_35235);
xnor U35404 (N_35404,N_35176,N_35001);
nor U35405 (N_35405,N_35086,N_35231);
or U35406 (N_35406,N_35213,N_35076);
or U35407 (N_35407,N_35177,N_35000);
nor U35408 (N_35408,N_35038,N_35111);
and U35409 (N_35409,N_35176,N_35106);
and U35410 (N_35410,N_35081,N_35190);
xor U35411 (N_35411,N_35092,N_35102);
xnor U35412 (N_35412,N_35006,N_35226);
and U35413 (N_35413,N_35172,N_35242);
nand U35414 (N_35414,N_35241,N_35010);
nand U35415 (N_35415,N_35155,N_35014);
nand U35416 (N_35416,N_35088,N_35087);
nand U35417 (N_35417,N_35070,N_35178);
xor U35418 (N_35418,N_35167,N_35130);
and U35419 (N_35419,N_35010,N_35164);
and U35420 (N_35420,N_35159,N_35105);
and U35421 (N_35421,N_35142,N_35016);
nor U35422 (N_35422,N_35009,N_35133);
and U35423 (N_35423,N_35144,N_35156);
and U35424 (N_35424,N_35016,N_35183);
or U35425 (N_35425,N_35031,N_35122);
nor U35426 (N_35426,N_35245,N_35041);
nor U35427 (N_35427,N_35178,N_35048);
and U35428 (N_35428,N_35038,N_35246);
and U35429 (N_35429,N_35091,N_35000);
nand U35430 (N_35430,N_35222,N_35119);
nor U35431 (N_35431,N_35091,N_35233);
nand U35432 (N_35432,N_35071,N_35109);
and U35433 (N_35433,N_35225,N_35053);
or U35434 (N_35434,N_35212,N_35101);
nand U35435 (N_35435,N_35216,N_35026);
nand U35436 (N_35436,N_35197,N_35068);
xor U35437 (N_35437,N_35131,N_35006);
nand U35438 (N_35438,N_35170,N_35177);
or U35439 (N_35439,N_35220,N_35002);
nand U35440 (N_35440,N_35182,N_35072);
xnor U35441 (N_35441,N_35123,N_35247);
nand U35442 (N_35442,N_35098,N_35025);
and U35443 (N_35443,N_35082,N_35211);
nor U35444 (N_35444,N_35029,N_35225);
nor U35445 (N_35445,N_35007,N_35238);
or U35446 (N_35446,N_35043,N_35212);
nor U35447 (N_35447,N_35070,N_35235);
nand U35448 (N_35448,N_35086,N_35113);
nor U35449 (N_35449,N_35139,N_35242);
nor U35450 (N_35450,N_35082,N_35216);
xor U35451 (N_35451,N_35162,N_35074);
nor U35452 (N_35452,N_35237,N_35235);
and U35453 (N_35453,N_35027,N_35012);
nand U35454 (N_35454,N_35064,N_35190);
xor U35455 (N_35455,N_35067,N_35053);
and U35456 (N_35456,N_35038,N_35242);
and U35457 (N_35457,N_35001,N_35086);
or U35458 (N_35458,N_35147,N_35060);
or U35459 (N_35459,N_35232,N_35111);
or U35460 (N_35460,N_35032,N_35220);
nor U35461 (N_35461,N_35172,N_35200);
nor U35462 (N_35462,N_35205,N_35221);
or U35463 (N_35463,N_35179,N_35022);
and U35464 (N_35464,N_35203,N_35233);
or U35465 (N_35465,N_35225,N_35064);
nand U35466 (N_35466,N_35155,N_35186);
and U35467 (N_35467,N_35114,N_35225);
or U35468 (N_35468,N_35161,N_35147);
xor U35469 (N_35469,N_35086,N_35059);
or U35470 (N_35470,N_35034,N_35102);
xnor U35471 (N_35471,N_35115,N_35117);
or U35472 (N_35472,N_35213,N_35229);
or U35473 (N_35473,N_35018,N_35059);
nand U35474 (N_35474,N_35139,N_35120);
xnor U35475 (N_35475,N_35097,N_35065);
nand U35476 (N_35476,N_35151,N_35016);
xor U35477 (N_35477,N_35113,N_35158);
nor U35478 (N_35478,N_35128,N_35004);
and U35479 (N_35479,N_35049,N_35153);
and U35480 (N_35480,N_35083,N_35168);
xnor U35481 (N_35481,N_35183,N_35022);
nor U35482 (N_35482,N_35145,N_35247);
and U35483 (N_35483,N_35199,N_35243);
nand U35484 (N_35484,N_35188,N_35149);
and U35485 (N_35485,N_35248,N_35222);
or U35486 (N_35486,N_35127,N_35078);
nand U35487 (N_35487,N_35030,N_35196);
nor U35488 (N_35488,N_35076,N_35101);
or U35489 (N_35489,N_35193,N_35161);
and U35490 (N_35490,N_35047,N_35039);
nor U35491 (N_35491,N_35064,N_35039);
or U35492 (N_35492,N_35156,N_35048);
and U35493 (N_35493,N_35006,N_35033);
and U35494 (N_35494,N_35194,N_35002);
and U35495 (N_35495,N_35177,N_35040);
or U35496 (N_35496,N_35010,N_35005);
or U35497 (N_35497,N_35028,N_35194);
and U35498 (N_35498,N_35049,N_35231);
or U35499 (N_35499,N_35247,N_35133);
xor U35500 (N_35500,N_35450,N_35363);
or U35501 (N_35501,N_35375,N_35297);
and U35502 (N_35502,N_35465,N_35290);
and U35503 (N_35503,N_35344,N_35417);
nor U35504 (N_35504,N_35447,N_35334);
xor U35505 (N_35505,N_35438,N_35341);
nor U35506 (N_35506,N_35361,N_35441);
and U35507 (N_35507,N_35291,N_35423);
or U35508 (N_35508,N_35296,N_35376);
nor U35509 (N_35509,N_35459,N_35373);
nor U35510 (N_35510,N_35427,N_35293);
nor U35511 (N_35511,N_35325,N_35322);
xnor U35512 (N_35512,N_35414,N_35491);
or U35513 (N_35513,N_35475,N_35300);
nor U35514 (N_35514,N_35284,N_35272);
xnor U35515 (N_35515,N_35370,N_35308);
xor U35516 (N_35516,N_35340,N_35330);
xor U35517 (N_35517,N_35401,N_35444);
and U35518 (N_35518,N_35371,N_35472);
or U35519 (N_35519,N_35271,N_35364);
and U35520 (N_35520,N_35396,N_35255);
nand U35521 (N_35521,N_35494,N_35306);
nor U35522 (N_35522,N_35392,N_35493);
or U35523 (N_35523,N_35400,N_35267);
or U35524 (N_35524,N_35264,N_35348);
nand U35525 (N_35525,N_35289,N_35424);
and U35526 (N_35526,N_35421,N_35425);
xnor U35527 (N_35527,N_35266,N_35324);
xor U35528 (N_35528,N_35256,N_35333);
nor U35529 (N_35529,N_35321,N_35426);
xor U35530 (N_35530,N_35270,N_35484);
and U35531 (N_35531,N_35467,N_35395);
xor U35532 (N_35532,N_35335,N_35442);
xor U35533 (N_35533,N_35253,N_35431);
and U35534 (N_35534,N_35269,N_35329);
or U35535 (N_35535,N_35303,N_35357);
nand U35536 (N_35536,N_35474,N_35299);
and U35537 (N_35537,N_35380,N_35323);
xnor U35538 (N_35538,N_35415,N_35430);
and U35539 (N_35539,N_35318,N_35295);
nor U35540 (N_35540,N_35485,N_35469);
nor U35541 (N_35541,N_35352,N_35368);
and U35542 (N_35542,N_35434,N_35405);
nor U35543 (N_35543,N_35429,N_35463);
nor U35544 (N_35544,N_35347,N_35327);
xor U35545 (N_35545,N_35268,N_35372);
or U35546 (N_35546,N_35495,N_35317);
or U35547 (N_35547,N_35278,N_35377);
or U35548 (N_35548,N_35470,N_35409);
and U35549 (N_35549,N_35359,N_35435);
xor U35550 (N_35550,N_35314,N_35259);
and U35551 (N_35551,N_35458,N_35407);
or U35552 (N_35552,N_35411,N_35262);
nand U35553 (N_35553,N_35384,N_35453);
nand U35554 (N_35554,N_35319,N_35446);
and U35555 (N_35555,N_35482,N_35286);
nand U35556 (N_35556,N_35263,N_35275);
and U35557 (N_35557,N_35346,N_35455);
nor U35558 (N_35558,N_35276,N_35331);
or U35559 (N_35559,N_35339,N_35403);
or U35560 (N_35560,N_35413,N_35422);
or U35561 (N_35561,N_35309,N_35287);
nand U35562 (N_35562,N_35252,N_35292);
nand U35563 (N_35563,N_35353,N_35457);
xor U35564 (N_35564,N_35261,N_35260);
nor U35565 (N_35565,N_35315,N_35285);
xor U35566 (N_35566,N_35477,N_35404);
nand U35567 (N_35567,N_35310,N_35320);
or U35568 (N_35568,N_35410,N_35449);
nand U35569 (N_35569,N_35419,N_35250);
xnor U35570 (N_35570,N_35356,N_35464);
and U35571 (N_35571,N_35490,N_35326);
or U35572 (N_35572,N_35265,N_35406);
nand U35573 (N_35573,N_35481,N_35349);
or U35574 (N_35574,N_35478,N_35279);
and U35575 (N_35575,N_35365,N_35468);
xor U35576 (N_35576,N_35328,N_35440);
nand U35577 (N_35577,N_35332,N_35358);
nand U35578 (N_35578,N_35342,N_35288);
xor U35579 (N_35579,N_35302,N_35311);
or U35580 (N_35580,N_35461,N_35312);
or U35581 (N_35581,N_35402,N_35277);
nor U35582 (N_35582,N_35462,N_35433);
or U35583 (N_35583,N_35393,N_35258);
or U35584 (N_35584,N_35369,N_35283);
xnor U35585 (N_35585,N_35350,N_35381);
xor U35586 (N_35586,N_35443,N_35351);
xor U35587 (N_35587,N_35366,N_35298);
or U35588 (N_35588,N_35489,N_35316);
and U35589 (N_35589,N_35378,N_35281);
xnor U35590 (N_35590,N_35394,N_35273);
xor U35591 (N_35591,N_35412,N_35445);
or U35592 (N_35592,N_35498,N_35362);
nor U35593 (N_35593,N_35354,N_35274);
nor U35594 (N_35594,N_35336,N_35471);
and U35595 (N_35595,N_35343,N_35456);
nor U35596 (N_35596,N_35473,N_35488);
or U35597 (N_35597,N_35496,N_35437);
nor U35598 (N_35598,N_35398,N_35428);
xor U35599 (N_35599,N_35388,N_35420);
and U35600 (N_35600,N_35487,N_35408);
or U35601 (N_35601,N_35355,N_35383);
xor U35602 (N_35602,N_35294,N_35466);
nor U35603 (N_35603,N_35476,N_35452);
xor U35604 (N_35604,N_35492,N_35454);
nor U35605 (N_35605,N_35399,N_35307);
xor U35606 (N_35606,N_35499,N_35432);
or U35607 (N_35607,N_35337,N_35374);
nand U35608 (N_35608,N_35390,N_35305);
and U35609 (N_35609,N_35313,N_35460);
nand U35610 (N_35610,N_35382,N_35367);
or U35611 (N_35611,N_35479,N_35385);
nand U35612 (N_35612,N_35280,N_35304);
nor U35613 (N_35613,N_35480,N_35338);
nand U35614 (N_35614,N_35418,N_35486);
xor U35615 (N_35615,N_35451,N_35345);
and U35616 (N_35616,N_35483,N_35251);
nand U35617 (N_35617,N_35448,N_35282);
nor U35618 (N_35618,N_35301,N_35257);
nor U35619 (N_35619,N_35397,N_35379);
nand U35620 (N_35620,N_35254,N_35389);
nor U35621 (N_35621,N_35416,N_35386);
xor U35622 (N_35622,N_35439,N_35436);
or U35623 (N_35623,N_35391,N_35497);
xor U35624 (N_35624,N_35387,N_35360);
nor U35625 (N_35625,N_35351,N_35493);
nor U35626 (N_35626,N_35490,N_35373);
nand U35627 (N_35627,N_35437,N_35450);
xnor U35628 (N_35628,N_35324,N_35342);
and U35629 (N_35629,N_35419,N_35372);
nand U35630 (N_35630,N_35480,N_35405);
nor U35631 (N_35631,N_35273,N_35363);
nand U35632 (N_35632,N_35264,N_35461);
or U35633 (N_35633,N_35405,N_35296);
nor U35634 (N_35634,N_35380,N_35287);
and U35635 (N_35635,N_35282,N_35470);
or U35636 (N_35636,N_35293,N_35497);
nand U35637 (N_35637,N_35267,N_35332);
nor U35638 (N_35638,N_35387,N_35359);
xor U35639 (N_35639,N_35383,N_35319);
or U35640 (N_35640,N_35432,N_35416);
xnor U35641 (N_35641,N_35411,N_35465);
and U35642 (N_35642,N_35401,N_35367);
xnor U35643 (N_35643,N_35492,N_35475);
nand U35644 (N_35644,N_35424,N_35382);
and U35645 (N_35645,N_35432,N_35453);
nor U35646 (N_35646,N_35472,N_35452);
or U35647 (N_35647,N_35437,N_35444);
nand U35648 (N_35648,N_35377,N_35380);
and U35649 (N_35649,N_35267,N_35395);
nand U35650 (N_35650,N_35295,N_35454);
xnor U35651 (N_35651,N_35346,N_35438);
nor U35652 (N_35652,N_35314,N_35422);
or U35653 (N_35653,N_35473,N_35277);
nor U35654 (N_35654,N_35393,N_35422);
nor U35655 (N_35655,N_35303,N_35371);
and U35656 (N_35656,N_35442,N_35351);
and U35657 (N_35657,N_35448,N_35267);
nor U35658 (N_35658,N_35439,N_35349);
and U35659 (N_35659,N_35474,N_35292);
or U35660 (N_35660,N_35316,N_35497);
xor U35661 (N_35661,N_35409,N_35418);
nand U35662 (N_35662,N_35306,N_35298);
or U35663 (N_35663,N_35374,N_35373);
and U35664 (N_35664,N_35289,N_35277);
nor U35665 (N_35665,N_35412,N_35403);
or U35666 (N_35666,N_35385,N_35410);
nor U35667 (N_35667,N_35302,N_35304);
and U35668 (N_35668,N_35330,N_35439);
xor U35669 (N_35669,N_35304,N_35263);
or U35670 (N_35670,N_35341,N_35370);
nor U35671 (N_35671,N_35415,N_35340);
nor U35672 (N_35672,N_35344,N_35437);
nand U35673 (N_35673,N_35322,N_35490);
xnor U35674 (N_35674,N_35272,N_35319);
or U35675 (N_35675,N_35402,N_35337);
and U35676 (N_35676,N_35284,N_35380);
and U35677 (N_35677,N_35305,N_35384);
and U35678 (N_35678,N_35269,N_35460);
xnor U35679 (N_35679,N_35314,N_35270);
and U35680 (N_35680,N_35450,N_35424);
or U35681 (N_35681,N_35411,N_35364);
nand U35682 (N_35682,N_35349,N_35253);
or U35683 (N_35683,N_35320,N_35398);
or U35684 (N_35684,N_35326,N_35489);
nand U35685 (N_35685,N_35270,N_35477);
xnor U35686 (N_35686,N_35488,N_35326);
or U35687 (N_35687,N_35282,N_35289);
nand U35688 (N_35688,N_35398,N_35381);
xnor U35689 (N_35689,N_35304,N_35268);
or U35690 (N_35690,N_35324,N_35487);
nor U35691 (N_35691,N_35424,N_35373);
xor U35692 (N_35692,N_35381,N_35273);
and U35693 (N_35693,N_35335,N_35336);
xor U35694 (N_35694,N_35405,N_35322);
nor U35695 (N_35695,N_35378,N_35343);
nor U35696 (N_35696,N_35260,N_35405);
and U35697 (N_35697,N_35343,N_35372);
nor U35698 (N_35698,N_35361,N_35468);
nand U35699 (N_35699,N_35251,N_35432);
nor U35700 (N_35700,N_35310,N_35366);
or U35701 (N_35701,N_35366,N_35378);
or U35702 (N_35702,N_35254,N_35488);
and U35703 (N_35703,N_35487,N_35463);
nor U35704 (N_35704,N_35420,N_35451);
nor U35705 (N_35705,N_35474,N_35451);
and U35706 (N_35706,N_35391,N_35330);
nor U35707 (N_35707,N_35336,N_35359);
nand U35708 (N_35708,N_35267,N_35406);
or U35709 (N_35709,N_35440,N_35438);
nor U35710 (N_35710,N_35342,N_35276);
nor U35711 (N_35711,N_35333,N_35348);
xor U35712 (N_35712,N_35304,N_35289);
or U35713 (N_35713,N_35303,N_35407);
nor U35714 (N_35714,N_35498,N_35274);
or U35715 (N_35715,N_35263,N_35315);
xor U35716 (N_35716,N_35417,N_35382);
nor U35717 (N_35717,N_35315,N_35388);
nand U35718 (N_35718,N_35338,N_35473);
xor U35719 (N_35719,N_35397,N_35266);
or U35720 (N_35720,N_35285,N_35437);
and U35721 (N_35721,N_35258,N_35461);
xor U35722 (N_35722,N_35436,N_35490);
and U35723 (N_35723,N_35284,N_35449);
or U35724 (N_35724,N_35375,N_35363);
nor U35725 (N_35725,N_35367,N_35275);
or U35726 (N_35726,N_35448,N_35304);
or U35727 (N_35727,N_35480,N_35320);
and U35728 (N_35728,N_35469,N_35404);
or U35729 (N_35729,N_35345,N_35357);
nor U35730 (N_35730,N_35288,N_35328);
and U35731 (N_35731,N_35326,N_35471);
xnor U35732 (N_35732,N_35313,N_35331);
or U35733 (N_35733,N_35308,N_35285);
nor U35734 (N_35734,N_35308,N_35307);
and U35735 (N_35735,N_35269,N_35428);
nor U35736 (N_35736,N_35259,N_35377);
nor U35737 (N_35737,N_35408,N_35484);
nor U35738 (N_35738,N_35312,N_35421);
xor U35739 (N_35739,N_35298,N_35361);
nor U35740 (N_35740,N_35466,N_35275);
and U35741 (N_35741,N_35477,N_35344);
xor U35742 (N_35742,N_35447,N_35378);
xor U35743 (N_35743,N_35333,N_35455);
nand U35744 (N_35744,N_35380,N_35474);
nand U35745 (N_35745,N_35261,N_35292);
xor U35746 (N_35746,N_35485,N_35468);
and U35747 (N_35747,N_35499,N_35261);
and U35748 (N_35748,N_35251,N_35475);
xor U35749 (N_35749,N_35486,N_35366);
xor U35750 (N_35750,N_35574,N_35716);
xor U35751 (N_35751,N_35596,N_35661);
xor U35752 (N_35752,N_35657,N_35723);
nor U35753 (N_35753,N_35659,N_35738);
xnor U35754 (N_35754,N_35650,N_35734);
and U35755 (N_35755,N_35603,N_35578);
xor U35756 (N_35756,N_35515,N_35740);
nand U35757 (N_35757,N_35531,N_35708);
and U35758 (N_35758,N_35538,N_35576);
nor U35759 (N_35759,N_35725,N_35730);
or U35760 (N_35760,N_35720,N_35581);
nor U35761 (N_35761,N_35672,N_35619);
xnor U35762 (N_35762,N_35658,N_35514);
nand U35763 (N_35763,N_35542,N_35742);
nor U35764 (N_35764,N_35605,N_35685);
nand U35765 (N_35765,N_35597,N_35541);
or U35766 (N_35766,N_35662,N_35620);
nor U35767 (N_35767,N_35736,N_35546);
or U35768 (N_35768,N_35711,N_35587);
and U35769 (N_35769,N_35528,N_35694);
and U35770 (N_35770,N_35526,N_35527);
nand U35771 (N_35771,N_35570,N_35640);
and U35772 (N_35772,N_35598,N_35618);
xnor U35773 (N_35773,N_35702,N_35675);
and U35774 (N_35774,N_35713,N_35556);
nor U35775 (N_35775,N_35554,N_35748);
nor U35776 (N_35776,N_35549,N_35586);
and U35777 (N_35777,N_35670,N_35565);
nor U35778 (N_35778,N_35705,N_35683);
or U35779 (N_35779,N_35545,N_35728);
xnor U35780 (N_35780,N_35577,N_35701);
nand U35781 (N_35781,N_35560,N_35647);
nor U35782 (N_35782,N_35590,N_35739);
nand U35783 (N_35783,N_35617,N_35592);
or U35784 (N_35784,N_35572,N_35712);
nor U35785 (N_35785,N_35682,N_35687);
nand U35786 (N_35786,N_35689,N_35709);
nor U35787 (N_35787,N_35536,N_35664);
or U35788 (N_35788,N_35699,N_35563);
nor U35789 (N_35789,N_35645,N_35706);
nand U35790 (N_35790,N_35669,N_35509);
or U35791 (N_35791,N_35743,N_35582);
or U35792 (N_35792,N_35544,N_35573);
nand U35793 (N_35793,N_35630,N_35585);
or U35794 (N_35794,N_35613,N_35506);
nand U35795 (N_35795,N_35633,N_35643);
or U35796 (N_35796,N_35501,N_35601);
xnor U35797 (N_35797,N_35673,N_35677);
nor U35798 (N_35798,N_35550,N_35690);
xnor U35799 (N_35799,N_35636,N_35535);
and U35800 (N_35800,N_35678,N_35626);
and U35801 (N_35801,N_35681,N_35567);
nand U35802 (N_35802,N_35552,N_35517);
or U35803 (N_35803,N_35641,N_35504);
and U35804 (N_35804,N_35609,N_35543);
nor U35805 (N_35805,N_35537,N_35516);
xor U35806 (N_35806,N_35533,N_35676);
xnor U35807 (N_35807,N_35558,N_35653);
xnor U35808 (N_35808,N_35651,N_35741);
and U35809 (N_35809,N_35594,N_35737);
xor U35810 (N_35810,N_35557,N_35732);
nor U35811 (N_35811,N_35566,N_35522);
nand U35812 (N_35812,N_35704,N_35666);
nand U35813 (N_35813,N_35726,N_35608);
xnor U35814 (N_35814,N_35511,N_35724);
or U35815 (N_35815,N_35642,N_35697);
nand U35816 (N_35816,N_35700,N_35513);
nor U35817 (N_35817,N_35680,N_35714);
nor U35818 (N_35818,N_35703,N_35564);
nor U35819 (N_35819,N_35621,N_35646);
and U35820 (N_35820,N_35744,N_35553);
and U35821 (N_35821,N_35721,N_35584);
and U35822 (N_35822,N_35644,N_35695);
or U35823 (N_35823,N_35717,N_35629);
nor U35824 (N_35824,N_35507,N_35634);
and U35825 (N_35825,N_35612,N_35523);
and U35826 (N_35826,N_35631,N_35632);
xor U35827 (N_35827,N_35600,N_35674);
nand U35828 (N_35828,N_35599,N_35604);
nand U35829 (N_35829,N_35745,N_35614);
nor U35830 (N_35830,N_35547,N_35551);
nand U35831 (N_35831,N_35692,N_35607);
nor U35832 (N_35832,N_35512,N_35655);
nor U35833 (N_35833,N_35638,N_35747);
or U35834 (N_35834,N_35671,N_35615);
nand U35835 (N_35835,N_35530,N_35532);
and U35836 (N_35836,N_35707,N_35519);
or U35837 (N_35837,N_35691,N_35505);
and U35838 (N_35838,N_35649,N_35580);
or U35839 (N_35839,N_35710,N_35698);
xor U35840 (N_35840,N_35559,N_35502);
nor U35841 (N_35841,N_35562,N_35568);
and U35842 (N_35842,N_35688,N_35525);
and U35843 (N_35843,N_35718,N_35591);
nand U35844 (N_35844,N_35715,N_35719);
nand U35845 (N_35845,N_35746,N_35555);
nor U35846 (N_35846,N_35654,N_35583);
xnor U35847 (N_35847,N_35733,N_35611);
xor U35848 (N_35848,N_35520,N_35602);
nand U35849 (N_35849,N_35521,N_35508);
nor U35850 (N_35850,N_35727,N_35500);
or U35851 (N_35851,N_35729,N_35595);
nor U35852 (N_35852,N_35665,N_35503);
xor U35853 (N_35853,N_35722,N_35625);
nand U35854 (N_35854,N_35524,N_35548);
nor U35855 (N_35855,N_35668,N_35696);
or U35856 (N_35856,N_35610,N_35623);
nor U35857 (N_35857,N_35606,N_35686);
xnor U35858 (N_35858,N_35684,N_35588);
and U35859 (N_35859,N_35593,N_35529);
or U35860 (N_35860,N_35616,N_35561);
nor U35861 (N_35861,N_35624,N_35652);
nor U35862 (N_35862,N_35627,N_35589);
or U35863 (N_35863,N_35571,N_35628);
and U35864 (N_35864,N_35518,N_35639);
xnor U35865 (N_35865,N_35663,N_35637);
nor U35866 (N_35866,N_35667,N_35534);
xor U35867 (N_35867,N_35648,N_35731);
or U35868 (N_35868,N_35510,N_35660);
nand U35869 (N_35869,N_35635,N_35539);
xnor U35870 (N_35870,N_35735,N_35575);
nand U35871 (N_35871,N_35622,N_35749);
or U35872 (N_35872,N_35656,N_35679);
or U35873 (N_35873,N_35579,N_35569);
or U35874 (N_35874,N_35540,N_35693);
and U35875 (N_35875,N_35575,N_35607);
nor U35876 (N_35876,N_35670,N_35742);
nor U35877 (N_35877,N_35581,N_35552);
and U35878 (N_35878,N_35535,N_35570);
or U35879 (N_35879,N_35707,N_35552);
nand U35880 (N_35880,N_35657,N_35730);
and U35881 (N_35881,N_35555,N_35695);
xor U35882 (N_35882,N_35610,N_35503);
nand U35883 (N_35883,N_35681,N_35603);
and U35884 (N_35884,N_35625,N_35520);
xnor U35885 (N_35885,N_35514,N_35634);
or U35886 (N_35886,N_35545,N_35562);
xnor U35887 (N_35887,N_35747,N_35706);
or U35888 (N_35888,N_35732,N_35733);
and U35889 (N_35889,N_35511,N_35500);
nand U35890 (N_35890,N_35677,N_35538);
or U35891 (N_35891,N_35702,N_35716);
nor U35892 (N_35892,N_35526,N_35634);
nor U35893 (N_35893,N_35508,N_35661);
and U35894 (N_35894,N_35536,N_35707);
and U35895 (N_35895,N_35529,N_35519);
nor U35896 (N_35896,N_35737,N_35692);
and U35897 (N_35897,N_35738,N_35588);
xnor U35898 (N_35898,N_35738,N_35699);
or U35899 (N_35899,N_35671,N_35538);
xor U35900 (N_35900,N_35685,N_35508);
xor U35901 (N_35901,N_35503,N_35561);
and U35902 (N_35902,N_35682,N_35500);
xor U35903 (N_35903,N_35606,N_35621);
and U35904 (N_35904,N_35531,N_35713);
or U35905 (N_35905,N_35516,N_35542);
or U35906 (N_35906,N_35565,N_35530);
nand U35907 (N_35907,N_35730,N_35655);
xnor U35908 (N_35908,N_35715,N_35555);
nor U35909 (N_35909,N_35589,N_35667);
xnor U35910 (N_35910,N_35712,N_35745);
xor U35911 (N_35911,N_35656,N_35533);
xnor U35912 (N_35912,N_35587,N_35657);
and U35913 (N_35913,N_35653,N_35711);
xnor U35914 (N_35914,N_35642,N_35595);
or U35915 (N_35915,N_35674,N_35508);
nor U35916 (N_35916,N_35636,N_35735);
nand U35917 (N_35917,N_35529,N_35744);
or U35918 (N_35918,N_35563,N_35649);
nand U35919 (N_35919,N_35703,N_35746);
and U35920 (N_35920,N_35656,N_35667);
nand U35921 (N_35921,N_35572,N_35521);
nor U35922 (N_35922,N_35643,N_35737);
xor U35923 (N_35923,N_35693,N_35556);
or U35924 (N_35924,N_35529,N_35609);
and U35925 (N_35925,N_35660,N_35617);
and U35926 (N_35926,N_35733,N_35717);
or U35927 (N_35927,N_35502,N_35657);
nor U35928 (N_35928,N_35703,N_35530);
and U35929 (N_35929,N_35504,N_35556);
or U35930 (N_35930,N_35699,N_35593);
nor U35931 (N_35931,N_35506,N_35601);
nand U35932 (N_35932,N_35500,N_35566);
nand U35933 (N_35933,N_35615,N_35706);
nand U35934 (N_35934,N_35548,N_35647);
or U35935 (N_35935,N_35738,N_35580);
or U35936 (N_35936,N_35563,N_35678);
and U35937 (N_35937,N_35501,N_35558);
or U35938 (N_35938,N_35681,N_35668);
or U35939 (N_35939,N_35575,N_35678);
or U35940 (N_35940,N_35521,N_35622);
nor U35941 (N_35941,N_35707,N_35557);
xor U35942 (N_35942,N_35631,N_35664);
nand U35943 (N_35943,N_35666,N_35553);
xor U35944 (N_35944,N_35572,N_35749);
nand U35945 (N_35945,N_35555,N_35576);
and U35946 (N_35946,N_35680,N_35722);
and U35947 (N_35947,N_35529,N_35541);
nand U35948 (N_35948,N_35565,N_35504);
and U35949 (N_35949,N_35564,N_35501);
nor U35950 (N_35950,N_35717,N_35653);
xnor U35951 (N_35951,N_35547,N_35742);
nor U35952 (N_35952,N_35682,N_35524);
xnor U35953 (N_35953,N_35587,N_35704);
or U35954 (N_35954,N_35601,N_35594);
xnor U35955 (N_35955,N_35637,N_35532);
or U35956 (N_35956,N_35688,N_35550);
xor U35957 (N_35957,N_35739,N_35619);
nand U35958 (N_35958,N_35648,N_35528);
nor U35959 (N_35959,N_35741,N_35586);
nor U35960 (N_35960,N_35686,N_35602);
and U35961 (N_35961,N_35538,N_35673);
or U35962 (N_35962,N_35581,N_35611);
and U35963 (N_35963,N_35627,N_35597);
nor U35964 (N_35964,N_35691,N_35581);
nand U35965 (N_35965,N_35732,N_35614);
xnor U35966 (N_35966,N_35665,N_35679);
or U35967 (N_35967,N_35681,N_35594);
xor U35968 (N_35968,N_35536,N_35728);
nand U35969 (N_35969,N_35748,N_35709);
xnor U35970 (N_35970,N_35685,N_35667);
and U35971 (N_35971,N_35639,N_35657);
xnor U35972 (N_35972,N_35680,N_35544);
xnor U35973 (N_35973,N_35656,N_35586);
xor U35974 (N_35974,N_35671,N_35627);
xor U35975 (N_35975,N_35569,N_35503);
nor U35976 (N_35976,N_35536,N_35661);
xnor U35977 (N_35977,N_35563,N_35644);
nand U35978 (N_35978,N_35570,N_35558);
and U35979 (N_35979,N_35537,N_35541);
or U35980 (N_35980,N_35520,N_35607);
nor U35981 (N_35981,N_35644,N_35555);
xnor U35982 (N_35982,N_35518,N_35592);
nand U35983 (N_35983,N_35717,N_35501);
nor U35984 (N_35984,N_35675,N_35667);
and U35985 (N_35985,N_35716,N_35695);
xnor U35986 (N_35986,N_35538,N_35614);
nor U35987 (N_35987,N_35642,N_35741);
xnor U35988 (N_35988,N_35599,N_35588);
and U35989 (N_35989,N_35739,N_35591);
nand U35990 (N_35990,N_35713,N_35665);
nor U35991 (N_35991,N_35614,N_35731);
and U35992 (N_35992,N_35730,N_35669);
nand U35993 (N_35993,N_35695,N_35651);
or U35994 (N_35994,N_35658,N_35511);
or U35995 (N_35995,N_35568,N_35545);
and U35996 (N_35996,N_35571,N_35666);
or U35997 (N_35997,N_35745,N_35735);
nand U35998 (N_35998,N_35654,N_35747);
nand U35999 (N_35999,N_35598,N_35596);
or U36000 (N_36000,N_35815,N_35875);
and U36001 (N_36001,N_35864,N_35774);
or U36002 (N_36002,N_35992,N_35894);
xor U36003 (N_36003,N_35803,N_35999);
and U36004 (N_36004,N_35760,N_35927);
nor U36005 (N_36005,N_35998,N_35898);
nand U36006 (N_36006,N_35833,N_35817);
nor U36007 (N_36007,N_35775,N_35758);
and U36008 (N_36008,N_35928,N_35938);
xor U36009 (N_36009,N_35850,N_35780);
or U36010 (N_36010,N_35810,N_35941);
or U36011 (N_36011,N_35954,N_35931);
xnor U36012 (N_36012,N_35914,N_35912);
or U36013 (N_36013,N_35878,N_35993);
and U36014 (N_36014,N_35777,N_35807);
nand U36015 (N_36015,N_35822,N_35759);
xnor U36016 (N_36016,N_35772,N_35788);
and U36017 (N_36017,N_35784,N_35986);
and U36018 (N_36018,N_35881,N_35769);
or U36019 (N_36019,N_35849,N_35861);
nand U36020 (N_36020,N_35791,N_35972);
nand U36021 (N_36021,N_35820,N_35761);
nor U36022 (N_36022,N_35805,N_35799);
nand U36023 (N_36023,N_35802,N_35856);
nand U36024 (N_36024,N_35766,N_35787);
nand U36025 (N_36025,N_35924,N_35955);
and U36026 (N_36026,N_35909,N_35841);
nand U36027 (N_36027,N_35773,N_35916);
nand U36028 (N_36028,N_35786,N_35907);
xnor U36029 (N_36029,N_35939,N_35763);
or U36030 (N_36030,N_35872,N_35838);
and U36031 (N_36031,N_35940,N_35923);
nor U36032 (N_36032,N_35771,N_35969);
nand U36033 (N_36033,N_35971,N_35997);
and U36034 (N_36034,N_35885,N_35982);
xnor U36035 (N_36035,N_35779,N_35935);
nor U36036 (N_36036,N_35855,N_35970);
nor U36037 (N_36037,N_35801,N_35937);
xor U36038 (N_36038,N_35858,N_35844);
nor U36039 (N_36039,N_35996,N_35988);
nand U36040 (N_36040,N_35756,N_35863);
or U36041 (N_36041,N_35889,N_35948);
and U36042 (N_36042,N_35910,N_35753);
and U36043 (N_36043,N_35843,N_35798);
or U36044 (N_36044,N_35950,N_35812);
nor U36045 (N_36045,N_35943,N_35831);
nand U36046 (N_36046,N_35977,N_35987);
nand U36047 (N_36047,N_35911,N_35897);
nor U36048 (N_36048,N_35949,N_35925);
nor U36049 (N_36049,N_35966,N_35946);
nor U36050 (N_36050,N_35917,N_35860);
or U36051 (N_36051,N_35837,N_35961);
or U36052 (N_36052,N_35976,N_35932);
or U36053 (N_36053,N_35904,N_35944);
and U36054 (N_36054,N_35962,N_35990);
xor U36055 (N_36055,N_35770,N_35785);
or U36056 (N_36056,N_35828,N_35752);
nor U36057 (N_36057,N_35884,N_35876);
nand U36058 (N_36058,N_35975,N_35792);
and U36059 (N_36059,N_35978,N_35765);
or U36060 (N_36060,N_35845,N_35768);
and U36061 (N_36061,N_35887,N_35930);
nand U36062 (N_36062,N_35965,N_35764);
and U36063 (N_36063,N_35933,N_35834);
nand U36064 (N_36064,N_35757,N_35981);
or U36065 (N_36065,N_35936,N_35958);
nand U36066 (N_36066,N_35879,N_35829);
and U36067 (N_36067,N_35794,N_35811);
or U36068 (N_36068,N_35918,N_35926);
and U36069 (N_36069,N_35960,N_35877);
and U36070 (N_36070,N_35821,N_35824);
nand U36071 (N_36071,N_35825,N_35797);
nand U36072 (N_36072,N_35813,N_35953);
nor U36073 (N_36073,N_35754,N_35886);
xnor U36074 (N_36074,N_35819,N_35985);
and U36075 (N_36075,N_35795,N_35854);
or U36076 (N_36076,N_35867,N_35900);
nor U36077 (N_36077,N_35891,N_35846);
or U36078 (N_36078,N_35852,N_35956);
xnor U36079 (N_36079,N_35903,N_35873);
xor U36080 (N_36080,N_35991,N_35751);
nor U36081 (N_36081,N_35832,N_35871);
and U36082 (N_36082,N_35967,N_35989);
nand U36083 (N_36083,N_35848,N_35806);
nor U36084 (N_36084,N_35951,N_35793);
and U36085 (N_36085,N_35823,N_35915);
or U36086 (N_36086,N_35826,N_35908);
xor U36087 (N_36087,N_35840,N_35893);
or U36088 (N_36088,N_35995,N_35776);
nand U36089 (N_36089,N_35870,N_35809);
or U36090 (N_36090,N_35974,N_35880);
nand U36091 (N_36091,N_35901,N_35851);
or U36092 (N_36092,N_35947,N_35892);
and U36093 (N_36093,N_35866,N_35919);
xnor U36094 (N_36094,N_35882,N_35913);
nor U36095 (N_36095,N_35808,N_35839);
xor U36096 (N_36096,N_35963,N_35862);
or U36097 (N_36097,N_35874,N_35964);
or U36098 (N_36098,N_35790,N_35781);
nor U36099 (N_36099,N_35869,N_35800);
nor U36100 (N_36100,N_35973,N_35994);
nand U36101 (N_36101,N_35929,N_35853);
xor U36102 (N_36102,N_35818,N_35783);
nand U36103 (N_36103,N_35762,N_35835);
and U36104 (N_36104,N_35827,N_35957);
nor U36105 (N_36105,N_35899,N_35814);
xor U36106 (N_36106,N_35921,N_35959);
or U36107 (N_36107,N_35984,N_35942);
or U36108 (N_36108,N_35842,N_35755);
xor U36109 (N_36109,N_35952,N_35934);
xnor U36110 (N_36110,N_35782,N_35906);
and U36111 (N_36111,N_35888,N_35902);
xnor U36112 (N_36112,N_35859,N_35750);
nor U36113 (N_36113,N_35890,N_35905);
nor U36114 (N_36114,N_35836,N_35922);
nor U36115 (N_36115,N_35896,N_35816);
or U36116 (N_36116,N_35980,N_35789);
nand U36117 (N_36117,N_35865,N_35857);
nand U36118 (N_36118,N_35945,N_35920);
and U36119 (N_36119,N_35847,N_35767);
and U36120 (N_36120,N_35883,N_35796);
and U36121 (N_36121,N_35830,N_35979);
or U36122 (N_36122,N_35804,N_35868);
or U36123 (N_36123,N_35983,N_35778);
or U36124 (N_36124,N_35895,N_35968);
or U36125 (N_36125,N_35927,N_35831);
or U36126 (N_36126,N_35876,N_35874);
and U36127 (N_36127,N_35784,N_35867);
xnor U36128 (N_36128,N_35751,N_35937);
xor U36129 (N_36129,N_35958,N_35867);
and U36130 (N_36130,N_35802,N_35852);
and U36131 (N_36131,N_35865,N_35903);
xor U36132 (N_36132,N_35855,N_35938);
or U36133 (N_36133,N_35878,N_35844);
or U36134 (N_36134,N_35780,N_35911);
or U36135 (N_36135,N_35782,N_35843);
nand U36136 (N_36136,N_35777,N_35939);
nor U36137 (N_36137,N_35869,N_35874);
xor U36138 (N_36138,N_35778,N_35920);
and U36139 (N_36139,N_35916,N_35887);
or U36140 (N_36140,N_35795,N_35953);
or U36141 (N_36141,N_35804,N_35979);
or U36142 (N_36142,N_35768,N_35879);
nand U36143 (N_36143,N_35815,N_35829);
nand U36144 (N_36144,N_35884,N_35825);
nor U36145 (N_36145,N_35866,N_35821);
and U36146 (N_36146,N_35878,N_35869);
and U36147 (N_36147,N_35957,N_35935);
nor U36148 (N_36148,N_35813,N_35926);
nor U36149 (N_36149,N_35930,N_35965);
nor U36150 (N_36150,N_35829,N_35855);
or U36151 (N_36151,N_35887,N_35816);
xnor U36152 (N_36152,N_35894,N_35930);
nand U36153 (N_36153,N_35936,N_35896);
xnor U36154 (N_36154,N_35851,N_35793);
nor U36155 (N_36155,N_35882,N_35808);
nand U36156 (N_36156,N_35899,N_35970);
or U36157 (N_36157,N_35803,N_35878);
xor U36158 (N_36158,N_35945,N_35931);
nor U36159 (N_36159,N_35800,N_35909);
nor U36160 (N_36160,N_35877,N_35853);
nand U36161 (N_36161,N_35824,N_35807);
nor U36162 (N_36162,N_35771,N_35850);
nand U36163 (N_36163,N_35986,N_35750);
or U36164 (N_36164,N_35864,N_35805);
nand U36165 (N_36165,N_35955,N_35940);
xnor U36166 (N_36166,N_35855,N_35797);
or U36167 (N_36167,N_35981,N_35972);
and U36168 (N_36168,N_35919,N_35822);
xor U36169 (N_36169,N_35790,N_35813);
xor U36170 (N_36170,N_35963,N_35895);
xor U36171 (N_36171,N_35892,N_35836);
xor U36172 (N_36172,N_35804,N_35782);
nand U36173 (N_36173,N_35816,N_35998);
or U36174 (N_36174,N_35995,N_35781);
xnor U36175 (N_36175,N_35790,N_35879);
nand U36176 (N_36176,N_35861,N_35800);
xor U36177 (N_36177,N_35845,N_35980);
nand U36178 (N_36178,N_35995,N_35993);
or U36179 (N_36179,N_35801,N_35802);
nand U36180 (N_36180,N_35942,N_35923);
xor U36181 (N_36181,N_35981,N_35803);
or U36182 (N_36182,N_35766,N_35881);
or U36183 (N_36183,N_35989,N_35768);
nand U36184 (N_36184,N_35768,N_35755);
and U36185 (N_36185,N_35809,N_35917);
or U36186 (N_36186,N_35905,N_35762);
or U36187 (N_36187,N_35889,N_35967);
and U36188 (N_36188,N_35849,N_35799);
and U36189 (N_36189,N_35816,N_35907);
or U36190 (N_36190,N_35832,N_35782);
xnor U36191 (N_36191,N_35825,N_35876);
or U36192 (N_36192,N_35811,N_35931);
nand U36193 (N_36193,N_35813,N_35969);
nor U36194 (N_36194,N_35938,N_35781);
and U36195 (N_36195,N_35830,N_35822);
xnor U36196 (N_36196,N_35902,N_35933);
nand U36197 (N_36197,N_35802,N_35945);
nor U36198 (N_36198,N_35971,N_35813);
nor U36199 (N_36199,N_35985,N_35785);
nor U36200 (N_36200,N_35775,N_35878);
nor U36201 (N_36201,N_35820,N_35759);
xor U36202 (N_36202,N_35772,N_35867);
nand U36203 (N_36203,N_35923,N_35892);
or U36204 (N_36204,N_35751,N_35994);
or U36205 (N_36205,N_35851,N_35751);
xor U36206 (N_36206,N_35911,N_35980);
xnor U36207 (N_36207,N_35766,N_35964);
and U36208 (N_36208,N_35766,N_35892);
xor U36209 (N_36209,N_35857,N_35830);
or U36210 (N_36210,N_35761,N_35837);
nor U36211 (N_36211,N_35859,N_35762);
or U36212 (N_36212,N_35994,N_35834);
or U36213 (N_36213,N_35862,N_35900);
or U36214 (N_36214,N_35764,N_35802);
nor U36215 (N_36215,N_35894,N_35805);
xnor U36216 (N_36216,N_35761,N_35910);
and U36217 (N_36217,N_35914,N_35750);
and U36218 (N_36218,N_35948,N_35773);
xor U36219 (N_36219,N_35868,N_35752);
xnor U36220 (N_36220,N_35759,N_35961);
or U36221 (N_36221,N_35936,N_35917);
xnor U36222 (N_36222,N_35938,N_35969);
or U36223 (N_36223,N_35899,N_35829);
or U36224 (N_36224,N_35777,N_35995);
nand U36225 (N_36225,N_35869,N_35762);
xnor U36226 (N_36226,N_35764,N_35918);
xor U36227 (N_36227,N_35916,N_35803);
nor U36228 (N_36228,N_35812,N_35887);
nor U36229 (N_36229,N_35811,N_35870);
and U36230 (N_36230,N_35762,N_35911);
nor U36231 (N_36231,N_35822,N_35816);
or U36232 (N_36232,N_35808,N_35961);
or U36233 (N_36233,N_35869,N_35766);
nor U36234 (N_36234,N_35760,N_35932);
xor U36235 (N_36235,N_35821,N_35975);
or U36236 (N_36236,N_35894,N_35777);
nand U36237 (N_36237,N_35929,N_35763);
nand U36238 (N_36238,N_35822,N_35761);
and U36239 (N_36239,N_35820,N_35888);
nor U36240 (N_36240,N_35985,N_35813);
nor U36241 (N_36241,N_35763,N_35765);
or U36242 (N_36242,N_35752,N_35895);
xnor U36243 (N_36243,N_35788,N_35880);
nand U36244 (N_36244,N_35878,N_35756);
xnor U36245 (N_36245,N_35980,N_35853);
nor U36246 (N_36246,N_35918,N_35762);
and U36247 (N_36247,N_35818,N_35881);
xnor U36248 (N_36248,N_35815,N_35941);
or U36249 (N_36249,N_35970,N_35912);
or U36250 (N_36250,N_36074,N_36141);
and U36251 (N_36251,N_36058,N_36092);
xnor U36252 (N_36252,N_36121,N_36117);
nand U36253 (N_36253,N_36203,N_36209);
nor U36254 (N_36254,N_36132,N_36054);
nor U36255 (N_36255,N_36165,N_36068);
nor U36256 (N_36256,N_36113,N_36157);
or U36257 (N_36257,N_36221,N_36156);
xor U36258 (N_36258,N_36016,N_36148);
and U36259 (N_36259,N_36226,N_36222);
xor U36260 (N_36260,N_36029,N_36109);
nor U36261 (N_36261,N_36015,N_36235);
xor U36262 (N_36262,N_36038,N_36133);
xnor U36263 (N_36263,N_36183,N_36005);
or U36264 (N_36264,N_36135,N_36212);
and U36265 (N_36265,N_36033,N_36245);
nand U36266 (N_36266,N_36006,N_36193);
nor U36267 (N_36267,N_36224,N_36014);
xor U36268 (N_36268,N_36030,N_36126);
nand U36269 (N_36269,N_36137,N_36067);
nor U36270 (N_36270,N_36198,N_36205);
nand U36271 (N_36271,N_36060,N_36150);
or U36272 (N_36272,N_36242,N_36097);
or U36273 (N_36273,N_36111,N_36227);
and U36274 (N_36274,N_36025,N_36059);
nor U36275 (N_36275,N_36062,N_36179);
nor U36276 (N_36276,N_36050,N_36238);
or U36277 (N_36277,N_36246,N_36065);
nand U36278 (N_36278,N_36087,N_36035);
xnor U36279 (N_36279,N_36241,N_36129);
nor U36280 (N_36280,N_36239,N_36151);
nor U36281 (N_36281,N_36194,N_36088);
nor U36282 (N_36282,N_36041,N_36237);
and U36283 (N_36283,N_36028,N_36158);
or U36284 (N_36284,N_36103,N_36191);
or U36285 (N_36285,N_36124,N_36098);
xor U36286 (N_36286,N_36223,N_36144);
and U36287 (N_36287,N_36002,N_36022);
or U36288 (N_36288,N_36176,N_36232);
and U36289 (N_36289,N_36108,N_36114);
and U36290 (N_36290,N_36130,N_36011);
or U36291 (N_36291,N_36163,N_36142);
and U36292 (N_36292,N_36192,N_36009);
xnor U36293 (N_36293,N_36112,N_36147);
nand U36294 (N_36294,N_36082,N_36159);
and U36295 (N_36295,N_36024,N_36136);
nand U36296 (N_36296,N_36043,N_36120);
xnor U36297 (N_36297,N_36013,N_36220);
and U36298 (N_36298,N_36155,N_36240);
nand U36299 (N_36299,N_36116,N_36107);
nor U36300 (N_36300,N_36243,N_36077);
xnor U36301 (N_36301,N_36021,N_36228);
nor U36302 (N_36302,N_36083,N_36233);
xnor U36303 (N_36303,N_36091,N_36230);
nor U36304 (N_36304,N_36064,N_36051);
xnor U36305 (N_36305,N_36036,N_36052);
and U36306 (N_36306,N_36076,N_36131);
and U36307 (N_36307,N_36018,N_36187);
nand U36308 (N_36308,N_36169,N_36095);
nand U36309 (N_36309,N_36061,N_36184);
xor U36310 (N_36310,N_36105,N_36219);
or U36311 (N_36311,N_36177,N_36081);
or U36312 (N_36312,N_36229,N_36185);
and U36313 (N_36313,N_36085,N_36110);
nor U36314 (N_36314,N_36249,N_36201);
nand U36315 (N_36315,N_36231,N_36215);
nor U36316 (N_36316,N_36166,N_36053);
or U36317 (N_36317,N_36217,N_36040);
nand U36318 (N_36318,N_36200,N_36034);
nand U36319 (N_36319,N_36216,N_36213);
and U36320 (N_36320,N_36047,N_36000);
xor U36321 (N_36321,N_36017,N_36099);
nand U36322 (N_36322,N_36075,N_36182);
and U36323 (N_36323,N_36211,N_36102);
nor U36324 (N_36324,N_36174,N_36004);
and U36325 (N_36325,N_36057,N_36045);
or U36326 (N_36326,N_36139,N_36196);
or U36327 (N_36327,N_36101,N_36180);
nand U36328 (N_36328,N_36001,N_36042);
nand U36329 (N_36329,N_36199,N_36072);
and U36330 (N_36330,N_36167,N_36093);
or U36331 (N_36331,N_36188,N_36078);
and U36332 (N_36332,N_36037,N_36080);
nor U36333 (N_36333,N_36066,N_36234);
or U36334 (N_36334,N_36032,N_36189);
or U36335 (N_36335,N_36170,N_36178);
nor U36336 (N_36336,N_36007,N_36044);
nand U36337 (N_36337,N_36162,N_36046);
nand U36338 (N_36338,N_36154,N_36063);
nor U36339 (N_36339,N_36161,N_36086);
xor U36340 (N_36340,N_36026,N_36008);
nand U36341 (N_36341,N_36190,N_36115);
nand U36342 (N_36342,N_36127,N_36084);
and U36343 (N_36343,N_36181,N_36244);
or U36344 (N_36344,N_36123,N_36056);
xor U36345 (N_36345,N_36225,N_36206);
or U36346 (N_36346,N_36248,N_36039);
xor U36347 (N_36347,N_36106,N_36145);
and U36348 (N_36348,N_36055,N_36010);
nand U36349 (N_36349,N_36027,N_36204);
or U36350 (N_36350,N_36100,N_36175);
xnor U36351 (N_36351,N_36143,N_36128);
and U36352 (N_36352,N_36079,N_36104);
nand U36353 (N_36353,N_36207,N_36247);
or U36354 (N_36354,N_36012,N_36171);
and U36355 (N_36355,N_36172,N_36149);
nand U36356 (N_36356,N_36089,N_36125);
xor U36357 (N_36357,N_36134,N_36094);
or U36358 (N_36358,N_36119,N_36214);
xnor U36359 (N_36359,N_36069,N_36023);
or U36360 (N_36360,N_36195,N_36073);
or U36361 (N_36361,N_36173,N_36122);
xor U36362 (N_36362,N_36202,N_36020);
or U36363 (N_36363,N_36218,N_36118);
and U36364 (N_36364,N_36146,N_36208);
nand U36365 (N_36365,N_36160,N_36186);
and U36366 (N_36366,N_36048,N_36168);
xor U36367 (N_36367,N_36003,N_36236);
and U36368 (N_36368,N_36152,N_36138);
xor U36369 (N_36369,N_36090,N_36153);
and U36370 (N_36370,N_36071,N_36070);
or U36371 (N_36371,N_36210,N_36049);
nor U36372 (N_36372,N_36197,N_36140);
and U36373 (N_36373,N_36164,N_36096);
or U36374 (N_36374,N_36019,N_36031);
nor U36375 (N_36375,N_36219,N_36161);
and U36376 (N_36376,N_36008,N_36135);
xnor U36377 (N_36377,N_36202,N_36209);
or U36378 (N_36378,N_36184,N_36020);
and U36379 (N_36379,N_36113,N_36137);
nand U36380 (N_36380,N_36051,N_36240);
nor U36381 (N_36381,N_36127,N_36182);
nand U36382 (N_36382,N_36234,N_36150);
nor U36383 (N_36383,N_36043,N_36073);
and U36384 (N_36384,N_36111,N_36182);
xnor U36385 (N_36385,N_36156,N_36155);
xnor U36386 (N_36386,N_36198,N_36246);
or U36387 (N_36387,N_36044,N_36196);
or U36388 (N_36388,N_36107,N_36109);
nor U36389 (N_36389,N_36157,N_36180);
and U36390 (N_36390,N_36116,N_36000);
xor U36391 (N_36391,N_36225,N_36122);
xor U36392 (N_36392,N_36196,N_36110);
and U36393 (N_36393,N_36177,N_36218);
nor U36394 (N_36394,N_36023,N_36214);
xnor U36395 (N_36395,N_36062,N_36003);
nand U36396 (N_36396,N_36163,N_36062);
nor U36397 (N_36397,N_36119,N_36077);
and U36398 (N_36398,N_36145,N_36050);
xnor U36399 (N_36399,N_36108,N_36166);
nor U36400 (N_36400,N_36138,N_36071);
or U36401 (N_36401,N_36157,N_36234);
nor U36402 (N_36402,N_36036,N_36048);
and U36403 (N_36403,N_36113,N_36134);
or U36404 (N_36404,N_36103,N_36193);
nor U36405 (N_36405,N_36070,N_36209);
xor U36406 (N_36406,N_36048,N_36155);
and U36407 (N_36407,N_36186,N_36180);
or U36408 (N_36408,N_36006,N_36249);
nand U36409 (N_36409,N_36009,N_36172);
and U36410 (N_36410,N_36077,N_36246);
nor U36411 (N_36411,N_36015,N_36048);
and U36412 (N_36412,N_36236,N_36030);
nor U36413 (N_36413,N_36231,N_36246);
xnor U36414 (N_36414,N_36085,N_36089);
or U36415 (N_36415,N_36204,N_36154);
or U36416 (N_36416,N_36108,N_36236);
nor U36417 (N_36417,N_36204,N_36069);
nor U36418 (N_36418,N_36205,N_36207);
nand U36419 (N_36419,N_36107,N_36117);
and U36420 (N_36420,N_36181,N_36164);
xnor U36421 (N_36421,N_36098,N_36118);
nand U36422 (N_36422,N_36152,N_36144);
nand U36423 (N_36423,N_36189,N_36022);
nor U36424 (N_36424,N_36100,N_36192);
nand U36425 (N_36425,N_36042,N_36009);
and U36426 (N_36426,N_36078,N_36122);
xnor U36427 (N_36427,N_36231,N_36180);
nor U36428 (N_36428,N_36085,N_36163);
nand U36429 (N_36429,N_36054,N_36009);
xnor U36430 (N_36430,N_36234,N_36196);
nor U36431 (N_36431,N_36239,N_36012);
nand U36432 (N_36432,N_36055,N_36035);
or U36433 (N_36433,N_36173,N_36149);
nor U36434 (N_36434,N_36130,N_36185);
or U36435 (N_36435,N_36247,N_36230);
nand U36436 (N_36436,N_36000,N_36106);
nand U36437 (N_36437,N_36177,N_36130);
and U36438 (N_36438,N_36001,N_36008);
and U36439 (N_36439,N_36060,N_36232);
xnor U36440 (N_36440,N_36143,N_36040);
nand U36441 (N_36441,N_36173,N_36086);
nor U36442 (N_36442,N_36041,N_36082);
xnor U36443 (N_36443,N_36069,N_36107);
nor U36444 (N_36444,N_36209,N_36161);
nand U36445 (N_36445,N_36170,N_36229);
nand U36446 (N_36446,N_36031,N_36005);
xnor U36447 (N_36447,N_36242,N_36001);
nand U36448 (N_36448,N_36168,N_36208);
xor U36449 (N_36449,N_36236,N_36010);
and U36450 (N_36450,N_36173,N_36132);
or U36451 (N_36451,N_36188,N_36111);
or U36452 (N_36452,N_36001,N_36193);
xor U36453 (N_36453,N_36167,N_36040);
xor U36454 (N_36454,N_36203,N_36089);
or U36455 (N_36455,N_36045,N_36244);
or U36456 (N_36456,N_36121,N_36073);
or U36457 (N_36457,N_36236,N_36201);
and U36458 (N_36458,N_36127,N_36244);
xor U36459 (N_36459,N_36066,N_36230);
and U36460 (N_36460,N_36070,N_36015);
nor U36461 (N_36461,N_36041,N_36167);
xnor U36462 (N_36462,N_36018,N_36152);
nand U36463 (N_36463,N_36123,N_36098);
or U36464 (N_36464,N_36022,N_36176);
and U36465 (N_36465,N_36197,N_36173);
or U36466 (N_36466,N_36179,N_36156);
or U36467 (N_36467,N_36011,N_36097);
and U36468 (N_36468,N_36163,N_36165);
and U36469 (N_36469,N_36241,N_36221);
and U36470 (N_36470,N_36041,N_36205);
nand U36471 (N_36471,N_36189,N_36143);
nand U36472 (N_36472,N_36026,N_36078);
or U36473 (N_36473,N_36243,N_36200);
nor U36474 (N_36474,N_36066,N_36140);
and U36475 (N_36475,N_36133,N_36190);
nor U36476 (N_36476,N_36105,N_36182);
or U36477 (N_36477,N_36220,N_36030);
or U36478 (N_36478,N_36208,N_36055);
nor U36479 (N_36479,N_36112,N_36176);
nand U36480 (N_36480,N_36056,N_36079);
or U36481 (N_36481,N_36244,N_36010);
nand U36482 (N_36482,N_36087,N_36148);
nor U36483 (N_36483,N_36129,N_36155);
nand U36484 (N_36484,N_36110,N_36020);
or U36485 (N_36485,N_36055,N_36192);
nor U36486 (N_36486,N_36113,N_36142);
or U36487 (N_36487,N_36102,N_36099);
and U36488 (N_36488,N_36053,N_36078);
nand U36489 (N_36489,N_36228,N_36174);
and U36490 (N_36490,N_36150,N_36010);
or U36491 (N_36491,N_36001,N_36144);
xnor U36492 (N_36492,N_36244,N_36202);
or U36493 (N_36493,N_36153,N_36217);
nor U36494 (N_36494,N_36081,N_36054);
nand U36495 (N_36495,N_36130,N_36023);
nand U36496 (N_36496,N_36068,N_36022);
xor U36497 (N_36497,N_36081,N_36214);
or U36498 (N_36498,N_36180,N_36236);
nand U36499 (N_36499,N_36112,N_36182);
nor U36500 (N_36500,N_36339,N_36482);
nor U36501 (N_36501,N_36471,N_36300);
and U36502 (N_36502,N_36402,N_36458);
nor U36503 (N_36503,N_36362,N_36307);
nand U36504 (N_36504,N_36407,N_36318);
and U36505 (N_36505,N_36381,N_36495);
nand U36506 (N_36506,N_36385,N_36480);
and U36507 (N_36507,N_36330,N_36391);
xor U36508 (N_36508,N_36282,N_36259);
nand U36509 (N_36509,N_36409,N_36323);
xnor U36510 (N_36510,N_36411,N_36379);
nor U36511 (N_36511,N_36461,N_36447);
nand U36512 (N_36512,N_36271,N_36489);
nand U36513 (N_36513,N_36256,N_36298);
xor U36514 (N_36514,N_36416,N_36451);
nor U36515 (N_36515,N_36436,N_36483);
nor U36516 (N_36516,N_36467,N_36493);
nand U36517 (N_36517,N_36358,N_36392);
and U36518 (N_36518,N_36291,N_36327);
xnor U36519 (N_36519,N_36341,N_36405);
xnor U36520 (N_36520,N_36315,N_36253);
and U36521 (N_36521,N_36410,N_36476);
nand U36522 (N_36522,N_36284,N_36338);
xnor U36523 (N_36523,N_36439,N_36463);
nand U36524 (N_36524,N_36262,N_36399);
and U36525 (N_36525,N_36430,N_36359);
nand U36526 (N_36526,N_36268,N_36373);
nor U36527 (N_36527,N_36316,N_36412);
xor U36528 (N_36528,N_36403,N_36478);
nor U36529 (N_36529,N_36277,N_36349);
or U36530 (N_36530,N_36365,N_36356);
xnor U36531 (N_36531,N_36440,N_36292);
or U36532 (N_36532,N_36374,N_36283);
and U36533 (N_36533,N_36433,N_36276);
and U36534 (N_36534,N_36331,N_36443);
nor U36535 (N_36535,N_36293,N_36345);
and U36536 (N_36536,N_36325,N_36352);
xnor U36537 (N_36537,N_36472,N_36322);
nand U36538 (N_36538,N_36372,N_36479);
and U36539 (N_36539,N_36384,N_36460);
or U36540 (N_36540,N_36360,N_36260);
xor U36541 (N_36541,N_36425,N_36441);
and U36542 (N_36542,N_36326,N_36272);
xnor U36543 (N_36543,N_36492,N_36438);
xnor U36544 (N_36544,N_36287,N_36328);
nor U36545 (N_36545,N_36367,N_36308);
and U36546 (N_36546,N_36361,N_36408);
or U36547 (N_36547,N_36387,N_36446);
nor U36548 (N_36548,N_36487,N_36305);
xor U36549 (N_36549,N_36275,N_36313);
nor U36550 (N_36550,N_36452,N_36497);
or U36551 (N_36551,N_36398,N_36469);
nor U36552 (N_36552,N_36484,N_36258);
and U36553 (N_36553,N_36317,N_36335);
nor U36554 (N_36554,N_36473,N_36429);
or U36555 (N_36555,N_36375,N_36422);
or U36556 (N_36556,N_36346,N_36355);
nor U36557 (N_36557,N_36454,N_36257);
nor U36558 (N_36558,N_36465,N_36432);
nand U36559 (N_36559,N_36336,N_36337);
nand U36560 (N_36560,N_36388,N_36296);
and U36561 (N_36561,N_36442,N_36394);
or U36562 (N_36562,N_36279,N_36295);
or U36563 (N_36563,N_36314,N_36414);
xor U36564 (N_36564,N_36380,N_36343);
xnor U36565 (N_36565,N_36290,N_36448);
and U36566 (N_36566,N_36265,N_36421);
nor U36567 (N_36567,N_36477,N_36406);
nand U36568 (N_36568,N_36459,N_36496);
or U36569 (N_36569,N_36423,N_36354);
nor U36570 (N_36570,N_36420,N_36310);
nand U36571 (N_36571,N_36289,N_36324);
nor U36572 (N_36572,N_36462,N_36404);
xnor U36573 (N_36573,N_36428,N_36347);
xor U36574 (N_36574,N_36263,N_36435);
xnor U36575 (N_36575,N_36393,N_36269);
and U36576 (N_36576,N_36464,N_36274);
and U36577 (N_36577,N_36306,N_36437);
nor U36578 (N_36578,N_36342,N_36424);
xnor U36579 (N_36579,N_36366,N_36395);
nor U36580 (N_36580,N_36449,N_36278);
and U36581 (N_36581,N_36383,N_36444);
nand U36582 (N_36582,N_36320,N_36332);
and U36583 (N_36583,N_36376,N_36390);
nor U36584 (N_36584,N_36369,N_36319);
or U36585 (N_36585,N_36485,N_36286);
xnor U36586 (N_36586,N_36252,N_36418);
or U36587 (N_36587,N_36297,N_36302);
and U36588 (N_36588,N_36417,N_36470);
nand U36589 (N_36589,N_36350,N_36445);
nand U36590 (N_36590,N_36431,N_36455);
nand U36591 (N_36591,N_36371,N_36281);
and U36592 (N_36592,N_36311,N_36386);
and U36593 (N_36593,N_36382,N_36481);
and U36594 (N_36594,N_36251,N_36486);
xor U36595 (N_36595,N_36427,N_36498);
nor U36596 (N_36596,N_36400,N_36363);
nand U36597 (N_36597,N_36321,N_36357);
xor U36598 (N_36598,N_36475,N_36254);
nor U36599 (N_36599,N_36401,N_36294);
xnor U36600 (N_36600,N_36453,N_36377);
or U36601 (N_36601,N_36426,N_36468);
or U36602 (N_36602,N_36474,N_36288);
xor U36603 (N_36603,N_36264,N_36353);
xnor U36604 (N_36604,N_36333,N_36389);
nor U36605 (N_36605,N_36499,N_36304);
or U36606 (N_36606,N_36303,N_36266);
nor U36607 (N_36607,N_36270,N_36413);
and U36608 (N_36608,N_36348,N_36255);
nand U36609 (N_36609,N_36299,N_36285);
nor U36610 (N_36610,N_36488,N_36491);
nor U36611 (N_36611,N_36301,N_36419);
xnor U36612 (N_36612,N_36415,N_36370);
and U36613 (N_36613,N_36364,N_36396);
nand U36614 (N_36614,N_36494,N_36456);
nor U36615 (N_36615,N_36457,N_36334);
nand U36616 (N_36616,N_36340,N_36344);
nand U36617 (N_36617,N_36309,N_36312);
or U36618 (N_36618,N_36250,N_36273);
nor U36619 (N_36619,N_36490,N_36378);
or U36620 (N_36620,N_36351,N_36368);
or U36621 (N_36621,N_36267,N_36329);
nand U36622 (N_36622,N_36450,N_36261);
or U36623 (N_36623,N_36466,N_36397);
nand U36624 (N_36624,N_36434,N_36280);
or U36625 (N_36625,N_36434,N_36361);
nor U36626 (N_36626,N_36477,N_36403);
and U36627 (N_36627,N_36468,N_36288);
and U36628 (N_36628,N_36497,N_36362);
nor U36629 (N_36629,N_36481,N_36455);
nand U36630 (N_36630,N_36312,N_36258);
nand U36631 (N_36631,N_36302,N_36447);
or U36632 (N_36632,N_36349,N_36450);
and U36633 (N_36633,N_36376,N_36263);
nor U36634 (N_36634,N_36472,N_36367);
or U36635 (N_36635,N_36327,N_36474);
or U36636 (N_36636,N_36460,N_36380);
or U36637 (N_36637,N_36458,N_36498);
or U36638 (N_36638,N_36448,N_36412);
nand U36639 (N_36639,N_36281,N_36261);
or U36640 (N_36640,N_36393,N_36392);
and U36641 (N_36641,N_36344,N_36493);
or U36642 (N_36642,N_36331,N_36271);
xnor U36643 (N_36643,N_36287,N_36378);
xnor U36644 (N_36644,N_36304,N_36328);
nand U36645 (N_36645,N_36366,N_36363);
nand U36646 (N_36646,N_36492,N_36423);
xnor U36647 (N_36647,N_36418,N_36310);
or U36648 (N_36648,N_36259,N_36357);
and U36649 (N_36649,N_36449,N_36422);
and U36650 (N_36650,N_36415,N_36349);
and U36651 (N_36651,N_36355,N_36415);
and U36652 (N_36652,N_36442,N_36450);
or U36653 (N_36653,N_36264,N_36349);
xnor U36654 (N_36654,N_36352,N_36374);
xor U36655 (N_36655,N_36466,N_36267);
and U36656 (N_36656,N_36262,N_36306);
or U36657 (N_36657,N_36374,N_36265);
nor U36658 (N_36658,N_36294,N_36372);
xor U36659 (N_36659,N_36383,N_36451);
nand U36660 (N_36660,N_36386,N_36377);
xor U36661 (N_36661,N_36490,N_36427);
or U36662 (N_36662,N_36254,N_36298);
nand U36663 (N_36663,N_36331,N_36308);
nand U36664 (N_36664,N_36458,N_36499);
nand U36665 (N_36665,N_36446,N_36440);
nor U36666 (N_36666,N_36378,N_36423);
nand U36667 (N_36667,N_36411,N_36296);
or U36668 (N_36668,N_36385,N_36288);
and U36669 (N_36669,N_36304,N_36479);
and U36670 (N_36670,N_36453,N_36375);
nand U36671 (N_36671,N_36482,N_36412);
nor U36672 (N_36672,N_36338,N_36484);
nor U36673 (N_36673,N_36415,N_36296);
xnor U36674 (N_36674,N_36416,N_36382);
or U36675 (N_36675,N_36406,N_36351);
or U36676 (N_36676,N_36427,N_36319);
xor U36677 (N_36677,N_36258,N_36301);
or U36678 (N_36678,N_36290,N_36458);
xnor U36679 (N_36679,N_36386,N_36454);
xnor U36680 (N_36680,N_36433,N_36432);
nand U36681 (N_36681,N_36420,N_36255);
xor U36682 (N_36682,N_36380,N_36367);
nand U36683 (N_36683,N_36428,N_36407);
nand U36684 (N_36684,N_36253,N_36320);
nor U36685 (N_36685,N_36285,N_36301);
nand U36686 (N_36686,N_36353,N_36437);
nor U36687 (N_36687,N_36270,N_36449);
xnor U36688 (N_36688,N_36492,N_36315);
or U36689 (N_36689,N_36433,N_36422);
nor U36690 (N_36690,N_36296,N_36458);
xor U36691 (N_36691,N_36361,N_36322);
nand U36692 (N_36692,N_36299,N_36273);
and U36693 (N_36693,N_36350,N_36373);
and U36694 (N_36694,N_36335,N_36458);
nor U36695 (N_36695,N_36349,N_36411);
or U36696 (N_36696,N_36498,N_36338);
xor U36697 (N_36697,N_36450,N_36437);
nor U36698 (N_36698,N_36383,N_36312);
nor U36699 (N_36699,N_36394,N_36334);
or U36700 (N_36700,N_36316,N_36487);
xor U36701 (N_36701,N_36283,N_36361);
nand U36702 (N_36702,N_36286,N_36463);
and U36703 (N_36703,N_36465,N_36347);
or U36704 (N_36704,N_36331,N_36366);
or U36705 (N_36705,N_36266,N_36251);
xnor U36706 (N_36706,N_36294,N_36489);
and U36707 (N_36707,N_36369,N_36264);
xnor U36708 (N_36708,N_36308,N_36438);
xor U36709 (N_36709,N_36403,N_36326);
nand U36710 (N_36710,N_36295,N_36285);
nor U36711 (N_36711,N_36413,N_36407);
nor U36712 (N_36712,N_36369,N_36353);
or U36713 (N_36713,N_36401,N_36450);
or U36714 (N_36714,N_36273,N_36308);
and U36715 (N_36715,N_36292,N_36287);
or U36716 (N_36716,N_36405,N_36290);
nor U36717 (N_36717,N_36479,N_36252);
nand U36718 (N_36718,N_36395,N_36435);
or U36719 (N_36719,N_36457,N_36347);
or U36720 (N_36720,N_36359,N_36306);
or U36721 (N_36721,N_36311,N_36257);
xor U36722 (N_36722,N_36443,N_36268);
xnor U36723 (N_36723,N_36406,N_36472);
nand U36724 (N_36724,N_36395,N_36388);
or U36725 (N_36725,N_36417,N_36430);
or U36726 (N_36726,N_36438,N_36430);
and U36727 (N_36727,N_36352,N_36443);
xnor U36728 (N_36728,N_36377,N_36435);
or U36729 (N_36729,N_36330,N_36341);
nor U36730 (N_36730,N_36316,N_36287);
nand U36731 (N_36731,N_36384,N_36252);
nand U36732 (N_36732,N_36497,N_36265);
xor U36733 (N_36733,N_36394,N_36477);
nand U36734 (N_36734,N_36348,N_36441);
and U36735 (N_36735,N_36319,N_36398);
xor U36736 (N_36736,N_36454,N_36463);
xor U36737 (N_36737,N_36495,N_36422);
and U36738 (N_36738,N_36349,N_36281);
xor U36739 (N_36739,N_36490,N_36393);
nand U36740 (N_36740,N_36293,N_36258);
nand U36741 (N_36741,N_36477,N_36400);
and U36742 (N_36742,N_36276,N_36332);
nand U36743 (N_36743,N_36495,N_36365);
nand U36744 (N_36744,N_36496,N_36430);
or U36745 (N_36745,N_36457,N_36397);
xnor U36746 (N_36746,N_36398,N_36294);
nor U36747 (N_36747,N_36423,N_36388);
nor U36748 (N_36748,N_36466,N_36409);
nor U36749 (N_36749,N_36312,N_36359);
nor U36750 (N_36750,N_36599,N_36502);
xnor U36751 (N_36751,N_36708,N_36731);
xor U36752 (N_36752,N_36650,N_36537);
and U36753 (N_36753,N_36557,N_36668);
and U36754 (N_36754,N_36654,N_36649);
xor U36755 (N_36755,N_36718,N_36694);
or U36756 (N_36756,N_36633,N_36715);
nand U36757 (N_36757,N_36723,N_36620);
or U36758 (N_36758,N_36680,N_36521);
or U36759 (N_36759,N_36690,N_36671);
xor U36760 (N_36760,N_36747,N_36735);
nand U36761 (N_36761,N_36583,N_36629);
nand U36762 (N_36762,N_36711,N_36721);
nor U36763 (N_36763,N_36677,N_36693);
or U36764 (N_36764,N_36553,N_36566);
nand U36765 (N_36765,N_36508,N_36555);
nor U36766 (N_36766,N_36554,N_36528);
and U36767 (N_36767,N_36641,N_36706);
xnor U36768 (N_36768,N_36591,N_36511);
nand U36769 (N_36769,N_36638,N_36709);
nor U36770 (N_36770,N_36504,N_36613);
nand U36771 (N_36771,N_36541,N_36597);
or U36772 (N_36772,N_36734,N_36743);
nor U36773 (N_36773,N_36701,N_36678);
or U36774 (N_36774,N_36660,N_36667);
nand U36775 (N_36775,N_36742,N_36600);
xnor U36776 (N_36776,N_36670,N_36609);
nand U36777 (N_36777,N_36643,N_36653);
or U36778 (N_36778,N_36601,N_36741);
and U36779 (N_36779,N_36563,N_36648);
xnor U36780 (N_36780,N_36740,N_36532);
nor U36781 (N_36781,N_36595,N_36669);
and U36782 (N_36782,N_36713,N_36561);
or U36783 (N_36783,N_36558,N_36500);
nor U36784 (N_36784,N_36515,N_36574);
or U36785 (N_36785,N_36501,N_36594);
and U36786 (N_36786,N_36642,N_36682);
xnor U36787 (N_36787,N_36540,N_36729);
and U36788 (N_36788,N_36587,N_36637);
and U36789 (N_36789,N_36738,N_36509);
nor U36790 (N_36790,N_36626,N_36749);
and U36791 (N_36791,N_36505,N_36610);
xnor U36792 (N_36792,N_36533,N_36665);
xnor U36793 (N_36793,N_36569,N_36512);
nand U36794 (N_36794,N_36549,N_36631);
nor U36795 (N_36795,N_36632,N_36546);
nor U36796 (N_36796,N_36535,N_36730);
nand U36797 (N_36797,N_36726,N_36679);
and U36798 (N_36798,N_36656,N_36581);
or U36799 (N_36799,N_36607,N_36618);
nand U36800 (N_36800,N_36615,N_36662);
nor U36801 (N_36801,N_36526,N_36586);
nor U36802 (N_36802,N_36733,N_36651);
nand U36803 (N_36803,N_36547,N_36705);
nand U36804 (N_36804,N_36534,N_36603);
nand U36805 (N_36805,N_36674,N_36612);
nor U36806 (N_36806,N_36699,N_36529);
nor U36807 (N_36807,N_36640,N_36722);
and U36808 (N_36808,N_36619,N_36578);
nor U36809 (N_36809,N_36565,N_36559);
or U36810 (N_36810,N_36687,N_36624);
xnor U36811 (N_36811,N_36698,N_36657);
or U36812 (N_36812,N_36530,N_36645);
or U36813 (N_36813,N_36545,N_36516);
or U36814 (N_36814,N_36696,N_36703);
or U36815 (N_36815,N_36577,N_36630);
nor U36816 (N_36816,N_36556,N_36514);
or U36817 (N_36817,N_36544,N_36623);
or U36818 (N_36818,N_36655,N_36606);
xnor U36819 (N_36819,N_36673,N_36621);
and U36820 (N_36820,N_36727,N_36634);
nor U36821 (N_36821,N_36683,N_36564);
nor U36822 (N_36822,N_36524,N_36745);
or U36823 (N_36823,N_36605,N_36614);
nor U36824 (N_36824,N_36608,N_36695);
and U36825 (N_36825,N_36716,N_36689);
and U36826 (N_36826,N_36604,N_36571);
or U36827 (N_36827,N_36746,N_36568);
xor U36828 (N_36828,N_36658,N_36617);
nor U36829 (N_36829,N_36732,N_36552);
nor U36830 (N_36830,N_36523,N_36580);
nand U36831 (N_36831,N_36704,N_36639);
xnor U36832 (N_36832,N_36710,N_36518);
nor U36833 (N_36833,N_36739,N_36550);
nor U36834 (N_36834,N_36560,N_36588);
nor U36835 (N_36835,N_36525,N_36531);
xor U36836 (N_36836,N_36592,N_36576);
and U36837 (N_36837,N_36539,N_36625);
and U36838 (N_36838,N_36507,N_36536);
nand U36839 (N_36839,N_36717,N_36644);
and U36840 (N_36840,N_36562,N_36622);
nand U36841 (N_36841,N_36519,N_36652);
xnor U36842 (N_36842,N_36712,N_36685);
xnor U36843 (N_36843,N_36702,N_36575);
nor U36844 (N_36844,N_36596,N_36725);
or U36845 (N_36845,N_36582,N_36548);
nand U36846 (N_36846,N_36513,N_36672);
nor U36847 (N_36847,N_36724,N_36748);
nand U36848 (N_36848,N_36567,N_36589);
xor U36849 (N_36849,N_36602,N_36666);
nor U36850 (N_36850,N_36659,N_36590);
nand U36851 (N_36851,N_36520,N_36684);
and U36852 (N_36852,N_36636,N_36635);
and U36853 (N_36853,N_36551,N_36538);
and U36854 (N_36854,N_36686,N_36664);
xnor U36855 (N_36855,N_36700,N_36707);
xnor U36856 (N_36856,N_36573,N_36681);
nor U36857 (N_36857,N_36506,N_36628);
nor U36858 (N_36858,N_36675,N_36598);
and U36859 (N_36859,N_36503,N_36527);
xor U36860 (N_36860,N_36691,N_36661);
nor U36861 (N_36861,N_36593,N_36720);
nor U36862 (N_36862,N_36744,N_36663);
nor U36863 (N_36863,N_36572,N_36579);
and U36864 (N_36864,N_36736,N_36616);
xor U36865 (N_36865,N_36688,N_36737);
nand U36866 (N_36866,N_36611,N_36692);
nor U36867 (N_36867,N_36585,N_36570);
and U36868 (N_36868,N_36627,N_36728);
nand U36869 (N_36869,N_36522,N_36697);
nand U36870 (N_36870,N_36542,N_36647);
nand U36871 (N_36871,N_36543,N_36517);
and U36872 (N_36872,N_36714,N_36676);
xor U36873 (N_36873,N_36510,N_36719);
nor U36874 (N_36874,N_36646,N_36584);
nand U36875 (N_36875,N_36512,N_36678);
nand U36876 (N_36876,N_36703,N_36649);
nor U36877 (N_36877,N_36719,N_36511);
or U36878 (N_36878,N_36633,N_36740);
or U36879 (N_36879,N_36508,N_36685);
nand U36880 (N_36880,N_36704,N_36576);
nand U36881 (N_36881,N_36677,N_36708);
and U36882 (N_36882,N_36565,N_36546);
or U36883 (N_36883,N_36720,N_36508);
nor U36884 (N_36884,N_36659,N_36512);
nor U36885 (N_36885,N_36654,N_36648);
or U36886 (N_36886,N_36564,N_36581);
nor U36887 (N_36887,N_36555,N_36697);
or U36888 (N_36888,N_36718,N_36567);
nor U36889 (N_36889,N_36562,N_36631);
nand U36890 (N_36890,N_36610,N_36568);
xnor U36891 (N_36891,N_36612,N_36695);
or U36892 (N_36892,N_36607,N_36506);
or U36893 (N_36893,N_36745,N_36608);
nand U36894 (N_36894,N_36730,N_36614);
and U36895 (N_36895,N_36720,N_36674);
or U36896 (N_36896,N_36686,N_36671);
or U36897 (N_36897,N_36554,N_36622);
or U36898 (N_36898,N_36628,N_36565);
nor U36899 (N_36899,N_36656,N_36749);
nand U36900 (N_36900,N_36637,N_36615);
nor U36901 (N_36901,N_36564,N_36746);
or U36902 (N_36902,N_36713,N_36738);
or U36903 (N_36903,N_36721,N_36618);
or U36904 (N_36904,N_36678,N_36607);
and U36905 (N_36905,N_36547,N_36595);
nor U36906 (N_36906,N_36731,N_36551);
nor U36907 (N_36907,N_36681,N_36584);
xnor U36908 (N_36908,N_36571,N_36643);
and U36909 (N_36909,N_36723,N_36643);
xor U36910 (N_36910,N_36590,N_36680);
xor U36911 (N_36911,N_36594,N_36572);
xor U36912 (N_36912,N_36511,N_36607);
and U36913 (N_36913,N_36531,N_36539);
nor U36914 (N_36914,N_36564,N_36695);
nor U36915 (N_36915,N_36689,N_36575);
or U36916 (N_36916,N_36723,N_36682);
nor U36917 (N_36917,N_36705,N_36697);
and U36918 (N_36918,N_36584,N_36643);
and U36919 (N_36919,N_36513,N_36600);
and U36920 (N_36920,N_36594,N_36578);
and U36921 (N_36921,N_36720,N_36571);
or U36922 (N_36922,N_36722,N_36623);
or U36923 (N_36923,N_36711,N_36661);
xor U36924 (N_36924,N_36668,N_36659);
xor U36925 (N_36925,N_36598,N_36510);
xnor U36926 (N_36926,N_36736,N_36749);
nor U36927 (N_36927,N_36571,N_36733);
and U36928 (N_36928,N_36523,N_36656);
xor U36929 (N_36929,N_36717,N_36626);
nand U36930 (N_36930,N_36726,N_36520);
xnor U36931 (N_36931,N_36716,N_36508);
nand U36932 (N_36932,N_36683,N_36558);
nor U36933 (N_36933,N_36577,N_36593);
and U36934 (N_36934,N_36728,N_36629);
xor U36935 (N_36935,N_36568,N_36714);
nor U36936 (N_36936,N_36544,N_36587);
xnor U36937 (N_36937,N_36722,N_36668);
xor U36938 (N_36938,N_36719,N_36621);
nor U36939 (N_36939,N_36710,N_36501);
nand U36940 (N_36940,N_36706,N_36719);
nand U36941 (N_36941,N_36604,N_36627);
xor U36942 (N_36942,N_36722,N_36657);
nor U36943 (N_36943,N_36663,N_36628);
nor U36944 (N_36944,N_36697,N_36714);
xnor U36945 (N_36945,N_36564,N_36658);
or U36946 (N_36946,N_36500,N_36632);
nor U36947 (N_36947,N_36718,N_36661);
nor U36948 (N_36948,N_36666,N_36636);
and U36949 (N_36949,N_36706,N_36609);
xor U36950 (N_36950,N_36658,N_36649);
nor U36951 (N_36951,N_36538,N_36714);
xnor U36952 (N_36952,N_36709,N_36644);
xor U36953 (N_36953,N_36505,N_36548);
and U36954 (N_36954,N_36538,N_36674);
or U36955 (N_36955,N_36629,N_36592);
or U36956 (N_36956,N_36632,N_36557);
nor U36957 (N_36957,N_36733,N_36736);
nand U36958 (N_36958,N_36550,N_36697);
and U36959 (N_36959,N_36612,N_36719);
xnor U36960 (N_36960,N_36696,N_36552);
or U36961 (N_36961,N_36561,N_36708);
or U36962 (N_36962,N_36533,N_36737);
xnor U36963 (N_36963,N_36708,N_36564);
xnor U36964 (N_36964,N_36542,N_36539);
nor U36965 (N_36965,N_36591,N_36560);
xnor U36966 (N_36966,N_36567,N_36749);
xor U36967 (N_36967,N_36521,N_36571);
and U36968 (N_36968,N_36744,N_36658);
xnor U36969 (N_36969,N_36595,N_36675);
nor U36970 (N_36970,N_36656,N_36670);
or U36971 (N_36971,N_36737,N_36535);
and U36972 (N_36972,N_36535,N_36629);
xor U36973 (N_36973,N_36680,N_36633);
and U36974 (N_36974,N_36650,N_36643);
and U36975 (N_36975,N_36519,N_36593);
nor U36976 (N_36976,N_36627,N_36538);
xor U36977 (N_36977,N_36565,N_36631);
or U36978 (N_36978,N_36669,N_36529);
nand U36979 (N_36979,N_36579,N_36705);
nand U36980 (N_36980,N_36557,N_36655);
xnor U36981 (N_36981,N_36638,N_36532);
nand U36982 (N_36982,N_36652,N_36687);
xor U36983 (N_36983,N_36608,N_36694);
nor U36984 (N_36984,N_36737,N_36698);
xnor U36985 (N_36985,N_36569,N_36685);
nor U36986 (N_36986,N_36648,N_36531);
xnor U36987 (N_36987,N_36698,N_36529);
nand U36988 (N_36988,N_36742,N_36718);
nor U36989 (N_36989,N_36602,N_36569);
nand U36990 (N_36990,N_36588,N_36744);
or U36991 (N_36991,N_36589,N_36659);
or U36992 (N_36992,N_36629,N_36748);
nand U36993 (N_36993,N_36508,N_36529);
or U36994 (N_36994,N_36668,N_36609);
nor U36995 (N_36995,N_36516,N_36694);
xor U36996 (N_36996,N_36585,N_36711);
xnor U36997 (N_36997,N_36537,N_36519);
or U36998 (N_36998,N_36653,N_36588);
nand U36999 (N_36999,N_36739,N_36677);
nor U37000 (N_37000,N_36922,N_36838);
or U37001 (N_37001,N_36908,N_36924);
nand U37002 (N_37002,N_36939,N_36974);
nand U37003 (N_37003,N_36828,N_36981);
nand U37004 (N_37004,N_36894,N_36871);
nor U37005 (N_37005,N_36841,N_36909);
and U37006 (N_37006,N_36952,N_36778);
or U37007 (N_37007,N_36886,N_36879);
nor U37008 (N_37008,N_36823,N_36809);
nand U37009 (N_37009,N_36784,N_36902);
or U37010 (N_37010,N_36934,N_36979);
xnor U37011 (N_37011,N_36956,N_36808);
xor U37012 (N_37012,N_36799,N_36750);
or U37013 (N_37013,N_36822,N_36966);
nor U37014 (N_37014,N_36954,N_36985);
nand U37015 (N_37015,N_36818,N_36906);
nand U37016 (N_37016,N_36949,N_36824);
nor U37017 (N_37017,N_36768,N_36868);
or U37018 (N_37018,N_36753,N_36834);
and U37019 (N_37019,N_36978,N_36913);
nor U37020 (N_37020,N_36904,N_36819);
nor U37021 (N_37021,N_36864,N_36811);
nand U37022 (N_37022,N_36788,N_36926);
xor U37023 (N_37023,N_36772,N_36994);
xnor U37024 (N_37024,N_36776,N_36989);
nor U37025 (N_37025,N_36987,N_36877);
and U37026 (N_37026,N_36795,N_36796);
nand U37027 (N_37027,N_36802,N_36854);
nand U37028 (N_37028,N_36999,N_36842);
or U37029 (N_37029,N_36980,N_36829);
xnor U37030 (N_37030,N_36907,N_36763);
or U37031 (N_37031,N_36805,N_36898);
and U37032 (N_37032,N_36767,N_36945);
and U37033 (N_37033,N_36967,N_36972);
nor U37034 (N_37034,N_36917,N_36831);
nor U37035 (N_37035,N_36865,N_36928);
and U37036 (N_37036,N_36844,N_36775);
nor U37037 (N_37037,N_36959,N_36996);
and U37038 (N_37038,N_36903,N_36777);
or U37039 (N_37039,N_36889,N_36845);
and U37040 (N_37040,N_36911,N_36754);
or U37041 (N_37041,N_36878,N_36849);
or U37042 (N_37042,N_36935,N_36881);
nor U37043 (N_37043,N_36783,N_36851);
xor U37044 (N_37044,N_36901,N_36764);
or U37045 (N_37045,N_36948,N_36986);
nand U37046 (N_37046,N_36997,N_36797);
and U37047 (N_37047,N_36860,N_36875);
and U37048 (N_37048,N_36968,N_36899);
and U37049 (N_37049,N_36887,N_36821);
nand U37050 (N_37050,N_36883,N_36755);
or U37051 (N_37051,N_36847,N_36983);
nand U37052 (N_37052,N_36803,N_36843);
nand U37053 (N_37053,N_36820,N_36814);
and U37054 (N_37054,N_36940,N_36957);
xnor U37055 (N_37055,N_36975,N_36798);
xnor U37056 (N_37056,N_36794,N_36888);
xor U37057 (N_37057,N_36977,N_36988);
and U37058 (N_37058,N_36905,N_36870);
nor U37059 (N_37059,N_36893,N_36992);
and U37060 (N_37060,N_36792,N_36833);
nor U37061 (N_37061,N_36846,N_36789);
and U37062 (N_37062,N_36770,N_36976);
xnor U37063 (N_37063,N_36855,N_36910);
xor U37064 (N_37064,N_36852,N_36766);
and U37065 (N_37065,N_36955,N_36816);
or U37066 (N_37066,N_36857,N_36812);
and U37067 (N_37067,N_36884,N_36961);
nand U37068 (N_37068,N_36859,N_36937);
or U37069 (N_37069,N_36872,N_36861);
nor U37070 (N_37070,N_36963,N_36781);
and U37071 (N_37071,N_36929,N_36752);
nor U37072 (N_37072,N_36951,N_36890);
and U37073 (N_37073,N_36895,N_36862);
and U37074 (N_37074,N_36953,N_36962);
nand U37075 (N_37075,N_36780,N_36827);
xnor U37076 (N_37076,N_36826,N_36931);
or U37077 (N_37077,N_36815,N_36982);
nor U37078 (N_37078,N_36970,N_36869);
nand U37079 (N_37079,N_36891,N_36876);
and U37080 (N_37080,N_36813,N_36944);
or U37081 (N_37081,N_36771,N_36810);
xnor U37082 (N_37082,N_36840,N_36760);
or U37083 (N_37083,N_36915,N_36925);
xor U37084 (N_37084,N_36995,N_36927);
nor U37085 (N_37085,N_36950,N_36836);
nor U37086 (N_37086,N_36946,N_36920);
nor U37087 (N_37087,N_36793,N_36762);
and U37088 (N_37088,N_36782,N_36751);
or U37089 (N_37089,N_36880,N_36765);
xor U37090 (N_37090,N_36964,N_36758);
or U37091 (N_37091,N_36853,N_36790);
nor U37092 (N_37092,N_36832,N_36807);
or U37093 (N_37093,N_36998,N_36761);
nand U37094 (N_37094,N_36900,N_36759);
xor U37095 (N_37095,N_36787,N_36856);
nor U37096 (N_37096,N_36791,N_36801);
xnor U37097 (N_37097,N_36779,N_36896);
or U37098 (N_37098,N_36993,N_36984);
xor U37099 (N_37099,N_36947,N_36941);
nand U37100 (N_37100,N_36932,N_36837);
nor U37101 (N_37101,N_36874,N_36973);
nand U37102 (N_37102,N_36971,N_36757);
and U37103 (N_37103,N_36866,N_36897);
and U37104 (N_37104,N_36942,N_36858);
or U37105 (N_37105,N_36804,N_36923);
nand U37106 (N_37106,N_36930,N_36863);
nand U37107 (N_37107,N_36965,N_36806);
and U37108 (N_37108,N_36921,N_36785);
xor U37109 (N_37109,N_36918,N_36916);
nor U37110 (N_37110,N_36933,N_36943);
xnor U37111 (N_37111,N_36867,N_36914);
nand U37112 (N_37112,N_36848,N_36839);
and U37113 (N_37113,N_36958,N_36817);
nor U37114 (N_37114,N_36969,N_36825);
xnor U37115 (N_37115,N_36885,N_36835);
and U37116 (N_37116,N_36873,N_36990);
xor U37117 (N_37117,N_36960,N_36830);
nor U37118 (N_37118,N_36773,N_36774);
and U37119 (N_37119,N_36882,N_36800);
and U37120 (N_37120,N_36850,N_36912);
and U37121 (N_37121,N_36991,N_36786);
or U37122 (N_37122,N_36938,N_36892);
nor U37123 (N_37123,N_36769,N_36919);
and U37124 (N_37124,N_36936,N_36756);
nand U37125 (N_37125,N_36854,N_36874);
and U37126 (N_37126,N_36792,N_36827);
nand U37127 (N_37127,N_36812,N_36908);
xor U37128 (N_37128,N_36907,N_36995);
xor U37129 (N_37129,N_36943,N_36834);
xor U37130 (N_37130,N_36803,N_36815);
and U37131 (N_37131,N_36838,N_36966);
xnor U37132 (N_37132,N_36989,N_36969);
nand U37133 (N_37133,N_36870,N_36791);
xnor U37134 (N_37134,N_36814,N_36962);
and U37135 (N_37135,N_36882,N_36941);
and U37136 (N_37136,N_36780,N_36930);
nor U37137 (N_37137,N_36883,N_36956);
or U37138 (N_37138,N_36963,N_36976);
xnor U37139 (N_37139,N_36866,N_36796);
nand U37140 (N_37140,N_36756,N_36834);
xor U37141 (N_37141,N_36800,N_36804);
or U37142 (N_37142,N_36880,N_36786);
nor U37143 (N_37143,N_36976,N_36878);
nand U37144 (N_37144,N_36990,N_36948);
or U37145 (N_37145,N_36903,N_36775);
nand U37146 (N_37146,N_36946,N_36907);
and U37147 (N_37147,N_36969,N_36974);
nor U37148 (N_37148,N_36947,N_36901);
xnor U37149 (N_37149,N_36886,N_36828);
or U37150 (N_37150,N_36816,N_36960);
or U37151 (N_37151,N_36963,N_36865);
or U37152 (N_37152,N_36995,N_36935);
xor U37153 (N_37153,N_36754,N_36927);
nand U37154 (N_37154,N_36865,N_36982);
and U37155 (N_37155,N_36805,N_36789);
nand U37156 (N_37156,N_36851,N_36812);
nor U37157 (N_37157,N_36964,N_36759);
or U37158 (N_37158,N_36886,N_36776);
nand U37159 (N_37159,N_36824,N_36754);
nor U37160 (N_37160,N_36929,N_36798);
and U37161 (N_37161,N_36784,N_36934);
xnor U37162 (N_37162,N_36950,N_36928);
nor U37163 (N_37163,N_36861,N_36857);
nand U37164 (N_37164,N_36846,N_36923);
or U37165 (N_37165,N_36895,N_36989);
xor U37166 (N_37166,N_36849,N_36940);
nor U37167 (N_37167,N_36924,N_36792);
xnor U37168 (N_37168,N_36805,N_36803);
xor U37169 (N_37169,N_36988,N_36995);
and U37170 (N_37170,N_36999,N_36822);
xnor U37171 (N_37171,N_36994,N_36914);
and U37172 (N_37172,N_36856,N_36983);
nor U37173 (N_37173,N_36788,N_36847);
or U37174 (N_37174,N_36871,N_36889);
xnor U37175 (N_37175,N_36814,N_36811);
nand U37176 (N_37176,N_36771,N_36844);
nand U37177 (N_37177,N_36905,N_36970);
nand U37178 (N_37178,N_36908,N_36803);
nand U37179 (N_37179,N_36937,N_36967);
and U37180 (N_37180,N_36865,N_36976);
nor U37181 (N_37181,N_36931,N_36762);
and U37182 (N_37182,N_36920,N_36988);
xnor U37183 (N_37183,N_36950,N_36940);
nor U37184 (N_37184,N_36763,N_36767);
and U37185 (N_37185,N_36862,N_36952);
xor U37186 (N_37186,N_36781,N_36755);
xor U37187 (N_37187,N_36880,N_36991);
xnor U37188 (N_37188,N_36804,N_36972);
and U37189 (N_37189,N_36904,N_36962);
xor U37190 (N_37190,N_36796,N_36938);
nor U37191 (N_37191,N_36789,N_36921);
xnor U37192 (N_37192,N_36879,N_36817);
xnor U37193 (N_37193,N_36961,N_36933);
and U37194 (N_37194,N_36970,N_36851);
and U37195 (N_37195,N_36987,N_36891);
xnor U37196 (N_37196,N_36810,N_36773);
and U37197 (N_37197,N_36870,N_36990);
and U37198 (N_37198,N_36827,N_36948);
xor U37199 (N_37199,N_36982,N_36850);
nand U37200 (N_37200,N_36830,N_36946);
xor U37201 (N_37201,N_36883,N_36902);
nor U37202 (N_37202,N_36996,N_36856);
nor U37203 (N_37203,N_36964,N_36880);
and U37204 (N_37204,N_36789,N_36911);
or U37205 (N_37205,N_36994,N_36867);
or U37206 (N_37206,N_36787,N_36973);
or U37207 (N_37207,N_36769,N_36766);
and U37208 (N_37208,N_36901,N_36980);
nor U37209 (N_37209,N_36946,N_36811);
or U37210 (N_37210,N_36772,N_36976);
or U37211 (N_37211,N_36961,N_36820);
nand U37212 (N_37212,N_36939,N_36870);
nor U37213 (N_37213,N_36773,N_36912);
nand U37214 (N_37214,N_36852,N_36805);
or U37215 (N_37215,N_36931,N_36880);
xor U37216 (N_37216,N_36847,N_36962);
and U37217 (N_37217,N_36986,N_36826);
or U37218 (N_37218,N_36864,N_36862);
and U37219 (N_37219,N_36992,N_36979);
or U37220 (N_37220,N_36828,N_36824);
nand U37221 (N_37221,N_36835,N_36800);
or U37222 (N_37222,N_36803,N_36790);
and U37223 (N_37223,N_36864,N_36833);
or U37224 (N_37224,N_36770,N_36979);
nor U37225 (N_37225,N_36989,N_36771);
or U37226 (N_37226,N_36838,N_36794);
and U37227 (N_37227,N_36973,N_36795);
nor U37228 (N_37228,N_36766,N_36889);
and U37229 (N_37229,N_36849,N_36819);
nor U37230 (N_37230,N_36803,N_36800);
and U37231 (N_37231,N_36980,N_36792);
nand U37232 (N_37232,N_36808,N_36895);
and U37233 (N_37233,N_36974,N_36981);
and U37234 (N_37234,N_36849,N_36836);
nor U37235 (N_37235,N_36914,N_36815);
xor U37236 (N_37236,N_36927,N_36948);
and U37237 (N_37237,N_36808,N_36976);
nor U37238 (N_37238,N_36969,N_36809);
nand U37239 (N_37239,N_36913,N_36908);
xnor U37240 (N_37240,N_36853,N_36890);
or U37241 (N_37241,N_36940,N_36935);
or U37242 (N_37242,N_36862,N_36756);
nor U37243 (N_37243,N_36817,N_36786);
nor U37244 (N_37244,N_36905,N_36940);
nand U37245 (N_37245,N_36895,N_36800);
nand U37246 (N_37246,N_36929,N_36852);
nor U37247 (N_37247,N_36864,N_36838);
or U37248 (N_37248,N_36755,N_36925);
or U37249 (N_37249,N_36917,N_36825);
nand U37250 (N_37250,N_37233,N_37218);
or U37251 (N_37251,N_37035,N_37051);
or U37252 (N_37252,N_37104,N_37075);
xnor U37253 (N_37253,N_37193,N_37129);
xor U37254 (N_37254,N_37067,N_37096);
xnor U37255 (N_37255,N_37020,N_37112);
nor U37256 (N_37256,N_37128,N_37071);
or U37257 (N_37257,N_37072,N_37231);
nand U37258 (N_37258,N_37153,N_37102);
or U37259 (N_37259,N_37182,N_37175);
and U37260 (N_37260,N_37042,N_37215);
or U37261 (N_37261,N_37239,N_37200);
and U37262 (N_37262,N_37119,N_37041);
or U37263 (N_37263,N_37143,N_37230);
xnor U37264 (N_37264,N_37079,N_37132);
nor U37265 (N_37265,N_37174,N_37146);
xnor U37266 (N_37266,N_37049,N_37190);
and U37267 (N_37267,N_37225,N_37066);
and U37268 (N_37268,N_37030,N_37220);
and U37269 (N_37269,N_37115,N_37198);
nand U37270 (N_37270,N_37163,N_37016);
or U37271 (N_37271,N_37179,N_37188);
xnor U37272 (N_37272,N_37080,N_37135);
nor U37273 (N_37273,N_37053,N_37183);
xor U37274 (N_37274,N_37249,N_37002);
and U37275 (N_37275,N_37158,N_37144);
and U37276 (N_37276,N_37162,N_37147);
xor U37277 (N_37277,N_37134,N_37003);
and U37278 (N_37278,N_37149,N_37076);
or U37279 (N_37279,N_37141,N_37055);
or U37280 (N_37280,N_37089,N_37095);
xor U37281 (N_37281,N_37232,N_37139);
nand U37282 (N_37282,N_37057,N_37054);
and U37283 (N_37283,N_37093,N_37116);
xnor U37284 (N_37284,N_37186,N_37148);
or U37285 (N_37285,N_37101,N_37137);
or U37286 (N_37286,N_37068,N_37222);
xnor U37287 (N_37287,N_37008,N_37063);
and U37288 (N_37288,N_37024,N_37056);
or U37289 (N_37289,N_37040,N_37140);
nor U37290 (N_37290,N_37125,N_37201);
nor U37291 (N_37291,N_37081,N_37018);
nor U37292 (N_37292,N_37037,N_37237);
or U37293 (N_37293,N_37109,N_37006);
and U37294 (N_37294,N_37133,N_37091);
nor U37295 (N_37295,N_37235,N_37214);
nand U37296 (N_37296,N_37159,N_37154);
nand U37297 (N_37297,N_37044,N_37191);
nand U37298 (N_37298,N_37113,N_37216);
xnor U37299 (N_37299,N_37009,N_37168);
or U37300 (N_37300,N_37221,N_37012);
nand U37301 (N_37301,N_37111,N_37114);
and U37302 (N_37302,N_37208,N_37181);
nand U37303 (N_37303,N_37050,N_37145);
xnor U37304 (N_37304,N_37107,N_37165);
or U37305 (N_37305,N_37138,N_37026);
nand U37306 (N_37306,N_37131,N_37155);
and U37307 (N_37307,N_37228,N_37209);
nor U37308 (N_37308,N_37203,N_37061);
nand U37309 (N_37309,N_37161,N_37078);
and U37310 (N_37310,N_37092,N_37205);
or U37311 (N_37311,N_37121,N_37192);
nor U37312 (N_37312,N_37094,N_37013);
or U37313 (N_37313,N_37234,N_37108);
nor U37314 (N_37314,N_37124,N_37167);
and U37315 (N_37315,N_37238,N_37087);
or U37316 (N_37316,N_37001,N_37136);
nand U37317 (N_37317,N_37025,N_37206);
nor U37318 (N_37318,N_37152,N_37015);
nand U37319 (N_37319,N_37226,N_37150);
or U37320 (N_37320,N_37097,N_37243);
and U37321 (N_37321,N_37156,N_37028);
or U37322 (N_37322,N_37039,N_37000);
and U37323 (N_37323,N_37069,N_37160);
nand U37324 (N_37324,N_37120,N_37100);
xor U37325 (N_37325,N_37177,N_37170);
or U37326 (N_37326,N_37219,N_37105);
nand U37327 (N_37327,N_37164,N_37077);
and U37328 (N_37328,N_37212,N_37127);
nand U37329 (N_37329,N_37059,N_37014);
nand U37330 (N_37330,N_37122,N_37248);
nor U37331 (N_37331,N_37058,N_37185);
nor U37332 (N_37332,N_37151,N_37036);
xnor U37333 (N_37333,N_37224,N_37047);
nor U37334 (N_37334,N_37062,N_37106);
and U37335 (N_37335,N_37244,N_37199);
and U37336 (N_37336,N_37245,N_37187);
and U37337 (N_37337,N_37033,N_37242);
nor U37338 (N_37338,N_37098,N_37088);
xor U37339 (N_37339,N_37227,N_37045);
nor U37340 (N_37340,N_37171,N_37110);
xor U37341 (N_37341,N_37046,N_37172);
nand U37342 (N_37342,N_37027,N_37083);
or U37343 (N_37343,N_37010,N_37213);
nand U37344 (N_37344,N_37180,N_37118);
or U37345 (N_37345,N_37166,N_37038);
xor U37346 (N_37346,N_37123,N_37207);
nand U37347 (N_37347,N_37240,N_37052);
and U37348 (N_37348,N_37202,N_37017);
xnor U37349 (N_37349,N_37195,N_37005);
xnor U37350 (N_37350,N_37032,N_37130);
xor U37351 (N_37351,N_37074,N_37034);
nand U37352 (N_37352,N_37157,N_37247);
or U37353 (N_37353,N_37204,N_37064);
and U37354 (N_37354,N_37184,N_37246);
nor U37355 (N_37355,N_37103,N_37070);
xnor U37356 (N_37356,N_37060,N_37073);
nand U37357 (N_37357,N_37019,N_37086);
and U37358 (N_37358,N_37007,N_37085);
nand U37359 (N_37359,N_37065,N_37023);
and U37360 (N_37360,N_37196,N_37210);
or U37361 (N_37361,N_37178,N_37099);
nand U37362 (N_37362,N_37217,N_37241);
nor U37363 (N_37363,N_37004,N_37082);
nor U37364 (N_37364,N_37031,N_37022);
or U37365 (N_37365,N_37173,N_37029);
xor U37366 (N_37366,N_37229,N_37021);
xor U37367 (N_37367,N_37189,N_37194);
or U37368 (N_37368,N_37117,N_37142);
xnor U37369 (N_37369,N_37169,N_37197);
nand U37370 (N_37370,N_37090,N_37223);
and U37371 (N_37371,N_37011,N_37211);
or U37372 (N_37372,N_37176,N_37236);
nor U37373 (N_37373,N_37048,N_37126);
nor U37374 (N_37374,N_37084,N_37043);
or U37375 (N_37375,N_37179,N_37232);
or U37376 (N_37376,N_37041,N_37042);
nor U37377 (N_37377,N_37115,N_37157);
and U37378 (N_37378,N_37113,N_37170);
and U37379 (N_37379,N_37186,N_37239);
nor U37380 (N_37380,N_37150,N_37032);
and U37381 (N_37381,N_37050,N_37166);
or U37382 (N_37382,N_37033,N_37244);
nor U37383 (N_37383,N_37069,N_37106);
and U37384 (N_37384,N_37057,N_37221);
xnor U37385 (N_37385,N_37014,N_37221);
xnor U37386 (N_37386,N_37046,N_37057);
nor U37387 (N_37387,N_37093,N_37170);
and U37388 (N_37388,N_37223,N_37150);
or U37389 (N_37389,N_37110,N_37117);
nand U37390 (N_37390,N_37194,N_37162);
nor U37391 (N_37391,N_37081,N_37190);
and U37392 (N_37392,N_37059,N_37140);
nor U37393 (N_37393,N_37095,N_37190);
and U37394 (N_37394,N_37156,N_37165);
and U37395 (N_37395,N_37212,N_37080);
xnor U37396 (N_37396,N_37212,N_37025);
and U37397 (N_37397,N_37004,N_37043);
and U37398 (N_37398,N_37071,N_37149);
xnor U37399 (N_37399,N_37131,N_37208);
or U37400 (N_37400,N_37188,N_37120);
xnor U37401 (N_37401,N_37028,N_37229);
or U37402 (N_37402,N_37185,N_37071);
nor U37403 (N_37403,N_37172,N_37247);
and U37404 (N_37404,N_37146,N_37028);
and U37405 (N_37405,N_37069,N_37228);
and U37406 (N_37406,N_37221,N_37102);
xnor U37407 (N_37407,N_37244,N_37243);
or U37408 (N_37408,N_37137,N_37181);
nor U37409 (N_37409,N_37115,N_37046);
nor U37410 (N_37410,N_37053,N_37044);
xnor U37411 (N_37411,N_37042,N_37224);
nor U37412 (N_37412,N_37109,N_37239);
nor U37413 (N_37413,N_37036,N_37237);
and U37414 (N_37414,N_37059,N_37049);
and U37415 (N_37415,N_37083,N_37018);
or U37416 (N_37416,N_37181,N_37203);
xnor U37417 (N_37417,N_37139,N_37064);
nor U37418 (N_37418,N_37087,N_37030);
nand U37419 (N_37419,N_37202,N_37226);
and U37420 (N_37420,N_37010,N_37172);
or U37421 (N_37421,N_37001,N_37205);
and U37422 (N_37422,N_37050,N_37185);
or U37423 (N_37423,N_37008,N_37101);
and U37424 (N_37424,N_37249,N_37003);
nand U37425 (N_37425,N_37101,N_37125);
nand U37426 (N_37426,N_37106,N_37171);
and U37427 (N_37427,N_37045,N_37211);
or U37428 (N_37428,N_37065,N_37227);
xor U37429 (N_37429,N_37019,N_37189);
xnor U37430 (N_37430,N_37172,N_37051);
or U37431 (N_37431,N_37183,N_37249);
and U37432 (N_37432,N_37128,N_37046);
nand U37433 (N_37433,N_37147,N_37206);
and U37434 (N_37434,N_37092,N_37048);
xnor U37435 (N_37435,N_37226,N_37206);
xnor U37436 (N_37436,N_37202,N_37210);
and U37437 (N_37437,N_37177,N_37090);
nand U37438 (N_37438,N_37083,N_37014);
nor U37439 (N_37439,N_37132,N_37142);
xnor U37440 (N_37440,N_37113,N_37054);
nand U37441 (N_37441,N_37153,N_37118);
or U37442 (N_37442,N_37005,N_37174);
nand U37443 (N_37443,N_37021,N_37213);
and U37444 (N_37444,N_37114,N_37139);
nand U37445 (N_37445,N_37083,N_37243);
and U37446 (N_37446,N_37183,N_37128);
nand U37447 (N_37447,N_37043,N_37167);
xor U37448 (N_37448,N_37224,N_37205);
nor U37449 (N_37449,N_37067,N_37116);
xor U37450 (N_37450,N_37098,N_37081);
or U37451 (N_37451,N_37085,N_37057);
or U37452 (N_37452,N_37058,N_37218);
and U37453 (N_37453,N_37242,N_37018);
or U37454 (N_37454,N_37190,N_37074);
xnor U37455 (N_37455,N_37136,N_37180);
nand U37456 (N_37456,N_37061,N_37092);
nand U37457 (N_37457,N_37056,N_37230);
nand U37458 (N_37458,N_37097,N_37068);
nand U37459 (N_37459,N_37192,N_37212);
or U37460 (N_37460,N_37116,N_37089);
and U37461 (N_37461,N_37238,N_37129);
and U37462 (N_37462,N_37142,N_37064);
nor U37463 (N_37463,N_37148,N_37006);
nor U37464 (N_37464,N_37206,N_37108);
nor U37465 (N_37465,N_37129,N_37078);
nor U37466 (N_37466,N_37237,N_37139);
xor U37467 (N_37467,N_37213,N_37066);
xnor U37468 (N_37468,N_37142,N_37065);
nor U37469 (N_37469,N_37011,N_37237);
nor U37470 (N_37470,N_37179,N_37060);
and U37471 (N_37471,N_37105,N_37036);
and U37472 (N_37472,N_37004,N_37060);
or U37473 (N_37473,N_37242,N_37034);
nor U37474 (N_37474,N_37174,N_37137);
nor U37475 (N_37475,N_37126,N_37116);
nor U37476 (N_37476,N_37216,N_37059);
or U37477 (N_37477,N_37057,N_37056);
xor U37478 (N_37478,N_37117,N_37057);
xnor U37479 (N_37479,N_37177,N_37043);
and U37480 (N_37480,N_37005,N_37045);
and U37481 (N_37481,N_37206,N_37018);
xor U37482 (N_37482,N_37197,N_37222);
and U37483 (N_37483,N_37142,N_37115);
xnor U37484 (N_37484,N_37207,N_37246);
nand U37485 (N_37485,N_37099,N_37134);
nand U37486 (N_37486,N_37050,N_37054);
and U37487 (N_37487,N_37035,N_37151);
xor U37488 (N_37488,N_37201,N_37110);
or U37489 (N_37489,N_37186,N_37224);
or U37490 (N_37490,N_37043,N_37062);
or U37491 (N_37491,N_37066,N_37043);
xor U37492 (N_37492,N_37160,N_37026);
xnor U37493 (N_37493,N_37151,N_37198);
nand U37494 (N_37494,N_37015,N_37218);
or U37495 (N_37495,N_37062,N_37016);
nor U37496 (N_37496,N_37162,N_37059);
xor U37497 (N_37497,N_37059,N_37113);
nand U37498 (N_37498,N_37243,N_37171);
or U37499 (N_37499,N_37136,N_37075);
or U37500 (N_37500,N_37481,N_37345);
and U37501 (N_37501,N_37381,N_37408);
and U37502 (N_37502,N_37322,N_37474);
xor U37503 (N_37503,N_37429,N_37483);
and U37504 (N_37504,N_37486,N_37342);
and U37505 (N_37505,N_37457,N_37441);
xnor U37506 (N_37506,N_37434,N_37276);
and U37507 (N_37507,N_37437,N_37360);
and U37508 (N_37508,N_37371,N_37301);
xor U37509 (N_37509,N_37422,N_37480);
and U37510 (N_37510,N_37375,N_37361);
xnor U37511 (N_37511,N_37449,N_37330);
or U37512 (N_37512,N_37485,N_37418);
nand U37513 (N_37513,N_37452,N_37430);
or U37514 (N_37514,N_37382,N_37320);
or U37515 (N_37515,N_37257,N_37315);
and U37516 (N_37516,N_37388,N_37324);
or U37517 (N_37517,N_37458,N_37451);
or U37518 (N_37518,N_37367,N_37396);
or U37519 (N_37519,N_37406,N_37411);
nand U37520 (N_37520,N_37392,N_37386);
nor U37521 (N_37521,N_37271,N_37393);
nand U37522 (N_37522,N_37472,N_37496);
and U37523 (N_37523,N_37385,N_37425);
and U37524 (N_37524,N_37407,N_37479);
xor U37525 (N_37525,N_37337,N_37369);
nand U37526 (N_37526,N_37468,N_37464);
or U37527 (N_37527,N_37387,N_37476);
nor U37528 (N_37528,N_37498,N_37269);
xor U37529 (N_37529,N_37357,N_37465);
nor U37530 (N_37530,N_37426,N_37350);
and U37531 (N_37531,N_37366,N_37376);
nor U37532 (N_37532,N_37277,N_37435);
or U37533 (N_37533,N_37318,N_37444);
xor U37534 (N_37534,N_37353,N_37492);
xnor U37535 (N_37535,N_37493,N_37478);
or U37536 (N_37536,N_37332,N_37497);
xor U37537 (N_37537,N_37368,N_37329);
xnor U37538 (N_37538,N_37292,N_37346);
or U37539 (N_37539,N_37298,N_37421);
nand U37540 (N_37540,N_37400,N_37370);
nor U37541 (N_37541,N_37340,N_37462);
nor U37542 (N_37542,N_37494,N_37454);
or U37543 (N_37543,N_37442,N_37440);
and U37544 (N_37544,N_37279,N_37309);
xor U37545 (N_37545,N_37267,N_37455);
and U37546 (N_37546,N_37383,N_37335);
or U37547 (N_37547,N_37352,N_37263);
or U37548 (N_37548,N_37287,N_37447);
nor U37549 (N_37549,N_37272,N_37488);
or U37550 (N_37550,N_37414,N_37365);
and U37551 (N_37551,N_37412,N_37373);
nor U37552 (N_37552,N_37323,N_37258);
nand U37553 (N_37553,N_37348,N_37372);
xor U37554 (N_37554,N_37261,N_37336);
xor U37555 (N_37555,N_37390,N_37326);
or U37556 (N_37556,N_37433,N_37300);
nor U37557 (N_37557,N_37467,N_37317);
nand U37558 (N_37558,N_37253,N_37311);
xor U37559 (N_37559,N_37351,N_37338);
nand U37560 (N_37560,N_37410,N_37450);
and U37561 (N_37561,N_37307,N_37379);
xor U37562 (N_37562,N_37297,N_37265);
or U37563 (N_37563,N_37423,N_37417);
or U37564 (N_37564,N_37347,N_37402);
nand U37565 (N_37565,N_37331,N_37349);
xor U37566 (N_37566,N_37362,N_37398);
xnor U37567 (N_37567,N_37397,N_37256);
and U37568 (N_37568,N_37487,N_37274);
and U37569 (N_37569,N_37254,N_37296);
nor U37570 (N_37570,N_37312,N_37355);
nor U37571 (N_37571,N_37270,N_37499);
or U37572 (N_37572,N_37252,N_37327);
and U37573 (N_37573,N_37358,N_37389);
and U37574 (N_37574,N_37466,N_37328);
or U37575 (N_37575,N_37319,N_37333);
nor U37576 (N_37576,N_37443,N_37284);
nor U37577 (N_37577,N_37461,N_37420);
nand U37578 (N_37578,N_37306,N_37334);
nand U37579 (N_37579,N_37294,N_37424);
and U37580 (N_37580,N_37446,N_37303);
nand U37581 (N_37581,N_37401,N_37282);
xor U37582 (N_37582,N_37290,N_37310);
nand U37583 (N_37583,N_37473,N_37490);
or U37584 (N_37584,N_37364,N_37439);
and U37585 (N_37585,N_37341,N_37374);
xor U37586 (N_37586,N_37302,N_37289);
nor U37587 (N_37587,N_37291,N_37495);
or U37588 (N_37588,N_37463,N_37308);
xnor U37589 (N_37589,N_37380,N_37384);
xor U37590 (N_37590,N_37286,N_37415);
and U37591 (N_37591,N_37268,N_37394);
nand U37592 (N_37592,N_37280,N_37399);
and U37593 (N_37593,N_37293,N_37343);
and U37594 (N_37594,N_37484,N_37344);
or U37595 (N_37595,N_37448,N_37438);
nor U37596 (N_37596,N_37339,N_37459);
nand U37597 (N_37597,N_37378,N_37391);
xnor U37598 (N_37598,N_37453,N_37471);
xor U37599 (N_37599,N_37470,N_37255);
nand U37600 (N_37600,N_37305,N_37285);
and U37601 (N_37601,N_37266,N_37404);
or U37602 (N_37602,N_37283,N_37288);
nand U37603 (N_37603,N_37419,N_37405);
xnor U37604 (N_37604,N_37356,N_37482);
or U37605 (N_37605,N_37445,N_37359);
and U37606 (N_37606,N_37363,N_37262);
and U37607 (N_37607,N_37477,N_37489);
nand U37608 (N_37608,N_37260,N_37409);
nand U37609 (N_37609,N_37259,N_37281);
xor U37610 (N_37610,N_37299,N_37431);
and U37611 (N_37611,N_37251,N_37395);
and U37612 (N_37612,N_37321,N_37436);
xnor U37613 (N_37613,N_37314,N_37273);
nand U37614 (N_37614,N_37377,N_37427);
nand U37615 (N_37615,N_37413,N_37460);
and U37616 (N_37616,N_37469,N_37250);
xnor U37617 (N_37617,N_37304,N_37313);
or U37618 (N_37618,N_37475,N_37416);
nor U37619 (N_37619,N_37428,N_37295);
nor U37620 (N_37620,N_37403,N_37354);
nand U37621 (N_37621,N_37264,N_37432);
nand U37622 (N_37622,N_37278,N_37275);
xor U37623 (N_37623,N_37456,N_37325);
nand U37624 (N_37624,N_37316,N_37491);
or U37625 (N_37625,N_37263,N_37283);
nand U37626 (N_37626,N_37452,N_37474);
xnor U37627 (N_37627,N_37261,N_37328);
and U37628 (N_37628,N_37483,N_37334);
and U37629 (N_37629,N_37268,N_37330);
and U37630 (N_37630,N_37264,N_37259);
nor U37631 (N_37631,N_37304,N_37459);
or U37632 (N_37632,N_37448,N_37437);
xnor U37633 (N_37633,N_37487,N_37429);
xor U37634 (N_37634,N_37451,N_37306);
nor U37635 (N_37635,N_37395,N_37400);
xor U37636 (N_37636,N_37466,N_37416);
or U37637 (N_37637,N_37255,N_37364);
xor U37638 (N_37638,N_37416,N_37425);
nand U37639 (N_37639,N_37413,N_37452);
xnor U37640 (N_37640,N_37324,N_37279);
or U37641 (N_37641,N_37282,N_37299);
xnor U37642 (N_37642,N_37367,N_37366);
or U37643 (N_37643,N_37346,N_37254);
xnor U37644 (N_37644,N_37315,N_37499);
and U37645 (N_37645,N_37328,N_37268);
or U37646 (N_37646,N_37471,N_37345);
or U37647 (N_37647,N_37356,N_37403);
xor U37648 (N_37648,N_37381,N_37422);
xor U37649 (N_37649,N_37328,N_37494);
or U37650 (N_37650,N_37341,N_37378);
nor U37651 (N_37651,N_37494,N_37457);
xor U37652 (N_37652,N_37353,N_37330);
nor U37653 (N_37653,N_37429,N_37497);
nor U37654 (N_37654,N_37359,N_37299);
nor U37655 (N_37655,N_37483,N_37423);
xnor U37656 (N_37656,N_37355,N_37378);
nand U37657 (N_37657,N_37432,N_37253);
or U37658 (N_37658,N_37428,N_37478);
nor U37659 (N_37659,N_37318,N_37442);
or U37660 (N_37660,N_37426,N_37250);
or U37661 (N_37661,N_37314,N_37463);
nor U37662 (N_37662,N_37254,N_37306);
and U37663 (N_37663,N_37418,N_37431);
xor U37664 (N_37664,N_37359,N_37422);
xor U37665 (N_37665,N_37451,N_37349);
and U37666 (N_37666,N_37314,N_37347);
or U37667 (N_37667,N_37464,N_37278);
xnor U37668 (N_37668,N_37329,N_37327);
xnor U37669 (N_37669,N_37395,N_37261);
and U37670 (N_37670,N_37426,N_37422);
or U37671 (N_37671,N_37434,N_37353);
xnor U37672 (N_37672,N_37303,N_37377);
xnor U37673 (N_37673,N_37272,N_37489);
nand U37674 (N_37674,N_37289,N_37381);
nand U37675 (N_37675,N_37317,N_37433);
or U37676 (N_37676,N_37453,N_37317);
or U37677 (N_37677,N_37287,N_37301);
nand U37678 (N_37678,N_37387,N_37468);
xor U37679 (N_37679,N_37462,N_37350);
nor U37680 (N_37680,N_37436,N_37383);
nand U37681 (N_37681,N_37259,N_37278);
nor U37682 (N_37682,N_37412,N_37366);
or U37683 (N_37683,N_37323,N_37376);
or U37684 (N_37684,N_37356,N_37490);
nor U37685 (N_37685,N_37293,N_37334);
nand U37686 (N_37686,N_37423,N_37288);
and U37687 (N_37687,N_37352,N_37359);
nor U37688 (N_37688,N_37397,N_37407);
xor U37689 (N_37689,N_37273,N_37274);
nand U37690 (N_37690,N_37372,N_37443);
nor U37691 (N_37691,N_37328,N_37325);
xnor U37692 (N_37692,N_37435,N_37328);
xnor U37693 (N_37693,N_37339,N_37269);
and U37694 (N_37694,N_37472,N_37447);
or U37695 (N_37695,N_37384,N_37338);
or U37696 (N_37696,N_37463,N_37386);
xor U37697 (N_37697,N_37455,N_37288);
nor U37698 (N_37698,N_37458,N_37284);
or U37699 (N_37699,N_37457,N_37412);
or U37700 (N_37700,N_37417,N_37266);
or U37701 (N_37701,N_37396,N_37314);
or U37702 (N_37702,N_37278,N_37331);
nor U37703 (N_37703,N_37340,N_37412);
and U37704 (N_37704,N_37291,N_37479);
or U37705 (N_37705,N_37317,N_37300);
and U37706 (N_37706,N_37338,N_37399);
and U37707 (N_37707,N_37494,N_37451);
or U37708 (N_37708,N_37302,N_37424);
nand U37709 (N_37709,N_37376,N_37377);
nand U37710 (N_37710,N_37391,N_37478);
nor U37711 (N_37711,N_37252,N_37456);
nand U37712 (N_37712,N_37323,N_37366);
and U37713 (N_37713,N_37413,N_37351);
nand U37714 (N_37714,N_37365,N_37387);
nand U37715 (N_37715,N_37450,N_37275);
xor U37716 (N_37716,N_37283,N_37337);
and U37717 (N_37717,N_37361,N_37455);
and U37718 (N_37718,N_37359,N_37428);
and U37719 (N_37719,N_37391,N_37276);
nor U37720 (N_37720,N_37313,N_37302);
xnor U37721 (N_37721,N_37296,N_37282);
xor U37722 (N_37722,N_37494,N_37259);
xnor U37723 (N_37723,N_37318,N_37301);
and U37724 (N_37724,N_37304,N_37276);
nor U37725 (N_37725,N_37347,N_37285);
or U37726 (N_37726,N_37430,N_37333);
xnor U37727 (N_37727,N_37447,N_37410);
xnor U37728 (N_37728,N_37491,N_37277);
xnor U37729 (N_37729,N_37425,N_37257);
xnor U37730 (N_37730,N_37440,N_37383);
nor U37731 (N_37731,N_37320,N_37281);
and U37732 (N_37732,N_37322,N_37413);
nor U37733 (N_37733,N_37451,N_37438);
xor U37734 (N_37734,N_37496,N_37274);
nor U37735 (N_37735,N_37479,N_37339);
or U37736 (N_37736,N_37444,N_37366);
xnor U37737 (N_37737,N_37342,N_37387);
or U37738 (N_37738,N_37265,N_37299);
xor U37739 (N_37739,N_37268,N_37374);
nand U37740 (N_37740,N_37367,N_37335);
xor U37741 (N_37741,N_37427,N_37478);
nand U37742 (N_37742,N_37269,N_37369);
nand U37743 (N_37743,N_37345,N_37268);
nor U37744 (N_37744,N_37265,N_37486);
or U37745 (N_37745,N_37363,N_37474);
nor U37746 (N_37746,N_37268,N_37314);
and U37747 (N_37747,N_37265,N_37292);
or U37748 (N_37748,N_37265,N_37444);
xor U37749 (N_37749,N_37404,N_37265);
nand U37750 (N_37750,N_37705,N_37728);
and U37751 (N_37751,N_37590,N_37628);
nand U37752 (N_37752,N_37617,N_37684);
xor U37753 (N_37753,N_37502,N_37651);
xnor U37754 (N_37754,N_37537,N_37587);
or U37755 (N_37755,N_37678,N_37719);
or U37756 (N_37756,N_37508,N_37646);
and U37757 (N_37757,N_37657,N_37515);
or U37758 (N_37758,N_37538,N_37732);
and U37759 (N_37759,N_37711,N_37606);
nor U37760 (N_37760,N_37668,N_37697);
xnor U37761 (N_37761,N_37607,N_37706);
and U37762 (N_37762,N_37681,N_37557);
xnor U37763 (N_37763,N_37644,N_37520);
xor U37764 (N_37764,N_37660,N_37730);
xnor U37765 (N_37765,N_37650,N_37688);
xor U37766 (N_37766,N_37709,N_37610);
xnor U37767 (N_37767,N_37589,N_37626);
nand U37768 (N_37768,N_37721,N_37613);
or U37769 (N_37769,N_37661,N_37726);
nor U37770 (N_37770,N_37528,N_37696);
nand U37771 (N_37771,N_37703,N_37655);
and U37772 (N_37772,N_37550,N_37682);
nor U37773 (N_37773,N_37566,N_37573);
nand U37774 (N_37774,N_37509,N_37531);
and U37775 (N_37775,N_37653,N_37600);
nor U37776 (N_37776,N_37586,N_37634);
nand U37777 (N_37777,N_37677,N_37629);
nand U37778 (N_37778,N_37574,N_37625);
or U37779 (N_37779,N_37701,N_37690);
nand U37780 (N_37780,N_37718,N_37627);
nor U37781 (N_37781,N_37720,N_37619);
and U37782 (N_37782,N_37702,N_37708);
or U37783 (N_37783,N_37689,N_37570);
nor U37784 (N_37784,N_37580,N_37740);
and U37785 (N_37785,N_37554,N_37680);
nor U37786 (N_37786,N_37699,N_37741);
nand U37787 (N_37787,N_37673,N_37547);
nor U37788 (N_37788,N_37665,N_37581);
and U37789 (N_37789,N_37608,N_37624);
nor U37790 (N_37790,N_37541,N_37659);
xor U37791 (N_37791,N_37664,N_37694);
xor U37792 (N_37792,N_37676,N_37739);
or U37793 (N_37793,N_37542,N_37748);
xnor U37794 (N_37794,N_37593,N_37723);
xnor U37795 (N_37795,N_37525,N_37743);
xor U37796 (N_37796,N_37514,N_37633);
nand U37797 (N_37797,N_37717,N_37507);
nor U37798 (N_37798,N_37545,N_37602);
or U37799 (N_37799,N_37631,N_37548);
nor U37800 (N_37800,N_37715,N_37724);
or U37801 (N_37801,N_37562,N_37618);
xnor U37802 (N_37802,N_37666,N_37506);
and U37803 (N_37803,N_37603,N_37518);
xor U37804 (N_37804,N_37579,N_37667);
nand U37805 (N_37805,N_37536,N_37539);
nand U37806 (N_37806,N_37577,N_37636);
xnor U37807 (N_37807,N_37745,N_37611);
nor U37808 (N_37808,N_37555,N_37513);
nand U37809 (N_37809,N_37713,N_37652);
and U37810 (N_37810,N_37549,N_37595);
and U37811 (N_37811,N_37698,N_37746);
nand U37812 (N_37812,N_37642,N_37516);
nor U37813 (N_37813,N_37686,N_37614);
xor U37814 (N_37814,N_37683,N_37558);
and U37815 (N_37815,N_37530,N_37532);
or U37816 (N_37816,N_37725,N_37576);
and U37817 (N_37817,N_37744,N_37575);
xnor U37818 (N_37818,N_37588,N_37523);
or U37819 (N_37819,N_37714,N_37687);
nor U37820 (N_37820,N_37679,N_37674);
nand U37821 (N_37821,N_37616,N_37529);
and U37822 (N_37822,N_37729,N_37567);
or U37823 (N_37823,N_37597,N_37630);
nand U37824 (N_37824,N_37716,N_37727);
nor U37825 (N_37825,N_37521,N_37583);
nand U37826 (N_37826,N_37691,N_37578);
nor U37827 (N_37827,N_37564,N_37737);
nand U37828 (N_37828,N_37571,N_37707);
and U37829 (N_37829,N_37585,N_37669);
nand U37830 (N_37830,N_37621,N_37734);
or U37831 (N_37831,N_37623,N_37556);
xor U37832 (N_37832,N_37722,N_37663);
xor U37833 (N_37833,N_37612,N_37569);
nand U37834 (N_37834,N_37662,N_37693);
xor U37835 (N_37835,N_37598,N_37543);
or U37836 (N_37836,N_37654,N_37533);
nand U37837 (N_37837,N_37637,N_37519);
nand U37838 (N_37838,N_37639,N_37517);
and U37839 (N_37839,N_37632,N_37710);
or U37840 (N_37840,N_37526,N_37648);
xor U37841 (N_37841,N_37671,N_37615);
or U37842 (N_37842,N_37700,N_37658);
nand U37843 (N_37843,N_37546,N_37609);
xnor U37844 (N_37844,N_37512,N_37604);
or U37845 (N_37845,N_37561,N_37647);
nand U37846 (N_37846,N_37511,N_37544);
nand U37847 (N_37847,N_37594,N_37656);
and U37848 (N_37848,N_37649,N_37692);
xor U37849 (N_37849,N_37524,N_37735);
and U37850 (N_37850,N_37638,N_37553);
or U37851 (N_37851,N_37572,N_37559);
nand U37852 (N_37852,N_37641,N_37584);
and U37853 (N_37853,N_37695,N_37596);
or U37854 (N_37854,N_37522,N_37563);
nor U37855 (N_37855,N_37599,N_37685);
and U37856 (N_37856,N_37568,N_37736);
nor U37857 (N_37857,N_37601,N_37582);
and U37858 (N_37858,N_37503,N_37704);
xnor U37859 (N_37859,N_37622,N_37505);
nor U37860 (N_37860,N_37670,N_37635);
or U37861 (N_37861,N_37672,N_37747);
nand U37862 (N_37862,N_37605,N_37738);
xor U37863 (N_37863,N_37500,N_37501);
nor U37864 (N_37864,N_37645,N_37712);
and U37865 (N_37865,N_37551,N_37560);
nor U37866 (N_37866,N_37675,N_37742);
nand U37867 (N_37867,N_37535,N_37749);
nor U37868 (N_37868,N_37731,N_37592);
nand U37869 (N_37869,N_37640,N_37534);
xor U37870 (N_37870,N_37504,N_37527);
xor U37871 (N_37871,N_37591,N_37510);
or U37872 (N_37872,N_37643,N_37540);
or U37873 (N_37873,N_37620,N_37733);
xor U37874 (N_37874,N_37565,N_37552);
nor U37875 (N_37875,N_37735,N_37507);
and U37876 (N_37876,N_37655,N_37606);
nor U37877 (N_37877,N_37599,N_37745);
or U37878 (N_37878,N_37571,N_37567);
or U37879 (N_37879,N_37749,N_37635);
xnor U37880 (N_37880,N_37708,N_37694);
nor U37881 (N_37881,N_37637,N_37730);
nand U37882 (N_37882,N_37603,N_37632);
nand U37883 (N_37883,N_37626,N_37564);
or U37884 (N_37884,N_37559,N_37585);
nand U37885 (N_37885,N_37547,N_37686);
and U37886 (N_37886,N_37685,N_37563);
or U37887 (N_37887,N_37703,N_37744);
nor U37888 (N_37888,N_37552,N_37690);
nand U37889 (N_37889,N_37638,N_37567);
and U37890 (N_37890,N_37601,N_37553);
and U37891 (N_37891,N_37532,N_37560);
nand U37892 (N_37892,N_37555,N_37663);
and U37893 (N_37893,N_37686,N_37611);
nand U37894 (N_37894,N_37564,N_37562);
xnor U37895 (N_37895,N_37695,N_37513);
nor U37896 (N_37896,N_37683,N_37524);
nor U37897 (N_37897,N_37724,N_37541);
and U37898 (N_37898,N_37713,N_37588);
nor U37899 (N_37899,N_37682,N_37563);
nor U37900 (N_37900,N_37742,N_37533);
or U37901 (N_37901,N_37599,N_37536);
nor U37902 (N_37902,N_37639,N_37528);
xnor U37903 (N_37903,N_37709,N_37559);
nand U37904 (N_37904,N_37639,N_37613);
nor U37905 (N_37905,N_37714,N_37559);
and U37906 (N_37906,N_37609,N_37516);
xor U37907 (N_37907,N_37638,N_37650);
and U37908 (N_37908,N_37520,N_37681);
and U37909 (N_37909,N_37572,N_37642);
xnor U37910 (N_37910,N_37527,N_37726);
xnor U37911 (N_37911,N_37626,N_37624);
and U37912 (N_37912,N_37528,N_37607);
and U37913 (N_37913,N_37699,N_37623);
xnor U37914 (N_37914,N_37620,N_37550);
xor U37915 (N_37915,N_37722,N_37677);
or U37916 (N_37916,N_37504,N_37612);
nand U37917 (N_37917,N_37653,N_37699);
nand U37918 (N_37918,N_37562,N_37599);
nand U37919 (N_37919,N_37668,N_37728);
and U37920 (N_37920,N_37723,N_37562);
and U37921 (N_37921,N_37587,N_37586);
nor U37922 (N_37922,N_37513,N_37745);
xnor U37923 (N_37923,N_37742,N_37703);
nand U37924 (N_37924,N_37657,N_37650);
and U37925 (N_37925,N_37619,N_37511);
nor U37926 (N_37926,N_37601,N_37658);
xor U37927 (N_37927,N_37693,N_37631);
nor U37928 (N_37928,N_37589,N_37614);
nand U37929 (N_37929,N_37557,N_37592);
or U37930 (N_37930,N_37566,N_37628);
nor U37931 (N_37931,N_37573,N_37541);
xor U37932 (N_37932,N_37609,N_37740);
and U37933 (N_37933,N_37536,N_37654);
and U37934 (N_37934,N_37667,N_37583);
nor U37935 (N_37935,N_37611,N_37733);
nor U37936 (N_37936,N_37694,N_37663);
xor U37937 (N_37937,N_37687,N_37540);
nand U37938 (N_37938,N_37741,N_37593);
and U37939 (N_37939,N_37638,N_37732);
xor U37940 (N_37940,N_37529,N_37639);
nor U37941 (N_37941,N_37739,N_37653);
nand U37942 (N_37942,N_37738,N_37717);
nor U37943 (N_37943,N_37708,N_37555);
nand U37944 (N_37944,N_37652,N_37632);
xor U37945 (N_37945,N_37717,N_37716);
or U37946 (N_37946,N_37689,N_37649);
or U37947 (N_37947,N_37566,N_37658);
or U37948 (N_37948,N_37714,N_37639);
nor U37949 (N_37949,N_37673,N_37694);
xor U37950 (N_37950,N_37686,N_37647);
nor U37951 (N_37951,N_37731,N_37582);
and U37952 (N_37952,N_37675,N_37570);
xor U37953 (N_37953,N_37749,N_37508);
nand U37954 (N_37954,N_37735,N_37652);
nand U37955 (N_37955,N_37711,N_37545);
nor U37956 (N_37956,N_37697,N_37698);
or U37957 (N_37957,N_37538,N_37625);
nor U37958 (N_37958,N_37550,N_37606);
nor U37959 (N_37959,N_37526,N_37607);
nor U37960 (N_37960,N_37741,N_37598);
and U37961 (N_37961,N_37719,N_37541);
nand U37962 (N_37962,N_37510,N_37564);
and U37963 (N_37963,N_37653,N_37567);
or U37964 (N_37964,N_37695,N_37508);
xnor U37965 (N_37965,N_37620,N_37605);
xnor U37966 (N_37966,N_37542,N_37572);
or U37967 (N_37967,N_37741,N_37627);
nor U37968 (N_37968,N_37645,N_37706);
nand U37969 (N_37969,N_37648,N_37742);
xor U37970 (N_37970,N_37738,N_37647);
and U37971 (N_37971,N_37737,N_37532);
nand U37972 (N_37972,N_37553,N_37623);
nand U37973 (N_37973,N_37742,N_37668);
and U37974 (N_37974,N_37653,N_37662);
or U37975 (N_37975,N_37712,N_37749);
or U37976 (N_37976,N_37680,N_37528);
nor U37977 (N_37977,N_37667,N_37524);
or U37978 (N_37978,N_37669,N_37722);
xor U37979 (N_37979,N_37664,N_37737);
xor U37980 (N_37980,N_37662,N_37609);
or U37981 (N_37981,N_37631,N_37543);
or U37982 (N_37982,N_37574,N_37668);
and U37983 (N_37983,N_37546,N_37577);
and U37984 (N_37984,N_37667,N_37737);
xnor U37985 (N_37985,N_37678,N_37692);
or U37986 (N_37986,N_37700,N_37562);
or U37987 (N_37987,N_37620,N_37734);
nand U37988 (N_37988,N_37636,N_37617);
or U37989 (N_37989,N_37539,N_37630);
nor U37990 (N_37990,N_37593,N_37661);
xnor U37991 (N_37991,N_37526,N_37560);
or U37992 (N_37992,N_37618,N_37509);
nor U37993 (N_37993,N_37630,N_37734);
and U37994 (N_37994,N_37712,N_37745);
and U37995 (N_37995,N_37610,N_37738);
xor U37996 (N_37996,N_37673,N_37619);
nand U37997 (N_37997,N_37726,N_37669);
and U37998 (N_37998,N_37557,N_37653);
or U37999 (N_37999,N_37605,N_37712);
nand U38000 (N_38000,N_37856,N_37974);
nor U38001 (N_38001,N_37801,N_37967);
xnor U38002 (N_38002,N_37898,N_37784);
and U38003 (N_38003,N_37899,N_37954);
nor U38004 (N_38004,N_37786,N_37972);
nand U38005 (N_38005,N_37829,N_37960);
xnor U38006 (N_38006,N_37939,N_37908);
xnor U38007 (N_38007,N_37971,N_37878);
or U38008 (N_38008,N_37812,N_37782);
and U38009 (N_38009,N_37894,N_37930);
and U38010 (N_38010,N_37839,N_37868);
or U38011 (N_38011,N_37961,N_37944);
xnor U38012 (N_38012,N_37857,N_37850);
nor U38013 (N_38013,N_37771,N_37854);
or U38014 (N_38014,N_37871,N_37869);
xnor U38015 (N_38015,N_37919,N_37800);
and U38016 (N_38016,N_37982,N_37835);
xor U38017 (N_38017,N_37807,N_37844);
or U38018 (N_38018,N_37912,N_37947);
or U38019 (N_38019,N_37918,N_37826);
nand U38020 (N_38020,N_37959,N_37872);
nand U38021 (N_38021,N_37762,N_37875);
nor U38022 (N_38022,N_37996,N_37905);
xor U38023 (N_38023,N_37775,N_37978);
xor U38024 (N_38024,N_37943,N_37805);
nor U38025 (N_38025,N_37847,N_37948);
or U38026 (N_38026,N_37825,N_37883);
nor U38027 (N_38027,N_37936,N_37979);
xor U38028 (N_38028,N_37777,N_37923);
and U38029 (N_38029,N_37901,N_37876);
nand U38030 (N_38030,N_37983,N_37897);
and U38031 (N_38031,N_37952,N_37984);
or U38032 (N_38032,N_37963,N_37796);
xor U38033 (N_38033,N_37773,N_37756);
nor U38034 (N_38034,N_37755,N_37836);
nor U38035 (N_38035,N_37933,N_37956);
or U38036 (N_38036,N_37833,N_37916);
and U38037 (N_38037,N_37750,N_37889);
and U38038 (N_38038,N_37892,N_37760);
or U38039 (N_38039,N_37880,N_37759);
xnor U38040 (N_38040,N_37764,N_37958);
xnor U38041 (N_38041,N_37957,N_37838);
nor U38042 (N_38042,N_37995,N_37953);
nor U38043 (N_38043,N_37998,N_37783);
nor U38044 (N_38044,N_37779,N_37965);
nand U38045 (N_38045,N_37904,N_37862);
xnor U38046 (N_38046,N_37822,N_37798);
nor U38047 (N_38047,N_37931,N_37781);
nand U38048 (N_38048,N_37917,N_37925);
and U38049 (N_38049,N_37962,N_37909);
xnor U38050 (N_38050,N_37840,N_37906);
nand U38051 (N_38051,N_37757,N_37885);
xor U38052 (N_38052,N_37991,N_37831);
nand U38053 (N_38053,N_37993,N_37951);
and U38054 (N_38054,N_37903,N_37942);
xor U38055 (N_38055,N_37858,N_37980);
nor U38056 (N_38056,N_37924,N_37828);
or U38057 (N_38057,N_37874,N_37821);
nand U38058 (N_38058,N_37927,N_37824);
xor U38059 (N_38059,N_37973,N_37846);
xnor U38060 (N_38060,N_37990,N_37830);
nand U38061 (N_38061,N_37761,N_37864);
and U38062 (N_38062,N_37884,N_37969);
and U38063 (N_38063,N_37770,N_37950);
nand U38064 (N_38064,N_37920,N_37819);
xor U38065 (N_38065,N_37992,N_37887);
and U38066 (N_38066,N_37911,N_37896);
and U38067 (N_38067,N_37792,N_37935);
nor U38068 (N_38068,N_37861,N_37852);
and U38069 (N_38069,N_37870,N_37774);
nand U38070 (N_38070,N_37849,N_37845);
or U38071 (N_38071,N_37902,N_37989);
or U38072 (N_38072,N_37976,N_37873);
and U38073 (N_38073,N_37814,N_37785);
or U38074 (N_38074,N_37928,N_37977);
xor U38075 (N_38075,N_37915,N_37809);
nor U38076 (N_38076,N_37769,N_37986);
nand U38077 (N_38077,N_37921,N_37900);
nor U38078 (N_38078,N_37910,N_37797);
xnor U38079 (N_38079,N_37968,N_37997);
or U38080 (N_38080,N_37799,N_37877);
or U38081 (N_38081,N_37981,N_37753);
nor U38082 (N_38082,N_37765,N_37941);
nand U38083 (N_38083,N_37964,N_37949);
and U38084 (N_38084,N_37832,N_37823);
nor U38085 (N_38085,N_37895,N_37865);
nand U38086 (N_38086,N_37780,N_37966);
nor U38087 (N_38087,N_37929,N_37751);
and U38088 (N_38088,N_37945,N_37934);
nand U38089 (N_38089,N_37820,N_37811);
nor U38090 (N_38090,N_37794,N_37818);
and U38091 (N_38091,N_37803,N_37914);
nand U38092 (N_38092,N_37763,N_37913);
nor U38093 (N_38093,N_37907,N_37866);
nand U38094 (N_38094,N_37938,N_37788);
nor U38095 (N_38095,N_37816,N_37975);
nor U38096 (N_38096,N_37817,N_37860);
or U38097 (N_38097,N_37890,N_37863);
and U38098 (N_38098,N_37837,N_37776);
or U38099 (N_38099,N_37787,N_37855);
xor U38100 (N_38100,N_37791,N_37827);
nor U38101 (N_38101,N_37790,N_37888);
and U38102 (N_38102,N_37802,N_37932);
xor U38103 (N_38103,N_37766,N_37795);
and U38104 (N_38104,N_37843,N_37886);
nand U38105 (N_38105,N_37851,N_37804);
or U38106 (N_38106,N_37999,N_37955);
xor U38107 (N_38107,N_37754,N_37859);
xor U38108 (N_38108,N_37772,N_37922);
nor U38109 (N_38109,N_37767,N_37842);
or U38110 (N_38110,N_37758,N_37985);
and U38111 (N_38111,N_37926,N_37994);
nand U38112 (N_38112,N_37937,N_37808);
nand U38113 (N_38113,N_37841,N_37893);
and U38114 (N_38114,N_37881,N_37853);
nor U38115 (N_38115,N_37879,N_37970);
and U38116 (N_38116,N_37810,N_37768);
xor U38117 (N_38117,N_37793,N_37752);
and U38118 (N_38118,N_37806,N_37778);
xor U38119 (N_38119,N_37891,N_37834);
nand U38120 (N_38120,N_37940,N_37813);
or U38121 (N_38121,N_37867,N_37946);
and U38122 (N_38122,N_37882,N_37987);
and U38123 (N_38123,N_37789,N_37988);
xnor U38124 (N_38124,N_37815,N_37848);
nand U38125 (N_38125,N_37781,N_37956);
nand U38126 (N_38126,N_37849,N_37988);
or U38127 (N_38127,N_37976,N_37900);
or U38128 (N_38128,N_37822,N_37766);
or U38129 (N_38129,N_37815,N_37897);
or U38130 (N_38130,N_37991,N_37899);
nand U38131 (N_38131,N_37836,N_37758);
nand U38132 (N_38132,N_37930,N_37893);
xor U38133 (N_38133,N_37821,N_37976);
or U38134 (N_38134,N_37779,N_37879);
or U38135 (N_38135,N_37996,N_37878);
or U38136 (N_38136,N_37822,N_37811);
and U38137 (N_38137,N_37861,N_37811);
or U38138 (N_38138,N_37871,N_37763);
nand U38139 (N_38139,N_37952,N_37789);
nand U38140 (N_38140,N_37899,N_37768);
nand U38141 (N_38141,N_37925,N_37824);
and U38142 (N_38142,N_37963,N_37819);
and U38143 (N_38143,N_37869,N_37896);
nor U38144 (N_38144,N_37995,N_37872);
and U38145 (N_38145,N_37795,N_37920);
nor U38146 (N_38146,N_37794,N_37850);
or U38147 (N_38147,N_37869,N_37850);
nor U38148 (N_38148,N_37916,N_37846);
and U38149 (N_38149,N_37825,N_37786);
nand U38150 (N_38150,N_37758,N_37864);
nand U38151 (N_38151,N_37787,N_37819);
or U38152 (N_38152,N_37902,N_37772);
and U38153 (N_38153,N_37781,N_37795);
nand U38154 (N_38154,N_37781,N_37916);
nand U38155 (N_38155,N_37951,N_37894);
and U38156 (N_38156,N_37927,N_37965);
xnor U38157 (N_38157,N_37835,N_37946);
or U38158 (N_38158,N_37783,N_37898);
nor U38159 (N_38159,N_37932,N_37761);
or U38160 (N_38160,N_37979,N_37973);
and U38161 (N_38161,N_37870,N_37816);
nand U38162 (N_38162,N_37793,N_37892);
nand U38163 (N_38163,N_37870,N_37934);
xor U38164 (N_38164,N_37943,N_37972);
nor U38165 (N_38165,N_37853,N_37816);
xor U38166 (N_38166,N_37828,N_37960);
xor U38167 (N_38167,N_37762,N_37886);
xnor U38168 (N_38168,N_37931,N_37840);
and U38169 (N_38169,N_37770,N_37776);
and U38170 (N_38170,N_37793,N_37975);
nor U38171 (N_38171,N_37939,N_37839);
xnor U38172 (N_38172,N_37973,N_37828);
and U38173 (N_38173,N_37939,N_37763);
or U38174 (N_38174,N_37904,N_37849);
nand U38175 (N_38175,N_37942,N_37926);
nor U38176 (N_38176,N_37862,N_37912);
nand U38177 (N_38177,N_37773,N_37922);
xnor U38178 (N_38178,N_37965,N_37782);
xor U38179 (N_38179,N_37786,N_37961);
nor U38180 (N_38180,N_37940,N_37865);
and U38181 (N_38181,N_37994,N_37764);
nand U38182 (N_38182,N_37887,N_37754);
and U38183 (N_38183,N_37896,N_37867);
nor U38184 (N_38184,N_37783,N_37757);
and U38185 (N_38185,N_37962,N_37768);
and U38186 (N_38186,N_37910,N_37945);
or U38187 (N_38187,N_37848,N_37970);
nand U38188 (N_38188,N_37898,N_37792);
xor U38189 (N_38189,N_37853,N_37775);
and U38190 (N_38190,N_37813,N_37896);
or U38191 (N_38191,N_37930,N_37987);
or U38192 (N_38192,N_37993,N_37983);
xor U38193 (N_38193,N_37808,N_37769);
xnor U38194 (N_38194,N_37832,N_37967);
or U38195 (N_38195,N_37902,N_37767);
or U38196 (N_38196,N_37791,N_37902);
xor U38197 (N_38197,N_37792,N_37850);
or U38198 (N_38198,N_37851,N_37854);
nand U38199 (N_38199,N_37954,N_37890);
nor U38200 (N_38200,N_37791,N_37874);
xnor U38201 (N_38201,N_37936,N_37757);
or U38202 (N_38202,N_37793,N_37845);
and U38203 (N_38203,N_37963,N_37924);
or U38204 (N_38204,N_37950,N_37876);
nand U38205 (N_38205,N_37826,N_37859);
xnor U38206 (N_38206,N_37924,N_37820);
or U38207 (N_38207,N_37846,N_37837);
and U38208 (N_38208,N_37773,N_37764);
and U38209 (N_38209,N_37786,N_37957);
xnor U38210 (N_38210,N_37967,N_37771);
nand U38211 (N_38211,N_37833,N_37875);
and U38212 (N_38212,N_37786,N_37849);
or U38213 (N_38213,N_37903,N_37768);
nor U38214 (N_38214,N_37959,N_37861);
or U38215 (N_38215,N_37752,N_37925);
or U38216 (N_38216,N_37964,N_37775);
xor U38217 (N_38217,N_37957,N_37916);
nor U38218 (N_38218,N_37793,N_37833);
and U38219 (N_38219,N_37816,N_37969);
and U38220 (N_38220,N_37872,N_37868);
nor U38221 (N_38221,N_37985,N_37794);
and U38222 (N_38222,N_37888,N_37767);
xnor U38223 (N_38223,N_37835,N_37898);
and U38224 (N_38224,N_37965,N_37869);
or U38225 (N_38225,N_37806,N_37985);
or U38226 (N_38226,N_37863,N_37874);
and U38227 (N_38227,N_37827,N_37841);
nand U38228 (N_38228,N_37877,N_37942);
xor U38229 (N_38229,N_37846,N_37790);
and U38230 (N_38230,N_37809,N_37887);
nand U38231 (N_38231,N_37979,N_37792);
or U38232 (N_38232,N_37965,N_37988);
or U38233 (N_38233,N_37808,N_37830);
xor U38234 (N_38234,N_37807,N_37770);
and U38235 (N_38235,N_37799,N_37988);
nand U38236 (N_38236,N_37853,N_37926);
and U38237 (N_38237,N_37907,N_37808);
nor U38238 (N_38238,N_37859,N_37799);
or U38239 (N_38239,N_37833,N_37755);
and U38240 (N_38240,N_37867,N_37898);
and U38241 (N_38241,N_37924,N_37787);
or U38242 (N_38242,N_37907,N_37998);
and U38243 (N_38243,N_37810,N_37985);
nand U38244 (N_38244,N_37871,N_37889);
nor U38245 (N_38245,N_37810,N_37833);
xor U38246 (N_38246,N_37925,N_37893);
and U38247 (N_38247,N_37830,N_37941);
nand U38248 (N_38248,N_37834,N_37928);
or U38249 (N_38249,N_37832,N_37752);
or U38250 (N_38250,N_38152,N_38179);
and U38251 (N_38251,N_38135,N_38106);
and U38252 (N_38252,N_38193,N_38025);
and U38253 (N_38253,N_38136,N_38236);
nand U38254 (N_38254,N_38017,N_38117);
nor U38255 (N_38255,N_38125,N_38061);
xor U38256 (N_38256,N_38227,N_38003);
xnor U38257 (N_38257,N_38123,N_38153);
nor U38258 (N_38258,N_38201,N_38062);
xor U38259 (N_38259,N_38079,N_38240);
xor U38260 (N_38260,N_38208,N_38203);
or U38261 (N_38261,N_38202,N_38118);
or U38262 (N_38262,N_38187,N_38165);
nor U38263 (N_38263,N_38073,N_38121);
or U38264 (N_38264,N_38213,N_38128);
or U38265 (N_38265,N_38210,N_38178);
nand U38266 (N_38266,N_38102,N_38022);
or U38267 (N_38267,N_38076,N_38075);
nor U38268 (N_38268,N_38027,N_38249);
or U38269 (N_38269,N_38081,N_38185);
nand U38270 (N_38270,N_38092,N_38232);
nand U38271 (N_38271,N_38130,N_38189);
and U38272 (N_38272,N_38028,N_38084);
and U38273 (N_38273,N_38148,N_38063);
nand U38274 (N_38274,N_38113,N_38037);
xor U38275 (N_38275,N_38188,N_38112);
xor U38276 (N_38276,N_38124,N_38209);
or U38277 (N_38277,N_38248,N_38205);
and U38278 (N_38278,N_38048,N_38020);
and U38279 (N_38279,N_38242,N_38064);
nand U38280 (N_38280,N_38096,N_38230);
xor U38281 (N_38281,N_38039,N_38035);
xor U38282 (N_38282,N_38216,N_38149);
and U38283 (N_38283,N_38002,N_38134);
xor U38284 (N_38284,N_38231,N_38158);
nand U38285 (N_38285,N_38145,N_38246);
or U38286 (N_38286,N_38168,N_38016);
or U38287 (N_38287,N_38157,N_38001);
nand U38288 (N_38288,N_38172,N_38186);
or U38289 (N_38289,N_38247,N_38045);
and U38290 (N_38290,N_38220,N_38103);
nand U38291 (N_38291,N_38226,N_38199);
and U38292 (N_38292,N_38054,N_38160);
nor U38293 (N_38293,N_38009,N_38067);
xor U38294 (N_38294,N_38049,N_38238);
nand U38295 (N_38295,N_38080,N_38085);
xnor U38296 (N_38296,N_38159,N_38083);
or U38297 (N_38297,N_38171,N_38132);
or U38298 (N_38298,N_38018,N_38047);
and U38299 (N_38299,N_38183,N_38107);
nor U38300 (N_38300,N_38089,N_38041);
nor U38301 (N_38301,N_38038,N_38173);
xor U38302 (N_38302,N_38223,N_38059);
nand U38303 (N_38303,N_38221,N_38243);
xor U38304 (N_38304,N_38244,N_38042);
and U38305 (N_38305,N_38099,N_38108);
xor U38306 (N_38306,N_38030,N_38177);
nor U38307 (N_38307,N_38215,N_38197);
nand U38308 (N_38308,N_38196,N_38139);
nor U38309 (N_38309,N_38077,N_38235);
and U38310 (N_38310,N_38225,N_38182);
nand U38311 (N_38311,N_38218,N_38091);
and U38312 (N_38312,N_38093,N_38180);
and U38313 (N_38313,N_38097,N_38147);
xnor U38314 (N_38314,N_38133,N_38074);
or U38315 (N_38315,N_38211,N_38044);
xor U38316 (N_38316,N_38011,N_38095);
or U38317 (N_38317,N_38090,N_38015);
nor U38318 (N_38318,N_38146,N_38200);
nand U38319 (N_38319,N_38154,N_38086);
nand U38320 (N_38320,N_38111,N_38023);
nor U38321 (N_38321,N_38144,N_38195);
and U38322 (N_38322,N_38101,N_38051);
nor U38323 (N_38323,N_38234,N_38013);
or U38324 (N_38324,N_38194,N_38237);
nor U38325 (N_38325,N_38008,N_38224);
xor U38326 (N_38326,N_38071,N_38105);
and U38327 (N_38327,N_38119,N_38116);
or U38328 (N_38328,N_38131,N_38245);
nor U38329 (N_38329,N_38120,N_38026);
or U38330 (N_38330,N_38229,N_38115);
or U38331 (N_38331,N_38207,N_38032);
and U38332 (N_38332,N_38175,N_38068);
nand U38333 (N_38333,N_38052,N_38241);
nor U38334 (N_38334,N_38050,N_38088);
xnor U38335 (N_38335,N_38004,N_38021);
nor U38336 (N_38336,N_38161,N_38053);
nor U38337 (N_38337,N_38162,N_38190);
xnor U38338 (N_38338,N_38137,N_38043);
xor U38339 (N_38339,N_38239,N_38005);
xnor U38340 (N_38340,N_38127,N_38110);
and U38341 (N_38341,N_38142,N_38104);
nor U38342 (N_38342,N_38014,N_38046);
and U38343 (N_38343,N_38036,N_38012);
and U38344 (N_38344,N_38163,N_38155);
and U38345 (N_38345,N_38141,N_38170);
or U38346 (N_38346,N_38143,N_38058);
xnor U38347 (N_38347,N_38034,N_38033);
nor U38348 (N_38348,N_38057,N_38019);
nand U38349 (N_38349,N_38156,N_38214);
and U38350 (N_38350,N_38122,N_38184);
xnor U38351 (N_38351,N_38040,N_38031);
and U38352 (N_38352,N_38010,N_38166);
xor U38353 (N_38353,N_38151,N_38176);
nand U38354 (N_38354,N_38212,N_38060);
and U38355 (N_38355,N_38167,N_38024);
xnor U38356 (N_38356,N_38029,N_38192);
and U38357 (N_38357,N_38066,N_38114);
nand U38358 (N_38358,N_38065,N_38204);
and U38359 (N_38359,N_38198,N_38164);
nand U38360 (N_38360,N_38056,N_38109);
and U38361 (N_38361,N_38222,N_38174);
nor U38362 (N_38362,N_38181,N_38070);
nor U38363 (N_38363,N_38006,N_38055);
or U38364 (N_38364,N_38098,N_38078);
or U38365 (N_38365,N_38072,N_38129);
nor U38366 (N_38366,N_38007,N_38169);
or U38367 (N_38367,N_38138,N_38126);
xor U38368 (N_38368,N_38082,N_38228);
nor U38369 (N_38369,N_38150,N_38100);
nand U38370 (N_38370,N_38000,N_38140);
and U38371 (N_38371,N_38094,N_38219);
or U38372 (N_38372,N_38069,N_38191);
nor U38373 (N_38373,N_38206,N_38217);
or U38374 (N_38374,N_38233,N_38087);
nand U38375 (N_38375,N_38121,N_38019);
or U38376 (N_38376,N_38092,N_38223);
xor U38377 (N_38377,N_38033,N_38115);
and U38378 (N_38378,N_38249,N_38199);
xor U38379 (N_38379,N_38110,N_38236);
nand U38380 (N_38380,N_38084,N_38142);
nor U38381 (N_38381,N_38145,N_38131);
xnor U38382 (N_38382,N_38129,N_38056);
and U38383 (N_38383,N_38057,N_38193);
nand U38384 (N_38384,N_38087,N_38147);
nor U38385 (N_38385,N_38238,N_38184);
nor U38386 (N_38386,N_38197,N_38161);
nand U38387 (N_38387,N_38170,N_38200);
and U38388 (N_38388,N_38211,N_38032);
nand U38389 (N_38389,N_38057,N_38024);
xnor U38390 (N_38390,N_38022,N_38051);
nand U38391 (N_38391,N_38016,N_38115);
and U38392 (N_38392,N_38056,N_38051);
nor U38393 (N_38393,N_38050,N_38013);
or U38394 (N_38394,N_38069,N_38242);
xor U38395 (N_38395,N_38131,N_38019);
nand U38396 (N_38396,N_38141,N_38136);
nand U38397 (N_38397,N_38230,N_38035);
xnor U38398 (N_38398,N_38017,N_38103);
and U38399 (N_38399,N_38069,N_38024);
nand U38400 (N_38400,N_38059,N_38043);
nor U38401 (N_38401,N_38020,N_38074);
and U38402 (N_38402,N_38023,N_38210);
nand U38403 (N_38403,N_38193,N_38195);
nor U38404 (N_38404,N_38165,N_38177);
and U38405 (N_38405,N_38023,N_38169);
and U38406 (N_38406,N_38059,N_38217);
nor U38407 (N_38407,N_38091,N_38142);
and U38408 (N_38408,N_38146,N_38000);
nor U38409 (N_38409,N_38203,N_38172);
nand U38410 (N_38410,N_38173,N_38184);
or U38411 (N_38411,N_38099,N_38000);
xnor U38412 (N_38412,N_38105,N_38011);
nor U38413 (N_38413,N_38030,N_38194);
nand U38414 (N_38414,N_38114,N_38021);
and U38415 (N_38415,N_38067,N_38045);
nand U38416 (N_38416,N_38068,N_38153);
nor U38417 (N_38417,N_38077,N_38211);
nor U38418 (N_38418,N_38062,N_38163);
or U38419 (N_38419,N_38075,N_38026);
xor U38420 (N_38420,N_38203,N_38102);
nor U38421 (N_38421,N_38241,N_38224);
nor U38422 (N_38422,N_38140,N_38139);
xnor U38423 (N_38423,N_38042,N_38249);
nor U38424 (N_38424,N_38225,N_38159);
nor U38425 (N_38425,N_38204,N_38052);
nand U38426 (N_38426,N_38059,N_38027);
nor U38427 (N_38427,N_38139,N_38023);
xnor U38428 (N_38428,N_38178,N_38209);
or U38429 (N_38429,N_38089,N_38130);
nand U38430 (N_38430,N_38028,N_38140);
nor U38431 (N_38431,N_38034,N_38025);
and U38432 (N_38432,N_38040,N_38010);
or U38433 (N_38433,N_38031,N_38097);
xnor U38434 (N_38434,N_38098,N_38073);
xnor U38435 (N_38435,N_38007,N_38217);
and U38436 (N_38436,N_38118,N_38179);
or U38437 (N_38437,N_38073,N_38008);
and U38438 (N_38438,N_38175,N_38219);
and U38439 (N_38439,N_38105,N_38126);
and U38440 (N_38440,N_38009,N_38129);
xnor U38441 (N_38441,N_38047,N_38231);
nand U38442 (N_38442,N_38193,N_38227);
xnor U38443 (N_38443,N_38153,N_38195);
and U38444 (N_38444,N_38078,N_38217);
and U38445 (N_38445,N_38024,N_38142);
and U38446 (N_38446,N_38101,N_38197);
and U38447 (N_38447,N_38244,N_38200);
or U38448 (N_38448,N_38046,N_38047);
and U38449 (N_38449,N_38103,N_38201);
and U38450 (N_38450,N_38043,N_38104);
xnor U38451 (N_38451,N_38201,N_38175);
nor U38452 (N_38452,N_38037,N_38187);
nor U38453 (N_38453,N_38014,N_38049);
nand U38454 (N_38454,N_38244,N_38183);
or U38455 (N_38455,N_38124,N_38204);
nand U38456 (N_38456,N_38037,N_38179);
or U38457 (N_38457,N_38206,N_38239);
and U38458 (N_38458,N_38199,N_38122);
xnor U38459 (N_38459,N_38136,N_38058);
nor U38460 (N_38460,N_38166,N_38180);
xor U38461 (N_38461,N_38017,N_38041);
nor U38462 (N_38462,N_38044,N_38024);
or U38463 (N_38463,N_38084,N_38137);
xor U38464 (N_38464,N_38015,N_38161);
or U38465 (N_38465,N_38248,N_38235);
nor U38466 (N_38466,N_38184,N_38032);
nor U38467 (N_38467,N_38233,N_38084);
nand U38468 (N_38468,N_38160,N_38063);
xor U38469 (N_38469,N_38150,N_38162);
nand U38470 (N_38470,N_38102,N_38221);
xor U38471 (N_38471,N_38172,N_38091);
and U38472 (N_38472,N_38071,N_38095);
or U38473 (N_38473,N_38225,N_38053);
nand U38474 (N_38474,N_38112,N_38003);
xnor U38475 (N_38475,N_38157,N_38056);
nor U38476 (N_38476,N_38001,N_38071);
and U38477 (N_38477,N_38230,N_38107);
or U38478 (N_38478,N_38152,N_38103);
nand U38479 (N_38479,N_38238,N_38018);
nand U38480 (N_38480,N_38068,N_38049);
xor U38481 (N_38481,N_38207,N_38065);
and U38482 (N_38482,N_38173,N_38165);
nand U38483 (N_38483,N_38195,N_38145);
nand U38484 (N_38484,N_38237,N_38201);
or U38485 (N_38485,N_38115,N_38170);
xnor U38486 (N_38486,N_38197,N_38038);
nand U38487 (N_38487,N_38016,N_38199);
nand U38488 (N_38488,N_38163,N_38106);
or U38489 (N_38489,N_38237,N_38216);
or U38490 (N_38490,N_38218,N_38024);
or U38491 (N_38491,N_38051,N_38077);
or U38492 (N_38492,N_38051,N_38098);
and U38493 (N_38493,N_38069,N_38134);
xnor U38494 (N_38494,N_38025,N_38106);
xor U38495 (N_38495,N_38012,N_38068);
and U38496 (N_38496,N_38032,N_38120);
xor U38497 (N_38497,N_38093,N_38201);
nor U38498 (N_38498,N_38155,N_38180);
or U38499 (N_38499,N_38186,N_38235);
nor U38500 (N_38500,N_38335,N_38378);
nor U38501 (N_38501,N_38443,N_38267);
xor U38502 (N_38502,N_38453,N_38421);
nor U38503 (N_38503,N_38465,N_38423);
nor U38504 (N_38504,N_38276,N_38445);
nor U38505 (N_38505,N_38367,N_38451);
xnor U38506 (N_38506,N_38337,N_38417);
nand U38507 (N_38507,N_38481,N_38472);
nor U38508 (N_38508,N_38455,N_38459);
or U38509 (N_38509,N_38364,N_38292);
and U38510 (N_38510,N_38313,N_38409);
nand U38511 (N_38511,N_38374,N_38330);
and U38512 (N_38512,N_38268,N_38482);
and U38513 (N_38513,N_38376,N_38258);
nor U38514 (N_38514,N_38396,N_38473);
or U38515 (N_38515,N_38355,N_38408);
nor U38516 (N_38516,N_38478,N_38372);
or U38517 (N_38517,N_38283,N_38363);
nand U38518 (N_38518,N_38358,N_38306);
or U38519 (N_38519,N_38256,N_38407);
or U38520 (N_38520,N_38304,N_38395);
and U38521 (N_38521,N_38490,N_38498);
or U38522 (N_38522,N_38323,N_38348);
nor U38523 (N_38523,N_38264,N_38310);
nor U38524 (N_38524,N_38270,N_38334);
nand U38525 (N_38525,N_38415,N_38432);
or U38526 (N_38526,N_38320,N_38491);
or U38527 (N_38527,N_38300,N_38377);
and U38528 (N_38528,N_38286,N_38379);
nand U38529 (N_38529,N_38279,N_38383);
or U38530 (N_38530,N_38312,N_38289);
nor U38531 (N_38531,N_38251,N_38483);
nand U38532 (N_38532,N_38284,N_38365);
or U38533 (N_38533,N_38303,N_38499);
nor U38534 (N_38534,N_38280,N_38275);
or U38535 (N_38535,N_38281,N_38411);
xor U38536 (N_38536,N_38413,N_38393);
nor U38537 (N_38537,N_38366,N_38474);
and U38538 (N_38538,N_38344,N_38288);
nor U38539 (N_38539,N_38476,N_38360);
nor U38540 (N_38540,N_38406,N_38349);
nand U38541 (N_38541,N_38397,N_38311);
nand U38542 (N_38542,N_38353,N_38308);
xor U38543 (N_38543,N_38250,N_38471);
nand U38544 (N_38544,N_38296,N_38361);
nand U38545 (N_38545,N_38368,N_38257);
or U38546 (N_38546,N_38418,N_38391);
or U38547 (N_38547,N_38392,N_38394);
xor U38548 (N_38548,N_38357,N_38435);
nand U38549 (N_38549,N_38362,N_38430);
xnor U38550 (N_38550,N_38429,N_38318);
and U38551 (N_38551,N_38266,N_38354);
and U38552 (N_38552,N_38384,N_38433);
and U38553 (N_38553,N_38326,N_38340);
xor U38554 (N_38554,N_38262,N_38420);
or U38555 (N_38555,N_38446,N_38449);
nor U38556 (N_38556,N_38448,N_38437);
nor U38557 (N_38557,N_38381,N_38434);
nand U38558 (N_38558,N_38333,N_38475);
and U38559 (N_38559,N_38489,N_38271);
or U38560 (N_38560,N_38464,N_38410);
nand U38561 (N_38561,N_38496,N_38497);
nor U38562 (N_38562,N_38338,N_38468);
xor U38563 (N_38563,N_38439,N_38467);
xor U38564 (N_38564,N_38398,N_38359);
nor U38565 (N_38565,N_38322,N_38371);
or U38566 (N_38566,N_38466,N_38382);
or U38567 (N_38567,N_38427,N_38404);
nor U38568 (N_38568,N_38331,N_38375);
or U38569 (N_38569,N_38454,N_38492);
nor U38570 (N_38570,N_38325,N_38493);
nand U38571 (N_38571,N_38324,N_38255);
nor U38572 (N_38572,N_38463,N_38419);
nor U38573 (N_38573,N_38297,N_38317);
nor U38574 (N_38574,N_38462,N_38412);
or U38575 (N_38575,N_38336,N_38380);
nand U38576 (N_38576,N_38345,N_38461);
nor U38577 (N_38577,N_38253,N_38456);
nand U38578 (N_38578,N_38477,N_38480);
nor U38579 (N_38579,N_38431,N_38261);
nor U38580 (N_38580,N_38401,N_38469);
nor U38581 (N_38581,N_38351,N_38341);
and U38582 (N_38582,N_38342,N_38263);
nor U38583 (N_38583,N_38479,N_38450);
nor U38584 (N_38584,N_38295,N_38447);
nand U38585 (N_38585,N_38441,N_38287);
and U38586 (N_38586,N_38347,N_38422);
and U38587 (N_38587,N_38316,N_38329);
nor U38588 (N_38588,N_38350,N_38259);
or U38589 (N_38589,N_38302,N_38402);
or U38590 (N_38590,N_38301,N_38485);
xnor U38591 (N_38591,N_38274,N_38272);
xnor U38592 (N_38592,N_38315,N_38457);
or U38593 (N_38593,N_38385,N_38495);
xor U38594 (N_38594,N_38440,N_38307);
and U38595 (N_38595,N_38314,N_38369);
nor U38596 (N_38596,N_38282,N_38319);
and U38597 (N_38597,N_38332,N_38400);
xnor U38598 (N_38598,N_38327,N_38339);
and U38599 (N_38599,N_38290,N_38277);
nor U38600 (N_38600,N_38273,N_38386);
and U38601 (N_38601,N_38278,N_38298);
and U38602 (N_38602,N_38438,N_38444);
or U38603 (N_38603,N_38414,N_38425);
or U38604 (N_38604,N_38484,N_38254);
and U38605 (N_38605,N_38424,N_38426);
nor U38606 (N_38606,N_38486,N_38388);
and U38607 (N_38607,N_38321,N_38293);
xor U38608 (N_38608,N_38265,N_38436);
nand U38609 (N_38609,N_38269,N_38405);
or U38610 (N_38610,N_38389,N_38309);
or U38611 (N_38611,N_38260,N_38487);
nor U38612 (N_38612,N_38399,N_38470);
or U38613 (N_38613,N_38416,N_38458);
xor U38614 (N_38614,N_38328,N_38488);
xor U38615 (N_38615,N_38387,N_38299);
nor U38616 (N_38616,N_38343,N_38346);
or U38617 (N_38617,N_38305,N_38291);
and U38618 (N_38618,N_38370,N_38494);
xor U38619 (N_38619,N_38294,N_38373);
or U38620 (N_38620,N_38460,N_38428);
nor U38621 (N_38621,N_38403,N_38356);
nand U38622 (N_38622,N_38442,N_38452);
and U38623 (N_38623,N_38352,N_38285);
nand U38624 (N_38624,N_38390,N_38252);
and U38625 (N_38625,N_38285,N_38442);
xnor U38626 (N_38626,N_38464,N_38471);
nand U38627 (N_38627,N_38317,N_38330);
nor U38628 (N_38628,N_38301,N_38394);
and U38629 (N_38629,N_38453,N_38445);
nor U38630 (N_38630,N_38366,N_38354);
nand U38631 (N_38631,N_38473,N_38354);
nor U38632 (N_38632,N_38461,N_38328);
or U38633 (N_38633,N_38496,N_38410);
and U38634 (N_38634,N_38288,N_38471);
nor U38635 (N_38635,N_38361,N_38388);
or U38636 (N_38636,N_38479,N_38283);
xnor U38637 (N_38637,N_38250,N_38268);
xor U38638 (N_38638,N_38475,N_38262);
xnor U38639 (N_38639,N_38434,N_38471);
and U38640 (N_38640,N_38422,N_38379);
and U38641 (N_38641,N_38276,N_38419);
xor U38642 (N_38642,N_38472,N_38379);
or U38643 (N_38643,N_38428,N_38280);
nor U38644 (N_38644,N_38283,N_38421);
nor U38645 (N_38645,N_38418,N_38415);
or U38646 (N_38646,N_38431,N_38393);
nor U38647 (N_38647,N_38427,N_38498);
and U38648 (N_38648,N_38457,N_38361);
xnor U38649 (N_38649,N_38468,N_38431);
nand U38650 (N_38650,N_38381,N_38393);
xor U38651 (N_38651,N_38293,N_38374);
xor U38652 (N_38652,N_38275,N_38405);
nor U38653 (N_38653,N_38403,N_38471);
nor U38654 (N_38654,N_38371,N_38379);
xor U38655 (N_38655,N_38270,N_38420);
or U38656 (N_38656,N_38398,N_38415);
xor U38657 (N_38657,N_38265,N_38274);
and U38658 (N_38658,N_38396,N_38418);
nor U38659 (N_38659,N_38460,N_38419);
and U38660 (N_38660,N_38478,N_38371);
or U38661 (N_38661,N_38275,N_38417);
or U38662 (N_38662,N_38293,N_38487);
nand U38663 (N_38663,N_38419,N_38432);
nand U38664 (N_38664,N_38307,N_38437);
xnor U38665 (N_38665,N_38322,N_38492);
or U38666 (N_38666,N_38324,N_38317);
nor U38667 (N_38667,N_38380,N_38303);
xor U38668 (N_38668,N_38251,N_38264);
or U38669 (N_38669,N_38262,N_38350);
and U38670 (N_38670,N_38386,N_38473);
nor U38671 (N_38671,N_38376,N_38437);
nand U38672 (N_38672,N_38399,N_38401);
and U38673 (N_38673,N_38414,N_38435);
nand U38674 (N_38674,N_38271,N_38438);
xnor U38675 (N_38675,N_38458,N_38330);
xnor U38676 (N_38676,N_38484,N_38297);
xor U38677 (N_38677,N_38489,N_38460);
or U38678 (N_38678,N_38333,N_38467);
nor U38679 (N_38679,N_38385,N_38440);
nand U38680 (N_38680,N_38488,N_38449);
nand U38681 (N_38681,N_38469,N_38286);
nand U38682 (N_38682,N_38406,N_38264);
and U38683 (N_38683,N_38274,N_38336);
xnor U38684 (N_38684,N_38364,N_38373);
or U38685 (N_38685,N_38361,N_38434);
nor U38686 (N_38686,N_38256,N_38318);
and U38687 (N_38687,N_38482,N_38488);
and U38688 (N_38688,N_38341,N_38407);
xor U38689 (N_38689,N_38313,N_38262);
nand U38690 (N_38690,N_38306,N_38366);
and U38691 (N_38691,N_38440,N_38287);
nand U38692 (N_38692,N_38317,N_38451);
nor U38693 (N_38693,N_38293,N_38471);
nor U38694 (N_38694,N_38316,N_38434);
nor U38695 (N_38695,N_38328,N_38452);
xnor U38696 (N_38696,N_38368,N_38484);
and U38697 (N_38697,N_38403,N_38259);
and U38698 (N_38698,N_38490,N_38464);
and U38699 (N_38699,N_38448,N_38413);
or U38700 (N_38700,N_38468,N_38453);
or U38701 (N_38701,N_38422,N_38391);
and U38702 (N_38702,N_38342,N_38399);
xnor U38703 (N_38703,N_38390,N_38361);
and U38704 (N_38704,N_38489,N_38426);
xnor U38705 (N_38705,N_38307,N_38495);
or U38706 (N_38706,N_38382,N_38455);
xnor U38707 (N_38707,N_38442,N_38383);
nand U38708 (N_38708,N_38370,N_38353);
or U38709 (N_38709,N_38483,N_38486);
xor U38710 (N_38710,N_38353,N_38294);
nand U38711 (N_38711,N_38416,N_38466);
nor U38712 (N_38712,N_38265,N_38387);
nor U38713 (N_38713,N_38471,N_38400);
nand U38714 (N_38714,N_38263,N_38254);
nand U38715 (N_38715,N_38348,N_38469);
nand U38716 (N_38716,N_38318,N_38307);
or U38717 (N_38717,N_38389,N_38491);
and U38718 (N_38718,N_38436,N_38356);
or U38719 (N_38719,N_38408,N_38315);
xnor U38720 (N_38720,N_38283,N_38437);
and U38721 (N_38721,N_38394,N_38271);
and U38722 (N_38722,N_38428,N_38476);
and U38723 (N_38723,N_38369,N_38410);
or U38724 (N_38724,N_38481,N_38325);
and U38725 (N_38725,N_38450,N_38495);
nand U38726 (N_38726,N_38492,N_38490);
nand U38727 (N_38727,N_38422,N_38357);
xnor U38728 (N_38728,N_38452,N_38476);
xnor U38729 (N_38729,N_38346,N_38389);
or U38730 (N_38730,N_38370,N_38323);
and U38731 (N_38731,N_38455,N_38343);
and U38732 (N_38732,N_38327,N_38451);
or U38733 (N_38733,N_38391,N_38386);
or U38734 (N_38734,N_38266,N_38411);
nor U38735 (N_38735,N_38390,N_38394);
or U38736 (N_38736,N_38261,N_38318);
nor U38737 (N_38737,N_38432,N_38282);
and U38738 (N_38738,N_38372,N_38345);
or U38739 (N_38739,N_38464,N_38375);
or U38740 (N_38740,N_38381,N_38404);
nand U38741 (N_38741,N_38250,N_38374);
and U38742 (N_38742,N_38359,N_38447);
nor U38743 (N_38743,N_38375,N_38419);
nand U38744 (N_38744,N_38302,N_38350);
and U38745 (N_38745,N_38424,N_38468);
nor U38746 (N_38746,N_38325,N_38346);
nor U38747 (N_38747,N_38269,N_38479);
or U38748 (N_38748,N_38495,N_38442);
nor U38749 (N_38749,N_38268,N_38370);
and U38750 (N_38750,N_38725,N_38591);
xnor U38751 (N_38751,N_38531,N_38545);
nor U38752 (N_38752,N_38730,N_38714);
xor U38753 (N_38753,N_38561,N_38580);
nand U38754 (N_38754,N_38676,N_38681);
xnor U38755 (N_38755,N_38719,N_38721);
nand U38756 (N_38756,N_38646,N_38550);
nor U38757 (N_38757,N_38657,N_38606);
xor U38758 (N_38758,N_38678,N_38524);
xor U38759 (N_38759,N_38510,N_38648);
nor U38760 (N_38760,N_38549,N_38604);
and U38761 (N_38761,N_38644,N_38742);
or U38762 (N_38762,N_38512,N_38519);
or U38763 (N_38763,N_38669,N_38611);
nor U38764 (N_38764,N_38596,N_38692);
nand U38765 (N_38765,N_38502,N_38666);
and U38766 (N_38766,N_38699,N_38553);
nor U38767 (N_38767,N_38564,N_38621);
or U38768 (N_38768,N_38537,N_38680);
nor U38769 (N_38769,N_38641,N_38506);
xor U38770 (N_38770,N_38533,N_38636);
or U38771 (N_38771,N_38590,N_38557);
xor U38772 (N_38772,N_38707,N_38713);
xor U38773 (N_38773,N_38541,N_38527);
xor U38774 (N_38774,N_38677,N_38691);
and U38775 (N_38775,N_38602,N_38736);
nand U38776 (N_38776,N_38599,N_38538);
and U38777 (N_38777,N_38521,N_38662);
nand U38778 (N_38778,N_38608,N_38740);
nand U38779 (N_38779,N_38555,N_38560);
or U38780 (N_38780,N_38520,N_38695);
nor U38781 (N_38781,N_38569,N_38552);
nor U38782 (N_38782,N_38565,N_38503);
and U38783 (N_38783,N_38637,N_38624);
and U38784 (N_38784,N_38747,N_38743);
nor U38785 (N_38785,N_38661,N_38528);
nand U38786 (N_38786,N_38544,N_38696);
or U38787 (N_38787,N_38732,N_38693);
xor U38788 (N_38788,N_38612,N_38532);
xnor U38789 (N_38789,N_38704,N_38711);
xnor U38790 (N_38790,N_38749,N_38726);
nand U38791 (N_38791,N_38650,N_38507);
and U38792 (N_38792,N_38735,N_38586);
xnor U38793 (N_38793,N_38543,N_38744);
and U38794 (N_38794,N_38523,N_38582);
or U38795 (N_38795,N_38578,N_38595);
and U38796 (N_38796,N_38518,N_38654);
or U38797 (N_38797,N_38605,N_38665);
nand U38798 (N_38798,N_38597,N_38628);
or U38799 (N_38799,N_38514,N_38540);
or U38800 (N_38800,N_38500,N_38640);
xnor U38801 (N_38801,N_38664,N_38535);
nand U38802 (N_38802,N_38504,N_38575);
nor U38803 (N_38803,N_38568,N_38690);
or U38804 (N_38804,N_38708,N_38579);
nand U38805 (N_38805,N_38513,N_38618);
and U38806 (N_38806,N_38728,N_38516);
nor U38807 (N_38807,N_38505,N_38729);
xor U38808 (N_38808,N_38694,N_38584);
and U38809 (N_38809,N_38589,N_38656);
xor U38810 (N_38810,N_38558,N_38703);
nor U38811 (N_38811,N_38702,N_38610);
nand U38812 (N_38812,N_38614,N_38723);
or U38813 (N_38813,N_38551,N_38734);
nand U38814 (N_38814,N_38609,N_38688);
or U38815 (N_38815,N_38554,N_38642);
nor U38816 (N_38816,N_38556,N_38745);
nor U38817 (N_38817,N_38718,N_38722);
and U38818 (N_38818,N_38689,N_38567);
nand U38819 (N_38819,N_38583,N_38570);
xor U38820 (N_38820,N_38737,N_38630);
and U38821 (N_38821,N_38660,N_38594);
xnor U38822 (N_38822,N_38668,N_38629);
or U38823 (N_38823,N_38542,N_38673);
xnor U38824 (N_38824,N_38539,N_38515);
or U38825 (N_38825,N_38731,N_38546);
nor U38826 (N_38826,N_38717,N_38577);
xor U38827 (N_38827,N_38563,N_38600);
nand U38828 (N_38828,N_38571,N_38639);
xnor U38829 (N_38829,N_38508,N_38727);
and U38830 (N_38830,N_38572,N_38529);
xnor U38831 (N_38831,N_38682,N_38585);
xnor U38832 (N_38832,N_38525,N_38622);
xor U38833 (N_38833,N_38653,N_38670);
and U38834 (N_38834,N_38709,N_38626);
xor U38835 (N_38835,N_38672,N_38562);
and U38836 (N_38836,N_38739,N_38526);
xor U38837 (N_38837,N_38593,N_38603);
or U38838 (N_38838,N_38566,N_38697);
nand U38839 (N_38839,N_38638,N_38733);
nor U38840 (N_38840,N_38592,N_38633);
or U38841 (N_38841,N_38511,N_38655);
and U38842 (N_38842,N_38679,N_38635);
nand U38843 (N_38843,N_38522,N_38675);
or U38844 (N_38844,N_38616,N_38746);
xor U38845 (N_38845,N_38617,N_38643);
and U38846 (N_38846,N_38705,N_38738);
xnor U38847 (N_38847,N_38509,N_38598);
xnor U38848 (N_38848,N_38517,N_38620);
or U38849 (N_38849,N_38651,N_38501);
xor U38850 (N_38850,N_38698,N_38659);
xnor U38851 (N_38851,N_38701,N_38674);
xnor U38852 (N_38852,N_38574,N_38536);
nor U38853 (N_38853,N_38685,N_38631);
nand U38854 (N_38854,N_38647,N_38671);
nand U38855 (N_38855,N_38724,N_38615);
or U38856 (N_38856,N_38625,N_38613);
xnor U38857 (N_38857,N_38715,N_38741);
nand U38858 (N_38858,N_38683,N_38658);
nor U38859 (N_38859,N_38706,N_38710);
nor U38860 (N_38860,N_38720,N_38700);
xnor U38861 (N_38861,N_38619,N_38601);
xor U38862 (N_38862,N_38748,N_38587);
and U38863 (N_38863,N_38581,N_38627);
nor U38864 (N_38864,N_38712,N_38686);
nor U38865 (N_38865,N_38652,N_38559);
nor U38866 (N_38866,N_38573,N_38645);
nor U38867 (N_38867,N_38634,N_38534);
xnor U38868 (N_38868,N_38684,N_38649);
nand U38869 (N_38869,N_38667,N_38663);
and U38870 (N_38870,N_38632,N_38687);
nand U38871 (N_38871,N_38530,N_38576);
and U38872 (N_38872,N_38588,N_38548);
or U38873 (N_38873,N_38607,N_38716);
or U38874 (N_38874,N_38547,N_38623);
or U38875 (N_38875,N_38726,N_38700);
nand U38876 (N_38876,N_38631,N_38684);
nor U38877 (N_38877,N_38502,N_38554);
nand U38878 (N_38878,N_38531,N_38621);
xnor U38879 (N_38879,N_38661,N_38641);
and U38880 (N_38880,N_38622,N_38702);
or U38881 (N_38881,N_38521,N_38597);
or U38882 (N_38882,N_38670,N_38553);
nor U38883 (N_38883,N_38532,N_38611);
or U38884 (N_38884,N_38658,N_38544);
xor U38885 (N_38885,N_38747,N_38594);
or U38886 (N_38886,N_38652,N_38662);
xor U38887 (N_38887,N_38630,N_38582);
xnor U38888 (N_38888,N_38733,N_38723);
and U38889 (N_38889,N_38604,N_38563);
nor U38890 (N_38890,N_38681,N_38663);
nand U38891 (N_38891,N_38654,N_38660);
xor U38892 (N_38892,N_38614,N_38500);
xor U38893 (N_38893,N_38666,N_38707);
nor U38894 (N_38894,N_38585,N_38727);
and U38895 (N_38895,N_38504,N_38552);
xor U38896 (N_38896,N_38719,N_38672);
nand U38897 (N_38897,N_38561,N_38505);
xnor U38898 (N_38898,N_38713,N_38606);
nand U38899 (N_38899,N_38592,N_38636);
nand U38900 (N_38900,N_38674,N_38573);
and U38901 (N_38901,N_38737,N_38531);
nand U38902 (N_38902,N_38588,N_38586);
or U38903 (N_38903,N_38526,N_38614);
nor U38904 (N_38904,N_38550,N_38724);
nor U38905 (N_38905,N_38673,N_38539);
or U38906 (N_38906,N_38531,N_38588);
and U38907 (N_38907,N_38576,N_38693);
and U38908 (N_38908,N_38705,N_38718);
and U38909 (N_38909,N_38540,N_38522);
and U38910 (N_38910,N_38699,N_38732);
nor U38911 (N_38911,N_38503,N_38585);
nor U38912 (N_38912,N_38517,N_38543);
nor U38913 (N_38913,N_38536,N_38586);
nor U38914 (N_38914,N_38587,N_38606);
nor U38915 (N_38915,N_38595,N_38700);
or U38916 (N_38916,N_38570,N_38532);
and U38917 (N_38917,N_38697,N_38650);
nand U38918 (N_38918,N_38606,N_38531);
and U38919 (N_38919,N_38723,N_38669);
or U38920 (N_38920,N_38703,N_38676);
xnor U38921 (N_38921,N_38508,N_38634);
nand U38922 (N_38922,N_38629,N_38602);
xor U38923 (N_38923,N_38527,N_38520);
xnor U38924 (N_38924,N_38638,N_38549);
and U38925 (N_38925,N_38544,N_38581);
nand U38926 (N_38926,N_38578,N_38730);
nor U38927 (N_38927,N_38651,N_38649);
nor U38928 (N_38928,N_38602,N_38626);
nor U38929 (N_38929,N_38634,N_38510);
nor U38930 (N_38930,N_38649,N_38704);
nor U38931 (N_38931,N_38603,N_38724);
nor U38932 (N_38932,N_38698,N_38656);
or U38933 (N_38933,N_38616,N_38598);
xor U38934 (N_38934,N_38676,N_38748);
and U38935 (N_38935,N_38561,N_38576);
nor U38936 (N_38936,N_38663,N_38531);
xnor U38937 (N_38937,N_38614,N_38512);
xnor U38938 (N_38938,N_38573,N_38742);
nand U38939 (N_38939,N_38655,N_38694);
nor U38940 (N_38940,N_38735,N_38524);
or U38941 (N_38941,N_38707,N_38511);
nor U38942 (N_38942,N_38500,N_38591);
nor U38943 (N_38943,N_38723,N_38663);
or U38944 (N_38944,N_38669,N_38698);
nand U38945 (N_38945,N_38724,N_38533);
nand U38946 (N_38946,N_38712,N_38739);
and U38947 (N_38947,N_38616,N_38619);
nor U38948 (N_38948,N_38589,N_38713);
nand U38949 (N_38949,N_38545,N_38674);
nor U38950 (N_38950,N_38674,N_38500);
nand U38951 (N_38951,N_38747,N_38742);
and U38952 (N_38952,N_38716,N_38657);
nand U38953 (N_38953,N_38660,N_38714);
xnor U38954 (N_38954,N_38508,N_38562);
and U38955 (N_38955,N_38610,N_38527);
and U38956 (N_38956,N_38697,N_38593);
xnor U38957 (N_38957,N_38712,N_38565);
nand U38958 (N_38958,N_38532,N_38522);
nand U38959 (N_38959,N_38731,N_38654);
or U38960 (N_38960,N_38610,N_38641);
xnor U38961 (N_38961,N_38575,N_38580);
nand U38962 (N_38962,N_38577,N_38716);
nor U38963 (N_38963,N_38551,N_38562);
and U38964 (N_38964,N_38742,N_38684);
xor U38965 (N_38965,N_38516,N_38588);
or U38966 (N_38966,N_38578,N_38508);
and U38967 (N_38967,N_38510,N_38560);
or U38968 (N_38968,N_38609,N_38636);
or U38969 (N_38969,N_38656,N_38509);
nand U38970 (N_38970,N_38712,N_38528);
nor U38971 (N_38971,N_38564,N_38528);
and U38972 (N_38972,N_38715,N_38558);
xor U38973 (N_38973,N_38533,N_38672);
nor U38974 (N_38974,N_38525,N_38696);
or U38975 (N_38975,N_38657,N_38667);
and U38976 (N_38976,N_38525,N_38621);
nand U38977 (N_38977,N_38704,N_38512);
nand U38978 (N_38978,N_38678,N_38630);
or U38979 (N_38979,N_38686,N_38566);
nor U38980 (N_38980,N_38555,N_38713);
or U38981 (N_38981,N_38734,N_38630);
and U38982 (N_38982,N_38627,N_38595);
xnor U38983 (N_38983,N_38723,N_38655);
and U38984 (N_38984,N_38651,N_38600);
nand U38985 (N_38985,N_38552,N_38549);
nand U38986 (N_38986,N_38538,N_38603);
nand U38987 (N_38987,N_38511,N_38569);
nand U38988 (N_38988,N_38606,N_38584);
xnor U38989 (N_38989,N_38744,N_38517);
nand U38990 (N_38990,N_38523,N_38588);
and U38991 (N_38991,N_38529,N_38628);
nor U38992 (N_38992,N_38669,N_38515);
nor U38993 (N_38993,N_38615,N_38652);
xor U38994 (N_38994,N_38736,N_38672);
and U38995 (N_38995,N_38739,N_38554);
and U38996 (N_38996,N_38745,N_38602);
xnor U38997 (N_38997,N_38734,N_38612);
nor U38998 (N_38998,N_38733,N_38543);
and U38999 (N_38999,N_38722,N_38643);
and U39000 (N_39000,N_38863,N_38843);
xnor U39001 (N_39001,N_38799,N_38865);
nor U39002 (N_39002,N_38876,N_38870);
and U39003 (N_39003,N_38976,N_38925);
nand U39004 (N_39004,N_38827,N_38834);
xnor U39005 (N_39005,N_38817,N_38983);
nand U39006 (N_39006,N_38883,N_38967);
nand U39007 (N_39007,N_38982,N_38949);
nand U39008 (N_39008,N_38904,N_38791);
xor U39009 (N_39009,N_38935,N_38936);
nand U39010 (N_39010,N_38898,N_38897);
nand U39011 (N_39011,N_38909,N_38836);
nor U39012 (N_39012,N_38813,N_38758);
or U39013 (N_39013,N_38889,N_38753);
and U39014 (N_39014,N_38990,N_38939);
nand U39015 (N_39015,N_38933,N_38912);
nand U39016 (N_39016,N_38916,N_38964);
or U39017 (N_39017,N_38954,N_38968);
and U39018 (N_39018,N_38887,N_38953);
and U39019 (N_39019,N_38807,N_38772);
and U39020 (N_39020,N_38833,N_38891);
nor U39021 (N_39021,N_38784,N_38970);
and U39022 (N_39022,N_38929,N_38989);
or U39023 (N_39023,N_38960,N_38957);
and U39024 (N_39024,N_38795,N_38878);
nor U39025 (N_39025,N_38808,N_38906);
nor U39026 (N_39026,N_38852,N_38835);
nor U39027 (N_39027,N_38928,N_38862);
or U39028 (N_39028,N_38905,N_38775);
or U39029 (N_39029,N_38941,N_38776);
or U39030 (N_39030,N_38815,N_38944);
xnor U39031 (N_39031,N_38942,N_38850);
xnor U39032 (N_39032,N_38771,N_38977);
nand U39033 (N_39033,N_38848,N_38777);
or U39034 (N_39034,N_38931,N_38804);
or U39035 (N_39035,N_38860,N_38763);
nor U39036 (N_39036,N_38806,N_38913);
nand U39037 (N_39037,N_38782,N_38902);
xnor U39038 (N_39038,N_38959,N_38781);
or U39039 (N_39039,N_38765,N_38858);
and U39040 (N_39040,N_38766,N_38893);
xnor U39041 (N_39041,N_38985,N_38903);
and U39042 (N_39042,N_38797,N_38757);
nor U39043 (N_39043,N_38831,N_38769);
xnor U39044 (N_39044,N_38864,N_38770);
nand U39045 (N_39045,N_38823,N_38945);
nand U39046 (N_39046,N_38886,N_38842);
nand U39047 (N_39047,N_38786,N_38962);
nor U39048 (N_39048,N_38875,N_38851);
nor U39049 (N_39049,N_38762,N_38927);
nor U39050 (N_39050,N_38930,N_38882);
nand U39051 (N_39051,N_38973,N_38873);
nand U39052 (N_39052,N_38859,N_38993);
or U39053 (N_39053,N_38783,N_38940);
nand U39054 (N_39054,N_38779,N_38952);
nand U39055 (N_39055,N_38794,N_38885);
or U39056 (N_39056,N_38790,N_38840);
nor U39057 (N_39057,N_38932,N_38999);
or U39058 (N_39058,N_38974,N_38961);
nor U39059 (N_39059,N_38921,N_38761);
nand U39060 (N_39060,N_38924,N_38796);
nor U39061 (N_39061,N_38778,N_38880);
nand U39062 (N_39062,N_38955,N_38789);
nand U39063 (N_39063,N_38901,N_38895);
nand U39064 (N_39064,N_38839,N_38995);
or U39065 (N_39065,N_38820,N_38764);
or U39066 (N_39066,N_38853,N_38812);
xnor U39067 (N_39067,N_38947,N_38829);
and U39068 (N_39068,N_38760,N_38826);
nand U39069 (N_39069,N_38946,N_38867);
and U39070 (N_39070,N_38915,N_38950);
xor U39071 (N_39071,N_38896,N_38756);
nor U39072 (N_39072,N_38972,N_38838);
nor U39073 (N_39073,N_38822,N_38785);
nor U39074 (N_39074,N_38984,N_38979);
nor U39075 (N_39075,N_38752,N_38926);
or U39076 (N_39076,N_38818,N_38956);
nand U39077 (N_39077,N_38814,N_38787);
or U39078 (N_39078,N_38907,N_38934);
nand U39079 (N_39079,N_38750,N_38802);
nor U39080 (N_39080,N_38793,N_38997);
nor U39081 (N_39081,N_38899,N_38809);
or U39082 (N_39082,N_38856,N_38996);
nor U39083 (N_39083,N_38780,N_38980);
or U39084 (N_39084,N_38894,N_38811);
and U39085 (N_39085,N_38881,N_38849);
nor U39086 (N_39086,N_38845,N_38998);
xor U39087 (N_39087,N_38992,N_38801);
nor U39088 (N_39088,N_38837,N_38841);
nor U39089 (N_39089,N_38986,N_38800);
nor U39090 (N_39090,N_38792,N_38888);
or U39091 (N_39091,N_38969,N_38773);
nand U39092 (N_39092,N_38910,N_38861);
nand U39093 (N_39093,N_38900,N_38825);
xor U39094 (N_39094,N_38892,N_38923);
or U39095 (N_39095,N_38846,N_38874);
or U39096 (N_39096,N_38994,N_38871);
or U39097 (N_39097,N_38803,N_38844);
nor U39098 (N_39098,N_38872,N_38751);
nand U39099 (N_39099,N_38918,N_38810);
nand U39100 (N_39100,N_38869,N_38919);
and U39101 (N_39101,N_38917,N_38816);
nor U39102 (N_39102,N_38788,N_38988);
or U39103 (N_39103,N_38911,N_38975);
nand U39104 (N_39104,N_38920,N_38978);
nor U39105 (N_39105,N_38866,N_38971);
nand U39106 (N_39106,N_38868,N_38914);
nor U39107 (N_39107,N_38981,N_38937);
or U39108 (N_39108,N_38857,N_38877);
nor U39109 (N_39109,N_38922,N_38948);
and U39110 (N_39110,N_38767,N_38943);
or U39111 (N_39111,N_38991,N_38832);
nand U39112 (N_39112,N_38966,N_38798);
nor U39113 (N_39113,N_38805,N_38963);
or U39114 (N_39114,N_38759,N_38830);
nand U39115 (N_39115,N_38890,N_38951);
nor U39116 (N_39116,N_38774,N_38938);
and U39117 (N_39117,N_38879,N_38965);
and U39118 (N_39118,N_38908,N_38819);
xor U39119 (N_39119,N_38958,N_38847);
nand U39120 (N_39120,N_38854,N_38768);
nor U39121 (N_39121,N_38824,N_38755);
nor U39122 (N_39122,N_38754,N_38821);
nand U39123 (N_39123,N_38855,N_38884);
nor U39124 (N_39124,N_38987,N_38828);
nand U39125 (N_39125,N_38896,N_38979);
or U39126 (N_39126,N_38808,N_38901);
nor U39127 (N_39127,N_38752,N_38958);
or U39128 (N_39128,N_38943,N_38911);
nand U39129 (N_39129,N_38956,N_38927);
nand U39130 (N_39130,N_38825,N_38939);
nand U39131 (N_39131,N_38908,N_38754);
or U39132 (N_39132,N_38893,N_38982);
xor U39133 (N_39133,N_38862,N_38841);
nand U39134 (N_39134,N_38933,N_38900);
nand U39135 (N_39135,N_38806,N_38957);
or U39136 (N_39136,N_38884,N_38836);
or U39137 (N_39137,N_38947,N_38820);
xnor U39138 (N_39138,N_38871,N_38902);
and U39139 (N_39139,N_38760,N_38856);
nor U39140 (N_39140,N_38975,N_38811);
or U39141 (N_39141,N_38780,N_38981);
nor U39142 (N_39142,N_38955,N_38860);
and U39143 (N_39143,N_38786,N_38876);
or U39144 (N_39144,N_38854,N_38933);
nor U39145 (N_39145,N_38933,N_38780);
nand U39146 (N_39146,N_38920,N_38830);
nand U39147 (N_39147,N_38791,N_38946);
and U39148 (N_39148,N_38902,N_38920);
xnor U39149 (N_39149,N_38758,N_38878);
nor U39150 (N_39150,N_38951,N_38979);
xor U39151 (N_39151,N_38752,N_38948);
nor U39152 (N_39152,N_38851,N_38808);
or U39153 (N_39153,N_38824,N_38976);
nand U39154 (N_39154,N_38767,N_38889);
nand U39155 (N_39155,N_38865,N_38821);
nor U39156 (N_39156,N_38966,N_38867);
nor U39157 (N_39157,N_38932,N_38822);
and U39158 (N_39158,N_38780,N_38783);
xor U39159 (N_39159,N_38921,N_38945);
and U39160 (N_39160,N_38960,N_38980);
nand U39161 (N_39161,N_38847,N_38773);
and U39162 (N_39162,N_38869,N_38865);
or U39163 (N_39163,N_38930,N_38878);
nor U39164 (N_39164,N_38982,N_38857);
xnor U39165 (N_39165,N_38781,N_38859);
xnor U39166 (N_39166,N_38799,N_38891);
nand U39167 (N_39167,N_38970,N_38830);
xor U39168 (N_39168,N_38840,N_38795);
nor U39169 (N_39169,N_38934,N_38870);
and U39170 (N_39170,N_38809,N_38881);
xnor U39171 (N_39171,N_38941,N_38855);
nand U39172 (N_39172,N_38755,N_38827);
nand U39173 (N_39173,N_38870,N_38871);
and U39174 (N_39174,N_38855,N_38804);
nand U39175 (N_39175,N_38787,N_38852);
or U39176 (N_39176,N_38796,N_38985);
nor U39177 (N_39177,N_38752,N_38930);
or U39178 (N_39178,N_38937,N_38853);
nor U39179 (N_39179,N_38941,N_38860);
or U39180 (N_39180,N_38990,N_38853);
nand U39181 (N_39181,N_38875,N_38817);
nand U39182 (N_39182,N_38872,N_38764);
nand U39183 (N_39183,N_38832,N_38932);
xor U39184 (N_39184,N_38785,N_38881);
xor U39185 (N_39185,N_38955,N_38889);
xnor U39186 (N_39186,N_38944,N_38881);
nand U39187 (N_39187,N_38877,N_38850);
xor U39188 (N_39188,N_38917,N_38833);
nand U39189 (N_39189,N_38779,N_38915);
or U39190 (N_39190,N_38794,N_38909);
xnor U39191 (N_39191,N_38970,N_38751);
nand U39192 (N_39192,N_38925,N_38984);
and U39193 (N_39193,N_38961,N_38771);
and U39194 (N_39194,N_38805,N_38841);
nor U39195 (N_39195,N_38885,N_38905);
or U39196 (N_39196,N_38854,N_38804);
xnor U39197 (N_39197,N_38919,N_38920);
or U39198 (N_39198,N_38920,N_38868);
xnor U39199 (N_39199,N_38778,N_38978);
xor U39200 (N_39200,N_38885,N_38974);
nor U39201 (N_39201,N_38955,N_38861);
nor U39202 (N_39202,N_38934,N_38871);
nor U39203 (N_39203,N_38887,N_38947);
or U39204 (N_39204,N_38915,N_38773);
or U39205 (N_39205,N_38869,N_38762);
or U39206 (N_39206,N_38854,N_38834);
and U39207 (N_39207,N_38967,N_38755);
and U39208 (N_39208,N_38782,N_38844);
xor U39209 (N_39209,N_38780,N_38840);
nor U39210 (N_39210,N_38997,N_38941);
xnor U39211 (N_39211,N_38915,N_38883);
xor U39212 (N_39212,N_38855,N_38969);
and U39213 (N_39213,N_38971,N_38978);
nand U39214 (N_39214,N_38866,N_38767);
nand U39215 (N_39215,N_38968,N_38880);
xor U39216 (N_39216,N_38985,N_38845);
and U39217 (N_39217,N_38762,N_38834);
nor U39218 (N_39218,N_38943,N_38881);
xor U39219 (N_39219,N_38919,N_38971);
nor U39220 (N_39220,N_38910,N_38858);
nand U39221 (N_39221,N_38803,N_38951);
and U39222 (N_39222,N_38840,N_38766);
nand U39223 (N_39223,N_38751,N_38797);
and U39224 (N_39224,N_38915,N_38952);
nor U39225 (N_39225,N_38867,N_38981);
xor U39226 (N_39226,N_38878,N_38816);
xnor U39227 (N_39227,N_38883,N_38852);
xor U39228 (N_39228,N_38930,N_38903);
nand U39229 (N_39229,N_38865,N_38751);
nand U39230 (N_39230,N_38826,N_38930);
nor U39231 (N_39231,N_38750,N_38868);
nand U39232 (N_39232,N_38785,N_38819);
and U39233 (N_39233,N_38801,N_38890);
xor U39234 (N_39234,N_38889,N_38865);
and U39235 (N_39235,N_38879,N_38894);
nand U39236 (N_39236,N_38895,N_38947);
and U39237 (N_39237,N_38785,N_38767);
nand U39238 (N_39238,N_38881,N_38885);
and U39239 (N_39239,N_38886,N_38773);
nand U39240 (N_39240,N_38932,N_38808);
or U39241 (N_39241,N_38848,N_38753);
nor U39242 (N_39242,N_38807,N_38856);
nor U39243 (N_39243,N_38777,N_38866);
or U39244 (N_39244,N_38882,N_38795);
xor U39245 (N_39245,N_38750,N_38837);
nand U39246 (N_39246,N_38882,N_38768);
or U39247 (N_39247,N_38879,N_38770);
xnor U39248 (N_39248,N_38910,N_38973);
and U39249 (N_39249,N_38923,N_38828);
nand U39250 (N_39250,N_39036,N_39097);
nand U39251 (N_39251,N_39080,N_39004);
nand U39252 (N_39252,N_39152,N_39211);
xor U39253 (N_39253,N_39062,N_39047);
and U39254 (N_39254,N_39221,N_39196);
and U39255 (N_39255,N_39111,N_39161);
nand U39256 (N_39256,N_39157,N_39213);
or U39257 (N_39257,N_39116,N_39020);
nor U39258 (N_39258,N_39076,N_39089);
xor U39259 (N_39259,N_39141,N_39171);
or U39260 (N_39260,N_39095,N_39085);
nand U39261 (N_39261,N_39023,N_39185);
xnor U39262 (N_39262,N_39203,N_39146);
nand U39263 (N_39263,N_39094,N_39025);
and U39264 (N_39264,N_39043,N_39104);
and U39265 (N_39265,N_39195,N_39125);
xor U39266 (N_39266,N_39138,N_39083);
or U39267 (N_39267,N_39038,N_39106);
nor U39268 (N_39268,N_39077,N_39242);
nand U39269 (N_39269,N_39016,N_39150);
or U39270 (N_39270,N_39073,N_39059);
nor U39271 (N_39271,N_39246,N_39173);
nor U39272 (N_39272,N_39117,N_39164);
nor U39273 (N_39273,N_39218,N_39057);
or U39274 (N_39274,N_39122,N_39001);
or U39275 (N_39275,N_39209,N_39159);
nor U39276 (N_39276,N_39224,N_39119);
or U39277 (N_39277,N_39028,N_39108);
or U39278 (N_39278,N_39132,N_39039);
and U39279 (N_39279,N_39230,N_39005);
nand U39280 (N_39280,N_39100,N_39056);
nand U39281 (N_39281,N_39178,N_39133);
xnor U39282 (N_39282,N_39172,N_39228);
or U39283 (N_39283,N_39029,N_39088);
and U39284 (N_39284,N_39035,N_39170);
and U39285 (N_39285,N_39024,N_39129);
nand U39286 (N_39286,N_39033,N_39053);
and U39287 (N_39287,N_39099,N_39091);
or U39288 (N_39288,N_39012,N_39189);
nand U39289 (N_39289,N_39009,N_39019);
nand U39290 (N_39290,N_39183,N_39032);
or U39291 (N_39291,N_39049,N_39214);
and U39292 (N_39292,N_39194,N_39151);
or U39293 (N_39293,N_39118,N_39014);
nand U39294 (N_39294,N_39115,N_39234);
nor U39295 (N_39295,N_39237,N_39148);
nor U39296 (N_39296,N_39075,N_39134);
and U39297 (N_39297,N_39041,N_39092);
or U39298 (N_39298,N_39210,N_39040);
xor U39299 (N_39299,N_39105,N_39034);
nor U39300 (N_39300,N_39205,N_39238);
xnor U39301 (N_39301,N_39090,N_39065);
and U39302 (N_39302,N_39160,N_39082);
or U39303 (N_39303,N_39165,N_39081);
nand U39304 (N_39304,N_39193,N_39169);
xor U39305 (N_39305,N_39204,N_39154);
nor U39306 (N_39306,N_39113,N_39231);
or U39307 (N_39307,N_39120,N_39236);
xor U39308 (N_39308,N_39124,N_39008);
nand U39309 (N_39309,N_39128,N_39098);
or U39310 (N_39310,N_39068,N_39147);
nand U39311 (N_39311,N_39158,N_39137);
nor U39312 (N_39312,N_39051,N_39144);
and U39313 (N_39313,N_39191,N_39072);
xnor U39314 (N_39314,N_39084,N_39067);
and U39315 (N_39315,N_39217,N_39123);
or U39316 (N_39316,N_39149,N_39070);
nand U39317 (N_39317,N_39121,N_39168);
xor U39318 (N_39318,N_39010,N_39215);
xnor U39319 (N_39319,N_39079,N_39223);
xor U39320 (N_39320,N_39011,N_39006);
nor U39321 (N_39321,N_39015,N_39227);
nor U39322 (N_39322,N_39000,N_39240);
xor U39323 (N_39323,N_39248,N_39187);
nand U39324 (N_39324,N_39199,N_39101);
xnor U39325 (N_39325,N_39037,N_39096);
nor U39326 (N_39326,N_39044,N_39109);
nor U39327 (N_39327,N_39190,N_39167);
and U39328 (N_39328,N_39114,N_39163);
nor U39329 (N_39329,N_39078,N_39206);
or U39330 (N_39330,N_39130,N_39245);
or U39331 (N_39331,N_39233,N_39143);
and U39332 (N_39332,N_39186,N_39179);
and U39333 (N_39333,N_39232,N_39042);
and U39334 (N_39334,N_39060,N_39162);
nand U39335 (N_39335,N_39244,N_39155);
xnor U39336 (N_39336,N_39027,N_39064);
or U39337 (N_39337,N_39007,N_39021);
and U39338 (N_39338,N_39048,N_39071);
nor U39339 (N_39339,N_39140,N_39127);
nor U39340 (N_39340,N_39142,N_39181);
or U39341 (N_39341,N_39184,N_39241);
nor U39342 (N_39342,N_39022,N_39017);
or U39343 (N_39343,N_39107,N_39093);
and U39344 (N_39344,N_39074,N_39202);
xor U39345 (N_39345,N_39239,N_39102);
nand U39346 (N_39346,N_39026,N_39201);
xor U39347 (N_39347,N_39243,N_39139);
xor U39348 (N_39348,N_39112,N_39063);
xor U39349 (N_39349,N_39131,N_39153);
and U39350 (N_39350,N_39003,N_39054);
xnor U39351 (N_39351,N_39249,N_39197);
nor U39352 (N_39352,N_39175,N_39086);
xnor U39353 (N_39353,N_39013,N_39050);
nand U39354 (N_39354,N_39055,N_39216);
xor U39355 (N_39355,N_39200,N_39136);
and U39356 (N_39356,N_39002,N_39247);
nor U39357 (N_39357,N_39058,N_39069);
xor U39358 (N_39358,N_39198,N_39235);
and U39359 (N_39359,N_39045,N_39110);
nand U39360 (N_39360,N_39225,N_39212);
or U39361 (N_39361,N_39176,N_39220);
nand U39362 (N_39362,N_39222,N_39103);
and U39363 (N_39363,N_39219,N_39166);
xor U39364 (N_39364,N_39177,N_39207);
and U39365 (N_39365,N_39174,N_39018);
and U39366 (N_39366,N_39226,N_39030);
and U39367 (N_39367,N_39208,N_39046);
nand U39368 (N_39368,N_39061,N_39087);
xnor U39369 (N_39369,N_39229,N_39188);
nand U39370 (N_39370,N_39182,N_39031);
nand U39371 (N_39371,N_39192,N_39126);
and U39372 (N_39372,N_39180,N_39066);
nand U39373 (N_39373,N_39135,N_39145);
xor U39374 (N_39374,N_39156,N_39052);
and U39375 (N_39375,N_39192,N_39230);
nor U39376 (N_39376,N_39037,N_39212);
nor U39377 (N_39377,N_39215,N_39138);
xor U39378 (N_39378,N_39185,N_39133);
xor U39379 (N_39379,N_39056,N_39124);
nor U39380 (N_39380,N_39169,N_39119);
and U39381 (N_39381,N_39062,N_39209);
or U39382 (N_39382,N_39175,N_39242);
or U39383 (N_39383,N_39010,N_39180);
nand U39384 (N_39384,N_39245,N_39239);
xor U39385 (N_39385,N_39229,N_39026);
xor U39386 (N_39386,N_39118,N_39163);
or U39387 (N_39387,N_39115,N_39177);
or U39388 (N_39388,N_39045,N_39128);
xor U39389 (N_39389,N_39125,N_39035);
xor U39390 (N_39390,N_39062,N_39085);
nor U39391 (N_39391,N_39006,N_39059);
or U39392 (N_39392,N_39247,N_39169);
and U39393 (N_39393,N_39026,N_39008);
xor U39394 (N_39394,N_39068,N_39204);
and U39395 (N_39395,N_39205,N_39004);
xnor U39396 (N_39396,N_39101,N_39085);
nand U39397 (N_39397,N_39206,N_39153);
xnor U39398 (N_39398,N_39038,N_39143);
nor U39399 (N_39399,N_39024,N_39044);
and U39400 (N_39400,N_39025,N_39088);
nand U39401 (N_39401,N_39134,N_39010);
and U39402 (N_39402,N_39174,N_39044);
nand U39403 (N_39403,N_39068,N_39055);
nand U39404 (N_39404,N_39112,N_39080);
xnor U39405 (N_39405,N_39156,N_39090);
xnor U39406 (N_39406,N_39161,N_39100);
or U39407 (N_39407,N_39146,N_39097);
or U39408 (N_39408,N_39061,N_39083);
nand U39409 (N_39409,N_39132,N_39003);
xnor U39410 (N_39410,N_39119,N_39154);
nand U39411 (N_39411,N_39196,N_39074);
or U39412 (N_39412,N_39223,N_39141);
and U39413 (N_39413,N_39012,N_39106);
nor U39414 (N_39414,N_39107,N_39133);
xnor U39415 (N_39415,N_39165,N_39092);
and U39416 (N_39416,N_39139,N_39133);
and U39417 (N_39417,N_39046,N_39158);
nor U39418 (N_39418,N_39111,N_39030);
nor U39419 (N_39419,N_39230,N_39167);
or U39420 (N_39420,N_39124,N_39130);
and U39421 (N_39421,N_39005,N_39147);
nand U39422 (N_39422,N_39064,N_39247);
xor U39423 (N_39423,N_39062,N_39123);
and U39424 (N_39424,N_39005,N_39187);
and U39425 (N_39425,N_39077,N_39199);
or U39426 (N_39426,N_39005,N_39176);
and U39427 (N_39427,N_39046,N_39224);
nor U39428 (N_39428,N_39135,N_39065);
and U39429 (N_39429,N_39060,N_39105);
or U39430 (N_39430,N_39136,N_39002);
or U39431 (N_39431,N_39238,N_39103);
nand U39432 (N_39432,N_39087,N_39235);
xnor U39433 (N_39433,N_39207,N_39003);
nand U39434 (N_39434,N_39019,N_39046);
and U39435 (N_39435,N_39140,N_39085);
nor U39436 (N_39436,N_39110,N_39057);
nand U39437 (N_39437,N_39194,N_39035);
and U39438 (N_39438,N_39082,N_39178);
and U39439 (N_39439,N_39218,N_39140);
or U39440 (N_39440,N_39236,N_39032);
xnor U39441 (N_39441,N_39010,N_39020);
or U39442 (N_39442,N_39179,N_39079);
nand U39443 (N_39443,N_39183,N_39170);
nand U39444 (N_39444,N_39244,N_39111);
and U39445 (N_39445,N_39179,N_39026);
or U39446 (N_39446,N_39116,N_39119);
nor U39447 (N_39447,N_39057,N_39224);
xnor U39448 (N_39448,N_39222,N_39042);
nor U39449 (N_39449,N_39058,N_39018);
xor U39450 (N_39450,N_39155,N_39086);
xor U39451 (N_39451,N_39146,N_39211);
and U39452 (N_39452,N_39098,N_39019);
xnor U39453 (N_39453,N_39012,N_39158);
and U39454 (N_39454,N_39220,N_39050);
xnor U39455 (N_39455,N_39134,N_39199);
nor U39456 (N_39456,N_39051,N_39244);
or U39457 (N_39457,N_39130,N_39244);
or U39458 (N_39458,N_39205,N_39206);
nand U39459 (N_39459,N_39193,N_39214);
or U39460 (N_39460,N_39182,N_39040);
or U39461 (N_39461,N_39216,N_39116);
or U39462 (N_39462,N_39040,N_39095);
and U39463 (N_39463,N_39057,N_39210);
nand U39464 (N_39464,N_39248,N_39119);
nor U39465 (N_39465,N_39139,N_39053);
and U39466 (N_39466,N_39237,N_39089);
nor U39467 (N_39467,N_39004,N_39158);
and U39468 (N_39468,N_39041,N_39039);
nor U39469 (N_39469,N_39026,N_39120);
nand U39470 (N_39470,N_39076,N_39193);
nor U39471 (N_39471,N_39045,N_39048);
nor U39472 (N_39472,N_39143,N_39162);
nor U39473 (N_39473,N_39005,N_39175);
and U39474 (N_39474,N_39150,N_39000);
or U39475 (N_39475,N_39089,N_39228);
nor U39476 (N_39476,N_39019,N_39013);
and U39477 (N_39477,N_39072,N_39210);
nor U39478 (N_39478,N_39011,N_39030);
nor U39479 (N_39479,N_39047,N_39024);
and U39480 (N_39480,N_39144,N_39142);
nor U39481 (N_39481,N_39045,N_39093);
and U39482 (N_39482,N_39023,N_39014);
nor U39483 (N_39483,N_39210,N_39024);
and U39484 (N_39484,N_39120,N_39208);
or U39485 (N_39485,N_39015,N_39007);
or U39486 (N_39486,N_39049,N_39073);
xor U39487 (N_39487,N_39068,N_39189);
or U39488 (N_39488,N_39098,N_39126);
nor U39489 (N_39489,N_39203,N_39090);
nand U39490 (N_39490,N_39062,N_39071);
or U39491 (N_39491,N_39245,N_39148);
xor U39492 (N_39492,N_39245,N_39177);
and U39493 (N_39493,N_39022,N_39122);
and U39494 (N_39494,N_39161,N_39050);
xnor U39495 (N_39495,N_39072,N_39220);
and U39496 (N_39496,N_39096,N_39114);
nor U39497 (N_39497,N_39122,N_39119);
and U39498 (N_39498,N_39074,N_39084);
nor U39499 (N_39499,N_39138,N_39197);
and U39500 (N_39500,N_39421,N_39330);
xnor U39501 (N_39501,N_39306,N_39459);
nor U39502 (N_39502,N_39352,N_39473);
nand U39503 (N_39503,N_39284,N_39420);
nor U39504 (N_39504,N_39364,N_39267);
xnor U39505 (N_39505,N_39400,N_39261);
xnor U39506 (N_39506,N_39262,N_39436);
nand U39507 (N_39507,N_39403,N_39431);
xor U39508 (N_39508,N_39369,N_39456);
or U39509 (N_39509,N_39366,N_39353);
nor U39510 (N_39510,N_39370,N_39299);
nor U39511 (N_39511,N_39355,N_39308);
or U39512 (N_39512,N_39418,N_39401);
or U39513 (N_39513,N_39336,N_39331);
or U39514 (N_39514,N_39452,N_39263);
or U39515 (N_39515,N_39309,N_39435);
nand U39516 (N_39516,N_39256,N_39254);
or U39517 (N_39517,N_39340,N_39354);
xor U39518 (N_39518,N_39408,N_39350);
xnor U39519 (N_39519,N_39455,N_39493);
nor U39520 (N_39520,N_39314,N_39379);
xnor U39521 (N_39521,N_39425,N_39441);
nor U39522 (N_39522,N_39499,N_39342);
xnor U39523 (N_39523,N_39270,N_39358);
xnor U39524 (N_39524,N_39332,N_39334);
or U39525 (N_39525,N_39383,N_39414);
xnor U39526 (N_39526,N_39470,N_39395);
xnor U39527 (N_39527,N_39349,N_39496);
nor U39528 (N_39528,N_39384,N_39329);
nor U39529 (N_39529,N_39326,N_39438);
and U39530 (N_39530,N_39323,N_39391);
nor U39531 (N_39531,N_39333,N_39375);
nand U39532 (N_39532,N_39345,N_39365);
nor U39533 (N_39533,N_39362,N_39347);
xor U39534 (N_39534,N_39392,N_39396);
nor U39535 (N_39535,N_39250,N_39387);
nor U39536 (N_39536,N_39399,N_39462);
and U39537 (N_39537,N_39491,N_39446);
or U39538 (N_39538,N_39293,N_39419);
and U39539 (N_39539,N_39337,N_39386);
and U39540 (N_39540,N_39477,N_39482);
nand U39541 (N_39541,N_39259,N_39339);
nand U39542 (N_39542,N_39453,N_39351);
xnor U39543 (N_39543,N_39382,N_39405);
nor U39544 (N_39544,N_39252,N_39303);
xnor U39545 (N_39545,N_39480,N_39372);
xor U39546 (N_39546,N_39301,N_39494);
nand U39547 (N_39547,N_39285,N_39363);
xnor U39548 (N_39548,N_39427,N_39497);
nor U39549 (N_39549,N_39495,N_39286);
nand U39550 (N_39550,N_39412,N_39317);
nand U39551 (N_39551,N_39447,N_39279);
nand U39552 (N_39552,N_39321,N_39422);
nand U39553 (N_39553,N_39458,N_39492);
nor U39554 (N_39554,N_39442,N_39268);
nor U39555 (N_39555,N_39433,N_39484);
nand U39556 (N_39556,N_39343,N_39440);
nand U39557 (N_39557,N_39388,N_39402);
nand U39558 (N_39558,N_39476,N_39302);
xnor U39559 (N_39559,N_39416,N_39269);
xor U39560 (N_39560,N_39457,N_39428);
nand U39561 (N_39561,N_39292,N_39485);
and U39562 (N_39562,N_39407,N_39315);
or U39563 (N_39563,N_39487,N_39469);
nor U39564 (N_39564,N_39411,N_39390);
nor U39565 (N_39565,N_39255,N_39460);
xnor U39566 (N_39566,N_39335,N_39277);
nand U39567 (N_39567,N_39313,N_39472);
nor U39568 (N_39568,N_39280,N_39371);
xor U39569 (N_39569,N_39409,N_39320);
nor U39570 (N_39570,N_39311,N_39291);
nand U39571 (N_39571,N_39264,N_39278);
xnor U39572 (N_39572,N_39271,N_39415);
xor U39573 (N_39573,N_39486,N_39294);
xor U39574 (N_39574,N_39310,N_39474);
and U39575 (N_39575,N_39430,N_39410);
nor U39576 (N_39576,N_39361,N_39376);
or U39577 (N_39577,N_39283,N_39467);
or U39578 (N_39578,N_39489,N_39468);
and U39579 (N_39579,N_39348,N_39318);
xnor U39580 (N_39580,N_39341,N_39454);
and U39581 (N_39581,N_39377,N_39439);
nor U39582 (N_39582,N_39295,N_39258);
nand U39583 (N_39583,N_39378,N_39338);
or U39584 (N_39584,N_39464,N_39297);
nand U39585 (N_39585,N_39393,N_39305);
nor U39586 (N_39586,N_39466,N_39406);
nor U39587 (N_39587,N_39296,N_39450);
or U39588 (N_39588,N_39479,N_39451);
nor U39589 (N_39589,N_39275,N_39394);
xor U39590 (N_39590,N_39488,N_39423);
nor U39591 (N_39591,N_39304,N_39312);
xor U39592 (N_39592,N_39287,N_39265);
or U39593 (N_39593,N_39322,N_39298);
xor U39594 (N_39594,N_39381,N_39385);
xor U39595 (N_39595,N_39290,N_39253);
nor U39596 (N_39596,N_39344,N_39357);
nand U39597 (N_39597,N_39274,N_39319);
and U39598 (N_39598,N_39404,N_39398);
or U39599 (N_39599,N_39374,N_39368);
xnor U39600 (N_39600,N_39373,N_39465);
xnor U39601 (N_39601,N_39498,N_39424);
xor U39602 (N_39602,N_39443,N_39445);
and U39603 (N_39603,N_39356,N_39281);
xor U39604 (N_39604,N_39300,N_39448);
and U39605 (N_39605,N_39449,N_39346);
nor U39606 (N_39606,N_39316,N_39413);
nor U39607 (N_39607,N_39273,N_39324);
nor U39608 (N_39608,N_39434,N_39266);
nand U39609 (N_39609,N_39282,N_39389);
nor U39610 (N_39610,N_39481,N_39307);
and U39611 (N_39611,N_39478,N_39463);
or U39612 (N_39612,N_39461,N_39328);
xor U39613 (N_39613,N_39367,N_39417);
and U39614 (N_39614,N_39251,N_39380);
nor U39615 (N_39615,N_39490,N_39429);
nor U39616 (N_39616,N_39471,N_39257);
and U39617 (N_39617,N_39288,N_39426);
nand U39618 (N_39618,N_39444,N_39325);
nor U39619 (N_39619,N_39437,N_39327);
nand U39620 (N_39620,N_39397,N_39272);
nor U39621 (N_39621,N_39260,N_39432);
nor U39622 (N_39622,N_39475,N_39359);
nand U39623 (N_39623,N_39289,N_39483);
xor U39624 (N_39624,N_39276,N_39360);
nor U39625 (N_39625,N_39448,N_39477);
nor U39626 (N_39626,N_39361,N_39404);
or U39627 (N_39627,N_39456,N_39446);
xor U39628 (N_39628,N_39377,N_39469);
nand U39629 (N_39629,N_39311,N_39339);
nor U39630 (N_39630,N_39429,N_39341);
nand U39631 (N_39631,N_39270,N_39257);
xnor U39632 (N_39632,N_39271,N_39366);
and U39633 (N_39633,N_39470,N_39355);
nand U39634 (N_39634,N_39351,N_39408);
nor U39635 (N_39635,N_39296,N_39491);
nor U39636 (N_39636,N_39421,N_39351);
or U39637 (N_39637,N_39476,N_39410);
nand U39638 (N_39638,N_39253,N_39373);
or U39639 (N_39639,N_39267,N_39494);
xor U39640 (N_39640,N_39338,N_39479);
nor U39641 (N_39641,N_39284,N_39351);
or U39642 (N_39642,N_39318,N_39269);
and U39643 (N_39643,N_39293,N_39333);
or U39644 (N_39644,N_39473,N_39397);
xnor U39645 (N_39645,N_39357,N_39410);
and U39646 (N_39646,N_39392,N_39489);
nor U39647 (N_39647,N_39441,N_39439);
xnor U39648 (N_39648,N_39313,N_39444);
nor U39649 (N_39649,N_39307,N_39495);
nor U39650 (N_39650,N_39404,N_39367);
xor U39651 (N_39651,N_39376,N_39252);
and U39652 (N_39652,N_39425,N_39261);
and U39653 (N_39653,N_39289,N_39317);
nor U39654 (N_39654,N_39469,N_39351);
nor U39655 (N_39655,N_39324,N_39436);
nand U39656 (N_39656,N_39319,N_39384);
or U39657 (N_39657,N_39372,N_39413);
or U39658 (N_39658,N_39269,N_39405);
xnor U39659 (N_39659,N_39303,N_39308);
or U39660 (N_39660,N_39330,N_39285);
xor U39661 (N_39661,N_39463,N_39450);
nor U39662 (N_39662,N_39280,N_39282);
nor U39663 (N_39663,N_39380,N_39334);
and U39664 (N_39664,N_39336,N_39283);
xnor U39665 (N_39665,N_39255,N_39441);
or U39666 (N_39666,N_39412,N_39355);
nor U39667 (N_39667,N_39398,N_39363);
nor U39668 (N_39668,N_39379,N_39424);
and U39669 (N_39669,N_39491,N_39428);
and U39670 (N_39670,N_39368,N_39272);
nor U39671 (N_39671,N_39414,N_39313);
and U39672 (N_39672,N_39423,N_39366);
nand U39673 (N_39673,N_39259,N_39328);
and U39674 (N_39674,N_39438,N_39452);
xnor U39675 (N_39675,N_39283,N_39418);
xnor U39676 (N_39676,N_39496,N_39318);
xnor U39677 (N_39677,N_39358,N_39454);
or U39678 (N_39678,N_39307,N_39489);
xor U39679 (N_39679,N_39384,N_39426);
nor U39680 (N_39680,N_39381,N_39474);
nand U39681 (N_39681,N_39256,N_39498);
nand U39682 (N_39682,N_39335,N_39367);
and U39683 (N_39683,N_39462,N_39310);
nor U39684 (N_39684,N_39435,N_39417);
and U39685 (N_39685,N_39484,N_39415);
or U39686 (N_39686,N_39259,N_39457);
nor U39687 (N_39687,N_39486,N_39439);
nor U39688 (N_39688,N_39380,N_39324);
and U39689 (N_39689,N_39332,N_39260);
or U39690 (N_39690,N_39433,N_39350);
xnor U39691 (N_39691,N_39343,N_39425);
or U39692 (N_39692,N_39343,N_39477);
xor U39693 (N_39693,N_39379,N_39366);
xnor U39694 (N_39694,N_39330,N_39448);
and U39695 (N_39695,N_39394,N_39316);
and U39696 (N_39696,N_39278,N_39461);
and U39697 (N_39697,N_39349,N_39292);
nor U39698 (N_39698,N_39388,N_39410);
or U39699 (N_39699,N_39374,N_39409);
nor U39700 (N_39700,N_39463,N_39465);
nand U39701 (N_39701,N_39329,N_39451);
xor U39702 (N_39702,N_39294,N_39295);
and U39703 (N_39703,N_39329,N_39455);
or U39704 (N_39704,N_39361,N_39464);
and U39705 (N_39705,N_39439,N_39472);
nand U39706 (N_39706,N_39406,N_39334);
xnor U39707 (N_39707,N_39408,N_39487);
nor U39708 (N_39708,N_39482,N_39286);
and U39709 (N_39709,N_39288,N_39460);
nor U39710 (N_39710,N_39456,N_39471);
and U39711 (N_39711,N_39498,N_39448);
and U39712 (N_39712,N_39335,N_39315);
xor U39713 (N_39713,N_39374,N_39459);
and U39714 (N_39714,N_39398,N_39492);
and U39715 (N_39715,N_39310,N_39371);
xor U39716 (N_39716,N_39412,N_39453);
xor U39717 (N_39717,N_39253,N_39388);
nand U39718 (N_39718,N_39489,N_39371);
nand U39719 (N_39719,N_39478,N_39253);
nand U39720 (N_39720,N_39275,N_39316);
nor U39721 (N_39721,N_39317,N_39343);
xnor U39722 (N_39722,N_39404,N_39351);
xnor U39723 (N_39723,N_39347,N_39386);
xor U39724 (N_39724,N_39415,N_39253);
xnor U39725 (N_39725,N_39327,N_39307);
nor U39726 (N_39726,N_39339,N_39498);
or U39727 (N_39727,N_39282,N_39457);
and U39728 (N_39728,N_39488,N_39334);
or U39729 (N_39729,N_39447,N_39318);
xor U39730 (N_39730,N_39316,N_39308);
nand U39731 (N_39731,N_39268,N_39312);
nor U39732 (N_39732,N_39290,N_39263);
xnor U39733 (N_39733,N_39396,N_39399);
xnor U39734 (N_39734,N_39459,N_39318);
nor U39735 (N_39735,N_39438,N_39316);
nand U39736 (N_39736,N_39348,N_39469);
xor U39737 (N_39737,N_39435,N_39495);
nand U39738 (N_39738,N_39481,N_39290);
nand U39739 (N_39739,N_39339,N_39334);
nand U39740 (N_39740,N_39356,N_39263);
or U39741 (N_39741,N_39488,N_39353);
xor U39742 (N_39742,N_39362,N_39258);
xor U39743 (N_39743,N_39447,N_39377);
or U39744 (N_39744,N_39361,N_39289);
xnor U39745 (N_39745,N_39466,N_39376);
nor U39746 (N_39746,N_39293,N_39301);
or U39747 (N_39747,N_39260,N_39308);
or U39748 (N_39748,N_39425,N_39333);
xor U39749 (N_39749,N_39468,N_39339);
nor U39750 (N_39750,N_39693,N_39527);
xnor U39751 (N_39751,N_39697,N_39701);
xor U39752 (N_39752,N_39638,N_39535);
nand U39753 (N_39753,N_39529,N_39664);
xnor U39754 (N_39754,N_39680,N_39665);
nand U39755 (N_39755,N_39602,N_39647);
nor U39756 (N_39756,N_39604,N_39713);
or U39757 (N_39757,N_39532,N_39674);
or U39758 (N_39758,N_39575,N_39518);
or U39759 (N_39759,N_39623,N_39534);
nand U39760 (N_39760,N_39550,N_39513);
nand U39761 (N_39761,N_39576,N_39606);
nor U39762 (N_39762,N_39577,N_39642);
and U39763 (N_39763,N_39671,N_39511);
and U39764 (N_39764,N_39591,N_39553);
nand U39765 (N_39765,N_39627,N_39525);
nand U39766 (N_39766,N_39578,N_39698);
nand U39767 (N_39767,N_39676,N_39547);
and U39768 (N_39768,N_39569,N_39579);
nand U39769 (N_39769,N_39669,N_39572);
nor U39770 (N_39770,N_39708,N_39560);
nand U39771 (N_39771,N_39558,N_39537);
nor U39772 (N_39772,N_39666,N_39538);
xnor U39773 (N_39773,N_39622,N_39555);
and U39774 (N_39774,N_39519,N_39749);
and U39775 (N_39775,N_39733,N_39641);
nand U39776 (N_39776,N_39643,N_39636);
or U39777 (N_39777,N_39726,N_39611);
nor U39778 (N_39778,N_39719,N_39565);
and U39779 (N_39779,N_39546,N_39710);
nor U39780 (N_39780,N_39603,N_39645);
nand U39781 (N_39781,N_39735,N_39600);
nor U39782 (N_39782,N_39514,N_39656);
nand U39783 (N_39783,N_39615,N_39651);
and U39784 (N_39784,N_39703,N_39571);
nand U39785 (N_39785,N_39542,N_39630);
and U39786 (N_39786,N_39731,N_39712);
nand U39787 (N_39787,N_39617,N_39631);
xor U39788 (N_39788,N_39556,N_39704);
and U39789 (N_39789,N_39748,N_39644);
and U39790 (N_39790,N_39567,N_39573);
and U39791 (N_39791,N_39747,N_39706);
or U39792 (N_39792,N_39725,N_39738);
nor U39793 (N_39793,N_39740,N_39681);
nand U39794 (N_39794,N_39728,N_39718);
nand U39795 (N_39795,N_39677,N_39654);
or U39796 (N_39796,N_39689,N_39683);
and U39797 (N_39797,N_39709,N_39563);
nor U39798 (N_39798,N_39614,N_39715);
and U39799 (N_39799,N_39522,N_39690);
or U39800 (N_39800,N_39520,N_39545);
and U39801 (N_39801,N_39661,N_39646);
nor U39802 (N_39802,N_39505,N_39652);
nor U39803 (N_39803,N_39516,N_39593);
and U39804 (N_39804,N_39620,N_39566);
nor U39805 (N_39805,N_39580,N_39624);
or U39806 (N_39806,N_39616,N_39730);
or U39807 (N_39807,N_39588,N_39509);
and U39808 (N_39808,N_39552,N_39720);
and U39809 (N_39809,N_39657,N_39632);
or U39810 (N_39810,N_39524,N_39668);
xnor U39811 (N_39811,N_39702,N_39549);
nand U39812 (N_39812,N_39705,N_39587);
nor U39813 (N_39813,N_39590,N_39727);
nand U39814 (N_39814,N_39692,N_39714);
and U39815 (N_39815,N_39598,N_39621);
xnor U39816 (N_39816,N_39619,N_39679);
and U39817 (N_39817,N_39515,N_39732);
nor U39818 (N_39818,N_39739,N_39530);
xnor U39819 (N_39819,N_39521,N_39557);
nand U39820 (N_39820,N_39673,N_39559);
nand U39821 (N_39821,N_39684,N_39607);
and U39822 (N_39822,N_39648,N_39536);
and U39823 (N_39823,N_39551,N_39517);
nand U39824 (N_39824,N_39586,N_39584);
nand U39825 (N_39825,N_39601,N_39554);
and U39826 (N_39826,N_39734,N_39629);
and U39827 (N_39827,N_39533,N_39548);
or U39828 (N_39828,N_39543,N_39723);
and U39829 (N_39829,N_39599,N_39507);
nor U39830 (N_39830,N_39508,N_39682);
and U39831 (N_39831,N_39628,N_39539);
or U39832 (N_39832,N_39717,N_39564);
nor U39833 (N_39833,N_39592,N_39695);
and U39834 (N_39834,N_39523,N_39596);
nor U39835 (N_39835,N_39688,N_39626);
and U39836 (N_39836,N_39687,N_39736);
or U39837 (N_39837,N_39594,N_39568);
nand U39838 (N_39838,N_39583,N_39658);
and U39839 (N_39839,N_39605,N_39589);
and U39840 (N_39840,N_39561,N_39581);
xnor U39841 (N_39841,N_39653,N_39640);
nor U39842 (N_39842,N_39613,N_39526);
xor U39843 (N_39843,N_39650,N_39597);
nor U39844 (N_39844,N_39649,N_39585);
nand U39845 (N_39845,N_39667,N_39562);
and U39846 (N_39846,N_39729,N_39741);
or U39847 (N_39847,N_39694,N_39541);
nor U39848 (N_39848,N_39659,N_39686);
and U39849 (N_39849,N_39672,N_39696);
nand U39850 (N_39850,N_39582,N_39500);
xor U39851 (N_39851,N_39711,N_39707);
or U39852 (N_39852,N_39612,N_39528);
xnor U39853 (N_39853,N_39506,N_39743);
or U39854 (N_39854,N_39721,N_39663);
nor U39855 (N_39855,N_39510,N_39512);
nand U39856 (N_39856,N_39540,N_39746);
and U39857 (N_39857,N_39501,N_39724);
xnor U39858 (N_39858,N_39716,N_39531);
nor U39859 (N_39859,N_39634,N_39744);
xor U39860 (N_39860,N_39675,N_39662);
xor U39861 (N_39861,N_39670,N_39633);
and U39862 (N_39862,N_39503,N_39618);
and U39863 (N_39863,N_39742,N_39639);
and U39864 (N_39864,N_39737,N_39637);
or U39865 (N_39865,N_39595,N_39660);
xor U39866 (N_39866,N_39655,N_39700);
and U39867 (N_39867,N_39699,N_39570);
xor U39868 (N_39868,N_39678,N_39574);
or U39869 (N_39869,N_39609,N_39544);
or U39870 (N_39870,N_39502,N_39745);
xor U39871 (N_39871,N_39685,N_39608);
or U39872 (N_39872,N_39691,N_39625);
and U39873 (N_39873,N_39722,N_39504);
nand U39874 (N_39874,N_39610,N_39635);
xor U39875 (N_39875,N_39621,N_39538);
nor U39876 (N_39876,N_39628,N_39712);
xnor U39877 (N_39877,N_39609,N_39716);
nand U39878 (N_39878,N_39671,N_39556);
xnor U39879 (N_39879,N_39632,N_39578);
and U39880 (N_39880,N_39530,N_39595);
or U39881 (N_39881,N_39635,N_39743);
nand U39882 (N_39882,N_39747,N_39649);
nand U39883 (N_39883,N_39521,N_39631);
xor U39884 (N_39884,N_39547,N_39563);
or U39885 (N_39885,N_39642,N_39569);
nor U39886 (N_39886,N_39728,N_39663);
xnor U39887 (N_39887,N_39699,N_39569);
xnor U39888 (N_39888,N_39550,N_39644);
and U39889 (N_39889,N_39675,N_39720);
nand U39890 (N_39890,N_39711,N_39620);
xor U39891 (N_39891,N_39625,N_39624);
or U39892 (N_39892,N_39731,N_39525);
nand U39893 (N_39893,N_39543,N_39545);
and U39894 (N_39894,N_39694,N_39695);
nor U39895 (N_39895,N_39721,N_39704);
or U39896 (N_39896,N_39598,N_39741);
nand U39897 (N_39897,N_39668,N_39576);
or U39898 (N_39898,N_39571,N_39726);
and U39899 (N_39899,N_39740,N_39636);
and U39900 (N_39900,N_39729,N_39531);
and U39901 (N_39901,N_39742,N_39743);
xor U39902 (N_39902,N_39726,N_39643);
nor U39903 (N_39903,N_39661,N_39582);
and U39904 (N_39904,N_39602,N_39626);
and U39905 (N_39905,N_39679,N_39713);
and U39906 (N_39906,N_39592,N_39521);
nor U39907 (N_39907,N_39535,N_39703);
nor U39908 (N_39908,N_39586,N_39521);
and U39909 (N_39909,N_39637,N_39623);
xnor U39910 (N_39910,N_39515,N_39528);
xnor U39911 (N_39911,N_39582,N_39613);
and U39912 (N_39912,N_39610,N_39724);
nor U39913 (N_39913,N_39659,N_39661);
or U39914 (N_39914,N_39571,N_39716);
nand U39915 (N_39915,N_39514,N_39601);
nand U39916 (N_39916,N_39572,N_39542);
nand U39917 (N_39917,N_39745,N_39732);
or U39918 (N_39918,N_39528,N_39585);
nand U39919 (N_39919,N_39589,N_39661);
xor U39920 (N_39920,N_39609,N_39524);
nor U39921 (N_39921,N_39687,N_39583);
and U39922 (N_39922,N_39744,N_39632);
xnor U39923 (N_39923,N_39609,N_39523);
nor U39924 (N_39924,N_39550,N_39606);
or U39925 (N_39925,N_39529,N_39582);
xor U39926 (N_39926,N_39550,N_39682);
nor U39927 (N_39927,N_39627,N_39581);
and U39928 (N_39928,N_39644,N_39721);
nand U39929 (N_39929,N_39591,N_39648);
xnor U39930 (N_39930,N_39701,N_39512);
xnor U39931 (N_39931,N_39647,N_39600);
or U39932 (N_39932,N_39642,N_39662);
and U39933 (N_39933,N_39696,N_39563);
or U39934 (N_39934,N_39638,N_39672);
xor U39935 (N_39935,N_39524,N_39642);
xnor U39936 (N_39936,N_39615,N_39575);
nor U39937 (N_39937,N_39556,N_39523);
nand U39938 (N_39938,N_39748,N_39713);
and U39939 (N_39939,N_39572,N_39742);
and U39940 (N_39940,N_39689,N_39631);
or U39941 (N_39941,N_39598,N_39638);
nor U39942 (N_39942,N_39708,N_39565);
nand U39943 (N_39943,N_39690,N_39537);
nor U39944 (N_39944,N_39645,N_39538);
or U39945 (N_39945,N_39680,N_39717);
and U39946 (N_39946,N_39604,N_39631);
nand U39947 (N_39947,N_39613,N_39663);
xnor U39948 (N_39948,N_39502,N_39637);
nor U39949 (N_39949,N_39568,N_39576);
nor U39950 (N_39950,N_39721,N_39561);
and U39951 (N_39951,N_39529,N_39718);
nor U39952 (N_39952,N_39597,N_39694);
or U39953 (N_39953,N_39681,N_39731);
and U39954 (N_39954,N_39641,N_39597);
xor U39955 (N_39955,N_39719,N_39541);
nor U39956 (N_39956,N_39591,N_39698);
nor U39957 (N_39957,N_39696,N_39688);
and U39958 (N_39958,N_39639,N_39739);
nor U39959 (N_39959,N_39743,N_39745);
nand U39960 (N_39960,N_39638,N_39686);
nand U39961 (N_39961,N_39551,N_39595);
nand U39962 (N_39962,N_39639,N_39644);
nand U39963 (N_39963,N_39605,N_39525);
or U39964 (N_39964,N_39576,N_39529);
or U39965 (N_39965,N_39737,N_39644);
xnor U39966 (N_39966,N_39627,N_39629);
xnor U39967 (N_39967,N_39576,N_39548);
nand U39968 (N_39968,N_39691,N_39513);
or U39969 (N_39969,N_39747,N_39556);
and U39970 (N_39970,N_39717,N_39567);
and U39971 (N_39971,N_39734,N_39540);
nand U39972 (N_39972,N_39501,N_39716);
nor U39973 (N_39973,N_39560,N_39550);
nand U39974 (N_39974,N_39658,N_39586);
or U39975 (N_39975,N_39702,N_39672);
nand U39976 (N_39976,N_39688,N_39655);
nor U39977 (N_39977,N_39547,N_39692);
xor U39978 (N_39978,N_39697,N_39540);
or U39979 (N_39979,N_39526,N_39659);
nand U39980 (N_39980,N_39746,N_39711);
and U39981 (N_39981,N_39688,N_39614);
nand U39982 (N_39982,N_39550,N_39724);
nand U39983 (N_39983,N_39593,N_39691);
nand U39984 (N_39984,N_39510,N_39557);
and U39985 (N_39985,N_39715,N_39670);
nor U39986 (N_39986,N_39656,N_39557);
xnor U39987 (N_39987,N_39628,N_39593);
nand U39988 (N_39988,N_39682,N_39592);
and U39989 (N_39989,N_39734,N_39739);
xnor U39990 (N_39990,N_39664,N_39671);
and U39991 (N_39991,N_39676,N_39728);
nand U39992 (N_39992,N_39555,N_39590);
nor U39993 (N_39993,N_39647,N_39689);
xor U39994 (N_39994,N_39720,N_39534);
and U39995 (N_39995,N_39593,N_39655);
xnor U39996 (N_39996,N_39533,N_39749);
xor U39997 (N_39997,N_39572,N_39515);
xor U39998 (N_39998,N_39547,N_39643);
and U39999 (N_39999,N_39511,N_39707);
nor U40000 (N_40000,N_39846,N_39923);
nand U40001 (N_40001,N_39910,N_39807);
or U40002 (N_40002,N_39904,N_39992);
and U40003 (N_40003,N_39890,N_39965);
or U40004 (N_40004,N_39871,N_39840);
nor U40005 (N_40005,N_39841,N_39766);
nor U40006 (N_40006,N_39800,N_39974);
and U40007 (N_40007,N_39945,N_39813);
xor U40008 (N_40008,N_39791,N_39858);
and U40009 (N_40009,N_39801,N_39816);
nand U40010 (N_40010,N_39775,N_39787);
or U40011 (N_40011,N_39872,N_39966);
or U40012 (N_40012,N_39764,N_39919);
or U40013 (N_40013,N_39826,N_39790);
xnor U40014 (N_40014,N_39932,N_39848);
nor U40015 (N_40015,N_39782,N_39753);
or U40016 (N_40016,N_39893,N_39933);
and U40017 (N_40017,N_39950,N_39752);
nand U40018 (N_40018,N_39998,N_39986);
xor U40019 (N_40019,N_39833,N_39759);
xnor U40020 (N_40020,N_39776,N_39984);
nand U40021 (N_40021,N_39810,N_39806);
and U40022 (N_40022,N_39997,N_39903);
and U40023 (N_40023,N_39771,N_39980);
or U40024 (N_40024,N_39856,N_39809);
or U40025 (N_40025,N_39751,N_39795);
xnor U40026 (N_40026,N_39981,N_39934);
and U40027 (N_40027,N_39837,N_39947);
nor U40028 (N_40028,N_39881,N_39915);
nor U40029 (N_40029,N_39769,N_39843);
and U40030 (N_40030,N_39865,N_39835);
xor U40031 (N_40031,N_39943,N_39983);
and U40032 (N_40032,N_39949,N_39773);
or U40033 (N_40033,N_39851,N_39811);
nor U40034 (N_40034,N_39999,N_39867);
nand U40035 (N_40035,N_39798,N_39862);
xor U40036 (N_40036,N_39880,N_39956);
nor U40037 (N_40037,N_39789,N_39887);
nor U40038 (N_40038,N_39948,N_39975);
xnor U40039 (N_40039,N_39939,N_39977);
or U40040 (N_40040,N_39823,N_39886);
nor U40041 (N_40041,N_39818,N_39860);
or U40042 (N_40042,N_39873,N_39828);
or U40043 (N_40043,N_39899,N_39821);
nand U40044 (N_40044,N_39889,N_39778);
nor U40045 (N_40045,N_39854,N_39750);
or U40046 (N_40046,N_39785,N_39829);
nand U40047 (N_40047,N_39946,N_39802);
nand U40048 (N_40048,N_39883,N_39781);
nor U40049 (N_40049,N_39913,N_39849);
nand U40050 (N_40050,N_39885,N_39784);
and U40051 (N_40051,N_39783,N_39879);
nor U40052 (N_40052,N_39814,N_39900);
xor U40053 (N_40053,N_39831,N_39892);
xnor U40054 (N_40054,N_39815,N_39988);
nand U40055 (N_40055,N_39768,N_39960);
and U40056 (N_40056,N_39901,N_39925);
xnor U40057 (N_40057,N_39857,N_39982);
nor U40058 (N_40058,N_39792,N_39779);
nand U40059 (N_40059,N_39930,N_39808);
nor U40060 (N_40060,N_39842,N_39918);
nand U40061 (N_40061,N_39796,N_39874);
nand U40062 (N_40062,N_39898,N_39907);
xor U40063 (N_40063,N_39963,N_39968);
nand U40064 (N_40064,N_39812,N_39911);
nor U40065 (N_40065,N_39869,N_39859);
nor U40066 (N_40066,N_39866,N_39761);
nor U40067 (N_40067,N_39989,N_39928);
nand U40068 (N_40068,N_39969,N_39971);
and U40069 (N_40069,N_39780,N_39820);
and U40070 (N_40070,N_39875,N_39902);
and U40071 (N_40071,N_39952,N_39935);
nand U40072 (N_40072,N_39877,N_39978);
nand U40073 (N_40073,N_39894,N_39944);
or U40074 (N_40074,N_39870,N_39774);
nand U40075 (N_40075,N_39996,N_39805);
or U40076 (N_40076,N_39839,N_39936);
or U40077 (N_40077,N_39868,N_39942);
or U40078 (N_40078,N_39760,N_39845);
nand U40079 (N_40079,N_39850,N_39827);
or U40080 (N_40080,N_39838,N_39804);
nor U40081 (N_40081,N_39767,N_39793);
xor U40082 (N_40082,N_39962,N_39987);
nor U40083 (N_40083,N_39799,N_39991);
nand U40084 (N_40084,N_39803,N_39931);
or U40085 (N_40085,N_39852,N_39884);
nor U40086 (N_40086,N_39921,N_39937);
nand U40087 (N_40087,N_39967,N_39832);
nand U40088 (N_40088,N_39916,N_39959);
nand U40089 (N_40089,N_39878,N_39955);
nor U40090 (N_40090,N_39888,N_39929);
nand U40091 (N_40091,N_39906,N_39770);
and U40092 (N_40092,N_39927,N_39876);
and U40093 (N_40093,N_39788,N_39979);
nor U40094 (N_40094,N_39758,N_39917);
xor U40095 (N_40095,N_39920,N_39822);
nor U40096 (N_40096,N_39957,N_39961);
xor U40097 (N_40097,N_39914,N_39905);
or U40098 (N_40098,N_39861,N_39924);
and U40099 (N_40099,N_39844,N_39972);
nand U40100 (N_40100,N_39976,N_39756);
xor U40101 (N_40101,N_39819,N_39786);
or U40102 (N_40102,N_39762,N_39954);
xor U40103 (N_40103,N_39755,N_39990);
or U40104 (N_40104,N_39964,N_39940);
xnor U40105 (N_40105,N_39825,N_39757);
xor U40106 (N_40106,N_39777,N_39882);
and U40107 (N_40107,N_39863,N_39853);
and U40108 (N_40108,N_39765,N_39834);
xor U40109 (N_40109,N_39985,N_39909);
xnor U40110 (N_40110,N_39855,N_39993);
nand U40111 (N_40111,N_39941,N_39754);
nand U40112 (N_40112,N_39895,N_39973);
nand U40113 (N_40113,N_39938,N_39922);
and U40114 (N_40114,N_39896,N_39830);
xnor U40115 (N_40115,N_39958,N_39995);
xnor U40116 (N_40116,N_39824,N_39763);
nor U40117 (N_40117,N_39953,N_39970);
nand U40118 (N_40118,N_39926,N_39912);
and U40119 (N_40119,N_39908,N_39847);
xnor U40120 (N_40120,N_39836,N_39891);
nand U40121 (N_40121,N_39797,N_39951);
and U40122 (N_40122,N_39994,N_39817);
nor U40123 (N_40123,N_39772,N_39864);
and U40124 (N_40124,N_39897,N_39794);
nor U40125 (N_40125,N_39806,N_39779);
or U40126 (N_40126,N_39782,N_39874);
nand U40127 (N_40127,N_39835,N_39755);
and U40128 (N_40128,N_39846,N_39924);
or U40129 (N_40129,N_39933,N_39783);
xor U40130 (N_40130,N_39757,N_39871);
xnor U40131 (N_40131,N_39952,N_39873);
or U40132 (N_40132,N_39800,N_39924);
nand U40133 (N_40133,N_39989,N_39965);
and U40134 (N_40134,N_39960,N_39760);
nor U40135 (N_40135,N_39948,N_39790);
or U40136 (N_40136,N_39954,N_39779);
xnor U40137 (N_40137,N_39927,N_39790);
nor U40138 (N_40138,N_39977,N_39910);
nand U40139 (N_40139,N_39836,N_39852);
nand U40140 (N_40140,N_39874,N_39818);
xnor U40141 (N_40141,N_39917,N_39880);
nand U40142 (N_40142,N_39934,N_39943);
nand U40143 (N_40143,N_39999,N_39900);
or U40144 (N_40144,N_39840,N_39878);
and U40145 (N_40145,N_39924,N_39963);
nand U40146 (N_40146,N_39899,N_39910);
or U40147 (N_40147,N_39943,N_39946);
xnor U40148 (N_40148,N_39974,N_39802);
xor U40149 (N_40149,N_39899,N_39789);
xnor U40150 (N_40150,N_39872,N_39945);
or U40151 (N_40151,N_39997,N_39843);
or U40152 (N_40152,N_39945,N_39931);
nand U40153 (N_40153,N_39846,N_39779);
or U40154 (N_40154,N_39801,N_39759);
nor U40155 (N_40155,N_39970,N_39850);
or U40156 (N_40156,N_39782,N_39921);
or U40157 (N_40157,N_39926,N_39754);
and U40158 (N_40158,N_39789,N_39787);
nand U40159 (N_40159,N_39831,N_39762);
or U40160 (N_40160,N_39806,N_39924);
nor U40161 (N_40161,N_39893,N_39834);
and U40162 (N_40162,N_39941,N_39809);
or U40163 (N_40163,N_39859,N_39914);
and U40164 (N_40164,N_39794,N_39812);
xnor U40165 (N_40165,N_39994,N_39877);
nand U40166 (N_40166,N_39922,N_39861);
or U40167 (N_40167,N_39862,N_39834);
nand U40168 (N_40168,N_39948,N_39980);
xor U40169 (N_40169,N_39849,N_39923);
nand U40170 (N_40170,N_39906,N_39868);
and U40171 (N_40171,N_39849,N_39863);
nor U40172 (N_40172,N_39965,N_39988);
and U40173 (N_40173,N_39869,N_39804);
xor U40174 (N_40174,N_39840,N_39779);
xor U40175 (N_40175,N_39978,N_39783);
or U40176 (N_40176,N_39883,N_39939);
and U40177 (N_40177,N_39871,N_39944);
and U40178 (N_40178,N_39997,N_39794);
nor U40179 (N_40179,N_39912,N_39758);
nand U40180 (N_40180,N_39816,N_39862);
nand U40181 (N_40181,N_39912,N_39917);
nand U40182 (N_40182,N_39952,N_39980);
and U40183 (N_40183,N_39792,N_39997);
xnor U40184 (N_40184,N_39984,N_39950);
or U40185 (N_40185,N_39757,N_39949);
nand U40186 (N_40186,N_39757,N_39914);
and U40187 (N_40187,N_39871,N_39919);
or U40188 (N_40188,N_39794,N_39830);
nand U40189 (N_40189,N_39934,N_39860);
nand U40190 (N_40190,N_39907,N_39827);
and U40191 (N_40191,N_39833,N_39824);
and U40192 (N_40192,N_39750,N_39995);
and U40193 (N_40193,N_39985,N_39892);
nor U40194 (N_40194,N_39810,N_39981);
and U40195 (N_40195,N_39953,N_39807);
or U40196 (N_40196,N_39753,N_39827);
xor U40197 (N_40197,N_39983,N_39976);
nor U40198 (N_40198,N_39967,N_39956);
nor U40199 (N_40199,N_39900,N_39899);
nor U40200 (N_40200,N_39913,N_39999);
nor U40201 (N_40201,N_39820,N_39854);
or U40202 (N_40202,N_39876,N_39820);
nor U40203 (N_40203,N_39947,N_39783);
nor U40204 (N_40204,N_39814,N_39769);
nand U40205 (N_40205,N_39893,N_39981);
nor U40206 (N_40206,N_39981,N_39932);
xnor U40207 (N_40207,N_39854,N_39773);
and U40208 (N_40208,N_39998,N_39863);
or U40209 (N_40209,N_39886,N_39975);
or U40210 (N_40210,N_39896,N_39871);
nand U40211 (N_40211,N_39977,N_39755);
nand U40212 (N_40212,N_39850,N_39785);
and U40213 (N_40213,N_39763,N_39963);
nand U40214 (N_40214,N_39978,N_39979);
nor U40215 (N_40215,N_39841,N_39878);
nand U40216 (N_40216,N_39916,N_39888);
xor U40217 (N_40217,N_39847,N_39929);
nor U40218 (N_40218,N_39838,N_39839);
xnor U40219 (N_40219,N_39992,N_39976);
nand U40220 (N_40220,N_39808,N_39955);
or U40221 (N_40221,N_39911,N_39789);
nand U40222 (N_40222,N_39855,N_39991);
or U40223 (N_40223,N_39780,N_39798);
or U40224 (N_40224,N_39916,N_39961);
xnor U40225 (N_40225,N_39890,N_39899);
nor U40226 (N_40226,N_39766,N_39797);
and U40227 (N_40227,N_39944,N_39961);
or U40228 (N_40228,N_39869,N_39904);
and U40229 (N_40229,N_39801,N_39893);
nand U40230 (N_40230,N_39933,N_39965);
nor U40231 (N_40231,N_39912,N_39995);
nor U40232 (N_40232,N_39837,N_39930);
and U40233 (N_40233,N_39917,N_39779);
nor U40234 (N_40234,N_39783,N_39949);
or U40235 (N_40235,N_39792,N_39920);
and U40236 (N_40236,N_39843,N_39926);
nand U40237 (N_40237,N_39750,N_39923);
or U40238 (N_40238,N_39873,N_39943);
or U40239 (N_40239,N_39873,N_39928);
nor U40240 (N_40240,N_39839,N_39889);
xnor U40241 (N_40241,N_39803,N_39856);
xor U40242 (N_40242,N_39902,N_39995);
and U40243 (N_40243,N_39888,N_39774);
xor U40244 (N_40244,N_39978,N_39815);
or U40245 (N_40245,N_39792,N_39972);
or U40246 (N_40246,N_39941,N_39935);
nand U40247 (N_40247,N_39923,N_39756);
or U40248 (N_40248,N_39751,N_39871);
xnor U40249 (N_40249,N_39842,N_39922);
or U40250 (N_40250,N_40132,N_40027);
or U40251 (N_40251,N_40015,N_40220);
xor U40252 (N_40252,N_40213,N_40142);
xor U40253 (N_40253,N_40094,N_40036);
xor U40254 (N_40254,N_40209,N_40065);
or U40255 (N_40255,N_40188,N_40055);
and U40256 (N_40256,N_40054,N_40051);
nor U40257 (N_40257,N_40157,N_40138);
xnor U40258 (N_40258,N_40079,N_40146);
and U40259 (N_40259,N_40085,N_40217);
nand U40260 (N_40260,N_40178,N_40204);
or U40261 (N_40261,N_40057,N_40060);
xor U40262 (N_40262,N_40147,N_40042);
or U40263 (N_40263,N_40134,N_40096);
xor U40264 (N_40264,N_40122,N_40189);
nor U40265 (N_40265,N_40007,N_40068);
xor U40266 (N_40266,N_40185,N_40210);
or U40267 (N_40267,N_40212,N_40044);
nor U40268 (N_40268,N_40089,N_40218);
and U40269 (N_40269,N_40140,N_40121);
or U40270 (N_40270,N_40219,N_40227);
nand U40271 (N_40271,N_40012,N_40148);
or U40272 (N_40272,N_40025,N_40017);
xor U40273 (N_40273,N_40013,N_40221);
and U40274 (N_40274,N_40166,N_40098);
nor U40275 (N_40275,N_40206,N_40101);
nor U40276 (N_40276,N_40043,N_40002);
and U40277 (N_40277,N_40056,N_40088);
or U40278 (N_40278,N_40075,N_40129);
nor U40279 (N_40279,N_40248,N_40111);
nand U40280 (N_40280,N_40026,N_40229);
and U40281 (N_40281,N_40164,N_40243);
and U40282 (N_40282,N_40171,N_40153);
and U40283 (N_40283,N_40082,N_40128);
nor U40284 (N_40284,N_40024,N_40064);
and U40285 (N_40285,N_40126,N_40203);
xor U40286 (N_40286,N_40003,N_40176);
and U40287 (N_40287,N_40154,N_40069);
nor U40288 (N_40288,N_40110,N_40021);
nor U40289 (N_40289,N_40087,N_40011);
xor U40290 (N_40290,N_40141,N_40034);
xnor U40291 (N_40291,N_40086,N_40105);
nor U40292 (N_40292,N_40127,N_40097);
and U40293 (N_40293,N_40230,N_40090);
nand U40294 (N_40294,N_40245,N_40237);
and U40295 (N_40295,N_40133,N_40039);
nor U40296 (N_40296,N_40031,N_40067);
nand U40297 (N_40297,N_40196,N_40233);
xor U40298 (N_40298,N_40214,N_40103);
and U40299 (N_40299,N_40181,N_40050);
xor U40300 (N_40300,N_40131,N_40223);
nor U40301 (N_40301,N_40238,N_40143);
xor U40302 (N_40302,N_40118,N_40099);
nand U40303 (N_40303,N_40023,N_40072);
nor U40304 (N_40304,N_40152,N_40063);
nand U40305 (N_40305,N_40194,N_40040);
or U40306 (N_40306,N_40108,N_40113);
xnor U40307 (N_40307,N_40222,N_40074);
nand U40308 (N_40308,N_40041,N_40183);
xnor U40309 (N_40309,N_40006,N_40130);
or U40310 (N_40310,N_40092,N_40163);
nor U40311 (N_40311,N_40192,N_40173);
xnor U40312 (N_40312,N_40215,N_40100);
or U40313 (N_40313,N_40177,N_40018);
and U40314 (N_40314,N_40073,N_40106);
or U40315 (N_40315,N_40200,N_40016);
xnor U40316 (N_40316,N_40193,N_40095);
and U40317 (N_40317,N_40228,N_40124);
and U40318 (N_40318,N_40052,N_40107);
nand U40319 (N_40319,N_40071,N_40249);
nand U40320 (N_40320,N_40145,N_40004);
nor U40321 (N_40321,N_40080,N_40125);
nor U40322 (N_40322,N_40158,N_40165);
nand U40323 (N_40323,N_40116,N_40109);
or U40324 (N_40324,N_40211,N_40208);
xnor U40325 (N_40325,N_40202,N_40058);
and U40326 (N_40326,N_40046,N_40049);
xnor U40327 (N_40327,N_40005,N_40240);
or U40328 (N_40328,N_40084,N_40000);
nor U40329 (N_40329,N_40201,N_40137);
or U40330 (N_40330,N_40235,N_40170);
or U40331 (N_40331,N_40066,N_40241);
and U40332 (N_40332,N_40231,N_40029);
nor U40333 (N_40333,N_40246,N_40115);
nor U40334 (N_40334,N_40186,N_40008);
or U40335 (N_40335,N_40195,N_40184);
nand U40336 (N_40336,N_40150,N_40123);
nand U40337 (N_40337,N_40117,N_40168);
and U40338 (N_40338,N_40236,N_40239);
nand U40339 (N_40339,N_40199,N_40028);
and U40340 (N_40340,N_40216,N_40190);
nor U40341 (N_40341,N_40047,N_40062);
xor U40342 (N_40342,N_40135,N_40032);
and U40343 (N_40343,N_40242,N_40155);
nand U40344 (N_40344,N_40205,N_40119);
nand U40345 (N_40345,N_40224,N_40225);
or U40346 (N_40346,N_40247,N_40179);
nand U40347 (N_40347,N_40120,N_40207);
nand U40348 (N_40348,N_40139,N_40030);
nor U40349 (N_40349,N_40112,N_40197);
nand U40350 (N_40350,N_40059,N_40182);
or U40351 (N_40351,N_40187,N_40180);
or U40352 (N_40352,N_40014,N_40104);
or U40353 (N_40353,N_40151,N_40136);
or U40354 (N_40354,N_40009,N_40114);
xor U40355 (N_40355,N_40078,N_40019);
xnor U40356 (N_40356,N_40091,N_40102);
nand U40357 (N_40357,N_40144,N_40001);
nand U40358 (N_40358,N_40035,N_40232);
nand U40359 (N_40359,N_40077,N_40093);
xor U40360 (N_40360,N_40033,N_40061);
nand U40361 (N_40361,N_40162,N_40172);
xor U40362 (N_40362,N_40198,N_40226);
xor U40363 (N_40363,N_40010,N_40161);
and U40364 (N_40364,N_40081,N_40167);
nor U40365 (N_40365,N_40037,N_40160);
nand U40366 (N_40366,N_40053,N_40083);
or U40367 (N_40367,N_40159,N_40169);
and U40368 (N_40368,N_40174,N_40022);
or U40369 (N_40369,N_40191,N_40038);
nand U40370 (N_40370,N_40244,N_40234);
xnor U40371 (N_40371,N_40149,N_40076);
and U40372 (N_40372,N_40156,N_40020);
nand U40373 (N_40373,N_40048,N_40045);
xnor U40374 (N_40374,N_40070,N_40175);
and U40375 (N_40375,N_40244,N_40004);
xor U40376 (N_40376,N_40142,N_40127);
and U40377 (N_40377,N_40096,N_40006);
nor U40378 (N_40378,N_40080,N_40029);
and U40379 (N_40379,N_40012,N_40221);
nor U40380 (N_40380,N_40060,N_40087);
nand U40381 (N_40381,N_40204,N_40217);
and U40382 (N_40382,N_40022,N_40056);
nand U40383 (N_40383,N_40058,N_40135);
xnor U40384 (N_40384,N_40221,N_40180);
nand U40385 (N_40385,N_40177,N_40092);
and U40386 (N_40386,N_40074,N_40011);
nand U40387 (N_40387,N_40152,N_40195);
nand U40388 (N_40388,N_40033,N_40127);
xor U40389 (N_40389,N_40223,N_40058);
nand U40390 (N_40390,N_40112,N_40100);
nand U40391 (N_40391,N_40092,N_40094);
or U40392 (N_40392,N_40237,N_40155);
nor U40393 (N_40393,N_40170,N_40169);
nor U40394 (N_40394,N_40037,N_40072);
or U40395 (N_40395,N_40099,N_40053);
nand U40396 (N_40396,N_40188,N_40089);
nor U40397 (N_40397,N_40113,N_40155);
nor U40398 (N_40398,N_40041,N_40147);
nor U40399 (N_40399,N_40000,N_40228);
nand U40400 (N_40400,N_40001,N_40074);
and U40401 (N_40401,N_40221,N_40100);
xnor U40402 (N_40402,N_40237,N_40165);
and U40403 (N_40403,N_40117,N_40155);
and U40404 (N_40404,N_40164,N_40129);
nand U40405 (N_40405,N_40063,N_40038);
and U40406 (N_40406,N_40197,N_40126);
xor U40407 (N_40407,N_40171,N_40180);
or U40408 (N_40408,N_40191,N_40032);
nor U40409 (N_40409,N_40111,N_40097);
nand U40410 (N_40410,N_40018,N_40041);
xor U40411 (N_40411,N_40120,N_40186);
or U40412 (N_40412,N_40036,N_40243);
xor U40413 (N_40413,N_40078,N_40001);
xnor U40414 (N_40414,N_40114,N_40092);
or U40415 (N_40415,N_40143,N_40144);
nand U40416 (N_40416,N_40177,N_40044);
xor U40417 (N_40417,N_40027,N_40035);
xnor U40418 (N_40418,N_40168,N_40103);
or U40419 (N_40419,N_40180,N_40126);
or U40420 (N_40420,N_40041,N_40182);
or U40421 (N_40421,N_40129,N_40223);
and U40422 (N_40422,N_40027,N_40230);
nor U40423 (N_40423,N_40217,N_40044);
nand U40424 (N_40424,N_40090,N_40192);
and U40425 (N_40425,N_40041,N_40140);
nor U40426 (N_40426,N_40053,N_40206);
or U40427 (N_40427,N_40115,N_40025);
xnor U40428 (N_40428,N_40085,N_40038);
xnor U40429 (N_40429,N_40247,N_40164);
xor U40430 (N_40430,N_40015,N_40081);
nand U40431 (N_40431,N_40151,N_40168);
or U40432 (N_40432,N_40226,N_40118);
nor U40433 (N_40433,N_40219,N_40228);
nand U40434 (N_40434,N_40128,N_40200);
or U40435 (N_40435,N_40064,N_40131);
nand U40436 (N_40436,N_40148,N_40092);
nor U40437 (N_40437,N_40120,N_40109);
or U40438 (N_40438,N_40052,N_40155);
nor U40439 (N_40439,N_40045,N_40148);
xor U40440 (N_40440,N_40174,N_40000);
nor U40441 (N_40441,N_40131,N_40090);
nor U40442 (N_40442,N_40038,N_40249);
nand U40443 (N_40443,N_40084,N_40152);
or U40444 (N_40444,N_40156,N_40194);
and U40445 (N_40445,N_40210,N_40026);
xor U40446 (N_40446,N_40202,N_40178);
or U40447 (N_40447,N_40204,N_40193);
and U40448 (N_40448,N_40056,N_40008);
and U40449 (N_40449,N_40137,N_40212);
xor U40450 (N_40450,N_40119,N_40040);
xor U40451 (N_40451,N_40074,N_40004);
xor U40452 (N_40452,N_40019,N_40065);
nand U40453 (N_40453,N_40046,N_40014);
xnor U40454 (N_40454,N_40114,N_40040);
nor U40455 (N_40455,N_40018,N_40091);
nand U40456 (N_40456,N_40170,N_40186);
or U40457 (N_40457,N_40060,N_40163);
nand U40458 (N_40458,N_40055,N_40155);
xor U40459 (N_40459,N_40053,N_40006);
nor U40460 (N_40460,N_40001,N_40118);
or U40461 (N_40461,N_40192,N_40189);
xor U40462 (N_40462,N_40125,N_40206);
and U40463 (N_40463,N_40040,N_40135);
or U40464 (N_40464,N_40043,N_40074);
and U40465 (N_40465,N_40163,N_40056);
xor U40466 (N_40466,N_40024,N_40192);
nor U40467 (N_40467,N_40196,N_40042);
and U40468 (N_40468,N_40126,N_40129);
nand U40469 (N_40469,N_40174,N_40135);
nor U40470 (N_40470,N_40039,N_40090);
or U40471 (N_40471,N_40076,N_40000);
or U40472 (N_40472,N_40153,N_40184);
and U40473 (N_40473,N_40083,N_40207);
xnor U40474 (N_40474,N_40196,N_40244);
nor U40475 (N_40475,N_40241,N_40242);
and U40476 (N_40476,N_40147,N_40227);
xnor U40477 (N_40477,N_40224,N_40010);
xor U40478 (N_40478,N_40020,N_40207);
xnor U40479 (N_40479,N_40173,N_40042);
or U40480 (N_40480,N_40191,N_40125);
or U40481 (N_40481,N_40199,N_40220);
nor U40482 (N_40482,N_40050,N_40201);
nand U40483 (N_40483,N_40029,N_40169);
xor U40484 (N_40484,N_40159,N_40188);
nand U40485 (N_40485,N_40047,N_40120);
or U40486 (N_40486,N_40188,N_40213);
nand U40487 (N_40487,N_40155,N_40018);
and U40488 (N_40488,N_40031,N_40216);
or U40489 (N_40489,N_40166,N_40218);
nor U40490 (N_40490,N_40196,N_40069);
nor U40491 (N_40491,N_40197,N_40243);
xnor U40492 (N_40492,N_40223,N_40161);
and U40493 (N_40493,N_40063,N_40233);
or U40494 (N_40494,N_40030,N_40193);
and U40495 (N_40495,N_40012,N_40103);
nand U40496 (N_40496,N_40199,N_40180);
nor U40497 (N_40497,N_40059,N_40107);
xor U40498 (N_40498,N_40144,N_40241);
nand U40499 (N_40499,N_40243,N_40223);
and U40500 (N_40500,N_40388,N_40421);
nor U40501 (N_40501,N_40264,N_40321);
xnor U40502 (N_40502,N_40477,N_40274);
xnor U40503 (N_40503,N_40387,N_40426);
nor U40504 (N_40504,N_40458,N_40309);
or U40505 (N_40505,N_40437,N_40395);
or U40506 (N_40506,N_40286,N_40324);
nand U40507 (N_40507,N_40420,N_40406);
or U40508 (N_40508,N_40339,N_40455);
xnor U40509 (N_40509,N_40391,N_40498);
nand U40510 (N_40510,N_40438,N_40463);
xnor U40511 (N_40511,N_40349,N_40374);
nand U40512 (N_40512,N_40469,N_40460);
nor U40513 (N_40513,N_40356,N_40468);
nand U40514 (N_40514,N_40330,N_40358);
or U40515 (N_40515,N_40450,N_40289);
xnor U40516 (N_40516,N_40383,N_40342);
or U40517 (N_40517,N_40390,N_40490);
and U40518 (N_40518,N_40352,N_40363);
or U40519 (N_40519,N_40250,N_40254);
nor U40520 (N_40520,N_40290,N_40305);
xnor U40521 (N_40521,N_40275,N_40291);
or U40522 (N_40522,N_40351,N_40367);
or U40523 (N_40523,N_40328,N_40268);
or U40524 (N_40524,N_40440,N_40467);
nand U40525 (N_40525,N_40287,N_40435);
xor U40526 (N_40526,N_40439,N_40353);
and U40527 (N_40527,N_40340,N_40251);
or U40528 (N_40528,N_40302,N_40281);
nor U40529 (N_40529,N_40255,N_40313);
or U40530 (N_40530,N_40412,N_40372);
nand U40531 (N_40531,N_40346,N_40292);
nor U40532 (N_40532,N_40447,N_40394);
nor U40533 (N_40533,N_40369,N_40345);
and U40534 (N_40534,N_40419,N_40402);
nand U40535 (N_40535,N_40263,N_40474);
and U40536 (N_40536,N_40496,N_40401);
xnor U40537 (N_40537,N_40441,N_40389);
xnor U40538 (N_40538,N_40259,N_40365);
nor U40539 (N_40539,N_40267,N_40261);
or U40540 (N_40540,N_40444,N_40443);
nor U40541 (N_40541,N_40473,N_40308);
nand U40542 (N_40542,N_40300,N_40491);
xor U40543 (N_40543,N_40271,N_40283);
and U40544 (N_40544,N_40288,N_40445);
nor U40545 (N_40545,N_40347,N_40385);
or U40546 (N_40546,N_40428,N_40379);
nor U40547 (N_40547,N_40269,N_40258);
nor U40548 (N_40548,N_40343,N_40362);
or U40549 (N_40549,N_40284,N_40430);
xnor U40550 (N_40550,N_40465,N_40457);
nand U40551 (N_40551,N_40282,N_40382);
and U40552 (N_40552,N_40252,N_40418);
nand U40553 (N_40553,N_40436,N_40484);
xnor U40554 (N_40554,N_40331,N_40320);
and U40555 (N_40555,N_40427,N_40304);
nor U40556 (N_40556,N_40381,N_40470);
or U40557 (N_40557,N_40480,N_40318);
and U40558 (N_40558,N_40335,N_40376);
xnor U40559 (N_40559,N_40285,N_40314);
nand U40560 (N_40560,N_40280,N_40425);
xnor U40561 (N_40561,N_40273,N_40429);
nand U40562 (N_40562,N_40414,N_40446);
nand U40563 (N_40563,N_40298,N_40262);
nor U40564 (N_40564,N_40393,N_40453);
or U40565 (N_40565,N_40434,N_40378);
and U40566 (N_40566,N_40479,N_40448);
or U40567 (N_40567,N_40296,N_40432);
nor U40568 (N_40568,N_40253,N_40483);
and U40569 (N_40569,N_40497,N_40471);
nor U40570 (N_40570,N_40452,N_40424);
nor U40571 (N_40571,N_40317,N_40404);
xnor U40572 (N_40572,N_40478,N_40431);
nor U40573 (N_40573,N_40310,N_40279);
nor U40574 (N_40574,N_40475,N_40472);
xnor U40575 (N_40575,N_40396,N_40326);
or U40576 (N_40576,N_40486,N_40355);
nor U40577 (N_40577,N_40322,N_40277);
nand U40578 (N_40578,N_40293,N_40299);
xnor U40579 (N_40579,N_40466,N_40265);
xnor U40580 (N_40580,N_40312,N_40333);
nand U40581 (N_40581,N_40357,N_40398);
and U40582 (N_40582,N_40462,N_40433);
or U40583 (N_40583,N_40370,N_40368);
nor U40584 (N_40584,N_40366,N_40482);
nand U40585 (N_40585,N_40332,N_40325);
and U40586 (N_40586,N_40336,N_40454);
xnor U40587 (N_40587,N_40423,N_40295);
and U40588 (N_40588,N_40485,N_40495);
nor U40589 (N_40589,N_40409,N_40413);
nor U40590 (N_40590,N_40371,N_40359);
and U40591 (N_40591,N_40405,N_40461);
xor U40592 (N_40592,N_40407,N_40338);
or U40593 (N_40593,N_40494,N_40492);
nor U40594 (N_40594,N_40459,N_40341);
or U40595 (N_40595,N_40373,N_40306);
xnor U40596 (N_40596,N_40417,N_40400);
nand U40597 (N_40597,N_40377,N_40256);
nor U40598 (N_40598,N_40399,N_40364);
nand U40599 (N_40599,N_40488,N_40294);
or U40600 (N_40600,N_40276,N_40272);
nor U40601 (N_40601,N_40451,N_40323);
nor U40602 (N_40602,N_40456,N_40408);
xor U40603 (N_40603,N_40315,N_40493);
nor U40604 (N_40604,N_40499,N_40386);
nand U40605 (N_40605,N_40360,N_40354);
nand U40606 (N_40606,N_40403,N_40266);
and U40607 (N_40607,N_40487,N_40361);
xnor U40608 (N_40608,N_40442,N_40278);
nor U40609 (N_40609,N_40311,N_40327);
and U40610 (N_40610,N_40375,N_40337);
or U40611 (N_40611,N_40392,N_40449);
or U40612 (N_40612,N_40260,N_40257);
and U40613 (N_40613,N_40380,N_40301);
and U40614 (N_40614,N_40316,N_40411);
nor U40615 (N_40615,N_40319,N_40410);
or U40616 (N_40616,N_40464,N_40348);
nor U40617 (N_40617,N_40481,N_40415);
xnor U40618 (N_40618,N_40422,N_40329);
nor U40619 (N_40619,N_40350,N_40416);
xor U40620 (N_40620,N_40303,N_40334);
xnor U40621 (N_40621,N_40476,N_40489);
nor U40622 (N_40622,N_40397,N_40297);
and U40623 (N_40623,N_40344,N_40384);
nand U40624 (N_40624,N_40270,N_40307);
nor U40625 (N_40625,N_40446,N_40453);
nand U40626 (N_40626,N_40279,N_40381);
nand U40627 (N_40627,N_40409,N_40268);
or U40628 (N_40628,N_40328,N_40411);
and U40629 (N_40629,N_40444,N_40267);
nand U40630 (N_40630,N_40334,N_40484);
and U40631 (N_40631,N_40493,N_40384);
xor U40632 (N_40632,N_40300,N_40281);
and U40633 (N_40633,N_40332,N_40315);
nand U40634 (N_40634,N_40257,N_40294);
xor U40635 (N_40635,N_40346,N_40262);
nand U40636 (N_40636,N_40467,N_40418);
xor U40637 (N_40637,N_40268,N_40316);
or U40638 (N_40638,N_40358,N_40365);
and U40639 (N_40639,N_40264,N_40402);
and U40640 (N_40640,N_40317,N_40430);
or U40641 (N_40641,N_40353,N_40312);
xnor U40642 (N_40642,N_40289,N_40299);
and U40643 (N_40643,N_40458,N_40267);
and U40644 (N_40644,N_40276,N_40312);
or U40645 (N_40645,N_40412,N_40323);
nor U40646 (N_40646,N_40430,N_40474);
or U40647 (N_40647,N_40408,N_40302);
xor U40648 (N_40648,N_40362,N_40410);
nor U40649 (N_40649,N_40494,N_40475);
and U40650 (N_40650,N_40327,N_40486);
xnor U40651 (N_40651,N_40373,N_40260);
nor U40652 (N_40652,N_40286,N_40419);
and U40653 (N_40653,N_40490,N_40268);
and U40654 (N_40654,N_40433,N_40358);
xor U40655 (N_40655,N_40338,N_40347);
or U40656 (N_40656,N_40393,N_40488);
nor U40657 (N_40657,N_40376,N_40476);
or U40658 (N_40658,N_40446,N_40270);
and U40659 (N_40659,N_40288,N_40299);
xor U40660 (N_40660,N_40270,N_40418);
nor U40661 (N_40661,N_40275,N_40286);
or U40662 (N_40662,N_40443,N_40397);
or U40663 (N_40663,N_40448,N_40301);
nand U40664 (N_40664,N_40330,N_40364);
or U40665 (N_40665,N_40427,N_40394);
xor U40666 (N_40666,N_40477,N_40483);
and U40667 (N_40667,N_40497,N_40368);
nor U40668 (N_40668,N_40332,N_40290);
or U40669 (N_40669,N_40474,N_40297);
nor U40670 (N_40670,N_40274,N_40426);
nor U40671 (N_40671,N_40434,N_40442);
or U40672 (N_40672,N_40290,N_40277);
and U40673 (N_40673,N_40375,N_40358);
nor U40674 (N_40674,N_40476,N_40419);
and U40675 (N_40675,N_40411,N_40433);
or U40676 (N_40676,N_40350,N_40258);
and U40677 (N_40677,N_40307,N_40364);
or U40678 (N_40678,N_40455,N_40416);
xnor U40679 (N_40679,N_40361,N_40272);
xnor U40680 (N_40680,N_40418,N_40365);
and U40681 (N_40681,N_40285,N_40355);
nand U40682 (N_40682,N_40288,N_40413);
and U40683 (N_40683,N_40432,N_40305);
nand U40684 (N_40684,N_40464,N_40435);
nand U40685 (N_40685,N_40294,N_40464);
nor U40686 (N_40686,N_40324,N_40394);
nor U40687 (N_40687,N_40313,N_40450);
or U40688 (N_40688,N_40309,N_40437);
xor U40689 (N_40689,N_40255,N_40381);
xnor U40690 (N_40690,N_40304,N_40283);
or U40691 (N_40691,N_40377,N_40392);
xor U40692 (N_40692,N_40377,N_40366);
xnor U40693 (N_40693,N_40445,N_40337);
xnor U40694 (N_40694,N_40290,N_40433);
xor U40695 (N_40695,N_40366,N_40382);
nor U40696 (N_40696,N_40387,N_40465);
or U40697 (N_40697,N_40354,N_40464);
or U40698 (N_40698,N_40418,N_40309);
or U40699 (N_40699,N_40440,N_40386);
xnor U40700 (N_40700,N_40458,N_40405);
xor U40701 (N_40701,N_40446,N_40468);
or U40702 (N_40702,N_40282,N_40383);
xnor U40703 (N_40703,N_40264,N_40482);
nand U40704 (N_40704,N_40327,N_40405);
or U40705 (N_40705,N_40422,N_40454);
nor U40706 (N_40706,N_40260,N_40255);
nand U40707 (N_40707,N_40317,N_40429);
nand U40708 (N_40708,N_40497,N_40461);
xor U40709 (N_40709,N_40390,N_40443);
nand U40710 (N_40710,N_40285,N_40403);
nand U40711 (N_40711,N_40370,N_40438);
nor U40712 (N_40712,N_40475,N_40435);
xor U40713 (N_40713,N_40428,N_40269);
xnor U40714 (N_40714,N_40263,N_40337);
nor U40715 (N_40715,N_40358,N_40329);
nor U40716 (N_40716,N_40451,N_40474);
and U40717 (N_40717,N_40288,N_40268);
and U40718 (N_40718,N_40474,N_40435);
and U40719 (N_40719,N_40295,N_40324);
and U40720 (N_40720,N_40296,N_40361);
and U40721 (N_40721,N_40490,N_40330);
and U40722 (N_40722,N_40286,N_40471);
xor U40723 (N_40723,N_40358,N_40356);
or U40724 (N_40724,N_40353,N_40279);
and U40725 (N_40725,N_40276,N_40265);
or U40726 (N_40726,N_40456,N_40436);
xnor U40727 (N_40727,N_40345,N_40278);
or U40728 (N_40728,N_40447,N_40354);
or U40729 (N_40729,N_40459,N_40283);
or U40730 (N_40730,N_40478,N_40330);
or U40731 (N_40731,N_40427,N_40415);
nor U40732 (N_40732,N_40384,N_40418);
nand U40733 (N_40733,N_40277,N_40425);
or U40734 (N_40734,N_40436,N_40427);
and U40735 (N_40735,N_40457,N_40475);
xnor U40736 (N_40736,N_40331,N_40277);
nand U40737 (N_40737,N_40292,N_40252);
nor U40738 (N_40738,N_40259,N_40254);
xnor U40739 (N_40739,N_40372,N_40253);
nand U40740 (N_40740,N_40284,N_40410);
nand U40741 (N_40741,N_40326,N_40263);
xnor U40742 (N_40742,N_40275,N_40432);
nand U40743 (N_40743,N_40280,N_40369);
nor U40744 (N_40744,N_40274,N_40281);
nand U40745 (N_40745,N_40352,N_40406);
xor U40746 (N_40746,N_40318,N_40295);
nor U40747 (N_40747,N_40401,N_40355);
and U40748 (N_40748,N_40333,N_40387);
and U40749 (N_40749,N_40486,N_40291);
and U40750 (N_40750,N_40571,N_40509);
nor U40751 (N_40751,N_40671,N_40656);
xnor U40752 (N_40752,N_40582,N_40738);
nor U40753 (N_40753,N_40601,N_40732);
xnor U40754 (N_40754,N_40619,N_40520);
xnor U40755 (N_40755,N_40537,N_40620);
and U40756 (N_40756,N_40706,N_40640);
or U40757 (N_40757,N_40668,N_40748);
and U40758 (N_40758,N_40648,N_40585);
xnor U40759 (N_40759,N_40575,N_40628);
nand U40760 (N_40760,N_40641,N_40680);
or U40761 (N_40761,N_40534,N_40697);
nand U40762 (N_40762,N_40649,N_40610);
nand U40763 (N_40763,N_40744,N_40699);
and U40764 (N_40764,N_40664,N_40580);
xnor U40765 (N_40765,N_40579,N_40665);
xnor U40766 (N_40766,N_40702,N_40513);
xor U40767 (N_40767,N_40530,N_40677);
nand U40768 (N_40768,N_40675,N_40511);
nand U40769 (N_40769,N_40714,N_40632);
nor U40770 (N_40770,N_40540,N_40647);
xor U40771 (N_40771,N_40569,N_40586);
nand U40772 (N_40772,N_40507,N_40578);
and U40773 (N_40773,N_40704,N_40521);
xnor U40774 (N_40774,N_40636,N_40556);
nor U40775 (N_40775,N_40514,N_40595);
or U40776 (N_40776,N_40739,N_40735);
and U40777 (N_40777,N_40560,N_40554);
xnor U40778 (N_40778,N_40599,N_40631);
and U40779 (N_40779,N_40666,N_40613);
nand U40780 (N_40780,N_40519,N_40728);
or U40781 (N_40781,N_40550,N_40701);
xnor U40782 (N_40782,N_40713,N_40532);
nor U40783 (N_40783,N_40724,N_40542);
or U40784 (N_40784,N_40705,N_40510);
nor U40785 (N_40785,N_40626,N_40673);
and U40786 (N_40786,N_40747,N_40711);
nand U40787 (N_40787,N_40527,N_40546);
nand U40788 (N_40788,N_40726,N_40564);
xnor U40789 (N_40789,N_40691,N_40515);
nor U40790 (N_40790,N_40574,N_40525);
nand U40791 (N_40791,N_40565,N_40722);
and U40792 (N_40792,N_40531,N_40555);
nor U40793 (N_40793,N_40566,N_40584);
and U40794 (N_40794,N_40616,N_40737);
or U40795 (N_40795,N_40541,N_40740);
and U40796 (N_40796,N_40674,N_40643);
xnor U40797 (N_40797,N_40516,N_40591);
and U40798 (N_40798,N_40553,N_40588);
nor U40799 (N_40799,N_40590,N_40716);
or U40800 (N_40800,N_40614,N_40681);
xor U40801 (N_40801,N_40634,N_40551);
or U40802 (N_40802,N_40646,N_40710);
nand U40803 (N_40803,N_40608,N_40504);
or U40804 (N_40804,N_40611,N_40659);
and U40805 (N_40805,N_40749,N_40559);
xor U40806 (N_40806,N_40695,N_40615);
nand U40807 (N_40807,N_40743,N_40645);
nand U40808 (N_40808,N_40624,N_40644);
xor U40809 (N_40809,N_40731,N_40625);
xor U40810 (N_40810,N_40598,N_40517);
nand U40811 (N_40811,N_40725,N_40745);
nand U40812 (N_40812,N_40686,N_40600);
and U40813 (N_40813,N_40729,N_40720);
or U40814 (N_40814,N_40623,N_40606);
or U40815 (N_40815,N_40633,N_40561);
nand U40816 (N_40816,N_40672,N_40662);
nand U40817 (N_40817,N_40661,N_40573);
or U40818 (N_40818,N_40607,N_40593);
or U40819 (N_40819,N_40501,N_40602);
nor U40820 (N_40820,N_40552,N_40654);
xor U40821 (N_40821,N_40736,N_40694);
and U40822 (N_40822,N_40679,N_40651);
or U40823 (N_40823,N_40549,N_40508);
or U40824 (N_40824,N_40529,N_40597);
nand U40825 (N_40825,N_40690,N_40503);
and U40826 (N_40826,N_40518,N_40653);
xor U40827 (N_40827,N_40577,N_40627);
or U40828 (N_40828,N_40708,N_40689);
nand U40829 (N_40829,N_40715,N_40730);
xnor U40830 (N_40830,N_40558,N_40719);
and U40831 (N_40831,N_40660,N_40594);
nor U40832 (N_40832,N_40563,N_40617);
nor U40833 (N_40833,N_40655,N_40570);
nor U40834 (N_40834,N_40548,N_40533);
xnor U40835 (N_40835,N_40592,N_40603);
or U40836 (N_40836,N_40547,N_40717);
nand U40837 (N_40837,N_40639,N_40630);
and U40838 (N_40838,N_40536,N_40670);
nand U40839 (N_40839,N_40688,N_40746);
xor U40840 (N_40840,N_40657,N_40696);
nand U40841 (N_40841,N_40721,N_40635);
xor U40842 (N_40842,N_40581,N_40621);
nand U40843 (N_40843,N_40572,N_40663);
or U40844 (N_40844,N_40589,N_40524);
or U40845 (N_40845,N_40687,N_40596);
xnor U40846 (N_40846,N_40568,N_40723);
xor U40847 (N_40847,N_40742,N_40678);
nor U40848 (N_40848,N_40733,N_40604);
nand U40849 (N_40849,N_40622,N_40502);
or U40850 (N_40850,N_40583,N_40512);
or U40851 (N_40851,N_40684,N_40506);
or U40852 (N_40852,N_40576,N_40727);
nor U40853 (N_40853,N_40605,N_40698);
xnor U40854 (N_40854,N_40652,N_40676);
nor U40855 (N_40855,N_40526,N_40500);
nand U40856 (N_40856,N_40629,N_40567);
nand U40857 (N_40857,N_40692,N_40562);
nor U40858 (N_40858,N_40650,N_40523);
xnor U40859 (N_40859,N_40612,N_40557);
nor U40860 (N_40860,N_40703,N_40544);
nand U40861 (N_40861,N_40528,N_40505);
nand U40862 (N_40862,N_40539,N_40709);
or U40863 (N_40863,N_40538,N_40638);
nor U40864 (N_40864,N_40707,N_40618);
xor U40865 (N_40865,N_40522,N_40683);
nor U40866 (N_40866,N_40682,N_40642);
xor U40867 (N_40867,N_40658,N_40535);
xnor U40868 (N_40868,N_40587,N_40693);
nor U40869 (N_40869,N_40712,N_40685);
or U40870 (N_40870,N_40637,N_40669);
and U40871 (N_40871,N_40543,N_40741);
or U40872 (N_40872,N_40609,N_40700);
nand U40873 (N_40873,N_40545,N_40718);
and U40874 (N_40874,N_40734,N_40667);
and U40875 (N_40875,N_40673,N_40540);
and U40876 (N_40876,N_40543,N_40739);
nor U40877 (N_40877,N_40592,N_40723);
nor U40878 (N_40878,N_40639,N_40624);
nand U40879 (N_40879,N_40557,N_40619);
nor U40880 (N_40880,N_40508,N_40593);
nor U40881 (N_40881,N_40629,N_40714);
nand U40882 (N_40882,N_40616,N_40745);
nor U40883 (N_40883,N_40520,N_40625);
xor U40884 (N_40884,N_40630,N_40560);
and U40885 (N_40885,N_40671,N_40746);
nor U40886 (N_40886,N_40617,N_40644);
and U40887 (N_40887,N_40585,N_40638);
or U40888 (N_40888,N_40737,N_40619);
nand U40889 (N_40889,N_40721,N_40556);
and U40890 (N_40890,N_40539,N_40650);
nand U40891 (N_40891,N_40556,N_40626);
or U40892 (N_40892,N_40576,N_40703);
or U40893 (N_40893,N_40615,N_40735);
and U40894 (N_40894,N_40612,N_40627);
nand U40895 (N_40895,N_40743,N_40538);
or U40896 (N_40896,N_40617,N_40742);
nor U40897 (N_40897,N_40682,N_40531);
xnor U40898 (N_40898,N_40739,N_40566);
or U40899 (N_40899,N_40571,N_40670);
nor U40900 (N_40900,N_40532,N_40700);
and U40901 (N_40901,N_40663,N_40721);
or U40902 (N_40902,N_40656,N_40549);
and U40903 (N_40903,N_40646,N_40507);
nand U40904 (N_40904,N_40520,N_40540);
xor U40905 (N_40905,N_40528,N_40560);
nand U40906 (N_40906,N_40736,N_40668);
nand U40907 (N_40907,N_40644,N_40726);
xor U40908 (N_40908,N_40533,N_40512);
nor U40909 (N_40909,N_40600,N_40735);
xnor U40910 (N_40910,N_40618,N_40572);
xor U40911 (N_40911,N_40699,N_40671);
xor U40912 (N_40912,N_40531,N_40705);
xnor U40913 (N_40913,N_40728,N_40632);
and U40914 (N_40914,N_40636,N_40672);
nor U40915 (N_40915,N_40537,N_40541);
or U40916 (N_40916,N_40701,N_40634);
or U40917 (N_40917,N_40623,N_40617);
nor U40918 (N_40918,N_40730,N_40747);
and U40919 (N_40919,N_40736,N_40561);
xor U40920 (N_40920,N_40731,N_40722);
and U40921 (N_40921,N_40746,N_40545);
xor U40922 (N_40922,N_40579,N_40705);
and U40923 (N_40923,N_40577,N_40564);
and U40924 (N_40924,N_40546,N_40638);
nand U40925 (N_40925,N_40506,N_40549);
xnor U40926 (N_40926,N_40564,N_40663);
or U40927 (N_40927,N_40710,N_40531);
or U40928 (N_40928,N_40532,N_40729);
xnor U40929 (N_40929,N_40693,N_40664);
nor U40930 (N_40930,N_40608,N_40741);
and U40931 (N_40931,N_40703,N_40639);
nor U40932 (N_40932,N_40591,N_40529);
nand U40933 (N_40933,N_40622,N_40653);
or U40934 (N_40934,N_40735,N_40650);
and U40935 (N_40935,N_40536,N_40502);
xnor U40936 (N_40936,N_40740,N_40679);
and U40937 (N_40937,N_40719,N_40614);
nor U40938 (N_40938,N_40745,N_40507);
nand U40939 (N_40939,N_40737,N_40696);
or U40940 (N_40940,N_40723,N_40510);
xnor U40941 (N_40941,N_40739,N_40540);
xnor U40942 (N_40942,N_40578,N_40566);
and U40943 (N_40943,N_40652,N_40615);
xnor U40944 (N_40944,N_40632,N_40691);
or U40945 (N_40945,N_40658,N_40588);
and U40946 (N_40946,N_40589,N_40695);
or U40947 (N_40947,N_40739,N_40720);
xnor U40948 (N_40948,N_40529,N_40652);
xnor U40949 (N_40949,N_40597,N_40596);
nor U40950 (N_40950,N_40647,N_40557);
and U40951 (N_40951,N_40527,N_40613);
and U40952 (N_40952,N_40688,N_40564);
xor U40953 (N_40953,N_40575,N_40515);
nor U40954 (N_40954,N_40513,N_40654);
or U40955 (N_40955,N_40741,N_40501);
and U40956 (N_40956,N_40554,N_40548);
nor U40957 (N_40957,N_40572,N_40659);
xor U40958 (N_40958,N_40721,N_40550);
xnor U40959 (N_40959,N_40633,N_40543);
or U40960 (N_40960,N_40706,N_40518);
and U40961 (N_40961,N_40675,N_40707);
and U40962 (N_40962,N_40698,N_40659);
or U40963 (N_40963,N_40677,N_40690);
xor U40964 (N_40964,N_40729,N_40523);
nor U40965 (N_40965,N_40501,N_40535);
or U40966 (N_40966,N_40714,N_40532);
or U40967 (N_40967,N_40536,N_40539);
nor U40968 (N_40968,N_40727,N_40509);
nand U40969 (N_40969,N_40621,N_40623);
nor U40970 (N_40970,N_40738,N_40598);
and U40971 (N_40971,N_40623,N_40639);
or U40972 (N_40972,N_40656,N_40681);
and U40973 (N_40973,N_40582,N_40658);
nand U40974 (N_40974,N_40648,N_40546);
or U40975 (N_40975,N_40538,N_40723);
nand U40976 (N_40976,N_40621,N_40625);
xor U40977 (N_40977,N_40605,N_40703);
nor U40978 (N_40978,N_40503,N_40686);
or U40979 (N_40979,N_40591,N_40519);
or U40980 (N_40980,N_40712,N_40574);
nor U40981 (N_40981,N_40547,N_40721);
nor U40982 (N_40982,N_40522,N_40582);
xor U40983 (N_40983,N_40620,N_40558);
xnor U40984 (N_40984,N_40718,N_40705);
xnor U40985 (N_40985,N_40528,N_40671);
nand U40986 (N_40986,N_40650,N_40561);
nand U40987 (N_40987,N_40621,N_40669);
xor U40988 (N_40988,N_40710,N_40656);
xnor U40989 (N_40989,N_40615,N_40578);
or U40990 (N_40990,N_40661,N_40509);
nor U40991 (N_40991,N_40675,N_40589);
nand U40992 (N_40992,N_40517,N_40707);
nand U40993 (N_40993,N_40533,N_40570);
and U40994 (N_40994,N_40595,N_40506);
nor U40995 (N_40995,N_40745,N_40523);
nand U40996 (N_40996,N_40743,N_40728);
nand U40997 (N_40997,N_40512,N_40684);
nand U40998 (N_40998,N_40680,N_40577);
nand U40999 (N_40999,N_40670,N_40729);
or U41000 (N_41000,N_40975,N_40937);
nor U41001 (N_41001,N_40934,N_40930);
nand U41002 (N_41002,N_40892,N_40883);
nor U41003 (N_41003,N_40756,N_40905);
and U41004 (N_41004,N_40970,N_40872);
nor U41005 (N_41005,N_40847,N_40819);
nor U41006 (N_41006,N_40920,N_40950);
and U41007 (N_41007,N_40820,N_40759);
xor U41008 (N_41008,N_40923,N_40757);
and U41009 (N_41009,N_40853,N_40781);
and U41010 (N_41010,N_40981,N_40867);
nand U41011 (N_41011,N_40809,N_40871);
xor U41012 (N_41012,N_40824,N_40774);
or U41013 (N_41013,N_40861,N_40878);
and U41014 (N_41014,N_40944,N_40841);
and U41015 (N_41015,N_40885,N_40795);
or U41016 (N_41016,N_40904,N_40899);
xor U41017 (N_41017,N_40791,N_40895);
xor U41018 (N_41018,N_40833,N_40898);
nor U41019 (N_41019,N_40831,N_40973);
and U41020 (N_41020,N_40894,N_40976);
nor U41021 (N_41021,N_40974,N_40830);
nor U41022 (N_41022,N_40818,N_40764);
and U41023 (N_41023,N_40804,N_40760);
xnor U41024 (N_41024,N_40928,N_40953);
or U41025 (N_41025,N_40915,N_40787);
and U41026 (N_41026,N_40960,N_40860);
xor U41027 (N_41027,N_40826,N_40812);
nor U41028 (N_41028,N_40992,N_40922);
and U41029 (N_41029,N_40941,N_40825);
nor U41030 (N_41030,N_40963,N_40838);
nor U41031 (N_41031,N_40879,N_40806);
nor U41032 (N_41032,N_40877,N_40768);
and U41033 (N_41033,N_40888,N_40817);
nor U41034 (N_41034,N_40775,N_40897);
or U41035 (N_41035,N_40839,N_40776);
and U41036 (N_41036,N_40751,N_40750);
nand U41037 (N_41037,N_40926,N_40880);
or U41038 (N_41038,N_40837,N_40956);
or U41039 (N_41039,N_40789,N_40990);
nor U41040 (N_41040,N_40844,N_40802);
and U41041 (N_41041,N_40790,N_40961);
and U41042 (N_41042,N_40783,N_40942);
and U41043 (N_41043,N_40908,N_40996);
nor U41044 (N_41044,N_40785,N_40929);
or U41045 (N_41045,N_40868,N_40932);
xnor U41046 (N_41046,N_40952,N_40919);
xor U41047 (N_41047,N_40921,N_40840);
or U41048 (N_41048,N_40752,N_40805);
nand U41049 (N_41049,N_40913,N_40858);
xnor U41050 (N_41050,N_40792,N_40900);
nand U41051 (N_41051,N_40784,N_40829);
nor U41052 (N_41052,N_40959,N_40855);
or U41053 (N_41053,N_40814,N_40991);
nand U41054 (N_41054,N_40978,N_40857);
nor U41055 (N_41055,N_40874,N_40995);
nand U41056 (N_41056,N_40999,N_40964);
or U41057 (N_41057,N_40917,N_40886);
or U41058 (N_41058,N_40754,N_40997);
nand U41059 (N_41059,N_40912,N_40933);
xor U41060 (N_41060,N_40935,N_40916);
or U41061 (N_41061,N_40778,N_40994);
nor U41062 (N_41062,N_40786,N_40862);
nand U41063 (N_41063,N_40769,N_40870);
xor U41064 (N_41064,N_40998,N_40985);
and U41065 (N_41065,N_40815,N_40780);
or U41066 (N_41066,N_40755,N_40796);
or U41067 (N_41067,N_40821,N_40763);
or U41068 (N_41068,N_40967,N_40850);
nor U41069 (N_41069,N_40906,N_40864);
nand U41070 (N_41070,N_40810,N_40925);
nand U41071 (N_41071,N_40852,N_40771);
and U41072 (N_41072,N_40955,N_40972);
or U41073 (N_41073,N_40758,N_40836);
xnor U41074 (N_41074,N_40968,N_40827);
and U41075 (N_41075,N_40834,N_40986);
and U41076 (N_41076,N_40987,N_40966);
or U41077 (N_41077,N_40767,N_40958);
or U41078 (N_41078,N_40842,N_40993);
xor U41079 (N_41079,N_40803,N_40800);
and U41080 (N_41080,N_40984,N_40766);
or U41081 (N_41081,N_40938,N_40980);
xor U41082 (N_41082,N_40924,N_40801);
or U41083 (N_41083,N_40949,N_40969);
and U41084 (N_41084,N_40909,N_40946);
and U41085 (N_41085,N_40765,N_40873);
and U41086 (N_41086,N_40798,N_40943);
or U41087 (N_41087,N_40761,N_40927);
or U41088 (N_41088,N_40843,N_40965);
nand U41089 (N_41089,N_40945,N_40807);
or U41090 (N_41090,N_40910,N_40866);
nor U41091 (N_41091,N_40859,N_40782);
nand U41092 (N_41092,N_40887,N_40988);
nor U41093 (N_41093,N_40890,N_40939);
nor U41094 (N_41094,N_40957,N_40875);
and U41095 (N_41095,N_40936,N_40777);
nor U41096 (N_41096,N_40848,N_40876);
xnor U41097 (N_41097,N_40889,N_40779);
or U41098 (N_41098,N_40903,N_40891);
or U41099 (N_41099,N_40753,N_40822);
nor U41100 (N_41100,N_40989,N_40799);
nor U41101 (N_41101,N_40901,N_40845);
or U41102 (N_41102,N_40951,N_40856);
xnor U41103 (N_41103,N_40911,N_40907);
xnor U41104 (N_41104,N_40797,N_40811);
xor U41105 (N_41105,N_40948,N_40971);
or U41106 (N_41106,N_40849,N_40881);
and U41107 (N_41107,N_40914,N_40931);
and U41108 (N_41108,N_40770,N_40773);
or U41109 (N_41109,N_40954,N_40828);
or U41110 (N_41110,N_40947,N_40962);
and U41111 (N_41111,N_40832,N_40808);
nor U41112 (N_41112,N_40846,N_40882);
nand U41113 (N_41113,N_40918,N_40979);
xnor U41114 (N_41114,N_40793,N_40982);
or U41115 (N_41115,N_40896,N_40902);
nor U41116 (N_41116,N_40977,N_40788);
nand U41117 (N_41117,N_40772,N_40813);
and U41118 (N_41118,N_40884,N_40869);
and U41119 (N_41119,N_40893,N_40823);
nor U41120 (N_41120,N_40863,N_40816);
nor U41121 (N_41121,N_40940,N_40794);
nor U41122 (N_41122,N_40854,N_40851);
nor U41123 (N_41123,N_40835,N_40983);
xor U41124 (N_41124,N_40762,N_40865);
or U41125 (N_41125,N_40754,N_40782);
nand U41126 (N_41126,N_40785,N_40891);
nor U41127 (N_41127,N_40979,N_40780);
xnor U41128 (N_41128,N_40826,N_40923);
nand U41129 (N_41129,N_40891,N_40981);
and U41130 (N_41130,N_40754,N_40774);
nand U41131 (N_41131,N_40803,N_40875);
nand U41132 (N_41132,N_40901,N_40788);
and U41133 (N_41133,N_40767,N_40921);
xnor U41134 (N_41134,N_40797,N_40947);
and U41135 (N_41135,N_40957,N_40946);
or U41136 (N_41136,N_40861,N_40811);
xnor U41137 (N_41137,N_40770,N_40778);
nor U41138 (N_41138,N_40908,N_40799);
and U41139 (N_41139,N_40996,N_40901);
xor U41140 (N_41140,N_40846,N_40792);
and U41141 (N_41141,N_40915,N_40831);
xor U41142 (N_41142,N_40796,N_40999);
and U41143 (N_41143,N_40883,N_40917);
xor U41144 (N_41144,N_40755,N_40812);
or U41145 (N_41145,N_40971,N_40872);
nand U41146 (N_41146,N_40985,N_40968);
or U41147 (N_41147,N_40799,N_40872);
xnor U41148 (N_41148,N_40836,N_40869);
or U41149 (N_41149,N_40856,N_40996);
nand U41150 (N_41150,N_40990,N_40760);
nand U41151 (N_41151,N_40843,N_40804);
or U41152 (N_41152,N_40751,N_40875);
nand U41153 (N_41153,N_40981,N_40773);
xor U41154 (N_41154,N_40779,N_40958);
or U41155 (N_41155,N_40909,N_40788);
or U41156 (N_41156,N_40825,N_40802);
or U41157 (N_41157,N_40859,N_40999);
and U41158 (N_41158,N_40981,N_40840);
or U41159 (N_41159,N_40811,N_40884);
nor U41160 (N_41160,N_40973,N_40965);
nand U41161 (N_41161,N_40762,N_40879);
nand U41162 (N_41162,N_40987,N_40996);
xnor U41163 (N_41163,N_40856,N_40997);
nand U41164 (N_41164,N_40932,N_40894);
xor U41165 (N_41165,N_40805,N_40896);
xnor U41166 (N_41166,N_40971,N_40843);
nand U41167 (N_41167,N_40856,N_40962);
xnor U41168 (N_41168,N_40894,N_40979);
and U41169 (N_41169,N_40989,N_40896);
and U41170 (N_41170,N_40755,N_40969);
and U41171 (N_41171,N_40900,N_40870);
xor U41172 (N_41172,N_40933,N_40892);
or U41173 (N_41173,N_40811,N_40755);
nor U41174 (N_41174,N_40871,N_40860);
and U41175 (N_41175,N_40893,N_40818);
or U41176 (N_41176,N_40842,N_40780);
nor U41177 (N_41177,N_40964,N_40797);
nor U41178 (N_41178,N_40750,N_40983);
xnor U41179 (N_41179,N_40760,N_40772);
nor U41180 (N_41180,N_40905,N_40941);
or U41181 (N_41181,N_40773,N_40779);
nand U41182 (N_41182,N_40933,N_40921);
xnor U41183 (N_41183,N_40906,N_40990);
or U41184 (N_41184,N_40932,N_40909);
nand U41185 (N_41185,N_40823,N_40905);
xor U41186 (N_41186,N_40859,N_40934);
nor U41187 (N_41187,N_40978,N_40869);
nor U41188 (N_41188,N_40834,N_40761);
nor U41189 (N_41189,N_40750,N_40861);
xor U41190 (N_41190,N_40853,N_40966);
xor U41191 (N_41191,N_40843,N_40907);
and U41192 (N_41192,N_40870,N_40925);
or U41193 (N_41193,N_40932,N_40895);
xnor U41194 (N_41194,N_40927,N_40991);
and U41195 (N_41195,N_40832,N_40904);
nand U41196 (N_41196,N_40788,N_40808);
nand U41197 (N_41197,N_40995,N_40923);
and U41198 (N_41198,N_40867,N_40879);
or U41199 (N_41199,N_40913,N_40898);
and U41200 (N_41200,N_40917,N_40876);
or U41201 (N_41201,N_40978,N_40780);
nand U41202 (N_41202,N_40823,N_40910);
nor U41203 (N_41203,N_40974,N_40765);
nand U41204 (N_41204,N_40759,N_40758);
and U41205 (N_41205,N_40934,N_40784);
or U41206 (N_41206,N_40845,N_40775);
or U41207 (N_41207,N_40833,N_40892);
nor U41208 (N_41208,N_40857,N_40931);
or U41209 (N_41209,N_40863,N_40754);
nand U41210 (N_41210,N_40918,N_40769);
or U41211 (N_41211,N_40817,N_40826);
xor U41212 (N_41212,N_40899,N_40970);
xnor U41213 (N_41213,N_40893,N_40972);
xnor U41214 (N_41214,N_40990,N_40898);
xor U41215 (N_41215,N_40873,N_40904);
and U41216 (N_41216,N_40902,N_40757);
or U41217 (N_41217,N_40894,N_40938);
nor U41218 (N_41218,N_40862,N_40918);
and U41219 (N_41219,N_40906,N_40773);
nand U41220 (N_41220,N_40981,N_40882);
and U41221 (N_41221,N_40953,N_40821);
and U41222 (N_41222,N_40837,N_40959);
nand U41223 (N_41223,N_40774,N_40977);
nand U41224 (N_41224,N_40926,N_40894);
xor U41225 (N_41225,N_40870,N_40818);
and U41226 (N_41226,N_40867,N_40942);
nor U41227 (N_41227,N_40907,N_40852);
nand U41228 (N_41228,N_40838,N_40789);
or U41229 (N_41229,N_40773,N_40997);
and U41230 (N_41230,N_40761,N_40756);
nand U41231 (N_41231,N_40841,N_40825);
or U41232 (N_41232,N_40872,N_40899);
and U41233 (N_41233,N_40995,N_40769);
or U41234 (N_41234,N_40875,N_40964);
and U41235 (N_41235,N_40886,N_40912);
and U41236 (N_41236,N_40771,N_40923);
nor U41237 (N_41237,N_40802,N_40909);
nand U41238 (N_41238,N_40955,N_40834);
nand U41239 (N_41239,N_40870,N_40919);
or U41240 (N_41240,N_40855,N_40977);
or U41241 (N_41241,N_40817,N_40911);
xor U41242 (N_41242,N_40886,N_40962);
nand U41243 (N_41243,N_40944,N_40785);
nand U41244 (N_41244,N_40812,N_40842);
nor U41245 (N_41245,N_40778,N_40974);
nor U41246 (N_41246,N_40910,N_40766);
and U41247 (N_41247,N_40872,N_40868);
xor U41248 (N_41248,N_40850,N_40874);
or U41249 (N_41249,N_40927,N_40875);
xor U41250 (N_41250,N_41039,N_41021);
xor U41251 (N_41251,N_41203,N_41199);
xnor U41252 (N_41252,N_41042,N_41201);
nor U41253 (N_41253,N_41006,N_41023);
nor U41254 (N_41254,N_41118,N_41171);
nand U41255 (N_41255,N_41078,N_41004);
nor U41256 (N_41256,N_41168,N_41073);
xor U41257 (N_41257,N_41018,N_41154);
nand U41258 (N_41258,N_41147,N_41099);
nor U41259 (N_41259,N_41238,N_41156);
or U41260 (N_41260,N_41145,N_41107);
or U41261 (N_41261,N_41207,N_41182);
nor U41262 (N_41262,N_41159,N_41214);
and U41263 (N_41263,N_41114,N_41081);
and U41264 (N_41264,N_41197,N_41029);
nand U41265 (N_41265,N_41053,N_41057);
or U41266 (N_41266,N_41041,N_41067);
or U41267 (N_41267,N_41125,N_41005);
xnor U41268 (N_41268,N_41208,N_41120);
xnor U41269 (N_41269,N_41216,N_41229);
or U41270 (N_41270,N_41150,N_41158);
nand U41271 (N_41271,N_41247,N_41188);
xor U41272 (N_41272,N_41065,N_41213);
and U41273 (N_41273,N_41079,N_41091);
xnor U41274 (N_41274,N_41027,N_41051);
or U41275 (N_41275,N_41024,N_41209);
or U41276 (N_41276,N_41122,N_41245);
and U41277 (N_41277,N_41052,N_41043);
or U41278 (N_41278,N_41045,N_41186);
nor U41279 (N_41279,N_41038,N_41222);
xnor U41280 (N_41280,N_41032,N_41096);
nand U41281 (N_41281,N_41172,N_41135);
or U41282 (N_41282,N_41133,N_41204);
or U41283 (N_41283,N_41000,N_41028);
xnor U41284 (N_41284,N_41049,N_41176);
nand U41285 (N_41285,N_41189,N_41180);
xor U41286 (N_41286,N_41058,N_41152);
and U41287 (N_41287,N_41046,N_41218);
or U41288 (N_41288,N_41055,N_41221);
and U41289 (N_41289,N_41181,N_41115);
nand U41290 (N_41290,N_41086,N_41111);
and U41291 (N_41291,N_41183,N_41202);
and U41292 (N_41292,N_41211,N_41170);
xor U41293 (N_41293,N_41236,N_41161);
xnor U41294 (N_41294,N_41178,N_41031);
nor U41295 (N_41295,N_41121,N_41192);
or U41296 (N_41296,N_41080,N_41090);
or U41297 (N_41297,N_41131,N_41116);
and U41298 (N_41298,N_41113,N_41015);
nand U41299 (N_41299,N_41095,N_41127);
xnor U41300 (N_41300,N_41084,N_41009);
xnor U41301 (N_41301,N_41160,N_41134);
and U41302 (N_41302,N_41132,N_41011);
xnor U41303 (N_41303,N_41034,N_41026);
nand U41304 (N_41304,N_41234,N_41085);
nor U41305 (N_41305,N_41016,N_41100);
nor U41306 (N_41306,N_41230,N_41056);
or U41307 (N_41307,N_41003,N_41193);
nor U41308 (N_41308,N_41179,N_41059);
nand U41309 (N_41309,N_41146,N_41089);
and U41310 (N_41310,N_41144,N_41190);
and U41311 (N_41311,N_41167,N_41092);
and U41312 (N_41312,N_41169,N_41074);
xnor U41313 (N_41313,N_41164,N_41037);
xnor U41314 (N_41314,N_41228,N_41063);
nand U41315 (N_41315,N_41174,N_41030);
xnor U41316 (N_41316,N_41112,N_41019);
xnor U41317 (N_41317,N_41149,N_41136);
or U41318 (N_41318,N_41071,N_41173);
nor U41319 (N_41319,N_41035,N_41163);
xor U41320 (N_41320,N_41217,N_41076);
or U41321 (N_41321,N_41175,N_41130);
and U41322 (N_41322,N_41249,N_41097);
nand U41323 (N_41323,N_41103,N_41142);
nor U41324 (N_41324,N_41094,N_41119);
nor U41325 (N_41325,N_41040,N_41194);
nand U41326 (N_41326,N_41246,N_41226);
or U41327 (N_41327,N_41123,N_41126);
nand U41328 (N_41328,N_41117,N_41148);
xor U41329 (N_41329,N_41017,N_41137);
nor U41330 (N_41330,N_41224,N_41070);
and U41331 (N_41331,N_41022,N_41072);
nand U41332 (N_41332,N_41036,N_41061);
xnor U41333 (N_41333,N_41162,N_41184);
and U41334 (N_41334,N_41157,N_41069);
and U41335 (N_41335,N_41001,N_41185);
nor U41336 (N_41336,N_41064,N_41048);
and U41337 (N_41337,N_41215,N_41151);
or U41338 (N_41338,N_41010,N_41232);
and U41339 (N_41339,N_41206,N_41240);
nor U41340 (N_41340,N_41233,N_41177);
or U41341 (N_41341,N_41165,N_41143);
xor U41342 (N_41342,N_41187,N_41093);
or U41343 (N_41343,N_41200,N_41066);
nor U41344 (N_41344,N_41013,N_41008);
and U41345 (N_41345,N_41166,N_41068);
nor U41346 (N_41346,N_41242,N_41198);
or U41347 (N_41347,N_41025,N_41044);
xnor U41348 (N_41348,N_41105,N_41235);
xor U41349 (N_41349,N_41098,N_41196);
and U41350 (N_41350,N_41106,N_41138);
nand U41351 (N_41351,N_41075,N_41104);
nor U41352 (N_41352,N_41205,N_41129);
and U41353 (N_41353,N_41219,N_41191);
or U41354 (N_41354,N_41220,N_41239);
or U41355 (N_41355,N_41054,N_41109);
xnor U41356 (N_41356,N_41244,N_41139);
nor U41357 (N_41357,N_41060,N_41210);
or U41358 (N_41358,N_41077,N_41102);
nand U41359 (N_41359,N_41227,N_41083);
nor U41360 (N_41360,N_41237,N_41231);
or U41361 (N_41361,N_41014,N_41033);
nand U41362 (N_41362,N_41140,N_41050);
nand U41363 (N_41363,N_41225,N_41153);
nor U41364 (N_41364,N_41110,N_41141);
xor U41365 (N_41365,N_41108,N_41101);
or U41366 (N_41366,N_41087,N_41195);
and U41367 (N_41367,N_41243,N_41020);
nor U41368 (N_41368,N_41241,N_41223);
nor U41369 (N_41369,N_41155,N_41062);
or U41370 (N_41370,N_41248,N_41047);
or U41371 (N_41371,N_41088,N_41212);
xnor U41372 (N_41372,N_41002,N_41012);
nor U41373 (N_41373,N_41128,N_41007);
xor U41374 (N_41374,N_41082,N_41124);
and U41375 (N_41375,N_41081,N_41158);
or U41376 (N_41376,N_41091,N_41174);
xnor U41377 (N_41377,N_41205,N_41149);
xnor U41378 (N_41378,N_41116,N_41187);
nand U41379 (N_41379,N_41199,N_41101);
nand U41380 (N_41380,N_41044,N_41221);
xnor U41381 (N_41381,N_41144,N_41246);
and U41382 (N_41382,N_41193,N_41184);
and U41383 (N_41383,N_41151,N_41023);
and U41384 (N_41384,N_41039,N_41181);
nand U41385 (N_41385,N_41038,N_41105);
xnor U41386 (N_41386,N_41055,N_41009);
xor U41387 (N_41387,N_41163,N_41126);
nor U41388 (N_41388,N_41123,N_41016);
or U41389 (N_41389,N_41157,N_41097);
nand U41390 (N_41390,N_41208,N_41038);
or U41391 (N_41391,N_41066,N_41164);
xnor U41392 (N_41392,N_41014,N_41109);
or U41393 (N_41393,N_41185,N_41226);
or U41394 (N_41394,N_41027,N_41083);
or U41395 (N_41395,N_41079,N_41099);
xnor U41396 (N_41396,N_41000,N_41211);
and U41397 (N_41397,N_41108,N_41168);
and U41398 (N_41398,N_41225,N_41147);
nor U41399 (N_41399,N_41055,N_41046);
or U41400 (N_41400,N_41045,N_41096);
or U41401 (N_41401,N_41032,N_41047);
nand U41402 (N_41402,N_41108,N_41203);
xor U41403 (N_41403,N_41161,N_41061);
and U41404 (N_41404,N_41079,N_41155);
and U41405 (N_41405,N_41235,N_41213);
nand U41406 (N_41406,N_41158,N_41179);
nor U41407 (N_41407,N_41087,N_41069);
nor U41408 (N_41408,N_41198,N_41095);
and U41409 (N_41409,N_41128,N_41064);
and U41410 (N_41410,N_41229,N_41225);
and U41411 (N_41411,N_41147,N_41136);
or U41412 (N_41412,N_41179,N_41116);
nand U41413 (N_41413,N_41127,N_41177);
nor U41414 (N_41414,N_41086,N_41113);
xnor U41415 (N_41415,N_41050,N_41183);
or U41416 (N_41416,N_41135,N_41024);
nor U41417 (N_41417,N_41208,N_41151);
and U41418 (N_41418,N_41082,N_41119);
nor U41419 (N_41419,N_41198,N_41234);
or U41420 (N_41420,N_41087,N_41212);
and U41421 (N_41421,N_41237,N_41062);
or U41422 (N_41422,N_41190,N_41151);
and U41423 (N_41423,N_41207,N_41063);
or U41424 (N_41424,N_41203,N_41208);
nor U41425 (N_41425,N_41188,N_41084);
or U41426 (N_41426,N_41025,N_41245);
xor U41427 (N_41427,N_41248,N_41230);
and U41428 (N_41428,N_41226,N_41245);
nand U41429 (N_41429,N_41207,N_41144);
nor U41430 (N_41430,N_41205,N_41138);
nor U41431 (N_41431,N_41201,N_41209);
or U41432 (N_41432,N_41001,N_41122);
nor U41433 (N_41433,N_41120,N_41244);
xnor U41434 (N_41434,N_41167,N_41234);
and U41435 (N_41435,N_41112,N_41078);
nor U41436 (N_41436,N_41176,N_41249);
xor U41437 (N_41437,N_41063,N_41041);
and U41438 (N_41438,N_41123,N_41098);
or U41439 (N_41439,N_41198,N_41053);
or U41440 (N_41440,N_41080,N_41122);
nor U41441 (N_41441,N_41192,N_41156);
nand U41442 (N_41442,N_41240,N_41234);
xor U41443 (N_41443,N_41069,N_41150);
nand U41444 (N_41444,N_41021,N_41019);
nor U41445 (N_41445,N_41084,N_41230);
and U41446 (N_41446,N_41249,N_41216);
nor U41447 (N_41447,N_41123,N_41248);
or U41448 (N_41448,N_41227,N_41166);
nand U41449 (N_41449,N_41118,N_41193);
nand U41450 (N_41450,N_41228,N_41210);
nor U41451 (N_41451,N_41230,N_41101);
and U41452 (N_41452,N_41248,N_41133);
nor U41453 (N_41453,N_41169,N_41192);
or U41454 (N_41454,N_41207,N_41225);
xnor U41455 (N_41455,N_41049,N_41071);
xor U41456 (N_41456,N_41145,N_41050);
xor U41457 (N_41457,N_41061,N_41108);
nand U41458 (N_41458,N_41011,N_41237);
or U41459 (N_41459,N_41056,N_41193);
and U41460 (N_41460,N_41079,N_41002);
or U41461 (N_41461,N_41096,N_41172);
nand U41462 (N_41462,N_41025,N_41083);
nor U41463 (N_41463,N_41214,N_41007);
nor U41464 (N_41464,N_41207,N_41192);
xor U41465 (N_41465,N_41212,N_41217);
or U41466 (N_41466,N_41191,N_41111);
nand U41467 (N_41467,N_41097,N_41225);
and U41468 (N_41468,N_41056,N_41130);
nor U41469 (N_41469,N_41115,N_41136);
xnor U41470 (N_41470,N_41117,N_41152);
or U41471 (N_41471,N_41016,N_41107);
nand U41472 (N_41472,N_41233,N_41237);
xor U41473 (N_41473,N_41109,N_41011);
or U41474 (N_41474,N_41174,N_41111);
and U41475 (N_41475,N_41030,N_41112);
nor U41476 (N_41476,N_41128,N_41240);
xnor U41477 (N_41477,N_41063,N_41001);
nand U41478 (N_41478,N_41214,N_41146);
and U41479 (N_41479,N_41142,N_41125);
and U41480 (N_41480,N_41047,N_41050);
xor U41481 (N_41481,N_41143,N_41243);
nand U41482 (N_41482,N_41031,N_41106);
and U41483 (N_41483,N_41149,N_41001);
xnor U41484 (N_41484,N_41209,N_41191);
and U41485 (N_41485,N_41161,N_41007);
nand U41486 (N_41486,N_41108,N_41025);
and U41487 (N_41487,N_41128,N_41206);
or U41488 (N_41488,N_41144,N_41028);
or U41489 (N_41489,N_41025,N_41190);
or U41490 (N_41490,N_41092,N_41062);
and U41491 (N_41491,N_41239,N_41177);
xnor U41492 (N_41492,N_41143,N_41063);
nor U41493 (N_41493,N_41173,N_41127);
nor U41494 (N_41494,N_41064,N_41037);
nor U41495 (N_41495,N_41005,N_41246);
xor U41496 (N_41496,N_41102,N_41194);
nor U41497 (N_41497,N_41047,N_41242);
and U41498 (N_41498,N_41018,N_41128);
nor U41499 (N_41499,N_41233,N_41106);
xor U41500 (N_41500,N_41456,N_41362);
or U41501 (N_41501,N_41288,N_41336);
or U41502 (N_41502,N_41319,N_41269);
nand U41503 (N_41503,N_41344,N_41333);
or U41504 (N_41504,N_41354,N_41423);
or U41505 (N_41505,N_41260,N_41364);
nor U41506 (N_41506,N_41496,N_41353);
nor U41507 (N_41507,N_41339,N_41419);
nand U41508 (N_41508,N_41273,N_41360);
xor U41509 (N_41509,N_41426,N_41386);
or U41510 (N_41510,N_41286,N_41349);
nand U41511 (N_41511,N_41313,N_41402);
or U41512 (N_41512,N_41284,N_41359);
xnor U41513 (N_41513,N_41250,N_41293);
nand U41514 (N_41514,N_41425,N_41299);
nand U41515 (N_41515,N_41338,N_41468);
and U41516 (N_41516,N_41469,N_41395);
xor U41517 (N_41517,N_41461,N_41436);
nand U41518 (N_41518,N_41438,N_41381);
or U41519 (N_41519,N_41429,N_41376);
nor U41520 (N_41520,N_41358,N_41356);
and U41521 (N_41521,N_41397,N_41321);
and U41522 (N_41522,N_41311,N_41498);
and U41523 (N_41523,N_41332,N_41322);
xnor U41524 (N_41524,N_41261,N_41365);
xor U41525 (N_41525,N_41279,N_41309);
nand U41526 (N_41526,N_41453,N_41324);
and U41527 (N_41527,N_41383,N_41331);
nor U41528 (N_41528,N_41280,N_41351);
or U41529 (N_41529,N_41435,N_41482);
nand U41530 (N_41530,N_41282,N_41492);
and U41531 (N_41531,N_41442,N_41297);
or U41532 (N_41532,N_41465,N_41346);
nor U41533 (N_41533,N_41263,N_41471);
and U41534 (N_41534,N_41254,N_41272);
xor U41535 (N_41535,N_41384,N_41320);
or U41536 (N_41536,N_41427,N_41252);
nor U41537 (N_41537,N_41390,N_41345);
xnor U41538 (N_41538,N_41387,N_41296);
and U41539 (N_41539,N_41460,N_41437);
and U41540 (N_41540,N_41315,N_41458);
or U41541 (N_41541,N_41366,N_41416);
xnor U41542 (N_41542,N_41418,N_41411);
and U41543 (N_41543,N_41481,N_41317);
and U41544 (N_41544,N_41497,N_41447);
nor U41545 (N_41545,N_41323,N_41457);
or U41546 (N_41546,N_41396,N_41255);
or U41547 (N_41547,N_41372,N_41477);
and U41548 (N_41548,N_41414,N_41413);
nor U41549 (N_41549,N_41377,N_41434);
xnor U41550 (N_41550,N_41277,N_41350);
nor U41551 (N_41551,N_41478,N_41483);
nand U41552 (N_41552,N_41473,N_41415);
nor U41553 (N_41553,N_41334,N_41303);
xor U41554 (N_41554,N_41287,N_41424);
nand U41555 (N_41555,N_41256,N_41337);
and U41556 (N_41556,N_41389,N_41432);
nand U41557 (N_41557,N_41441,N_41258);
nand U41558 (N_41558,N_41369,N_41433);
and U41559 (N_41559,N_41392,N_41420);
nor U41560 (N_41560,N_41289,N_41479);
nor U41561 (N_41561,N_41499,N_41398);
and U41562 (N_41562,N_41271,N_41304);
nor U41563 (N_41563,N_41448,N_41253);
or U41564 (N_41564,N_41300,N_41444);
and U41565 (N_41565,N_41443,N_41307);
nor U41566 (N_41566,N_41391,N_41276);
nand U41567 (N_41567,N_41343,N_41452);
or U41568 (N_41568,N_41295,N_41417);
nor U41569 (N_41569,N_41476,N_41480);
and U41570 (N_41570,N_41302,N_41363);
nor U41571 (N_41571,N_41290,N_41318);
or U41572 (N_41572,N_41445,N_41262);
or U41573 (N_41573,N_41488,N_41410);
xnor U41574 (N_41574,N_41373,N_41306);
nor U41575 (N_41575,N_41401,N_41474);
nand U41576 (N_41576,N_41409,N_41379);
nor U41577 (N_41577,N_41327,N_41405);
and U41578 (N_41578,N_41259,N_41371);
nor U41579 (N_41579,N_41305,N_41407);
nor U41580 (N_41580,N_41325,N_41341);
nor U41581 (N_41581,N_41294,N_41470);
xnor U41582 (N_41582,N_41285,N_41385);
nand U41583 (N_41583,N_41340,N_41264);
nand U41584 (N_41584,N_41430,N_41489);
or U41585 (N_41585,N_41493,N_41451);
nand U41586 (N_41586,N_41399,N_41495);
xor U41587 (N_41587,N_41265,N_41472);
nor U41588 (N_41588,N_41310,N_41278);
and U41589 (N_41589,N_41459,N_41494);
xor U41590 (N_41590,N_41403,N_41404);
or U41591 (N_41591,N_41291,N_41274);
or U41592 (N_41592,N_41335,N_41467);
xor U41593 (N_41593,N_41475,N_41266);
xnor U41594 (N_41594,N_41388,N_41355);
and U41595 (N_41595,N_41281,N_41370);
or U41596 (N_41596,N_41454,N_41400);
nor U41597 (N_41597,N_41440,N_41257);
nor U41598 (N_41598,N_41342,N_41330);
nand U41599 (N_41599,N_41394,N_41375);
nor U41600 (N_41600,N_41347,N_41368);
nand U41601 (N_41601,N_41357,N_41464);
or U41602 (N_41602,N_41301,N_41270);
or U41603 (N_41603,N_41484,N_41268);
or U41604 (N_41604,N_41283,N_41406);
or U41605 (N_41605,N_41462,N_41267);
and U41606 (N_41606,N_41491,N_41422);
nor U41607 (N_41607,N_41361,N_41367);
nand U41608 (N_41608,N_41393,N_41329);
or U41609 (N_41609,N_41275,N_41374);
and U41610 (N_41610,N_41490,N_41312);
nand U41611 (N_41611,N_41378,N_41292);
and U41612 (N_41612,N_41298,N_41463);
xor U41613 (N_41613,N_41431,N_41408);
xnor U41614 (N_41614,N_41412,N_41326);
or U41615 (N_41615,N_41308,N_41485);
or U41616 (N_41616,N_41316,N_41314);
nand U41617 (N_41617,N_41486,N_41466);
and U41618 (N_41618,N_41449,N_41352);
or U41619 (N_41619,N_41251,N_41380);
nand U41620 (N_41620,N_41382,N_41328);
xnor U41621 (N_41621,N_41421,N_41487);
or U41622 (N_41622,N_41446,N_41455);
and U41623 (N_41623,N_41428,N_41348);
or U41624 (N_41624,N_41439,N_41450);
or U41625 (N_41625,N_41265,N_41356);
nand U41626 (N_41626,N_41332,N_41359);
and U41627 (N_41627,N_41295,N_41479);
nor U41628 (N_41628,N_41329,N_41442);
xor U41629 (N_41629,N_41359,N_41313);
nor U41630 (N_41630,N_41317,N_41457);
and U41631 (N_41631,N_41267,N_41319);
xor U41632 (N_41632,N_41434,N_41288);
and U41633 (N_41633,N_41391,N_41368);
xor U41634 (N_41634,N_41299,N_41314);
nor U41635 (N_41635,N_41428,N_41305);
nor U41636 (N_41636,N_41346,N_41466);
or U41637 (N_41637,N_41288,N_41369);
nor U41638 (N_41638,N_41332,N_41310);
or U41639 (N_41639,N_41497,N_41382);
nor U41640 (N_41640,N_41319,N_41446);
xnor U41641 (N_41641,N_41472,N_41281);
or U41642 (N_41642,N_41475,N_41473);
and U41643 (N_41643,N_41463,N_41479);
xor U41644 (N_41644,N_41475,N_41466);
nand U41645 (N_41645,N_41277,N_41377);
xor U41646 (N_41646,N_41271,N_41408);
xor U41647 (N_41647,N_41392,N_41385);
or U41648 (N_41648,N_41347,N_41278);
or U41649 (N_41649,N_41411,N_41389);
nor U41650 (N_41650,N_41314,N_41326);
xnor U41651 (N_41651,N_41252,N_41481);
and U41652 (N_41652,N_41409,N_41420);
nand U41653 (N_41653,N_41493,N_41494);
or U41654 (N_41654,N_41431,N_41421);
and U41655 (N_41655,N_41301,N_41372);
xnor U41656 (N_41656,N_41258,N_41263);
and U41657 (N_41657,N_41393,N_41415);
xnor U41658 (N_41658,N_41424,N_41392);
or U41659 (N_41659,N_41460,N_41289);
xor U41660 (N_41660,N_41384,N_41427);
nand U41661 (N_41661,N_41412,N_41433);
xnor U41662 (N_41662,N_41315,N_41365);
and U41663 (N_41663,N_41499,N_41324);
and U41664 (N_41664,N_41465,N_41378);
nor U41665 (N_41665,N_41252,N_41452);
nand U41666 (N_41666,N_41397,N_41461);
or U41667 (N_41667,N_41336,N_41332);
nand U41668 (N_41668,N_41266,N_41328);
and U41669 (N_41669,N_41451,N_41465);
nand U41670 (N_41670,N_41451,N_41488);
and U41671 (N_41671,N_41499,N_41492);
or U41672 (N_41672,N_41412,N_41262);
or U41673 (N_41673,N_41445,N_41282);
or U41674 (N_41674,N_41395,N_41267);
xnor U41675 (N_41675,N_41497,N_41342);
xor U41676 (N_41676,N_41362,N_41404);
or U41677 (N_41677,N_41361,N_41307);
and U41678 (N_41678,N_41254,N_41425);
nand U41679 (N_41679,N_41268,N_41409);
or U41680 (N_41680,N_41303,N_41293);
nand U41681 (N_41681,N_41274,N_41393);
xor U41682 (N_41682,N_41348,N_41297);
and U41683 (N_41683,N_41251,N_41317);
or U41684 (N_41684,N_41278,N_41403);
nor U41685 (N_41685,N_41488,N_41441);
or U41686 (N_41686,N_41430,N_41434);
or U41687 (N_41687,N_41428,N_41409);
or U41688 (N_41688,N_41388,N_41255);
nor U41689 (N_41689,N_41414,N_41495);
nand U41690 (N_41690,N_41462,N_41484);
xor U41691 (N_41691,N_41480,N_41427);
and U41692 (N_41692,N_41488,N_41301);
xnor U41693 (N_41693,N_41319,N_41449);
or U41694 (N_41694,N_41325,N_41462);
xor U41695 (N_41695,N_41278,N_41385);
and U41696 (N_41696,N_41490,N_41294);
and U41697 (N_41697,N_41269,N_41474);
nor U41698 (N_41698,N_41256,N_41316);
or U41699 (N_41699,N_41352,N_41345);
or U41700 (N_41700,N_41380,N_41479);
nor U41701 (N_41701,N_41264,N_41466);
or U41702 (N_41702,N_41291,N_41365);
or U41703 (N_41703,N_41414,N_41295);
nor U41704 (N_41704,N_41272,N_41463);
xnor U41705 (N_41705,N_41343,N_41309);
or U41706 (N_41706,N_41282,N_41362);
xnor U41707 (N_41707,N_41363,N_41489);
and U41708 (N_41708,N_41344,N_41432);
xor U41709 (N_41709,N_41402,N_41444);
and U41710 (N_41710,N_41493,N_41256);
nand U41711 (N_41711,N_41424,N_41276);
nand U41712 (N_41712,N_41358,N_41357);
nand U41713 (N_41713,N_41402,N_41410);
and U41714 (N_41714,N_41406,N_41306);
or U41715 (N_41715,N_41251,N_41366);
and U41716 (N_41716,N_41488,N_41393);
nor U41717 (N_41717,N_41273,N_41468);
nand U41718 (N_41718,N_41324,N_41429);
and U41719 (N_41719,N_41286,N_41329);
nand U41720 (N_41720,N_41413,N_41321);
and U41721 (N_41721,N_41408,N_41332);
or U41722 (N_41722,N_41264,N_41414);
xor U41723 (N_41723,N_41431,N_41305);
nand U41724 (N_41724,N_41356,N_41281);
nor U41725 (N_41725,N_41424,N_41367);
xor U41726 (N_41726,N_41401,N_41346);
or U41727 (N_41727,N_41353,N_41284);
nand U41728 (N_41728,N_41448,N_41331);
and U41729 (N_41729,N_41318,N_41405);
nand U41730 (N_41730,N_41379,N_41256);
xor U41731 (N_41731,N_41291,N_41328);
and U41732 (N_41732,N_41273,N_41400);
nand U41733 (N_41733,N_41312,N_41250);
nand U41734 (N_41734,N_41331,N_41336);
or U41735 (N_41735,N_41348,N_41360);
nor U41736 (N_41736,N_41470,N_41358);
and U41737 (N_41737,N_41276,N_41495);
xor U41738 (N_41738,N_41315,N_41327);
or U41739 (N_41739,N_41470,N_41383);
and U41740 (N_41740,N_41261,N_41263);
and U41741 (N_41741,N_41322,N_41440);
nand U41742 (N_41742,N_41439,N_41350);
and U41743 (N_41743,N_41448,N_41428);
or U41744 (N_41744,N_41488,N_41347);
or U41745 (N_41745,N_41407,N_41477);
nand U41746 (N_41746,N_41493,N_41310);
nor U41747 (N_41747,N_41412,N_41398);
or U41748 (N_41748,N_41280,N_41375);
xor U41749 (N_41749,N_41351,N_41345);
nor U41750 (N_41750,N_41504,N_41550);
nor U41751 (N_41751,N_41744,N_41510);
and U41752 (N_41752,N_41544,N_41673);
xor U41753 (N_41753,N_41503,N_41569);
xnor U41754 (N_41754,N_41685,N_41654);
nor U41755 (N_41755,N_41626,N_41649);
and U41756 (N_41756,N_41529,N_41730);
xor U41757 (N_41757,N_41682,N_41525);
xnor U41758 (N_41758,N_41506,N_41552);
xor U41759 (N_41759,N_41665,N_41636);
nor U41760 (N_41760,N_41566,N_41624);
nand U41761 (N_41761,N_41656,N_41708);
nand U41762 (N_41762,N_41746,N_41704);
or U41763 (N_41763,N_41633,N_41526);
nand U41764 (N_41764,N_41729,N_41643);
or U41765 (N_41765,N_41639,N_41748);
nor U41766 (N_41766,N_41533,N_41672);
or U41767 (N_41767,N_41630,N_41507);
or U41768 (N_41768,N_41647,N_41585);
nand U41769 (N_41769,N_41631,N_41515);
or U41770 (N_41770,N_41578,N_41535);
or U41771 (N_41771,N_41701,N_41727);
nand U41772 (N_41772,N_41595,N_41745);
nand U41773 (N_41773,N_41551,N_41628);
or U41774 (N_41774,N_41739,N_41537);
and U41775 (N_41775,N_41646,N_41596);
nand U41776 (N_41776,N_41680,N_41725);
and U41777 (N_41777,N_41553,N_41686);
and U41778 (N_41778,N_41611,N_41565);
nand U41779 (N_41779,N_41681,N_41549);
xnor U41780 (N_41780,N_41653,N_41668);
and U41781 (N_41781,N_41700,N_41502);
xor U41782 (N_41782,N_41530,N_41664);
nand U41783 (N_41783,N_41677,N_41547);
and U41784 (N_41784,N_41568,N_41548);
and U41785 (N_41785,N_41742,N_41574);
or U41786 (N_41786,N_41598,N_41661);
nor U41787 (N_41787,N_41678,N_41606);
nand U41788 (N_41788,N_41500,N_41592);
xnor U41789 (N_41789,N_41726,N_41732);
and U41790 (N_41790,N_41718,N_41733);
or U41791 (N_41791,N_41579,N_41512);
and U41792 (N_41792,N_41545,N_41737);
xor U41793 (N_41793,N_41534,N_41714);
and U41794 (N_41794,N_41676,N_41591);
xor U41795 (N_41795,N_41590,N_41543);
nand U41796 (N_41796,N_41617,N_41683);
and U41797 (N_41797,N_41696,N_41669);
nand U41798 (N_41798,N_41694,N_41555);
nor U41799 (N_41799,N_41671,N_41687);
nor U41800 (N_41800,N_41554,N_41740);
nor U41801 (N_41801,N_41514,N_41542);
nor U41802 (N_41802,N_41717,N_41675);
nand U41803 (N_41803,N_41662,N_41575);
and U41804 (N_41804,N_41721,N_41702);
and U41805 (N_41805,N_41527,N_41616);
xor U41806 (N_41806,N_41508,N_41651);
nand U41807 (N_41807,N_41667,N_41528);
and U41808 (N_41808,N_41621,N_41659);
or U41809 (N_41809,N_41559,N_41524);
or U41810 (N_41810,N_41658,N_41699);
nand U41811 (N_41811,N_41716,N_41541);
and U41812 (N_41812,N_41517,N_41720);
or U41813 (N_41813,N_41622,N_41655);
nor U41814 (N_41814,N_41632,N_41738);
xor U41815 (N_41815,N_41713,N_41724);
and U41816 (N_41816,N_41600,N_41638);
nor U41817 (N_41817,N_41560,N_41712);
nand U41818 (N_41818,N_41580,N_41516);
nand U41819 (N_41819,N_41657,N_41693);
or U41820 (N_41820,N_41610,N_41731);
xor U41821 (N_41821,N_41557,N_41520);
nor U41822 (N_41822,N_41625,N_41599);
nor U41823 (N_41823,N_41623,N_41640);
or U41824 (N_41824,N_41715,N_41609);
or U41825 (N_41825,N_41531,N_41518);
or U41826 (N_41826,N_41695,N_41741);
and U41827 (N_41827,N_41523,N_41743);
and U41828 (N_41828,N_41567,N_41619);
and U41829 (N_41829,N_41586,N_41573);
and U41830 (N_41830,N_41703,N_41674);
or U41831 (N_41831,N_41536,N_41690);
or U41832 (N_41832,N_41735,N_41612);
nand U41833 (N_41833,N_41634,N_41571);
nand U41834 (N_41834,N_41644,N_41540);
and U41835 (N_41835,N_41577,N_41584);
and U41836 (N_41836,N_41581,N_41509);
nand U41837 (N_41837,N_41546,N_41607);
xnor U41838 (N_41838,N_41629,N_41707);
xnor U41839 (N_41839,N_41601,N_41710);
nor U41840 (N_41840,N_41692,N_41719);
nor U41841 (N_41841,N_41522,N_41562);
and U41842 (N_41842,N_41602,N_41635);
xor U41843 (N_41843,N_41637,N_41604);
and U41844 (N_41844,N_41594,N_41615);
or U41845 (N_41845,N_41572,N_41728);
nor U41846 (N_41846,N_41722,N_41582);
nor U41847 (N_41847,N_41561,N_41709);
xnor U41848 (N_41848,N_41642,N_41576);
nor U41849 (N_41849,N_41705,N_41597);
or U41850 (N_41850,N_41605,N_41660);
or U41851 (N_41851,N_41652,N_41641);
or U41852 (N_41852,N_41670,N_41688);
and U41853 (N_41853,N_41645,N_41505);
nand U41854 (N_41854,N_41501,N_41583);
or U41855 (N_41855,N_41539,N_41723);
nor U41856 (N_41856,N_41558,N_41538);
nor U41857 (N_41857,N_41734,N_41618);
or U41858 (N_41858,N_41747,N_41521);
and U41859 (N_41859,N_41614,N_41613);
and U41860 (N_41860,N_41697,N_41511);
xnor U41861 (N_41861,N_41679,N_41706);
and U41862 (N_41862,N_41532,N_41648);
nor U41863 (N_41863,N_41563,N_41620);
nor U41864 (N_41864,N_41564,N_41603);
and U41865 (N_41865,N_41749,N_41666);
nor U41866 (N_41866,N_41556,N_41570);
and U41867 (N_41867,N_41513,N_41608);
or U41868 (N_41868,N_41691,N_41711);
or U41869 (N_41869,N_41587,N_41698);
xor U41870 (N_41870,N_41589,N_41650);
xor U41871 (N_41871,N_41736,N_41689);
nor U41872 (N_41872,N_41663,N_41519);
nand U41873 (N_41873,N_41588,N_41593);
nand U41874 (N_41874,N_41627,N_41684);
nor U41875 (N_41875,N_41703,N_41607);
and U41876 (N_41876,N_41686,N_41671);
or U41877 (N_41877,N_41648,N_41568);
nor U41878 (N_41878,N_41522,N_41587);
xnor U41879 (N_41879,N_41730,N_41553);
xor U41880 (N_41880,N_41604,N_41661);
nand U41881 (N_41881,N_41501,N_41664);
xnor U41882 (N_41882,N_41714,N_41589);
and U41883 (N_41883,N_41660,N_41692);
and U41884 (N_41884,N_41675,N_41500);
nand U41885 (N_41885,N_41618,N_41659);
xor U41886 (N_41886,N_41734,N_41655);
xor U41887 (N_41887,N_41593,N_41525);
nor U41888 (N_41888,N_41516,N_41684);
or U41889 (N_41889,N_41569,N_41586);
nor U41890 (N_41890,N_41575,N_41678);
and U41891 (N_41891,N_41721,N_41741);
or U41892 (N_41892,N_41530,N_41541);
nor U41893 (N_41893,N_41626,N_41693);
xnor U41894 (N_41894,N_41514,N_41738);
nor U41895 (N_41895,N_41569,N_41742);
xor U41896 (N_41896,N_41693,N_41524);
and U41897 (N_41897,N_41575,N_41742);
nor U41898 (N_41898,N_41561,N_41539);
xnor U41899 (N_41899,N_41603,N_41552);
or U41900 (N_41900,N_41528,N_41631);
nand U41901 (N_41901,N_41559,N_41570);
xnor U41902 (N_41902,N_41591,N_41627);
and U41903 (N_41903,N_41566,N_41695);
xor U41904 (N_41904,N_41549,N_41685);
xor U41905 (N_41905,N_41648,N_41617);
and U41906 (N_41906,N_41680,N_41705);
or U41907 (N_41907,N_41732,N_41613);
and U41908 (N_41908,N_41641,N_41685);
nor U41909 (N_41909,N_41645,N_41715);
nor U41910 (N_41910,N_41709,N_41546);
nand U41911 (N_41911,N_41662,N_41663);
nand U41912 (N_41912,N_41737,N_41687);
nand U41913 (N_41913,N_41672,N_41721);
and U41914 (N_41914,N_41563,N_41699);
and U41915 (N_41915,N_41546,N_41664);
or U41916 (N_41916,N_41694,N_41596);
nor U41917 (N_41917,N_41708,N_41610);
nand U41918 (N_41918,N_41643,N_41607);
and U41919 (N_41919,N_41724,N_41690);
and U41920 (N_41920,N_41744,N_41678);
and U41921 (N_41921,N_41564,N_41647);
xor U41922 (N_41922,N_41629,N_41512);
nand U41923 (N_41923,N_41562,N_41551);
nand U41924 (N_41924,N_41609,N_41524);
and U41925 (N_41925,N_41656,N_41507);
or U41926 (N_41926,N_41733,N_41702);
nand U41927 (N_41927,N_41629,N_41598);
xor U41928 (N_41928,N_41572,N_41634);
or U41929 (N_41929,N_41703,N_41550);
nor U41930 (N_41930,N_41621,N_41510);
xnor U41931 (N_41931,N_41557,N_41660);
and U41932 (N_41932,N_41556,N_41727);
nand U41933 (N_41933,N_41655,N_41720);
and U41934 (N_41934,N_41592,N_41632);
xnor U41935 (N_41935,N_41537,N_41713);
nor U41936 (N_41936,N_41727,N_41708);
nand U41937 (N_41937,N_41616,N_41519);
or U41938 (N_41938,N_41668,N_41599);
and U41939 (N_41939,N_41690,N_41571);
nand U41940 (N_41940,N_41566,N_41707);
and U41941 (N_41941,N_41510,N_41636);
nor U41942 (N_41942,N_41539,N_41628);
or U41943 (N_41943,N_41654,N_41671);
xor U41944 (N_41944,N_41715,N_41711);
and U41945 (N_41945,N_41519,N_41593);
nand U41946 (N_41946,N_41633,N_41601);
or U41947 (N_41947,N_41619,N_41527);
and U41948 (N_41948,N_41522,N_41559);
nand U41949 (N_41949,N_41655,N_41510);
xor U41950 (N_41950,N_41733,N_41680);
and U41951 (N_41951,N_41709,N_41603);
or U41952 (N_41952,N_41555,N_41724);
or U41953 (N_41953,N_41651,N_41515);
nand U41954 (N_41954,N_41747,N_41736);
nand U41955 (N_41955,N_41702,N_41555);
and U41956 (N_41956,N_41600,N_41729);
nor U41957 (N_41957,N_41702,N_41617);
or U41958 (N_41958,N_41632,N_41591);
nand U41959 (N_41959,N_41632,N_41715);
xor U41960 (N_41960,N_41667,N_41592);
nand U41961 (N_41961,N_41531,N_41506);
or U41962 (N_41962,N_41681,N_41637);
xor U41963 (N_41963,N_41545,N_41671);
nand U41964 (N_41964,N_41504,N_41532);
nand U41965 (N_41965,N_41725,N_41598);
nor U41966 (N_41966,N_41510,N_41694);
and U41967 (N_41967,N_41607,N_41709);
nand U41968 (N_41968,N_41671,N_41626);
or U41969 (N_41969,N_41535,N_41582);
nor U41970 (N_41970,N_41717,N_41633);
and U41971 (N_41971,N_41671,N_41594);
xor U41972 (N_41972,N_41660,N_41730);
and U41973 (N_41973,N_41504,N_41693);
nor U41974 (N_41974,N_41717,N_41683);
nand U41975 (N_41975,N_41607,N_41684);
xnor U41976 (N_41976,N_41713,N_41587);
and U41977 (N_41977,N_41546,N_41674);
nand U41978 (N_41978,N_41689,N_41540);
and U41979 (N_41979,N_41734,N_41590);
and U41980 (N_41980,N_41736,N_41691);
nand U41981 (N_41981,N_41520,N_41658);
nand U41982 (N_41982,N_41595,N_41556);
nor U41983 (N_41983,N_41656,N_41645);
nor U41984 (N_41984,N_41541,N_41623);
nand U41985 (N_41985,N_41580,N_41744);
xnor U41986 (N_41986,N_41737,N_41706);
nand U41987 (N_41987,N_41671,N_41523);
or U41988 (N_41988,N_41520,N_41534);
and U41989 (N_41989,N_41743,N_41739);
or U41990 (N_41990,N_41569,N_41558);
nand U41991 (N_41991,N_41526,N_41579);
nand U41992 (N_41992,N_41733,N_41600);
and U41993 (N_41993,N_41575,N_41714);
and U41994 (N_41994,N_41735,N_41667);
nand U41995 (N_41995,N_41547,N_41682);
nand U41996 (N_41996,N_41629,N_41670);
nand U41997 (N_41997,N_41702,N_41708);
nor U41998 (N_41998,N_41536,N_41625);
xnor U41999 (N_41999,N_41606,N_41665);
xnor U42000 (N_42000,N_41793,N_41973);
nand U42001 (N_42001,N_41895,N_41751);
or U42002 (N_42002,N_41885,N_41981);
nand U42003 (N_42003,N_41819,N_41823);
nand U42004 (N_42004,N_41852,N_41923);
xor U42005 (N_42005,N_41889,N_41908);
nor U42006 (N_42006,N_41925,N_41864);
xnor U42007 (N_42007,N_41972,N_41865);
nor U42008 (N_42008,N_41843,N_41994);
xor U42009 (N_42009,N_41919,N_41977);
xnor U42010 (N_42010,N_41763,N_41820);
nand U42011 (N_42011,N_41928,N_41935);
nand U42012 (N_42012,N_41980,N_41797);
xor U42013 (N_42013,N_41888,N_41880);
or U42014 (N_42014,N_41943,N_41815);
and U42015 (N_42015,N_41999,N_41831);
and U42016 (N_42016,N_41760,N_41958);
nand U42017 (N_42017,N_41940,N_41936);
and U42018 (N_42018,N_41877,N_41764);
xnor U42019 (N_42019,N_41870,N_41768);
or U42020 (N_42020,N_41765,N_41961);
nand U42021 (N_42021,N_41757,N_41884);
or U42022 (N_42022,N_41761,N_41986);
or U42023 (N_42023,N_41845,N_41868);
nand U42024 (N_42024,N_41812,N_41901);
or U42025 (N_42025,N_41946,N_41783);
or U42026 (N_42026,N_41938,N_41910);
xor U42027 (N_42027,N_41891,N_41902);
nand U42028 (N_42028,N_41835,N_41930);
or U42029 (N_42029,N_41838,N_41966);
or U42030 (N_42030,N_41849,N_41776);
or U42031 (N_42031,N_41773,N_41970);
or U42032 (N_42032,N_41933,N_41967);
nor U42033 (N_42033,N_41953,N_41903);
nor U42034 (N_42034,N_41784,N_41878);
and U42035 (N_42035,N_41990,N_41769);
and U42036 (N_42036,N_41787,N_41813);
or U42037 (N_42037,N_41792,N_41968);
nand U42038 (N_42038,N_41817,N_41912);
nor U42039 (N_42039,N_41844,N_41841);
nand U42040 (N_42040,N_41979,N_41959);
nand U42041 (N_42041,N_41978,N_41882);
nand U42042 (N_42042,N_41834,N_41932);
nand U42043 (N_42043,N_41833,N_41807);
xor U42044 (N_42044,N_41816,N_41927);
and U42045 (N_42045,N_41995,N_41922);
or U42046 (N_42046,N_41975,N_41893);
nand U42047 (N_42047,N_41754,N_41904);
nor U42048 (N_42048,N_41857,N_41971);
and U42049 (N_42049,N_41756,N_41992);
or U42050 (N_42050,N_41906,N_41851);
nand U42051 (N_42051,N_41991,N_41824);
nand U42052 (N_42052,N_41942,N_41795);
or U42053 (N_42053,N_41926,N_41881);
xnor U42054 (N_42054,N_41918,N_41790);
xnor U42055 (N_42055,N_41855,N_41771);
and U42056 (N_42056,N_41766,N_41955);
nand U42057 (N_42057,N_41862,N_41860);
nor U42058 (N_42058,N_41875,N_41772);
nor U42059 (N_42059,N_41755,N_41989);
nand U42060 (N_42060,N_41794,N_41876);
and U42061 (N_42061,N_41883,N_41802);
xnor U42062 (N_42062,N_41915,N_41898);
xor U42063 (N_42063,N_41993,N_41956);
nand U42064 (N_42064,N_41803,N_41778);
xor U42065 (N_42065,N_41900,N_41848);
or U42066 (N_42066,N_41811,N_41842);
nor U42067 (N_42067,N_41879,N_41810);
xor U42068 (N_42068,N_41905,N_41806);
xor U42069 (N_42069,N_41988,N_41775);
xnor U42070 (N_42070,N_41866,N_41872);
xnor U42071 (N_42071,N_41798,N_41832);
or U42072 (N_42072,N_41779,N_41921);
nand U42073 (N_42073,N_41856,N_41924);
xor U42074 (N_42074,N_41853,N_41894);
nand U42075 (N_42075,N_41752,N_41847);
nor U42076 (N_42076,N_41809,N_41916);
nand U42077 (N_42077,N_41801,N_41854);
xor U42078 (N_42078,N_41987,N_41780);
nor U42079 (N_42079,N_41861,N_41774);
or U42080 (N_42080,N_41788,N_41837);
xnor U42081 (N_42081,N_41758,N_41937);
or U42082 (N_42082,N_41871,N_41781);
and U42083 (N_42083,N_41964,N_41873);
and U42084 (N_42084,N_41799,N_41828);
nor U42085 (N_42085,N_41826,N_41914);
nand U42086 (N_42086,N_41983,N_41920);
and U42087 (N_42087,N_41957,N_41846);
xor U42088 (N_42088,N_41796,N_41947);
nor U42089 (N_42089,N_41952,N_41770);
and U42090 (N_42090,N_41939,N_41836);
and U42091 (N_42091,N_41974,N_41897);
xor U42092 (N_42092,N_41911,N_41997);
nand U42093 (N_42093,N_41839,N_41982);
and U42094 (N_42094,N_41886,N_41985);
nor U42095 (N_42095,N_41814,N_41874);
xor U42096 (N_42096,N_41996,N_41791);
nand U42097 (N_42097,N_41777,N_41858);
nor U42098 (N_42098,N_41998,N_41954);
or U42099 (N_42099,N_41825,N_41869);
or U42100 (N_42100,N_41867,N_41762);
xor U42101 (N_42101,N_41913,N_41785);
or U42102 (N_42102,N_41969,N_41840);
nor U42103 (N_42103,N_41805,N_41944);
xnor U42104 (N_42104,N_41850,N_41984);
xnor U42105 (N_42105,N_41759,N_41945);
xor U42106 (N_42106,N_41896,N_41976);
nor U42107 (N_42107,N_41821,N_41822);
or U42108 (N_42108,N_41808,N_41934);
nor U42109 (N_42109,N_41890,N_41818);
nand U42110 (N_42110,N_41949,N_41917);
xor U42111 (N_42111,N_41829,N_41960);
or U42112 (N_42112,N_41800,N_41899);
xnor U42113 (N_42113,N_41782,N_41963);
nand U42114 (N_42114,N_41892,N_41804);
xor U42115 (N_42115,N_41962,N_41786);
nor U42116 (N_42116,N_41789,N_41859);
nand U42117 (N_42117,N_41907,N_41931);
nor U42118 (N_42118,N_41767,N_41909);
nor U42119 (N_42119,N_41830,N_41951);
nor U42120 (N_42120,N_41929,N_41887);
nor U42121 (N_42121,N_41863,N_41965);
or U42122 (N_42122,N_41827,N_41941);
or U42123 (N_42123,N_41753,N_41750);
xnor U42124 (N_42124,N_41948,N_41950);
nand U42125 (N_42125,N_41911,N_41827);
or U42126 (N_42126,N_41784,N_41847);
xnor U42127 (N_42127,N_41894,N_41786);
or U42128 (N_42128,N_41866,N_41813);
or U42129 (N_42129,N_41831,N_41940);
nand U42130 (N_42130,N_41936,N_41860);
xnor U42131 (N_42131,N_41952,N_41816);
or U42132 (N_42132,N_41987,N_41985);
xnor U42133 (N_42133,N_41974,N_41850);
nor U42134 (N_42134,N_41830,N_41805);
xnor U42135 (N_42135,N_41777,N_41837);
nand U42136 (N_42136,N_41918,N_41862);
and U42137 (N_42137,N_41882,N_41855);
nor U42138 (N_42138,N_41976,N_41847);
nand U42139 (N_42139,N_41783,N_41775);
or U42140 (N_42140,N_41900,N_41932);
or U42141 (N_42141,N_41860,N_41887);
or U42142 (N_42142,N_41816,N_41943);
xnor U42143 (N_42143,N_41913,N_41941);
or U42144 (N_42144,N_41964,N_41838);
nand U42145 (N_42145,N_41822,N_41921);
nor U42146 (N_42146,N_41964,N_41764);
nand U42147 (N_42147,N_41914,N_41878);
xor U42148 (N_42148,N_41773,N_41795);
xor U42149 (N_42149,N_41824,N_41907);
xor U42150 (N_42150,N_41938,N_41925);
nor U42151 (N_42151,N_41865,N_41798);
nand U42152 (N_42152,N_41977,N_41891);
xnor U42153 (N_42153,N_41796,N_41750);
xnor U42154 (N_42154,N_41846,N_41928);
or U42155 (N_42155,N_41997,N_41956);
nand U42156 (N_42156,N_41936,N_41759);
and U42157 (N_42157,N_41824,N_41795);
and U42158 (N_42158,N_41775,N_41970);
or U42159 (N_42159,N_41819,N_41752);
xor U42160 (N_42160,N_41825,N_41751);
and U42161 (N_42161,N_41782,N_41996);
and U42162 (N_42162,N_41960,N_41819);
and U42163 (N_42163,N_41773,N_41937);
and U42164 (N_42164,N_41797,N_41785);
or U42165 (N_42165,N_41885,N_41933);
nand U42166 (N_42166,N_41774,N_41800);
nor U42167 (N_42167,N_41990,N_41787);
nor U42168 (N_42168,N_41963,N_41985);
or U42169 (N_42169,N_41917,N_41816);
nand U42170 (N_42170,N_41867,N_41893);
or U42171 (N_42171,N_41819,N_41788);
xor U42172 (N_42172,N_41819,N_41846);
and U42173 (N_42173,N_41896,N_41891);
and U42174 (N_42174,N_41775,N_41776);
xnor U42175 (N_42175,N_41805,N_41775);
xnor U42176 (N_42176,N_41825,N_41951);
xor U42177 (N_42177,N_41972,N_41789);
or U42178 (N_42178,N_41956,N_41919);
nor U42179 (N_42179,N_41797,N_41976);
or U42180 (N_42180,N_41968,N_41812);
nor U42181 (N_42181,N_41987,N_41774);
or U42182 (N_42182,N_41847,N_41992);
nor U42183 (N_42183,N_41908,N_41881);
xor U42184 (N_42184,N_41777,N_41874);
or U42185 (N_42185,N_41769,N_41871);
nor U42186 (N_42186,N_41844,N_41805);
and U42187 (N_42187,N_41969,N_41952);
nor U42188 (N_42188,N_41993,N_41863);
xor U42189 (N_42189,N_41920,N_41824);
nor U42190 (N_42190,N_41953,N_41847);
or U42191 (N_42191,N_41835,N_41924);
or U42192 (N_42192,N_41751,N_41857);
and U42193 (N_42193,N_41920,N_41754);
nor U42194 (N_42194,N_41879,N_41940);
or U42195 (N_42195,N_41922,N_41833);
nand U42196 (N_42196,N_41757,N_41914);
nor U42197 (N_42197,N_41776,N_41819);
and U42198 (N_42198,N_41799,N_41921);
xor U42199 (N_42199,N_41781,N_41758);
xnor U42200 (N_42200,N_41912,N_41852);
nand U42201 (N_42201,N_41963,N_41898);
nor U42202 (N_42202,N_41948,N_41988);
nor U42203 (N_42203,N_41842,N_41765);
xnor U42204 (N_42204,N_41752,N_41803);
or U42205 (N_42205,N_41907,N_41954);
or U42206 (N_42206,N_41890,N_41770);
xnor U42207 (N_42207,N_41781,N_41826);
and U42208 (N_42208,N_41771,N_41947);
nor U42209 (N_42209,N_41876,N_41957);
and U42210 (N_42210,N_41986,N_41793);
nand U42211 (N_42211,N_41845,N_41853);
xor U42212 (N_42212,N_41996,N_41939);
nand U42213 (N_42213,N_41982,N_41949);
xnor U42214 (N_42214,N_41757,N_41841);
nand U42215 (N_42215,N_41965,N_41931);
nand U42216 (N_42216,N_41855,N_41844);
xnor U42217 (N_42217,N_41975,N_41824);
xor U42218 (N_42218,N_41907,N_41830);
xor U42219 (N_42219,N_41792,N_41803);
nand U42220 (N_42220,N_41769,N_41808);
xor U42221 (N_42221,N_41965,N_41774);
xnor U42222 (N_42222,N_41932,N_41759);
xor U42223 (N_42223,N_41751,N_41854);
and U42224 (N_42224,N_41891,N_41957);
xnor U42225 (N_42225,N_41906,N_41954);
xor U42226 (N_42226,N_41933,N_41864);
nor U42227 (N_42227,N_41957,N_41845);
nor U42228 (N_42228,N_41795,N_41836);
nor U42229 (N_42229,N_41999,N_41813);
or U42230 (N_42230,N_41773,N_41999);
nor U42231 (N_42231,N_41858,N_41867);
nor U42232 (N_42232,N_41953,N_41859);
xor U42233 (N_42233,N_41910,N_41872);
nor U42234 (N_42234,N_41839,N_41771);
nor U42235 (N_42235,N_41924,N_41842);
and U42236 (N_42236,N_41919,N_41836);
or U42237 (N_42237,N_41757,N_41938);
or U42238 (N_42238,N_41905,N_41868);
and U42239 (N_42239,N_41901,N_41943);
or U42240 (N_42240,N_41993,N_41757);
or U42241 (N_42241,N_41810,N_41831);
nand U42242 (N_42242,N_41903,N_41998);
and U42243 (N_42243,N_41789,N_41753);
or U42244 (N_42244,N_41854,N_41919);
nor U42245 (N_42245,N_41816,N_41998);
or U42246 (N_42246,N_41922,N_41959);
nor U42247 (N_42247,N_41943,N_41806);
nand U42248 (N_42248,N_41800,N_41912);
xnor U42249 (N_42249,N_41958,N_41785);
or U42250 (N_42250,N_42199,N_42182);
or U42251 (N_42251,N_42055,N_42205);
or U42252 (N_42252,N_42193,N_42085);
xnor U42253 (N_42253,N_42113,N_42101);
nor U42254 (N_42254,N_42249,N_42143);
and U42255 (N_42255,N_42062,N_42059);
xor U42256 (N_42256,N_42134,N_42244);
and U42257 (N_42257,N_42165,N_42149);
or U42258 (N_42258,N_42160,N_42031);
xnor U42259 (N_42259,N_42078,N_42198);
nand U42260 (N_42260,N_42240,N_42129);
xor U42261 (N_42261,N_42222,N_42245);
nand U42262 (N_42262,N_42127,N_42103);
xor U42263 (N_42263,N_42000,N_42157);
or U42264 (N_42264,N_42166,N_42006);
xnor U42265 (N_42265,N_42045,N_42024);
and U42266 (N_42266,N_42186,N_42147);
xor U42267 (N_42267,N_42139,N_42048);
xnor U42268 (N_42268,N_42184,N_42188);
nor U42269 (N_42269,N_42014,N_42227);
or U42270 (N_42270,N_42230,N_42190);
and U42271 (N_42271,N_42096,N_42039);
nand U42272 (N_42272,N_42215,N_42154);
and U42273 (N_42273,N_42047,N_42213);
xor U42274 (N_42274,N_42159,N_42088);
nor U42275 (N_42275,N_42248,N_42191);
nor U42276 (N_42276,N_42017,N_42108);
or U42277 (N_42277,N_42203,N_42064);
or U42278 (N_42278,N_42219,N_42171);
nor U42279 (N_42279,N_42179,N_42034);
and U42280 (N_42280,N_42138,N_42226);
nand U42281 (N_42281,N_42217,N_42172);
nand U42282 (N_42282,N_42100,N_42004);
and U42283 (N_42283,N_42112,N_42210);
xnor U42284 (N_42284,N_42214,N_42162);
nand U42285 (N_42285,N_42207,N_42056);
xnor U42286 (N_42286,N_42043,N_42211);
nand U42287 (N_42287,N_42135,N_42035);
nor U42288 (N_42288,N_42099,N_42177);
or U42289 (N_42289,N_42015,N_42090);
nor U42290 (N_42290,N_42170,N_42019);
or U42291 (N_42291,N_42054,N_42042);
nand U42292 (N_42292,N_42029,N_42003);
nor U42293 (N_42293,N_42241,N_42163);
xor U42294 (N_42294,N_42049,N_42235);
nor U42295 (N_42295,N_42218,N_42225);
nand U42296 (N_42296,N_42052,N_42033);
nand U42297 (N_42297,N_42136,N_42077);
and U42298 (N_42298,N_42137,N_42046);
nor U42299 (N_42299,N_42093,N_42124);
and U42300 (N_42300,N_42246,N_42117);
xnor U42301 (N_42301,N_42122,N_42074);
and U42302 (N_42302,N_42153,N_42018);
nor U42303 (N_42303,N_42067,N_42178);
nor U42304 (N_42304,N_42234,N_42102);
xor U42305 (N_42305,N_42183,N_42009);
nand U42306 (N_42306,N_42168,N_42083);
nand U42307 (N_42307,N_42080,N_42239);
nor U42308 (N_42308,N_42126,N_42152);
nand U42309 (N_42309,N_42229,N_42180);
nor U42310 (N_42310,N_42023,N_42236);
nand U42311 (N_42311,N_42041,N_42176);
and U42312 (N_42312,N_42087,N_42011);
or U42313 (N_42313,N_42120,N_42075);
nor U42314 (N_42314,N_42247,N_42005);
or U42315 (N_42315,N_42189,N_42022);
nor U42316 (N_42316,N_42107,N_42237);
nand U42317 (N_42317,N_42145,N_42084);
nand U42318 (N_42318,N_42012,N_42216);
nor U42319 (N_42319,N_42013,N_42060);
or U42320 (N_42320,N_42231,N_42094);
nor U42321 (N_42321,N_42032,N_42142);
nand U42322 (N_42322,N_42140,N_42144);
xnor U42323 (N_42323,N_42146,N_42202);
and U42324 (N_42324,N_42050,N_42082);
nand U42325 (N_42325,N_42116,N_42155);
nor U42326 (N_42326,N_42095,N_42020);
or U42327 (N_42327,N_42111,N_42133);
and U42328 (N_42328,N_42086,N_42233);
nand U42329 (N_42329,N_42175,N_42030);
and U42330 (N_42330,N_42164,N_42001);
or U42331 (N_42331,N_42070,N_42174);
nor U42332 (N_42332,N_42148,N_42027);
nand U42333 (N_42333,N_42200,N_42156);
nor U42334 (N_42334,N_42118,N_42040);
and U42335 (N_42335,N_42097,N_42053);
xnor U42336 (N_42336,N_42195,N_42092);
nand U42337 (N_42337,N_42232,N_42242);
or U42338 (N_42338,N_42106,N_42010);
nor U42339 (N_42339,N_42091,N_42197);
nand U42340 (N_42340,N_42026,N_42194);
xor U42341 (N_42341,N_42187,N_42063);
nor U42342 (N_42342,N_42221,N_42130);
nor U42343 (N_42343,N_42044,N_42016);
nor U42344 (N_42344,N_42057,N_42228);
and U42345 (N_42345,N_42051,N_42204);
nor U42346 (N_42346,N_42132,N_42028);
or U42347 (N_42347,N_42151,N_42089);
nor U42348 (N_42348,N_42105,N_42220);
xor U42349 (N_42349,N_42150,N_42038);
nor U42350 (N_42350,N_42131,N_42181);
xnor U42351 (N_42351,N_42098,N_42058);
nor U42352 (N_42352,N_42068,N_42167);
nand U42353 (N_42353,N_42073,N_42071);
or U42354 (N_42354,N_42079,N_42238);
nor U42355 (N_42355,N_42119,N_42185);
nand U42356 (N_42356,N_42223,N_42201);
or U42357 (N_42357,N_42072,N_42169);
xor U42358 (N_42358,N_42109,N_42173);
and U42359 (N_42359,N_42224,N_42212);
nand U42360 (N_42360,N_42123,N_42141);
xor U42361 (N_42361,N_42206,N_42104);
or U42362 (N_42362,N_42025,N_42209);
nor U42363 (N_42363,N_42121,N_42125);
xnor U42364 (N_42364,N_42128,N_42002);
and U42365 (N_42365,N_42161,N_42037);
and U42366 (N_42366,N_42208,N_42069);
xnor U42367 (N_42367,N_42192,N_42114);
and U42368 (N_42368,N_42036,N_42158);
xnor U42369 (N_42369,N_42066,N_42061);
nor U42370 (N_42370,N_42110,N_42076);
nor U42371 (N_42371,N_42007,N_42008);
and U42372 (N_42372,N_42021,N_42081);
nand U42373 (N_42373,N_42115,N_42065);
xor U42374 (N_42374,N_42196,N_42243);
and U42375 (N_42375,N_42136,N_42003);
and U42376 (N_42376,N_42222,N_42177);
and U42377 (N_42377,N_42070,N_42001);
and U42378 (N_42378,N_42024,N_42180);
nand U42379 (N_42379,N_42064,N_42037);
xor U42380 (N_42380,N_42050,N_42101);
and U42381 (N_42381,N_42229,N_42233);
nor U42382 (N_42382,N_42148,N_42209);
nor U42383 (N_42383,N_42156,N_42076);
or U42384 (N_42384,N_42153,N_42220);
xor U42385 (N_42385,N_42241,N_42091);
nor U42386 (N_42386,N_42095,N_42183);
or U42387 (N_42387,N_42087,N_42107);
nand U42388 (N_42388,N_42088,N_42038);
or U42389 (N_42389,N_42106,N_42226);
and U42390 (N_42390,N_42205,N_42085);
xnor U42391 (N_42391,N_42180,N_42123);
nor U42392 (N_42392,N_42009,N_42004);
xnor U42393 (N_42393,N_42096,N_42019);
and U42394 (N_42394,N_42189,N_42249);
or U42395 (N_42395,N_42097,N_42246);
nor U42396 (N_42396,N_42200,N_42234);
nand U42397 (N_42397,N_42028,N_42009);
and U42398 (N_42398,N_42054,N_42210);
and U42399 (N_42399,N_42205,N_42065);
nand U42400 (N_42400,N_42069,N_42031);
nor U42401 (N_42401,N_42063,N_42218);
xor U42402 (N_42402,N_42022,N_42150);
and U42403 (N_42403,N_42128,N_42018);
xnor U42404 (N_42404,N_42188,N_42152);
and U42405 (N_42405,N_42143,N_42111);
nand U42406 (N_42406,N_42222,N_42195);
nor U42407 (N_42407,N_42022,N_42083);
or U42408 (N_42408,N_42131,N_42163);
nor U42409 (N_42409,N_42038,N_42229);
nand U42410 (N_42410,N_42076,N_42022);
nand U42411 (N_42411,N_42078,N_42014);
and U42412 (N_42412,N_42072,N_42170);
and U42413 (N_42413,N_42176,N_42059);
nand U42414 (N_42414,N_42232,N_42224);
nor U42415 (N_42415,N_42157,N_42027);
nor U42416 (N_42416,N_42156,N_42188);
and U42417 (N_42417,N_42048,N_42211);
nand U42418 (N_42418,N_42125,N_42222);
xnor U42419 (N_42419,N_42168,N_42217);
xor U42420 (N_42420,N_42007,N_42096);
nand U42421 (N_42421,N_42070,N_42165);
or U42422 (N_42422,N_42163,N_42217);
or U42423 (N_42423,N_42019,N_42181);
or U42424 (N_42424,N_42016,N_42033);
nor U42425 (N_42425,N_42189,N_42196);
xnor U42426 (N_42426,N_42120,N_42154);
nand U42427 (N_42427,N_42118,N_42184);
nand U42428 (N_42428,N_42142,N_42088);
nand U42429 (N_42429,N_42062,N_42223);
nand U42430 (N_42430,N_42134,N_42054);
or U42431 (N_42431,N_42059,N_42106);
or U42432 (N_42432,N_42230,N_42146);
nand U42433 (N_42433,N_42179,N_42071);
xor U42434 (N_42434,N_42159,N_42176);
nor U42435 (N_42435,N_42163,N_42166);
xor U42436 (N_42436,N_42017,N_42023);
or U42437 (N_42437,N_42173,N_42181);
or U42438 (N_42438,N_42135,N_42238);
or U42439 (N_42439,N_42055,N_42014);
or U42440 (N_42440,N_42051,N_42110);
xnor U42441 (N_42441,N_42058,N_42049);
and U42442 (N_42442,N_42155,N_42112);
or U42443 (N_42443,N_42128,N_42180);
xor U42444 (N_42444,N_42086,N_42104);
and U42445 (N_42445,N_42188,N_42050);
or U42446 (N_42446,N_42178,N_42209);
nand U42447 (N_42447,N_42232,N_42132);
and U42448 (N_42448,N_42194,N_42077);
nor U42449 (N_42449,N_42072,N_42201);
nand U42450 (N_42450,N_42020,N_42057);
nand U42451 (N_42451,N_42117,N_42239);
xnor U42452 (N_42452,N_42054,N_42065);
and U42453 (N_42453,N_42022,N_42182);
nand U42454 (N_42454,N_42013,N_42006);
nand U42455 (N_42455,N_42154,N_42163);
xnor U42456 (N_42456,N_42062,N_42204);
or U42457 (N_42457,N_42183,N_42085);
xor U42458 (N_42458,N_42069,N_42120);
and U42459 (N_42459,N_42074,N_42116);
xor U42460 (N_42460,N_42187,N_42212);
nor U42461 (N_42461,N_42100,N_42170);
xnor U42462 (N_42462,N_42240,N_42179);
nor U42463 (N_42463,N_42102,N_42038);
and U42464 (N_42464,N_42149,N_42163);
or U42465 (N_42465,N_42207,N_42180);
or U42466 (N_42466,N_42056,N_42088);
nand U42467 (N_42467,N_42112,N_42137);
or U42468 (N_42468,N_42124,N_42069);
or U42469 (N_42469,N_42152,N_42091);
and U42470 (N_42470,N_42047,N_42183);
and U42471 (N_42471,N_42128,N_42200);
nor U42472 (N_42472,N_42211,N_42000);
or U42473 (N_42473,N_42181,N_42003);
or U42474 (N_42474,N_42217,N_42192);
xor U42475 (N_42475,N_42242,N_42018);
xnor U42476 (N_42476,N_42197,N_42152);
nand U42477 (N_42477,N_42083,N_42104);
and U42478 (N_42478,N_42187,N_42110);
xnor U42479 (N_42479,N_42035,N_42187);
or U42480 (N_42480,N_42035,N_42240);
nor U42481 (N_42481,N_42121,N_42069);
nand U42482 (N_42482,N_42226,N_42164);
xnor U42483 (N_42483,N_42203,N_42099);
and U42484 (N_42484,N_42078,N_42230);
and U42485 (N_42485,N_42102,N_42168);
xor U42486 (N_42486,N_42184,N_42098);
or U42487 (N_42487,N_42246,N_42087);
nor U42488 (N_42488,N_42184,N_42069);
nand U42489 (N_42489,N_42036,N_42150);
or U42490 (N_42490,N_42024,N_42227);
nor U42491 (N_42491,N_42008,N_42071);
and U42492 (N_42492,N_42174,N_42161);
xor U42493 (N_42493,N_42045,N_42070);
xnor U42494 (N_42494,N_42135,N_42095);
or U42495 (N_42495,N_42008,N_42158);
nor U42496 (N_42496,N_42080,N_42071);
or U42497 (N_42497,N_42146,N_42031);
and U42498 (N_42498,N_42233,N_42083);
nand U42499 (N_42499,N_42025,N_42135);
or U42500 (N_42500,N_42345,N_42434);
and U42501 (N_42501,N_42461,N_42317);
or U42502 (N_42502,N_42385,N_42423);
and U42503 (N_42503,N_42499,N_42495);
xor U42504 (N_42504,N_42453,N_42337);
and U42505 (N_42505,N_42472,N_42302);
or U42506 (N_42506,N_42422,N_42272);
xnor U42507 (N_42507,N_42456,N_42477);
nor U42508 (N_42508,N_42288,N_42384);
xnor U42509 (N_42509,N_42498,N_42439);
and U42510 (N_42510,N_42448,N_42250);
or U42511 (N_42511,N_42271,N_42310);
xnor U42512 (N_42512,N_42287,N_42471);
nor U42513 (N_42513,N_42350,N_42486);
and U42514 (N_42514,N_42364,N_42413);
nand U42515 (N_42515,N_42263,N_42280);
and U42516 (N_42516,N_42268,N_42432);
or U42517 (N_42517,N_42262,N_42397);
nor U42518 (N_42518,N_42341,N_42301);
nand U42519 (N_42519,N_42438,N_42484);
and U42520 (N_42520,N_42464,N_42319);
nor U42521 (N_42521,N_42264,N_42400);
nor U42522 (N_42522,N_42362,N_42418);
and U42523 (N_42523,N_42318,N_42440);
or U42524 (N_42524,N_42433,N_42382);
or U42525 (N_42525,N_42463,N_42386);
and U42526 (N_42526,N_42332,N_42445);
or U42527 (N_42527,N_42387,N_42305);
nand U42528 (N_42528,N_42348,N_42489);
nand U42529 (N_42529,N_42474,N_42366);
nor U42530 (N_42530,N_42333,N_42275);
nand U42531 (N_42531,N_42267,N_42378);
or U42532 (N_42532,N_42443,N_42313);
nor U42533 (N_42533,N_42295,N_42361);
or U42534 (N_42534,N_42425,N_42342);
nor U42535 (N_42535,N_42292,N_42259);
xnor U42536 (N_42536,N_42444,N_42420);
and U42537 (N_42537,N_42395,N_42373);
and U42538 (N_42538,N_42493,N_42253);
or U42539 (N_42539,N_42339,N_42276);
xnor U42540 (N_42540,N_42405,N_42431);
or U42541 (N_42541,N_42468,N_42383);
or U42542 (N_42542,N_42258,N_42465);
and U42543 (N_42543,N_42478,N_42407);
or U42544 (N_42544,N_42283,N_42408);
nor U42545 (N_42545,N_42412,N_42426);
xnor U42546 (N_42546,N_42459,N_42330);
xor U42547 (N_42547,N_42490,N_42307);
nor U42548 (N_42548,N_42488,N_42308);
nand U42549 (N_42549,N_42349,N_42452);
nand U42550 (N_42550,N_42297,N_42331);
xor U42551 (N_42551,N_42446,N_42360);
and U42552 (N_42552,N_42316,N_42251);
and U42553 (N_42553,N_42303,N_42314);
nand U42554 (N_42554,N_42254,N_42340);
or U42555 (N_42555,N_42496,N_42401);
xor U42556 (N_42556,N_42325,N_42327);
xor U42557 (N_42557,N_42458,N_42300);
nor U42558 (N_42558,N_42389,N_42381);
xor U42559 (N_42559,N_42450,N_42380);
or U42560 (N_42560,N_42285,N_42483);
nor U42561 (N_42561,N_42487,N_42375);
or U42562 (N_42562,N_42286,N_42352);
nand U42563 (N_42563,N_42255,N_42353);
xor U42564 (N_42564,N_42334,N_42261);
xor U42565 (N_42565,N_42289,N_42277);
or U42566 (N_42566,N_42479,N_42372);
or U42567 (N_42567,N_42451,N_42343);
nand U42568 (N_42568,N_42299,N_42256);
and U42569 (N_42569,N_42390,N_42291);
nand U42570 (N_42570,N_42398,N_42417);
nor U42571 (N_42571,N_42290,N_42491);
and U42572 (N_42572,N_42306,N_42257);
nor U42573 (N_42573,N_42419,N_42281);
nand U42574 (N_42574,N_42480,N_42335);
nand U42575 (N_42575,N_42475,N_42329);
xnor U42576 (N_42576,N_42324,N_42466);
nand U42577 (N_42577,N_42323,N_42315);
and U42578 (N_42578,N_42406,N_42411);
or U42579 (N_42579,N_42435,N_42494);
nor U42580 (N_42580,N_42436,N_42326);
nand U42581 (N_42581,N_42346,N_42402);
xnor U42582 (N_42582,N_42363,N_42338);
or U42583 (N_42583,N_42428,N_42368);
xor U42584 (N_42584,N_42376,N_42266);
nand U42585 (N_42585,N_42358,N_42322);
nor U42586 (N_42586,N_42476,N_42367);
and U42587 (N_42587,N_42377,N_42447);
nor U42588 (N_42588,N_42365,N_42351);
nor U42589 (N_42589,N_42492,N_42355);
nor U42590 (N_42590,N_42356,N_42274);
nor U42591 (N_42591,N_42293,N_42415);
or U42592 (N_42592,N_42320,N_42457);
xor U42593 (N_42593,N_42311,N_42359);
or U42594 (N_42594,N_42442,N_42462);
or U42595 (N_42595,N_42429,N_42441);
xnor U42596 (N_42596,N_42421,N_42344);
or U42597 (N_42597,N_42270,N_42449);
nand U42598 (N_42598,N_42427,N_42460);
nand U42599 (N_42599,N_42404,N_42485);
nor U42600 (N_42600,N_42357,N_42403);
and U42601 (N_42601,N_42399,N_42328);
xor U42602 (N_42602,N_42455,N_42279);
xor U42603 (N_42603,N_42312,N_42391);
and U42604 (N_42604,N_42396,N_42410);
nand U42605 (N_42605,N_42298,N_42482);
nand U42606 (N_42606,N_42473,N_42265);
nor U42607 (N_42607,N_42336,N_42269);
nand U42608 (N_42608,N_42252,N_42371);
nor U42609 (N_42609,N_42392,N_42278);
and U42610 (N_42610,N_42388,N_42321);
and U42611 (N_42611,N_42354,N_42294);
nand U42612 (N_42612,N_42470,N_42260);
and U42613 (N_42613,N_42347,N_42467);
or U42614 (N_42614,N_42414,N_42393);
nor U42615 (N_42615,N_42454,N_42273);
nor U42616 (N_42616,N_42309,N_42409);
nand U42617 (N_42617,N_42416,N_42379);
nor U42618 (N_42618,N_42394,N_42282);
and U42619 (N_42619,N_42304,N_42424);
xnor U42620 (N_42620,N_42284,N_42369);
or U42621 (N_42621,N_42437,N_42430);
and U42622 (N_42622,N_42374,N_42469);
nor U42623 (N_42623,N_42497,N_42370);
nor U42624 (N_42624,N_42296,N_42481);
nor U42625 (N_42625,N_42373,N_42451);
or U42626 (N_42626,N_42488,N_42349);
nand U42627 (N_42627,N_42399,N_42279);
xnor U42628 (N_42628,N_42316,N_42491);
and U42629 (N_42629,N_42465,N_42445);
and U42630 (N_42630,N_42273,N_42487);
nor U42631 (N_42631,N_42417,N_42425);
nor U42632 (N_42632,N_42487,N_42477);
xnor U42633 (N_42633,N_42332,N_42480);
or U42634 (N_42634,N_42285,N_42386);
xor U42635 (N_42635,N_42470,N_42482);
nor U42636 (N_42636,N_42282,N_42388);
or U42637 (N_42637,N_42405,N_42482);
xnor U42638 (N_42638,N_42411,N_42362);
nand U42639 (N_42639,N_42327,N_42377);
xnor U42640 (N_42640,N_42429,N_42409);
nor U42641 (N_42641,N_42301,N_42305);
and U42642 (N_42642,N_42316,N_42433);
nand U42643 (N_42643,N_42457,N_42396);
nand U42644 (N_42644,N_42351,N_42467);
and U42645 (N_42645,N_42412,N_42303);
xnor U42646 (N_42646,N_42360,N_42392);
or U42647 (N_42647,N_42496,N_42320);
nor U42648 (N_42648,N_42374,N_42479);
and U42649 (N_42649,N_42433,N_42390);
xor U42650 (N_42650,N_42464,N_42317);
xor U42651 (N_42651,N_42387,N_42348);
xnor U42652 (N_42652,N_42348,N_42305);
or U42653 (N_42653,N_42469,N_42319);
xor U42654 (N_42654,N_42291,N_42422);
or U42655 (N_42655,N_42266,N_42308);
and U42656 (N_42656,N_42307,N_42397);
nand U42657 (N_42657,N_42308,N_42372);
nand U42658 (N_42658,N_42432,N_42306);
and U42659 (N_42659,N_42442,N_42362);
or U42660 (N_42660,N_42386,N_42427);
or U42661 (N_42661,N_42483,N_42251);
or U42662 (N_42662,N_42368,N_42410);
or U42663 (N_42663,N_42490,N_42354);
and U42664 (N_42664,N_42425,N_42263);
xor U42665 (N_42665,N_42473,N_42411);
or U42666 (N_42666,N_42334,N_42462);
nand U42667 (N_42667,N_42276,N_42420);
and U42668 (N_42668,N_42451,N_42470);
nor U42669 (N_42669,N_42325,N_42360);
xnor U42670 (N_42670,N_42378,N_42480);
xor U42671 (N_42671,N_42469,N_42459);
nand U42672 (N_42672,N_42477,N_42498);
nand U42673 (N_42673,N_42337,N_42261);
nand U42674 (N_42674,N_42283,N_42356);
nand U42675 (N_42675,N_42353,N_42282);
and U42676 (N_42676,N_42486,N_42442);
and U42677 (N_42677,N_42467,N_42357);
nor U42678 (N_42678,N_42404,N_42469);
xor U42679 (N_42679,N_42486,N_42373);
or U42680 (N_42680,N_42316,N_42373);
nand U42681 (N_42681,N_42419,N_42473);
nand U42682 (N_42682,N_42283,N_42365);
nand U42683 (N_42683,N_42271,N_42438);
nor U42684 (N_42684,N_42493,N_42303);
nand U42685 (N_42685,N_42308,N_42462);
and U42686 (N_42686,N_42366,N_42349);
and U42687 (N_42687,N_42282,N_42484);
xor U42688 (N_42688,N_42402,N_42479);
or U42689 (N_42689,N_42393,N_42278);
nor U42690 (N_42690,N_42320,N_42433);
nand U42691 (N_42691,N_42462,N_42413);
xnor U42692 (N_42692,N_42280,N_42371);
nand U42693 (N_42693,N_42252,N_42341);
or U42694 (N_42694,N_42319,N_42490);
xnor U42695 (N_42695,N_42370,N_42380);
or U42696 (N_42696,N_42269,N_42323);
xnor U42697 (N_42697,N_42364,N_42317);
and U42698 (N_42698,N_42259,N_42397);
and U42699 (N_42699,N_42334,N_42264);
nor U42700 (N_42700,N_42341,N_42337);
and U42701 (N_42701,N_42370,N_42309);
xnor U42702 (N_42702,N_42317,N_42328);
nand U42703 (N_42703,N_42305,N_42400);
xnor U42704 (N_42704,N_42392,N_42481);
nand U42705 (N_42705,N_42447,N_42477);
or U42706 (N_42706,N_42349,N_42319);
nand U42707 (N_42707,N_42431,N_42473);
nand U42708 (N_42708,N_42374,N_42344);
nor U42709 (N_42709,N_42276,N_42351);
and U42710 (N_42710,N_42467,N_42474);
or U42711 (N_42711,N_42457,N_42299);
nand U42712 (N_42712,N_42399,N_42498);
nand U42713 (N_42713,N_42376,N_42482);
or U42714 (N_42714,N_42345,N_42289);
nor U42715 (N_42715,N_42416,N_42432);
xnor U42716 (N_42716,N_42408,N_42332);
or U42717 (N_42717,N_42293,N_42454);
or U42718 (N_42718,N_42415,N_42440);
nor U42719 (N_42719,N_42496,N_42375);
or U42720 (N_42720,N_42496,N_42361);
nor U42721 (N_42721,N_42263,N_42270);
and U42722 (N_42722,N_42477,N_42318);
nand U42723 (N_42723,N_42380,N_42293);
nand U42724 (N_42724,N_42338,N_42322);
xor U42725 (N_42725,N_42258,N_42430);
nand U42726 (N_42726,N_42407,N_42418);
nand U42727 (N_42727,N_42314,N_42438);
nand U42728 (N_42728,N_42466,N_42497);
xnor U42729 (N_42729,N_42333,N_42311);
or U42730 (N_42730,N_42342,N_42312);
or U42731 (N_42731,N_42357,N_42267);
xnor U42732 (N_42732,N_42282,N_42289);
xnor U42733 (N_42733,N_42472,N_42276);
nor U42734 (N_42734,N_42429,N_42283);
or U42735 (N_42735,N_42380,N_42455);
nand U42736 (N_42736,N_42324,N_42283);
nand U42737 (N_42737,N_42412,N_42424);
nand U42738 (N_42738,N_42284,N_42328);
or U42739 (N_42739,N_42496,N_42425);
xnor U42740 (N_42740,N_42411,N_42386);
nand U42741 (N_42741,N_42417,N_42410);
or U42742 (N_42742,N_42461,N_42485);
or U42743 (N_42743,N_42295,N_42351);
xnor U42744 (N_42744,N_42356,N_42302);
and U42745 (N_42745,N_42317,N_42470);
and U42746 (N_42746,N_42458,N_42328);
nand U42747 (N_42747,N_42320,N_42288);
and U42748 (N_42748,N_42253,N_42495);
nand U42749 (N_42749,N_42300,N_42356);
nor U42750 (N_42750,N_42532,N_42735);
nand U42751 (N_42751,N_42627,N_42500);
or U42752 (N_42752,N_42545,N_42587);
and U42753 (N_42753,N_42660,N_42634);
or U42754 (N_42754,N_42667,N_42629);
xor U42755 (N_42755,N_42569,N_42559);
nand U42756 (N_42756,N_42523,N_42624);
and U42757 (N_42757,N_42598,N_42720);
nor U42758 (N_42758,N_42636,N_42704);
nand U42759 (N_42759,N_42588,N_42746);
nand U42760 (N_42760,N_42533,N_42726);
or U42761 (N_42761,N_42561,N_42616);
or U42762 (N_42762,N_42652,N_42540);
nor U42763 (N_42763,N_42713,N_42515);
or U42764 (N_42764,N_42644,N_42661);
and U42765 (N_42765,N_42641,N_42676);
and U42766 (N_42766,N_42510,N_42630);
nand U42767 (N_42767,N_42653,N_42613);
and U42768 (N_42768,N_42712,N_42586);
xnor U42769 (N_42769,N_42589,N_42606);
or U42770 (N_42770,N_42575,N_42709);
nand U42771 (N_42771,N_42679,N_42579);
and U42772 (N_42772,N_42680,N_42734);
nor U42773 (N_42773,N_42529,N_42541);
xor U42774 (N_42774,N_42693,N_42608);
xnor U42775 (N_42775,N_42674,N_42650);
xor U42776 (N_42776,N_42549,N_42711);
nor U42777 (N_42777,N_42505,N_42691);
nor U42778 (N_42778,N_42619,N_42595);
or U42779 (N_42779,N_42651,N_42565);
or U42780 (N_42780,N_42517,N_42550);
nand U42781 (N_42781,N_42640,N_42701);
or U42782 (N_42782,N_42542,N_42527);
and U42783 (N_42783,N_42690,N_42719);
nor U42784 (N_42784,N_42738,N_42714);
nor U42785 (N_42785,N_42553,N_42556);
and U42786 (N_42786,N_42747,N_42605);
or U42787 (N_42787,N_42507,N_42673);
nor U42788 (N_42788,N_42695,N_42737);
xnor U42789 (N_42789,N_42597,N_42551);
or U42790 (N_42790,N_42741,N_42548);
xnor U42791 (N_42791,N_42703,N_42566);
and U42792 (N_42792,N_42546,N_42521);
xor U42793 (N_42793,N_42731,N_42718);
nor U42794 (N_42794,N_42684,N_42508);
nor U42795 (N_42795,N_42562,N_42614);
nor U42796 (N_42796,N_42727,N_42648);
nand U42797 (N_42797,N_42518,N_42740);
or U42798 (N_42798,N_42672,N_42600);
xnor U42799 (N_42799,N_42531,N_42683);
nor U42800 (N_42800,N_42632,N_42604);
nor U42801 (N_42801,N_42519,N_42729);
and U42802 (N_42802,N_42601,N_42697);
xnor U42803 (N_42803,N_42593,N_42513);
and U42804 (N_42804,N_42547,N_42621);
nor U42805 (N_42805,N_42620,N_42723);
or U42806 (N_42806,N_42563,N_42639);
or U42807 (N_42807,N_42524,N_42707);
nand U42808 (N_42808,N_42615,N_42692);
xnor U42809 (N_42809,N_42658,N_42520);
nor U42810 (N_42810,N_42631,N_42696);
xnor U42811 (N_42811,N_42728,N_42682);
nor U42812 (N_42812,N_42539,N_42612);
nor U42813 (N_42813,N_42638,N_42526);
nor U42814 (N_42814,N_42689,N_42739);
nand U42815 (N_42815,N_42623,N_42670);
xnor U42816 (N_42816,N_42509,N_42716);
xor U42817 (N_42817,N_42555,N_42654);
and U42818 (N_42818,N_42617,N_42686);
and U42819 (N_42819,N_42585,N_42592);
or U42820 (N_42820,N_42669,N_42576);
nand U42821 (N_42821,N_42677,N_42665);
xnor U42822 (N_42822,N_42705,N_42688);
or U42823 (N_42823,N_42602,N_42732);
or U42824 (N_42824,N_42618,N_42571);
xor U42825 (N_42825,N_42584,N_42647);
and U42826 (N_42826,N_42649,N_42748);
nor U42827 (N_42827,N_42744,N_42708);
xor U42828 (N_42828,N_42702,N_42512);
and U42829 (N_42829,N_42666,N_42570);
xnor U42830 (N_42830,N_42698,N_42599);
and U42831 (N_42831,N_42504,N_42749);
nor U42832 (N_42832,N_42646,N_42678);
and U42833 (N_42833,N_42645,N_42578);
and U42834 (N_42834,N_42668,N_42730);
nand U42835 (N_42835,N_42567,N_42596);
or U42836 (N_42836,N_42511,N_42560);
nand U42837 (N_42837,N_42554,N_42516);
xor U42838 (N_42838,N_42558,N_42552);
nor U42839 (N_42839,N_42706,N_42610);
nand U42840 (N_42840,N_42543,N_42642);
nor U42841 (N_42841,N_42710,N_42611);
or U42842 (N_42842,N_42503,N_42564);
nand U42843 (N_42843,N_42671,N_42534);
nand U42844 (N_42844,N_42607,N_42528);
nand U42845 (N_42845,N_42685,N_42538);
xnor U42846 (N_42846,N_42525,N_42609);
xnor U42847 (N_42847,N_42501,N_42514);
xor U42848 (N_42848,N_42643,N_42694);
xor U42849 (N_42849,N_42577,N_42681);
xor U42850 (N_42850,N_42568,N_42742);
or U42851 (N_42851,N_42715,N_42721);
nor U42852 (N_42852,N_42743,N_42535);
nor U42853 (N_42853,N_42522,N_42700);
nor U42854 (N_42854,N_42675,N_42574);
or U42855 (N_42855,N_42502,N_42662);
xnor U42856 (N_42856,N_42506,N_42724);
and U42857 (N_42857,N_42733,N_42536);
and U42858 (N_42858,N_42583,N_42687);
nand U42859 (N_42859,N_42580,N_42628);
nor U42860 (N_42860,N_42635,N_42656);
xor U42861 (N_42861,N_42657,N_42622);
nor U42862 (N_42862,N_42582,N_42663);
xnor U42863 (N_42863,N_42725,N_42745);
nand U42864 (N_42864,N_42626,N_42625);
nand U42865 (N_42865,N_42655,N_42544);
nand U42866 (N_42866,N_42699,N_42537);
nand U42867 (N_42867,N_42633,N_42572);
nor U42868 (N_42868,N_42717,N_42659);
xor U42869 (N_42869,N_42581,N_42594);
nand U42870 (N_42870,N_42530,N_42590);
xor U42871 (N_42871,N_42573,N_42557);
nor U42872 (N_42872,N_42637,N_42603);
or U42873 (N_42873,N_42591,N_42664);
xnor U42874 (N_42874,N_42722,N_42736);
and U42875 (N_42875,N_42719,N_42575);
xnor U42876 (N_42876,N_42617,N_42663);
xnor U42877 (N_42877,N_42528,N_42533);
nor U42878 (N_42878,N_42700,N_42699);
and U42879 (N_42879,N_42621,N_42742);
and U42880 (N_42880,N_42565,N_42694);
and U42881 (N_42881,N_42722,N_42634);
and U42882 (N_42882,N_42659,N_42558);
xor U42883 (N_42883,N_42732,N_42648);
nand U42884 (N_42884,N_42607,N_42570);
and U42885 (N_42885,N_42634,N_42544);
or U42886 (N_42886,N_42686,N_42502);
and U42887 (N_42887,N_42656,N_42547);
nand U42888 (N_42888,N_42733,N_42665);
nand U42889 (N_42889,N_42505,N_42707);
and U42890 (N_42890,N_42683,N_42609);
nand U42891 (N_42891,N_42530,N_42601);
xnor U42892 (N_42892,N_42552,N_42645);
xnor U42893 (N_42893,N_42508,N_42698);
nand U42894 (N_42894,N_42628,N_42668);
or U42895 (N_42895,N_42683,N_42693);
or U42896 (N_42896,N_42572,N_42618);
and U42897 (N_42897,N_42522,N_42595);
nor U42898 (N_42898,N_42724,N_42533);
and U42899 (N_42899,N_42542,N_42707);
nand U42900 (N_42900,N_42593,N_42606);
nor U42901 (N_42901,N_42710,N_42649);
nor U42902 (N_42902,N_42586,N_42634);
nor U42903 (N_42903,N_42581,N_42532);
and U42904 (N_42904,N_42531,N_42557);
and U42905 (N_42905,N_42741,N_42642);
xnor U42906 (N_42906,N_42709,N_42549);
xnor U42907 (N_42907,N_42537,N_42738);
nor U42908 (N_42908,N_42703,N_42593);
nand U42909 (N_42909,N_42641,N_42523);
xnor U42910 (N_42910,N_42663,N_42509);
xor U42911 (N_42911,N_42517,N_42536);
nand U42912 (N_42912,N_42566,N_42720);
or U42913 (N_42913,N_42570,N_42746);
and U42914 (N_42914,N_42658,N_42709);
nand U42915 (N_42915,N_42645,N_42617);
and U42916 (N_42916,N_42695,N_42518);
xor U42917 (N_42917,N_42571,N_42512);
or U42918 (N_42918,N_42685,N_42614);
nor U42919 (N_42919,N_42626,N_42737);
nor U42920 (N_42920,N_42536,N_42567);
nor U42921 (N_42921,N_42560,N_42698);
xor U42922 (N_42922,N_42692,N_42632);
nor U42923 (N_42923,N_42565,N_42653);
or U42924 (N_42924,N_42602,N_42705);
or U42925 (N_42925,N_42656,N_42723);
or U42926 (N_42926,N_42704,N_42748);
xnor U42927 (N_42927,N_42582,N_42697);
and U42928 (N_42928,N_42580,N_42640);
nor U42929 (N_42929,N_42592,N_42530);
and U42930 (N_42930,N_42621,N_42654);
and U42931 (N_42931,N_42551,N_42718);
xnor U42932 (N_42932,N_42640,N_42509);
nand U42933 (N_42933,N_42568,N_42578);
xnor U42934 (N_42934,N_42696,N_42665);
or U42935 (N_42935,N_42644,N_42662);
and U42936 (N_42936,N_42705,N_42556);
nand U42937 (N_42937,N_42538,N_42516);
xor U42938 (N_42938,N_42712,N_42695);
nor U42939 (N_42939,N_42671,N_42685);
nand U42940 (N_42940,N_42567,N_42591);
nor U42941 (N_42941,N_42589,N_42500);
nand U42942 (N_42942,N_42603,N_42672);
and U42943 (N_42943,N_42708,N_42581);
nand U42944 (N_42944,N_42519,N_42515);
xor U42945 (N_42945,N_42637,N_42682);
xor U42946 (N_42946,N_42614,N_42648);
nor U42947 (N_42947,N_42578,N_42691);
or U42948 (N_42948,N_42697,N_42600);
or U42949 (N_42949,N_42633,N_42553);
xnor U42950 (N_42950,N_42652,N_42648);
or U42951 (N_42951,N_42585,N_42548);
or U42952 (N_42952,N_42637,N_42549);
nand U42953 (N_42953,N_42716,N_42700);
nand U42954 (N_42954,N_42520,N_42529);
or U42955 (N_42955,N_42618,N_42749);
nor U42956 (N_42956,N_42719,N_42560);
and U42957 (N_42957,N_42710,N_42561);
nand U42958 (N_42958,N_42532,N_42585);
or U42959 (N_42959,N_42674,N_42644);
nor U42960 (N_42960,N_42595,N_42713);
or U42961 (N_42961,N_42534,N_42606);
nor U42962 (N_42962,N_42703,N_42713);
or U42963 (N_42963,N_42590,N_42620);
xnor U42964 (N_42964,N_42518,N_42684);
and U42965 (N_42965,N_42675,N_42578);
nor U42966 (N_42966,N_42612,N_42641);
nand U42967 (N_42967,N_42650,N_42608);
or U42968 (N_42968,N_42741,N_42533);
or U42969 (N_42969,N_42597,N_42504);
nor U42970 (N_42970,N_42559,N_42644);
nor U42971 (N_42971,N_42745,N_42733);
and U42972 (N_42972,N_42502,N_42543);
xnor U42973 (N_42973,N_42666,N_42625);
nor U42974 (N_42974,N_42542,N_42623);
and U42975 (N_42975,N_42610,N_42679);
or U42976 (N_42976,N_42684,N_42742);
and U42977 (N_42977,N_42577,N_42685);
nor U42978 (N_42978,N_42725,N_42587);
or U42979 (N_42979,N_42665,N_42707);
and U42980 (N_42980,N_42596,N_42580);
nor U42981 (N_42981,N_42691,N_42513);
xnor U42982 (N_42982,N_42692,N_42651);
xnor U42983 (N_42983,N_42542,N_42737);
nor U42984 (N_42984,N_42719,N_42559);
nand U42985 (N_42985,N_42527,N_42513);
nand U42986 (N_42986,N_42575,N_42547);
and U42987 (N_42987,N_42595,N_42628);
or U42988 (N_42988,N_42664,N_42740);
nand U42989 (N_42989,N_42655,N_42576);
nor U42990 (N_42990,N_42648,N_42620);
xnor U42991 (N_42991,N_42553,N_42512);
or U42992 (N_42992,N_42543,N_42744);
nand U42993 (N_42993,N_42678,N_42692);
and U42994 (N_42994,N_42651,N_42598);
nor U42995 (N_42995,N_42533,N_42641);
nor U42996 (N_42996,N_42606,N_42613);
nand U42997 (N_42997,N_42733,N_42691);
or U42998 (N_42998,N_42569,N_42630);
xor U42999 (N_42999,N_42585,N_42658);
nor U43000 (N_43000,N_42968,N_42990);
nor U43001 (N_43001,N_42893,N_42870);
and U43002 (N_43002,N_42826,N_42825);
nand U43003 (N_43003,N_42984,N_42814);
and U43004 (N_43004,N_42944,N_42800);
nor U43005 (N_43005,N_42900,N_42985);
nand U43006 (N_43006,N_42788,N_42999);
nand U43007 (N_43007,N_42861,N_42883);
nor U43008 (N_43008,N_42763,N_42879);
and U43009 (N_43009,N_42928,N_42810);
nor U43010 (N_43010,N_42891,N_42764);
nand U43011 (N_43011,N_42817,N_42804);
nor U43012 (N_43012,N_42751,N_42915);
xnor U43013 (N_43013,N_42770,N_42762);
and U43014 (N_43014,N_42924,N_42809);
and U43015 (N_43015,N_42778,N_42941);
and U43016 (N_43016,N_42802,N_42898);
or U43017 (N_43017,N_42859,N_42953);
and U43018 (N_43018,N_42949,N_42828);
and U43019 (N_43019,N_42851,N_42858);
or U43020 (N_43020,N_42995,N_42831);
and U43021 (N_43021,N_42906,N_42962);
xor U43022 (N_43022,N_42926,N_42756);
xnor U43023 (N_43023,N_42881,N_42799);
xor U43024 (N_43024,N_42836,N_42753);
xor U43025 (N_43025,N_42913,N_42946);
nand U43026 (N_43026,N_42773,N_42854);
nor U43027 (N_43027,N_42954,N_42860);
and U43028 (N_43028,N_42922,N_42960);
or U43029 (N_43029,N_42779,N_42867);
nor U43030 (N_43030,N_42925,N_42772);
nand U43031 (N_43031,N_42961,N_42996);
nor U43032 (N_43032,N_42818,N_42793);
or U43033 (N_43033,N_42843,N_42899);
nor U43034 (N_43034,N_42987,N_42821);
nand U43035 (N_43035,N_42761,N_42963);
xnor U43036 (N_43036,N_42872,N_42873);
and U43037 (N_43037,N_42816,N_42903);
and U43038 (N_43038,N_42973,N_42839);
nand U43039 (N_43039,N_42886,N_42937);
nand U43040 (N_43040,N_42787,N_42908);
nor U43041 (N_43041,N_42754,N_42874);
and U43042 (N_43042,N_42940,N_42864);
and U43043 (N_43043,N_42786,N_42827);
nand U43044 (N_43044,N_42783,N_42796);
nor U43045 (N_43045,N_42977,N_42853);
nor U43046 (N_43046,N_42840,N_42884);
nand U43047 (N_43047,N_42855,N_42997);
or U43048 (N_43048,N_42998,N_42808);
and U43049 (N_43049,N_42824,N_42780);
xnor U43050 (N_43050,N_42907,N_42849);
and U43051 (N_43051,N_42807,N_42852);
and U43052 (N_43052,N_42904,N_42757);
and U43053 (N_43053,N_42951,N_42958);
xor U43054 (N_43054,N_42847,N_42834);
or U43055 (N_43055,N_42755,N_42994);
xor U43056 (N_43056,N_42803,N_42919);
nor U43057 (N_43057,N_42797,N_42813);
xnor U43058 (N_43058,N_42896,N_42866);
and U43059 (N_43059,N_42805,N_42939);
or U43060 (N_43060,N_42917,N_42911);
and U43061 (N_43061,N_42776,N_42869);
and U43062 (N_43062,N_42765,N_42811);
and U43063 (N_43063,N_42857,N_42932);
and U43064 (N_43064,N_42856,N_42912);
and U43065 (N_43065,N_42892,N_42947);
nor U43066 (N_43066,N_42875,N_42974);
or U43067 (N_43067,N_42838,N_42914);
or U43068 (N_43068,N_42952,N_42823);
nor U43069 (N_43069,N_42981,N_42822);
xnor U43070 (N_43070,N_42850,N_42792);
or U43071 (N_43071,N_42905,N_42830);
nand U43072 (N_43072,N_42806,N_42833);
nand U43073 (N_43073,N_42901,N_42991);
and U43074 (N_43074,N_42832,N_42931);
and U43075 (N_43075,N_42895,N_42938);
or U43076 (N_43076,N_42978,N_42848);
nor U43077 (N_43077,N_42976,N_42888);
nor U43078 (N_43078,N_42777,N_42885);
nand U43079 (N_43079,N_42846,N_42945);
xnor U43080 (N_43080,N_42970,N_42837);
nand U43081 (N_43081,N_42880,N_42812);
and U43082 (N_43082,N_42815,N_42890);
xnor U43083 (N_43083,N_42784,N_42782);
and U43084 (N_43084,N_42750,N_42868);
nor U43085 (N_43085,N_42966,N_42933);
nor U43086 (N_43086,N_42781,N_42909);
or U43087 (N_43087,N_42835,N_42758);
nand U43088 (N_43088,N_42927,N_42790);
and U43089 (N_43089,N_42844,N_42829);
nand U43090 (N_43090,N_42877,N_42959);
or U43091 (N_43091,N_42986,N_42794);
or U43092 (N_43092,N_42955,N_42916);
and U43093 (N_43093,N_42766,N_42775);
nor U43094 (N_43094,N_42948,N_42935);
nor U43095 (N_43095,N_42863,N_42887);
nor U43096 (N_43096,N_42820,N_42920);
nand U43097 (N_43097,N_42801,N_42982);
nand U43098 (N_43098,N_42956,N_42865);
xor U43099 (N_43099,N_42983,N_42992);
nand U43100 (N_43100,N_42921,N_42930);
or U43101 (N_43101,N_42845,N_42798);
nand U43102 (N_43102,N_42943,N_42934);
nand U43103 (N_43103,N_42871,N_42878);
xor U43104 (N_43104,N_42936,N_42842);
and U43105 (N_43105,N_42980,N_42993);
nand U43106 (N_43106,N_42942,N_42910);
nor U43107 (N_43107,N_42918,N_42972);
or U43108 (N_43108,N_42771,N_42795);
or U43109 (N_43109,N_42768,N_42862);
nand U43110 (N_43110,N_42774,N_42929);
and U43111 (N_43111,N_42897,N_42967);
xor U43112 (N_43112,N_42894,N_42760);
nor U43113 (N_43113,N_42979,N_42950);
or U43114 (N_43114,N_42965,N_42882);
xor U43115 (N_43115,N_42819,N_42989);
nor U43116 (N_43116,N_42923,N_42964);
and U43117 (N_43117,N_42767,N_42785);
or U43118 (N_43118,N_42969,N_42769);
nor U43119 (N_43119,N_42789,N_42752);
or U43120 (N_43120,N_42791,N_42889);
or U43121 (N_43121,N_42759,N_42988);
xor U43122 (N_43122,N_42957,N_42902);
xnor U43123 (N_43123,N_42841,N_42971);
or U43124 (N_43124,N_42876,N_42975);
xnor U43125 (N_43125,N_42945,N_42920);
and U43126 (N_43126,N_42787,N_42910);
or U43127 (N_43127,N_42773,N_42780);
nor U43128 (N_43128,N_42806,N_42791);
nor U43129 (N_43129,N_42775,N_42861);
and U43130 (N_43130,N_42853,N_42840);
nand U43131 (N_43131,N_42969,N_42877);
nor U43132 (N_43132,N_42986,N_42863);
xor U43133 (N_43133,N_42976,N_42844);
or U43134 (N_43134,N_42917,N_42864);
nor U43135 (N_43135,N_42948,N_42823);
nand U43136 (N_43136,N_42872,N_42869);
or U43137 (N_43137,N_42764,N_42876);
and U43138 (N_43138,N_42879,N_42835);
xor U43139 (N_43139,N_42845,N_42751);
xor U43140 (N_43140,N_42975,N_42839);
or U43141 (N_43141,N_42782,N_42860);
nor U43142 (N_43142,N_42935,N_42754);
nand U43143 (N_43143,N_42971,N_42866);
xor U43144 (N_43144,N_42797,N_42927);
nand U43145 (N_43145,N_42976,N_42890);
xnor U43146 (N_43146,N_42926,N_42797);
nand U43147 (N_43147,N_42907,N_42905);
or U43148 (N_43148,N_42849,N_42879);
nand U43149 (N_43149,N_42954,N_42999);
or U43150 (N_43150,N_42877,N_42876);
nand U43151 (N_43151,N_42754,N_42912);
nor U43152 (N_43152,N_42932,N_42820);
nand U43153 (N_43153,N_42988,N_42787);
nor U43154 (N_43154,N_42836,N_42763);
xnor U43155 (N_43155,N_42762,N_42999);
xnor U43156 (N_43156,N_42797,N_42964);
nand U43157 (N_43157,N_42851,N_42857);
nor U43158 (N_43158,N_42873,N_42972);
nand U43159 (N_43159,N_42854,N_42765);
nor U43160 (N_43160,N_42971,N_42905);
or U43161 (N_43161,N_42880,N_42860);
and U43162 (N_43162,N_42791,N_42953);
or U43163 (N_43163,N_42766,N_42774);
nor U43164 (N_43164,N_42857,N_42891);
nor U43165 (N_43165,N_42889,N_42994);
nand U43166 (N_43166,N_42794,N_42811);
or U43167 (N_43167,N_42764,N_42976);
xnor U43168 (N_43168,N_42993,N_42761);
nand U43169 (N_43169,N_42994,N_42775);
nand U43170 (N_43170,N_42927,N_42841);
and U43171 (N_43171,N_42841,N_42953);
or U43172 (N_43172,N_42853,N_42818);
xor U43173 (N_43173,N_42770,N_42854);
or U43174 (N_43174,N_42790,N_42771);
nand U43175 (N_43175,N_42851,N_42754);
and U43176 (N_43176,N_42981,N_42971);
and U43177 (N_43177,N_42957,N_42784);
xnor U43178 (N_43178,N_42894,N_42858);
nand U43179 (N_43179,N_42869,N_42859);
xnor U43180 (N_43180,N_42889,N_42913);
nand U43181 (N_43181,N_42771,N_42864);
or U43182 (N_43182,N_42779,N_42937);
and U43183 (N_43183,N_42757,N_42905);
or U43184 (N_43184,N_42896,N_42891);
nand U43185 (N_43185,N_42910,N_42926);
and U43186 (N_43186,N_42856,N_42832);
or U43187 (N_43187,N_42758,N_42856);
and U43188 (N_43188,N_42931,N_42891);
xor U43189 (N_43189,N_42982,N_42878);
or U43190 (N_43190,N_42888,N_42753);
nor U43191 (N_43191,N_42814,N_42834);
nand U43192 (N_43192,N_42831,N_42888);
and U43193 (N_43193,N_42809,N_42901);
nand U43194 (N_43194,N_42774,N_42965);
nor U43195 (N_43195,N_42914,N_42939);
or U43196 (N_43196,N_42826,N_42970);
and U43197 (N_43197,N_42889,N_42764);
nor U43198 (N_43198,N_42839,N_42936);
nor U43199 (N_43199,N_42932,N_42869);
nor U43200 (N_43200,N_42815,N_42886);
nand U43201 (N_43201,N_42783,N_42888);
and U43202 (N_43202,N_42883,N_42935);
xor U43203 (N_43203,N_42937,N_42917);
nor U43204 (N_43204,N_42856,N_42819);
xnor U43205 (N_43205,N_42830,N_42859);
nand U43206 (N_43206,N_42776,N_42885);
xor U43207 (N_43207,N_42764,N_42859);
xnor U43208 (N_43208,N_42932,N_42771);
nand U43209 (N_43209,N_42776,N_42815);
and U43210 (N_43210,N_42751,N_42855);
nor U43211 (N_43211,N_42923,N_42948);
nor U43212 (N_43212,N_42964,N_42799);
and U43213 (N_43213,N_42785,N_42876);
and U43214 (N_43214,N_42944,N_42839);
nor U43215 (N_43215,N_42829,N_42968);
xnor U43216 (N_43216,N_42842,N_42955);
or U43217 (N_43217,N_42769,N_42944);
nand U43218 (N_43218,N_42853,N_42780);
nand U43219 (N_43219,N_42971,N_42888);
nor U43220 (N_43220,N_42826,N_42965);
and U43221 (N_43221,N_42873,N_42841);
or U43222 (N_43222,N_42868,N_42895);
xnor U43223 (N_43223,N_42929,N_42831);
nor U43224 (N_43224,N_42767,N_42801);
nor U43225 (N_43225,N_42754,N_42989);
nand U43226 (N_43226,N_42910,N_42846);
nor U43227 (N_43227,N_42975,N_42805);
nor U43228 (N_43228,N_42869,N_42965);
xnor U43229 (N_43229,N_42854,N_42786);
nor U43230 (N_43230,N_42980,N_42977);
xor U43231 (N_43231,N_42790,N_42776);
or U43232 (N_43232,N_42844,N_42936);
and U43233 (N_43233,N_42765,N_42882);
nand U43234 (N_43234,N_42763,N_42930);
and U43235 (N_43235,N_42770,N_42824);
or U43236 (N_43236,N_42962,N_42839);
xor U43237 (N_43237,N_42858,N_42782);
and U43238 (N_43238,N_42818,N_42836);
or U43239 (N_43239,N_42870,N_42941);
or U43240 (N_43240,N_42871,N_42956);
xnor U43241 (N_43241,N_42779,N_42944);
nand U43242 (N_43242,N_42993,N_42841);
xor U43243 (N_43243,N_42862,N_42994);
xor U43244 (N_43244,N_42989,N_42930);
or U43245 (N_43245,N_42830,N_42870);
xor U43246 (N_43246,N_42860,N_42871);
xor U43247 (N_43247,N_42837,N_42756);
and U43248 (N_43248,N_42778,N_42760);
nor U43249 (N_43249,N_42787,N_42972);
xor U43250 (N_43250,N_43011,N_43083);
and U43251 (N_43251,N_43107,N_43120);
nor U43252 (N_43252,N_43000,N_43150);
nand U43253 (N_43253,N_43144,N_43181);
and U43254 (N_43254,N_43093,N_43089);
and U43255 (N_43255,N_43080,N_43192);
and U43256 (N_43256,N_43166,N_43173);
xnor U43257 (N_43257,N_43197,N_43194);
xor U43258 (N_43258,N_43189,N_43196);
nor U43259 (N_43259,N_43004,N_43233);
and U43260 (N_43260,N_43147,N_43100);
and U43261 (N_43261,N_43244,N_43112);
nand U43262 (N_43262,N_43175,N_43047);
and U43263 (N_43263,N_43180,N_43161);
nor U43264 (N_43264,N_43246,N_43230);
xor U43265 (N_43265,N_43241,N_43232);
xnor U43266 (N_43266,N_43245,N_43101);
nor U43267 (N_43267,N_43206,N_43212);
and U43268 (N_43268,N_43062,N_43159);
xor U43269 (N_43269,N_43037,N_43091);
nor U43270 (N_43270,N_43121,N_43139);
or U43271 (N_43271,N_43013,N_43220);
and U43272 (N_43272,N_43242,N_43015);
nor U43273 (N_43273,N_43009,N_43012);
nand U43274 (N_43274,N_43050,N_43155);
or U43275 (N_43275,N_43191,N_43014);
nor U43276 (N_43276,N_43209,N_43026);
or U43277 (N_43277,N_43193,N_43207);
or U43278 (N_43278,N_43141,N_43236);
xor U43279 (N_43279,N_43152,N_43127);
xor U43280 (N_43280,N_43137,N_43095);
nand U43281 (N_43281,N_43199,N_43118);
and U43282 (N_43282,N_43184,N_43059);
or U43283 (N_43283,N_43163,N_43016);
nor U43284 (N_43284,N_43198,N_43102);
and U43285 (N_43285,N_43052,N_43222);
nand U43286 (N_43286,N_43087,N_43098);
or U43287 (N_43287,N_43129,N_43188);
or U43288 (N_43288,N_43224,N_43051);
or U43289 (N_43289,N_43125,N_43097);
and U43290 (N_43290,N_43063,N_43092);
nand U43291 (N_43291,N_43170,N_43067);
nor U43292 (N_43292,N_43130,N_43044);
nand U43293 (N_43293,N_43049,N_43056);
xnor U43294 (N_43294,N_43231,N_43070);
or U43295 (N_43295,N_43162,N_43226);
or U43296 (N_43296,N_43034,N_43061);
xor U43297 (N_43297,N_43024,N_43133);
nor U43298 (N_43298,N_43001,N_43234);
nand U43299 (N_43299,N_43073,N_43079);
nor U43300 (N_43300,N_43023,N_43158);
xnor U43301 (N_43301,N_43138,N_43058);
and U43302 (N_43302,N_43060,N_43221);
xnor U43303 (N_43303,N_43142,N_43208);
xnor U43304 (N_43304,N_43126,N_43081);
nor U43305 (N_43305,N_43041,N_43183);
and U43306 (N_43306,N_43178,N_43240);
or U43307 (N_43307,N_43187,N_43154);
or U43308 (N_43308,N_43005,N_43134);
xnor U43309 (N_43309,N_43140,N_43036);
xor U43310 (N_43310,N_43085,N_43168);
nand U43311 (N_43311,N_43177,N_43109);
and U43312 (N_43312,N_43190,N_43035);
or U43313 (N_43313,N_43099,N_43008);
nor U43314 (N_43314,N_43103,N_43119);
or U43315 (N_43315,N_43186,N_43243);
xnor U43316 (N_43316,N_43007,N_43223);
and U43317 (N_43317,N_43071,N_43045);
nor U43318 (N_43318,N_43110,N_43135);
nand U43319 (N_43319,N_43055,N_43238);
nor U43320 (N_43320,N_43022,N_43149);
and U43321 (N_43321,N_43157,N_43040);
or U43322 (N_43322,N_43048,N_43179);
and U43323 (N_43323,N_43115,N_43124);
xor U43324 (N_43324,N_43104,N_43195);
nand U43325 (N_43325,N_43172,N_43042);
nand U43326 (N_43326,N_43122,N_43165);
and U43327 (N_43327,N_43148,N_43164);
and U43328 (N_43328,N_43169,N_43068);
or U43329 (N_43329,N_43201,N_43053);
and U43330 (N_43330,N_43249,N_43219);
and U43331 (N_43331,N_43108,N_43145);
xnor U43332 (N_43332,N_43146,N_43054);
nand U43333 (N_43333,N_43182,N_43235);
nand U43334 (N_43334,N_43229,N_43132);
xor U43335 (N_43335,N_43200,N_43176);
nand U43336 (N_43336,N_43114,N_43174);
or U43337 (N_43337,N_43028,N_43239);
and U43338 (N_43338,N_43202,N_43151);
xor U43339 (N_43339,N_43215,N_43030);
xnor U43340 (N_43340,N_43003,N_43143);
or U43341 (N_43341,N_43006,N_43153);
or U43342 (N_43342,N_43064,N_43077);
nand U43343 (N_43343,N_43069,N_43237);
nor U43344 (N_43344,N_43248,N_43094);
and U43345 (N_43345,N_43228,N_43074);
and U43346 (N_43346,N_43203,N_43086);
nor U43347 (N_43347,N_43002,N_43078);
nor U43348 (N_43348,N_43117,N_43227);
nor U43349 (N_43349,N_43160,N_43010);
and U43350 (N_43350,N_43072,N_43123);
and U43351 (N_43351,N_43020,N_43019);
nor U43352 (N_43352,N_43027,N_43106);
xnor U43353 (N_43353,N_43156,N_43216);
or U43354 (N_43354,N_43084,N_43167);
or U43355 (N_43355,N_43032,N_43205);
and U43356 (N_43356,N_43214,N_43043);
nor U43357 (N_43357,N_43031,N_43075);
nor U43358 (N_43358,N_43128,N_43211);
and U43359 (N_43359,N_43210,N_43033);
and U43360 (N_43360,N_43046,N_43105);
and U43361 (N_43361,N_43171,N_43038);
nor U43362 (N_43362,N_43136,N_43113);
and U43363 (N_43363,N_43017,N_43090);
and U43364 (N_43364,N_43185,N_43131);
and U43365 (N_43365,N_43213,N_43029);
and U43366 (N_43366,N_43065,N_43057);
nor U43367 (N_43367,N_43247,N_43088);
nand U43368 (N_43368,N_43225,N_43025);
nor U43369 (N_43369,N_43039,N_43082);
nor U43370 (N_43370,N_43218,N_43111);
or U43371 (N_43371,N_43204,N_43116);
xor U43372 (N_43372,N_43066,N_43018);
xnor U43373 (N_43373,N_43096,N_43076);
and U43374 (N_43374,N_43217,N_43021);
or U43375 (N_43375,N_43176,N_43174);
nor U43376 (N_43376,N_43003,N_43191);
or U43377 (N_43377,N_43179,N_43050);
xnor U43378 (N_43378,N_43103,N_43024);
nand U43379 (N_43379,N_43089,N_43000);
nor U43380 (N_43380,N_43227,N_43136);
xnor U43381 (N_43381,N_43242,N_43167);
and U43382 (N_43382,N_43131,N_43012);
or U43383 (N_43383,N_43215,N_43142);
xor U43384 (N_43384,N_43049,N_43021);
xnor U43385 (N_43385,N_43163,N_43045);
and U43386 (N_43386,N_43038,N_43229);
xor U43387 (N_43387,N_43190,N_43080);
or U43388 (N_43388,N_43055,N_43005);
nand U43389 (N_43389,N_43145,N_43110);
xor U43390 (N_43390,N_43191,N_43223);
nor U43391 (N_43391,N_43021,N_43047);
nand U43392 (N_43392,N_43105,N_43216);
and U43393 (N_43393,N_43004,N_43136);
and U43394 (N_43394,N_43156,N_43020);
nand U43395 (N_43395,N_43070,N_43172);
nand U43396 (N_43396,N_43171,N_43096);
xor U43397 (N_43397,N_43013,N_43041);
nor U43398 (N_43398,N_43191,N_43118);
nand U43399 (N_43399,N_43118,N_43037);
and U43400 (N_43400,N_43106,N_43217);
nand U43401 (N_43401,N_43209,N_43178);
nand U43402 (N_43402,N_43185,N_43020);
nor U43403 (N_43403,N_43168,N_43062);
xor U43404 (N_43404,N_43000,N_43112);
nor U43405 (N_43405,N_43019,N_43124);
nor U43406 (N_43406,N_43154,N_43168);
or U43407 (N_43407,N_43043,N_43094);
nor U43408 (N_43408,N_43245,N_43242);
nor U43409 (N_43409,N_43171,N_43066);
or U43410 (N_43410,N_43168,N_43188);
nand U43411 (N_43411,N_43150,N_43076);
xnor U43412 (N_43412,N_43162,N_43153);
nor U43413 (N_43413,N_43100,N_43094);
nor U43414 (N_43414,N_43109,N_43187);
nor U43415 (N_43415,N_43154,N_43150);
nor U43416 (N_43416,N_43075,N_43051);
nand U43417 (N_43417,N_43077,N_43021);
xnor U43418 (N_43418,N_43088,N_43160);
or U43419 (N_43419,N_43218,N_43086);
and U43420 (N_43420,N_43056,N_43220);
and U43421 (N_43421,N_43182,N_43217);
nor U43422 (N_43422,N_43249,N_43176);
nand U43423 (N_43423,N_43038,N_43200);
nand U43424 (N_43424,N_43015,N_43172);
nor U43425 (N_43425,N_43242,N_43050);
xnor U43426 (N_43426,N_43148,N_43120);
or U43427 (N_43427,N_43071,N_43091);
xor U43428 (N_43428,N_43143,N_43127);
xnor U43429 (N_43429,N_43166,N_43027);
or U43430 (N_43430,N_43185,N_43127);
and U43431 (N_43431,N_43122,N_43015);
and U43432 (N_43432,N_43166,N_43005);
and U43433 (N_43433,N_43237,N_43187);
xnor U43434 (N_43434,N_43058,N_43126);
and U43435 (N_43435,N_43119,N_43124);
xnor U43436 (N_43436,N_43209,N_43243);
nor U43437 (N_43437,N_43059,N_43115);
xnor U43438 (N_43438,N_43200,N_43006);
nor U43439 (N_43439,N_43186,N_43190);
and U43440 (N_43440,N_43065,N_43200);
or U43441 (N_43441,N_43194,N_43129);
nor U43442 (N_43442,N_43126,N_43038);
or U43443 (N_43443,N_43101,N_43019);
and U43444 (N_43444,N_43150,N_43243);
and U43445 (N_43445,N_43212,N_43174);
and U43446 (N_43446,N_43241,N_43246);
and U43447 (N_43447,N_43179,N_43108);
nand U43448 (N_43448,N_43032,N_43046);
or U43449 (N_43449,N_43055,N_43038);
nand U43450 (N_43450,N_43151,N_43180);
or U43451 (N_43451,N_43115,N_43211);
xor U43452 (N_43452,N_43240,N_43170);
nor U43453 (N_43453,N_43226,N_43127);
nor U43454 (N_43454,N_43193,N_43064);
nor U43455 (N_43455,N_43209,N_43137);
xor U43456 (N_43456,N_43211,N_43168);
xnor U43457 (N_43457,N_43092,N_43240);
xor U43458 (N_43458,N_43224,N_43111);
nand U43459 (N_43459,N_43159,N_43061);
xor U43460 (N_43460,N_43147,N_43182);
and U43461 (N_43461,N_43141,N_43123);
or U43462 (N_43462,N_43228,N_43191);
nand U43463 (N_43463,N_43072,N_43084);
nor U43464 (N_43464,N_43202,N_43166);
and U43465 (N_43465,N_43220,N_43207);
xnor U43466 (N_43466,N_43107,N_43103);
nor U43467 (N_43467,N_43217,N_43018);
nor U43468 (N_43468,N_43089,N_43075);
nor U43469 (N_43469,N_43079,N_43136);
nor U43470 (N_43470,N_43093,N_43185);
xor U43471 (N_43471,N_43249,N_43158);
nor U43472 (N_43472,N_43037,N_43021);
nor U43473 (N_43473,N_43064,N_43214);
or U43474 (N_43474,N_43237,N_43031);
nor U43475 (N_43475,N_43147,N_43165);
xor U43476 (N_43476,N_43141,N_43148);
or U43477 (N_43477,N_43155,N_43032);
nand U43478 (N_43478,N_43020,N_43177);
nand U43479 (N_43479,N_43067,N_43136);
and U43480 (N_43480,N_43046,N_43181);
nor U43481 (N_43481,N_43174,N_43196);
and U43482 (N_43482,N_43133,N_43007);
nand U43483 (N_43483,N_43208,N_43139);
or U43484 (N_43484,N_43108,N_43067);
nor U43485 (N_43485,N_43159,N_43167);
nand U43486 (N_43486,N_43199,N_43194);
nor U43487 (N_43487,N_43030,N_43129);
xor U43488 (N_43488,N_43231,N_43064);
nand U43489 (N_43489,N_43171,N_43030);
or U43490 (N_43490,N_43006,N_43191);
xnor U43491 (N_43491,N_43246,N_43204);
nand U43492 (N_43492,N_43135,N_43047);
nand U43493 (N_43493,N_43155,N_43188);
nor U43494 (N_43494,N_43220,N_43039);
and U43495 (N_43495,N_43047,N_43138);
and U43496 (N_43496,N_43091,N_43035);
and U43497 (N_43497,N_43065,N_43097);
or U43498 (N_43498,N_43094,N_43068);
and U43499 (N_43499,N_43055,N_43060);
nor U43500 (N_43500,N_43263,N_43269);
or U43501 (N_43501,N_43357,N_43377);
nor U43502 (N_43502,N_43259,N_43449);
and U43503 (N_43503,N_43329,N_43379);
nand U43504 (N_43504,N_43389,N_43468);
nor U43505 (N_43505,N_43312,N_43437);
xnor U43506 (N_43506,N_43302,N_43253);
nor U43507 (N_43507,N_43361,N_43447);
and U43508 (N_43508,N_43427,N_43484);
nor U43509 (N_43509,N_43303,N_43395);
or U43510 (N_43510,N_43463,N_43338);
nand U43511 (N_43511,N_43425,N_43494);
or U43512 (N_43512,N_43301,N_43290);
nor U43513 (N_43513,N_43268,N_43281);
and U43514 (N_43514,N_43260,N_43460);
nand U43515 (N_43515,N_43383,N_43288);
nand U43516 (N_43516,N_43470,N_43400);
and U43517 (N_43517,N_43336,N_43252);
and U43518 (N_43518,N_43315,N_43355);
or U43519 (N_43519,N_43490,N_43304);
or U43520 (N_43520,N_43365,N_43384);
nor U43521 (N_43521,N_43310,N_43420);
nand U43522 (N_43522,N_43471,N_43405);
xor U43523 (N_43523,N_43408,N_43331);
nand U43524 (N_43524,N_43495,N_43353);
nand U43525 (N_43525,N_43485,N_43350);
or U43526 (N_43526,N_43323,N_43373);
nand U43527 (N_43527,N_43345,N_43398);
and U43528 (N_43528,N_43300,N_43295);
or U43529 (N_43529,N_43363,N_43452);
xnor U43530 (N_43530,N_43284,N_43273);
xor U43531 (N_43531,N_43349,N_43382);
nand U43532 (N_43532,N_43407,N_43251);
xor U43533 (N_43533,N_43311,N_43413);
xor U43534 (N_43534,N_43326,N_43298);
xnor U43535 (N_43535,N_43374,N_43309);
nor U43536 (N_43536,N_43472,N_43354);
nor U43537 (N_43537,N_43411,N_43476);
nand U43538 (N_43538,N_43324,N_43313);
and U43539 (N_43539,N_43285,N_43428);
or U43540 (N_43540,N_43319,N_43487);
and U43541 (N_43541,N_43299,N_43258);
and U43542 (N_43542,N_43417,N_43335);
xnor U43543 (N_43543,N_43414,N_43360);
xor U43544 (N_43544,N_43435,N_43334);
nor U43545 (N_43545,N_43403,N_43356);
xor U43546 (N_43546,N_43318,N_43271);
and U43547 (N_43547,N_43364,N_43402);
nor U43548 (N_43548,N_43339,N_43283);
xnor U43549 (N_43549,N_43386,N_43483);
nor U43550 (N_43550,N_43482,N_43293);
or U43551 (N_43551,N_43279,N_43453);
and U43552 (N_43552,N_43296,N_43343);
nor U43553 (N_43553,N_43404,N_43486);
nand U43554 (N_43554,N_43394,N_43358);
or U43555 (N_43555,N_43488,N_43433);
and U43556 (N_43556,N_43458,N_43392);
or U43557 (N_43557,N_43421,N_43305);
nor U43558 (N_43558,N_43391,N_43254);
xor U43559 (N_43559,N_43367,N_43352);
nand U43560 (N_43560,N_43390,N_43274);
nand U43561 (N_43561,N_43262,N_43492);
nor U43562 (N_43562,N_43321,N_43297);
xor U43563 (N_43563,N_43448,N_43286);
nand U43564 (N_43564,N_43399,N_43451);
nor U43565 (N_43565,N_43489,N_43479);
nand U43566 (N_43566,N_43368,N_43340);
nor U43567 (N_43567,N_43422,N_43325);
xnor U43568 (N_43568,N_43426,N_43307);
nand U43569 (N_43569,N_43409,N_43292);
nor U43570 (N_43570,N_43278,N_43261);
and U43571 (N_43571,N_43450,N_43378);
nand U43572 (N_43572,N_43445,N_43276);
or U43573 (N_43573,N_43369,N_43475);
nor U43574 (N_43574,N_43320,N_43385);
xnor U43575 (N_43575,N_43439,N_43306);
and U43576 (N_43576,N_43346,N_43282);
and U43577 (N_43577,N_43491,N_43443);
and U43578 (N_43578,N_43376,N_43366);
or U43579 (N_43579,N_43255,N_43289);
and U43580 (N_43580,N_43351,N_43381);
nand U43581 (N_43581,N_43387,N_43478);
and U43582 (N_43582,N_43280,N_43308);
nand U43583 (N_43583,N_43322,N_43436);
and U43584 (N_43584,N_43375,N_43457);
and U43585 (N_43585,N_43393,N_43481);
and U43586 (N_43586,N_43294,N_43419);
nand U43587 (N_43587,N_43465,N_43431);
or U43588 (N_43588,N_43459,N_43477);
nor U43589 (N_43589,N_43498,N_43257);
nand U43590 (N_43590,N_43412,N_43497);
or U43591 (N_43591,N_43442,N_43397);
and U43592 (N_43592,N_43473,N_43444);
and U43593 (N_43593,N_43372,N_43332);
xor U43594 (N_43594,N_43266,N_43474);
xor U43595 (N_43595,N_43496,N_43330);
or U43596 (N_43596,N_43446,N_43359);
nor U43597 (N_43597,N_43440,N_43480);
xnor U43598 (N_43598,N_43270,N_43429);
nand U43599 (N_43599,N_43441,N_43423);
nor U43600 (N_43600,N_43265,N_43327);
nand U43601 (N_43601,N_43461,N_43410);
xor U43602 (N_43602,N_43264,N_43370);
xnor U43603 (N_43603,N_43462,N_43342);
xnor U43604 (N_43604,N_43316,N_43256);
nor U43605 (N_43605,N_43464,N_43499);
nand U43606 (N_43606,N_43467,N_43314);
nor U43607 (N_43607,N_43380,N_43493);
nand U43608 (N_43608,N_43416,N_43291);
xor U43609 (N_43609,N_43401,N_43424);
or U43610 (N_43610,N_43434,N_43347);
and U43611 (N_43611,N_43469,N_43348);
nand U43612 (N_43612,N_43415,N_43275);
xnor U43613 (N_43613,N_43277,N_43456);
nor U43614 (N_43614,N_43267,N_43328);
nor U43615 (N_43615,N_43396,N_43371);
nor U43616 (N_43616,N_43250,N_43344);
xnor U43617 (N_43617,N_43430,N_43406);
and U43618 (N_43618,N_43454,N_43333);
nand U43619 (N_43619,N_43455,N_43272);
or U43620 (N_43620,N_43362,N_43466);
and U43621 (N_43621,N_43418,N_43432);
nor U43622 (N_43622,N_43287,N_43317);
nor U43623 (N_43623,N_43438,N_43341);
or U43624 (N_43624,N_43388,N_43337);
nor U43625 (N_43625,N_43396,N_43353);
or U43626 (N_43626,N_43355,N_43470);
nand U43627 (N_43627,N_43420,N_43416);
and U43628 (N_43628,N_43466,N_43266);
nor U43629 (N_43629,N_43491,N_43372);
and U43630 (N_43630,N_43495,N_43478);
xor U43631 (N_43631,N_43366,N_43381);
and U43632 (N_43632,N_43418,N_43426);
xor U43633 (N_43633,N_43451,N_43325);
nand U43634 (N_43634,N_43438,N_43268);
and U43635 (N_43635,N_43253,N_43371);
nand U43636 (N_43636,N_43424,N_43341);
xor U43637 (N_43637,N_43364,N_43392);
nor U43638 (N_43638,N_43438,N_43308);
xor U43639 (N_43639,N_43407,N_43329);
or U43640 (N_43640,N_43306,N_43285);
nor U43641 (N_43641,N_43268,N_43258);
and U43642 (N_43642,N_43491,N_43301);
or U43643 (N_43643,N_43298,N_43344);
or U43644 (N_43644,N_43348,N_43344);
and U43645 (N_43645,N_43327,N_43345);
nor U43646 (N_43646,N_43428,N_43345);
or U43647 (N_43647,N_43405,N_43358);
nor U43648 (N_43648,N_43265,N_43470);
or U43649 (N_43649,N_43310,N_43404);
or U43650 (N_43650,N_43467,N_43301);
xor U43651 (N_43651,N_43348,N_43317);
and U43652 (N_43652,N_43448,N_43379);
and U43653 (N_43653,N_43397,N_43363);
nand U43654 (N_43654,N_43474,N_43499);
nor U43655 (N_43655,N_43345,N_43336);
or U43656 (N_43656,N_43450,N_43264);
nor U43657 (N_43657,N_43466,N_43341);
or U43658 (N_43658,N_43442,N_43411);
nor U43659 (N_43659,N_43295,N_43476);
nor U43660 (N_43660,N_43256,N_43497);
nor U43661 (N_43661,N_43428,N_43250);
and U43662 (N_43662,N_43272,N_43481);
nor U43663 (N_43663,N_43303,N_43287);
or U43664 (N_43664,N_43265,N_43437);
nand U43665 (N_43665,N_43338,N_43467);
or U43666 (N_43666,N_43411,N_43377);
nor U43667 (N_43667,N_43327,N_43277);
nor U43668 (N_43668,N_43365,N_43279);
nor U43669 (N_43669,N_43467,N_43326);
and U43670 (N_43670,N_43401,N_43302);
or U43671 (N_43671,N_43425,N_43311);
or U43672 (N_43672,N_43390,N_43438);
nand U43673 (N_43673,N_43256,N_43493);
nor U43674 (N_43674,N_43276,N_43396);
nand U43675 (N_43675,N_43385,N_43343);
and U43676 (N_43676,N_43433,N_43409);
or U43677 (N_43677,N_43333,N_43361);
or U43678 (N_43678,N_43389,N_43345);
or U43679 (N_43679,N_43331,N_43431);
and U43680 (N_43680,N_43310,N_43313);
or U43681 (N_43681,N_43299,N_43320);
xnor U43682 (N_43682,N_43359,N_43395);
and U43683 (N_43683,N_43280,N_43323);
nand U43684 (N_43684,N_43251,N_43412);
xor U43685 (N_43685,N_43447,N_43331);
and U43686 (N_43686,N_43499,N_43257);
nor U43687 (N_43687,N_43437,N_43264);
nor U43688 (N_43688,N_43494,N_43464);
xor U43689 (N_43689,N_43497,N_43435);
xnor U43690 (N_43690,N_43379,N_43432);
nor U43691 (N_43691,N_43265,N_43374);
xnor U43692 (N_43692,N_43468,N_43483);
or U43693 (N_43693,N_43305,N_43349);
xnor U43694 (N_43694,N_43389,N_43460);
and U43695 (N_43695,N_43362,N_43477);
nand U43696 (N_43696,N_43297,N_43459);
nor U43697 (N_43697,N_43268,N_43351);
xor U43698 (N_43698,N_43494,N_43296);
and U43699 (N_43699,N_43389,N_43271);
and U43700 (N_43700,N_43323,N_43263);
nor U43701 (N_43701,N_43284,N_43375);
xnor U43702 (N_43702,N_43464,N_43429);
and U43703 (N_43703,N_43250,N_43385);
or U43704 (N_43704,N_43423,N_43452);
and U43705 (N_43705,N_43466,N_43483);
nor U43706 (N_43706,N_43428,N_43452);
and U43707 (N_43707,N_43421,N_43440);
or U43708 (N_43708,N_43499,N_43416);
or U43709 (N_43709,N_43274,N_43474);
and U43710 (N_43710,N_43387,N_43274);
nor U43711 (N_43711,N_43365,N_43259);
and U43712 (N_43712,N_43454,N_43463);
nor U43713 (N_43713,N_43261,N_43447);
xor U43714 (N_43714,N_43484,N_43277);
nand U43715 (N_43715,N_43464,N_43348);
nor U43716 (N_43716,N_43475,N_43440);
and U43717 (N_43717,N_43278,N_43299);
and U43718 (N_43718,N_43259,N_43305);
nand U43719 (N_43719,N_43344,N_43296);
or U43720 (N_43720,N_43323,N_43312);
nand U43721 (N_43721,N_43499,N_43443);
and U43722 (N_43722,N_43378,N_43451);
xor U43723 (N_43723,N_43389,N_43344);
or U43724 (N_43724,N_43335,N_43293);
nand U43725 (N_43725,N_43363,N_43416);
and U43726 (N_43726,N_43429,N_43419);
nor U43727 (N_43727,N_43338,N_43445);
and U43728 (N_43728,N_43394,N_43367);
nand U43729 (N_43729,N_43353,N_43390);
nor U43730 (N_43730,N_43487,N_43310);
or U43731 (N_43731,N_43442,N_43370);
nand U43732 (N_43732,N_43348,N_43318);
and U43733 (N_43733,N_43322,N_43264);
and U43734 (N_43734,N_43288,N_43475);
nand U43735 (N_43735,N_43468,N_43335);
and U43736 (N_43736,N_43434,N_43474);
and U43737 (N_43737,N_43295,N_43343);
or U43738 (N_43738,N_43435,N_43403);
and U43739 (N_43739,N_43486,N_43450);
nand U43740 (N_43740,N_43383,N_43316);
xor U43741 (N_43741,N_43250,N_43468);
and U43742 (N_43742,N_43266,N_43383);
or U43743 (N_43743,N_43279,N_43384);
or U43744 (N_43744,N_43456,N_43428);
xor U43745 (N_43745,N_43458,N_43350);
or U43746 (N_43746,N_43449,N_43430);
or U43747 (N_43747,N_43314,N_43461);
nor U43748 (N_43748,N_43356,N_43317);
xnor U43749 (N_43749,N_43450,N_43276);
and U43750 (N_43750,N_43579,N_43670);
nand U43751 (N_43751,N_43689,N_43710);
xor U43752 (N_43752,N_43701,N_43527);
and U43753 (N_43753,N_43624,N_43682);
and U43754 (N_43754,N_43547,N_43673);
xor U43755 (N_43755,N_43655,N_43734);
or U43756 (N_43756,N_43525,N_43517);
nand U43757 (N_43757,N_43724,N_43551);
nor U43758 (N_43758,N_43535,N_43740);
or U43759 (N_43759,N_43668,N_43585);
xor U43760 (N_43760,N_43735,N_43694);
or U43761 (N_43761,N_43667,N_43516);
nand U43762 (N_43762,N_43588,N_43610);
and U43763 (N_43763,N_43681,N_43567);
or U43764 (N_43764,N_43559,N_43660);
and U43765 (N_43765,N_43538,N_43548);
nand U43766 (N_43766,N_43648,N_43572);
nor U43767 (N_43767,N_43631,N_43731);
or U43768 (N_43768,N_43738,N_43522);
or U43769 (N_43769,N_43571,N_43613);
or U43770 (N_43770,N_43537,N_43569);
nand U43771 (N_43771,N_43565,N_43623);
nand U43772 (N_43772,N_43545,N_43530);
xor U43773 (N_43773,N_43601,N_43683);
xnor U43774 (N_43774,N_43626,N_43697);
nand U43775 (N_43775,N_43594,N_43739);
and U43776 (N_43776,N_43533,N_43662);
nand U43777 (N_43777,N_43659,N_43730);
nor U43778 (N_43778,N_43645,N_43728);
nand U43779 (N_43779,N_43519,N_43581);
and U43780 (N_43780,N_43737,N_43675);
or U43781 (N_43781,N_43540,N_43693);
nor U43782 (N_43782,N_43564,N_43696);
or U43783 (N_43783,N_43621,N_43712);
and U43784 (N_43784,N_43709,N_43688);
nand U43785 (N_43785,N_43653,N_43515);
nor U43786 (N_43786,N_43713,N_43629);
nor U43787 (N_43787,N_43513,N_43566);
or U43788 (N_43788,N_43642,N_43619);
or U43789 (N_43789,N_43534,N_43528);
and U43790 (N_43790,N_43622,N_43598);
nor U43791 (N_43791,N_43716,N_43707);
xor U43792 (N_43792,N_43720,N_43555);
and U43793 (N_43793,N_43586,N_43666);
and U43794 (N_43794,N_43607,N_43634);
and U43795 (N_43795,N_43736,N_43745);
or U43796 (N_43796,N_43741,N_43557);
nor U43797 (N_43797,N_43597,N_43544);
or U43798 (N_43798,N_43742,N_43643);
nand U43799 (N_43799,N_43507,N_43531);
nor U43800 (N_43800,N_43636,N_43714);
and U43801 (N_43801,N_43614,N_43690);
xnor U43802 (N_43802,N_43568,N_43608);
nor U43803 (N_43803,N_43606,N_43502);
nor U43804 (N_43804,N_43590,N_43706);
and U43805 (N_43805,N_43529,N_43524);
nor U43806 (N_43806,N_43503,N_43677);
xor U43807 (N_43807,N_43721,N_43605);
or U43808 (N_43808,N_43576,N_43685);
nor U43809 (N_43809,N_43536,N_43695);
or U43810 (N_43810,N_43687,N_43711);
xnor U43811 (N_43811,N_43616,N_43518);
nor U43812 (N_43812,N_43640,N_43583);
and U43813 (N_43813,N_43592,N_43595);
xor U43814 (N_43814,N_43722,N_43725);
nand U43815 (N_43815,N_43599,N_43647);
or U43816 (N_43816,N_43663,N_43617);
or U43817 (N_43817,N_43732,N_43674);
xor U43818 (N_43818,N_43541,N_43676);
nor U43819 (N_43819,N_43542,N_43618);
nand U43820 (N_43820,N_43678,N_43723);
or U43821 (N_43821,N_43729,N_43644);
or U43822 (N_43822,N_43641,N_43703);
or U43823 (N_43823,N_43671,N_43661);
and U43824 (N_43824,N_43632,N_43511);
or U43825 (N_43825,N_43539,N_43749);
nand U43826 (N_43826,N_43684,N_43506);
nand U43827 (N_43827,N_43546,N_43652);
nand U43828 (N_43828,N_43727,N_43635);
nor U43829 (N_43829,N_43702,N_43639);
and U43830 (N_43830,N_43733,N_43554);
nor U43831 (N_43831,N_43698,N_43620);
nor U43832 (N_43832,N_43672,N_43669);
and U43833 (N_43833,N_43726,N_43532);
or U43834 (N_43834,N_43514,N_43501);
xor U43835 (N_43835,N_43549,N_43521);
xor U43836 (N_43836,N_43637,N_43717);
nor U43837 (N_43837,N_43651,N_43649);
or U43838 (N_43838,N_43657,N_43664);
nor U43839 (N_43839,N_43591,N_43679);
and U43840 (N_43840,N_43578,N_43561);
and U43841 (N_43841,N_43719,N_43615);
or U43842 (N_43842,N_43680,N_43705);
xor U43843 (N_43843,N_43563,N_43558);
xnor U43844 (N_43844,N_43743,N_43509);
and U43845 (N_43845,N_43704,N_43500);
nand U43846 (N_43846,N_43612,N_43654);
and U43847 (N_43847,N_43747,N_43505);
and U43848 (N_43848,N_43604,N_43589);
and U43849 (N_43849,N_43570,N_43746);
nor U43850 (N_43850,N_43718,N_43627);
xnor U43851 (N_43851,N_43552,N_43600);
xor U43852 (N_43852,N_43638,N_43510);
nor U43853 (N_43853,N_43625,N_43611);
nor U43854 (N_43854,N_43609,N_43512);
xor U43855 (N_43855,N_43692,N_43504);
xnor U43856 (N_43856,N_43577,N_43575);
nand U43857 (N_43857,N_43584,N_43656);
nor U43858 (N_43858,N_43553,N_43650);
nand U43859 (N_43859,N_43646,N_43665);
and U43860 (N_43860,N_43562,N_43630);
or U43861 (N_43861,N_43658,N_43526);
or U43862 (N_43862,N_43523,N_43596);
nand U43863 (N_43863,N_43580,N_43715);
or U43864 (N_43864,N_43633,N_43520);
nand U43865 (N_43865,N_43593,N_43744);
and U43866 (N_43866,N_43708,N_43602);
nand U43867 (N_43867,N_43700,N_43587);
or U43868 (N_43868,N_43691,N_43574);
xnor U43869 (N_43869,N_43582,N_43686);
xor U43870 (N_43870,N_43699,N_43748);
and U43871 (N_43871,N_43628,N_43560);
xor U43872 (N_43872,N_43573,N_43543);
and U43873 (N_43873,N_43603,N_43508);
xor U43874 (N_43874,N_43556,N_43550);
xnor U43875 (N_43875,N_43739,N_43515);
xnor U43876 (N_43876,N_43735,N_43610);
nor U43877 (N_43877,N_43717,N_43531);
and U43878 (N_43878,N_43573,N_43656);
nand U43879 (N_43879,N_43595,N_43562);
or U43880 (N_43880,N_43571,N_43537);
xor U43881 (N_43881,N_43540,N_43649);
nand U43882 (N_43882,N_43633,N_43643);
and U43883 (N_43883,N_43738,N_43589);
nand U43884 (N_43884,N_43615,N_43503);
nand U43885 (N_43885,N_43687,N_43673);
and U43886 (N_43886,N_43670,N_43711);
nand U43887 (N_43887,N_43572,N_43615);
nor U43888 (N_43888,N_43642,N_43651);
or U43889 (N_43889,N_43570,N_43522);
nor U43890 (N_43890,N_43729,N_43654);
nor U43891 (N_43891,N_43521,N_43573);
nand U43892 (N_43892,N_43602,N_43526);
nand U43893 (N_43893,N_43679,N_43566);
and U43894 (N_43894,N_43530,N_43562);
xor U43895 (N_43895,N_43657,N_43665);
and U43896 (N_43896,N_43683,N_43655);
or U43897 (N_43897,N_43636,N_43700);
or U43898 (N_43898,N_43593,N_43640);
and U43899 (N_43899,N_43527,N_43541);
and U43900 (N_43900,N_43683,N_43504);
nand U43901 (N_43901,N_43728,N_43729);
nand U43902 (N_43902,N_43707,N_43586);
nand U43903 (N_43903,N_43522,N_43648);
and U43904 (N_43904,N_43716,N_43712);
xor U43905 (N_43905,N_43591,N_43647);
and U43906 (N_43906,N_43525,N_43585);
and U43907 (N_43907,N_43609,N_43614);
nand U43908 (N_43908,N_43596,N_43627);
or U43909 (N_43909,N_43696,N_43658);
xnor U43910 (N_43910,N_43578,N_43732);
nand U43911 (N_43911,N_43724,N_43648);
or U43912 (N_43912,N_43529,N_43723);
nand U43913 (N_43913,N_43552,N_43685);
nor U43914 (N_43914,N_43607,N_43736);
nor U43915 (N_43915,N_43698,N_43715);
and U43916 (N_43916,N_43698,N_43564);
and U43917 (N_43917,N_43637,N_43635);
nand U43918 (N_43918,N_43517,N_43674);
or U43919 (N_43919,N_43700,N_43620);
and U43920 (N_43920,N_43705,N_43590);
nor U43921 (N_43921,N_43692,N_43651);
and U43922 (N_43922,N_43681,N_43588);
nor U43923 (N_43923,N_43587,N_43723);
xor U43924 (N_43924,N_43561,N_43545);
xnor U43925 (N_43925,N_43748,N_43656);
nand U43926 (N_43926,N_43528,N_43745);
xnor U43927 (N_43927,N_43748,N_43517);
nand U43928 (N_43928,N_43636,N_43652);
nand U43929 (N_43929,N_43513,N_43613);
or U43930 (N_43930,N_43699,N_43700);
xnor U43931 (N_43931,N_43746,N_43563);
nor U43932 (N_43932,N_43658,N_43625);
nand U43933 (N_43933,N_43745,N_43698);
or U43934 (N_43934,N_43645,N_43615);
or U43935 (N_43935,N_43748,N_43593);
and U43936 (N_43936,N_43744,N_43552);
or U43937 (N_43937,N_43743,N_43745);
nand U43938 (N_43938,N_43629,N_43625);
or U43939 (N_43939,N_43528,N_43676);
or U43940 (N_43940,N_43675,N_43625);
nor U43941 (N_43941,N_43726,N_43600);
and U43942 (N_43942,N_43685,N_43584);
or U43943 (N_43943,N_43596,N_43726);
nand U43944 (N_43944,N_43540,N_43525);
or U43945 (N_43945,N_43646,N_43531);
or U43946 (N_43946,N_43673,N_43698);
and U43947 (N_43947,N_43710,N_43573);
and U43948 (N_43948,N_43731,N_43661);
nand U43949 (N_43949,N_43636,N_43598);
nor U43950 (N_43950,N_43739,N_43702);
or U43951 (N_43951,N_43504,N_43658);
nor U43952 (N_43952,N_43692,N_43622);
and U43953 (N_43953,N_43687,N_43723);
or U43954 (N_43954,N_43528,N_43657);
nand U43955 (N_43955,N_43599,N_43591);
and U43956 (N_43956,N_43714,N_43723);
xnor U43957 (N_43957,N_43737,N_43733);
or U43958 (N_43958,N_43670,N_43500);
nand U43959 (N_43959,N_43673,N_43522);
nor U43960 (N_43960,N_43578,N_43635);
and U43961 (N_43961,N_43673,N_43503);
or U43962 (N_43962,N_43575,N_43668);
nand U43963 (N_43963,N_43685,N_43664);
and U43964 (N_43964,N_43669,N_43706);
and U43965 (N_43965,N_43549,N_43500);
or U43966 (N_43966,N_43581,N_43573);
nor U43967 (N_43967,N_43643,N_43654);
xor U43968 (N_43968,N_43646,N_43546);
nor U43969 (N_43969,N_43715,N_43666);
xnor U43970 (N_43970,N_43572,N_43535);
xor U43971 (N_43971,N_43725,N_43529);
or U43972 (N_43972,N_43725,N_43727);
and U43973 (N_43973,N_43579,N_43644);
nand U43974 (N_43974,N_43551,N_43586);
nor U43975 (N_43975,N_43709,N_43735);
nor U43976 (N_43976,N_43566,N_43576);
nor U43977 (N_43977,N_43610,N_43745);
and U43978 (N_43978,N_43587,N_43544);
xnor U43979 (N_43979,N_43738,N_43616);
and U43980 (N_43980,N_43542,N_43640);
xor U43981 (N_43981,N_43582,N_43530);
and U43982 (N_43982,N_43562,N_43633);
xor U43983 (N_43983,N_43595,N_43706);
nor U43984 (N_43984,N_43544,N_43695);
and U43985 (N_43985,N_43645,N_43682);
nand U43986 (N_43986,N_43732,N_43613);
or U43987 (N_43987,N_43716,N_43528);
nor U43988 (N_43988,N_43623,N_43684);
nor U43989 (N_43989,N_43598,N_43561);
and U43990 (N_43990,N_43691,N_43590);
or U43991 (N_43991,N_43664,N_43749);
nor U43992 (N_43992,N_43729,N_43748);
nor U43993 (N_43993,N_43729,N_43570);
xnor U43994 (N_43994,N_43717,N_43713);
nand U43995 (N_43995,N_43623,N_43615);
nand U43996 (N_43996,N_43571,N_43717);
xor U43997 (N_43997,N_43700,N_43599);
nand U43998 (N_43998,N_43593,N_43626);
nand U43999 (N_43999,N_43644,N_43665);
nor U44000 (N_44000,N_43957,N_43821);
nor U44001 (N_44001,N_43994,N_43816);
and U44002 (N_44002,N_43893,N_43909);
or U44003 (N_44003,N_43908,N_43935);
nor U44004 (N_44004,N_43879,N_43896);
and U44005 (N_44005,N_43880,N_43905);
and U44006 (N_44006,N_43841,N_43850);
nand U44007 (N_44007,N_43882,N_43982);
nor U44008 (N_44008,N_43911,N_43779);
or U44009 (N_44009,N_43795,N_43825);
nor U44010 (N_44010,N_43966,N_43972);
and U44011 (N_44011,N_43798,N_43752);
nand U44012 (N_44012,N_43832,N_43860);
or U44013 (N_44013,N_43848,N_43789);
xor U44014 (N_44014,N_43954,N_43854);
and U44015 (N_44015,N_43773,N_43857);
xor U44016 (N_44016,N_43822,N_43987);
nand U44017 (N_44017,N_43877,N_43891);
and U44018 (N_44018,N_43840,N_43923);
xor U44019 (N_44019,N_43791,N_43842);
or U44020 (N_44020,N_43792,N_43947);
and U44021 (N_44021,N_43975,N_43813);
or U44022 (N_44022,N_43885,N_43776);
or U44023 (N_44023,N_43912,N_43777);
xnor U44024 (N_44024,N_43871,N_43936);
and U44025 (N_44025,N_43800,N_43919);
or U44026 (N_44026,N_43844,N_43888);
xor U44027 (N_44027,N_43875,N_43944);
nor U44028 (N_44028,N_43764,N_43775);
and U44029 (N_44029,N_43805,N_43938);
and U44030 (N_44030,N_43759,N_43894);
or U44031 (N_44031,N_43945,N_43804);
xor U44032 (N_44032,N_43801,N_43851);
nor U44033 (N_44033,N_43784,N_43767);
xnor U44034 (N_44034,N_43810,N_43788);
or U44035 (N_44035,N_43811,N_43992);
or U44036 (N_44036,N_43937,N_43790);
nand U44037 (N_44037,N_43998,N_43918);
xnor U44038 (N_44038,N_43806,N_43861);
nand U44039 (N_44039,N_43815,N_43899);
xnor U44040 (N_44040,N_43887,N_43958);
and U44041 (N_44041,N_43950,N_43755);
xnor U44042 (N_44042,N_43809,N_43866);
and U44043 (N_44043,N_43874,N_43847);
and U44044 (N_44044,N_43897,N_43942);
xor U44045 (N_44045,N_43981,N_43985);
nor U44046 (N_44046,N_43837,N_43962);
nand U44047 (N_44047,N_43983,N_43758);
or U44048 (N_44048,N_43794,N_43756);
and U44049 (N_44049,N_43898,N_43886);
and U44050 (N_44050,N_43914,N_43974);
xor U44051 (N_44051,N_43979,N_43906);
nand U44052 (N_44052,N_43892,N_43922);
xor U44053 (N_44053,N_43910,N_43916);
xor U44054 (N_44054,N_43830,N_43807);
or U44055 (N_44055,N_43820,N_43951);
or U44056 (N_44056,N_43873,N_43797);
or U44057 (N_44057,N_43913,N_43754);
nand U44058 (N_44058,N_43943,N_43863);
nor U44059 (N_44059,N_43890,N_43929);
nor U44060 (N_44060,N_43819,N_43903);
xor U44061 (N_44061,N_43836,N_43997);
nand U44062 (N_44062,N_43814,N_43931);
or U44063 (N_44063,N_43991,N_43964);
nor U44064 (N_44064,N_43940,N_43865);
and U44065 (N_44065,N_43852,N_43802);
and U44066 (N_44066,N_43925,N_43753);
nand U44067 (N_44067,N_43955,N_43963);
xor U44068 (N_44068,N_43995,N_43883);
or U44069 (N_44069,N_43833,N_43986);
and U44070 (N_44070,N_43969,N_43780);
or U44071 (N_44071,N_43928,N_43799);
and U44072 (N_44072,N_43920,N_43818);
nor U44073 (N_44073,N_43926,N_43976);
nor U44074 (N_44074,N_43881,N_43774);
nand U44075 (N_44075,N_43952,N_43824);
and U44076 (N_44076,N_43783,N_43872);
and U44077 (N_44077,N_43803,N_43941);
nor U44078 (N_44078,N_43859,N_43868);
and U44079 (N_44079,N_43927,N_43769);
nor U44080 (N_44080,N_43930,N_43766);
nand U44081 (N_44081,N_43970,N_43956);
nor U44082 (N_44082,N_43771,N_43838);
or U44083 (N_44083,N_43978,N_43812);
or U44084 (N_44084,N_43867,N_43864);
xnor U44085 (N_44085,N_43924,N_43751);
xor U44086 (N_44086,N_43835,N_43946);
and U44087 (N_44087,N_43761,N_43826);
and U44088 (N_44088,N_43884,N_43827);
nor U44089 (N_44089,N_43853,N_43862);
nor U44090 (N_44090,N_43980,N_43990);
or U44091 (N_44091,N_43902,N_43900);
nand U44092 (N_44092,N_43787,N_43953);
nor U44093 (N_44093,N_43968,N_43977);
xnor U44094 (N_44094,N_43939,N_43770);
xnor U44095 (N_44095,N_43949,N_43829);
nand U44096 (N_44096,N_43993,N_43870);
nand U44097 (N_44097,N_43961,N_43750);
xor U44098 (N_44098,N_43869,N_43907);
nor U44099 (N_44099,N_43996,N_43843);
and U44100 (N_44100,N_43855,N_43895);
or U44101 (N_44101,N_43967,N_43760);
and U44102 (N_44102,N_43782,N_43793);
xnor U44103 (N_44103,N_43834,N_43757);
xor U44104 (N_44104,N_43762,N_43889);
nand U44105 (N_44105,N_43901,N_43768);
or U44106 (N_44106,N_43878,N_43959);
and U44107 (N_44107,N_43989,N_43817);
nor U44108 (N_44108,N_43988,N_43763);
xor U44109 (N_44109,N_43858,N_43839);
nand U44110 (N_44110,N_43846,N_43781);
and U44111 (N_44111,N_43786,N_43856);
nor U44112 (N_44112,N_43831,N_43904);
nand U44113 (N_44113,N_43828,N_43845);
or U44114 (N_44114,N_43849,N_43915);
xnor U44115 (N_44115,N_43823,N_43772);
and U44116 (N_44116,N_43765,N_43917);
and U44117 (N_44117,N_43999,N_43934);
or U44118 (N_44118,N_43965,N_43808);
nor U44119 (N_44119,N_43785,N_43876);
xor U44120 (N_44120,N_43921,N_43971);
or U44121 (N_44121,N_43933,N_43984);
xnor U44122 (N_44122,N_43960,N_43948);
or U44123 (N_44123,N_43973,N_43778);
nor U44124 (N_44124,N_43796,N_43932);
xnor U44125 (N_44125,N_43767,N_43856);
nor U44126 (N_44126,N_43786,N_43808);
and U44127 (N_44127,N_43915,N_43930);
nand U44128 (N_44128,N_43826,N_43978);
xor U44129 (N_44129,N_43916,N_43879);
nor U44130 (N_44130,N_43891,N_43979);
and U44131 (N_44131,N_43979,N_43816);
nor U44132 (N_44132,N_43950,N_43964);
xor U44133 (N_44133,N_43921,N_43800);
xnor U44134 (N_44134,N_43955,N_43759);
xnor U44135 (N_44135,N_43811,N_43871);
xnor U44136 (N_44136,N_43919,N_43980);
or U44137 (N_44137,N_43878,N_43920);
xor U44138 (N_44138,N_43975,N_43855);
xor U44139 (N_44139,N_43862,N_43779);
nor U44140 (N_44140,N_43942,N_43991);
nand U44141 (N_44141,N_43759,N_43771);
nor U44142 (N_44142,N_43868,N_43925);
and U44143 (N_44143,N_43822,N_43763);
nand U44144 (N_44144,N_43907,N_43963);
nor U44145 (N_44145,N_43845,N_43754);
and U44146 (N_44146,N_43898,N_43948);
nand U44147 (N_44147,N_43977,N_43874);
nand U44148 (N_44148,N_43947,N_43790);
nor U44149 (N_44149,N_43815,N_43830);
nand U44150 (N_44150,N_43842,N_43841);
nor U44151 (N_44151,N_43921,N_43935);
xor U44152 (N_44152,N_43968,N_43974);
or U44153 (N_44153,N_43859,N_43759);
nand U44154 (N_44154,N_43910,N_43854);
nand U44155 (N_44155,N_43944,N_43852);
and U44156 (N_44156,N_43920,N_43872);
or U44157 (N_44157,N_43953,N_43950);
nand U44158 (N_44158,N_43839,N_43899);
xnor U44159 (N_44159,N_43784,N_43942);
and U44160 (N_44160,N_43776,N_43752);
xor U44161 (N_44161,N_43779,N_43904);
and U44162 (N_44162,N_43982,N_43976);
or U44163 (N_44163,N_43951,N_43783);
xnor U44164 (N_44164,N_43818,N_43946);
nand U44165 (N_44165,N_43970,N_43943);
nand U44166 (N_44166,N_43843,N_43905);
nor U44167 (N_44167,N_43884,N_43940);
nand U44168 (N_44168,N_43919,N_43982);
nand U44169 (N_44169,N_43865,N_43780);
or U44170 (N_44170,N_43789,N_43853);
xnor U44171 (N_44171,N_43870,N_43850);
or U44172 (N_44172,N_43895,N_43954);
nor U44173 (N_44173,N_43921,N_43765);
and U44174 (N_44174,N_43980,N_43837);
and U44175 (N_44175,N_43834,N_43898);
xor U44176 (N_44176,N_43815,N_43925);
xor U44177 (N_44177,N_43879,N_43757);
nor U44178 (N_44178,N_43978,N_43913);
or U44179 (N_44179,N_43911,N_43762);
nor U44180 (N_44180,N_43969,N_43761);
xor U44181 (N_44181,N_43927,N_43956);
xnor U44182 (N_44182,N_43819,N_43753);
nand U44183 (N_44183,N_43821,N_43877);
nand U44184 (N_44184,N_43919,N_43827);
or U44185 (N_44185,N_43855,N_43963);
xnor U44186 (N_44186,N_43810,N_43818);
xor U44187 (N_44187,N_43809,N_43770);
xor U44188 (N_44188,N_43945,N_43987);
or U44189 (N_44189,N_43992,N_43960);
nand U44190 (N_44190,N_43865,N_43967);
nand U44191 (N_44191,N_43918,N_43867);
nand U44192 (N_44192,N_43873,N_43912);
xnor U44193 (N_44193,N_43873,N_43841);
nor U44194 (N_44194,N_43805,N_43779);
or U44195 (N_44195,N_43788,N_43766);
nand U44196 (N_44196,N_43962,N_43981);
or U44197 (N_44197,N_43891,N_43759);
or U44198 (N_44198,N_43990,N_43898);
and U44199 (N_44199,N_43995,N_43814);
nor U44200 (N_44200,N_43867,N_43790);
nor U44201 (N_44201,N_43876,N_43954);
and U44202 (N_44202,N_43883,N_43921);
and U44203 (N_44203,N_43906,N_43883);
nor U44204 (N_44204,N_43791,N_43978);
and U44205 (N_44205,N_43958,N_43917);
xor U44206 (N_44206,N_43849,N_43789);
nor U44207 (N_44207,N_43913,N_43864);
or U44208 (N_44208,N_43827,N_43899);
xor U44209 (N_44209,N_43995,N_43925);
and U44210 (N_44210,N_43850,N_43765);
nand U44211 (N_44211,N_43859,N_43774);
or U44212 (N_44212,N_43836,N_43890);
and U44213 (N_44213,N_43852,N_43890);
and U44214 (N_44214,N_43858,N_43926);
nor U44215 (N_44215,N_43877,N_43941);
nor U44216 (N_44216,N_43797,N_43772);
nor U44217 (N_44217,N_43872,N_43762);
nor U44218 (N_44218,N_43786,N_43860);
nor U44219 (N_44219,N_43910,N_43870);
nand U44220 (N_44220,N_43873,N_43934);
nor U44221 (N_44221,N_43784,N_43937);
and U44222 (N_44222,N_43941,N_43866);
xor U44223 (N_44223,N_43912,N_43941);
and U44224 (N_44224,N_43820,N_43883);
nor U44225 (N_44225,N_43804,N_43839);
nor U44226 (N_44226,N_43800,N_43853);
and U44227 (N_44227,N_43779,N_43969);
nand U44228 (N_44228,N_43928,N_43939);
xnor U44229 (N_44229,N_43838,N_43874);
nor U44230 (N_44230,N_43864,N_43937);
nand U44231 (N_44231,N_43845,N_43773);
and U44232 (N_44232,N_43896,N_43831);
nor U44233 (N_44233,N_43947,N_43797);
or U44234 (N_44234,N_43794,N_43751);
nor U44235 (N_44235,N_43959,N_43913);
nor U44236 (N_44236,N_43935,N_43907);
nand U44237 (N_44237,N_43842,N_43875);
or U44238 (N_44238,N_43843,N_43790);
nand U44239 (N_44239,N_43805,N_43834);
or U44240 (N_44240,N_43904,N_43918);
nand U44241 (N_44241,N_43775,N_43902);
nor U44242 (N_44242,N_43798,N_43776);
xor U44243 (N_44243,N_43991,N_43866);
xnor U44244 (N_44244,N_43901,N_43937);
or U44245 (N_44245,N_43978,N_43888);
nand U44246 (N_44246,N_43869,N_43945);
nor U44247 (N_44247,N_43805,N_43955);
and U44248 (N_44248,N_43899,N_43775);
and U44249 (N_44249,N_43901,N_43984);
nand U44250 (N_44250,N_44155,N_44103);
nor U44251 (N_44251,N_44125,N_44063);
xor U44252 (N_44252,N_44009,N_44120);
and U44253 (N_44253,N_44080,N_44151);
and U44254 (N_44254,N_44026,N_44025);
xnor U44255 (N_44255,N_44156,N_44087);
or U44256 (N_44256,N_44070,N_44170);
or U44257 (N_44257,N_44169,N_44124);
xor U44258 (N_44258,N_44003,N_44013);
nor U44259 (N_44259,N_44232,N_44054);
xnor U44260 (N_44260,N_44006,N_44056);
xor U44261 (N_44261,N_44100,N_44012);
or U44262 (N_44262,N_44098,N_44053);
nor U44263 (N_44263,N_44188,N_44183);
nand U44264 (N_44264,N_44007,N_44243);
xnor U44265 (N_44265,N_44206,N_44186);
nand U44266 (N_44266,N_44229,N_44237);
xnor U44267 (N_44267,N_44238,N_44085);
xor U44268 (N_44268,N_44131,N_44236);
or U44269 (N_44269,N_44011,N_44205);
and U44270 (N_44270,N_44076,N_44217);
nor U44271 (N_44271,N_44211,N_44041);
xnor U44272 (N_44272,N_44051,N_44212);
xnor U44273 (N_44273,N_44153,N_44075);
and U44274 (N_44274,N_44079,N_44168);
xor U44275 (N_44275,N_44016,N_44047);
and U44276 (N_44276,N_44044,N_44144);
or U44277 (N_44277,N_44118,N_44189);
xor U44278 (N_44278,N_44089,N_44132);
nand U44279 (N_44279,N_44223,N_44067);
xnor U44280 (N_44280,N_44241,N_44152);
xnor U44281 (N_44281,N_44059,N_44107);
nand U44282 (N_44282,N_44127,N_44015);
or U44283 (N_44283,N_44071,N_44165);
nand U44284 (N_44284,N_44240,N_44064);
nand U44285 (N_44285,N_44210,N_44109);
nor U44286 (N_44286,N_44163,N_44197);
xnor U44287 (N_44287,N_44086,N_44145);
nand U44288 (N_44288,N_44134,N_44018);
nand U44289 (N_44289,N_44180,N_44062);
and U44290 (N_44290,N_44113,N_44014);
nand U44291 (N_44291,N_44005,N_44058);
nand U44292 (N_44292,N_44001,N_44245);
nor U44293 (N_44293,N_44072,N_44239);
and U44294 (N_44294,N_44166,N_44038);
and U44295 (N_44295,N_44081,N_44046);
nand U44296 (N_44296,N_44181,N_44004);
or U44297 (N_44297,N_44213,N_44111);
or U44298 (N_44298,N_44108,N_44050);
or U44299 (N_44299,N_44105,N_44036);
nor U44300 (N_44300,N_44164,N_44101);
and U44301 (N_44301,N_44022,N_44179);
xnor U44302 (N_44302,N_44192,N_44214);
nor U44303 (N_44303,N_44052,N_44216);
and U44304 (N_44304,N_44147,N_44073);
nand U44305 (N_44305,N_44154,N_44141);
and U44306 (N_44306,N_44031,N_44077);
nand U44307 (N_44307,N_44193,N_44099);
xnor U44308 (N_44308,N_44116,N_44097);
and U44309 (N_44309,N_44083,N_44035);
xor U44310 (N_44310,N_44066,N_44142);
nor U44311 (N_44311,N_44167,N_44045);
or U44312 (N_44312,N_44225,N_44221);
or U44313 (N_44313,N_44202,N_44247);
and U44314 (N_44314,N_44162,N_44178);
xnor U44315 (N_44315,N_44017,N_44078);
xnor U44316 (N_44316,N_44104,N_44235);
xor U44317 (N_44317,N_44122,N_44133);
nor U44318 (N_44318,N_44149,N_44000);
nor U44319 (N_44319,N_44119,N_44138);
and U44320 (N_44320,N_44126,N_44090);
nand U44321 (N_44321,N_44224,N_44249);
nand U44322 (N_44322,N_44042,N_44204);
or U44323 (N_44323,N_44176,N_44084);
nand U44324 (N_44324,N_44061,N_44049);
or U44325 (N_44325,N_44195,N_44002);
or U44326 (N_44326,N_44030,N_44033);
nand U44327 (N_44327,N_44222,N_44032);
or U44328 (N_44328,N_44121,N_44123);
xnor U44329 (N_44329,N_44117,N_44174);
and U44330 (N_44330,N_44194,N_44048);
or U44331 (N_44331,N_44023,N_44233);
nand U44332 (N_44332,N_44248,N_44208);
nand U44333 (N_44333,N_44029,N_44034);
xnor U44334 (N_44334,N_44203,N_44021);
nand U44335 (N_44335,N_44220,N_44093);
or U44336 (N_44336,N_44028,N_44008);
nand U44337 (N_44337,N_44110,N_44158);
xnor U44338 (N_44338,N_44175,N_44129);
nor U44339 (N_44339,N_44200,N_44037);
and U44340 (N_44340,N_44136,N_44057);
nor U44341 (N_44341,N_44039,N_44095);
or U44342 (N_44342,N_44231,N_44173);
and U44343 (N_44343,N_44019,N_44114);
nor U44344 (N_44344,N_44027,N_44201);
or U44345 (N_44345,N_44159,N_44112);
xnor U44346 (N_44346,N_44157,N_44160);
nand U44347 (N_44347,N_44148,N_44040);
nand U44348 (N_44348,N_44184,N_44199);
nand U44349 (N_44349,N_44092,N_44219);
xnor U44350 (N_44350,N_44172,N_44242);
xnor U44351 (N_44351,N_44177,N_44182);
or U44352 (N_44352,N_44185,N_44060);
nand U44353 (N_44353,N_44102,N_44140);
nand U44354 (N_44354,N_44010,N_44198);
nor U44355 (N_44355,N_44094,N_44082);
or U44356 (N_44356,N_44139,N_44146);
and U44357 (N_44357,N_44074,N_44043);
and U44358 (N_44358,N_44137,N_44128);
nor U44359 (N_44359,N_44069,N_44190);
or U44360 (N_44360,N_44096,N_44115);
or U44361 (N_44361,N_44191,N_44068);
or U44362 (N_44362,N_44088,N_44228);
nand U44363 (N_44363,N_44187,N_44246);
xor U44364 (N_44364,N_44234,N_44227);
or U44365 (N_44365,N_44130,N_44150);
nand U44366 (N_44366,N_44065,N_44024);
and U44367 (N_44367,N_44161,N_44091);
or U44368 (N_44368,N_44218,N_44230);
or U44369 (N_44369,N_44055,N_44171);
and U44370 (N_44370,N_44226,N_44135);
xnor U44371 (N_44371,N_44020,N_44244);
nor U44372 (N_44372,N_44196,N_44209);
or U44373 (N_44373,N_44106,N_44215);
nor U44374 (N_44374,N_44143,N_44207);
nand U44375 (N_44375,N_44239,N_44091);
nand U44376 (N_44376,N_44138,N_44125);
xor U44377 (N_44377,N_44049,N_44048);
nor U44378 (N_44378,N_44192,N_44099);
nor U44379 (N_44379,N_44213,N_44066);
and U44380 (N_44380,N_44088,N_44027);
and U44381 (N_44381,N_44005,N_44078);
xor U44382 (N_44382,N_44075,N_44088);
and U44383 (N_44383,N_44227,N_44171);
and U44384 (N_44384,N_44020,N_44077);
or U44385 (N_44385,N_44043,N_44135);
nor U44386 (N_44386,N_44017,N_44186);
nand U44387 (N_44387,N_44131,N_44094);
or U44388 (N_44388,N_44126,N_44135);
or U44389 (N_44389,N_44102,N_44120);
nand U44390 (N_44390,N_44134,N_44205);
nor U44391 (N_44391,N_44191,N_44177);
nor U44392 (N_44392,N_44229,N_44110);
nor U44393 (N_44393,N_44008,N_44121);
nor U44394 (N_44394,N_44249,N_44213);
and U44395 (N_44395,N_44194,N_44079);
xor U44396 (N_44396,N_44242,N_44162);
or U44397 (N_44397,N_44118,N_44138);
xnor U44398 (N_44398,N_44241,N_44146);
or U44399 (N_44399,N_44163,N_44048);
or U44400 (N_44400,N_44022,N_44018);
xnor U44401 (N_44401,N_44213,N_44048);
or U44402 (N_44402,N_44079,N_44074);
and U44403 (N_44403,N_44135,N_44011);
xnor U44404 (N_44404,N_44074,N_44195);
or U44405 (N_44405,N_44087,N_44221);
and U44406 (N_44406,N_44115,N_44192);
nor U44407 (N_44407,N_44028,N_44007);
nor U44408 (N_44408,N_44246,N_44153);
nand U44409 (N_44409,N_44044,N_44111);
nand U44410 (N_44410,N_44066,N_44045);
or U44411 (N_44411,N_44158,N_44213);
or U44412 (N_44412,N_44199,N_44087);
and U44413 (N_44413,N_44057,N_44047);
nor U44414 (N_44414,N_44212,N_44031);
or U44415 (N_44415,N_44063,N_44061);
nand U44416 (N_44416,N_44135,N_44109);
nand U44417 (N_44417,N_44114,N_44069);
and U44418 (N_44418,N_44075,N_44010);
nand U44419 (N_44419,N_44018,N_44213);
and U44420 (N_44420,N_44200,N_44245);
nand U44421 (N_44421,N_44209,N_44115);
or U44422 (N_44422,N_44200,N_44047);
or U44423 (N_44423,N_44067,N_44022);
or U44424 (N_44424,N_44093,N_44064);
and U44425 (N_44425,N_44047,N_44086);
nand U44426 (N_44426,N_44233,N_44101);
and U44427 (N_44427,N_44039,N_44053);
xnor U44428 (N_44428,N_44048,N_44223);
xnor U44429 (N_44429,N_44164,N_44002);
or U44430 (N_44430,N_44081,N_44225);
nand U44431 (N_44431,N_44191,N_44162);
nand U44432 (N_44432,N_44024,N_44196);
nand U44433 (N_44433,N_44073,N_44081);
nand U44434 (N_44434,N_44114,N_44021);
or U44435 (N_44435,N_44065,N_44220);
nor U44436 (N_44436,N_44114,N_44131);
nor U44437 (N_44437,N_44102,N_44174);
and U44438 (N_44438,N_44070,N_44243);
and U44439 (N_44439,N_44214,N_44018);
nand U44440 (N_44440,N_44162,N_44011);
and U44441 (N_44441,N_44042,N_44061);
xor U44442 (N_44442,N_44120,N_44061);
xnor U44443 (N_44443,N_44171,N_44145);
and U44444 (N_44444,N_44242,N_44166);
nand U44445 (N_44445,N_44003,N_44245);
nor U44446 (N_44446,N_44083,N_44007);
nand U44447 (N_44447,N_44225,N_44169);
nor U44448 (N_44448,N_44178,N_44059);
nand U44449 (N_44449,N_44100,N_44007);
nor U44450 (N_44450,N_44214,N_44068);
or U44451 (N_44451,N_44026,N_44113);
and U44452 (N_44452,N_44152,N_44056);
nand U44453 (N_44453,N_44108,N_44248);
or U44454 (N_44454,N_44000,N_44097);
or U44455 (N_44455,N_44096,N_44127);
nor U44456 (N_44456,N_44168,N_44186);
xor U44457 (N_44457,N_44137,N_44204);
and U44458 (N_44458,N_44094,N_44242);
and U44459 (N_44459,N_44178,N_44123);
or U44460 (N_44460,N_44144,N_44248);
xor U44461 (N_44461,N_44043,N_44001);
nor U44462 (N_44462,N_44086,N_44210);
nor U44463 (N_44463,N_44203,N_44194);
xnor U44464 (N_44464,N_44025,N_44177);
and U44465 (N_44465,N_44061,N_44228);
nand U44466 (N_44466,N_44027,N_44211);
nor U44467 (N_44467,N_44016,N_44225);
nor U44468 (N_44468,N_44124,N_44107);
nor U44469 (N_44469,N_44129,N_44200);
and U44470 (N_44470,N_44237,N_44086);
or U44471 (N_44471,N_44214,N_44051);
nor U44472 (N_44472,N_44030,N_44197);
and U44473 (N_44473,N_44161,N_44038);
nor U44474 (N_44474,N_44148,N_44089);
xnor U44475 (N_44475,N_44030,N_44053);
nor U44476 (N_44476,N_44248,N_44133);
and U44477 (N_44477,N_44230,N_44121);
and U44478 (N_44478,N_44236,N_44227);
nor U44479 (N_44479,N_44193,N_44073);
xnor U44480 (N_44480,N_44122,N_44148);
and U44481 (N_44481,N_44139,N_44148);
nand U44482 (N_44482,N_44159,N_44107);
nor U44483 (N_44483,N_44055,N_44187);
or U44484 (N_44484,N_44186,N_44013);
or U44485 (N_44485,N_44232,N_44213);
or U44486 (N_44486,N_44201,N_44066);
nand U44487 (N_44487,N_44131,N_44117);
xnor U44488 (N_44488,N_44062,N_44056);
xnor U44489 (N_44489,N_44089,N_44243);
xor U44490 (N_44490,N_44076,N_44046);
and U44491 (N_44491,N_44236,N_44048);
or U44492 (N_44492,N_44134,N_44176);
and U44493 (N_44493,N_44116,N_44009);
nor U44494 (N_44494,N_44207,N_44078);
nor U44495 (N_44495,N_44196,N_44076);
and U44496 (N_44496,N_44095,N_44137);
nor U44497 (N_44497,N_44142,N_44199);
or U44498 (N_44498,N_44209,N_44052);
and U44499 (N_44499,N_44179,N_44119);
nand U44500 (N_44500,N_44263,N_44333);
and U44501 (N_44501,N_44486,N_44373);
or U44502 (N_44502,N_44446,N_44378);
nor U44503 (N_44503,N_44377,N_44488);
and U44504 (N_44504,N_44418,N_44459);
or U44505 (N_44505,N_44390,N_44289);
or U44506 (N_44506,N_44465,N_44318);
nor U44507 (N_44507,N_44272,N_44487);
nand U44508 (N_44508,N_44323,N_44284);
nor U44509 (N_44509,N_44331,N_44384);
xor U44510 (N_44510,N_44281,N_44343);
and U44511 (N_44511,N_44416,N_44382);
nor U44512 (N_44512,N_44385,N_44461);
or U44513 (N_44513,N_44463,N_44429);
xor U44514 (N_44514,N_44267,N_44477);
nand U44515 (N_44515,N_44351,N_44296);
or U44516 (N_44516,N_44256,N_44271);
and U44517 (N_44517,N_44346,N_44264);
nor U44518 (N_44518,N_44406,N_44401);
xor U44519 (N_44519,N_44324,N_44374);
or U44520 (N_44520,N_44475,N_44472);
nor U44521 (N_44521,N_44259,N_44376);
and U44522 (N_44522,N_44262,N_44454);
nand U44523 (N_44523,N_44365,N_44492);
and U44524 (N_44524,N_44438,N_44295);
or U44525 (N_44525,N_44345,N_44303);
or U44526 (N_44526,N_44404,N_44260);
xor U44527 (N_44527,N_44291,N_44321);
and U44528 (N_44528,N_44478,N_44474);
xnor U44529 (N_44529,N_44290,N_44252);
and U44530 (N_44530,N_44356,N_44400);
nor U44531 (N_44531,N_44358,N_44336);
and U44532 (N_44532,N_44425,N_44276);
or U44533 (N_44533,N_44370,N_44350);
xor U44534 (N_44534,N_44379,N_44326);
nor U44535 (N_44535,N_44444,N_44411);
nand U44536 (N_44536,N_44298,N_44435);
and U44537 (N_44537,N_44481,N_44431);
xor U44538 (N_44538,N_44457,N_44419);
and U44539 (N_44539,N_44311,N_44352);
nand U44540 (N_44540,N_44410,N_44279);
or U44541 (N_44541,N_44493,N_44497);
nor U44542 (N_44542,N_44433,N_44287);
and U44543 (N_44543,N_44338,N_44375);
nand U44544 (N_44544,N_44427,N_44319);
xor U44545 (N_44545,N_44316,N_44470);
nand U44546 (N_44546,N_44313,N_44368);
and U44547 (N_44547,N_44282,N_44408);
nand U44548 (N_44548,N_44304,N_44437);
nand U44549 (N_44549,N_44403,N_44428);
and U44550 (N_44550,N_44270,N_44367);
nor U44551 (N_44551,N_44369,N_44462);
or U44552 (N_44552,N_44394,N_44332);
nand U44553 (N_44553,N_44450,N_44327);
nand U44554 (N_44554,N_44468,N_44342);
nor U44555 (N_44555,N_44417,N_44274);
or U44556 (N_44556,N_44329,N_44440);
nand U44557 (N_44557,N_44380,N_44415);
or U44558 (N_44558,N_44261,N_44467);
and U44559 (N_44559,N_44347,N_44473);
xnor U44560 (N_44560,N_44344,N_44341);
nand U44561 (N_44561,N_44458,N_44426);
nand U44562 (N_44562,N_44335,N_44466);
xor U44563 (N_44563,N_44294,N_44489);
nand U44564 (N_44564,N_44453,N_44476);
nand U44565 (N_44565,N_44330,N_44273);
nand U44566 (N_44566,N_44275,N_44254);
and U44567 (N_44567,N_44307,N_44443);
or U44568 (N_44568,N_44381,N_44317);
xor U44569 (N_44569,N_44285,N_44334);
xor U44570 (N_44570,N_44395,N_44269);
or U44571 (N_44571,N_44409,N_44283);
or U44572 (N_44572,N_44396,N_44360);
and U44573 (N_44573,N_44402,N_44366);
and U44574 (N_44574,N_44300,N_44340);
nand U44575 (N_44575,N_44460,N_44251);
or U44576 (N_44576,N_44257,N_44325);
or U44577 (N_44577,N_44253,N_44349);
nand U44578 (N_44578,N_44495,N_44482);
or U44579 (N_44579,N_44471,N_44388);
and U44580 (N_44580,N_44391,N_44439);
xor U44581 (N_44581,N_44387,N_44310);
xnor U44582 (N_44582,N_44452,N_44315);
or U44583 (N_44583,N_44372,N_44302);
or U44584 (N_44584,N_44469,N_44484);
nand U44585 (N_44585,N_44359,N_44434);
or U44586 (N_44586,N_44420,N_44265);
and U44587 (N_44587,N_44292,N_44353);
xor U44588 (N_44588,N_44490,N_44485);
nand U44589 (N_44589,N_44424,N_44496);
nor U44590 (N_44590,N_44308,N_44309);
xnor U44591 (N_44591,N_44479,N_44286);
nand U44592 (N_44592,N_44445,N_44266);
nor U44593 (N_44593,N_44357,N_44337);
nor U44594 (N_44594,N_44413,N_44430);
nor U44595 (N_44595,N_44442,N_44299);
nand U44596 (N_44596,N_44389,N_44364);
xor U44597 (N_44597,N_44464,N_44314);
xor U44598 (N_44598,N_44328,N_44399);
nand U44599 (N_44599,N_44354,N_44361);
nand U44600 (N_44600,N_44405,N_44268);
and U44601 (N_44601,N_44250,N_44397);
and U44602 (N_44602,N_44494,N_44498);
xor U44603 (N_44603,N_44355,N_44393);
xor U44604 (N_44604,N_44436,N_44407);
xor U44605 (N_44605,N_44423,N_44448);
nand U44606 (N_44606,N_44322,N_44305);
and U44607 (N_44607,N_44306,N_44386);
nor U44608 (N_44608,N_44348,N_44339);
or U44609 (N_44609,N_44414,N_44432);
xnor U44610 (N_44610,N_44412,N_44447);
nor U44611 (N_44611,N_44301,N_44293);
nor U44612 (N_44612,N_44449,N_44288);
nand U44613 (N_44613,N_44383,N_44362);
nor U44614 (N_44614,N_44398,N_44312);
xor U44615 (N_44615,N_44280,N_44455);
or U44616 (N_44616,N_44451,N_44277);
or U44617 (N_44617,N_44483,N_44491);
xnor U44618 (N_44618,N_44255,N_44363);
and U44619 (N_44619,N_44441,N_44499);
nor U44620 (N_44620,N_44456,N_44421);
and U44621 (N_44621,N_44278,N_44320);
xor U44622 (N_44622,N_44480,N_44258);
or U44623 (N_44623,N_44392,N_44371);
nand U44624 (N_44624,N_44297,N_44422);
and U44625 (N_44625,N_44499,N_44470);
or U44626 (N_44626,N_44393,N_44310);
nor U44627 (N_44627,N_44291,N_44269);
and U44628 (N_44628,N_44499,N_44346);
and U44629 (N_44629,N_44378,N_44291);
nor U44630 (N_44630,N_44472,N_44363);
nor U44631 (N_44631,N_44375,N_44309);
xnor U44632 (N_44632,N_44263,N_44289);
and U44633 (N_44633,N_44259,N_44430);
xnor U44634 (N_44634,N_44256,N_44341);
xnor U44635 (N_44635,N_44358,N_44357);
or U44636 (N_44636,N_44446,N_44322);
and U44637 (N_44637,N_44436,N_44493);
xor U44638 (N_44638,N_44356,N_44304);
nor U44639 (N_44639,N_44455,N_44325);
and U44640 (N_44640,N_44262,N_44456);
nor U44641 (N_44641,N_44334,N_44403);
nand U44642 (N_44642,N_44355,N_44427);
xor U44643 (N_44643,N_44363,N_44269);
nand U44644 (N_44644,N_44447,N_44330);
nand U44645 (N_44645,N_44463,N_44274);
nand U44646 (N_44646,N_44433,N_44448);
or U44647 (N_44647,N_44342,N_44409);
nor U44648 (N_44648,N_44423,N_44426);
or U44649 (N_44649,N_44261,N_44417);
or U44650 (N_44650,N_44305,N_44445);
nor U44651 (N_44651,N_44341,N_44493);
or U44652 (N_44652,N_44413,N_44400);
xnor U44653 (N_44653,N_44446,N_44424);
nor U44654 (N_44654,N_44259,N_44295);
or U44655 (N_44655,N_44363,N_44375);
and U44656 (N_44656,N_44333,N_44444);
or U44657 (N_44657,N_44357,N_44442);
xnor U44658 (N_44658,N_44282,N_44359);
or U44659 (N_44659,N_44388,N_44481);
xor U44660 (N_44660,N_44488,N_44405);
and U44661 (N_44661,N_44443,N_44471);
nand U44662 (N_44662,N_44433,N_44454);
nor U44663 (N_44663,N_44287,N_44408);
or U44664 (N_44664,N_44487,N_44489);
nor U44665 (N_44665,N_44284,N_44308);
nand U44666 (N_44666,N_44345,N_44392);
or U44667 (N_44667,N_44413,N_44360);
nor U44668 (N_44668,N_44354,N_44304);
nand U44669 (N_44669,N_44399,N_44435);
nor U44670 (N_44670,N_44470,N_44410);
xor U44671 (N_44671,N_44332,N_44271);
xnor U44672 (N_44672,N_44357,N_44284);
xnor U44673 (N_44673,N_44297,N_44482);
and U44674 (N_44674,N_44408,N_44327);
and U44675 (N_44675,N_44430,N_44469);
xnor U44676 (N_44676,N_44351,N_44350);
and U44677 (N_44677,N_44414,N_44348);
nand U44678 (N_44678,N_44414,N_44472);
nand U44679 (N_44679,N_44499,N_44437);
nor U44680 (N_44680,N_44345,N_44424);
nor U44681 (N_44681,N_44256,N_44477);
xnor U44682 (N_44682,N_44427,N_44250);
nor U44683 (N_44683,N_44477,N_44321);
nand U44684 (N_44684,N_44283,N_44313);
and U44685 (N_44685,N_44356,N_44424);
or U44686 (N_44686,N_44324,N_44342);
and U44687 (N_44687,N_44324,N_44358);
xor U44688 (N_44688,N_44305,N_44250);
nor U44689 (N_44689,N_44308,N_44368);
xor U44690 (N_44690,N_44378,N_44258);
and U44691 (N_44691,N_44250,N_44422);
nor U44692 (N_44692,N_44307,N_44493);
nand U44693 (N_44693,N_44426,N_44331);
nor U44694 (N_44694,N_44319,N_44434);
nor U44695 (N_44695,N_44420,N_44317);
xnor U44696 (N_44696,N_44488,N_44368);
nor U44697 (N_44697,N_44283,N_44351);
nand U44698 (N_44698,N_44491,N_44362);
or U44699 (N_44699,N_44311,N_44343);
and U44700 (N_44700,N_44299,N_44449);
and U44701 (N_44701,N_44486,N_44442);
nor U44702 (N_44702,N_44477,N_44422);
nand U44703 (N_44703,N_44324,N_44440);
nand U44704 (N_44704,N_44341,N_44320);
xnor U44705 (N_44705,N_44410,N_44351);
xor U44706 (N_44706,N_44400,N_44496);
or U44707 (N_44707,N_44488,N_44370);
xor U44708 (N_44708,N_44400,N_44487);
and U44709 (N_44709,N_44484,N_44491);
nor U44710 (N_44710,N_44279,N_44337);
and U44711 (N_44711,N_44452,N_44349);
nand U44712 (N_44712,N_44287,N_44278);
xnor U44713 (N_44713,N_44374,N_44308);
nand U44714 (N_44714,N_44365,N_44391);
xor U44715 (N_44715,N_44367,N_44485);
nor U44716 (N_44716,N_44340,N_44468);
nand U44717 (N_44717,N_44296,N_44313);
or U44718 (N_44718,N_44314,N_44396);
nand U44719 (N_44719,N_44426,N_44422);
xnor U44720 (N_44720,N_44272,N_44358);
nor U44721 (N_44721,N_44345,N_44347);
and U44722 (N_44722,N_44357,N_44268);
nor U44723 (N_44723,N_44456,N_44263);
nand U44724 (N_44724,N_44281,N_44418);
or U44725 (N_44725,N_44369,N_44402);
nor U44726 (N_44726,N_44382,N_44285);
xor U44727 (N_44727,N_44260,N_44377);
and U44728 (N_44728,N_44302,N_44332);
or U44729 (N_44729,N_44297,N_44382);
nand U44730 (N_44730,N_44368,N_44290);
xor U44731 (N_44731,N_44491,N_44278);
nand U44732 (N_44732,N_44484,N_44304);
or U44733 (N_44733,N_44327,N_44260);
xor U44734 (N_44734,N_44486,N_44490);
xnor U44735 (N_44735,N_44422,N_44418);
nor U44736 (N_44736,N_44406,N_44323);
xnor U44737 (N_44737,N_44387,N_44379);
nor U44738 (N_44738,N_44282,N_44258);
or U44739 (N_44739,N_44297,N_44329);
and U44740 (N_44740,N_44334,N_44294);
nor U44741 (N_44741,N_44465,N_44467);
xnor U44742 (N_44742,N_44386,N_44420);
nor U44743 (N_44743,N_44297,N_44319);
nor U44744 (N_44744,N_44272,N_44301);
nor U44745 (N_44745,N_44499,N_44384);
nor U44746 (N_44746,N_44481,N_44281);
xnor U44747 (N_44747,N_44403,N_44438);
nand U44748 (N_44748,N_44334,N_44262);
nand U44749 (N_44749,N_44422,N_44359);
xnor U44750 (N_44750,N_44594,N_44603);
xor U44751 (N_44751,N_44682,N_44739);
xor U44752 (N_44752,N_44704,N_44742);
or U44753 (N_44753,N_44506,N_44659);
nor U44754 (N_44754,N_44644,N_44694);
nor U44755 (N_44755,N_44699,N_44620);
xor U44756 (N_44756,N_44714,N_44532);
or U44757 (N_44757,N_44636,N_44664);
nor U44758 (N_44758,N_44679,N_44528);
nor U44759 (N_44759,N_44721,N_44634);
and U44760 (N_44760,N_44529,N_44525);
and U44761 (N_44761,N_44635,N_44545);
or U44762 (N_44762,N_44558,N_44629);
and U44763 (N_44763,N_44514,N_44573);
nor U44764 (N_44764,N_44560,N_44672);
nor U44765 (N_44765,N_44590,N_44702);
xor U44766 (N_44766,N_44625,N_44658);
xnor U44767 (N_44767,N_44515,N_44678);
nor U44768 (N_44768,N_44556,N_44684);
nor U44769 (N_44769,N_44568,N_44745);
and U44770 (N_44770,N_44656,N_44578);
or U44771 (N_44771,N_44744,N_44643);
or U44772 (N_44772,N_44536,N_44674);
or U44773 (N_44773,N_44649,N_44716);
and U44774 (N_44774,N_44588,N_44623);
xnor U44775 (N_44775,N_44709,N_44681);
or U44776 (N_44776,N_44612,N_44576);
nor U44777 (N_44777,N_44557,N_44530);
and U44778 (N_44778,N_44692,N_44523);
and U44779 (N_44779,N_44639,N_44626);
nand U44780 (N_44780,N_44687,N_44749);
xor U44781 (N_44781,N_44516,N_44577);
and U44782 (N_44782,N_44628,N_44501);
and U44783 (N_44783,N_44593,N_44707);
or U44784 (N_44784,N_44615,N_44518);
xnor U44785 (N_44785,N_44574,N_44503);
nand U44786 (N_44786,N_44517,N_44711);
nor U44787 (N_44787,N_44554,N_44559);
xnor U44788 (N_44788,N_44617,N_44539);
nand U44789 (N_44789,N_44641,N_44662);
xor U44790 (N_44790,N_44671,N_44748);
nand U44791 (N_44791,N_44719,N_44686);
nor U44792 (N_44792,N_44604,N_44653);
or U44793 (N_44793,N_44570,N_44710);
nand U44794 (N_44794,N_44632,N_44567);
nand U44795 (N_44795,N_44630,N_44543);
xnor U44796 (N_44796,N_44601,N_44552);
xor U44797 (N_44797,N_44747,N_44737);
or U44798 (N_44798,N_44726,N_44610);
nand U44799 (N_44799,N_44645,N_44696);
nand U44800 (N_44800,N_44579,N_44685);
or U44801 (N_44801,N_44531,N_44602);
and U44802 (N_44802,N_44728,N_44691);
nor U44803 (N_44803,N_44580,N_44589);
or U44804 (N_44804,N_44740,N_44540);
nor U44805 (N_44805,N_44718,N_44583);
xor U44806 (N_44806,N_44591,N_44638);
nand U44807 (N_44807,N_44587,N_44542);
nor U44808 (N_44808,N_44586,N_44675);
or U44809 (N_44809,N_44655,N_44534);
nand U44810 (N_44810,N_44614,N_44698);
nand U44811 (N_44811,N_44519,N_44670);
xor U44812 (N_44812,N_44533,N_44510);
nor U44813 (N_44813,N_44613,N_44688);
or U44814 (N_44814,N_44693,N_44703);
nand U44815 (N_44815,N_44727,N_44673);
or U44816 (N_44816,N_44551,N_44722);
or U44817 (N_44817,N_44584,N_44652);
nor U44818 (N_44818,N_44697,N_44596);
and U44819 (N_44819,N_44526,N_44705);
nor U44820 (N_44820,N_44566,N_44544);
nor U44821 (N_44821,N_44650,N_44733);
xor U44822 (N_44822,N_44668,N_44723);
xor U44823 (N_44823,N_44700,N_44665);
nand U44824 (N_44824,N_44695,N_44535);
or U44825 (N_44825,N_44732,N_44606);
nor U44826 (N_44826,N_44564,N_44595);
nor U44827 (N_44827,N_44717,N_44735);
nor U44828 (N_44828,N_44637,N_44605);
xor U44829 (N_44829,N_44500,N_44555);
nand U44830 (N_44830,N_44575,N_44657);
xnor U44831 (N_44831,N_44712,N_44627);
and U44832 (N_44832,N_44548,N_44508);
xnor U44833 (N_44833,N_44608,N_44522);
xor U44834 (N_44834,N_44585,N_44729);
nor U44835 (N_44835,N_44553,N_44538);
nand U44836 (N_44836,N_44611,N_44549);
nor U44837 (N_44837,N_44565,N_44677);
xor U44838 (N_44838,N_44646,N_44736);
nand U44839 (N_44839,N_44746,N_44661);
xor U44840 (N_44840,N_44738,N_44502);
nor U44841 (N_44841,N_44730,N_44546);
or U44842 (N_44842,N_44743,N_44524);
or U44843 (N_44843,N_44631,N_44509);
and U44844 (N_44844,N_44724,N_44648);
xor U44845 (N_44845,N_44701,N_44507);
xnor U44846 (N_44846,N_44642,N_44572);
nand U44847 (N_44847,N_44689,N_44633);
xnor U44848 (N_44848,N_44725,N_44547);
or U44849 (N_44849,N_44599,N_44521);
xnor U44850 (N_44850,N_44640,N_44563);
and U44851 (N_44851,N_44561,N_44537);
and U44852 (N_44852,N_44663,N_44741);
or U44853 (N_44853,N_44571,N_44680);
xnor U44854 (N_44854,N_44667,N_44731);
and U44855 (N_44855,N_44651,N_44715);
nand U44856 (N_44856,N_44734,N_44708);
xnor U44857 (N_44857,N_44660,N_44624);
or U44858 (N_44858,N_44616,N_44706);
and U44859 (N_44859,N_44582,N_44666);
nand U44860 (N_44860,N_44720,N_44597);
or U44861 (N_44861,N_44609,N_44512);
nand U44862 (N_44862,N_44600,N_44550);
nand U44863 (N_44863,N_44713,N_44504);
xnor U44864 (N_44864,N_44592,N_44621);
and U44865 (N_44865,N_44581,N_44513);
xnor U44866 (N_44866,N_44505,N_44676);
or U44867 (N_44867,N_44541,N_44527);
xor U44868 (N_44868,N_44669,N_44647);
nand U44869 (N_44869,N_44619,N_44562);
and U44870 (N_44870,N_44690,N_44618);
nand U44871 (N_44871,N_44683,N_44520);
or U44872 (N_44872,N_44598,N_44622);
nand U44873 (N_44873,N_44511,N_44569);
xor U44874 (N_44874,N_44654,N_44607);
xor U44875 (N_44875,N_44705,N_44591);
nand U44876 (N_44876,N_44634,N_44512);
nor U44877 (N_44877,N_44640,N_44564);
and U44878 (N_44878,N_44665,N_44702);
and U44879 (N_44879,N_44694,N_44663);
or U44880 (N_44880,N_44746,N_44518);
xnor U44881 (N_44881,N_44582,N_44724);
nor U44882 (N_44882,N_44506,N_44660);
xnor U44883 (N_44883,N_44740,N_44607);
or U44884 (N_44884,N_44667,N_44592);
nand U44885 (N_44885,N_44662,N_44599);
nand U44886 (N_44886,N_44610,N_44647);
and U44887 (N_44887,N_44528,N_44730);
nor U44888 (N_44888,N_44712,N_44536);
or U44889 (N_44889,N_44553,N_44583);
nor U44890 (N_44890,N_44649,N_44539);
nor U44891 (N_44891,N_44588,N_44556);
nor U44892 (N_44892,N_44710,N_44715);
nand U44893 (N_44893,N_44600,N_44542);
nand U44894 (N_44894,N_44578,N_44660);
or U44895 (N_44895,N_44526,N_44707);
nand U44896 (N_44896,N_44526,N_44595);
or U44897 (N_44897,N_44594,N_44526);
xnor U44898 (N_44898,N_44703,N_44591);
or U44899 (N_44899,N_44597,N_44625);
nand U44900 (N_44900,N_44548,N_44647);
xor U44901 (N_44901,N_44608,N_44688);
xnor U44902 (N_44902,N_44601,N_44536);
and U44903 (N_44903,N_44560,N_44549);
nand U44904 (N_44904,N_44720,N_44693);
nand U44905 (N_44905,N_44667,N_44573);
or U44906 (N_44906,N_44509,N_44733);
or U44907 (N_44907,N_44592,N_44639);
or U44908 (N_44908,N_44740,N_44532);
nand U44909 (N_44909,N_44602,N_44669);
nor U44910 (N_44910,N_44573,N_44672);
xnor U44911 (N_44911,N_44729,N_44511);
nor U44912 (N_44912,N_44505,N_44612);
or U44913 (N_44913,N_44634,N_44646);
and U44914 (N_44914,N_44727,N_44588);
or U44915 (N_44915,N_44601,N_44515);
or U44916 (N_44916,N_44642,N_44589);
or U44917 (N_44917,N_44710,N_44692);
nor U44918 (N_44918,N_44528,N_44527);
or U44919 (N_44919,N_44586,N_44664);
nor U44920 (N_44920,N_44553,N_44566);
xnor U44921 (N_44921,N_44587,N_44683);
and U44922 (N_44922,N_44532,N_44627);
nand U44923 (N_44923,N_44675,N_44520);
nand U44924 (N_44924,N_44702,N_44724);
nand U44925 (N_44925,N_44575,N_44636);
nand U44926 (N_44926,N_44737,N_44607);
xor U44927 (N_44927,N_44577,N_44588);
nor U44928 (N_44928,N_44667,N_44646);
and U44929 (N_44929,N_44733,N_44665);
nor U44930 (N_44930,N_44566,N_44648);
nand U44931 (N_44931,N_44714,N_44622);
and U44932 (N_44932,N_44697,N_44641);
nor U44933 (N_44933,N_44590,N_44693);
or U44934 (N_44934,N_44686,N_44582);
nand U44935 (N_44935,N_44658,N_44709);
nand U44936 (N_44936,N_44559,N_44585);
nand U44937 (N_44937,N_44609,N_44611);
or U44938 (N_44938,N_44559,N_44724);
nand U44939 (N_44939,N_44548,N_44649);
nor U44940 (N_44940,N_44635,N_44648);
nand U44941 (N_44941,N_44663,N_44613);
nand U44942 (N_44942,N_44599,N_44706);
and U44943 (N_44943,N_44743,N_44583);
and U44944 (N_44944,N_44551,N_44634);
nand U44945 (N_44945,N_44662,N_44500);
nand U44946 (N_44946,N_44564,N_44733);
nor U44947 (N_44947,N_44625,N_44599);
xnor U44948 (N_44948,N_44619,N_44682);
nor U44949 (N_44949,N_44529,N_44574);
or U44950 (N_44950,N_44500,N_44671);
xor U44951 (N_44951,N_44683,N_44618);
nand U44952 (N_44952,N_44666,N_44624);
xnor U44953 (N_44953,N_44545,N_44744);
and U44954 (N_44954,N_44669,N_44598);
nor U44955 (N_44955,N_44717,N_44688);
nor U44956 (N_44956,N_44561,N_44679);
nand U44957 (N_44957,N_44668,N_44667);
xor U44958 (N_44958,N_44704,N_44684);
and U44959 (N_44959,N_44561,N_44574);
nand U44960 (N_44960,N_44733,N_44676);
xnor U44961 (N_44961,N_44592,N_44690);
or U44962 (N_44962,N_44701,N_44532);
nor U44963 (N_44963,N_44647,N_44569);
nand U44964 (N_44964,N_44744,N_44667);
xor U44965 (N_44965,N_44718,N_44631);
and U44966 (N_44966,N_44516,N_44730);
or U44967 (N_44967,N_44627,N_44660);
or U44968 (N_44968,N_44510,N_44541);
or U44969 (N_44969,N_44545,N_44529);
or U44970 (N_44970,N_44744,N_44560);
nor U44971 (N_44971,N_44587,N_44676);
and U44972 (N_44972,N_44726,N_44555);
or U44973 (N_44973,N_44694,N_44600);
xor U44974 (N_44974,N_44697,N_44716);
xnor U44975 (N_44975,N_44635,N_44511);
nor U44976 (N_44976,N_44514,N_44742);
nor U44977 (N_44977,N_44592,N_44524);
nand U44978 (N_44978,N_44725,N_44559);
nor U44979 (N_44979,N_44698,N_44586);
and U44980 (N_44980,N_44643,N_44706);
nor U44981 (N_44981,N_44510,N_44674);
xor U44982 (N_44982,N_44529,N_44715);
nor U44983 (N_44983,N_44595,N_44513);
nor U44984 (N_44984,N_44596,N_44731);
and U44985 (N_44985,N_44561,N_44664);
nand U44986 (N_44986,N_44640,N_44635);
xor U44987 (N_44987,N_44509,N_44516);
and U44988 (N_44988,N_44530,N_44561);
or U44989 (N_44989,N_44688,N_44524);
xor U44990 (N_44990,N_44580,N_44662);
nand U44991 (N_44991,N_44531,N_44591);
xor U44992 (N_44992,N_44566,N_44615);
and U44993 (N_44993,N_44683,N_44676);
and U44994 (N_44994,N_44601,N_44645);
nand U44995 (N_44995,N_44685,N_44526);
and U44996 (N_44996,N_44615,N_44520);
nor U44997 (N_44997,N_44630,N_44564);
and U44998 (N_44998,N_44549,N_44600);
nand U44999 (N_44999,N_44697,N_44510);
xnor U45000 (N_45000,N_44839,N_44966);
and U45001 (N_45001,N_44787,N_44952);
xnor U45002 (N_45002,N_44784,N_44865);
or U45003 (N_45003,N_44941,N_44778);
and U45004 (N_45004,N_44956,N_44867);
xor U45005 (N_45005,N_44883,N_44832);
nor U45006 (N_45006,N_44848,N_44926);
nor U45007 (N_45007,N_44997,N_44798);
or U45008 (N_45008,N_44938,N_44946);
nor U45009 (N_45009,N_44897,N_44769);
or U45010 (N_45010,N_44836,N_44820);
or U45011 (N_45011,N_44974,N_44880);
xnor U45012 (N_45012,N_44984,N_44898);
and U45013 (N_45013,N_44765,N_44965);
xor U45014 (N_45014,N_44870,N_44768);
xnor U45015 (N_45015,N_44850,N_44936);
xnor U45016 (N_45016,N_44849,N_44821);
xnor U45017 (N_45017,N_44766,N_44904);
and U45018 (N_45018,N_44864,N_44872);
or U45019 (N_45019,N_44847,N_44942);
xnor U45020 (N_45020,N_44875,N_44841);
nand U45021 (N_45021,N_44976,N_44893);
and U45022 (N_45022,N_44978,N_44969);
nand U45023 (N_45023,N_44868,N_44774);
or U45024 (N_45024,N_44822,N_44773);
xor U45025 (N_45025,N_44771,N_44921);
xor U45026 (N_45026,N_44959,N_44980);
or U45027 (N_45027,N_44902,N_44948);
or U45028 (N_45028,N_44947,N_44783);
xnor U45029 (N_45029,N_44801,N_44983);
xnor U45030 (N_45030,N_44923,N_44842);
nand U45031 (N_45031,N_44757,N_44927);
nor U45032 (N_45032,N_44857,N_44852);
xnor U45033 (N_45033,N_44805,N_44862);
and U45034 (N_45034,N_44789,N_44887);
or U45035 (N_45035,N_44991,N_44866);
and U45036 (N_45036,N_44754,N_44800);
or U45037 (N_45037,N_44854,N_44780);
nor U45038 (N_45038,N_44896,N_44845);
nor U45039 (N_45039,N_44964,N_44752);
xnor U45040 (N_45040,N_44933,N_44861);
or U45041 (N_45041,N_44871,N_44929);
nor U45042 (N_45042,N_44788,N_44953);
nand U45043 (N_45043,N_44891,N_44992);
xor U45044 (N_45044,N_44775,N_44881);
nand U45045 (N_45045,N_44796,N_44855);
or U45046 (N_45046,N_44934,N_44909);
nand U45047 (N_45047,N_44834,N_44753);
xor U45048 (N_45048,N_44970,N_44901);
nand U45049 (N_45049,N_44791,N_44825);
or U45050 (N_45050,N_44751,N_44826);
nor U45051 (N_45051,N_44975,N_44818);
xor U45052 (N_45052,N_44988,N_44874);
nand U45053 (N_45053,N_44790,N_44932);
or U45054 (N_45054,N_44761,N_44890);
or U45055 (N_45055,N_44985,N_44915);
nor U45056 (N_45056,N_44910,N_44908);
nor U45057 (N_45057,N_44920,N_44799);
nand U45058 (N_45058,N_44814,N_44989);
or U45059 (N_45059,N_44835,N_44859);
or U45060 (N_45060,N_44758,N_44802);
nand U45061 (N_45061,N_44990,N_44767);
nor U45062 (N_45062,N_44914,N_44999);
xor U45063 (N_45063,N_44782,N_44957);
or U45064 (N_45064,N_44876,N_44777);
xnor U45065 (N_45065,N_44981,N_44763);
or U45066 (N_45066,N_44844,N_44928);
and U45067 (N_45067,N_44776,N_44961);
or U45068 (N_45068,N_44828,N_44779);
or U45069 (N_45069,N_44967,N_44892);
xor U45070 (N_45070,N_44954,N_44905);
or U45071 (N_45071,N_44772,N_44907);
nor U45072 (N_45072,N_44808,N_44869);
nor U45073 (N_45073,N_44994,N_44837);
or U45074 (N_45074,N_44903,N_44860);
or U45075 (N_45075,N_44795,N_44829);
and U45076 (N_45076,N_44807,N_44918);
and U45077 (N_45077,N_44797,N_44770);
nand U45078 (N_45078,N_44949,N_44815);
nor U45079 (N_45079,N_44943,N_44838);
nor U45080 (N_45080,N_44786,N_44911);
nand U45081 (N_45081,N_44856,N_44863);
xnor U45082 (N_45082,N_44906,N_44996);
or U45083 (N_45083,N_44900,N_44810);
and U45084 (N_45084,N_44960,N_44972);
nor U45085 (N_45085,N_44979,N_44950);
nor U45086 (N_45086,N_44889,N_44830);
or U45087 (N_45087,N_44878,N_44931);
or U45088 (N_45088,N_44987,N_44827);
xnor U45089 (N_45089,N_44944,N_44917);
xnor U45090 (N_45090,N_44809,N_44803);
and U45091 (N_45091,N_44824,N_44785);
nor U45092 (N_45092,N_44937,N_44924);
and U45093 (N_45093,N_44884,N_44916);
xnor U45094 (N_45094,N_44846,N_44888);
or U45095 (N_45095,N_44968,N_44806);
nor U45096 (N_45096,N_44963,N_44885);
xor U45097 (N_45097,N_44811,N_44895);
nor U45098 (N_45098,N_44819,N_44879);
nor U45099 (N_45099,N_44945,N_44913);
or U45100 (N_45100,N_44958,N_44781);
nand U45101 (N_45101,N_44977,N_44899);
nor U45102 (N_45102,N_44804,N_44750);
nand U45103 (N_45103,N_44840,N_44764);
nor U45104 (N_45104,N_44919,N_44882);
or U45105 (N_45105,N_44762,N_44939);
nand U45106 (N_45106,N_44971,N_44935);
nand U45107 (N_45107,N_44951,N_44794);
nand U45108 (N_45108,N_44925,N_44792);
nand U45109 (N_45109,N_44955,N_44886);
nand U45110 (N_45110,N_44993,N_44986);
and U45111 (N_45111,N_44853,N_44755);
xor U45112 (N_45112,N_44759,N_44831);
xor U45113 (N_45113,N_44817,N_44962);
and U45114 (N_45114,N_44793,N_44998);
nand U45115 (N_45115,N_44873,N_44816);
and U45116 (N_45116,N_44922,N_44930);
nor U45117 (N_45117,N_44894,N_44812);
or U45118 (N_45118,N_44982,N_44823);
nand U45119 (N_45119,N_44858,N_44813);
or U45120 (N_45120,N_44995,N_44877);
or U45121 (N_45121,N_44973,N_44760);
nand U45122 (N_45122,N_44833,N_44940);
and U45123 (N_45123,N_44912,N_44843);
nor U45124 (N_45124,N_44851,N_44756);
nor U45125 (N_45125,N_44843,N_44768);
nand U45126 (N_45126,N_44765,N_44752);
and U45127 (N_45127,N_44874,N_44760);
nor U45128 (N_45128,N_44983,N_44813);
and U45129 (N_45129,N_44927,N_44824);
and U45130 (N_45130,N_44839,N_44951);
nor U45131 (N_45131,N_44822,N_44806);
and U45132 (N_45132,N_44883,N_44789);
nand U45133 (N_45133,N_44787,N_44862);
and U45134 (N_45134,N_44880,N_44823);
or U45135 (N_45135,N_44846,N_44988);
and U45136 (N_45136,N_44912,N_44949);
or U45137 (N_45137,N_44909,N_44827);
xor U45138 (N_45138,N_44840,N_44887);
or U45139 (N_45139,N_44770,N_44984);
or U45140 (N_45140,N_44816,N_44803);
nand U45141 (N_45141,N_44973,N_44755);
xor U45142 (N_45142,N_44885,N_44961);
nor U45143 (N_45143,N_44813,N_44824);
and U45144 (N_45144,N_44920,N_44960);
nand U45145 (N_45145,N_44896,N_44818);
nand U45146 (N_45146,N_44852,N_44958);
and U45147 (N_45147,N_44837,N_44878);
xnor U45148 (N_45148,N_44884,N_44935);
nand U45149 (N_45149,N_44951,N_44827);
and U45150 (N_45150,N_44805,N_44850);
nand U45151 (N_45151,N_44978,N_44870);
xnor U45152 (N_45152,N_44777,N_44873);
xnor U45153 (N_45153,N_44877,N_44878);
and U45154 (N_45154,N_44762,N_44904);
nand U45155 (N_45155,N_44765,N_44763);
or U45156 (N_45156,N_44815,N_44805);
xnor U45157 (N_45157,N_44864,N_44988);
xnor U45158 (N_45158,N_44859,N_44781);
nand U45159 (N_45159,N_44804,N_44908);
xor U45160 (N_45160,N_44979,N_44842);
or U45161 (N_45161,N_44848,N_44821);
nand U45162 (N_45162,N_44759,N_44764);
nor U45163 (N_45163,N_44924,N_44969);
nand U45164 (N_45164,N_44902,N_44807);
nor U45165 (N_45165,N_44874,N_44820);
nand U45166 (N_45166,N_44845,N_44819);
and U45167 (N_45167,N_44951,N_44869);
nor U45168 (N_45168,N_44959,N_44958);
nor U45169 (N_45169,N_44798,N_44805);
or U45170 (N_45170,N_44877,N_44915);
and U45171 (N_45171,N_44811,N_44752);
nor U45172 (N_45172,N_44870,N_44954);
and U45173 (N_45173,N_44826,N_44801);
nor U45174 (N_45174,N_44813,N_44935);
or U45175 (N_45175,N_44814,N_44798);
or U45176 (N_45176,N_44917,N_44849);
and U45177 (N_45177,N_44849,N_44855);
and U45178 (N_45178,N_44821,N_44990);
nor U45179 (N_45179,N_44814,N_44913);
nand U45180 (N_45180,N_44996,N_44821);
or U45181 (N_45181,N_44973,N_44851);
and U45182 (N_45182,N_44969,N_44910);
and U45183 (N_45183,N_44976,N_44751);
or U45184 (N_45184,N_44843,N_44971);
nand U45185 (N_45185,N_44981,N_44973);
xnor U45186 (N_45186,N_44921,N_44852);
or U45187 (N_45187,N_44778,N_44784);
nand U45188 (N_45188,N_44899,N_44761);
and U45189 (N_45189,N_44789,N_44875);
and U45190 (N_45190,N_44930,N_44841);
or U45191 (N_45191,N_44777,N_44768);
and U45192 (N_45192,N_44850,N_44952);
xor U45193 (N_45193,N_44861,N_44905);
xor U45194 (N_45194,N_44804,N_44809);
and U45195 (N_45195,N_44884,N_44780);
nor U45196 (N_45196,N_44759,N_44988);
nand U45197 (N_45197,N_44861,N_44815);
and U45198 (N_45198,N_44771,N_44982);
xnor U45199 (N_45199,N_44833,N_44891);
nand U45200 (N_45200,N_44891,N_44965);
xor U45201 (N_45201,N_44790,N_44902);
xnor U45202 (N_45202,N_44768,N_44818);
nand U45203 (N_45203,N_44996,N_44780);
nor U45204 (N_45204,N_44964,N_44852);
nor U45205 (N_45205,N_44942,N_44757);
xnor U45206 (N_45206,N_44966,N_44936);
or U45207 (N_45207,N_44813,N_44833);
xnor U45208 (N_45208,N_44995,N_44798);
and U45209 (N_45209,N_44881,N_44934);
nor U45210 (N_45210,N_44874,N_44862);
nand U45211 (N_45211,N_44942,N_44900);
xnor U45212 (N_45212,N_44775,N_44882);
and U45213 (N_45213,N_44962,N_44963);
xor U45214 (N_45214,N_44878,N_44966);
xnor U45215 (N_45215,N_44916,N_44933);
nor U45216 (N_45216,N_44853,N_44849);
and U45217 (N_45217,N_44753,N_44985);
or U45218 (N_45218,N_44962,N_44911);
and U45219 (N_45219,N_44857,N_44987);
nand U45220 (N_45220,N_44763,N_44967);
nand U45221 (N_45221,N_44876,N_44877);
xnor U45222 (N_45222,N_44997,N_44759);
or U45223 (N_45223,N_44811,N_44935);
or U45224 (N_45224,N_44907,N_44881);
or U45225 (N_45225,N_44961,N_44941);
xnor U45226 (N_45226,N_44765,N_44937);
nand U45227 (N_45227,N_44901,N_44914);
or U45228 (N_45228,N_44832,N_44793);
and U45229 (N_45229,N_44891,N_44984);
or U45230 (N_45230,N_44797,N_44923);
or U45231 (N_45231,N_44927,N_44931);
nor U45232 (N_45232,N_44934,N_44832);
xnor U45233 (N_45233,N_44896,N_44806);
and U45234 (N_45234,N_44949,N_44875);
or U45235 (N_45235,N_44913,N_44770);
xnor U45236 (N_45236,N_44776,N_44883);
or U45237 (N_45237,N_44873,N_44930);
xnor U45238 (N_45238,N_44823,N_44910);
nor U45239 (N_45239,N_44753,N_44917);
nor U45240 (N_45240,N_44831,N_44946);
or U45241 (N_45241,N_44922,N_44839);
nor U45242 (N_45242,N_44766,N_44824);
nor U45243 (N_45243,N_44780,N_44808);
nand U45244 (N_45244,N_44762,N_44985);
nand U45245 (N_45245,N_44965,N_44918);
or U45246 (N_45246,N_44808,N_44788);
or U45247 (N_45247,N_44894,N_44994);
xor U45248 (N_45248,N_44998,N_44981);
and U45249 (N_45249,N_44946,N_44875);
nand U45250 (N_45250,N_45063,N_45236);
xor U45251 (N_45251,N_45167,N_45068);
or U45252 (N_45252,N_45238,N_45042);
or U45253 (N_45253,N_45224,N_45216);
xnor U45254 (N_45254,N_45096,N_45044);
nor U45255 (N_45255,N_45230,N_45102);
xor U45256 (N_45256,N_45240,N_45060);
and U45257 (N_45257,N_45222,N_45225);
nand U45258 (N_45258,N_45032,N_45119);
and U45259 (N_45259,N_45145,N_45055);
xnor U45260 (N_45260,N_45004,N_45171);
and U45261 (N_45261,N_45066,N_45117);
and U45262 (N_45262,N_45116,N_45121);
nor U45263 (N_45263,N_45029,N_45056);
and U45264 (N_45264,N_45202,N_45003);
and U45265 (N_45265,N_45020,N_45192);
xor U45266 (N_45266,N_45128,N_45177);
xor U45267 (N_45267,N_45026,N_45181);
and U45268 (N_45268,N_45195,N_45191);
or U45269 (N_45269,N_45174,N_45212);
nor U45270 (N_45270,N_45111,N_45185);
or U45271 (N_45271,N_45197,N_45118);
xor U45272 (N_45272,N_45085,N_45069);
xor U45273 (N_45273,N_45126,N_45215);
or U45274 (N_45274,N_45208,N_45053);
nor U45275 (N_45275,N_45206,N_45107);
or U45276 (N_45276,N_45245,N_45156);
xor U45277 (N_45277,N_45144,N_45237);
nand U45278 (N_45278,N_45164,N_45048);
or U45279 (N_45279,N_45217,N_45084);
and U45280 (N_45280,N_45075,N_45155);
xnor U45281 (N_45281,N_45163,N_45140);
xnor U45282 (N_45282,N_45006,N_45039);
or U45283 (N_45283,N_45244,N_45194);
and U45284 (N_45284,N_45213,N_45046);
and U45285 (N_45285,N_45204,N_45227);
nand U45286 (N_45286,N_45147,N_45043);
xnor U45287 (N_45287,N_45207,N_45073);
and U45288 (N_45288,N_45114,N_45218);
nor U45289 (N_45289,N_45170,N_45062);
or U45290 (N_45290,N_45077,N_45049);
nand U45291 (N_45291,N_45072,N_45235);
or U45292 (N_45292,N_45078,N_45115);
nand U45293 (N_45293,N_45157,N_45133);
xor U45294 (N_45294,N_45221,N_45086);
xor U45295 (N_45295,N_45038,N_45205);
nand U45296 (N_45296,N_45033,N_45120);
and U45297 (N_45297,N_45027,N_45190);
and U45298 (N_45298,N_45247,N_45219);
and U45299 (N_45299,N_45008,N_45059);
nand U45300 (N_45300,N_45127,N_45090);
nand U45301 (N_45301,N_45129,N_45015);
and U45302 (N_45302,N_45154,N_45179);
nor U45303 (N_45303,N_45071,N_45249);
xnor U45304 (N_45304,N_45124,N_45143);
nor U45305 (N_45305,N_45104,N_45226);
nor U45306 (N_45306,N_45000,N_45100);
nand U45307 (N_45307,N_45248,N_45141);
or U45308 (N_45308,N_45138,N_45021);
xnor U45309 (N_45309,N_45035,N_45097);
and U45310 (N_45310,N_45011,N_45018);
and U45311 (N_45311,N_45228,N_45101);
and U45312 (N_45312,N_45074,N_45229);
nand U45313 (N_45313,N_45110,N_45223);
xor U45314 (N_45314,N_45178,N_45024);
xor U45315 (N_45315,N_45031,N_45176);
xor U45316 (N_45316,N_45189,N_45082);
xnor U45317 (N_45317,N_45007,N_45175);
nor U45318 (N_45318,N_45045,N_45095);
nor U45319 (N_45319,N_45054,N_45234);
or U45320 (N_45320,N_45025,N_45094);
nand U45321 (N_45321,N_45131,N_45040);
and U45322 (N_45322,N_45211,N_45142);
xnor U45323 (N_45323,N_45152,N_45182);
and U45324 (N_45324,N_45098,N_45162);
nor U45325 (N_45325,N_45091,N_45137);
xnor U45326 (N_45326,N_45123,N_45001);
nor U45327 (N_45327,N_45081,N_45243);
nor U45328 (N_45328,N_45186,N_45037);
nand U45329 (N_45329,N_45023,N_45231);
nor U45330 (N_45330,N_45013,N_45002);
xor U45331 (N_45331,N_45173,N_45028);
nor U45332 (N_45332,N_45076,N_45148);
and U45333 (N_45333,N_45187,N_45087);
nor U45334 (N_45334,N_45198,N_45088);
and U45335 (N_45335,N_45165,N_45122);
and U45336 (N_45336,N_45246,N_45103);
nor U45337 (N_45337,N_45161,N_45080);
nand U45338 (N_45338,N_45052,N_45134);
nand U45339 (N_45339,N_45064,N_45130);
xnor U45340 (N_45340,N_45005,N_45019);
or U45341 (N_45341,N_45172,N_45108);
and U45342 (N_45342,N_45201,N_45180);
xor U45343 (N_45343,N_45199,N_45022);
nor U45344 (N_45344,N_45188,N_45132);
nor U45345 (N_45345,N_45093,N_45061);
and U45346 (N_45346,N_45149,N_45193);
xnor U45347 (N_45347,N_45099,N_45051);
nor U45348 (N_45348,N_45214,N_45113);
xnor U45349 (N_45349,N_45158,N_45030);
xor U45350 (N_45350,N_45241,N_45233);
nor U45351 (N_45351,N_45196,N_45183);
or U45352 (N_45352,N_45017,N_45012);
nor U45353 (N_45353,N_45057,N_45210);
nor U45354 (N_45354,N_45112,N_45166);
nand U45355 (N_45355,N_45079,N_45016);
and U45356 (N_45356,N_45067,N_45200);
nor U45357 (N_45357,N_45047,N_45150);
nand U45358 (N_45358,N_45203,N_45050);
or U45359 (N_45359,N_45220,N_45036);
and U45360 (N_45360,N_45089,N_45065);
nand U45361 (N_45361,N_45151,N_45010);
xnor U45362 (N_45362,N_45034,N_45184);
and U45363 (N_45363,N_45058,N_45239);
nor U45364 (N_45364,N_45070,N_45153);
nand U45365 (N_45365,N_45160,N_45136);
nand U45366 (N_45366,N_45168,N_45209);
and U45367 (N_45367,N_45092,N_45009);
xnor U45368 (N_45368,N_45105,N_45106);
nand U45369 (N_45369,N_45242,N_45159);
nand U45370 (N_45370,N_45232,N_45169);
or U45371 (N_45371,N_45146,N_45041);
nand U45372 (N_45372,N_45014,N_45109);
xor U45373 (N_45373,N_45125,N_45139);
nand U45374 (N_45374,N_45135,N_45083);
or U45375 (N_45375,N_45150,N_45171);
and U45376 (N_45376,N_45202,N_45105);
nor U45377 (N_45377,N_45066,N_45184);
or U45378 (N_45378,N_45031,N_45206);
nor U45379 (N_45379,N_45089,N_45196);
and U45380 (N_45380,N_45180,N_45200);
nand U45381 (N_45381,N_45148,N_45050);
xnor U45382 (N_45382,N_45170,N_45156);
and U45383 (N_45383,N_45226,N_45016);
and U45384 (N_45384,N_45099,N_45142);
and U45385 (N_45385,N_45171,N_45196);
xnor U45386 (N_45386,N_45238,N_45101);
nor U45387 (N_45387,N_45183,N_45067);
nand U45388 (N_45388,N_45008,N_45009);
xnor U45389 (N_45389,N_45104,N_45010);
nand U45390 (N_45390,N_45177,N_45190);
or U45391 (N_45391,N_45118,N_45086);
or U45392 (N_45392,N_45030,N_45230);
nand U45393 (N_45393,N_45147,N_45067);
nand U45394 (N_45394,N_45066,N_45155);
and U45395 (N_45395,N_45031,N_45218);
nor U45396 (N_45396,N_45097,N_45221);
or U45397 (N_45397,N_45223,N_45192);
nand U45398 (N_45398,N_45036,N_45175);
nor U45399 (N_45399,N_45019,N_45060);
xor U45400 (N_45400,N_45234,N_45240);
nand U45401 (N_45401,N_45190,N_45078);
or U45402 (N_45402,N_45093,N_45043);
xnor U45403 (N_45403,N_45045,N_45213);
or U45404 (N_45404,N_45216,N_45075);
or U45405 (N_45405,N_45171,N_45060);
or U45406 (N_45406,N_45020,N_45004);
nor U45407 (N_45407,N_45045,N_45232);
xor U45408 (N_45408,N_45122,N_45215);
and U45409 (N_45409,N_45049,N_45217);
nor U45410 (N_45410,N_45180,N_45112);
or U45411 (N_45411,N_45172,N_45103);
and U45412 (N_45412,N_45129,N_45181);
xnor U45413 (N_45413,N_45012,N_45191);
nand U45414 (N_45414,N_45151,N_45067);
and U45415 (N_45415,N_45154,N_45160);
xor U45416 (N_45416,N_45249,N_45123);
xor U45417 (N_45417,N_45134,N_45012);
xnor U45418 (N_45418,N_45197,N_45211);
or U45419 (N_45419,N_45086,N_45232);
nand U45420 (N_45420,N_45051,N_45248);
and U45421 (N_45421,N_45105,N_45236);
nor U45422 (N_45422,N_45244,N_45030);
xor U45423 (N_45423,N_45041,N_45065);
nor U45424 (N_45424,N_45056,N_45124);
or U45425 (N_45425,N_45030,N_45108);
xor U45426 (N_45426,N_45231,N_45032);
or U45427 (N_45427,N_45045,N_45173);
and U45428 (N_45428,N_45244,N_45224);
nand U45429 (N_45429,N_45170,N_45146);
nand U45430 (N_45430,N_45025,N_45142);
and U45431 (N_45431,N_45177,N_45097);
or U45432 (N_45432,N_45149,N_45170);
and U45433 (N_45433,N_45078,N_45113);
nand U45434 (N_45434,N_45151,N_45156);
nor U45435 (N_45435,N_45021,N_45112);
and U45436 (N_45436,N_45196,N_45026);
nand U45437 (N_45437,N_45228,N_45024);
nand U45438 (N_45438,N_45136,N_45038);
or U45439 (N_45439,N_45209,N_45205);
xor U45440 (N_45440,N_45038,N_45213);
nand U45441 (N_45441,N_45199,N_45014);
or U45442 (N_45442,N_45117,N_45174);
xor U45443 (N_45443,N_45023,N_45142);
or U45444 (N_45444,N_45209,N_45077);
nor U45445 (N_45445,N_45104,N_45219);
or U45446 (N_45446,N_45018,N_45051);
and U45447 (N_45447,N_45248,N_45188);
xor U45448 (N_45448,N_45070,N_45060);
or U45449 (N_45449,N_45020,N_45110);
nand U45450 (N_45450,N_45054,N_45202);
or U45451 (N_45451,N_45152,N_45201);
xor U45452 (N_45452,N_45169,N_45036);
and U45453 (N_45453,N_45118,N_45016);
nor U45454 (N_45454,N_45205,N_45129);
xor U45455 (N_45455,N_45028,N_45122);
xor U45456 (N_45456,N_45154,N_45027);
and U45457 (N_45457,N_45096,N_45200);
or U45458 (N_45458,N_45044,N_45034);
xor U45459 (N_45459,N_45138,N_45228);
or U45460 (N_45460,N_45194,N_45128);
nand U45461 (N_45461,N_45163,N_45204);
or U45462 (N_45462,N_45227,N_45202);
xnor U45463 (N_45463,N_45171,N_45063);
nor U45464 (N_45464,N_45227,N_45198);
nor U45465 (N_45465,N_45247,N_45190);
and U45466 (N_45466,N_45061,N_45236);
xnor U45467 (N_45467,N_45006,N_45167);
xnor U45468 (N_45468,N_45116,N_45189);
nor U45469 (N_45469,N_45125,N_45032);
nor U45470 (N_45470,N_45037,N_45036);
xnor U45471 (N_45471,N_45196,N_45210);
nor U45472 (N_45472,N_45131,N_45048);
nand U45473 (N_45473,N_45191,N_45109);
xnor U45474 (N_45474,N_45235,N_45052);
nand U45475 (N_45475,N_45114,N_45171);
xnor U45476 (N_45476,N_45194,N_45010);
nor U45477 (N_45477,N_45112,N_45104);
nor U45478 (N_45478,N_45112,N_45128);
xnor U45479 (N_45479,N_45009,N_45220);
xnor U45480 (N_45480,N_45131,N_45090);
nand U45481 (N_45481,N_45220,N_45024);
and U45482 (N_45482,N_45187,N_45118);
or U45483 (N_45483,N_45085,N_45011);
nor U45484 (N_45484,N_45092,N_45241);
nand U45485 (N_45485,N_45215,N_45133);
nor U45486 (N_45486,N_45029,N_45064);
nand U45487 (N_45487,N_45234,N_45051);
or U45488 (N_45488,N_45213,N_45122);
and U45489 (N_45489,N_45039,N_45224);
nand U45490 (N_45490,N_45245,N_45241);
and U45491 (N_45491,N_45053,N_45100);
and U45492 (N_45492,N_45019,N_45227);
or U45493 (N_45493,N_45183,N_45079);
xnor U45494 (N_45494,N_45205,N_45220);
xor U45495 (N_45495,N_45170,N_45057);
xnor U45496 (N_45496,N_45249,N_45182);
xor U45497 (N_45497,N_45139,N_45131);
or U45498 (N_45498,N_45104,N_45193);
and U45499 (N_45499,N_45216,N_45120);
nand U45500 (N_45500,N_45338,N_45438);
xor U45501 (N_45501,N_45483,N_45266);
xnor U45502 (N_45502,N_45412,N_45420);
and U45503 (N_45503,N_45311,N_45271);
or U45504 (N_45504,N_45439,N_45335);
nor U45505 (N_45505,N_45470,N_45262);
nor U45506 (N_45506,N_45275,N_45449);
or U45507 (N_45507,N_45488,N_45278);
and U45508 (N_45508,N_45277,N_45291);
and U45509 (N_45509,N_45458,N_45253);
xnor U45510 (N_45510,N_45379,N_45364);
or U45511 (N_45511,N_45425,N_45313);
nor U45512 (N_45512,N_45382,N_45414);
and U45513 (N_45513,N_45497,N_45415);
or U45514 (N_45514,N_45268,N_45336);
nand U45515 (N_45515,N_45448,N_45442);
xor U45516 (N_45516,N_45484,N_45340);
xor U45517 (N_45517,N_45365,N_45467);
nor U45518 (N_45518,N_45490,N_45452);
and U45519 (N_45519,N_45304,N_45384);
nor U45520 (N_45520,N_45369,N_45295);
xor U45521 (N_45521,N_45276,N_45435);
nand U45522 (N_45522,N_45389,N_45451);
nand U45523 (N_45523,N_45477,N_45487);
and U45524 (N_45524,N_45440,N_45436);
nor U45525 (N_45525,N_45399,N_45310);
xor U45526 (N_45526,N_45334,N_45454);
xor U45527 (N_45527,N_45355,N_45348);
and U45528 (N_45528,N_45468,N_45472);
nand U45529 (N_45529,N_45402,N_45288);
xor U45530 (N_45530,N_45377,N_45281);
nand U45531 (N_45531,N_45492,N_45498);
nor U45532 (N_45532,N_45471,N_45250);
or U45533 (N_45533,N_45428,N_45434);
nor U45534 (N_45534,N_45322,N_45359);
nor U45535 (N_45535,N_45342,N_45330);
xor U45536 (N_45536,N_45318,N_45489);
nor U45537 (N_45537,N_45282,N_45352);
nand U45538 (N_45538,N_45427,N_45473);
or U45539 (N_45539,N_45287,N_45392);
nor U45540 (N_45540,N_45430,N_45475);
and U45541 (N_45541,N_45432,N_45286);
nand U45542 (N_45542,N_45418,N_45368);
xor U45543 (N_45543,N_45270,N_45301);
nand U45544 (N_45544,N_45387,N_45419);
nand U45545 (N_45545,N_45398,N_45491);
nor U45546 (N_45546,N_45325,N_45372);
and U45547 (N_45547,N_45395,N_45457);
or U45548 (N_45548,N_45424,N_45366);
xor U45549 (N_45549,N_45361,N_45303);
and U45550 (N_45550,N_45486,N_45423);
or U45551 (N_45551,N_45417,N_45476);
or U45552 (N_45552,N_45341,N_45347);
and U45553 (N_45553,N_45259,N_45307);
nor U45554 (N_45554,N_45328,N_45380);
or U45555 (N_45555,N_45280,N_45279);
nor U45556 (N_45556,N_45273,N_45465);
nor U45557 (N_45557,N_45381,N_45474);
xor U45558 (N_45558,N_45413,N_45390);
and U45559 (N_45559,N_45421,N_45370);
or U45560 (N_45560,N_45292,N_45385);
nand U45561 (N_45561,N_45314,N_45378);
nor U45562 (N_45562,N_45332,N_45496);
nand U45563 (N_45563,N_45263,N_45409);
nor U45564 (N_45564,N_45479,N_45437);
or U45565 (N_45565,N_45351,N_45255);
or U45566 (N_45566,N_45302,N_45323);
nand U45567 (N_45567,N_45422,N_45481);
xor U45568 (N_45568,N_45265,N_45353);
or U45569 (N_45569,N_45494,N_45499);
xor U45570 (N_45570,N_45356,N_45388);
or U45571 (N_45571,N_45459,N_45463);
and U45572 (N_45572,N_45290,N_45403);
nand U45573 (N_45573,N_45257,N_45344);
nand U45574 (N_45574,N_45357,N_45445);
xnor U45575 (N_45575,N_45376,N_45469);
nand U45576 (N_45576,N_45345,N_45408);
xnor U45577 (N_45577,N_45256,N_45383);
xnor U45578 (N_45578,N_45293,N_45315);
nor U45579 (N_45579,N_45316,N_45251);
and U45580 (N_45580,N_45258,N_45411);
xor U45581 (N_45581,N_45326,N_45349);
nor U45582 (N_45582,N_45444,N_45308);
nand U45583 (N_45583,N_45269,N_45324);
nand U45584 (N_45584,N_45371,N_45309);
xor U45585 (N_45585,N_45312,N_45297);
nor U45586 (N_45586,N_45289,N_45429);
and U45587 (N_45587,N_45393,N_45410);
nand U45588 (N_45588,N_45354,N_45358);
nand U45589 (N_45589,N_45296,N_45272);
nand U45590 (N_45590,N_45446,N_45493);
nand U45591 (N_45591,N_45329,N_45367);
nand U45592 (N_45592,N_45485,N_45337);
or U45593 (N_45593,N_45252,N_45283);
and U45594 (N_45594,N_45305,N_45274);
xnor U45595 (N_45595,N_45363,N_45455);
and U45596 (N_45596,N_45350,N_45401);
xnor U45597 (N_45597,N_45339,N_45396);
nand U45598 (N_45598,N_45298,N_45450);
or U45599 (N_45599,N_45333,N_45404);
and U45600 (N_45600,N_45306,N_45346);
and U45601 (N_45601,N_45285,N_45461);
and U45602 (N_45602,N_45391,N_45441);
xor U45603 (N_45603,N_45327,N_45299);
nand U45604 (N_45604,N_45362,N_45431);
or U45605 (N_45605,N_45447,N_45478);
xor U45606 (N_45606,N_45260,N_45453);
or U45607 (N_45607,N_45261,N_45406);
or U45608 (N_45608,N_45264,N_45375);
nand U45609 (N_45609,N_45300,N_45400);
and U45610 (N_45610,N_45394,N_45482);
nor U45611 (N_45611,N_45433,N_45407);
xnor U45612 (N_45612,N_45464,N_45374);
nand U45613 (N_45613,N_45320,N_45405);
xor U45614 (N_45614,N_45373,N_45386);
and U45615 (N_45615,N_45416,N_45466);
nor U45616 (N_45616,N_45294,N_45456);
xnor U45617 (N_45617,N_45321,N_45254);
nand U45618 (N_45618,N_45360,N_45317);
nand U45619 (N_45619,N_45443,N_45495);
nand U45620 (N_45620,N_45426,N_45460);
nor U45621 (N_45621,N_45397,N_45480);
nor U45622 (N_45622,N_45284,N_45267);
nor U45623 (N_45623,N_45331,N_45319);
nor U45624 (N_45624,N_45462,N_45343);
nor U45625 (N_45625,N_45258,N_45282);
nand U45626 (N_45626,N_45459,N_45397);
nor U45627 (N_45627,N_45453,N_45372);
xnor U45628 (N_45628,N_45312,N_45459);
nand U45629 (N_45629,N_45490,N_45288);
nor U45630 (N_45630,N_45270,N_45278);
nor U45631 (N_45631,N_45268,N_45294);
or U45632 (N_45632,N_45364,N_45257);
or U45633 (N_45633,N_45389,N_45429);
xnor U45634 (N_45634,N_45297,N_45355);
and U45635 (N_45635,N_45473,N_45485);
nor U45636 (N_45636,N_45327,N_45320);
nand U45637 (N_45637,N_45288,N_45499);
nor U45638 (N_45638,N_45265,N_45350);
nand U45639 (N_45639,N_45259,N_45494);
or U45640 (N_45640,N_45472,N_45451);
nor U45641 (N_45641,N_45316,N_45323);
nand U45642 (N_45642,N_45421,N_45453);
nor U45643 (N_45643,N_45308,N_45312);
nor U45644 (N_45644,N_45440,N_45327);
or U45645 (N_45645,N_45423,N_45354);
nand U45646 (N_45646,N_45345,N_45471);
nor U45647 (N_45647,N_45412,N_45368);
nand U45648 (N_45648,N_45301,N_45389);
nand U45649 (N_45649,N_45445,N_45295);
and U45650 (N_45650,N_45388,N_45484);
nand U45651 (N_45651,N_45488,N_45397);
xnor U45652 (N_45652,N_45422,N_45491);
nor U45653 (N_45653,N_45332,N_45292);
and U45654 (N_45654,N_45497,N_45492);
nand U45655 (N_45655,N_45402,N_45474);
nand U45656 (N_45656,N_45319,N_45442);
nand U45657 (N_45657,N_45319,N_45278);
nand U45658 (N_45658,N_45386,N_45365);
and U45659 (N_45659,N_45315,N_45488);
and U45660 (N_45660,N_45362,N_45254);
or U45661 (N_45661,N_45340,N_45466);
and U45662 (N_45662,N_45259,N_45381);
and U45663 (N_45663,N_45409,N_45267);
nor U45664 (N_45664,N_45295,N_45470);
nor U45665 (N_45665,N_45396,N_45466);
and U45666 (N_45666,N_45343,N_45428);
nand U45667 (N_45667,N_45298,N_45479);
xnor U45668 (N_45668,N_45476,N_45486);
and U45669 (N_45669,N_45446,N_45288);
xor U45670 (N_45670,N_45334,N_45399);
nor U45671 (N_45671,N_45498,N_45266);
xor U45672 (N_45672,N_45326,N_45488);
nor U45673 (N_45673,N_45434,N_45288);
and U45674 (N_45674,N_45328,N_45403);
nor U45675 (N_45675,N_45264,N_45330);
xnor U45676 (N_45676,N_45431,N_45449);
and U45677 (N_45677,N_45449,N_45457);
xnor U45678 (N_45678,N_45478,N_45446);
nor U45679 (N_45679,N_45353,N_45396);
and U45680 (N_45680,N_45438,N_45251);
nand U45681 (N_45681,N_45348,N_45304);
or U45682 (N_45682,N_45385,N_45313);
xor U45683 (N_45683,N_45271,N_45418);
nand U45684 (N_45684,N_45277,N_45468);
and U45685 (N_45685,N_45280,N_45464);
or U45686 (N_45686,N_45373,N_45313);
nand U45687 (N_45687,N_45354,N_45300);
nand U45688 (N_45688,N_45328,N_45497);
and U45689 (N_45689,N_45268,N_45483);
or U45690 (N_45690,N_45343,N_45315);
nor U45691 (N_45691,N_45328,N_45330);
and U45692 (N_45692,N_45495,N_45378);
nand U45693 (N_45693,N_45351,N_45309);
nand U45694 (N_45694,N_45349,N_45470);
nor U45695 (N_45695,N_45372,N_45366);
xor U45696 (N_45696,N_45476,N_45464);
xor U45697 (N_45697,N_45381,N_45461);
and U45698 (N_45698,N_45453,N_45279);
and U45699 (N_45699,N_45462,N_45487);
nor U45700 (N_45700,N_45427,N_45334);
and U45701 (N_45701,N_45345,N_45304);
or U45702 (N_45702,N_45464,N_45396);
and U45703 (N_45703,N_45399,N_45491);
nand U45704 (N_45704,N_45402,N_45408);
or U45705 (N_45705,N_45257,N_45327);
or U45706 (N_45706,N_45339,N_45281);
xor U45707 (N_45707,N_45348,N_45339);
xor U45708 (N_45708,N_45425,N_45302);
or U45709 (N_45709,N_45282,N_45460);
or U45710 (N_45710,N_45448,N_45397);
nand U45711 (N_45711,N_45295,N_45333);
nor U45712 (N_45712,N_45427,N_45405);
xnor U45713 (N_45713,N_45344,N_45326);
and U45714 (N_45714,N_45285,N_45392);
and U45715 (N_45715,N_45371,N_45301);
and U45716 (N_45716,N_45488,N_45417);
and U45717 (N_45717,N_45425,N_45456);
nor U45718 (N_45718,N_45478,N_45253);
xor U45719 (N_45719,N_45336,N_45309);
xnor U45720 (N_45720,N_45361,N_45294);
or U45721 (N_45721,N_45487,N_45292);
nand U45722 (N_45722,N_45277,N_45308);
or U45723 (N_45723,N_45398,N_45390);
nor U45724 (N_45724,N_45351,N_45488);
nor U45725 (N_45725,N_45272,N_45365);
xnor U45726 (N_45726,N_45382,N_45404);
or U45727 (N_45727,N_45433,N_45375);
nor U45728 (N_45728,N_45398,N_45427);
xor U45729 (N_45729,N_45402,N_45329);
nor U45730 (N_45730,N_45343,N_45423);
and U45731 (N_45731,N_45328,N_45320);
and U45732 (N_45732,N_45383,N_45456);
nand U45733 (N_45733,N_45319,N_45479);
and U45734 (N_45734,N_45499,N_45320);
xor U45735 (N_45735,N_45439,N_45267);
nor U45736 (N_45736,N_45252,N_45250);
nand U45737 (N_45737,N_45398,N_45293);
nor U45738 (N_45738,N_45407,N_45409);
or U45739 (N_45739,N_45251,N_45263);
or U45740 (N_45740,N_45451,N_45441);
nand U45741 (N_45741,N_45468,N_45381);
nor U45742 (N_45742,N_45435,N_45257);
nor U45743 (N_45743,N_45358,N_45394);
nor U45744 (N_45744,N_45377,N_45376);
and U45745 (N_45745,N_45415,N_45447);
and U45746 (N_45746,N_45350,N_45309);
nand U45747 (N_45747,N_45470,N_45494);
or U45748 (N_45748,N_45432,N_45463);
xor U45749 (N_45749,N_45364,N_45289);
nand U45750 (N_45750,N_45732,N_45627);
nand U45751 (N_45751,N_45731,N_45668);
nor U45752 (N_45752,N_45559,N_45584);
nand U45753 (N_45753,N_45666,N_45691);
nor U45754 (N_45754,N_45594,N_45625);
nor U45755 (N_45755,N_45516,N_45682);
or U45756 (N_45756,N_45500,N_45717);
and U45757 (N_45757,N_45733,N_45591);
nand U45758 (N_45758,N_45725,N_45607);
nand U45759 (N_45759,N_45694,N_45530);
nor U45760 (N_45760,N_45542,N_45609);
or U45761 (N_45761,N_45679,N_45661);
nand U45762 (N_45762,N_45599,N_45673);
nor U45763 (N_45763,N_45509,N_45653);
nand U45764 (N_45764,N_45512,N_45543);
xnor U45765 (N_45765,N_45616,N_45522);
and U45766 (N_45766,N_45620,N_45590);
nand U45767 (N_45767,N_45716,N_45748);
nor U45768 (N_45768,N_45556,N_45665);
xnor U45769 (N_45769,N_45645,N_45728);
xnor U45770 (N_45770,N_45592,N_45720);
nand U45771 (N_45771,N_45572,N_45739);
and U45772 (N_45772,N_45685,N_45528);
xnor U45773 (N_45773,N_45545,N_45547);
xor U45774 (N_45774,N_45686,N_45549);
xnor U45775 (N_45775,N_45575,N_45576);
nor U45776 (N_45776,N_45521,N_45713);
nand U45777 (N_45777,N_45611,N_45657);
xor U45778 (N_45778,N_45567,N_45714);
and U45779 (N_45779,N_45703,N_45568);
nand U45780 (N_45780,N_45631,N_45589);
nand U45781 (N_45781,N_45630,N_45534);
or U45782 (N_45782,N_45704,N_45747);
nand U45783 (N_45783,N_45532,N_45648);
nor U45784 (N_45784,N_45517,N_45523);
and U45785 (N_45785,N_45582,N_45684);
or U45786 (N_45786,N_45565,N_45636);
or U45787 (N_45787,N_45745,N_45535);
nand U45788 (N_45788,N_45672,N_45604);
nor U45789 (N_45789,N_45724,N_45707);
nor U45790 (N_45790,N_45678,N_45735);
and U45791 (N_45791,N_45730,N_45680);
nor U45792 (N_45792,N_45538,N_45554);
and U45793 (N_45793,N_45702,N_45524);
nand U45794 (N_45794,N_45660,N_45566);
nor U45795 (N_45795,N_45681,N_45629);
xnor U45796 (N_45796,N_45526,N_45688);
nand U45797 (N_45797,N_45581,N_45583);
nor U45798 (N_45798,N_45525,N_45573);
or U45799 (N_45799,N_45612,N_45708);
nor U45800 (N_45800,N_45503,N_45588);
and U45801 (N_45801,N_45706,N_45709);
nand U45802 (N_45802,N_45741,N_45555);
and U45803 (N_45803,N_45738,N_45608);
xnor U45804 (N_45804,N_45734,N_45676);
xor U45805 (N_45805,N_45654,N_45718);
or U45806 (N_45806,N_45602,N_45638);
nor U45807 (N_45807,N_45721,N_45643);
or U45808 (N_45808,N_45647,N_45719);
and U45809 (N_45809,N_45603,N_45705);
xnor U45810 (N_45810,N_45619,N_45670);
nand U45811 (N_45811,N_45507,N_45557);
xnor U45812 (N_45812,N_45552,N_45696);
nor U45813 (N_45813,N_45618,N_45729);
or U45814 (N_45814,N_45649,N_45511);
or U45815 (N_45815,N_45744,N_45628);
nand U45816 (N_45816,N_45715,N_45641);
or U45817 (N_45817,N_45737,N_45560);
or U45818 (N_45818,N_45674,N_45632);
xnor U45819 (N_45819,N_45601,N_45655);
xnor U45820 (N_45820,N_45743,N_45587);
nor U45821 (N_45821,N_45669,N_45656);
xor U45822 (N_45822,N_45699,N_45536);
xor U45823 (N_45823,N_45651,N_45692);
nand U45824 (N_45824,N_45546,N_45723);
nand U45825 (N_45825,N_45652,N_45659);
nor U45826 (N_45826,N_45623,N_45639);
and U45827 (N_45827,N_45613,N_45677);
nand U45828 (N_45828,N_45558,N_45675);
or U45829 (N_45829,N_45598,N_45504);
or U45830 (N_45830,N_45527,N_45640);
or U45831 (N_45831,N_45614,N_45501);
or U45832 (N_45832,N_45606,N_45624);
or U45833 (N_45833,N_45749,N_45510);
nand U45834 (N_45834,N_45637,N_45569);
nand U45835 (N_45835,N_45736,N_45615);
nand U45836 (N_45836,N_45626,N_45635);
nor U45837 (N_45837,N_45548,N_45617);
and U45838 (N_45838,N_45700,N_45701);
nor U45839 (N_45839,N_45519,N_45663);
or U45840 (N_45840,N_45553,N_45742);
nor U45841 (N_45841,N_45570,N_45710);
nand U45842 (N_45842,N_45574,N_45513);
nor U45843 (N_45843,N_45664,N_45506);
nor U45844 (N_45844,N_45667,N_45689);
xnor U45845 (N_45845,N_45644,N_45515);
or U45846 (N_45846,N_45502,N_45658);
xor U45847 (N_45847,N_45562,N_45621);
or U45848 (N_45848,N_45746,N_45633);
or U45849 (N_45849,N_45561,N_45508);
and U45850 (N_45850,N_45650,N_45726);
xnor U45851 (N_45851,N_45622,N_45571);
or U45852 (N_45852,N_45595,N_45693);
nand U45853 (N_45853,N_45520,N_45687);
and U45854 (N_45854,N_45531,N_45518);
or U45855 (N_45855,N_45533,N_45662);
or U45856 (N_45856,N_45697,N_45539);
nor U45857 (N_45857,N_45727,N_45540);
nand U45858 (N_45858,N_45605,N_45722);
xor U45859 (N_45859,N_45646,N_45579);
xor U45860 (N_45860,N_45695,N_45585);
or U45861 (N_45861,N_45580,N_45544);
and U45862 (N_45862,N_45537,N_45740);
nor U45863 (N_45863,N_45577,N_45642);
nor U45864 (N_45864,N_45593,N_45596);
nand U45865 (N_45865,N_45610,N_45550);
xor U45866 (N_45866,N_45711,N_45505);
nand U45867 (N_45867,N_45597,N_45634);
and U45868 (N_45868,N_45671,N_45683);
and U45869 (N_45869,N_45564,N_45578);
or U45870 (N_45870,N_45690,N_45514);
nand U45871 (N_45871,N_45551,N_45712);
nand U45872 (N_45872,N_45698,N_45541);
xor U45873 (N_45873,N_45529,N_45563);
xor U45874 (N_45874,N_45586,N_45600);
nor U45875 (N_45875,N_45733,N_45713);
xnor U45876 (N_45876,N_45654,N_45612);
or U45877 (N_45877,N_45611,N_45605);
nand U45878 (N_45878,N_45656,N_45745);
xnor U45879 (N_45879,N_45657,N_45503);
xnor U45880 (N_45880,N_45696,N_45560);
and U45881 (N_45881,N_45517,N_45583);
and U45882 (N_45882,N_45631,N_45744);
nand U45883 (N_45883,N_45540,N_45648);
nand U45884 (N_45884,N_45537,N_45670);
or U45885 (N_45885,N_45689,N_45603);
or U45886 (N_45886,N_45730,N_45698);
nor U45887 (N_45887,N_45504,N_45562);
and U45888 (N_45888,N_45584,N_45732);
nor U45889 (N_45889,N_45502,N_45653);
nor U45890 (N_45890,N_45595,N_45539);
or U45891 (N_45891,N_45568,N_45722);
nor U45892 (N_45892,N_45607,N_45648);
or U45893 (N_45893,N_45594,N_45545);
and U45894 (N_45894,N_45624,N_45670);
xor U45895 (N_45895,N_45608,N_45603);
nor U45896 (N_45896,N_45722,N_45567);
nand U45897 (N_45897,N_45636,N_45603);
nor U45898 (N_45898,N_45734,N_45571);
and U45899 (N_45899,N_45535,N_45621);
nand U45900 (N_45900,N_45593,N_45685);
xor U45901 (N_45901,N_45693,N_45623);
nand U45902 (N_45902,N_45627,N_45713);
or U45903 (N_45903,N_45586,N_45510);
xor U45904 (N_45904,N_45696,N_45592);
nor U45905 (N_45905,N_45654,N_45745);
nor U45906 (N_45906,N_45558,N_45544);
nor U45907 (N_45907,N_45566,N_45578);
nand U45908 (N_45908,N_45642,N_45716);
or U45909 (N_45909,N_45743,N_45573);
or U45910 (N_45910,N_45749,N_45594);
xnor U45911 (N_45911,N_45743,N_45588);
or U45912 (N_45912,N_45607,N_45621);
or U45913 (N_45913,N_45530,N_45617);
or U45914 (N_45914,N_45563,N_45550);
or U45915 (N_45915,N_45677,N_45618);
xor U45916 (N_45916,N_45577,N_45731);
nand U45917 (N_45917,N_45583,N_45597);
nand U45918 (N_45918,N_45725,N_45593);
or U45919 (N_45919,N_45503,N_45548);
nand U45920 (N_45920,N_45564,N_45737);
and U45921 (N_45921,N_45616,N_45512);
nor U45922 (N_45922,N_45652,N_45516);
xnor U45923 (N_45923,N_45629,N_45736);
and U45924 (N_45924,N_45720,N_45673);
xnor U45925 (N_45925,N_45559,N_45542);
and U45926 (N_45926,N_45513,N_45644);
nor U45927 (N_45927,N_45666,N_45673);
or U45928 (N_45928,N_45578,N_45595);
and U45929 (N_45929,N_45509,N_45522);
nand U45930 (N_45930,N_45526,N_45663);
nor U45931 (N_45931,N_45619,N_45738);
nand U45932 (N_45932,N_45573,N_45648);
nand U45933 (N_45933,N_45505,N_45666);
xnor U45934 (N_45934,N_45662,N_45577);
nand U45935 (N_45935,N_45577,N_45508);
xor U45936 (N_45936,N_45574,N_45524);
or U45937 (N_45937,N_45551,N_45542);
xnor U45938 (N_45938,N_45706,N_45575);
or U45939 (N_45939,N_45503,N_45641);
xor U45940 (N_45940,N_45528,N_45696);
and U45941 (N_45941,N_45663,N_45660);
and U45942 (N_45942,N_45545,N_45544);
xor U45943 (N_45943,N_45696,N_45642);
or U45944 (N_45944,N_45534,N_45526);
nor U45945 (N_45945,N_45643,N_45579);
nand U45946 (N_45946,N_45734,N_45749);
and U45947 (N_45947,N_45578,N_45742);
nand U45948 (N_45948,N_45629,N_45531);
nand U45949 (N_45949,N_45665,N_45502);
and U45950 (N_45950,N_45612,N_45698);
xor U45951 (N_45951,N_45647,N_45593);
nor U45952 (N_45952,N_45692,N_45711);
nand U45953 (N_45953,N_45685,N_45558);
or U45954 (N_45954,N_45510,N_45742);
nand U45955 (N_45955,N_45601,N_45618);
xor U45956 (N_45956,N_45726,N_45596);
xnor U45957 (N_45957,N_45544,N_45557);
nor U45958 (N_45958,N_45613,N_45557);
xnor U45959 (N_45959,N_45744,N_45528);
and U45960 (N_45960,N_45594,N_45627);
nand U45961 (N_45961,N_45733,N_45715);
or U45962 (N_45962,N_45581,N_45512);
and U45963 (N_45963,N_45711,N_45555);
or U45964 (N_45964,N_45513,N_45730);
and U45965 (N_45965,N_45617,N_45684);
xnor U45966 (N_45966,N_45672,N_45522);
xnor U45967 (N_45967,N_45629,N_45580);
xnor U45968 (N_45968,N_45709,N_45652);
or U45969 (N_45969,N_45737,N_45563);
and U45970 (N_45970,N_45575,N_45568);
xor U45971 (N_45971,N_45748,N_45615);
or U45972 (N_45972,N_45745,N_45718);
or U45973 (N_45973,N_45688,N_45534);
xnor U45974 (N_45974,N_45507,N_45663);
nor U45975 (N_45975,N_45551,N_45697);
and U45976 (N_45976,N_45737,N_45630);
xnor U45977 (N_45977,N_45571,N_45705);
nor U45978 (N_45978,N_45593,N_45598);
xnor U45979 (N_45979,N_45533,N_45648);
and U45980 (N_45980,N_45580,N_45741);
and U45981 (N_45981,N_45638,N_45691);
nor U45982 (N_45982,N_45731,N_45695);
nand U45983 (N_45983,N_45551,N_45596);
nor U45984 (N_45984,N_45611,N_45569);
or U45985 (N_45985,N_45691,N_45547);
nor U45986 (N_45986,N_45742,N_45512);
or U45987 (N_45987,N_45648,N_45512);
nor U45988 (N_45988,N_45709,N_45609);
and U45989 (N_45989,N_45703,N_45577);
nor U45990 (N_45990,N_45612,N_45676);
xnor U45991 (N_45991,N_45537,N_45746);
nor U45992 (N_45992,N_45510,N_45672);
and U45993 (N_45993,N_45715,N_45598);
nand U45994 (N_45994,N_45527,N_45611);
nor U45995 (N_45995,N_45527,N_45671);
or U45996 (N_45996,N_45605,N_45638);
nand U45997 (N_45997,N_45596,N_45731);
or U45998 (N_45998,N_45526,N_45737);
nand U45999 (N_45999,N_45599,N_45514);
nand U46000 (N_46000,N_45767,N_45908);
xnor U46001 (N_46001,N_45809,N_45762);
nor U46002 (N_46002,N_45931,N_45919);
and U46003 (N_46003,N_45753,N_45990);
and U46004 (N_46004,N_45832,N_45947);
or U46005 (N_46005,N_45840,N_45995);
xnor U46006 (N_46006,N_45813,N_45776);
xor U46007 (N_46007,N_45978,N_45921);
or U46008 (N_46008,N_45785,N_45885);
nor U46009 (N_46009,N_45872,N_45871);
or U46010 (N_46010,N_45792,N_45831);
xor U46011 (N_46011,N_45877,N_45865);
nand U46012 (N_46012,N_45864,N_45754);
nor U46013 (N_46013,N_45876,N_45909);
or U46014 (N_46014,N_45834,N_45996);
nor U46015 (N_46015,N_45860,N_45856);
or U46016 (N_46016,N_45882,N_45838);
nand U46017 (N_46017,N_45906,N_45853);
nor U46018 (N_46018,N_45970,N_45936);
nor U46019 (N_46019,N_45868,N_45966);
or U46020 (N_46020,N_45958,N_45823);
nand U46021 (N_46021,N_45752,N_45955);
or U46022 (N_46022,N_45957,N_45902);
nand U46023 (N_46023,N_45982,N_45769);
xor U46024 (N_46024,N_45898,N_45825);
xor U46025 (N_46025,N_45869,N_45822);
nand U46026 (N_46026,N_45848,N_45758);
or U46027 (N_46027,N_45858,N_45866);
and U46028 (N_46028,N_45784,N_45878);
xnor U46029 (N_46029,N_45816,N_45922);
xor U46030 (N_46030,N_45941,N_45857);
and U46031 (N_46031,N_45756,N_45818);
and U46032 (N_46032,N_45952,N_45802);
or U46033 (N_46033,N_45779,N_45992);
xnor U46034 (N_46034,N_45806,N_45965);
xnor U46035 (N_46035,N_45914,N_45988);
xor U46036 (N_46036,N_45855,N_45826);
and U46037 (N_46037,N_45974,N_45928);
nand U46038 (N_46038,N_45751,N_45913);
nor U46039 (N_46039,N_45789,N_45893);
nor U46040 (N_46040,N_45967,N_45994);
nor U46041 (N_46041,N_45973,N_45798);
and U46042 (N_46042,N_45963,N_45962);
and U46043 (N_46043,N_45803,N_45904);
or U46044 (N_46044,N_45924,N_45833);
and U46045 (N_46045,N_45900,N_45907);
nand U46046 (N_46046,N_45760,N_45911);
xor U46047 (N_46047,N_45766,N_45780);
and U46048 (N_46048,N_45942,N_45821);
nor U46049 (N_46049,N_45964,N_45937);
or U46050 (N_46050,N_45808,N_45793);
xnor U46051 (N_46051,N_45845,N_45873);
xor U46052 (N_46052,N_45997,N_45901);
nand U46053 (N_46053,N_45770,N_45917);
nand U46054 (N_46054,N_45910,N_45984);
or U46055 (N_46055,N_45943,N_45915);
and U46056 (N_46056,N_45815,N_45972);
or U46057 (N_46057,N_45875,N_45849);
xor U46058 (N_46058,N_45890,N_45774);
and U46059 (N_46059,N_45805,N_45899);
nor U46060 (N_46060,N_45926,N_45986);
or U46061 (N_46061,N_45794,N_45861);
nand U46062 (N_46062,N_45850,N_45896);
or U46063 (N_46063,N_45956,N_45842);
or U46064 (N_46064,N_45836,N_45847);
and U46065 (N_46065,N_45960,N_45980);
or U46066 (N_46066,N_45903,N_45920);
or U46067 (N_46067,N_45863,N_45940);
nand U46068 (N_46068,N_45773,N_45959);
nand U46069 (N_46069,N_45945,N_45880);
and U46070 (N_46070,N_45979,N_45824);
nand U46071 (N_46071,N_45837,N_45891);
xor U46072 (N_46072,N_45887,N_45846);
xor U46073 (N_46073,N_45985,N_45781);
xnor U46074 (N_46074,N_45918,N_45807);
or U46075 (N_46075,N_45987,N_45791);
xor U46076 (N_46076,N_45999,N_45977);
xor U46077 (N_46077,N_45843,N_45783);
nand U46078 (N_46078,N_45755,N_45835);
nand U46079 (N_46079,N_45870,N_45777);
nor U46080 (N_46080,N_45812,N_45881);
nand U46081 (N_46081,N_45796,N_45787);
xor U46082 (N_46082,N_45771,N_45772);
nand U46083 (N_46083,N_45892,N_45930);
and U46084 (N_46084,N_45757,N_45961);
nor U46085 (N_46085,N_45819,N_45799);
or U46086 (N_46086,N_45981,N_45932);
and U46087 (N_46087,N_45814,N_45968);
nor U46088 (N_46088,N_45929,N_45925);
nor U46089 (N_46089,N_45933,N_45879);
xnor U46090 (N_46090,N_45759,N_45804);
nor U46091 (N_46091,N_45829,N_45852);
and U46092 (N_46092,N_45788,N_45938);
and U46093 (N_46093,N_45927,N_45888);
xor U46094 (N_46094,N_45874,N_45763);
nor U46095 (N_46095,N_45976,N_45820);
nor U46096 (N_46096,N_45828,N_45750);
xnor U46097 (N_46097,N_45817,N_45889);
nand U46098 (N_46098,N_45948,N_45949);
and U46099 (N_46099,N_45884,N_45768);
or U46100 (N_46100,N_45954,N_45944);
nor U46101 (N_46101,N_45971,N_45934);
xor U46102 (N_46102,N_45867,N_45993);
nor U46103 (N_46103,N_45786,N_45883);
nor U46104 (N_46104,N_45841,N_45897);
and U46105 (N_46105,N_45991,N_45795);
or U46106 (N_46106,N_45946,N_45797);
and U46107 (N_46107,N_45975,N_45939);
nand U46108 (N_46108,N_45801,N_45839);
or U46109 (N_46109,N_45844,N_45905);
and U46110 (N_46110,N_45790,N_45827);
xnor U46111 (N_46111,N_45830,N_45859);
nor U46112 (N_46112,N_45778,N_45765);
and U46113 (N_46113,N_45761,N_45998);
nand U46114 (N_46114,N_45810,N_45912);
nand U46115 (N_46115,N_45951,N_45935);
nand U46116 (N_46116,N_45916,N_45775);
nor U46117 (N_46117,N_45764,N_45851);
xnor U46118 (N_46118,N_45894,N_45969);
nor U46119 (N_46119,N_45923,N_45989);
nand U46120 (N_46120,N_45953,N_45950);
xnor U46121 (N_46121,N_45886,N_45782);
xor U46122 (N_46122,N_45862,N_45854);
and U46123 (N_46123,N_45983,N_45800);
xnor U46124 (N_46124,N_45895,N_45811);
or U46125 (N_46125,N_45934,N_45820);
nand U46126 (N_46126,N_45988,N_45852);
nand U46127 (N_46127,N_45867,N_45989);
xnor U46128 (N_46128,N_45844,N_45773);
and U46129 (N_46129,N_45821,N_45813);
or U46130 (N_46130,N_45844,N_45792);
or U46131 (N_46131,N_45769,N_45978);
or U46132 (N_46132,N_45799,N_45863);
xor U46133 (N_46133,N_45927,N_45856);
or U46134 (N_46134,N_45939,N_45785);
nand U46135 (N_46135,N_45765,N_45831);
nor U46136 (N_46136,N_45856,N_45840);
and U46137 (N_46137,N_45848,N_45942);
nor U46138 (N_46138,N_45938,N_45877);
nand U46139 (N_46139,N_45831,N_45784);
and U46140 (N_46140,N_45804,N_45893);
and U46141 (N_46141,N_45899,N_45897);
nand U46142 (N_46142,N_45915,N_45768);
nand U46143 (N_46143,N_45790,N_45750);
nand U46144 (N_46144,N_45923,N_45790);
or U46145 (N_46145,N_45914,N_45774);
or U46146 (N_46146,N_45826,N_45986);
xnor U46147 (N_46147,N_45884,N_45772);
nand U46148 (N_46148,N_45853,N_45952);
nor U46149 (N_46149,N_45786,N_45917);
and U46150 (N_46150,N_45786,N_45851);
nor U46151 (N_46151,N_45783,N_45859);
nand U46152 (N_46152,N_45971,N_45859);
nand U46153 (N_46153,N_45840,N_45961);
and U46154 (N_46154,N_45844,N_45848);
xor U46155 (N_46155,N_45804,N_45927);
and U46156 (N_46156,N_45931,N_45962);
nand U46157 (N_46157,N_45918,N_45949);
nand U46158 (N_46158,N_45803,N_45929);
and U46159 (N_46159,N_45849,N_45923);
and U46160 (N_46160,N_45880,N_45909);
nand U46161 (N_46161,N_45975,N_45913);
nand U46162 (N_46162,N_45784,N_45817);
and U46163 (N_46163,N_45979,N_45814);
nand U46164 (N_46164,N_45970,N_45842);
and U46165 (N_46165,N_45957,N_45824);
and U46166 (N_46166,N_45981,N_45938);
nand U46167 (N_46167,N_45949,N_45871);
nand U46168 (N_46168,N_45858,N_45902);
nor U46169 (N_46169,N_45763,N_45906);
and U46170 (N_46170,N_45882,N_45840);
nor U46171 (N_46171,N_45974,N_45896);
xor U46172 (N_46172,N_45907,N_45910);
xor U46173 (N_46173,N_45886,N_45824);
xnor U46174 (N_46174,N_45914,N_45908);
or U46175 (N_46175,N_45964,N_45893);
nor U46176 (N_46176,N_45998,N_45936);
nor U46177 (N_46177,N_45894,N_45842);
nand U46178 (N_46178,N_45817,N_45756);
xnor U46179 (N_46179,N_45759,N_45764);
nor U46180 (N_46180,N_45762,N_45779);
xor U46181 (N_46181,N_45872,N_45840);
nand U46182 (N_46182,N_45886,N_45833);
nor U46183 (N_46183,N_45932,N_45800);
xnor U46184 (N_46184,N_45878,N_45753);
nor U46185 (N_46185,N_45939,N_45913);
nand U46186 (N_46186,N_45951,N_45868);
or U46187 (N_46187,N_45796,N_45837);
nand U46188 (N_46188,N_45981,N_45903);
nand U46189 (N_46189,N_45945,N_45827);
nand U46190 (N_46190,N_45752,N_45855);
xnor U46191 (N_46191,N_45771,N_45954);
nor U46192 (N_46192,N_45959,N_45991);
or U46193 (N_46193,N_45951,N_45913);
xor U46194 (N_46194,N_45858,N_45833);
nand U46195 (N_46195,N_45791,N_45853);
or U46196 (N_46196,N_45777,N_45784);
or U46197 (N_46197,N_45909,N_45851);
nor U46198 (N_46198,N_45967,N_45845);
xor U46199 (N_46199,N_45938,N_45787);
nand U46200 (N_46200,N_45886,N_45784);
and U46201 (N_46201,N_45901,N_45780);
or U46202 (N_46202,N_45862,N_45905);
xnor U46203 (N_46203,N_45981,N_45899);
and U46204 (N_46204,N_45921,N_45910);
and U46205 (N_46205,N_45789,N_45788);
or U46206 (N_46206,N_45764,N_45945);
nand U46207 (N_46207,N_45851,N_45773);
xnor U46208 (N_46208,N_45989,N_45886);
or U46209 (N_46209,N_45975,N_45824);
or U46210 (N_46210,N_45785,N_45948);
xnor U46211 (N_46211,N_45982,N_45966);
nor U46212 (N_46212,N_45976,N_45977);
and U46213 (N_46213,N_45824,N_45816);
or U46214 (N_46214,N_45798,N_45947);
xor U46215 (N_46215,N_45965,N_45890);
nand U46216 (N_46216,N_45800,N_45756);
and U46217 (N_46217,N_45923,N_45940);
xnor U46218 (N_46218,N_45942,N_45897);
nor U46219 (N_46219,N_45912,N_45963);
xor U46220 (N_46220,N_45927,N_45754);
nand U46221 (N_46221,N_45994,N_45996);
xor U46222 (N_46222,N_45815,N_45977);
nand U46223 (N_46223,N_45801,N_45799);
and U46224 (N_46224,N_45843,N_45991);
and U46225 (N_46225,N_45834,N_45891);
xor U46226 (N_46226,N_45860,N_45847);
nand U46227 (N_46227,N_45932,N_45831);
nor U46228 (N_46228,N_45756,N_45963);
or U46229 (N_46229,N_45943,N_45779);
nand U46230 (N_46230,N_45822,N_45913);
and U46231 (N_46231,N_45890,N_45855);
or U46232 (N_46232,N_45854,N_45815);
nor U46233 (N_46233,N_45957,N_45990);
nand U46234 (N_46234,N_45883,N_45840);
and U46235 (N_46235,N_45981,N_45781);
or U46236 (N_46236,N_45835,N_45897);
or U46237 (N_46237,N_45990,N_45817);
xnor U46238 (N_46238,N_45765,N_45793);
xor U46239 (N_46239,N_45905,N_45969);
or U46240 (N_46240,N_45763,N_45815);
nand U46241 (N_46241,N_45896,N_45842);
nand U46242 (N_46242,N_45888,N_45875);
and U46243 (N_46243,N_45871,N_45905);
nand U46244 (N_46244,N_45962,N_45783);
and U46245 (N_46245,N_45784,N_45824);
xnor U46246 (N_46246,N_45775,N_45853);
xnor U46247 (N_46247,N_45787,N_45782);
nor U46248 (N_46248,N_45979,N_45905);
xor U46249 (N_46249,N_45978,N_45967);
nor U46250 (N_46250,N_46061,N_46110);
nand U46251 (N_46251,N_46094,N_46066);
nor U46252 (N_46252,N_46068,N_46018);
nand U46253 (N_46253,N_46037,N_46085);
or U46254 (N_46254,N_46234,N_46141);
xnor U46255 (N_46255,N_46045,N_46025);
xor U46256 (N_46256,N_46000,N_46127);
nor U46257 (N_46257,N_46001,N_46034);
and U46258 (N_46258,N_46225,N_46239);
xor U46259 (N_46259,N_46184,N_46087);
or U46260 (N_46260,N_46121,N_46090);
or U46261 (N_46261,N_46003,N_46243);
nor U46262 (N_46262,N_46204,N_46229);
nand U46263 (N_46263,N_46168,N_46054);
and U46264 (N_46264,N_46048,N_46213);
xor U46265 (N_46265,N_46143,N_46084);
or U46266 (N_46266,N_46049,N_46091);
and U46267 (N_46267,N_46079,N_46189);
xnor U46268 (N_46268,N_46187,N_46010);
xor U46269 (N_46269,N_46019,N_46224);
nor U46270 (N_46270,N_46052,N_46044);
nand U46271 (N_46271,N_46013,N_46060);
and U46272 (N_46272,N_46152,N_46180);
nand U46273 (N_46273,N_46002,N_46161);
or U46274 (N_46274,N_46240,N_46073);
nor U46275 (N_46275,N_46122,N_46147);
nor U46276 (N_46276,N_46020,N_46162);
and U46277 (N_46277,N_46205,N_46065);
xnor U46278 (N_46278,N_46062,N_46132);
nor U46279 (N_46279,N_46177,N_46117);
or U46280 (N_46280,N_46153,N_46181);
or U46281 (N_46281,N_46179,N_46194);
or U46282 (N_46282,N_46157,N_46138);
and U46283 (N_46283,N_46191,N_46098);
or U46284 (N_46284,N_46118,N_46145);
nor U46285 (N_46285,N_46130,N_46160);
and U46286 (N_46286,N_46211,N_46072);
nand U46287 (N_46287,N_46057,N_46173);
and U46288 (N_46288,N_46102,N_46174);
or U46289 (N_46289,N_46111,N_46218);
or U46290 (N_46290,N_46030,N_46163);
nor U46291 (N_46291,N_46182,N_46144);
nor U46292 (N_46292,N_46176,N_46208);
xor U46293 (N_46293,N_46200,N_46217);
and U46294 (N_46294,N_46017,N_46185);
nand U46295 (N_46295,N_46101,N_46129);
nor U46296 (N_46296,N_46026,N_46228);
and U46297 (N_46297,N_46126,N_46146);
nor U46298 (N_46298,N_46159,N_46190);
and U46299 (N_46299,N_46096,N_46188);
nor U46300 (N_46300,N_46064,N_46199);
xnor U46301 (N_46301,N_46175,N_46036);
xnor U46302 (N_46302,N_46105,N_46056);
and U46303 (N_46303,N_46220,N_46095);
nor U46304 (N_46304,N_46137,N_46083);
nand U46305 (N_46305,N_46082,N_46043);
nor U46306 (N_46306,N_46133,N_46119);
or U46307 (N_46307,N_46023,N_46156);
nor U46308 (N_46308,N_46093,N_46123);
and U46309 (N_46309,N_46212,N_46046);
and U46310 (N_46310,N_46042,N_46109);
and U46311 (N_46311,N_46125,N_46216);
and U46312 (N_46312,N_46202,N_46136);
xor U46313 (N_46313,N_46222,N_46086);
nor U46314 (N_46314,N_46055,N_46230);
nor U46315 (N_46315,N_46214,N_46245);
and U46316 (N_46316,N_46032,N_46140);
nand U46317 (N_46317,N_46124,N_46027);
xor U46318 (N_46318,N_46165,N_46007);
nor U46319 (N_46319,N_46248,N_46235);
nand U46320 (N_46320,N_46081,N_46155);
nand U46321 (N_46321,N_46022,N_46024);
nor U46322 (N_46322,N_46195,N_46172);
nor U46323 (N_46323,N_46009,N_46120);
nand U46324 (N_46324,N_46236,N_46115);
nor U46325 (N_46325,N_46135,N_46150);
xnor U46326 (N_46326,N_46004,N_46131);
and U46327 (N_46327,N_46051,N_46231);
xor U46328 (N_46328,N_46186,N_46053);
or U46329 (N_46329,N_46154,N_46008);
and U46330 (N_46330,N_46192,N_46108);
xor U46331 (N_46331,N_46099,N_46067);
nand U46332 (N_46332,N_46233,N_46167);
xnor U46333 (N_46333,N_46171,N_46203);
nand U46334 (N_46334,N_46050,N_46005);
xor U46335 (N_46335,N_46219,N_46075);
or U46336 (N_46336,N_46031,N_46241);
nor U46337 (N_46337,N_46114,N_46232);
xnor U46338 (N_46338,N_46078,N_46242);
xor U46339 (N_46339,N_46104,N_46029);
or U46340 (N_46340,N_46151,N_46058);
or U46341 (N_46341,N_46198,N_46021);
and U46342 (N_46342,N_46201,N_46092);
or U46343 (N_46343,N_46100,N_46074);
xnor U46344 (N_46344,N_46196,N_46039);
and U46345 (N_46345,N_46209,N_46041);
and U46346 (N_46346,N_46089,N_46040);
xor U46347 (N_46347,N_46106,N_46069);
nor U46348 (N_46348,N_46016,N_46206);
xnor U46349 (N_46349,N_46227,N_46149);
nor U46350 (N_46350,N_46103,N_46088);
xnor U46351 (N_46351,N_46193,N_46197);
nand U46352 (N_46352,N_46047,N_46028);
nor U46353 (N_46353,N_46170,N_46221);
or U46354 (N_46354,N_46169,N_46166);
xor U46355 (N_46355,N_46063,N_46237);
and U46356 (N_46356,N_46015,N_46038);
xnor U46357 (N_46357,N_46178,N_46033);
xnor U46358 (N_46358,N_46011,N_46249);
xnor U46359 (N_46359,N_46070,N_46116);
or U46360 (N_46360,N_46148,N_46006);
nor U46361 (N_46361,N_46207,N_46210);
or U46362 (N_46362,N_46158,N_46014);
nor U46363 (N_46363,N_46080,N_46097);
xor U46364 (N_46364,N_46113,N_46226);
nor U46365 (N_46365,N_46134,N_46223);
xor U46366 (N_46366,N_46035,N_46247);
nor U46367 (N_46367,N_46139,N_46244);
or U46368 (N_46368,N_46238,N_46071);
xor U46369 (N_46369,N_46183,N_46215);
and U46370 (N_46370,N_46077,N_46012);
nor U46371 (N_46371,N_46164,N_46246);
nand U46372 (N_46372,N_46128,N_46112);
nor U46373 (N_46373,N_46107,N_46142);
nor U46374 (N_46374,N_46059,N_46076);
nor U46375 (N_46375,N_46233,N_46218);
xor U46376 (N_46376,N_46204,N_46003);
nand U46377 (N_46377,N_46202,N_46012);
nor U46378 (N_46378,N_46097,N_46098);
and U46379 (N_46379,N_46136,N_46090);
nand U46380 (N_46380,N_46179,N_46024);
nor U46381 (N_46381,N_46185,N_46022);
or U46382 (N_46382,N_46023,N_46123);
and U46383 (N_46383,N_46181,N_46033);
or U46384 (N_46384,N_46212,N_46197);
nand U46385 (N_46385,N_46137,N_46063);
nand U46386 (N_46386,N_46019,N_46057);
nor U46387 (N_46387,N_46027,N_46030);
xnor U46388 (N_46388,N_46206,N_46109);
or U46389 (N_46389,N_46140,N_46137);
nor U46390 (N_46390,N_46136,N_46074);
and U46391 (N_46391,N_46138,N_46113);
and U46392 (N_46392,N_46068,N_46057);
or U46393 (N_46393,N_46031,N_46197);
nor U46394 (N_46394,N_46203,N_46015);
nor U46395 (N_46395,N_46083,N_46225);
nand U46396 (N_46396,N_46147,N_46074);
and U46397 (N_46397,N_46125,N_46227);
and U46398 (N_46398,N_46059,N_46144);
nand U46399 (N_46399,N_46202,N_46086);
xnor U46400 (N_46400,N_46239,N_46132);
nor U46401 (N_46401,N_46037,N_46236);
xor U46402 (N_46402,N_46160,N_46223);
and U46403 (N_46403,N_46077,N_46245);
and U46404 (N_46404,N_46005,N_46186);
nor U46405 (N_46405,N_46105,N_46005);
nor U46406 (N_46406,N_46106,N_46167);
and U46407 (N_46407,N_46079,N_46172);
or U46408 (N_46408,N_46242,N_46001);
and U46409 (N_46409,N_46073,N_46173);
xor U46410 (N_46410,N_46095,N_46026);
nor U46411 (N_46411,N_46240,N_46157);
or U46412 (N_46412,N_46138,N_46024);
nor U46413 (N_46413,N_46236,N_46056);
nor U46414 (N_46414,N_46243,N_46154);
nand U46415 (N_46415,N_46232,N_46149);
or U46416 (N_46416,N_46151,N_46215);
nand U46417 (N_46417,N_46033,N_46247);
xor U46418 (N_46418,N_46096,N_46222);
or U46419 (N_46419,N_46208,N_46071);
nand U46420 (N_46420,N_46158,N_46079);
nand U46421 (N_46421,N_46171,N_46033);
or U46422 (N_46422,N_46015,N_46214);
xor U46423 (N_46423,N_46049,N_46223);
and U46424 (N_46424,N_46029,N_46102);
and U46425 (N_46425,N_46188,N_46121);
nor U46426 (N_46426,N_46192,N_46036);
nor U46427 (N_46427,N_46124,N_46164);
nor U46428 (N_46428,N_46054,N_46071);
and U46429 (N_46429,N_46241,N_46061);
nand U46430 (N_46430,N_46062,N_46164);
nor U46431 (N_46431,N_46229,N_46034);
nand U46432 (N_46432,N_46032,N_46121);
nor U46433 (N_46433,N_46141,N_46110);
nand U46434 (N_46434,N_46229,N_46094);
or U46435 (N_46435,N_46051,N_46149);
nand U46436 (N_46436,N_46031,N_46059);
nor U46437 (N_46437,N_46236,N_46023);
xor U46438 (N_46438,N_46197,N_46113);
and U46439 (N_46439,N_46036,N_46130);
or U46440 (N_46440,N_46101,N_46080);
or U46441 (N_46441,N_46247,N_46108);
nand U46442 (N_46442,N_46009,N_46051);
or U46443 (N_46443,N_46089,N_46244);
nor U46444 (N_46444,N_46203,N_46222);
or U46445 (N_46445,N_46200,N_46008);
or U46446 (N_46446,N_46020,N_46098);
nor U46447 (N_46447,N_46148,N_46159);
or U46448 (N_46448,N_46053,N_46076);
xor U46449 (N_46449,N_46155,N_46110);
or U46450 (N_46450,N_46095,N_46082);
or U46451 (N_46451,N_46158,N_46150);
and U46452 (N_46452,N_46131,N_46211);
or U46453 (N_46453,N_46189,N_46145);
nand U46454 (N_46454,N_46220,N_46185);
nor U46455 (N_46455,N_46232,N_46229);
xnor U46456 (N_46456,N_46213,N_46169);
and U46457 (N_46457,N_46055,N_46056);
and U46458 (N_46458,N_46223,N_46020);
xor U46459 (N_46459,N_46152,N_46197);
nor U46460 (N_46460,N_46096,N_46204);
and U46461 (N_46461,N_46086,N_46181);
xnor U46462 (N_46462,N_46175,N_46077);
xor U46463 (N_46463,N_46128,N_46085);
and U46464 (N_46464,N_46012,N_46118);
and U46465 (N_46465,N_46086,N_46034);
xnor U46466 (N_46466,N_46144,N_46109);
xor U46467 (N_46467,N_46071,N_46246);
or U46468 (N_46468,N_46128,N_46061);
or U46469 (N_46469,N_46091,N_46225);
and U46470 (N_46470,N_46093,N_46111);
xnor U46471 (N_46471,N_46145,N_46149);
nor U46472 (N_46472,N_46185,N_46033);
and U46473 (N_46473,N_46136,N_46131);
nand U46474 (N_46474,N_46004,N_46058);
xnor U46475 (N_46475,N_46087,N_46236);
and U46476 (N_46476,N_46215,N_46021);
nand U46477 (N_46477,N_46202,N_46163);
nor U46478 (N_46478,N_46116,N_46194);
or U46479 (N_46479,N_46246,N_46043);
xnor U46480 (N_46480,N_46102,N_46249);
and U46481 (N_46481,N_46239,N_46060);
or U46482 (N_46482,N_46066,N_46077);
nand U46483 (N_46483,N_46072,N_46185);
xor U46484 (N_46484,N_46233,N_46011);
and U46485 (N_46485,N_46214,N_46157);
or U46486 (N_46486,N_46083,N_46050);
or U46487 (N_46487,N_46178,N_46102);
nor U46488 (N_46488,N_46208,N_46084);
nor U46489 (N_46489,N_46059,N_46088);
nand U46490 (N_46490,N_46125,N_46128);
nand U46491 (N_46491,N_46207,N_46024);
nor U46492 (N_46492,N_46030,N_46152);
xnor U46493 (N_46493,N_46018,N_46035);
and U46494 (N_46494,N_46027,N_46182);
nor U46495 (N_46495,N_46049,N_46217);
nor U46496 (N_46496,N_46233,N_46178);
and U46497 (N_46497,N_46184,N_46202);
and U46498 (N_46498,N_46182,N_46011);
xor U46499 (N_46499,N_46219,N_46052);
and U46500 (N_46500,N_46429,N_46465);
nand U46501 (N_46501,N_46498,N_46410);
xnor U46502 (N_46502,N_46360,N_46334);
xnor U46503 (N_46503,N_46361,N_46304);
or U46504 (N_46504,N_46496,N_46457);
or U46505 (N_46505,N_46411,N_46466);
xnor U46506 (N_46506,N_46415,N_46341);
or U46507 (N_46507,N_46329,N_46495);
or U46508 (N_46508,N_46285,N_46374);
xor U46509 (N_46509,N_46264,N_46376);
or U46510 (N_46510,N_46395,N_46409);
or U46511 (N_46511,N_46354,N_46402);
xnor U46512 (N_46512,N_46363,N_46288);
or U46513 (N_46513,N_46451,N_46336);
nand U46514 (N_46514,N_46393,N_46293);
nand U46515 (N_46515,N_46487,N_46419);
nor U46516 (N_46516,N_46477,N_46428);
or U46517 (N_46517,N_46328,N_46353);
nand U46518 (N_46518,N_46407,N_46283);
nor U46519 (N_46519,N_46260,N_46417);
nor U46520 (N_46520,N_46269,N_46322);
nand U46521 (N_46521,N_46330,N_46326);
xor U46522 (N_46522,N_46434,N_46358);
xnor U46523 (N_46523,N_46398,N_46327);
nand U46524 (N_46524,N_46416,N_46379);
and U46525 (N_46525,N_46312,N_46406);
xnor U46526 (N_46526,N_46383,N_46473);
or U46527 (N_46527,N_46308,N_46297);
nand U46528 (N_46528,N_46386,N_46436);
and U46529 (N_46529,N_46381,N_46268);
and U46530 (N_46530,N_46408,N_46489);
nand U46531 (N_46531,N_46305,N_46342);
nand U46532 (N_46532,N_46266,N_46454);
or U46533 (N_46533,N_46366,N_46464);
nor U46534 (N_46534,N_46396,N_46413);
nor U46535 (N_46535,N_46338,N_46418);
nor U46536 (N_46536,N_46491,N_46332);
xnor U46537 (N_46537,N_46488,N_46340);
or U46538 (N_46538,N_46325,N_46291);
xor U46539 (N_46539,N_46346,N_46294);
nand U46540 (N_46540,N_46368,N_46401);
or U46541 (N_46541,N_46323,N_46314);
nor U46542 (N_46542,N_46492,N_46310);
nor U46543 (N_46543,N_46382,N_46482);
nor U46544 (N_46544,N_46320,N_46385);
or U46545 (N_46545,N_46319,N_46399);
nand U46546 (N_46546,N_46378,N_46420);
and U46547 (N_46547,N_46261,N_46271);
xnor U46548 (N_46548,N_46472,N_46371);
nor U46549 (N_46549,N_46459,N_46256);
or U46550 (N_46550,N_46315,N_46377);
nand U46551 (N_46551,N_46469,N_46425);
and U46552 (N_46552,N_46499,N_46391);
nor U46553 (N_46553,N_46474,N_46296);
nor U46554 (N_46554,N_46485,N_46276);
nand U46555 (N_46555,N_46370,N_46460);
or U46556 (N_46556,N_46448,N_46380);
nor U46557 (N_46557,N_46311,N_46337);
nor U46558 (N_46558,N_46307,N_46352);
or U46559 (N_46559,N_46470,N_46253);
nand U46560 (N_46560,N_46343,N_46445);
and U46561 (N_46561,N_46375,N_46287);
or U46562 (N_46562,N_46486,N_46412);
nor U46563 (N_46563,N_46278,N_46452);
nor U46564 (N_46564,N_46422,N_46316);
or U46565 (N_46565,N_46282,N_46279);
and U46566 (N_46566,N_46462,N_46455);
nand U46567 (N_46567,N_46481,N_46479);
nor U46568 (N_46568,N_46347,N_46397);
and U46569 (N_46569,N_46444,N_46387);
and U46570 (N_46570,N_46372,N_46456);
xnor U46571 (N_46571,N_46333,N_46480);
nand U46572 (N_46572,N_46438,N_46306);
nor U46573 (N_46573,N_46369,N_46257);
nand U46574 (N_46574,N_46476,N_46405);
and U46575 (N_46575,N_46389,N_46453);
nand U46576 (N_46576,N_46384,N_46403);
or U46577 (N_46577,N_46356,N_46439);
or U46578 (N_46578,N_46446,N_46289);
xnor U46579 (N_46579,N_46259,N_46345);
nand U46580 (N_46580,N_46440,N_46357);
and U46581 (N_46581,N_46394,N_46494);
or U46582 (N_46582,N_46478,N_46351);
xor U46583 (N_46583,N_46303,N_46295);
xor U46584 (N_46584,N_46251,N_46292);
nor U46585 (N_46585,N_46280,N_46490);
nand U46586 (N_46586,N_46335,N_46258);
xnor U46587 (N_46587,N_46267,N_46302);
or U46588 (N_46588,N_46367,N_46467);
nor U46589 (N_46589,N_46364,N_46450);
xnor U46590 (N_46590,N_46265,N_46350);
and U46591 (N_46591,N_46437,N_46252);
nand U46592 (N_46592,N_46468,N_46449);
and U46593 (N_46593,N_46263,N_46497);
nor U46594 (N_46594,N_46359,N_46426);
and U46595 (N_46595,N_46388,N_46349);
nor U46596 (N_46596,N_46484,N_46390);
and U46597 (N_46597,N_46281,N_46299);
xor U46598 (N_46598,N_46273,N_46493);
nor U46599 (N_46599,N_46321,N_46318);
xnor U46600 (N_46600,N_46461,N_46404);
xor U46601 (N_46601,N_46317,N_46301);
and U46602 (N_46602,N_46254,N_46421);
or U46603 (N_46603,N_46471,N_46284);
nand U46604 (N_46604,N_46442,N_46331);
nand U46605 (N_46605,N_46423,N_46339);
xnor U46606 (N_46606,N_46277,N_46443);
or U46607 (N_46607,N_46355,N_46324);
nor U46608 (N_46608,N_46365,N_46447);
and U46609 (N_46609,N_46373,N_46458);
nand U46610 (N_46610,N_46392,N_46250);
nor U46611 (N_46611,N_46431,N_46344);
xnor U46612 (N_46612,N_46262,N_46255);
nor U46613 (N_46613,N_46275,N_46427);
nor U46614 (N_46614,N_46298,N_46424);
xnor U46615 (N_46615,N_46313,N_46274);
nor U46616 (N_46616,N_46430,N_46414);
xor U46617 (N_46617,N_46463,N_46309);
or U46618 (N_46618,N_46483,N_46290);
and U46619 (N_46619,N_46400,N_46435);
or U46620 (N_46620,N_46432,N_46441);
nand U46621 (N_46621,N_46270,N_46286);
xor U46622 (N_46622,N_46348,N_46433);
or U46623 (N_46623,N_46362,N_46272);
and U46624 (N_46624,N_46300,N_46475);
or U46625 (N_46625,N_46359,N_46453);
or U46626 (N_46626,N_46293,N_46297);
and U46627 (N_46627,N_46268,N_46366);
xnor U46628 (N_46628,N_46398,N_46402);
and U46629 (N_46629,N_46382,N_46408);
and U46630 (N_46630,N_46257,N_46436);
or U46631 (N_46631,N_46411,N_46376);
nand U46632 (N_46632,N_46389,N_46492);
nor U46633 (N_46633,N_46317,N_46487);
nand U46634 (N_46634,N_46375,N_46472);
and U46635 (N_46635,N_46298,N_46350);
xor U46636 (N_46636,N_46475,N_46495);
nand U46637 (N_46637,N_46397,N_46325);
xor U46638 (N_46638,N_46337,N_46396);
xnor U46639 (N_46639,N_46357,N_46324);
nand U46640 (N_46640,N_46388,N_46442);
xnor U46641 (N_46641,N_46430,N_46425);
and U46642 (N_46642,N_46422,N_46475);
nand U46643 (N_46643,N_46410,N_46489);
xor U46644 (N_46644,N_46484,N_46318);
and U46645 (N_46645,N_46290,N_46446);
or U46646 (N_46646,N_46487,N_46376);
nand U46647 (N_46647,N_46478,N_46383);
and U46648 (N_46648,N_46400,N_46284);
and U46649 (N_46649,N_46321,N_46462);
nor U46650 (N_46650,N_46380,N_46481);
or U46651 (N_46651,N_46478,N_46448);
nand U46652 (N_46652,N_46390,N_46294);
nor U46653 (N_46653,N_46386,N_46416);
nand U46654 (N_46654,N_46271,N_46425);
or U46655 (N_46655,N_46486,N_46471);
xnor U46656 (N_46656,N_46492,N_46338);
nor U46657 (N_46657,N_46379,N_46397);
and U46658 (N_46658,N_46278,N_46297);
xor U46659 (N_46659,N_46388,N_46317);
nand U46660 (N_46660,N_46356,N_46456);
or U46661 (N_46661,N_46320,N_46293);
nand U46662 (N_46662,N_46383,N_46341);
nor U46663 (N_46663,N_46487,N_46337);
or U46664 (N_46664,N_46368,N_46252);
nor U46665 (N_46665,N_46430,N_46443);
and U46666 (N_46666,N_46381,N_46346);
nor U46667 (N_46667,N_46259,N_46359);
nor U46668 (N_46668,N_46394,N_46353);
nor U46669 (N_46669,N_46351,N_46474);
nor U46670 (N_46670,N_46482,N_46301);
nor U46671 (N_46671,N_46337,N_46481);
xor U46672 (N_46672,N_46403,N_46365);
and U46673 (N_46673,N_46438,N_46402);
nor U46674 (N_46674,N_46301,N_46321);
nor U46675 (N_46675,N_46480,N_46387);
and U46676 (N_46676,N_46332,N_46272);
or U46677 (N_46677,N_46428,N_46437);
or U46678 (N_46678,N_46495,N_46421);
nor U46679 (N_46679,N_46327,N_46286);
nand U46680 (N_46680,N_46344,N_46477);
nor U46681 (N_46681,N_46337,N_46467);
xor U46682 (N_46682,N_46281,N_46386);
or U46683 (N_46683,N_46304,N_46420);
and U46684 (N_46684,N_46333,N_46325);
nor U46685 (N_46685,N_46397,N_46388);
nand U46686 (N_46686,N_46301,N_46471);
or U46687 (N_46687,N_46409,N_46447);
nor U46688 (N_46688,N_46358,N_46314);
and U46689 (N_46689,N_46285,N_46308);
and U46690 (N_46690,N_46404,N_46293);
nand U46691 (N_46691,N_46428,N_46423);
nor U46692 (N_46692,N_46302,N_46273);
or U46693 (N_46693,N_46370,N_46376);
nor U46694 (N_46694,N_46426,N_46254);
nand U46695 (N_46695,N_46419,N_46409);
or U46696 (N_46696,N_46495,N_46274);
xnor U46697 (N_46697,N_46406,N_46415);
nand U46698 (N_46698,N_46397,N_46251);
nand U46699 (N_46699,N_46260,N_46269);
xor U46700 (N_46700,N_46365,N_46343);
xnor U46701 (N_46701,N_46391,N_46312);
and U46702 (N_46702,N_46306,N_46370);
or U46703 (N_46703,N_46386,N_46253);
nand U46704 (N_46704,N_46351,N_46266);
xnor U46705 (N_46705,N_46263,N_46352);
xnor U46706 (N_46706,N_46399,N_46292);
nor U46707 (N_46707,N_46396,N_46494);
or U46708 (N_46708,N_46293,N_46348);
and U46709 (N_46709,N_46258,N_46274);
and U46710 (N_46710,N_46369,N_46308);
nand U46711 (N_46711,N_46472,N_46260);
or U46712 (N_46712,N_46470,N_46344);
and U46713 (N_46713,N_46469,N_46266);
nor U46714 (N_46714,N_46498,N_46312);
nor U46715 (N_46715,N_46279,N_46434);
nand U46716 (N_46716,N_46411,N_46432);
nor U46717 (N_46717,N_46499,N_46297);
nand U46718 (N_46718,N_46295,N_46461);
nand U46719 (N_46719,N_46255,N_46462);
xnor U46720 (N_46720,N_46282,N_46259);
nor U46721 (N_46721,N_46446,N_46336);
nand U46722 (N_46722,N_46334,N_46443);
nor U46723 (N_46723,N_46288,N_46465);
and U46724 (N_46724,N_46470,N_46408);
xor U46725 (N_46725,N_46448,N_46497);
or U46726 (N_46726,N_46388,N_46262);
and U46727 (N_46727,N_46450,N_46446);
and U46728 (N_46728,N_46289,N_46469);
or U46729 (N_46729,N_46420,N_46414);
and U46730 (N_46730,N_46447,N_46372);
nand U46731 (N_46731,N_46346,N_46308);
and U46732 (N_46732,N_46393,N_46266);
xor U46733 (N_46733,N_46334,N_46363);
nand U46734 (N_46734,N_46340,N_46271);
and U46735 (N_46735,N_46420,N_46334);
or U46736 (N_46736,N_46315,N_46403);
and U46737 (N_46737,N_46420,N_46391);
nand U46738 (N_46738,N_46327,N_46321);
or U46739 (N_46739,N_46357,N_46497);
or U46740 (N_46740,N_46464,N_46272);
nor U46741 (N_46741,N_46405,N_46322);
nor U46742 (N_46742,N_46400,N_46260);
nor U46743 (N_46743,N_46495,N_46319);
or U46744 (N_46744,N_46329,N_46473);
nand U46745 (N_46745,N_46464,N_46372);
or U46746 (N_46746,N_46456,N_46399);
and U46747 (N_46747,N_46294,N_46399);
or U46748 (N_46748,N_46266,N_46441);
or U46749 (N_46749,N_46272,N_46343);
nor U46750 (N_46750,N_46540,N_46636);
nor U46751 (N_46751,N_46715,N_46727);
xor U46752 (N_46752,N_46654,N_46609);
nor U46753 (N_46753,N_46622,N_46619);
nor U46754 (N_46754,N_46680,N_46613);
and U46755 (N_46755,N_46561,N_46629);
or U46756 (N_46756,N_46749,N_46621);
nand U46757 (N_46757,N_46598,N_46604);
or U46758 (N_46758,N_46558,N_46548);
nand U46759 (N_46759,N_46515,N_46568);
nor U46760 (N_46760,N_46575,N_46646);
nor U46761 (N_46761,N_46579,N_46655);
xor U46762 (N_46762,N_46511,N_46625);
xor U46763 (N_46763,N_46701,N_46537);
xnor U46764 (N_46764,N_46617,N_46616);
xnor U46765 (N_46765,N_46664,N_46674);
nor U46766 (N_46766,N_46641,N_46581);
nor U46767 (N_46767,N_46662,N_46530);
or U46768 (N_46768,N_46531,N_46524);
xnor U46769 (N_46769,N_46670,N_46536);
and U46770 (N_46770,N_46620,N_46716);
nand U46771 (N_46771,N_46563,N_46572);
xor U46772 (N_46772,N_46696,N_46667);
or U46773 (N_46773,N_46506,N_46505);
and U46774 (N_46774,N_46585,N_46658);
xor U46775 (N_46775,N_46605,N_46736);
nand U46776 (N_46776,N_46692,N_46565);
xnor U46777 (N_46777,N_46747,N_46699);
nor U46778 (N_46778,N_46547,N_46597);
xnor U46779 (N_46779,N_46612,N_46669);
or U46780 (N_46780,N_46591,N_46666);
or U46781 (N_46781,N_46576,N_46726);
nand U46782 (N_46782,N_46649,N_46746);
nor U46783 (N_46783,N_46628,N_46732);
and U46784 (N_46784,N_46638,N_46551);
nand U46785 (N_46785,N_46714,N_46627);
xor U46786 (N_46786,N_46682,N_46508);
nor U46787 (N_46787,N_46721,N_46707);
nor U46788 (N_46788,N_46639,N_46539);
or U46789 (N_46789,N_46559,N_46644);
nor U46790 (N_46790,N_46672,N_46724);
or U46791 (N_46791,N_46740,N_46693);
and U46792 (N_46792,N_46648,N_46584);
xor U46793 (N_46793,N_46560,N_46719);
nor U46794 (N_46794,N_46510,N_46618);
or U46795 (N_46795,N_46587,N_46643);
and U46796 (N_46796,N_46683,N_46574);
or U46797 (N_46797,N_46708,N_46642);
nor U46798 (N_46798,N_46668,N_46728);
nor U46799 (N_46799,N_46634,N_46653);
and U46800 (N_46800,N_46573,N_46562);
nand U46801 (N_46801,N_46599,N_46671);
xor U46802 (N_46802,N_46734,N_46608);
or U46803 (N_46803,N_46723,N_46606);
xnor U46804 (N_46804,N_46645,N_46571);
or U46805 (N_46805,N_46543,N_46514);
and U46806 (N_46806,N_46545,N_46603);
xnor U46807 (N_46807,N_46748,N_46718);
nand U46808 (N_46808,N_46615,N_46731);
nand U46809 (N_46809,N_46556,N_46651);
nor U46810 (N_46810,N_46677,N_46730);
xnor U46811 (N_46811,N_46709,N_46700);
or U46812 (N_46812,N_46712,N_46513);
or U46813 (N_46813,N_46503,N_46583);
xnor U46814 (N_46814,N_46741,N_46702);
nor U46815 (N_46815,N_46637,N_46555);
xnor U46816 (N_46816,N_46713,N_46656);
nor U46817 (N_46817,N_46659,N_46652);
or U46818 (N_46818,N_46532,N_46742);
and U46819 (N_46819,N_46553,N_46518);
and U46820 (N_46820,N_46594,N_46527);
or U46821 (N_46821,N_46690,N_46733);
nor U46822 (N_46822,N_46665,N_46504);
or U46823 (N_46823,N_46661,N_46717);
and U46824 (N_46824,N_46509,N_46507);
xor U46825 (N_46825,N_46737,N_46704);
xor U46826 (N_46826,N_46688,N_46600);
nand U46827 (N_46827,N_46577,N_46590);
and U46828 (N_46828,N_46694,N_46650);
nor U46829 (N_46829,N_46678,N_46624);
or U46830 (N_46830,N_46541,N_46578);
or U46831 (N_46831,N_46517,N_46711);
nor U46832 (N_46832,N_46729,N_46550);
or U46833 (N_46833,N_46695,N_46533);
or U46834 (N_46834,N_46601,N_46607);
nor U46835 (N_46835,N_46687,N_46534);
nor U46836 (N_46836,N_46679,N_46725);
nand U46837 (N_46837,N_46595,N_46640);
nand U46838 (N_46838,N_46739,N_46697);
nand U46839 (N_46839,N_46720,N_46520);
and U46840 (N_46840,N_46567,N_46744);
and U46841 (N_46841,N_46554,N_46611);
nor U46842 (N_46842,N_46544,N_46516);
nor U46843 (N_46843,N_46525,N_46586);
or U46844 (N_46844,N_46675,N_46522);
or U46845 (N_46845,N_46592,N_46582);
xor U46846 (N_46846,N_46569,N_46738);
or U46847 (N_46847,N_46500,N_46542);
nor U46848 (N_46848,N_46593,N_46689);
xor U46849 (N_46849,N_46676,N_46686);
xnor U46850 (N_46850,N_46546,N_46663);
or U46851 (N_46851,N_46703,N_46626);
nor U46852 (N_46852,N_46528,N_46529);
xor U46853 (N_46853,N_46589,N_46631);
or U46854 (N_46854,N_46580,N_46557);
nor U46855 (N_46855,N_46632,N_46521);
or U46856 (N_46856,N_46710,N_46630);
and U46857 (N_46857,N_46633,N_46566);
nor U46858 (N_46858,N_46523,N_46745);
xor U46859 (N_46859,N_46623,N_46681);
and U46860 (N_46860,N_46588,N_46564);
nand U46861 (N_46861,N_46549,N_46635);
and U46862 (N_46862,N_46519,N_46691);
or U46863 (N_46863,N_46657,N_46647);
nor U46864 (N_46864,N_46535,N_46684);
and U46865 (N_46865,N_46596,N_46501);
xnor U46866 (N_46866,N_46743,N_46526);
or U46867 (N_46867,N_46735,N_46685);
nand U46868 (N_46868,N_46698,N_46706);
or U46869 (N_46869,N_46512,N_46673);
nor U46870 (N_46870,N_46538,N_46722);
and U46871 (N_46871,N_46705,N_46614);
or U46872 (N_46872,N_46660,N_46570);
nand U46873 (N_46873,N_46602,N_46502);
and U46874 (N_46874,N_46552,N_46610);
nor U46875 (N_46875,N_46679,N_46650);
nand U46876 (N_46876,N_46559,N_46739);
nor U46877 (N_46877,N_46531,N_46652);
xnor U46878 (N_46878,N_46582,N_46641);
nor U46879 (N_46879,N_46558,N_46501);
or U46880 (N_46880,N_46706,N_46582);
and U46881 (N_46881,N_46636,N_46694);
xor U46882 (N_46882,N_46670,N_46514);
xnor U46883 (N_46883,N_46501,N_46719);
or U46884 (N_46884,N_46654,N_46610);
nand U46885 (N_46885,N_46730,N_46609);
nor U46886 (N_46886,N_46604,N_46621);
or U46887 (N_46887,N_46677,N_46644);
and U46888 (N_46888,N_46617,N_46567);
or U46889 (N_46889,N_46542,N_46525);
and U46890 (N_46890,N_46553,N_46505);
nor U46891 (N_46891,N_46692,N_46629);
nor U46892 (N_46892,N_46566,N_46725);
or U46893 (N_46893,N_46746,N_46735);
xnor U46894 (N_46894,N_46584,N_46718);
and U46895 (N_46895,N_46613,N_46592);
nand U46896 (N_46896,N_46544,N_46746);
and U46897 (N_46897,N_46523,N_46573);
nand U46898 (N_46898,N_46686,N_46721);
nand U46899 (N_46899,N_46677,N_46617);
nor U46900 (N_46900,N_46582,N_46716);
or U46901 (N_46901,N_46670,N_46618);
nor U46902 (N_46902,N_46691,N_46556);
nor U46903 (N_46903,N_46576,N_46512);
nand U46904 (N_46904,N_46556,N_46540);
or U46905 (N_46905,N_46545,N_46563);
nor U46906 (N_46906,N_46700,N_46663);
nor U46907 (N_46907,N_46599,N_46743);
and U46908 (N_46908,N_46711,N_46645);
xor U46909 (N_46909,N_46725,N_46634);
nand U46910 (N_46910,N_46697,N_46628);
nor U46911 (N_46911,N_46688,N_46531);
nand U46912 (N_46912,N_46729,N_46534);
or U46913 (N_46913,N_46592,N_46720);
nor U46914 (N_46914,N_46658,N_46603);
nand U46915 (N_46915,N_46721,N_46724);
nand U46916 (N_46916,N_46707,N_46658);
or U46917 (N_46917,N_46656,N_46608);
or U46918 (N_46918,N_46710,N_46732);
or U46919 (N_46919,N_46543,N_46518);
nand U46920 (N_46920,N_46505,N_46581);
xor U46921 (N_46921,N_46664,N_46576);
or U46922 (N_46922,N_46603,N_46624);
and U46923 (N_46923,N_46570,N_46649);
or U46924 (N_46924,N_46631,N_46692);
nor U46925 (N_46925,N_46510,N_46580);
and U46926 (N_46926,N_46598,N_46526);
xnor U46927 (N_46927,N_46714,N_46607);
xnor U46928 (N_46928,N_46718,N_46568);
nand U46929 (N_46929,N_46667,N_46613);
and U46930 (N_46930,N_46623,N_46565);
nand U46931 (N_46931,N_46599,N_46619);
xnor U46932 (N_46932,N_46630,N_46695);
nand U46933 (N_46933,N_46640,N_46691);
nand U46934 (N_46934,N_46708,N_46598);
or U46935 (N_46935,N_46674,N_46584);
and U46936 (N_46936,N_46693,N_46650);
or U46937 (N_46937,N_46729,N_46507);
nand U46938 (N_46938,N_46629,N_46691);
or U46939 (N_46939,N_46719,N_46744);
xor U46940 (N_46940,N_46748,N_46704);
xor U46941 (N_46941,N_46679,N_46602);
nand U46942 (N_46942,N_46598,N_46745);
xnor U46943 (N_46943,N_46740,N_46562);
and U46944 (N_46944,N_46733,N_46669);
xor U46945 (N_46945,N_46568,N_46669);
nor U46946 (N_46946,N_46665,N_46724);
and U46947 (N_46947,N_46590,N_46586);
nor U46948 (N_46948,N_46582,N_46512);
xor U46949 (N_46949,N_46648,N_46741);
nor U46950 (N_46950,N_46698,N_46636);
and U46951 (N_46951,N_46580,N_46586);
nor U46952 (N_46952,N_46526,N_46661);
nand U46953 (N_46953,N_46608,N_46593);
nand U46954 (N_46954,N_46624,N_46512);
and U46955 (N_46955,N_46653,N_46717);
nand U46956 (N_46956,N_46607,N_46506);
or U46957 (N_46957,N_46562,N_46554);
nand U46958 (N_46958,N_46511,N_46681);
nor U46959 (N_46959,N_46569,N_46667);
or U46960 (N_46960,N_46692,N_46606);
and U46961 (N_46961,N_46652,N_46525);
nand U46962 (N_46962,N_46570,N_46538);
nand U46963 (N_46963,N_46636,N_46651);
or U46964 (N_46964,N_46719,N_46676);
xor U46965 (N_46965,N_46684,N_46736);
and U46966 (N_46966,N_46715,N_46599);
xor U46967 (N_46967,N_46695,N_46651);
and U46968 (N_46968,N_46639,N_46690);
xnor U46969 (N_46969,N_46656,N_46518);
nor U46970 (N_46970,N_46582,N_46568);
nor U46971 (N_46971,N_46726,N_46659);
nand U46972 (N_46972,N_46639,N_46688);
nand U46973 (N_46973,N_46619,N_46660);
or U46974 (N_46974,N_46726,N_46645);
xnor U46975 (N_46975,N_46562,N_46698);
nand U46976 (N_46976,N_46705,N_46621);
nor U46977 (N_46977,N_46742,N_46724);
or U46978 (N_46978,N_46741,N_46742);
nand U46979 (N_46979,N_46636,N_46634);
and U46980 (N_46980,N_46555,N_46681);
nor U46981 (N_46981,N_46599,N_46647);
nor U46982 (N_46982,N_46746,N_46572);
nor U46983 (N_46983,N_46594,N_46618);
nand U46984 (N_46984,N_46735,N_46520);
xor U46985 (N_46985,N_46501,N_46539);
or U46986 (N_46986,N_46579,N_46546);
nor U46987 (N_46987,N_46555,N_46624);
nor U46988 (N_46988,N_46623,N_46581);
and U46989 (N_46989,N_46693,N_46598);
nor U46990 (N_46990,N_46736,N_46677);
or U46991 (N_46991,N_46519,N_46554);
or U46992 (N_46992,N_46538,N_46587);
and U46993 (N_46993,N_46658,N_46625);
nor U46994 (N_46994,N_46621,N_46567);
nor U46995 (N_46995,N_46618,N_46533);
and U46996 (N_46996,N_46582,N_46573);
or U46997 (N_46997,N_46620,N_46580);
xnor U46998 (N_46998,N_46733,N_46619);
xnor U46999 (N_46999,N_46606,N_46704);
nand U47000 (N_47000,N_46906,N_46915);
and U47001 (N_47001,N_46754,N_46821);
nor U47002 (N_47002,N_46984,N_46833);
and U47003 (N_47003,N_46830,N_46903);
or U47004 (N_47004,N_46989,N_46755);
nor U47005 (N_47005,N_46796,N_46857);
nand U47006 (N_47006,N_46949,N_46855);
or U47007 (N_47007,N_46874,N_46935);
nand U47008 (N_47008,N_46832,N_46768);
nor U47009 (N_47009,N_46823,N_46788);
nand U47010 (N_47010,N_46801,N_46946);
and U47011 (N_47011,N_46793,N_46907);
xnor U47012 (N_47012,N_46815,N_46846);
nor U47013 (N_47013,N_46980,N_46879);
nor U47014 (N_47014,N_46818,N_46831);
nand U47015 (N_47015,N_46763,N_46923);
nor U47016 (N_47016,N_46953,N_46994);
nor U47017 (N_47017,N_46863,N_46985);
nor U47018 (N_47018,N_46890,N_46804);
and U47019 (N_47019,N_46967,N_46955);
or U47020 (N_47020,N_46940,N_46993);
nand U47021 (N_47021,N_46780,N_46848);
nand U47022 (N_47022,N_46811,N_46800);
xor U47023 (N_47023,N_46850,N_46892);
and U47024 (N_47024,N_46789,N_46996);
and U47025 (N_47025,N_46834,N_46901);
and U47026 (N_47026,N_46962,N_46939);
nor U47027 (N_47027,N_46774,N_46757);
and U47028 (N_47028,N_46767,N_46979);
xnor U47029 (N_47029,N_46816,N_46988);
and U47030 (N_47030,N_46961,N_46797);
xor U47031 (N_47031,N_46924,N_46778);
nand U47032 (N_47032,N_46758,N_46752);
or U47033 (N_47033,N_46847,N_46875);
and U47034 (N_47034,N_46813,N_46838);
nand U47035 (N_47035,N_46826,N_46934);
or U47036 (N_47036,N_46889,N_46992);
xnor U47037 (N_47037,N_46837,N_46897);
nor U47038 (N_47038,N_46779,N_46808);
nand U47039 (N_47039,N_46922,N_46877);
nor U47040 (N_47040,N_46963,N_46771);
nor U47041 (N_47041,N_46756,N_46978);
xnor U47042 (N_47042,N_46829,N_46944);
nor U47043 (N_47043,N_46870,N_46910);
and U47044 (N_47044,N_46853,N_46881);
xnor U47045 (N_47045,N_46769,N_46931);
or U47046 (N_47046,N_46927,N_46895);
or U47047 (N_47047,N_46845,N_46941);
nor U47048 (N_47048,N_46835,N_46840);
nor U47049 (N_47049,N_46882,N_46957);
xnor U47050 (N_47050,N_46990,N_46803);
nor U47051 (N_47051,N_46849,N_46921);
or U47052 (N_47052,N_46969,N_46886);
nor U47053 (N_47053,N_46760,N_46973);
nand U47054 (N_47054,N_46759,N_46937);
nand U47055 (N_47055,N_46820,N_46805);
and U47056 (N_47056,N_46861,N_46948);
xor U47057 (N_47057,N_46960,N_46983);
nand U47058 (N_47058,N_46851,N_46887);
nand U47059 (N_47059,N_46764,N_46807);
and U47060 (N_47060,N_46824,N_46928);
nand U47061 (N_47061,N_46856,N_46860);
or U47062 (N_47062,N_46958,N_46896);
xnor U47063 (N_47063,N_46867,N_46753);
or U47064 (N_47064,N_46884,N_46812);
and U47065 (N_47065,N_46792,N_46844);
or U47066 (N_47066,N_46914,N_46864);
xnor U47067 (N_47067,N_46965,N_46950);
or U47068 (N_47068,N_46968,N_46970);
xnor U47069 (N_47069,N_46770,N_46975);
nor U47070 (N_47070,N_46972,N_46932);
or U47071 (N_47071,N_46902,N_46819);
or U47072 (N_47072,N_46827,N_46795);
nand U47073 (N_47073,N_46951,N_46974);
xor U47074 (N_47074,N_46883,N_46933);
or U47075 (N_47075,N_46791,N_46995);
and U47076 (N_47076,N_46899,N_46912);
or U47077 (N_47077,N_46817,N_46894);
and U47078 (N_47078,N_46904,N_46885);
nor U47079 (N_47079,N_46891,N_46913);
or U47080 (N_47080,N_46859,N_46880);
nor U47081 (N_47081,N_46783,N_46872);
or U47082 (N_47082,N_46828,N_46761);
xor U47083 (N_47083,N_46938,N_46772);
and U47084 (N_47084,N_46936,N_46929);
and U47085 (N_47085,N_46987,N_46842);
nand U47086 (N_47086,N_46911,N_46858);
or U47087 (N_47087,N_46750,N_46919);
or U47088 (N_47088,N_46776,N_46836);
xnor U47089 (N_47089,N_46809,N_46998);
xnor U47090 (N_47090,N_46982,N_46873);
nor U47091 (N_47091,N_46917,N_46773);
nand U47092 (N_47092,N_46777,N_46841);
or U47093 (N_47093,N_46930,N_46916);
xnor U47094 (N_47094,N_46839,N_46966);
nor U47095 (N_47095,N_46942,N_46888);
or U47096 (N_47096,N_46810,N_46806);
nand U47097 (N_47097,N_46964,N_46997);
or U47098 (N_47098,N_46865,N_46814);
nor U47099 (N_47099,N_46876,N_46900);
and U47100 (N_47100,N_46898,N_46751);
or U47101 (N_47101,N_46871,N_46794);
nand U47102 (N_47102,N_46775,N_46799);
nor U47103 (N_47103,N_46765,N_46976);
nor U47104 (N_47104,N_46787,N_46868);
xor U47105 (N_47105,N_46918,N_46766);
nand U47106 (N_47106,N_46905,N_46908);
nand U47107 (N_47107,N_46999,N_46986);
nand U47108 (N_47108,N_46825,N_46786);
and U47109 (N_47109,N_46843,N_46959);
nand U47110 (N_47110,N_46945,N_46854);
and U47111 (N_47111,N_46947,N_46981);
and U47112 (N_47112,N_46762,N_46971);
or U47113 (N_47113,N_46954,N_46952);
nand U47114 (N_47114,N_46943,N_46862);
and U47115 (N_47115,N_46909,N_46822);
xnor U47116 (N_47116,N_46869,N_46781);
or U47117 (N_47117,N_46802,N_46991);
nor U47118 (N_47118,N_46893,N_46866);
or U47119 (N_47119,N_46925,N_46977);
xnor U47120 (N_47120,N_46956,N_46782);
xor U47121 (N_47121,N_46878,N_46920);
or U47122 (N_47122,N_46785,N_46784);
nand U47123 (N_47123,N_46798,N_46852);
xor U47124 (N_47124,N_46790,N_46926);
xor U47125 (N_47125,N_46991,N_46858);
nand U47126 (N_47126,N_46802,N_46961);
xnor U47127 (N_47127,N_46988,N_46936);
xor U47128 (N_47128,N_46874,N_46789);
xnor U47129 (N_47129,N_46753,N_46926);
and U47130 (N_47130,N_46833,N_46790);
and U47131 (N_47131,N_46996,N_46750);
xor U47132 (N_47132,N_46884,N_46975);
nand U47133 (N_47133,N_46800,N_46843);
nor U47134 (N_47134,N_46816,N_46789);
or U47135 (N_47135,N_46841,N_46916);
nand U47136 (N_47136,N_46906,N_46893);
and U47137 (N_47137,N_46911,N_46933);
xor U47138 (N_47138,N_46898,N_46939);
nor U47139 (N_47139,N_46963,N_46751);
nor U47140 (N_47140,N_46795,N_46778);
nor U47141 (N_47141,N_46807,N_46941);
and U47142 (N_47142,N_46970,N_46935);
or U47143 (N_47143,N_46918,N_46839);
nand U47144 (N_47144,N_46929,N_46782);
or U47145 (N_47145,N_46832,N_46837);
and U47146 (N_47146,N_46958,N_46862);
xor U47147 (N_47147,N_46940,N_46768);
nor U47148 (N_47148,N_46752,N_46877);
nand U47149 (N_47149,N_46886,N_46917);
nand U47150 (N_47150,N_46836,N_46898);
and U47151 (N_47151,N_46922,N_46910);
xnor U47152 (N_47152,N_46865,N_46843);
xnor U47153 (N_47153,N_46851,N_46879);
and U47154 (N_47154,N_46937,N_46816);
nor U47155 (N_47155,N_46770,N_46868);
nor U47156 (N_47156,N_46919,N_46904);
xnor U47157 (N_47157,N_46963,N_46790);
or U47158 (N_47158,N_46757,N_46985);
nand U47159 (N_47159,N_46933,N_46839);
and U47160 (N_47160,N_46896,N_46932);
nand U47161 (N_47161,N_46841,N_46786);
nor U47162 (N_47162,N_46868,N_46996);
nand U47163 (N_47163,N_46955,N_46975);
xnor U47164 (N_47164,N_46785,N_46790);
nor U47165 (N_47165,N_46966,N_46994);
xnor U47166 (N_47166,N_46819,N_46941);
nor U47167 (N_47167,N_46850,N_46969);
or U47168 (N_47168,N_46943,N_46955);
xor U47169 (N_47169,N_46918,N_46958);
nand U47170 (N_47170,N_46850,N_46911);
nor U47171 (N_47171,N_46781,N_46806);
and U47172 (N_47172,N_46789,N_46917);
and U47173 (N_47173,N_46776,N_46975);
and U47174 (N_47174,N_46949,N_46877);
nand U47175 (N_47175,N_46834,N_46991);
xor U47176 (N_47176,N_46799,N_46872);
xnor U47177 (N_47177,N_46787,N_46977);
and U47178 (N_47178,N_46773,N_46775);
nor U47179 (N_47179,N_46852,N_46824);
nor U47180 (N_47180,N_46864,N_46807);
or U47181 (N_47181,N_46868,N_46762);
and U47182 (N_47182,N_46891,N_46922);
xor U47183 (N_47183,N_46874,N_46758);
or U47184 (N_47184,N_46842,N_46780);
or U47185 (N_47185,N_46883,N_46988);
nor U47186 (N_47186,N_46795,N_46772);
or U47187 (N_47187,N_46945,N_46850);
and U47188 (N_47188,N_46871,N_46926);
and U47189 (N_47189,N_46919,N_46934);
and U47190 (N_47190,N_46961,N_46838);
nand U47191 (N_47191,N_46858,N_46815);
xor U47192 (N_47192,N_46786,N_46902);
xor U47193 (N_47193,N_46814,N_46844);
nand U47194 (N_47194,N_46844,N_46769);
or U47195 (N_47195,N_46751,N_46917);
and U47196 (N_47196,N_46867,N_46761);
and U47197 (N_47197,N_46777,N_46769);
nand U47198 (N_47198,N_46784,N_46880);
xnor U47199 (N_47199,N_46959,N_46955);
nand U47200 (N_47200,N_46949,N_46900);
xnor U47201 (N_47201,N_46887,N_46931);
and U47202 (N_47202,N_46788,N_46981);
xor U47203 (N_47203,N_46950,N_46806);
and U47204 (N_47204,N_46987,N_46994);
nor U47205 (N_47205,N_46832,N_46796);
nor U47206 (N_47206,N_46943,N_46917);
nand U47207 (N_47207,N_46785,N_46982);
or U47208 (N_47208,N_46785,N_46913);
and U47209 (N_47209,N_46907,N_46767);
nor U47210 (N_47210,N_46856,N_46886);
and U47211 (N_47211,N_46799,N_46804);
nor U47212 (N_47212,N_46865,N_46944);
xor U47213 (N_47213,N_46938,N_46866);
or U47214 (N_47214,N_46919,N_46972);
nor U47215 (N_47215,N_46753,N_46967);
or U47216 (N_47216,N_46936,N_46831);
and U47217 (N_47217,N_46776,N_46838);
xor U47218 (N_47218,N_46865,N_46848);
or U47219 (N_47219,N_46779,N_46906);
nand U47220 (N_47220,N_46862,N_46857);
and U47221 (N_47221,N_46863,N_46960);
nand U47222 (N_47222,N_46939,N_46864);
and U47223 (N_47223,N_46761,N_46785);
xnor U47224 (N_47224,N_46772,N_46915);
and U47225 (N_47225,N_46783,N_46988);
and U47226 (N_47226,N_46976,N_46925);
nor U47227 (N_47227,N_46976,N_46763);
xor U47228 (N_47228,N_46802,N_46943);
nor U47229 (N_47229,N_46853,N_46830);
xnor U47230 (N_47230,N_46953,N_46917);
or U47231 (N_47231,N_46939,N_46953);
xnor U47232 (N_47232,N_46977,N_46914);
nand U47233 (N_47233,N_46922,N_46991);
nand U47234 (N_47234,N_46792,N_46752);
nand U47235 (N_47235,N_46796,N_46960);
nand U47236 (N_47236,N_46919,N_46812);
xor U47237 (N_47237,N_46908,N_46856);
and U47238 (N_47238,N_46842,N_46832);
nand U47239 (N_47239,N_46887,N_46946);
nand U47240 (N_47240,N_46758,N_46767);
nand U47241 (N_47241,N_46959,N_46769);
and U47242 (N_47242,N_46934,N_46939);
nand U47243 (N_47243,N_46966,N_46950);
and U47244 (N_47244,N_46942,N_46752);
xor U47245 (N_47245,N_46966,N_46986);
and U47246 (N_47246,N_46983,N_46859);
nand U47247 (N_47247,N_46837,N_46885);
xor U47248 (N_47248,N_46782,N_46799);
and U47249 (N_47249,N_46894,N_46776);
or U47250 (N_47250,N_47067,N_47049);
nand U47251 (N_47251,N_47144,N_47219);
or U47252 (N_47252,N_47040,N_47082);
nor U47253 (N_47253,N_47051,N_47202);
or U47254 (N_47254,N_47118,N_47187);
and U47255 (N_47255,N_47087,N_47193);
nand U47256 (N_47256,N_47150,N_47146);
and U47257 (N_47257,N_47047,N_47085);
xnor U47258 (N_47258,N_47230,N_47141);
or U47259 (N_47259,N_47209,N_47083);
nand U47260 (N_47260,N_47204,N_47052);
xor U47261 (N_47261,N_47149,N_47200);
and U47262 (N_47262,N_47115,N_47017);
xnor U47263 (N_47263,N_47130,N_47246);
or U47264 (N_47264,N_47211,N_47007);
nand U47265 (N_47265,N_47030,N_47080);
or U47266 (N_47266,N_47213,N_47244);
nor U47267 (N_47267,N_47164,N_47172);
or U47268 (N_47268,N_47233,N_47046);
or U47269 (N_47269,N_47135,N_47038);
xnor U47270 (N_47270,N_47162,N_47026);
nor U47271 (N_47271,N_47196,N_47055);
or U47272 (N_47272,N_47020,N_47088);
or U47273 (N_47273,N_47116,N_47237);
or U47274 (N_47274,N_47003,N_47195);
nor U47275 (N_47275,N_47142,N_47104);
and U47276 (N_47276,N_47097,N_47053);
xor U47277 (N_47277,N_47064,N_47176);
nor U47278 (N_47278,N_47159,N_47245);
nor U47279 (N_47279,N_47073,N_47199);
nand U47280 (N_47280,N_47101,N_47133);
and U47281 (N_47281,N_47121,N_47173);
or U47282 (N_47282,N_47190,N_47109);
or U47283 (N_47283,N_47151,N_47189);
xor U47284 (N_47284,N_47216,N_47100);
and U47285 (N_47285,N_47113,N_47015);
xnor U47286 (N_47286,N_47169,N_47134);
or U47287 (N_47287,N_47210,N_47156);
or U47288 (N_47288,N_47110,N_47090);
xnor U47289 (N_47289,N_47066,N_47241);
nand U47290 (N_47290,N_47005,N_47132);
xnor U47291 (N_47291,N_47065,N_47112);
nand U47292 (N_47292,N_47039,N_47054);
xor U47293 (N_47293,N_47106,N_47183);
or U47294 (N_47294,N_47179,N_47035);
or U47295 (N_47295,N_47212,N_47084);
and U47296 (N_47296,N_47036,N_47182);
or U47297 (N_47297,N_47057,N_47102);
nor U47298 (N_47298,N_47229,N_47208);
nand U47299 (N_47299,N_47016,N_47238);
and U47300 (N_47300,N_47075,N_47062);
nand U47301 (N_47301,N_47158,N_47068);
nand U47302 (N_47302,N_47095,N_47143);
or U47303 (N_47303,N_47091,N_47032);
xnor U47304 (N_47304,N_47019,N_47050);
and U47305 (N_47305,N_47081,N_47247);
xor U47306 (N_47306,N_47166,N_47221);
xnor U47307 (N_47307,N_47181,N_47157);
nor U47308 (N_47308,N_47044,N_47224);
nor U47309 (N_47309,N_47000,N_47077);
nand U47310 (N_47310,N_47098,N_47206);
xor U47311 (N_47311,N_47027,N_47155);
and U47312 (N_47312,N_47009,N_47160);
xnor U47313 (N_47313,N_47072,N_47093);
nand U47314 (N_47314,N_47174,N_47033);
nand U47315 (N_47315,N_47177,N_47226);
nand U47316 (N_47316,N_47028,N_47041);
or U47317 (N_47317,N_47243,N_47010);
nand U47318 (N_47318,N_47127,N_47071);
or U47319 (N_47319,N_47004,N_47048);
or U47320 (N_47320,N_47096,N_47001);
nor U47321 (N_47321,N_47188,N_47167);
nor U47322 (N_47322,N_47214,N_47205);
xnor U47323 (N_47323,N_47207,N_47171);
nor U47324 (N_47324,N_47234,N_47013);
xnor U47325 (N_47325,N_47043,N_47203);
nor U47326 (N_47326,N_47056,N_47140);
and U47327 (N_47327,N_47006,N_47008);
and U47328 (N_47328,N_47059,N_47147);
and U47329 (N_47329,N_47227,N_47185);
or U47330 (N_47330,N_47022,N_47076);
nand U47331 (N_47331,N_47126,N_47103);
nand U47332 (N_47332,N_47105,N_47011);
and U47333 (N_47333,N_47094,N_47045);
nor U47334 (N_47334,N_47037,N_47058);
xnor U47335 (N_47335,N_47218,N_47069);
xor U47336 (N_47336,N_47184,N_47031);
and U47337 (N_47337,N_47239,N_47201);
nand U47338 (N_47338,N_47024,N_47197);
xnor U47339 (N_47339,N_47078,N_47192);
and U47340 (N_47340,N_47136,N_47242);
xnor U47341 (N_47341,N_47119,N_47099);
xnor U47342 (N_47342,N_47152,N_47021);
and U47343 (N_47343,N_47225,N_47180);
or U47344 (N_47344,N_47215,N_47042);
nand U47345 (N_47345,N_47198,N_47074);
nand U47346 (N_47346,N_47232,N_47079);
and U47347 (N_47347,N_47236,N_47148);
nand U47348 (N_47348,N_47153,N_47018);
nor U47349 (N_47349,N_47168,N_47108);
nor U47350 (N_47350,N_47002,N_47154);
xnor U47351 (N_47351,N_47235,N_47139);
nand U47352 (N_47352,N_47114,N_47060);
nor U47353 (N_47353,N_47240,N_47170);
xor U47354 (N_47354,N_47249,N_47029);
and U47355 (N_47355,N_47186,N_47117);
or U47356 (N_47356,N_47231,N_47138);
nor U47357 (N_47357,N_47161,N_47128);
or U47358 (N_47358,N_47086,N_47063);
or U47359 (N_47359,N_47178,N_47191);
xor U47360 (N_47360,N_47222,N_47194);
and U47361 (N_47361,N_47122,N_47089);
nand U47362 (N_47362,N_47107,N_47023);
nor U47363 (N_47363,N_47111,N_47120);
or U47364 (N_47364,N_47220,N_47217);
nand U47365 (N_47365,N_47025,N_47175);
nand U47366 (N_47366,N_47145,N_47124);
nor U47367 (N_47367,N_47131,N_47014);
nand U47368 (N_47368,N_47137,N_47163);
nand U47369 (N_47369,N_47123,N_47034);
and U47370 (N_47370,N_47228,N_47223);
nand U47371 (N_47371,N_47129,N_47012);
xor U47372 (N_47372,N_47092,N_47248);
nor U47373 (N_47373,N_47061,N_47070);
nor U47374 (N_47374,N_47125,N_47165);
or U47375 (N_47375,N_47027,N_47168);
and U47376 (N_47376,N_47021,N_47241);
xnor U47377 (N_47377,N_47020,N_47033);
nand U47378 (N_47378,N_47145,N_47122);
nand U47379 (N_47379,N_47115,N_47049);
and U47380 (N_47380,N_47202,N_47079);
nor U47381 (N_47381,N_47091,N_47184);
nand U47382 (N_47382,N_47061,N_47125);
nand U47383 (N_47383,N_47145,N_47189);
and U47384 (N_47384,N_47247,N_47156);
xnor U47385 (N_47385,N_47154,N_47157);
or U47386 (N_47386,N_47174,N_47247);
nor U47387 (N_47387,N_47010,N_47000);
or U47388 (N_47388,N_47067,N_47188);
or U47389 (N_47389,N_47194,N_47004);
xnor U47390 (N_47390,N_47152,N_47120);
xnor U47391 (N_47391,N_47077,N_47016);
xnor U47392 (N_47392,N_47037,N_47020);
nor U47393 (N_47393,N_47167,N_47025);
xor U47394 (N_47394,N_47188,N_47099);
nand U47395 (N_47395,N_47138,N_47037);
and U47396 (N_47396,N_47021,N_47060);
or U47397 (N_47397,N_47215,N_47191);
nand U47398 (N_47398,N_47176,N_47076);
or U47399 (N_47399,N_47226,N_47129);
or U47400 (N_47400,N_47131,N_47225);
xnor U47401 (N_47401,N_47018,N_47226);
and U47402 (N_47402,N_47245,N_47177);
nand U47403 (N_47403,N_47046,N_47080);
xnor U47404 (N_47404,N_47208,N_47202);
nor U47405 (N_47405,N_47181,N_47120);
nand U47406 (N_47406,N_47112,N_47074);
xor U47407 (N_47407,N_47001,N_47041);
nor U47408 (N_47408,N_47196,N_47038);
and U47409 (N_47409,N_47098,N_47105);
and U47410 (N_47410,N_47129,N_47241);
or U47411 (N_47411,N_47033,N_47114);
or U47412 (N_47412,N_47156,N_47074);
xnor U47413 (N_47413,N_47037,N_47063);
nand U47414 (N_47414,N_47157,N_47024);
or U47415 (N_47415,N_47115,N_47028);
nor U47416 (N_47416,N_47055,N_47106);
and U47417 (N_47417,N_47194,N_47120);
and U47418 (N_47418,N_47143,N_47185);
xor U47419 (N_47419,N_47160,N_47089);
nor U47420 (N_47420,N_47223,N_47161);
nand U47421 (N_47421,N_47116,N_47123);
nand U47422 (N_47422,N_47075,N_47097);
nand U47423 (N_47423,N_47188,N_47063);
xor U47424 (N_47424,N_47246,N_47038);
xor U47425 (N_47425,N_47007,N_47012);
nand U47426 (N_47426,N_47128,N_47199);
and U47427 (N_47427,N_47222,N_47167);
nand U47428 (N_47428,N_47166,N_47114);
xor U47429 (N_47429,N_47171,N_47053);
nand U47430 (N_47430,N_47074,N_47200);
nand U47431 (N_47431,N_47199,N_47086);
and U47432 (N_47432,N_47155,N_47113);
and U47433 (N_47433,N_47050,N_47076);
nand U47434 (N_47434,N_47192,N_47043);
and U47435 (N_47435,N_47237,N_47076);
nand U47436 (N_47436,N_47072,N_47095);
and U47437 (N_47437,N_47248,N_47018);
xor U47438 (N_47438,N_47018,N_47157);
nor U47439 (N_47439,N_47056,N_47210);
xor U47440 (N_47440,N_47067,N_47201);
and U47441 (N_47441,N_47195,N_47222);
xor U47442 (N_47442,N_47161,N_47164);
xnor U47443 (N_47443,N_47186,N_47230);
and U47444 (N_47444,N_47085,N_47021);
xnor U47445 (N_47445,N_47046,N_47165);
xnor U47446 (N_47446,N_47092,N_47034);
and U47447 (N_47447,N_47142,N_47001);
nor U47448 (N_47448,N_47163,N_47135);
or U47449 (N_47449,N_47113,N_47160);
nand U47450 (N_47450,N_47158,N_47153);
nor U47451 (N_47451,N_47155,N_47239);
and U47452 (N_47452,N_47008,N_47192);
nor U47453 (N_47453,N_47106,N_47194);
nor U47454 (N_47454,N_47162,N_47025);
and U47455 (N_47455,N_47198,N_47086);
nand U47456 (N_47456,N_47103,N_47185);
nor U47457 (N_47457,N_47003,N_47137);
nor U47458 (N_47458,N_47188,N_47139);
xor U47459 (N_47459,N_47147,N_47210);
nand U47460 (N_47460,N_47060,N_47219);
and U47461 (N_47461,N_47033,N_47127);
or U47462 (N_47462,N_47111,N_47173);
or U47463 (N_47463,N_47215,N_47175);
nor U47464 (N_47464,N_47123,N_47056);
nand U47465 (N_47465,N_47150,N_47174);
nand U47466 (N_47466,N_47203,N_47017);
nand U47467 (N_47467,N_47173,N_47248);
nand U47468 (N_47468,N_47047,N_47112);
nand U47469 (N_47469,N_47087,N_47061);
or U47470 (N_47470,N_47142,N_47209);
nand U47471 (N_47471,N_47210,N_47191);
or U47472 (N_47472,N_47104,N_47040);
xor U47473 (N_47473,N_47088,N_47094);
and U47474 (N_47474,N_47050,N_47143);
and U47475 (N_47475,N_47189,N_47175);
and U47476 (N_47476,N_47218,N_47187);
and U47477 (N_47477,N_47013,N_47038);
and U47478 (N_47478,N_47173,N_47196);
or U47479 (N_47479,N_47092,N_47176);
and U47480 (N_47480,N_47146,N_47110);
nand U47481 (N_47481,N_47104,N_47092);
and U47482 (N_47482,N_47142,N_47107);
or U47483 (N_47483,N_47211,N_47130);
and U47484 (N_47484,N_47208,N_47028);
nand U47485 (N_47485,N_47093,N_47248);
nor U47486 (N_47486,N_47098,N_47157);
or U47487 (N_47487,N_47144,N_47212);
nand U47488 (N_47488,N_47095,N_47118);
xnor U47489 (N_47489,N_47236,N_47068);
or U47490 (N_47490,N_47003,N_47064);
or U47491 (N_47491,N_47215,N_47135);
nand U47492 (N_47492,N_47183,N_47086);
nor U47493 (N_47493,N_47087,N_47228);
xor U47494 (N_47494,N_47108,N_47236);
or U47495 (N_47495,N_47197,N_47068);
or U47496 (N_47496,N_47058,N_47034);
or U47497 (N_47497,N_47063,N_47146);
or U47498 (N_47498,N_47224,N_47240);
and U47499 (N_47499,N_47226,N_47168);
nor U47500 (N_47500,N_47334,N_47472);
and U47501 (N_47501,N_47347,N_47362);
xor U47502 (N_47502,N_47368,N_47402);
nand U47503 (N_47503,N_47441,N_47426);
and U47504 (N_47504,N_47346,N_47263);
nor U47505 (N_47505,N_47342,N_47376);
xnor U47506 (N_47506,N_47388,N_47470);
and U47507 (N_47507,N_47438,N_47449);
xnor U47508 (N_47508,N_47399,N_47297);
and U47509 (N_47509,N_47279,N_47433);
or U47510 (N_47510,N_47428,N_47341);
or U47511 (N_47511,N_47284,N_47272);
nand U47512 (N_47512,N_47309,N_47316);
and U47513 (N_47513,N_47325,N_47253);
xnor U47514 (N_47514,N_47375,N_47252);
nor U47515 (N_47515,N_47384,N_47398);
and U47516 (N_47516,N_47442,N_47327);
or U47517 (N_47517,N_47370,N_47357);
nor U47518 (N_47518,N_47372,N_47411);
nand U47519 (N_47519,N_47269,N_47460);
nand U47520 (N_47520,N_47331,N_47478);
and U47521 (N_47521,N_47355,N_47482);
xnor U47522 (N_47522,N_47320,N_47349);
nand U47523 (N_47523,N_47280,N_47466);
xor U47524 (N_47524,N_47359,N_47312);
or U47525 (N_47525,N_47400,N_47311);
nor U47526 (N_47526,N_47344,N_47407);
and U47527 (N_47527,N_47406,N_47317);
xor U47528 (N_47528,N_47439,N_47386);
xnor U47529 (N_47529,N_47454,N_47389);
xnor U47530 (N_47530,N_47260,N_47250);
and U47531 (N_47531,N_47262,N_47488);
xnor U47532 (N_47532,N_47358,N_47390);
and U47533 (N_47533,N_47274,N_47401);
nand U47534 (N_47534,N_47416,N_47427);
and U47535 (N_47535,N_47420,N_47373);
or U47536 (N_47536,N_47415,N_47292);
or U47537 (N_47537,N_47363,N_47458);
xnor U47538 (N_47538,N_47330,N_47383);
and U47539 (N_47539,N_47304,N_47282);
and U47540 (N_47540,N_47305,N_47483);
xor U47541 (N_47541,N_47385,N_47409);
nor U47542 (N_47542,N_47319,N_47289);
nand U47543 (N_47543,N_47307,N_47414);
and U47544 (N_47544,N_47417,N_47366);
or U47545 (N_47545,N_47369,N_47264);
xnor U47546 (N_47546,N_47410,N_47485);
nor U47547 (N_47547,N_47322,N_47294);
nand U47548 (N_47548,N_47451,N_47408);
and U47549 (N_47549,N_47403,N_47476);
or U47550 (N_47550,N_47266,N_47293);
nand U47551 (N_47551,N_47352,N_47382);
or U47552 (N_47552,N_47473,N_47450);
xnor U47553 (N_47553,N_47323,N_47397);
xnor U47554 (N_47554,N_47361,N_47469);
and U47555 (N_47555,N_47419,N_47437);
nand U47556 (N_47556,N_47275,N_47393);
xor U47557 (N_47557,N_47436,N_47475);
xor U47558 (N_47558,N_47430,N_47374);
and U47559 (N_47559,N_47423,N_47378);
xor U47560 (N_47560,N_47492,N_47429);
or U47561 (N_47561,N_47413,N_47295);
nand U47562 (N_47562,N_47455,N_47452);
nand U47563 (N_47563,N_47302,N_47300);
nor U47564 (N_47564,N_47490,N_47443);
xnor U47565 (N_47565,N_47281,N_47315);
xnor U47566 (N_47566,N_47259,N_47354);
and U47567 (N_47567,N_47424,N_47387);
or U47568 (N_47568,N_47299,N_47474);
and U47569 (N_47569,N_47444,N_47265);
and U47570 (N_47570,N_47287,N_47467);
nor U47571 (N_47571,N_47495,N_47425);
or U47572 (N_47572,N_47268,N_47360);
nor U47573 (N_47573,N_47493,N_47432);
and U47574 (N_47574,N_47499,N_47464);
or U47575 (N_47575,N_47498,N_47336);
and U47576 (N_47576,N_47494,N_47481);
xor U47577 (N_47577,N_47326,N_47343);
or U47578 (N_47578,N_47446,N_47258);
xnor U47579 (N_47579,N_47380,N_47276);
xor U47580 (N_47580,N_47285,N_47434);
xnor U47581 (N_47581,N_47313,N_47395);
or U47582 (N_47582,N_47487,N_47468);
or U47583 (N_47583,N_47496,N_47283);
xnor U47584 (N_47584,N_47333,N_47477);
and U47585 (N_47585,N_47457,N_47350);
xnor U47586 (N_47586,N_47277,N_47394);
or U47587 (N_47587,N_47271,N_47306);
nand U47588 (N_47588,N_47356,N_47270);
nor U47589 (N_47589,N_47301,N_47412);
and U47590 (N_47590,N_47445,N_47261);
or U47591 (N_47591,N_47329,N_47337);
nand U47592 (N_47592,N_47340,N_47456);
or U47593 (N_47593,N_47435,N_47484);
xor U47594 (N_47594,N_47377,N_47291);
nor U47595 (N_47595,N_47254,N_47440);
xnor U47596 (N_47596,N_47364,N_47480);
xnor U47597 (N_47597,N_47345,N_47491);
or U47598 (N_47598,N_47486,N_47328);
nor U47599 (N_47599,N_47351,N_47256);
nand U47600 (N_47600,N_47404,N_47296);
nor U47601 (N_47601,N_47267,N_47257);
or U47602 (N_47602,N_47339,N_47396);
or U47603 (N_47603,N_47353,N_47465);
and U47604 (N_47604,N_47303,N_47453);
or U47605 (N_47605,N_47286,N_47288);
xnor U47606 (N_47606,N_47418,N_47462);
nand U47607 (N_47607,N_47371,N_47290);
and U47608 (N_47608,N_47459,N_47391);
nand U47609 (N_47609,N_47447,N_47421);
nor U47610 (N_47610,N_47367,N_47348);
nor U47611 (N_47611,N_47278,N_47463);
or U47612 (N_47612,N_47431,N_47310);
and U47613 (N_47613,N_47324,N_47379);
or U47614 (N_47614,N_47365,N_47471);
nand U47615 (N_47615,N_47298,N_47255);
xnor U47616 (N_47616,N_47479,N_47318);
and U47617 (N_47617,N_47448,N_47338);
and U47618 (N_47618,N_47251,N_47321);
and U47619 (N_47619,N_47461,N_47497);
nand U47620 (N_47620,N_47273,N_47308);
or U47621 (N_47621,N_47392,N_47422);
nor U47622 (N_47622,N_47405,N_47335);
and U47623 (N_47623,N_47381,N_47489);
or U47624 (N_47624,N_47314,N_47332);
nor U47625 (N_47625,N_47258,N_47402);
and U47626 (N_47626,N_47277,N_47453);
or U47627 (N_47627,N_47463,N_47327);
xnor U47628 (N_47628,N_47467,N_47284);
or U47629 (N_47629,N_47442,N_47374);
nand U47630 (N_47630,N_47328,N_47367);
nor U47631 (N_47631,N_47499,N_47462);
or U47632 (N_47632,N_47451,N_47406);
and U47633 (N_47633,N_47376,N_47417);
nand U47634 (N_47634,N_47294,N_47343);
nor U47635 (N_47635,N_47327,N_47271);
or U47636 (N_47636,N_47433,N_47301);
nor U47637 (N_47637,N_47304,N_47311);
or U47638 (N_47638,N_47454,N_47327);
or U47639 (N_47639,N_47251,N_47404);
nand U47640 (N_47640,N_47359,N_47408);
and U47641 (N_47641,N_47390,N_47253);
nand U47642 (N_47642,N_47369,N_47259);
and U47643 (N_47643,N_47429,N_47362);
nand U47644 (N_47644,N_47366,N_47478);
nand U47645 (N_47645,N_47472,N_47366);
nor U47646 (N_47646,N_47256,N_47412);
or U47647 (N_47647,N_47478,N_47291);
nand U47648 (N_47648,N_47474,N_47311);
or U47649 (N_47649,N_47299,N_47259);
nor U47650 (N_47650,N_47461,N_47398);
nand U47651 (N_47651,N_47284,N_47489);
nand U47652 (N_47652,N_47263,N_47449);
or U47653 (N_47653,N_47358,N_47290);
or U47654 (N_47654,N_47363,N_47428);
xor U47655 (N_47655,N_47476,N_47260);
nand U47656 (N_47656,N_47420,N_47333);
and U47657 (N_47657,N_47465,N_47412);
xor U47658 (N_47658,N_47313,N_47322);
nor U47659 (N_47659,N_47334,N_47361);
nand U47660 (N_47660,N_47488,N_47456);
and U47661 (N_47661,N_47382,N_47475);
nand U47662 (N_47662,N_47393,N_47385);
or U47663 (N_47663,N_47483,N_47319);
xor U47664 (N_47664,N_47388,N_47264);
nand U47665 (N_47665,N_47318,N_47471);
nor U47666 (N_47666,N_47451,N_47476);
and U47667 (N_47667,N_47356,N_47268);
and U47668 (N_47668,N_47487,N_47316);
and U47669 (N_47669,N_47314,N_47337);
nor U47670 (N_47670,N_47412,N_47451);
or U47671 (N_47671,N_47385,N_47397);
and U47672 (N_47672,N_47402,N_47455);
nand U47673 (N_47673,N_47413,N_47443);
and U47674 (N_47674,N_47333,N_47331);
nor U47675 (N_47675,N_47485,N_47425);
or U47676 (N_47676,N_47492,N_47259);
nor U47677 (N_47677,N_47431,N_47278);
and U47678 (N_47678,N_47272,N_47287);
and U47679 (N_47679,N_47369,N_47291);
xnor U47680 (N_47680,N_47363,N_47378);
xnor U47681 (N_47681,N_47331,N_47321);
nand U47682 (N_47682,N_47268,N_47498);
xnor U47683 (N_47683,N_47300,N_47343);
xor U47684 (N_47684,N_47449,N_47402);
and U47685 (N_47685,N_47354,N_47376);
xnor U47686 (N_47686,N_47435,N_47309);
and U47687 (N_47687,N_47483,N_47369);
and U47688 (N_47688,N_47430,N_47433);
or U47689 (N_47689,N_47466,N_47481);
nor U47690 (N_47690,N_47260,N_47380);
nor U47691 (N_47691,N_47448,N_47380);
xor U47692 (N_47692,N_47277,N_47445);
nand U47693 (N_47693,N_47484,N_47457);
nor U47694 (N_47694,N_47483,N_47263);
nand U47695 (N_47695,N_47473,N_47311);
nor U47696 (N_47696,N_47479,N_47315);
nor U47697 (N_47697,N_47360,N_47281);
nor U47698 (N_47698,N_47458,N_47412);
nor U47699 (N_47699,N_47483,N_47285);
nor U47700 (N_47700,N_47367,N_47493);
or U47701 (N_47701,N_47357,N_47486);
and U47702 (N_47702,N_47497,N_47452);
nor U47703 (N_47703,N_47322,N_47254);
or U47704 (N_47704,N_47330,N_47362);
or U47705 (N_47705,N_47333,N_47362);
and U47706 (N_47706,N_47307,N_47441);
or U47707 (N_47707,N_47273,N_47318);
nand U47708 (N_47708,N_47273,N_47491);
or U47709 (N_47709,N_47458,N_47250);
and U47710 (N_47710,N_47281,N_47276);
and U47711 (N_47711,N_47350,N_47276);
xor U47712 (N_47712,N_47404,N_47490);
and U47713 (N_47713,N_47381,N_47328);
nor U47714 (N_47714,N_47470,N_47341);
or U47715 (N_47715,N_47393,N_47316);
or U47716 (N_47716,N_47474,N_47446);
nor U47717 (N_47717,N_47314,N_47471);
nand U47718 (N_47718,N_47413,N_47345);
nor U47719 (N_47719,N_47371,N_47390);
nor U47720 (N_47720,N_47261,N_47326);
or U47721 (N_47721,N_47292,N_47393);
nor U47722 (N_47722,N_47390,N_47491);
and U47723 (N_47723,N_47499,N_47254);
nand U47724 (N_47724,N_47449,N_47491);
nor U47725 (N_47725,N_47361,N_47270);
and U47726 (N_47726,N_47410,N_47495);
or U47727 (N_47727,N_47392,N_47435);
and U47728 (N_47728,N_47398,N_47416);
or U47729 (N_47729,N_47364,N_47348);
nand U47730 (N_47730,N_47490,N_47347);
nand U47731 (N_47731,N_47342,N_47421);
or U47732 (N_47732,N_47327,N_47435);
and U47733 (N_47733,N_47482,N_47436);
and U47734 (N_47734,N_47258,N_47404);
and U47735 (N_47735,N_47352,N_47366);
xnor U47736 (N_47736,N_47407,N_47391);
and U47737 (N_47737,N_47385,N_47434);
and U47738 (N_47738,N_47387,N_47272);
or U47739 (N_47739,N_47440,N_47251);
nor U47740 (N_47740,N_47446,N_47404);
nor U47741 (N_47741,N_47388,N_47302);
xnor U47742 (N_47742,N_47315,N_47401);
xor U47743 (N_47743,N_47250,N_47418);
nor U47744 (N_47744,N_47408,N_47281);
xnor U47745 (N_47745,N_47482,N_47258);
nand U47746 (N_47746,N_47418,N_47271);
or U47747 (N_47747,N_47318,N_47278);
xnor U47748 (N_47748,N_47439,N_47421);
and U47749 (N_47749,N_47496,N_47355);
and U47750 (N_47750,N_47665,N_47522);
and U47751 (N_47751,N_47738,N_47671);
xor U47752 (N_47752,N_47623,N_47592);
xnor U47753 (N_47753,N_47547,N_47652);
nor U47754 (N_47754,N_47563,N_47667);
nor U47755 (N_47755,N_47698,N_47719);
nor U47756 (N_47756,N_47553,N_47622);
xnor U47757 (N_47757,N_47700,N_47525);
xor U47758 (N_47758,N_47554,N_47741);
nand U47759 (N_47759,N_47678,N_47580);
nand U47760 (N_47760,N_47558,N_47636);
xnor U47761 (N_47761,N_47718,N_47562);
nand U47762 (N_47762,N_47735,N_47542);
and U47763 (N_47763,N_47617,N_47722);
nand U47764 (N_47764,N_47744,N_47520);
xnor U47765 (N_47765,N_47610,N_47612);
or U47766 (N_47766,N_47635,N_47535);
nand U47767 (N_47767,N_47666,N_47685);
xnor U47768 (N_47768,N_47658,N_47601);
or U47769 (N_47769,N_47515,N_47697);
and U47770 (N_47770,N_47591,N_47713);
nor U47771 (N_47771,N_47573,N_47587);
nor U47772 (N_47772,N_47729,N_47651);
xnor U47773 (N_47773,N_47707,N_47672);
and U47774 (N_47774,N_47708,N_47680);
nor U47775 (N_47775,N_47543,N_47732);
or U47776 (N_47776,N_47711,N_47557);
or U47777 (N_47777,N_47609,N_47699);
nor U47778 (N_47778,N_47584,N_47546);
and U47779 (N_47779,N_47613,N_47724);
and U47780 (N_47780,N_47510,N_47620);
and U47781 (N_47781,N_47728,N_47602);
xor U47782 (N_47782,N_47673,N_47508);
nand U47783 (N_47783,N_47717,N_47626);
nor U47784 (N_47784,N_47649,N_47749);
xor U47785 (N_47785,N_47569,N_47637);
and U47786 (N_47786,N_47507,N_47643);
and U47787 (N_47787,N_47502,N_47551);
and U47788 (N_47788,N_47527,N_47555);
and U47789 (N_47789,N_47536,N_47568);
and U47790 (N_47790,N_47632,N_47593);
nor U47791 (N_47791,N_47571,N_47677);
or U47792 (N_47792,N_47605,N_47552);
xnor U47793 (N_47793,N_47648,N_47519);
xnor U47794 (N_47794,N_47664,N_47606);
or U47795 (N_47795,N_47681,N_47630);
nand U47796 (N_47796,N_47682,N_47726);
xnor U47797 (N_47797,N_47559,N_47505);
nor U47798 (N_47798,N_47514,N_47663);
or U47799 (N_47799,N_47687,N_47572);
xnor U47800 (N_47800,N_47598,N_47590);
and U47801 (N_47801,N_47742,N_47692);
xnor U47802 (N_47802,N_47529,N_47662);
and U47803 (N_47803,N_47588,N_47720);
nor U47804 (N_47804,N_47675,N_47693);
or U47805 (N_47805,N_47701,N_47653);
nor U47806 (N_47806,N_47511,N_47631);
nand U47807 (N_47807,N_47556,N_47704);
or U47808 (N_47808,N_47585,N_47595);
nor U47809 (N_47809,N_47688,N_47731);
nor U47810 (N_47810,N_47624,N_47594);
and U47811 (N_47811,N_47538,N_47570);
nor U47812 (N_47812,N_47560,N_47581);
and U47813 (N_47813,N_47628,N_47714);
nor U47814 (N_47814,N_47725,N_47577);
and U47815 (N_47815,N_47616,N_47670);
xnor U47816 (N_47816,N_47621,N_47625);
and U47817 (N_47817,N_47712,N_47716);
nand U47818 (N_47818,N_47524,N_47549);
or U47819 (N_47819,N_47539,N_47545);
nor U47820 (N_47820,N_47639,N_47506);
and U47821 (N_47821,N_47574,N_47611);
xor U47822 (N_47822,N_47661,N_47565);
nand U47823 (N_47823,N_47743,N_47509);
nand U47824 (N_47824,N_47532,N_47674);
or U47825 (N_47825,N_47596,N_47597);
xnor U47826 (N_47826,N_47721,N_47575);
and U47827 (N_47827,N_47702,N_47715);
xor U47828 (N_47828,N_47654,N_47646);
xor U47829 (N_47829,N_47534,N_47660);
nand U47830 (N_47830,N_47600,N_47736);
xnor U47831 (N_47831,N_47608,N_47541);
and U47832 (N_47832,N_47684,N_47727);
nand U47833 (N_47833,N_47676,N_47504);
nand U47834 (N_47834,N_47564,N_47657);
nand U47835 (N_47835,N_47691,N_47523);
and U47836 (N_47836,N_47544,N_47537);
nand U47837 (N_47837,N_47740,N_47583);
nand U47838 (N_47838,N_47703,N_47747);
nand U47839 (N_47839,N_47530,N_47513);
nor U47840 (N_47840,N_47690,N_47645);
nand U47841 (N_47841,N_47618,N_47614);
nor U47842 (N_47842,N_47650,N_47589);
nor U47843 (N_47843,N_47723,N_47501);
nand U47844 (N_47844,N_47655,N_47533);
nand U47845 (N_47845,N_47604,N_47512);
or U47846 (N_47846,N_47550,N_47500);
nor U47847 (N_47847,N_47634,N_47709);
and U47848 (N_47848,N_47582,N_47696);
or U47849 (N_47849,N_47705,N_47516);
or U47850 (N_47850,N_47710,N_47633);
and U47851 (N_47851,N_47668,N_47615);
or U47852 (N_47852,N_47734,N_47517);
and U47853 (N_47853,N_47642,N_47521);
nand U47854 (N_47854,N_47518,N_47683);
and U47855 (N_47855,N_47561,N_47733);
or U47856 (N_47856,N_47566,N_47638);
xor U47857 (N_47857,N_47540,N_47689);
xor U47858 (N_47858,N_47586,N_47579);
nor U47859 (N_47859,N_47627,N_47619);
nor U47860 (N_47860,N_47548,N_47531);
or U47861 (N_47861,N_47739,N_47503);
nor U47862 (N_47862,N_47640,N_47746);
and U47863 (N_47863,N_47686,N_47695);
nand U47864 (N_47864,N_47730,N_47603);
xnor U47865 (N_47865,N_47659,N_47706);
xnor U47866 (N_47866,N_47679,N_47528);
or U47867 (N_47867,N_47644,N_47526);
nand U47868 (N_47868,N_47629,N_47656);
or U47869 (N_47869,N_47599,N_47578);
or U47870 (N_47870,N_47748,N_47641);
nor U47871 (N_47871,N_47567,N_47647);
or U47872 (N_47872,N_47669,N_47745);
and U47873 (N_47873,N_47576,N_47607);
nand U47874 (N_47874,N_47694,N_47737);
or U47875 (N_47875,N_47644,N_47746);
or U47876 (N_47876,N_47726,N_47511);
nand U47877 (N_47877,N_47594,N_47614);
nor U47878 (N_47878,N_47570,N_47670);
or U47879 (N_47879,N_47577,N_47589);
xnor U47880 (N_47880,N_47527,N_47586);
and U47881 (N_47881,N_47717,N_47594);
nand U47882 (N_47882,N_47536,N_47639);
xnor U47883 (N_47883,N_47628,N_47710);
or U47884 (N_47884,N_47656,N_47675);
xor U47885 (N_47885,N_47697,N_47724);
nand U47886 (N_47886,N_47604,N_47594);
nand U47887 (N_47887,N_47574,N_47624);
nand U47888 (N_47888,N_47638,N_47608);
or U47889 (N_47889,N_47579,N_47748);
and U47890 (N_47890,N_47710,N_47539);
or U47891 (N_47891,N_47588,N_47547);
and U47892 (N_47892,N_47749,N_47614);
nor U47893 (N_47893,N_47705,N_47713);
xor U47894 (N_47894,N_47600,N_47574);
or U47895 (N_47895,N_47698,N_47740);
and U47896 (N_47896,N_47689,N_47635);
nand U47897 (N_47897,N_47570,N_47633);
xnor U47898 (N_47898,N_47605,N_47622);
xnor U47899 (N_47899,N_47519,N_47618);
nand U47900 (N_47900,N_47739,N_47666);
nor U47901 (N_47901,N_47639,N_47541);
nor U47902 (N_47902,N_47503,N_47737);
or U47903 (N_47903,N_47523,N_47714);
nor U47904 (N_47904,N_47518,N_47667);
nand U47905 (N_47905,N_47664,N_47651);
or U47906 (N_47906,N_47511,N_47677);
and U47907 (N_47907,N_47598,N_47719);
and U47908 (N_47908,N_47724,N_47741);
nand U47909 (N_47909,N_47569,N_47573);
nand U47910 (N_47910,N_47691,N_47638);
or U47911 (N_47911,N_47739,N_47516);
and U47912 (N_47912,N_47560,N_47508);
and U47913 (N_47913,N_47564,N_47735);
xor U47914 (N_47914,N_47722,N_47665);
xnor U47915 (N_47915,N_47556,N_47653);
and U47916 (N_47916,N_47680,N_47546);
nand U47917 (N_47917,N_47558,N_47631);
or U47918 (N_47918,N_47593,N_47718);
or U47919 (N_47919,N_47652,N_47662);
nand U47920 (N_47920,N_47698,N_47516);
xnor U47921 (N_47921,N_47657,N_47573);
nor U47922 (N_47922,N_47589,N_47715);
and U47923 (N_47923,N_47721,N_47742);
nor U47924 (N_47924,N_47505,N_47682);
nor U47925 (N_47925,N_47736,N_47570);
and U47926 (N_47926,N_47615,N_47744);
or U47927 (N_47927,N_47747,N_47551);
xor U47928 (N_47928,N_47706,N_47554);
nand U47929 (N_47929,N_47607,N_47543);
xnor U47930 (N_47930,N_47577,N_47641);
and U47931 (N_47931,N_47662,N_47570);
nand U47932 (N_47932,N_47553,N_47621);
nand U47933 (N_47933,N_47538,N_47621);
nand U47934 (N_47934,N_47738,N_47517);
nand U47935 (N_47935,N_47719,N_47691);
and U47936 (N_47936,N_47714,N_47710);
and U47937 (N_47937,N_47701,N_47597);
nand U47938 (N_47938,N_47629,N_47718);
nor U47939 (N_47939,N_47667,N_47619);
and U47940 (N_47940,N_47521,N_47612);
and U47941 (N_47941,N_47638,N_47557);
nand U47942 (N_47942,N_47742,N_47597);
and U47943 (N_47943,N_47702,N_47708);
or U47944 (N_47944,N_47614,N_47613);
xor U47945 (N_47945,N_47646,N_47554);
or U47946 (N_47946,N_47678,N_47725);
and U47947 (N_47947,N_47559,N_47655);
nor U47948 (N_47948,N_47611,N_47625);
or U47949 (N_47949,N_47528,N_47537);
nor U47950 (N_47950,N_47560,N_47698);
and U47951 (N_47951,N_47703,N_47723);
nand U47952 (N_47952,N_47500,N_47554);
or U47953 (N_47953,N_47698,N_47726);
and U47954 (N_47954,N_47608,N_47566);
or U47955 (N_47955,N_47660,N_47590);
nor U47956 (N_47956,N_47584,N_47626);
xor U47957 (N_47957,N_47747,N_47669);
nand U47958 (N_47958,N_47679,N_47702);
xnor U47959 (N_47959,N_47525,N_47602);
nor U47960 (N_47960,N_47599,N_47678);
nand U47961 (N_47961,N_47570,N_47706);
or U47962 (N_47962,N_47671,N_47559);
or U47963 (N_47963,N_47544,N_47594);
xnor U47964 (N_47964,N_47682,N_47737);
xnor U47965 (N_47965,N_47579,N_47603);
nor U47966 (N_47966,N_47678,N_47526);
xor U47967 (N_47967,N_47647,N_47565);
or U47968 (N_47968,N_47504,N_47614);
xor U47969 (N_47969,N_47579,N_47720);
nand U47970 (N_47970,N_47644,N_47583);
nand U47971 (N_47971,N_47548,N_47663);
xnor U47972 (N_47972,N_47737,N_47723);
or U47973 (N_47973,N_47528,N_47697);
nor U47974 (N_47974,N_47532,N_47672);
nand U47975 (N_47975,N_47703,N_47591);
nand U47976 (N_47976,N_47650,N_47734);
and U47977 (N_47977,N_47745,N_47505);
nor U47978 (N_47978,N_47711,N_47531);
xor U47979 (N_47979,N_47511,N_47500);
and U47980 (N_47980,N_47532,N_47692);
nor U47981 (N_47981,N_47562,N_47685);
and U47982 (N_47982,N_47581,N_47528);
nor U47983 (N_47983,N_47581,N_47539);
or U47984 (N_47984,N_47679,N_47688);
nor U47985 (N_47985,N_47548,N_47673);
or U47986 (N_47986,N_47681,N_47552);
nor U47987 (N_47987,N_47650,N_47513);
or U47988 (N_47988,N_47682,N_47687);
or U47989 (N_47989,N_47709,N_47600);
nand U47990 (N_47990,N_47617,N_47644);
and U47991 (N_47991,N_47558,N_47672);
nor U47992 (N_47992,N_47687,N_47684);
nor U47993 (N_47993,N_47626,N_47557);
nand U47994 (N_47994,N_47636,N_47675);
or U47995 (N_47995,N_47516,N_47710);
nand U47996 (N_47996,N_47550,N_47622);
nand U47997 (N_47997,N_47649,N_47508);
nand U47998 (N_47998,N_47674,N_47672);
and U47999 (N_47999,N_47608,N_47639);
nor U48000 (N_48000,N_47777,N_47947);
nor U48001 (N_48001,N_47902,N_47849);
xor U48002 (N_48002,N_47806,N_47984);
xnor U48003 (N_48003,N_47916,N_47889);
xnor U48004 (N_48004,N_47758,N_47816);
nor U48005 (N_48005,N_47990,N_47839);
and U48006 (N_48006,N_47956,N_47786);
and U48007 (N_48007,N_47830,N_47815);
nand U48008 (N_48008,N_47941,N_47986);
xor U48009 (N_48009,N_47919,N_47912);
or U48010 (N_48010,N_47923,N_47868);
and U48011 (N_48011,N_47996,N_47794);
and U48012 (N_48012,N_47904,N_47826);
nand U48013 (N_48013,N_47999,N_47860);
or U48014 (N_48014,N_47811,N_47775);
nor U48015 (N_48015,N_47994,N_47952);
or U48016 (N_48016,N_47931,N_47778);
nor U48017 (N_48017,N_47870,N_47782);
xor U48018 (N_48018,N_47836,N_47971);
nor U48019 (N_48019,N_47965,N_47881);
nand U48020 (N_48020,N_47762,N_47877);
or U48021 (N_48021,N_47873,N_47938);
xnor U48022 (N_48022,N_47825,N_47822);
or U48023 (N_48023,N_47942,N_47917);
nor U48024 (N_48024,N_47897,N_47759);
and U48025 (N_48025,N_47765,N_47903);
nand U48026 (N_48026,N_47973,N_47892);
and U48027 (N_48027,N_47751,N_47878);
nand U48028 (N_48028,N_47769,N_47954);
nand U48029 (N_48029,N_47953,N_47851);
nor U48030 (N_48030,N_47850,N_47812);
or U48031 (N_48031,N_47933,N_47977);
nand U48032 (N_48032,N_47930,N_47779);
nand U48033 (N_48033,N_47798,N_47987);
and U48034 (N_48034,N_47966,N_47792);
or U48035 (N_48035,N_47885,N_47799);
nor U48036 (N_48036,N_47863,N_47985);
nor U48037 (N_48037,N_47837,N_47832);
nor U48038 (N_48038,N_47752,N_47879);
xnor U48039 (N_48039,N_47796,N_47784);
and U48040 (N_48040,N_47886,N_47962);
nor U48041 (N_48041,N_47963,N_47924);
and U48042 (N_48042,N_47970,N_47757);
xnor U48043 (N_48043,N_47833,N_47835);
xnor U48044 (N_48044,N_47969,N_47838);
nor U48045 (N_48045,N_47896,N_47937);
and U48046 (N_48046,N_47857,N_47859);
or U48047 (N_48047,N_47880,N_47824);
nand U48048 (N_48048,N_47895,N_47867);
nor U48049 (N_48049,N_47927,N_47913);
or U48050 (N_48050,N_47972,N_47831);
and U48051 (N_48051,N_47813,N_47773);
nor U48052 (N_48052,N_47866,N_47855);
xnor U48053 (N_48053,N_47764,N_47852);
or U48054 (N_48054,N_47906,N_47801);
and U48055 (N_48055,N_47891,N_47774);
and U48056 (N_48056,N_47894,N_47959);
and U48057 (N_48057,N_47958,N_47793);
nor U48058 (N_48058,N_47946,N_47900);
or U48059 (N_48059,N_47795,N_47817);
and U48060 (N_48060,N_47797,N_47898);
nand U48061 (N_48061,N_47763,N_47842);
nand U48062 (N_48062,N_47772,N_47928);
xor U48063 (N_48063,N_47869,N_47935);
xnor U48064 (N_48064,N_47968,N_47908);
and U48065 (N_48065,N_47940,N_47929);
nor U48066 (N_48066,N_47858,N_47805);
xnor U48067 (N_48067,N_47945,N_47809);
and U48068 (N_48068,N_47800,N_47808);
nand U48069 (N_48069,N_47883,N_47993);
xnor U48070 (N_48070,N_47807,N_47767);
and U48071 (N_48071,N_47934,N_47997);
xor U48072 (N_48072,N_47982,N_47820);
or U48073 (N_48073,N_47932,N_47888);
nand U48074 (N_48074,N_47964,N_47846);
and U48075 (N_48075,N_47814,N_47834);
or U48076 (N_48076,N_47939,N_47998);
xnor U48077 (N_48077,N_47770,N_47988);
nand U48078 (N_48078,N_47991,N_47979);
xor U48079 (N_48079,N_47871,N_47949);
nor U48080 (N_48080,N_47862,N_47865);
xnor U48081 (N_48081,N_47890,N_47948);
xnor U48082 (N_48082,N_47915,N_47944);
and U48083 (N_48083,N_47783,N_47840);
and U48084 (N_48084,N_47844,N_47901);
nor U48085 (N_48085,N_47776,N_47920);
xor U48086 (N_48086,N_47887,N_47950);
nor U48087 (N_48087,N_47914,N_47847);
or U48088 (N_48088,N_47899,N_47853);
or U48089 (N_48089,N_47926,N_47874);
nand U48090 (N_48090,N_47961,N_47995);
nand U48091 (N_48091,N_47976,N_47921);
nor U48092 (N_48092,N_47829,N_47967);
nand U48093 (N_48093,N_47856,N_47756);
nand U48094 (N_48094,N_47978,N_47909);
nor U48095 (N_48095,N_47980,N_47754);
and U48096 (N_48096,N_47843,N_47788);
xnor U48097 (N_48097,N_47893,N_47781);
xor U48098 (N_48098,N_47876,N_47955);
and U48099 (N_48099,N_47848,N_47790);
or U48100 (N_48100,N_47760,N_47827);
and U48101 (N_48101,N_47755,N_47960);
nor U48102 (N_48102,N_47907,N_47828);
nand U48103 (N_48103,N_47753,N_47823);
or U48104 (N_48104,N_47802,N_47785);
or U48105 (N_48105,N_47943,N_47918);
xnor U48106 (N_48106,N_47936,N_47819);
nor U48107 (N_48107,N_47861,N_47818);
xnor U48108 (N_48108,N_47922,N_47974);
nor U48109 (N_48109,N_47791,N_47975);
nor U48110 (N_48110,N_47780,N_47951);
or U48111 (N_48111,N_47957,N_47821);
or U48112 (N_48112,N_47983,N_47804);
xor U48113 (N_48113,N_47925,N_47992);
xnor U48114 (N_48114,N_47989,N_47905);
or U48115 (N_48115,N_47981,N_47875);
nor U48116 (N_48116,N_47761,N_47771);
nor U48117 (N_48117,N_47910,N_47854);
nand U48118 (N_48118,N_47872,N_47884);
nor U48119 (N_48119,N_47911,N_47810);
nor U48120 (N_48120,N_47768,N_47766);
nand U48121 (N_48121,N_47789,N_47864);
xnor U48122 (N_48122,N_47882,N_47841);
and U48123 (N_48123,N_47845,N_47787);
and U48124 (N_48124,N_47750,N_47803);
nand U48125 (N_48125,N_47988,N_47920);
xor U48126 (N_48126,N_47911,N_47993);
nand U48127 (N_48127,N_47914,N_47765);
xnor U48128 (N_48128,N_47804,N_47846);
or U48129 (N_48129,N_47949,N_47823);
nor U48130 (N_48130,N_47757,N_47794);
and U48131 (N_48131,N_47820,N_47821);
nor U48132 (N_48132,N_47877,N_47858);
and U48133 (N_48133,N_47764,N_47888);
and U48134 (N_48134,N_47921,N_47788);
nor U48135 (N_48135,N_47912,N_47767);
nor U48136 (N_48136,N_47760,N_47992);
xnor U48137 (N_48137,N_47801,N_47802);
xor U48138 (N_48138,N_47958,N_47923);
nor U48139 (N_48139,N_47934,N_47939);
xor U48140 (N_48140,N_47888,N_47982);
or U48141 (N_48141,N_47795,N_47784);
nand U48142 (N_48142,N_47998,N_47982);
nor U48143 (N_48143,N_47923,N_47898);
xor U48144 (N_48144,N_47838,N_47918);
and U48145 (N_48145,N_47878,N_47872);
or U48146 (N_48146,N_47917,N_47944);
nand U48147 (N_48147,N_47957,N_47907);
nor U48148 (N_48148,N_47940,N_47992);
nor U48149 (N_48149,N_47869,N_47929);
xnor U48150 (N_48150,N_47878,N_47761);
or U48151 (N_48151,N_47771,N_47913);
nor U48152 (N_48152,N_47882,N_47759);
xor U48153 (N_48153,N_47870,N_47892);
nor U48154 (N_48154,N_47829,N_47804);
nand U48155 (N_48155,N_47784,N_47757);
and U48156 (N_48156,N_47773,N_47787);
nand U48157 (N_48157,N_47817,N_47909);
nand U48158 (N_48158,N_47974,N_47870);
nor U48159 (N_48159,N_47904,N_47887);
and U48160 (N_48160,N_47987,N_47981);
or U48161 (N_48161,N_47864,N_47820);
and U48162 (N_48162,N_47904,N_47869);
nor U48163 (N_48163,N_47783,N_47821);
nor U48164 (N_48164,N_47847,N_47890);
nand U48165 (N_48165,N_47793,N_47976);
xor U48166 (N_48166,N_47771,N_47793);
and U48167 (N_48167,N_47932,N_47845);
nor U48168 (N_48168,N_47810,N_47931);
xnor U48169 (N_48169,N_47766,N_47978);
xnor U48170 (N_48170,N_47891,N_47802);
and U48171 (N_48171,N_47879,N_47922);
nand U48172 (N_48172,N_47968,N_47901);
xor U48173 (N_48173,N_47778,N_47956);
and U48174 (N_48174,N_47956,N_47919);
nor U48175 (N_48175,N_47860,N_47925);
nand U48176 (N_48176,N_47871,N_47768);
nor U48177 (N_48177,N_47770,N_47994);
or U48178 (N_48178,N_47758,N_47824);
nand U48179 (N_48179,N_47902,N_47972);
or U48180 (N_48180,N_47771,N_47918);
nand U48181 (N_48181,N_47973,N_47912);
nor U48182 (N_48182,N_47965,N_47847);
xnor U48183 (N_48183,N_47855,N_47942);
xnor U48184 (N_48184,N_47928,N_47831);
xnor U48185 (N_48185,N_47860,N_47962);
xor U48186 (N_48186,N_47950,N_47992);
and U48187 (N_48187,N_47902,N_47863);
nand U48188 (N_48188,N_47898,N_47954);
nor U48189 (N_48189,N_47980,N_47875);
xnor U48190 (N_48190,N_47861,N_47881);
xnor U48191 (N_48191,N_47842,N_47753);
nand U48192 (N_48192,N_47849,N_47956);
nand U48193 (N_48193,N_47767,N_47819);
nand U48194 (N_48194,N_47805,N_47884);
or U48195 (N_48195,N_47781,N_47921);
and U48196 (N_48196,N_47938,N_47796);
nand U48197 (N_48197,N_47975,N_47843);
nand U48198 (N_48198,N_47952,N_47809);
and U48199 (N_48199,N_47963,N_47940);
nor U48200 (N_48200,N_47977,N_47904);
and U48201 (N_48201,N_47980,N_47837);
and U48202 (N_48202,N_47907,N_47855);
xnor U48203 (N_48203,N_47831,N_47821);
and U48204 (N_48204,N_47817,N_47812);
nand U48205 (N_48205,N_47809,N_47799);
nor U48206 (N_48206,N_47774,N_47783);
xnor U48207 (N_48207,N_47768,N_47855);
nor U48208 (N_48208,N_47848,N_47961);
and U48209 (N_48209,N_47871,N_47834);
nor U48210 (N_48210,N_47926,N_47989);
nor U48211 (N_48211,N_47884,N_47827);
xor U48212 (N_48212,N_47892,N_47943);
xnor U48213 (N_48213,N_47801,N_47769);
or U48214 (N_48214,N_47876,N_47999);
nand U48215 (N_48215,N_47754,N_47796);
or U48216 (N_48216,N_47828,N_47955);
nand U48217 (N_48217,N_47818,N_47821);
xor U48218 (N_48218,N_47921,N_47813);
nand U48219 (N_48219,N_47756,N_47787);
nand U48220 (N_48220,N_47872,N_47858);
and U48221 (N_48221,N_47974,N_47882);
nand U48222 (N_48222,N_47865,N_47874);
nand U48223 (N_48223,N_47945,N_47840);
nor U48224 (N_48224,N_47909,N_47756);
xnor U48225 (N_48225,N_47784,N_47765);
and U48226 (N_48226,N_47791,N_47984);
and U48227 (N_48227,N_47788,N_47760);
or U48228 (N_48228,N_47914,N_47797);
xor U48229 (N_48229,N_47980,N_47991);
or U48230 (N_48230,N_47860,N_47838);
nand U48231 (N_48231,N_47945,N_47977);
and U48232 (N_48232,N_47796,N_47801);
nand U48233 (N_48233,N_47763,N_47767);
and U48234 (N_48234,N_47995,N_47853);
or U48235 (N_48235,N_47997,N_47866);
and U48236 (N_48236,N_47940,N_47764);
xor U48237 (N_48237,N_47831,N_47769);
nand U48238 (N_48238,N_47757,N_47960);
and U48239 (N_48239,N_47959,N_47848);
nand U48240 (N_48240,N_47813,N_47812);
and U48241 (N_48241,N_47756,N_47997);
nor U48242 (N_48242,N_47752,N_47860);
xnor U48243 (N_48243,N_47855,N_47890);
and U48244 (N_48244,N_47989,N_47956);
nand U48245 (N_48245,N_47896,N_47798);
nand U48246 (N_48246,N_47847,N_47803);
nand U48247 (N_48247,N_47854,N_47878);
nor U48248 (N_48248,N_47811,N_47887);
and U48249 (N_48249,N_47926,N_47845);
and U48250 (N_48250,N_48096,N_48057);
and U48251 (N_48251,N_48054,N_48052);
nor U48252 (N_48252,N_48132,N_48009);
nor U48253 (N_48253,N_48138,N_48160);
nand U48254 (N_48254,N_48021,N_48166);
and U48255 (N_48255,N_48015,N_48190);
nor U48256 (N_48256,N_48192,N_48134);
nand U48257 (N_48257,N_48078,N_48083);
xnor U48258 (N_48258,N_48025,N_48189);
or U48259 (N_48259,N_48149,N_48048);
nand U48260 (N_48260,N_48196,N_48073);
and U48261 (N_48261,N_48191,N_48087);
nor U48262 (N_48262,N_48065,N_48042);
or U48263 (N_48263,N_48169,N_48067);
xor U48264 (N_48264,N_48049,N_48234);
nand U48265 (N_48265,N_48144,N_48116);
nor U48266 (N_48266,N_48123,N_48024);
and U48267 (N_48267,N_48075,N_48107);
or U48268 (N_48268,N_48247,N_48212);
nor U48269 (N_48269,N_48173,N_48245);
nand U48270 (N_48270,N_48017,N_48003);
nand U48271 (N_48271,N_48040,N_48037);
xor U48272 (N_48272,N_48239,N_48238);
or U48273 (N_48273,N_48027,N_48185);
xnor U48274 (N_48274,N_48181,N_48146);
nor U48275 (N_48275,N_48228,N_48224);
nor U48276 (N_48276,N_48214,N_48094);
or U48277 (N_48277,N_48063,N_48165);
nor U48278 (N_48278,N_48005,N_48104);
xor U48279 (N_48279,N_48120,N_48044);
nor U48280 (N_48280,N_48227,N_48151);
and U48281 (N_48281,N_48032,N_48202);
or U48282 (N_48282,N_48090,N_48208);
nand U48283 (N_48283,N_48117,N_48225);
nand U48284 (N_48284,N_48112,N_48204);
nor U48285 (N_48285,N_48122,N_48060);
and U48286 (N_48286,N_48100,N_48001);
nand U48287 (N_48287,N_48156,N_48176);
nor U48288 (N_48288,N_48193,N_48110);
and U48289 (N_48289,N_48220,N_48158);
xnor U48290 (N_48290,N_48233,N_48179);
and U48291 (N_48291,N_48168,N_48219);
nor U48292 (N_48292,N_48171,N_48079);
nor U48293 (N_48293,N_48127,N_48201);
nor U48294 (N_48294,N_48036,N_48035);
or U48295 (N_48295,N_48115,N_48246);
xor U48296 (N_48296,N_48126,N_48205);
xor U48297 (N_48297,N_48241,N_48231);
or U48298 (N_48298,N_48172,N_48153);
nand U48299 (N_48299,N_48125,N_48137);
and U48300 (N_48300,N_48199,N_48031);
xor U48301 (N_48301,N_48213,N_48047);
nand U48302 (N_48302,N_48098,N_48046);
nand U48303 (N_48303,N_48092,N_48142);
xor U48304 (N_48304,N_48119,N_48174);
and U48305 (N_48305,N_48053,N_48170);
nor U48306 (N_48306,N_48089,N_48136);
nor U48307 (N_48307,N_48108,N_48178);
or U48308 (N_48308,N_48121,N_48163);
and U48309 (N_48309,N_48041,N_48018);
nor U48310 (N_48310,N_48043,N_48050);
xor U48311 (N_48311,N_48081,N_48222);
and U48312 (N_48312,N_48091,N_48064);
nand U48313 (N_48313,N_48240,N_48097);
nor U48314 (N_48314,N_48135,N_48070);
xnor U48315 (N_48315,N_48210,N_48232);
nor U48316 (N_48316,N_48086,N_48131);
or U48317 (N_48317,N_48162,N_48159);
and U48318 (N_48318,N_48038,N_48129);
nand U48319 (N_48319,N_48128,N_48061);
nor U48320 (N_48320,N_48106,N_48074);
nand U48321 (N_48321,N_48195,N_48150);
xnor U48322 (N_48322,N_48184,N_48026);
xnor U48323 (N_48323,N_48130,N_48230);
and U48324 (N_48324,N_48167,N_48180);
xor U48325 (N_48325,N_48029,N_48010);
or U48326 (N_48326,N_48084,N_48071);
nor U48327 (N_48327,N_48113,N_48226);
nor U48328 (N_48328,N_48237,N_48243);
xor U48329 (N_48329,N_48218,N_48013);
nand U48330 (N_48330,N_48066,N_48101);
nand U48331 (N_48331,N_48088,N_48242);
and U48332 (N_48332,N_48068,N_48177);
and U48333 (N_48333,N_48055,N_48140);
nor U48334 (N_48334,N_48058,N_48248);
nor U48335 (N_48335,N_48207,N_48235);
or U48336 (N_48336,N_48229,N_48186);
xnor U48337 (N_48337,N_48152,N_48155);
and U48338 (N_48338,N_48102,N_48093);
or U48339 (N_48339,N_48188,N_48175);
and U48340 (N_48340,N_48076,N_48236);
xor U48341 (N_48341,N_48124,N_48016);
xnor U48342 (N_48342,N_48139,N_48011);
nand U48343 (N_48343,N_48069,N_48056);
nor U48344 (N_48344,N_48164,N_48085);
and U48345 (N_48345,N_48004,N_48039);
nor U48346 (N_48346,N_48203,N_48194);
or U48347 (N_48347,N_48062,N_48133);
and U48348 (N_48348,N_48157,N_48082);
or U48349 (N_48349,N_48217,N_48045);
nand U48350 (N_48350,N_48059,N_48118);
or U48351 (N_48351,N_48244,N_48182);
or U48352 (N_48352,N_48111,N_48154);
nand U48353 (N_48353,N_48077,N_48028);
nand U48354 (N_48354,N_48249,N_48187);
nand U48355 (N_48355,N_48209,N_48020);
or U48356 (N_48356,N_48023,N_48033);
xnor U48357 (N_48357,N_48072,N_48221);
and U48358 (N_48358,N_48215,N_48147);
or U48359 (N_48359,N_48080,N_48211);
or U48360 (N_48360,N_48216,N_48014);
xnor U48361 (N_48361,N_48109,N_48103);
nand U48362 (N_48362,N_48148,N_48019);
nor U48363 (N_48363,N_48022,N_48141);
nand U48364 (N_48364,N_48095,N_48000);
nor U48365 (N_48365,N_48012,N_48099);
and U48366 (N_48366,N_48105,N_48197);
xor U48367 (N_48367,N_48145,N_48006);
nor U48368 (N_48368,N_48002,N_48051);
xor U48369 (N_48369,N_48198,N_48223);
nor U48370 (N_48370,N_48114,N_48030);
xnor U48371 (N_48371,N_48206,N_48161);
or U48372 (N_48372,N_48008,N_48183);
and U48373 (N_48373,N_48034,N_48143);
or U48374 (N_48374,N_48200,N_48007);
or U48375 (N_48375,N_48064,N_48174);
xnor U48376 (N_48376,N_48021,N_48005);
nor U48377 (N_48377,N_48115,N_48107);
nor U48378 (N_48378,N_48138,N_48131);
nand U48379 (N_48379,N_48083,N_48024);
and U48380 (N_48380,N_48226,N_48245);
nand U48381 (N_48381,N_48040,N_48162);
and U48382 (N_48382,N_48226,N_48164);
or U48383 (N_48383,N_48159,N_48242);
xnor U48384 (N_48384,N_48180,N_48070);
and U48385 (N_48385,N_48037,N_48072);
nor U48386 (N_48386,N_48081,N_48046);
or U48387 (N_48387,N_48223,N_48038);
nor U48388 (N_48388,N_48070,N_48172);
xor U48389 (N_48389,N_48169,N_48218);
and U48390 (N_48390,N_48169,N_48244);
or U48391 (N_48391,N_48203,N_48231);
or U48392 (N_48392,N_48043,N_48009);
xor U48393 (N_48393,N_48244,N_48127);
nand U48394 (N_48394,N_48184,N_48135);
xor U48395 (N_48395,N_48018,N_48249);
and U48396 (N_48396,N_48158,N_48127);
xnor U48397 (N_48397,N_48047,N_48139);
or U48398 (N_48398,N_48200,N_48193);
nand U48399 (N_48399,N_48049,N_48225);
and U48400 (N_48400,N_48053,N_48240);
xor U48401 (N_48401,N_48082,N_48061);
and U48402 (N_48402,N_48134,N_48207);
and U48403 (N_48403,N_48119,N_48016);
nor U48404 (N_48404,N_48167,N_48007);
or U48405 (N_48405,N_48149,N_48244);
nand U48406 (N_48406,N_48086,N_48036);
nand U48407 (N_48407,N_48099,N_48132);
nand U48408 (N_48408,N_48230,N_48029);
xor U48409 (N_48409,N_48210,N_48244);
or U48410 (N_48410,N_48074,N_48039);
or U48411 (N_48411,N_48117,N_48158);
or U48412 (N_48412,N_48229,N_48172);
and U48413 (N_48413,N_48106,N_48006);
and U48414 (N_48414,N_48096,N_48123);
or U48415 (N_48415,N_48139,N_48101);
nor U48416 (N_48416,N_48222,N_48106);
nand U48417 (N_48417,N_48140,N_48211);
nor U48418 (N_48418,N_48184,N_48246);
nand U48419 (N_48419,N_48162,N_48037);
nand U48420 (N_48420,N_48189,N_48188);
nor U48421 (N_48421,N_48113,N_48243);
nor U48422 (N_48422,N_48052,N_48239);
or U48423 (N_48423,N_48187,N_48113);
nand U48424 (N_48424,N_48175,N_48181);
nand U48425 (N_48425,N_48064,N_48028);
or U48426 (N_48426,N_48197,N_48080);
and U48427 (N_48427,N_48236,N_48105);
and U48428 (N_48428,N_48030,N_48043);
nor U48429 (N_48429,N_48080,N_48051);
xnor U48430 (N_48430,N_48048,N_48160);
xnor U48431 (N_48431,N_48013,N_48060);
nand U48432 (N_48432,N_48194,N_48244);
xor U48433 (N_48433,N_48158,N_48093);
and U48434 (N_48434,N_48242,N_48204);
nand U48435 (N_48435,N_48111,N_48242);
nand U48436 (N_48436,N_48132,N_48047);
xnor U48437 (N_48437,N_48205,N_48183);
xor U48438 (N_48438,N_48179,N_48027);
or U48439 (N_48439,N_48165,N_48159);
and U48440 (N_48440,N_48206,N_48246);
nor U48441 (N_48441,N_48204,N_48166);
or U48442 (N_48442,N_48189,N_48174);
or U48443 (N_48443,N_48139,N_48030);
or U48444 (N_48444,N_48072,N_48090);
nor U48445 (N_48445,N_48087,N_48029);
nand U48446 (N_48446,N_48177,N_48110);
or U48447 (N_48447,N_48242,N_48068);
and U48448 (N_48448,N_48114,N_48015);
nor U48449 (N_48449,N_48134,N_48163);
nor U48450 (N_48450,N_48008,N_48174);
or U48451 (N_48451,N_48035,N_48123);
xnor U48452 (N_48452,N_48120,N_48015);
nand U48453 (N_48453,N_48109,N_48047);
nand U48454 (N_48454,N_48213,N_48003);
and U48455 (N_48455,N_48165,N_48214);
xnor U48456 (N_48456,N_48147,N_48176);
and U48457 (N_48457,N_48218,N_48228);
nand U48458 (N_48458,N_48004,N_48082);
xor U48459 (N_48459,N_48037,N_48120);
nand U48460 (N_48460,N_48118,N_48160);
nor U48461 (N_48461,N_48012,N_48163);
nand U48462 (N_48462,N_48020,N_48192);
nand U48463 (N_48463,N_48038,N_48152);
xor U48464 (N_48464,N_48213,N_48072);
xnor U48465 (N_48465,N_48173,N_48057);
or U48466 (N_48466,N_48207,N_48099);
and U48467 (N_48467,N_48075,N_48086);
xnor U48468 (N_48468,N_48139,N_48127);
nand U48469 (N_48469,N_48135,N_48106);
nor U48470 (N_48470,N_48230,N_48185);
nand U48471 (N_48471,N_48077,N_48092);
nor U48472 (N_48472,N_48040,N_48136);
or U48473 (N_48473,N_48011,N_48081);
or U48474 (N_48474,N_48207,N_48160);
xnor U48475 (N_48475,N_48202,N_48104);
or U48476 (N_48476,N_48061,N_48055);
or U48477 (N_48477,N_48065,N_48125);
and U48478 (N_48478,N_48146,N_48110);
nor U48479 (N_48479,N_48152,N_48077);
or U48480 (N_48480,N_48156,N_48239);
nor U48481 (N_48481,N_48247,N_48108);
and U48482 (N_48482,N_48069,N_48118);
nor U48483 (N_48483,N_48036,N_48121);
and U48484 (N_48484,N_48023,N_48043);
or U48485 (N_48485,N_48059,N_48060);
and U48486 (N_48486,N_48185,N_48202);
and U48487 (N_48487,N_48105,N_48181);
or U48488 (N_48488,N_48029,N_48246);
nand U48489 (N_48489,N_48206,N_48023);
nor U48490 (N_48490,N_48156,N_48174);
nand U48491 (N_48491,N_48058,N_48132);
and U48492 (N_48492,N_48212,N_48179);
and U48493 (N_48493,N_48099,N_48166);
xor U48494 (N_48494,N_48041,N_48150);
nor U48495 (N_48495,N_48000,N_48215);
and U48496 (N_48496,N_48044,N_48230);
xnor U48497 (N_48497,N_48020,N_48076);
and U48498 (N_48498,N_48180,N_48224);
or U48499 (N_48499,N_48169,N_48216);
nor U48500 (N_48500,N_48421,N_48455);
xor U48501 (N_48501,N_48335,N_48280);
and U48502 (N_48502,N_48487,N_48351);
or U48503 (N_48503,N_48386,N_48274);
xnor U48504 (N_48504,N_48460,N_48320);
xnor U48505 (N_48505,N_48411,N_48446);
xor U48506 (N_48506,N_48345,N_48358);
xnor U48507 (N_48507,N_48289,N_48474);
or U48508 (N_48508,N_48364,N_48251);
nand U48509 (N_48509,N_48448,N_48273);
xnor U48510 (N_48510,N_48481,N_48477);
nor U48511 (N_48511,N_48453,N_48257);
nand U48512 (N_48512,N_48388,N_48254);
xnor U48513 (N_48513,N_48431,N_48311);
xor U48514 (N_48514,N_48410,N_48301);
nand U48515 (N_48515,N_48265,N_48490);
or U48516 (N_48516,N_48295,N_48465);
or U48517 (N_48517,N_48483,N_48491);
nor U48518 (N_48518,N_48469,N_48437);
nand U48519 (N_48519,N_48258,N_48290);
nand U48520 (N_48520,N_48377,N_48312);
or U48521 (N_48521,N_48306,N_48407);
xor U48522 (N_48522,N_48489,N_48464);
nand U48523 (N_48523,N_48406,N_48346);
or U48524 (N_48524,N_48271,N_48396);
nor U48525 (N_48525,N_48359,N_48379);
nand U48526 (N_48526,N_48304,N_48409);
and U48527 (N_48527,N_48468,N_48263);
or U48528 (N_48528,N_48355,N_48319);
or U48529 (N_48529,N_48348,N_48314);
nor U48530 (N_48530,N_48292,N_48378);
nand U48531 (N_48531,N_48360,N_48447);
nand U48532 (N_48532,N_48485,N_48414);
and U48533 (N_48533,N_48401,N_48349);
xor U48534 (N_48534,N_48384,N_48370);
and U48535 (N_48535,N_48375,N_48357);
or U48536 (N_48536,N_48284,N_48342);
or U48537 (N_48537,N_48340,N_48293);
nor U48538 (N_48538,N_48374,N_48315);
nor U48539 (N_48539,N_48277,N_48253);
and U48540 (N_48540,N_48278,N_48463);
nor U48541 (N_48541,N_48443,N_48291);
nor U48542 (N_48542,N_48399,N_48405);
xor U48543 (N_48543,N_48495,N_48252);
or U48544 (N_48544,N_48478,N_48412);
or U48545 (N_48545,N_48272,N_48372);
xor U48546 (N_48546,N_48444,N_48362);
nand U48547 (N_48547,N_48452,N_48427);
xnor U48548 (N_48548,N_48492,N_48323);
xor U48549 (N_48549,N_48322,N_48339);
nor U48550 (N_48550,N_48398,N_48270);
xor U48551 (N_48551,N_48316,N_48385);
and U48552 (N_48552,N_48371,N_48425);
nand U48553 (N_48553,N_48390,N_48328);
nand U48554 (N_48554,N_48488,N_48423);
and U48555 (N_48555,N_48473,N_48420);
and U48556 (N_48556,N_48333,N_48476);
and U48557 (N_48557,N_48286,N_48461);
or U48558 (N_48558,N_48344,N_48361);
and U48559 (N_48559,N_48294,N_48300);
nor U48560 (N_48560,N_48424,N_48307);
or U48561 (N_48561,N_48445,N_48416);
nor U48562 (N_48562,N_48303,N_48264);
xor U48563 (N_48563,N_48366,N_48430);
xor U48564 (N_48564,N_48313,N_48404);
xnor U48565 (N_48565,N_48394,N_48268);
and U48566 (N_48566,N_48267,N_48347);
or U48567 (N_48567,N_48480,N_48317);
nor U48568 (N_48568,N_48305,N_48365);
nand U48569 (N_48569,N_48496,N_48353);
xor U48570 (N_48570,N_48454,N_48438);
nor U48571 (N_48571,N_48338,N_48497);
or U48572 (N_48572,N_48400,N_48299);
xor U48573 (N_48573,N_48493,N_48354);
nand U48574 (N_48574,N_48330,N_48451);
nand U48575 (N_48575,N_48415,N_48467);
or U48576 (N_48576,N_48391,N_48429);
or U48577 (N_48577,N_48288,N_48326);
nor U48578 (N_48578,N_48279,N_48392);
nand U48579 (N_48579,N_48318,N_48450);
nor U48580 (N_48580,N_48261,N_48260);
nand U48581 (N_48581,N_48442,N_48419);
nor U48582 (N_48582,N_48259,N_48285);
and U48583 (N_48583,N_48343,N_48324);
or U48584 (N_48584,N_48433,N_48486);
nor U48585 (N_48585,N_48275,N_48250);
nand U48586 (N_48586,N_48432,N_48381);
nor U48587 (N_48587,N_48352,N_48441);
nand U48588 (N_48588,N_48499,N_48276);
xor U48589 (N_48589,N_48256,N_48494);
and U48590 (N_48590,N_48393,N_48262);
or U48591 (N_48591,N_48302,N_48402);
or U48592 (N_48592,N_48321,N_48397);
nor U48593 (N_48593,N_48368,N_48403);
and U48594 (N_48594,N_48297,N_48298);
nor U48595 (N_48595,N_48466,N_48479);
nor U48596 (N_48596,N_48395,N_48434);
xnor U48597 (N_48597,N_48470,N_48331);
or U48598 (N_48598,N_48426,N_48389);
and U48599 (N_48599,N_48356,N_48281);
xnor U48600 (N_48600,N_48367,N_48337);
or U48601 (N_48601,N_48283,N_48422);
and U48602 (N_48602,N_48459,N_48449);
and U48603 (N_48603,N_48408,N_48458);
xnor U48604 (N_48604,N_48484,N_48255);
nor U48605 (N_48605,N_48336,N_48436);
or U48606 (N_48606,N_48498,N_48287);
nor U48607 (N_48607,N_48332,N_48428);
or U48608 (N_48608,N_48269,N_48309);
xor U48609 (N_48609,N_48413,N_48310);
nor U48610 (N_48610,N_48482,N_48471);
nor U48611 (N_48611,N_48383,N_48376);
or U48612 (N_48612,N_48472,N_48457);
or U48613 (N_48613,N_48435,N_48373);
or U48614 (N_48614,N_48308,N_48296);
nand U48615 (N_48615,N_48327,N_48282);
or U48616 (N_48616,N_48440,N_48439);
nor U48617 (N_48617,N_48329,N_48456);
and U48618 (N_48618,N_48387,N_48462);
and U48619 (N_48619,N_48382,N_48418);
and U48620 (N_48620,N_48363,N_48334);
nor U48621 (N_48621,N_48369,N_48417);
nand U48622 (N_48622,N_48325,N_48266);
xnor U48623 (N_48623,N_48475,N_48341);
and U48624 (N_48624,N_48380,N_48350);
or U48625 (N_48625,N_48366,N_48372);
xnor U48626 (N_48626,N_48456,N_48405);
or U48627 (N_48627,N_48433,N_48345);
and U48628 (N_48628,N_48479,N_48316);
xnor U48629 (N_48629,N_48359,N_48446);
xor U48630 (N_48630,N_48326,N_48387);
or U48631 (N_48631,N_48282,N_48315);
or U48632 (N_48632,N_48492,N_48307);
xor U48633 (N_48633,N_48370,N_48262);
xor U48634 (N_48634,N_48429,N_48465);
or U48635 (N_48635,N_48451,N_48360);
nor U48636 (N_48636,N_48337,N_48328);
and U48637 (N_48637,N_48416,N_48446);
or U48638 (N_48638,N_48381,N_48266);
xnor U48639 (N_48639,N_48291,N_48334);
xor U48640 (N_48640,N_48372,N_48297);
nand U48641 (N_48641,N_48452,N_48300);
nand U48642 (N_48642,N_48277,N_48367);
and U48643 (N_48643,N_48426,N_48460);
xor U48644 (N_48644,N_48496,N_48312);
or U48645 (N_48645,N_48377,N_48348);
xor U48646 (N_48646,N_48394,N_48332);
or U48647 (N_48647,N_48366,N_48261);
nand U48648 (N_48648,N_48340,N_48255);
nand U48649 (N_48649,N_48426,N_48367);
and U48650 (N_48650,N_48361,N_48447);
or U48651 (N_48651,N_48353,N_48461);
and U48652 (N_48652,N_48474,N_48257);
nor U48653 (N_48653,N_48450,N_48350);
xor U48654 (N_48654,N_48365,N_48433);
or U48655 (N_48655,N_48350,N_48381);
and U48656 (N_48656,N_48313,N_48357);
nand U48657 (N_48657,N_48288,N_48273);
nor U48658 (N_48658,N_48380,N_48393);
or U48659 (N_48659,N_48252,N_48295);
and U48660 (N_48660,N_48333,N_48468);
nand U48661 (N_48661,N_48358,N_48400);
xnor U48662 (N_48662,N_48297,N_48299);
or U48663 (N_48663,N_48373,N_48492);
xnor U48664 (N_48664,N_48284,N_48373);
or U48665 (N_48665,N_48332,N_48426);
nor U48666 (N_48666,N_48410,N_48390);
nand U48667 (N_48667,N_48378,N_48379);
or U48668 (N_48668,N_48360,N_48300);
nor U48669 (N_48669,N_48306,N_48418);
xor U48670 (N_48670,N_48343,N_48431);
and U48671 (N_48671,N_48381,N_48326);
and U48672 (N_48672,N_48409,N_48437);
and U48673 (N_48673,N_48477,N_48393);
and U48674 (N_48674,N_48388,N_48402);
and U48675 (N_48675,N_48348,N_48316);
and U48676 (N_48676,N_48411,N_48404);
nor U48677 (N_48677,N_48423,N_48363);
xnor U48678 (N_48678,N_48271,N_48487);
xnor U48679 (N_48679,N_48336,N_48406);
or U48680 (N_48680,N_48304,N_48275);
nand U48681 (N_48681,N_48386,N_48344);
and U48682 (N_48682,N_48348,N_48424);
and U48683 (N_48683,N_48354,N_48253);
nor U48684 (N_48684,N_48484,N_48312);
or U48685 (N_48685,N_48379,N_48381);
or U48686 (N_48686,N_48329,N_48479);
nor U48687 (N_48687,N_48382,N_48324);
xnor U48688 (N_48688,N_48371,N_48333);
nor U48689 (N_48689,N_48290,N_48438);
nor U48690 (N_48690,N_48390,N_48321);
nor U48691 (N_48691,N_48470,N_48371);
nor U48692 (N_48692,N_48349,N_48375);
xnor U48693 (N_48693,N_48263,N_48442);
or U48694 (N_48694,N_48272,N_48251);
nand U48695 (N_48695,N_48486,N_48344);
and U48696 (N_48696,N_48417,N_48352);
or U48697 (N_48697,N_48305,N_48383);
or U48698 (N_48698,N_48291,N_48499);
xnor U48699 (N_48699,N_48441,N_48417);
and U48700 (N_48700,N_48285,N_48424);
nand U48701 (N_48701,N_48331,N_48315);
nor U48702 (N_48702,N_48394,N_48493);
xor U48703 (N_48703,N_48433,N_48459);
xor U48704 (N_48704,N_48300,N_48354);
nand U48705 (N_48705,N_48388,N_48427);
or U48706 (N_48706,N_48273,N_48497);
and U48707 (N_48707,N_48257,N_48262);
nor U48708 (N_48708,N_48278,N_48316);
nor U48709 (N_48709,N_48334,N_48461);
nor U48710 (N_48710,N_48412,N_48295);
nand U48711 (N_48711,N_48302,N_48468);
nor U48712 (N_48712,N_48339,N_48380);
or U48713 (N_48713,N_48464,N_48392);
xor U48714 (N_48714,N_48255,N_48257);
nor U48715 (N_48715,N_48255,N_48366);
xnor U48716 (N_48716,N_48365,N_48436);
nand U48717 (N_48717,N_48476,N_48491);
and U48718 (N_48718,N_48413,N_48442);
and U48719 (N_48719,N_48499,N_48402);
or U48720 (N_48720,N_48315,N_48334);
nand U48721 (N_48721,N_48294,N_48376);
xnor U48722 (N_48722,N_48309,N_48325);
nand U48723 (N_48723,N_48294,N_48307);
or U48724 (N_48724,N_48267,N_48414);
and U48725 (N_48725,N_48446,N_48406);
nand U48726 (N_48726,N_48348,N_48360);
xor U48727 (N_48727,N_48495,N_48319);
nand U48728 (N_48728,N_48414,N_48304);
xnor U48729 (N_48729,N_48456,N_48413);
and U48730 (N_48730,N_48265,N_48298);
xnor U48731 (N_48731,N_48427,N_48499);
nor U48732 (N_48732,N_48453,N_48403);
nand U48733 (N_48733,N_48297,N_48487);
nand U48734 (N_48734,N_48326,N_48347);
xnor U48735 (N_48735,N_48276,N_48496);
nor U48736 (N_48736,N_48337,N_48293);
xnor U48737 (N_48737,N_48461,N_48322);
or U48738 (N_48738,N_48458,N_48486);
and U48739 (N_48739,N_48415,N_48435);
and U48740 (N_48740,N_48354,N_48385);
nand U48741 (N_48741,N_48480,N_48469);
and U48742 (N_48742,N_48381,N_48331);
and U48743 (N_48743,N_48499,N_48350);
nor U48744 (N_48744,N_48268,N_48381);
nand U48745 (N_48745,N_48385,N_48446);
nand U48746 (N_48746,N_48423,N_48309);
nand U48747 (N_48747,N_48426,N_48335);
nand U48748 (N_48748,N_48267,N_48443);
xnor U48749 (N_48749,N_48375,N_48346);
xor U48750 (N_48750,N_48502,N_48511);
xnor U48751 (N_48751,N_48659,N_48707);
and U48752 (N_48752,N_48570,N_48718);
nand U48753 (N_48753,N_48616,N_48706);
and U48754 (N_48754,N_48557,N_48742);
nand U48755 (N_48755,N_48641,N_48602);
nand U48756 (N_48756,N_48547,N_48552);
nand U48757 (N_48757,N_48627,N_48636);
or U48758 (N_48758,N_48509,N_48522);
nand U48759 (N_48759,N_48671,N_48741);
or U48760 (N_48760,N_48617,N_48716);
nand U48761 (N_48761,N_48505,N_48739);
and U48762 (N_48762,N_48645,N_48691);
or U48763 (N_48763,N_48536,N_48626);
xor U48764 (N_48764,N_48577,N_48532);
or U48765 (N_48765,N_48589,N_48693);
nand U48766 (N_48766,N_48531,N_48567);
and U48767 (N_48767,N_48639,N_48647);
nand U48768 (N_48768,N_48587,N_48580);
nand U48769 (N_48769,N_48603,N_48523);
nand U48770 (N_48770,N_48652,N_48649);
nand U48771 (N_48771,N_48554,N_48670);
and U48772 (N_48772,N_48528,N_48729);
or U48773 (N_48773,N_48747,N_48572);
and U48774 (N_48774,N_48703,N_48614);
and U48775 (N_48775,N_48598,N_48732);
xor U48776 (N_48776,N_48543,N_48500);
nand U48777 (N_48777,N_48524,N_48512);
nand U48778 (N_48778,N_48721,N_48573);
xor U48779 (N_48779,N_48674,N_48749);
or U48780 (N_48780,N_48628,N_48593);
and U48781 (N_48781,N_48658,N_48665);
nand U48782 (N_48782,N_48646,N_48591);
nand U48783 (N_48783,N_48681,N_48513);
or U48784 (N_48784,N_48568,N_48700);
xor U48785 (N_48785,N_48668,N_48734);
or U48786 (N_48786,N_48596,N_48613);
nor U48787 (N_48787,N_48683,N_48661);
or U48788 (N_48788,N_48560,N_48530);
nor U48789 (N_48789,N_48583,N_48704);
and U48790 (N_48790,N_48669,N_48542);
and U48791 (N_48791,N_48604,N_48605);
or U48792 (N_48792,N_48642,N_48620);
and U48793 (N_48793,N_48728,N_48526);
or U48794 (N_48794,N_48623,N_48534);
nand U48795 (N_48795,N_48566,N_48680);
or U48796 (N_48796,N_48651,N_48735);
nor U48797 (N_48797,N_48631,N_48696);
or U48798 (N_48798,N_48687,N_48684);
nor U48799 (N_48799,N_48612,N_48615);
xor U48800 (N_48800,N_48551,N_48719);
nand U48801 (N_48801,N_48535,N_48584);
xor U48802 (N_48802,N_48515,N_48638);
nand U48803 (N_48803,N_48541,N_48692);
and U48804 (N_48804,N_48608,N_48730);
xor U48805 (N_48805,N_48519,N_48640);
nor U48806 (N_48806,N_48514,N_48621);
nor U48807 (N_48807,N_48607,N_48571);
nand U48808 (N_48808,N_48624,N_48632);
nor U48809 (N_48809,N_48697,N_48501);
xnor U48810 (N_48810,N_48743,N_48520);
nand U48811 (N_48811,N_48618,N_48690);
or U48812 (N_48812,N_48565,N_48675);
and U48813 (N_48813,N_48725,N_48548);
or U48814 (N_48814,N_48699,N_48678);
nor U48815 (N_48815,N_48525,N_48714);
nor U48816 (N_48816,N_48654,N_48731);
nand U48817 (N_48817,N_48510,N_48679);
and U48818 (N_48818,N_48722,N_48744);
and U48819 (N_48819,N_48685,N_48736);
nand U48820 (N_48820,N_48702,N_48601);
nor U48821 (N_48821,N_48698,N_48677);
or U48822 (N_48822,N_48676,N_48592);
or U48823 (N_48823,N_48713,N_48715);
xor U48824 (N_48824,N_48569,N_48561);
or U48825 (N_48825,N_48517,N_48701);
nor U48826 (N_48826,N_48663,N_48610);
nor U48827 (N_48827,N_48644,N_48694);
nor U48828 (N_48828,N_48746,N_48667);
and U48829 (N_48829,N_48656,N_48559);
nor U48830 (N_48830,N_48720,N_48594);
nand U48831 (N_48831,N_48507,N_48688);
nand U48832 (N_48832,N_48586,N_48549);
nor U48833 (N_48833,N_48650,N_48562);
nand U48834 (N_48834,N_48558,N_48733);
nand U48835 (N_48835,N_48686,N_48712);
and U48836 (N_48836,N_48553,N_48695);
and U48837 (N_48837,N_48504,N_48539);
nor U48838 (N_48838,N_48506,N_48611);
nor U48839 (N_48839,N_48738,N_48574);
and U48840 (N_48840,N_48748,N_48556);
and U48841 (N_48841,N_48546,N_48563);
nor U48842 (N_48842,N_48582,N_48588);
or U48843 (N_48843,N_48516,N_48662);
and U48844 (N_48844,N_48708,N_48527);
nand U48845 (N_48845,N_48609,N_48625);
nor U48846 (N_48846,N_48666,N_48745);
or U48847 (N_48847,N_48633,N_48619);
xnor U48848 (N_48848,N_48710,N_48564);
nor U48849 (N_48849,N_48724,N_48637);
xnor U48850 (N_48850,N_48629,N_48597);
and U48851 (N_48851,N_48622,N_48585);
and U48852 (N_48852,N_48705,N_48682);
nor U48853 (N_48853,N_48655,N_48657);
and U48854 (N_48854,N_48643,N_48575);
xor U48855 (N_48855,N_48538,N_48664);
nor U48856 (N_48856,N_48576,N_48634);
xnor U48857 (N_48857,N_48673,N_48660);
nor U48858 (N_48858,N_48689,N_48595);
xnor U48859 (N_48859,N_48599,N_48717);
nor U48860 (N_48860,N_48521,N_48540);
nand U48861 (N_48861,N_48709,N_48550);
and U48862 (N_48862,N_48579,N_48740);
and U48863 (N_48863,N_48544,N_48503);
and U48864 (N_48864,N_48581,N_48606);
xnor U48865 (N_48865,N_48537,N_48545);
nor U48866 (N_48866,N_48578,N_48630);
xnor U48867 (N_48867,N_48600,N_48529);
nand U48868 (N_48868,N_48711,N_48737);
xnor U48869 (N_48869,N_48555,N_48672);
xnor U48870 (N_48870,N_48590,N_48726);
nand U48871 (N_48871,N_48533,N_48723);
nor U48872 (N_48872,N_48635,N_48518);
or U48873 (N_48873,N_48727,N_48648);
nor U48874 (N_48874,N_48508,N_48653);
xor U48875 (N_48875,N_48543,N_48687);
nand U48876 (N_48876,N_48509,N_48545);
xnor U48877 (N_48877,N_48538,N_48616);
or U48878 (N_48878,N_48703,N_48574);
xnor U48879 (N_48879,N_48586,N_48621);
xor U48880 (N_48880,N_48622,N_48745);
xor U48881 (N_48881,N_48660,N_48696);
and U48882 (N_48882,N_48519,N_48683);
nor U48883 (N_48883,N_48597,N_48689);
and U48884 (N_48884,N_48597,N_48711);
nand U48885 (N_48885,N_48667,N_48618);
or U48886 (N_48886,N_48538,N_48703);
and U48887 (N_48887,N_48680,N_48737);
nand U48888 (N_48888,N_48626,N_48578);
xor U48889 (N_48889,N_48736,N_48658);
and U48890 (N_48890,N_48735,N_48618);
and U48891 (N_48891,N_48560,N_48548);
and U48892 (N_48892,N_48646,N_48568);
and U48893 (N_48893,N_48626,N_48554);
and U48894 (N_48894,N_48718,N_48682);
xor U48895 (N_48895,N_48614,N_48570);
nand U48896 (N_48896,N_48523,N_48672);
and U48897 (N_48897,N_48735,N_48598);
or U48898 (N_48898,N_48591,N_48630);
nor U48899 (N_48899,N_48674,N_48725);
nor U48900 (N_48900,N_48538,N_48712);
or U48901 (N_48901,N_48718,N_48553);
and U48902 (N_48902,N_48517,N_48714);
nand U48903 (N_48903,N_48538,N_48559);
nor U48904 (N_48904,N_48541,N_48581);
or U48905 (N_48905,N_48716,N_48561);
xnor U48906 (N_48906,N_48642,N_48732);
or U48907 (N_48907,N_48592,N_48738);
and U48908 (N_48908,N_48542,N_48511);
and U48909 (N_48909,N_48557,N_48721);
and U48910 (N_48910,N_48635,N_48667);
xnor U48911 (N_48911,N_48547,N_48698);
nor U48912 (N_48912,N_48658,N_48696);
nor U48913 (N_48913,N_48501,N_48725);
or U48914 (N_48914,N_48577,N_48631);
nor U48915 (N_48915,N_48648,N_48507);
nor U48916 (N_48916,N_48550,N_48538);
or U48917 (N_48917,N_48724,N_48622);
and U48918 (N_48918,N_48535,N_48597);
xnor U48919 (N_48919,N_48564,N_48731);
nor U48920 (N_48920,N_48580,N_48600);
nand U48921 (N_48921,N_48648,N_48664);
or U48922 (N_48922,N_48695,N_48621);
nand U48923 (N_48923,N_48569,N_48730);
nor U48924 (N_48924,N_48673,N_48523);
and U48925 (N_48925,N_48568,N_48624);
and U48926 (N_48926,N_48718,N_48540);
or U48927 (N_48927,N_48710,N_48684);
xor U48928 (N_48928,N_48699,N_48646);
nand U48929 (N_48929,N_48659,N_48682);
nand U48930 (N_48930,N_48625,N_48724);
nand U48931 (N_48931,N_48606,N_48648);
nand U48932 (N_48932,N_48724,N_48711);
or U48933 (N_48933,N_48633,N_48671);
and U48934 (N_48934,N_48703,N_48526);
nor U48935 (N_48935,N_48681,N_48685);
nor U48936 (N_48936,N_48542,N_48644);
and U48937 (N_48937,N_48682,N_48749);
nand U48938 (N_48938,N_48731,N_48709);
nor U48939 (N_48939,N_48714,N_48632);
nand U48940 (N_48940,N_48583,N_48655);
and U48941 (N_48941,N_48704,N_48553);
nor U48942 (N_48942,N_48505,N_48689);
and U48943 (N_48943,N_48573,N_48725);
nand U48944 (N_48944,N_48731,N_48685);
xnor U48945 (N_48945,N_48720,N_48691);
and U48946 (N_48946,N_48714,N_48697);
or U48947 (N_48947,N_48627,N_48568);
nand U48948 (N_48948,N_48623,N_48523);
nor U48949 (N_48949,N_48512,N_48505);
and U48950 (N_48950,N_48705,N_48555);
xnor U48951 (N_48951,N_48618,N_48526);
nor U48952 (N_48952,N_48521,N_48652);
or U48953 (N_48953,N_48652,N_48593);
and U48954 (N_48954,N_48528,N_48721);
xor U48955 (N_48955,N_48576,N_48685);
and U48956 (N_48956,N_48734,N_48726);
and U48957 (N_48957,N_48745,N_48555);
xnor U48958 (N_48958,N_48599,N_48747);
and U48959 (N_48959,N_48526,N_48646);
xor U48960 (N_48960,N_48616,N_48622);
nand U48961 (N_48961,N_48667,N_48649);
and U48962 (N_48962,N_48516,N_48520);
xor U48963 (N_48963,N_48550,N_48743);
or U48964 (N_48964,N_48518,N_48521);
and U48965 (N_48965,N_48540,N_48574);
xor U48966 (N_48966,N_48600,N_48678);
and U48967 (N_48967,N_48689,N_48706);
xor U48968 (N_48968,N_48706,N_48529);
or U48969 (N_48969,N_48737,N_48571);
nor U48970 (N_48970,N_48597,N_48536);
xor U48971 (N_48971,N_48529,N_48748);
or U48972 (N_48972,N_48714,N_48586);
xor U48973 (N_48973,N_48700,N_48741);
xor U48974 (N_48974,N_48538,N_48576);
nor U48975 (N_48975,N_48689,N_48575);
and U48976 (N_48976,N_48711,N_48695);
or U48977 (N_48977,N_48594,N_48655);
nand U48978 (N_48978,N_48737,N_48513);
xor U48979 (N_48979,N_48595,N_48641);
or U48980 (N_48980,N_48712,N_48621);
nand U48981 (N_48981,N_48653,N_48574);
xnor U48982 (N_48982,N_48603,N_48563);
xnor U48983 (N_48983,N_48529,N_48746);
xnor U48984 (N_48984,N_48730,N_48537);
or U48985 (N_48985,N_48709,N_48524);
xor U48986 (N_48986,N_48663,N_48669);
nand U48987 (N_48987,N_48511,N_48658);
xor U48988 (N_48988,N_48740,N_48732);
nor U48989 (N_48989,N_48510,N_48657);
nand U48990 (N_48990,N_48629,N_48653);
nor U48991 (N_48991,N_48580,N_48643);
nor U48992 (N_48992,N_48528,N_48585);
nor U48993 (N_48993,N_48529,N_48715);
nor U48994 (N_48994,N_48605,N_48740);
and U48995 (N_48995,N_48522,N_48702);
and U48996 (N_48996,N_48609,N_48629);
xor U48997 (N_48997,N_48731,N_48599);
xor U48998 (N_48998,N_48517,N_48744);
and U48999 (N_48999,N_48627,N_48679);
nor U49000 (N_49000,N_48964,N_48784);
nor U49001 (N_49001,N_48812,N_48882);
and U49002 (N_49002,N_48813,N_48931);
or U49003 (N_49003,N_48835,N_48766);
and U49004 (N_49004,N_48963,N_48988);
or U49005 (N_49005,N_48929,N_48751);
and U49006 (N_49006,N_48854,N_48786);
nor U49007 (N_49007,N_48885,N_48891);
or U49008 (N_49008,N_48969,N_48905);
xnor U49009 (N_49009,N_48955,N_48761);
xor U49010 (N_49010,N_48961,N_48933);
nor U49011 (N_49011,N_48825,N_48972);
or U49012 (N_49012,N_48886,N_48977);
nor U49013 (N_49013,N_48934,N_48992);
nor U49014 (N_49014,N_48960,N_48864);
nand U49015 (N_49015,N_48878,N_48903);
xor U49016 (N_49016,N_48899,N_48846);
nand U49017 (N_49017,N_48954,N_48803);
and U49018 (N_49018,N_48862,N_48881);
and U49019 (N_49019,N_48917,N_48827);
nor U49020 (N_49020,N_48858,N_48884);
and U49021 (N_49021,N_48795,N_48853);
xor U49022 (N_49022,N_48906,N_48937);
xor U49023 (N_49023,N_48781,N_48856);
and U49024 (N_49024,N_48898,N_48867);
nor U49025 (N_49025,N_48798,N_48975);
and U49026 (N_49026,N_48945,N_48815);
or U49027 (N_49027,N_48894,N_48752);
or U49028 (N_49028,N_48998,N_48774);
nand U49029 (N_49029,N_48987,N_48783);
nand U49030 (N_49030,N_48978,N_48926);
nand U49031 (N_49031,N_48847,N_48757);
or U49032 (N_49032,N_48799,N_48822);
nand U49033 (N_49033,N_48823,N_48957);
and U49034 (N_49034,N_48909,N_48772);
nand U49035 (N_49035,N_48792,N_48838);
nor U49036 (N_49036,N_48765,N_48984);
and U49037 (N_49037,N_48908,N_48950);
and U49038 (N_49038,N_48956,N_48900);
nand U49039 (N_49039,N_48880,N_48875);
nand U49040 (N_49040,N_48976,N_48986);
nand U49041 (N_49041,N_48851,N_48943);
nor U49042 (N_49042,N_48840,N_48893);
xnor U49043 (N_49043,N_48990,N_48915);
or U49044 (N_49044,N_48768,N_48912);
xnor U49045 (N_49045,N_48980,N_48859);
and U49046 (N_49046,N_48802,N_48763);
xnor U49047 (N_49047,N_48979,N_48932);
and U49048 (N_49048,N_48800,N_48850);
and U49049 (N_49049,N_48995,N_48806);
nor U49050 (N_49050,N_48868,N_48902);
nor U49051 (N_49051,N_48824,N_48767);
nand U49052 (N_49052,N_48845,N_48778);
or U49053 (N_49053,N_48753,N_48870);
xnor U49054 (N_49054,N_48994,N_48951);
xnor U49055 (N_49055,N_48920,N_48936);
and U49056 (N_49056,N_48836,N_48892);
xor U49057 (N_49057,N_48958,N_48923);
or U49058 (N_49058,N_48816,N_48832);
and U49059 (N_49059,N_48811,N_48764);
xnor U49060 (N_49060,N_48996,N_48791);
and U49061 (N_49061,N_48896,N_48971);
xnor U49062 (N_49062,N_48843,N_48805);
nor U49063 (N_49063,N_48948,N_48769);
xor U49064 (N_49064,N_48944,N_48946);
nand U49065 (N_49065,N_48965,N_48949);
nor U49066 (N_49066,N_48930,N_48844);
nor U49067 (N_49067,N_48889,N_48869);
nand U49068 (N_49068,N_48871,N_48999);
nor U49069 (N_49069,N_48826,N_48833);
or U49070 (N_49070,N_48983,N_48848);
xor U49071 (N_49071,N_48834,N_48872);
or U49072 (N_49072,N_48907,N_48782);
nand U49073 (N_49073,N_48777,N_48967);
and U49074 (N_49074,N_48829,N_48918);
nand U49075 (N_49075,N_48922,N_48762);
nor U49076 (N_49076,N_48861,N_48921);
or U49077 (N_49077,N_48993,N_48857);
xor U49078 (N_49078,N_48952,N_48750);
xor U49079 (N_49079,N_48897,N_48962);
or U49080 (N_49080,N_48797,N_48855);
nand U49081 (N_49081,N_48860,N_48814);
nand U49082 (N_49082,N_48997,N_48793);
and U49083 (N_49083,N_48953,N_48818);
or U49084 (N_49084,N_48991,N_48925);
nand U49085 (N_49085,N_48947,N_48817);
xnor U49086 (N_49086,N_48890,N_48901);
nand U49087 (N_49087,N_48935,N_48831);
xnor U49088 (N_49088,N_48830,N_48873);
nor U49089 (N_49089,N_48879,N_48910);
and U49090 (N_49090,N_48974,N_48941);
xnor U49091 (N_49091,N_48924,N_48959);
or U49092 (N_49092,N_48771,N_48982);
xor U49093 (N_49093,N_48787,N_48779);
nor U49094 (N_49094,N_48754,N_48809);
xnor U49095 (N_49095,N_48914,N_48866);
xnor U49096 (N_49096,N_48940,N_48810);
or U49097 (N_49097,N_48852,N_48849);
nand U49098 (N_49098,N_48780,N_48928);
or U49099 (N_49099,N_48942,N_48916);
nor U49100 (N_49100,N_48760,N_48756);
xnor U49101 (N_49101,N_48865,N_48821);
or U49102 (N_49102,N_48785,N_48876);
nand U49103 (N_49103,N_48755,N_48841);
and U49104 (N_49104,N_48801,N_48913);
xor U49105 (N_49105,N_48895,N_48919);
nand U49106 (N_49106,N_48773,N_48939);
nand U49107 (N_49107,N_48790,N_48842);
or U49108 (N_49108,N_48828,N_48775);
nor U49109 (N_49109,N_48927,N_48883);
or U49110 (N_49110,N_48808,N_48759);
nor U49111 (N_49111,N_48758,N_48888);
nand U49112 (N_49112,N_48877,N_48904);
and U49113 (N_49113,N_48837,N_48794);
nand U49114 (N_49114,N_48911,N_48887);
and U49115 (N_49115,N_48819,N_48968);
xnor U49116 (N_49116,N_48985,N_48820);
xor U49117 (N_49117,N_48973,N_48804);
or U49118 (N_49118,N_48981,N_48796);
xnor U49119 (N_49119,N_48776,N_48863);
xor U49120 (N_49120,N_48938,N_48789);
or U49121 (N_49121,N_48966,N_48770);
or U49122 (N_49122,N_48989,N_48874);
xor U49123 (N_49123,N_48839,N_48970);
and U49124 (N_49124,N_48788,N_48807);
and U49125 (N_49125,N_48796,N_48961);
xor U49126 (N_49126,N_48938,N_48996);
or U49127 (N_49127,N_48842,N_48890);
nor U49128 (N_49128,N_48991,N_48963);
and U49129 (N_49129,N_48873,N_48954);
or U49130 (N_49130,N_48944,N_48839);
nand U49131 (N_49131,N_48852,N_48782);
xor U49132 (N_49132,N_48794,N_48959);
nor U49133 (N_49133,N_48974,N_48839);
and U49134 (N_49134,N_48997,N_48758);
or U49135 (N_49135,N_48766,N_48839);
xor U49136 (N_49136,N_48939,N_48957);
or U49137 (N_49137,N_48909,N_48851);
xnor U49138 (N_49138,N_48872,N_48994);
nor U49139 (N_49139,N_48963,N_48823);
nand U49140 (N_49140,N_48789,N_48754);
xnor U49141 (N_49141,N_48974,N_48805);
nor U49142 (N_49142,N_48865,N_48784);
and U49143 (N_49143,N_48906,N_48779);
nor U49144 (N_49144,N_48771,N_48992);
and U49145 (N_49145,N_48822,N_48859);
nand U49146 (N_49146,N_48953,N_48839);
nand U49147 (N_49147,N_48980,N_48922);
nand U49148 (N_49148,N_48886,N_48801);
xor U49149 (N_49149,N_48769,N_48868);
and U49150 (N_49150,N_48772,N_48890);
nor U49151 (N_49151,N_48984,N_48980);
nor U49152 (N_49152,N_48823,N_48857);
nor U49153 (N_49153,N_48891,N_48853);
nand U49154 (N_49154,N_48772,N_48826);
nor U49155 (N_49155,N_48991,N_48798);
and U49156 (N_49156,N_48985,N_48858);
or U49157 (N_49157,N_48940,N_48750);
or U49158 (N_49158,N_48770,N_48963);
and U49159 (N_49159,N_48976,N_48970);
xnor U49160 (N_49160,N_48805,N_48991);
nor U49161 (N_49161,N_48751,N_48852);
and U49162 (N_49162,N_48835,N_48790);
nand U49163 (N_49163,N_48829,N_48962);
nand U49164 (N_49164,N_48781,N_48811);
nor U49165 (N_49165,N_48861,N_48810);
xor U49166 (N_49166,N_48783,N_48756);
nor U49167 (N_49167,N_48814,N_48929);
nor U49168 (N_49168,N_48817,N_48804);
nor U49169 (N_49169,N_48900,N_48962);
xnor U49170 (N_49170,N_48879,N_48984);
and U49171 (N_49171,N_48897,N_48825);
and U49172 (N_49172,N_48931,N_48840);
nor U49173 (N_49173,N_48753,N_48875);
and U49174 (N_49174,N_48838,N_48770);
xnor U49175 (N_49175,N_48935,N_48784);
xor U49176 (N_49176,N_48861,N_48912);
and U49177 (N_49177,N_48854,N_48880);
xor U49178 (N_49178,N_48837,N_48978);
and U49179 (N_49179,N_48809,N_48914);
xnor U49180 (N_49180,N_48880,N_48802);
nand U49181 (N_49181,N_48975,N_48815);
nor U49182 (N_49182,N_48828,N_48766);
and U49183 (N_49183,N_48812,N_48815);
and U49184 (N_49184,N_48963,N_48959);
xnor U49185 (N_49185,N_48889,N_48959);
nor U49186 (N_49186,N_48951,N_48913);
xnor U49187 (N_49187,N_48915,N_48967);
and U49188 (N_49188,N_48893,N_48873);
nand U49189 (N_49189,N_48757,N_48936);
nor U49190 (N_49190,N_48987,N_48907);
and U49191 (N_49191,N_48938,N_48962);
nor U49192 (N_49192,N_48955,N_48919);
nand U49193 (N_49193,N_48757,N_48859);
nor U49194 (N_49194,N_48756,N_48896);
nor U49195 (N_49195,N_48834,N_48883);
xor U49196 (N_49196,N_48936,N_48961);
or U49197 (N_49197,N_48761,N_48772);
xnor U49198 (N_49198,N_48933,N_48798);
nand U49199 (N_49199,N_48984,N_48782);
and U49200 (N_49200,N_48890,N_48943);
nor U49201 (N_49201,N_48862,N_48878);
xnor U49202 (N_49202,N_48767,N_48965);
and U49203 (N_49203,N_48819,N_48889);
nand U49204 (N_49204,N_48777,N_48894);
nand U49205 (N_49205,N_48894,N_48788);
and U49206 (N_49206,N_48765,N_48813);
xnor U49207 (N_49207,N_48943,N_48797);
and U49208 (N_49208,N_48892,N_48831);
and U49209 (N_49209,N_48924,N_48975);
nand U49210 (N_49210,N_48920,N_48824);
and U49211 (N_49211,N_48824,N_48836);
nand U49212 (N_49212,N_48962,N_48816);
or U49213 (N_49213,N_48913,N_48806);
nor U49214 (N_49214,N_48788,N_48902);
nor U49215 (N_49215,N_48848,N_48825);
and U49216 (N_49216,N_48924,N_48859);
nor U49217 (N_49217,N_48863,N_48835);
xor U49218 (N_49218,N_48859,N_48952);
nand U49219 (N_49219,N_48993,N_48761);
or U49220 (N_49220,N_48766,N_48763);
xnor U49221 (N_49221,N_48830,N_48950);
nand U49222 (N_49222,N_48965,N_48877);
xnor U49223 (N_49223,N_48958,N_48851);
or U49224 (N_49224,N_48792,N_48968);
or U49225 (N_49225,N_48843,N_48780);
xnor U49226 (N_49226,N_48890,N_48766);
nand U49227 (N_49227,N_48917,N_48953);
xor U49228 (N_49228,N_48900,N_48897);
xor U49229 (N_49229,N_48886,N_48920);
or U49230 (N_49230,N_48758,N_48862);
or U49231 (N_49231,N_48945,N_48784);
or U49232 (N_49232,N_48854,N_48876);
or U49233 (N_49233,N_48772,N_48953);
or U49234 (N_49234,N_48929,N_48815);
or U49235 (N_49235,N_48848,N_48856);
xor U49236 (N_49236,N_48800,N_48785);
xnor U49237 (N_49237,N_48857,N_48848);
nand U49238 (N_49238,N_48951,N_48938);
and U49239 (N_49239,N_48804,N_48783);
nand U49240 (N_49240,N_48875,N_48870);
nor U49241 (N_49241,N_48777,N_48826);
nor U49242 (N_49242,N_48972,N_48751);
nand U49243 (N_49243,N_48828,N_48878);
or U49244 (N_49244,N_48927,N_48859);
nand U49245 (N_49245,N_48797,N_48981);
xor U49246 (N_49246,N_48987,N_48940);
nand U49247 (N_49247,N_48757,N_48957);
nor U49248 (N_49248,N_48915,N_48836);
nor U49249 (N_49249,N_48924,N_48901);
and U49250 (N_49250,N_49068,N_49180);
nor U49251 (N_49251,N_49174,N_49207);
nor U49252 (N_49252,N_49248,N_49022);
and U49253 (N_49253,N_49192,N_49143);
nor U49254 (N_49254,N_49037,N_49050);
xor U49255 (N_49255,N_49246,N_49033);
and U49256 (N_49256,N_49157,N_49001);
nand U49257 (N_49257,N_49016,N_49231);
or U49258 (N_49258,N_49185,N_49079);
or U49259 (N_49259,N_49109,N_49166);
nor U49260 (N_49260,N_49142,N_49223);
and U49261 (N_49261,N_49034,N_49235);
or U49262 (N_49262,N_49072,N_49116);
xor U49263 (N_49263,N_49029,N_49010);
nand U49264 (N_49264,N_49169,N_49240);
or U49265 (N_49265,N_49154,N_49077);
nand U49266 (N_49266,N_49106,N_49130);
nor U49267 (N_49267,N_49242,N_49117);
xor U49268 (N_49268,N_49214,N_49136);
xor U49269 (N_49269,N_49119,N_49047);
and U49270 (N_49270,N_49186,N_49243);
xor U49271 (N_49271,N_49045,N_49151);
nand U49272 (N_49272,N_49206,N_49188);
xnor U49273 (N_49273,N_49177,N_49115);
nand U49274 (N_49274,N_49225,N_49201);
and U49275 (N_49275,N_49172,N_49126);
and U49276 (N_49276,N_49063,N_49167);
nor U49277 (N_49277,N_49113,N_49043);
or U49278 (N_49278,N_49114,N_49159);
nor U49279 (N_49279,N_49102,N_49165);
or U49280 (N_49280,N_49082,N_49057);
nor U49281 (N_49281,N_49039,N_49215);
or U49282 (N_49282,N_49135,N_49104);
xnor U49283 (N_49283,N_49048,N_49209);
and U49284 (N_49284,N_49232,N_49245);
nor U49285 (N_49285,N_49003,N_49128);
or U49286 (N_49286,N_49024,N_49226);
nor U49287 (N_49287,N_49171,N_49196);
xnor U49288 (N_49288,N_49153,N_49093);
nand U49289 (N_49289,N_49073,N_49121);
or U49290 (N_49290,N_49139,N_49069);
and U49291 (N_49291,N_49004,N_49228);
nor U49292 (N_49292,N_49056,N_49013);
xnor U49293 (N_49293,N_49198,N_49249);
or U49294 (N_49294,N_49229,N_49149);
nor U49295 (N_49295,N_49012,N_49061);
nor U49296 (N_49296,N_49161,N_49191);
or U49297 (N_49297,N_49091,N_49031);
nand U49298 (N_49298,N_49038,N_49125);
nor U49299 (N_49299,N_49233,N_49028);
or U49300 (N_49300,N_49118,N_49216);
nor U49301 (N_49301,N_49123,N_49182);
or U49302 (N_49302,N_49202,N_49213);
xnor U49303 (N_49303,N_49088,N_49076);
nand U49304 (N_49304,N_49129,N_49086);
and U49305 (N_49305,N_49236,N_49241);
xnor U49306 (N_49306,N_49194,N_49017);
xor U49307 (N_49307,N_49084,N_49224);
nor U49308 (N_49308,N_49127,N_49025);
or U49309 (N_49309,N_49140,N_49218);
nand U49310 (N_49310,N_49042,N_49211);
or U49311 (N_49311,N_49111,N_49176);
nand U49312 (N_49312,N_49200,N_49237);
nor U49313 (N_49313,N_49150,N_49217);
nor U49314 (N_49314,N_49005,N_49163);
nand U49315 (N_49315,N_49193,N_49011);
and U49316 (N_49316,N_49148,N_49099);
or U49317 (N_49317,N_49158,N_49179);
nand U49318 (N_49318,N_49002,N_49175);
nand U49319 (N_49319,N_49054,N_49009);
nand U49320 (N_49320,N_49044,N_49041);
or U49321 (N_49321,N_49210,N_49178);
nor U49322 (N_49322,N_49095,N_49107);
xor U49323 (N_49323,N_49134,N_49032);
xnor U49324 (N_49324,N_49103,N_49239);
or U49325 (N_49325,N_49083,N_49090);
xor U49326 (N_49326,N_49144,N_49085);
or U49327 (N_49327,N_49080,N_49051);
nor U49328 (N_49328,N_49059,N_49168);
or U49329 (N_49329,N_49014,N_49060);
nand U49330 (N_49330,N_49027,N_49105);
and U49331 (N_49331,N_49173,N_49058);
nor U49332 (N_49332,N_49049,N_49075);
nor U49333 (N_49333,N_49030,N_49074);
nand U49334 (N_49334,N_49081,N_49055);
or U49335 (N_49335,N_49067,N_49195);
xnor U49336 (N_49336,N_49170,N_49138);
and U49337 (N_49337,N_49124,N_49162);
nor U49338 (N_49338,N_49007,N_49197);
nor U49339 (N_49339,N_49087,N_49146);
or U49340 (N_49340,N_49208,N_49187);
xor U49341 (N_49341,N_49141,N_49244);
or U49342 (N_49342,N_49098,N_49108);
nand U49343 (N_49343,N_49203,N_49238);
or U49344 (N_49344,N_49147,N_49219);
and U49345 (N_49345,N_49184,N_49132);
nand U49346 (N_49346,N_49100,N_49052);
nor U49347 (N_49347,N_49092,N_49097);
or U49348 (N_49348,N_49040,N_49204);
or U49349 (N_49349,N_49078,N_49183);
or U49350 (N_49350,N_49120,N_49220);
or U49351 (N_49351,N_49131,N_49018);
xnor U49352 (N_49352,N_49221,N_49205);
nand U49353 (N_49353,N_49152,N_49015);
and U49354 (N_49354,N_49190,N_49019);
xor U49355 (N_49355,N_49234,N_49189);
nand U49356 (N_49356,N_49036,N_49156);
nor U49357 (N_49357,N_49008,N_49021);
and U49358 (N_49358,N_49006,N_49035);
nand U49359 (N_49359,N_49112,N_49096);
nor U49360 (N_49360,N_49094,N_49089);
nor U49361 (N_49361,N_49133,N_49023);
nor U49362 (N_49362,N_49145,N_49160);
xor U49363 (N_49363,N_49053,N_49046);
or U49364 (N_49364,N_49000,N_49181);
xor U49365 (N_49365,N_49064,N_49247);
nor U49366 (N_49366,N_49071,N_49020);
nor U49367 (N_49367,N_49066,N_49101);
and U49368 (N_49368,N_49227,N_49110);
or U49369 (N_49369,N_49222,N_49062);
xnor U49370 (N_49370,N_49137,N_49230);
nand U49371 (N_49371,N_49199,N_49155);
and U49372 (N_49372,N_49065,N_49026);
and U49373 (N_49373,N_49070,N_49122);
or U49374 (N_49374,N_49212,N_49164);
and U49375 (N_49375,N_49056,N_49188);
nor U49376 (N_49376,N_49132,N_49224);
nand U49377 (N_49377,N_49047,N_49176);
and U49378 (N_49378,N_49231,N_49116);
and U49379 (N_49379,N_49076,N_49072);
nand U49380 (N_49380,N_49097,N_49163);
nor U49381 (N_49381,N_49122,N_49084);
xnor U49382 (N_49382,N_49037,N_49153);
or U49383 (N_49383,N_49015,N_49112);
xnor U49384 (N_49384,N_49136,N_49028);
xnor U49385 (N_49385,N_49234,N_49155);
nor U49386 (N_49386,N_49136,N_49002);
nor U49387 (N_49387,N_49191,N_49215);
or U49388 (N_49388,N_49236,N_49024);
nor U49389 (N_49389,N_49060,N_49102);
or U49390 (N_49390,N_49059,N_49157);
and U49391 (N_49391,N_49167,N_49021);
or U49392 (N_49392,N_49186,N_49015);
and U49393 (N_49393,N_49217,N_49027);
and U49394 (N_49394,N_49226,N_49054);
nand U49395 (N_49395,N_49023,N_49164);
and U49396 (N_49396,N_49165,N_49204);
xnor U49397 (N_49397,N_49127,N_49136);
nor U49398 (N_49398,N_49246,N_49127);
nor U49399 (N_49399,N_49084,N_49062);
xnor U49400 (N_49400,N_49172,N_49009);
nor U49401 (N_49401,N_49158,N_49079);
and U49402 (N_49402,N_49134,N_49196);
xnor U49403 (N_49403,N_49154,N_49144);
xnor U49404 (N_49404,N_49142,N_49206);
nand U49405 (N_49405,N_49185,N_49094);
nor U49406 (N_49406,N_49024,N_49078);
or U49407 (N_49407,N_49132,N_49012);
xnor U49408 (N_49408,N_49004,N_49219);
nand U49409 (N_49409,N_49095,N_49149);
nand U49410 (N_49410,N_49020,N_49226);
nand U49411 (N_49411,N_49123,N_49149);
and U49412 (N_49412,N_49111,N_49032);
and U49413 (N_49413,N_49000,N_49077);
xor U49414 (N_49414,N_49073,N_49034);
xor U49415 (N_49415,N_49117,N_49012);
and U49416 (N_49416,N_49059,N_49011);
or U49417 (N_49417,N_49225,N_49085);
or U49418 (N_49418,N_49122,N_49033);
xor U49419 (N_49419,N_49160,N_49044);
nand U49420 (N_49420,N_49042,N_49191);
nor U49421 (N_49421,N_49000,N_49039);
nand U49422 (N_49422,N_49062,N_49177);
and U49423 (N_49423,N_49082,N_49166);
nor U49424 (N_49424,N_49116,N_49148);
xor U49425 (N_49425,N_49078,N_49055);
and U49426 (N_49426,N_49034,N_49169);
nand U49427 (N_49427,N_49214,N_49137);
and U49428 (N_49428,N_49190,N_49089);
xnor U49429 (N_49429,N_49212,N_49095);
and U49430 (N_49430,N_49065,N_49212);
xor U49431 (N_49431,N_49013,N_49038);
nor U49432 (N_49432,N_49123,N_49020);
nand U49433 (N_49433,N_49017,N_49163);
or U49434 (N_49434,N_49008,N_49116);
nor U49435 (N_49435,N_49091,N_49190);
nor U49436 (N_49436,N_49008,N_49214);
nand U49437 (N_49437,N_49032,N_49236);
xor U49438 (N_49438,N_49038,N_49184);
and U49439 (N_49439,N_49050,N_49064);
xnor U49440 (N_49440,N_49025,N_49029);
nor U49441 (N_49441,N_49065,N_49182);
nor U49442 (N_49442,N_49019,N_49171);
and U49443 (N_49443,N_49035,N_49172);
xor U49444 (N_49444,N_49203,N_49065);
nand U49445 (N_49445,N_49191,N_49130);
nand U49446 (N_49446,N_49177,N_49220);
xnor U49447 (N_49447,N_49195,N_49175);
nand U49448 (N_49448,N_49188,N_49111);
nor U49449 (N_49449,N_49053,N_49055);
nor U49450 (N_49450,N_49035,N_49193);
nor U49451 (N_49451,N_49139,N_49132);
nand U49452 (N_49452,N_49041,N_49169);
xor U49453 (N_49453,N_49024,N_49170);
xnor U49454 (N_49454,N_49037,N_49070);
or U49455 (N_49455,N_49173,N_49163);
nand U49456 (N_49456,N_49153,N_49064);
nand U49457 (N_49457,N_49159,N_49130);
and U49458 (N_49458,N_49060,N_49243);
nor U49459 (N_49459,N_49185,N_49089);
nor U49460 (N_49460,N_49060,N_49077);
nor U49461 (N_49461,N_49098,N_49247);
xnor U49462 (N_49462,N_49070,N_49170);
or U49463 (N_49463,N_49108,N_49134);
nand U49464 (N_49464,N_49067,N_49225);
xnor U49465 (N_49465,N_49247,N_49239);
nand U49466 (N_49466,N_49094,N_49067);
nor U49467 (N_49467,N_49024,N_49161);
xnor U49468 (N_49468,N_49067,N_49028);
nor U49469 (N_49469,N_49020,N_49238);
xnor U49470 (N_49470,N_49246,N_49151);
nand U49471 (N_49471,N_49021,N_49028);
nand U49472 (N_49472,N_49056,N_49201);
nand U49473 (N_49473,N_49181,N_49198);
nand U49474 (N_49474,N_49041,N_49115);
nor U49475 (N_49475,N_49085,N_49086);
xnor U49476 (N_49476,N_49233,N_49111);
nor U49477 (N_49477,N_49013,N_49168);
xor U49478 (N_49478,N_49158,N_49078);
and U49479 (N_49479,N_49102,N_49005);
and U49480 (N_49480,N_49089,N_49108);
and U49481 (N_49481,N_49146,N_49030);
and U49482 (N_49482,N_49185,N_49246);
nand U49483 (N_49483,N_49226,N_49233);
nand U49484 (N_49484,N_49225,N_49007);
xor U49485 (N_49485,N_49062,N_49226);
nor U49486 (N_49486,N_49160,N_49071);
nand U49487 (N_49487,N_49226,N_49075);
and U49488 (N_49488,N_49161,N_49230);
xnor U49489 (N_49489,N_49030,N_49153);
and U49490 (N_49490,N_49116,N_49218);
nand U49491 (N_49491,N_49105,N_49231);
or U49492 (N_49492,N_49084,N_49247);
xnor U49493 (N_49493,N_49173,N_49059);
xnor U49494 (N_49494,N_49060,N_49026);
and U49495 (N_49495,N_49104,N_49180);
nand U49496 (N_49496,N_49017,N_49054);
xnor U49497 (N_49497,N_49141,N_49229);
xnor U49498 (N_49498,N_49126,N_49133);
or U49499 (N_49499,N_49182,N_49169);
nor U49500 (N_49500,N_49329,N_49347);
and U49501 (N_49501,N_49322,N_49289);
xor U49502 (N_49502,N_49277,N_49465);
and U49503 (N_49503,N_49320,N_49354);
nand U49504 (N_49504,N_49263,N_49276);
and U49505 (N_49505,N_49379,N_49365);
and U49506 (N_49506,N_49472,N_49307);
or U49507 (N_49507,N_49324,N_49287);
xor U49508 (N_49508,N_49385,N_49291);
xor U49509 (N_49509,N_49351,N_49394);
or U49510 (N_49510,N_49398,N_49368);
xnor U49511 (N_49511,N_49313,N_49302);
or U49512 (N_49512,N_49382,N_49355);
xor U49513 (N_49513,N_49336,N_49334);
or U49514 (N_49514,N_49356,N_49498);
nor U49515 (N_49515,N_49434,N_49381);
nor U49516 (N_49516,N_49309,N_49428);
nand U49517 (N_49517,N_49339,N_49477);
or U49518 (N_49518,N_49429,N_49453);
nor U49519 (N_49519,N_49294,N_49257);
nor U49520 (N_49520,N_49449,N_49393);
nand U49521 (N_49521,N_49388,N_49284);
nor U49522 (N_49522,N_49425,N_49370);
or U49523 (N_49523,N_49481,N_49437);
or U49524 (N_49524,N_49312,N_49343);
and U49525 (N_49525,N_49488,N_49327);
or U49526 (N_49526,N_49269,N_49253);
xor U49527 (N_49527,N_49431,N_49358);
xnor U49528 (N_49528,N_49282,N_49461);
xor U49529 (N_49529,N_49409,N_49278);
or U49530 (N_49530,N_49340,N_49261);
nand U49531 (N_49531,N_49426,N_49457);
xor U49532 (N_49532,N_49468,N_49353);
nand U49533 (N_49533,N_49316,N_49366);
nand U49534 (N_49534,N_49485,N_49482);
xnor U49535 (N_49535,N_49396,N_49456);
nor U49536 (N_49536,N_49464,N_49346);
and U49537 (N_49537,N_49311,N_49293);
xor U49538 (N_49538,N_49386,N_49272);
xnor U49539 (N_49539,N_49273,N_49266);
and U49540 (N_49540,N_49331,N_49387);
xnor U49541 (N_49541,N_49421,N_49445);
nand U49542 (N_49542,N_49323,N_49254);
and U49543 (N_49543,N_49424,N_49330);
xor U49544 (N_49544,N_49443,N_49262);
or U49545 (N_49545,N_49268,N_49423);
and U49546 (N_49546,N_49321,N_49410);
and U49547 (N_49547,N_49275,N_49402);
and U49548 (N_49548,N_49484,N_49337);
and U49549 (N_49549,N_49487,N_49399);
nor U49550 (N_49550,N_49493,N_49486);
and U49551 (N_49551,N_49454,N_49474);
and U49552 (N_49552,N_49471,N_49460);
xnor U49553 (N_49553,N_49335,N_49427);
and U49554 (N_49554,N_49374,N_49391);
or U49555 (N_49555,N_49452,N_49436);
or U49556 (N_49556,N_49404,N_49397);
xor U49557 (N_49557,N_49299,N_49350);
nor U49558 (N_49558,N_49306,N_49314);
nor U49559 (N_49559,N_49480,N_49407);
xor U49560 (N_49560,N_49342,N_49304);
or U49561 (N_49561,N_49395,N_49414);
and U49562 (N_49562,N_49290,N_49280);
xnor U49563 (N_49563,N_49442,N_49352);
or U49564 (N_49564,N_49462,N_49440);
and U49565 (N_49565,N_49459,N_49470);
and U49566 (N_49566,N_49305,N_49378);
nand U49567 (N_49567,N_49258,N_49418);
or U49568 (N_49568,N_49412,N_49411);
nand U49569 (N_49569,N_49432,N_49372);
or U49570 (N_49570,N_49455,N_49435);
nor U49571 (N_49571,N_49271,N_49420);
xnor U49572 (N_49572,N_49341,N_49415);
and U49573 (N_49573,N_49458,N_49281);
and U49574 (N_49574,N_49315,N_49473);
nor U49575 (N_49575,N_49392,N_49450);
nor U49576 (N_49576,N_49466,N_49444);
and U49577 (N_49577,N_49446,N_49333);
or U49578 (N_49578,N_49403,N_49364);
xnor U49579 (N_49579,N_49361,N_49296);
nand U49580 (N_49580,N_49349,N_49298);
nand U49581 (N_49581,N_49300,N_49400);
and U49582 (N_49582,N_49463,N_49297);
nand U49583 (N_49583,N_49499,N_49325);
nand U49584 (N_49584,N_49492,N_49332);
or U49585 (N_49585,N_49360,N_49447);
and U49586 (N_49586,N_49359,N_49389);
nand U49587 (N_49587,N_49406,N_49338);
or U49588 (N_49588,N_49448,N_49274);
nor U49589 (N_49589,N_49256,N_49260);
nand U49590 (N_49590,N_49283,N_49483);
nor U49591 (N_49591,N_49362,N_49489);
and U49592 (N_49592,N_49496,N_49497);
nand U49593 (N_49593,N_49430,N_49417);
nand U49594 (N_49594,N_49250,N_49494);
xor U49595 (N_49595,N_49265,N_49288);
nor U49596 (N_49596,N_49326,N_49419);
nand U49597 (N_49597,N_49413,N_49408);
nor U49598 (N_49598,N_49390,N_49251);
nand U49599 (N_49599,N_49479,N_49467);
nor U49600 (N_49600,N_49348,N_49295);
nand U49601 (N_49601,N_49286,N_49317);
xnor U49602 (N_49602,N_49363,N_49375);
and U49603 (N_49603,N_49264,N_49345);
nand U49604 (N_49604,N_49369,N_49328);
nand U49605 (N_49605,N_49422,N_49367);
xnor U49606 (N_49606,N_49301,N_49469);
and U49607 (N_49607,N_49376,N_49371);
xor U49608 (N_49608,N_49308,N_49478);
nor U49609 (N_49609,N_49380,N_49270);
and U49610 (N_49610,N_49292,N_49303);
xnor U49611 (N_49611,N_49344,N_49475);
xor U49612 (N_49612,N_49319,N_49439);
nand U49613 (N_49613,N_49252,N_49255);
and U49614 (N_49614,N_49384,N_49310);
xor U49615 (N_49615,N_49401,N_49259);
or U49616 (N_49616,N_49405,N_49441);
xor U49617 (N_49617,N_49357,N_49495);
nor U49618 (N_49618,N_49491,N_49451);
or U49619 (N_49619,N_49279,N_49373);
xnor U49620 (N_49620,N_49416,N_49476);
xnor U49621 (N_49621,N_49490,N_49318);
xnor U49622 (N_49622,N_49267,N_49438);
xnor U49623 (N_49623,N_49377,N_49383);
and U49624 (N_49624,N_49433,N_49285);
or U49625 (N_49625,N_49476,N_49282);
xor U49626 (N_49626,N_49332,N_49416);
nand U49627 (N_49627,N_49298,N_49382);
xor U49628 (N_49628,N_49334,N_49446);
xnor U49629 (N_49629,N_49450,N_49416);
and U49630 (N_49630,N_49283,N_49467);
or U49631 (N_49631,N_49350,N_49437);
or U49632 (N_49632,N_49428,N_49383);
and U49633 (N_49633,N_49425,N_49399);
or U49634 (N_49634,N_49278,N_49410);
or U49635 (N_49635,N_49392,N_49333);
nand U49636 (N_49636,N_49460,N_49282);
and U49637 (N_49637,N_49467,N_49323);
and U49638 (N_49638,N_49470,N_49344);
nor U49639 (N_49639,N_49382,N_49499);
and U49640 (N_49640,N_49265,N_49449);
nand U49641 (N_49641,N_49277,N_49290);
nand U49642 (N_49642,N_49335,N_49385);
nand U49643 (N_49643,N_49342,N_49294);
nand U49644 (N_49644,N_49453,N_49418);
nor U49645 (N_49645,N_49373,N_49319);
nor U49646 (N_49646,N_49488,N_49262);
nor U49647 (N_49647,N_49380,N_49452);
xnor U49648 (N_49648,N_49369,N_49260);
nor U49649 (N_49649,N_49332,N_49338);
nor U49650 (N_49650,N_49387,N_49312);
nor U49651 (N_49651,N_49330,N_49454);
nor U49652 (N_49652,N_49393,N_49253);
and U49653 (N_49653,N_49398,N_49419);
nor U49654 (N_49654,N_49294,N_49498);
and U49655 (N_49655,N_49416,N_49438);
nor U49656 (N_49656,N_49363,N_49265);
nor U49657 (N_49657,N_49328,N_49429);
xor U49658 (N_49658,N_49387,N_49277);
xnor U49659 (N_49659,N_49380,N_49253);
or U49660 (N_49660,N_49367,N_49475);
or U49661 (N_49661,N_49329,N_49455);
nor U49662 (N_49662,N_49330,N_49285);
nor U49663 (N_49663,N_49292,N_49396);
or U49664 (N_49664,N_49291,N_49472);
nand U49665 (N_49665,N_49283,N_49471);
or U49666 (N_49666,N_49448,N_49376);
nand U49667 (N_49667,N_49365,N_49479);
and U49668 (N_49668,N_49400,N_49494);
and U49669 (N_49669,N_49328,N_49482);
and U49670 (N_49670,N_49389,N_49490);
and U49671 (N_49671,N_49429,N_49478);
nand U49672 (N_49672,N_49419,N_49261);
nand U49673 (N_49673,N_49388,N_49266);
nand U49674 (N_49674,N_49323,N_49496);
nor U49675 (N_49675,N_49497,N_49389);
xor U49676 (N_49676,N_49388,N_49374);
nor U49677 (N_49677,N_49478,N_49441);
xnor U49678 (N_49678,N_49281,N_49495);
xnor U49679 (N_49679,N_49268,N_49381);
xnor U49680 (N_49680,N_49310,N_49288);
nor U49681 (N_49681,N_49314,N_49301);
nand U49682 (N_49682,N_49357,N_49393);
and U49683 (N_49683,N_49300,N_49315);
or U49684 (N_49684,N_49447,N_49266);
and U49685 (N_49685,N_49481,N_49381);
and U49686 (N_49686,N_49387,N_49350);
and U49687 (N_49687,N_49428,N_49350);
xnor U49688 (N_49688,N_49381,N_49468);
nor U49689 (N_49689,N_49286,N_49410);
nor U49690 (N_49690,N_49356,N_49463);
and U49691 (N_49691,N_49398,N_49333);
nor U49692 (N_49692,N_49291,N_49303);
and U49693 (N_49693,N_49255,N_49417);
and U49694 (N_49694,N_49271,N_49424);
and U49695 (N_49695,N_49378,N_49467);
and U49696 (N_49696,N_49360,N_49427);
nand U49697 (N_49697,N_49491,N_49341);
or U49698 (N_49698,N_49253,N_49332);
nand U49699 (N_49699,N_49489,N_49306);
and U49700 (N_49700,N_49485,N_49442);
nor U49701 (N_49701,N_49327,N_49456);
xnor U49702 (N_49702,N_49448,N_49422);
nand U49703 (N_49703,N_49344,N_49375);
or U49704 (N_49704,N_49358,N_49329);
and U49705 (N_49705,N_49335,N_49428);
xnor U49706 (N_49706,N_49451,N_49380);
and U49707 (N_49707,N_49399,N_49344);
xor U49708 (N_49708,N_49440,N_49320);
nand U49709 (N_49709,N_49391,N_49282);
xor U49710 (N_49710,N_49449,N_49430);
and U49711 (N_49711,N_49260,N_49380);
and U49712 (N_49712,N_49353,N_49338);
xnor U49713 (N_49713,N_49377,N_49275);
nand U49714 (N_49714,N_49307,N_49331);
nand U49715 (N_49715,N_49330,N_49331);
nor U49716 (N_49716,N_49453,N_49416);
and U49717 (N_49717,N_49497,N_49449);
xnor U49718 (N_49718,N_49261,N_49287);
or U49719 (N_49719,N_49280,N_49346);
or U49720 (N_49720,N_49295,N_49310);
and U49721 (N_49721,N_49322,N_49317);
xor U49722 (N_49722,N_49466,N_49421);
nor U49723 (N_49723,N_49495,N_49450);
and U49724 (N_49724,N_49491,N_49494);
nand U49725 (N_49725,N_49320,N_49400);
or U49726 (N_49726,N_49405,N_49462);
or U49727 (N_49727,N_49434,N_49388);
or U49728 (N_49728,N_49417,N_49269);
nand U49729 (N_49729,N_49418,N_49491);
nand U49730 (N_49730,N_49366,N_49255);
nand U49731 (N_49731,N_49264,N_49250);
or U49732 (N_49732,N_49394,N_49303);
or U49733 (N_49733,N_49323,N_49424);
xnor U49734 (N_49734,N_49284,N_49435);
and U49735 (N_49735,N_49354,N_49393);
or U49736 (N_49736,N_49291,N_49466);
nor U49737 (N_49737,N_49358,N_49485);
and U49738 (N_49738,N_49347,N_49271);
or U49739 (N_49739,N_49314,N_49435);
nor U49740 (N_49740,N_49462,N_49491);
nand U49741 (N_49741,N_49411,N_49354);
and U49742 (N_49742,N_49456,N_49278);
or U49743 (N_49743,N_49295,N_49267);
xnor U49744 (N_49744,N_49464,N_49252);
xor U49745 (N_49745,N_49261,N_49368);
nor U49746 (N_49746,N_49324,N_49496);
nor U49747 (N_49747,N_49300,N_49254);
or U49748 (N_49748,N_49333,N_49481);
and U49749 (N_49749,N_49409,N_49463);
xnor U49750 (N_49750,N_49737,N_49676);
xnor U49751 (N_49751,N_49654,N_49646);
nand U49752 (N_49752,N_49740,N_49643);
and U49753 (N_49753,N_49633,N_49522);
and U49754 (N_49754,N_49559,N_49732);
or U49755 (N_49755,N_49506,N_49656);
nand U49756 (N_49756,N_49553,N_49583);
nand U49757 (N_49757,N_49550,N_49713);
xnor U49758 (N_49758,N_49743,N_49651);
nor U49759 (N_49759,N_49572,N_49710);
nor U49760 (N_49760,N_49671,N_49524);
nor U49761 (N_49761,N_49514,N_49597);
and U49762 (N_49762,N_49541,N_49575);
nand U49763 (N_49763,N_49700,N_49701);
or U49764 (N_49764,N_49703,N_49733);
nor U49765 (N_49765,N_49693,N_49558);
and U49766 (N_49766,N_49725,N_49730);
nand U49767 (N_49767,N_49606,N_49504);
or U49768 (N_49768,N_49557,N_49660);
or U49769 (N_49769,N_49711,N_49600);
or U49770 (N_49770,N_49515,N_49644);
xor U49771 (N_49771,N_49645,N_49578);
or U49772 (N_49772,N_49688,N_49636);
xnor U49773 (N_49773,N_49590,N_49562);
and U49774 (N_49774,N_49649,N_49702);
nor U49775 (N_49775,N_49637,N_49641);
xor U49776 (N_49776,N_49692,N_49610);
nand U49777 (N_49777,N_49502,N_49564);
xor U49778 (N_49778,N_49519,N_49736);
and U49779 (N_49779,N_49611,N_49563);
xnor U49780 (N_49780,N_49704,N_49567);
xor U49781 (N_49781,N_49532,N_49694);
and U49782 (N_49782,N_49531,N_49593);
nand U49783 (N_49783,N_49680,N_49708);
nand U49784 (N_49784,N_49674,N_49620);
xor U49785 (N_49785,N_49561,N_49690);
nor U49786 (N_49786,N_49626,N_49529);
xor U49787 (N_49787,N_49540,N_49536);
and U49788 (N_49788,N_49508,N_49679);
nor U49789 (N_49789,N_49566,N_49503);
nand U49790 (N_49790,N_49748,N_49568);
or U49791 (N_49791,N_49523,N_49603);
xor U49792 (N_49792,N_49683,N_49602);
xor U49793 (N_49793,N_49608,N_49618);
nor U49794 (N_49794,N_49580,N_49731);
nor U49795 (N_49795,N_49662,N_49554);
or U49796 (N_49796,N_49709,N_49509);
and U49797 (N_49797,N_49686,N_49664);
nand U49798 (N_49798,N_49623,N_49714);
and U49799 (N_49799,N_49621,N_49663);
nor U49800 (N_49800,N_49658,N_49587);
nor U49801 (N_49801,N_49517,N_49707);
nor U49802 (N_49802,N_49538,N_49742);
nand U49803 (N_49803,N_49601,N_49726);
and U49804 (N_49804,N_49581,N_49582);
and U49805 (N_49805,N_49729,N_49548);
and U49806 (N_49806,N_49652,N_49675);
and U49807 (N_49807,N_49560,N_49598);
xor U49808 (N_49808,N_49542,N_49642);
or U49809 (N_49809,N_49659,N_49571);
nand U49810 (N_49810,N_49589,N_49573);
xnor U49811 (N_49811,N_49706,N_49512);
nand U49812 (N_49812,N_49655,N_49591);
or U49813 (N_49813,N_49691,N_49661);
nand U49814 (N_49814,N_49697,N_49588);
xor U49815 (N_49815,N_49685,N_49635);
xor U49816 (N_49816,N_49716,N_49534);
xnor U49817 (N_49817,N_49634,N_49647);
xor U49818 (N_49818,N_49734,N_49715);
and U49819 (N_49819,N_49574,N_49594);
nand U49820 (N_49820,N_49695,N_49526);
nand U49821 (N_49821,N_49579,N_49551);
xnor U49822 (N_49822,N_49543,N_49595);
nor U49823 (N_49823,N_49552,N_49530);
or U49824 (N_49824,N_49576,N_49744);
xor U49825 (N_49825,N_49570,N_49681);
and U49826 (N_49826,N_49614,N_49630);
nand U49827 (N_49827,N_49741,N_49665);
nand U49828 (N_49828,N_49670,N_49705);
or U49829 (N_49829,N_49749,N_49516);
nand U49830 (N_49830,N_49500,N_49520);
or U49831 (N_49831,N_49527,N_49698);
xor U49832 (N_49832,N_49505,N_49632);
or U49833 (N_49833,N_49615,N_49546);
nand U49834 (N_49834,N_49604,N_49687);
xnor U49835 (N_49835,N_49616,N_49728);
nor U49836 (N_49836,N_49668,N_49617);
nor U49837 (N_49837,N_49510,N_49628);
or U49838 (N_49838,N_49682,N_49673);
nor U49839 (N_49839,N_49657,N_49556);
nand U49840 (N_49840,N_49545,N_49513);
xnor U49841 (N_49841,N_49719,N_49607);
nand U49842 (N_49842,N_49535,N_49577);
xnor U49843 (N_49843,N_49511,N_49605);
nand U49844 (N_49844,N_49738,N_49507);
nand U49845 (N_49845,N_49747,N_49565);
or U49846 (N_49846,N_49547,N_49625);
nor U49847 (N_49847,N_49569,N_49586);
xor U49848 (N_49848,N_49629,N_49599);
nor U49849 (N_49849,N_49739,N_49613);
or U49850 (N_49850,N_49684,N_49650);
nand U49851 (N_49851,N_49624,N_49735);
nor U49852 (N_49852,N_49678,N_49501);
and U49853 (N_49853,N_49727,N_49612);
and U49854 (N_49854,N_49622,N_49712);
or U49855 (N_49855,N_49746,N_49717);
or U49856 (N_49856,N_49585,N_49718);
nand U49857 (N_49857,N_49528,N_49592);
xnor U49858 (N_49858,N_49609,N_49584);
xnor U49859 (N_49859,N_49653,N_49539);
nor U49860 (N_49860,N_49537,N_49521);
and U49861 (N_49861,N_49555,N_49638);
and U49862 (N_49862,N_49720,N_49721);
nor U49863 (N_49863,N_49596,N_49631);
or U49864 (N_49864,N_49723,N_49648);
or U49865 (N_49865,N_49549,N_49666);
or U49866 (N_49866,N_49619,N_49639);
nor U49867 (N_49867,N_49669,N_49745);
or U49868 (N_49868,N_49667,N_49696);
or U49869 (N_49869,N_49722,N_49518);
xor U49870 (N_49870,N_49677,N_49724);
xnor U49871 (N_49871,N_49689,N_49525);
nand U49872 (N_49872,N_49544,N_49699);
or U49873 (N_49873,N_49672,N_49627);
nand U49874 (N_49874,N_49533,N_49640);
nor U49875 (N_49875,N_49602,N_49736);
xnor U49876 (N_49876,N_49515,N_49530);
nor U49877 (N_49877,N_49634,N_49655);
nor U49878 (N_49878,N_49591,N_49504);
nor U49879 (N_49879,N_49611,N_49666);
and U49880 (N_49880,N_49593,N_49731);
or U49881 (N_49881,N_49674,N_49740);
nor U49882 (N_49882,N_49596,N_49597);
or U49883 (N_49883,N_49718,N_49624);
or U49884 (N_49884,N_49533,N_49532);
and U49885 (N_49885,N_49628,N_49606);
xnor U49886 (N_49886,N_49633,N_49619);
nor U49887 (N_49887,N_49568,N_49671);
xor U49888 (N_49888,N_49676,N_49728);
or U49889 (N_49889,N_49505,N_49702);
or U49890 (N_49890,N_49508,N_49572);
nor U49891 (N_49891,N_49630,N_49731);
and U49892 (N_49892,N_49716,N_49656);
nor U49893 (N_49893,N_49662,N_49639);
nand U49894 (N_49894,N_49737,N_49522);
and U49895 (N_49895,N_49541,N_49504);
and U49896 (N_49896,N_49694,N_49673);
and U49897 (N_49897,N_49583,N_49721);
xor U49898 (N_49898,N_49534,N_49634);
nand U49899 (N_49899,N_49691,N_49517);
and U49900 (N_49900,N_49520,N_49521);
and U49901 (N_49901,N_49502,N_49727);
nand U49902 (N_49902,N_49508,N_49561);
or U49903 (N_49903,N_49612,N_49677);
xnor U49904 (N_49904,N_49608,N_49733);
and U49905 (N_49905,N_49571,N_49691);
nand U49906 (N_49906,N_49667,N_49523);
xnor U49907 (N_49907,N_49514,N_49522);
nand U49908 (N_49908,N_49519,N_49583);
or U49909 (N_49909,N_49532,N_49668);
nor U49910 (N_49910,N_49728,N_49583);
and U49911 (N_49911,N_49582,N_49602);
and U49912 (N_49912,N_49550,N_49556);
xor U49913 (N_49913,N_49509,N_49540);
nand U49914 (N_49914,N_49529,N_49570);
or U49915 (N_49915,N_49508,N_49741);
xnor U49916 (N_49916,N_49737,N_49715);
xnor U49917 (N_49917,N_49729,N_49542);
nor U49918 (N_49918,N_49608,N_49664);
or U49919 (N_49919,N_49590,N_49642);
or U49920 (N_49920,N_49653,N_49523);
xnor U49921 (N_49921,N_49672,N_49563);
and U49922 (N_49922,N_49662,N_49685);
xor U49923 (N_49923,N_49525,N_49730);
and U49924 (N_49924,N_49551,N_49643);
nand U49925 (N_49925,N_49660,N_49527);
nor U49926 (N_49926,N_49630,N_49682);
and U49927 (N_49927,N_49702,N_49566);
and U49928 (N_49928,N_49515,N_49665);
nor U49929 (N_49929,N_49701,N_49549);
nand U49930 (N_49930,N_49574,N_49716);
xor U49931 (N_49931,N_49726,N_49695);
xnor U49932 (N_49932,N_49679,N_49698);
nor U49933 (N_49933,N_49681,N_49540);
nor U49934 (N_49934,N_49680,N_49529);
or U49935 (N_49935,N_49631,N_49646);
xnor U49936 (N_49936,N_49692,N_49730);
or U49937 (N_49937,N_49615,N_49517);
and U49938 (N_49938,N_49688,N_49587);
and U49939 (N_49939,N_49552,N_49693);
nand U49940 (N_49940,N_49674,N_49501);
or U49941 (N_49941,N_49598,N_49747);
nand U49942 (N_49942,N_49729,N_49501);
or U49943 (N_49943,N_49546,N_49696);
and U49944 (N_49944,N_49614,N_49631);
nor U49945 (N_49945,N_49560,N_49701);
nand U49946 (N_49946,N_49553,N_49557);
nand U49947 (N_49947,N_49715,N_49606);
or U49948 (N_49948,N_49647,N_49617);
xor U49949 (N_49949,N_49702,N_49661);
nor U49950 (N_49950,N_49592,N_49744);
nor U49951 (N_49951,N_49737,N_49536);
nand U49952 (N_49952,N_49564,N_49571);
and U49953 (N_49953,N_49649,N_49743);
nor U49954 (N_49954,N_49556,N_49725);
and U49955 (N_49955,N_49605,N_49632);
nor U49956 (N_49956,N_49721,N_49614);
nor U49957 (N_49957,N_49703,N_49614);
nand U49958 (N_49958,N_49639,N_49527);
xor U49959 (N_49959,N_49701,N_49554);
or U49960 (N_49960,N_49512,N_49709);
and U49961 (N_49961,N_49539,N_49681);
nand U49962 (N_49962,N_49520,N_49643);
and U49963 (N_49963,N_49664,N_49641);
nand U49964 (N_49964,N_49642,N_49621);
nor U49965 (N_49965,N_49655,N_49738);
xnor U49966 (N_49966,N_49565,N_49745);
or U49967 (N_49967,N_49542,N_49597);
and U49968 (N_49968,N_49675,N_49678);
nand U49969 (N_49969,N_49612,N_49585);
nor U49970 (N_49970,N_49699,N_49670);
or U49971 (N_49971,N_49627,N_49650);
and U49972 (N_49972,N_49598,N_49739);
and U49973 (N_49973,N_49717,N_49544);
and U49974 (N_49974,N_49544,N_49504);
nor U49975 (N_49975,N_49696,N_49556);
and U49976 (N_49976,N_49740,N_49625);
or U49977 (N_49977,N_49646,N_49701);
xnor U49978 (N_49978,N_49629,N_49659);
and U49979 (N_49979,N_49632,N_49548);
and U49980 (N_49980,N_49640,N_49726);
and U49981 (N_49981,N_49725,N_49749);
or U49982 (N_49982,N_49502,N_49565);
or U49983 (N_49983,N_49718,N_49608);
and U49984 (N_49984,N_49730,N_49666);
and U49985 (N_49985,N_49643,N_49715);
xor U49986 (N_49986,N_49508,N_49646);
nand U49987 (N_49987,N_49651,N_49589);
nor U49988 (N_49988,N_49621,N_49631);
nand U49989 (N_49989,N_49626,N_49650);
xor U49990 (N_49990,N_49711,N_49725);
and U49991 (N_49991,N_49735,N_49507);
and U49992 (N_49992,N_49694,N_49668);
xor U49993 (N_49993,N_49568,N_49659);
nand U49994 (N_49994,N_49661,N_49606);
and U49995 (N_49995,N_49636,N_49631);
nor U49996 (N_49996,N_49588,N_49676);
xor U49997 (N_49997,N_49634,N_49739);
xnor U49998 (N_49998,N_49513,N_49692);
xnor U49999 (N_49999,N_49546,N_49617);
or UO_0 (O_0,N_49943,N_49805);
nor UO_1 (O_1,N_49879,N_49929);
nand UO_2 (O_2,N_49979,N_49931);
or UO_3 (O_3,N_49985,N_49843);
nand UO_4 (O_4,N_49803,N_49952);
nor UO_5 (O_5,N_49864,N_49983);
or UO_6 (O_6,N_49834,N_49961);
nand UO_7 (O_7,N_49772,N_49957);
nand UO_8 (O_8,N_49824,N_49756);
nand UO_9 (O_9,N_49764,N_49938);
nand UO_10 (O_10,N_49826,N_49838);
nor UO_11 (O_11,N_49862,N_49987);
nand UO_12 (O_12,N_49832,N_49883);
nand UO_13 (O_13,N_49982,N_49912);
nand UO_14 (O_14,N_49853,N_49860);
and UO_15 (O_15,N_49777,N_49954);
xor UO_16 (O_16,N_49973,N_49876);
or UO_17 (O_17,N_49924,N_49874);
or UO_18 (O_18,N_49820,N_49833);
or UO_19 (O_19,N_49950,N_49995);
nand UO_20 (O_20,N_49927,N_49873);
and UO_21 (O_21,N_49844,N_49845);
xor UO_22 (O_22,N_49786,N_49768);
xor UO_23 (O_23,N_49794,N_49932);
xnor UO_24 (O_24,N_49795,N_49866);
xnor UO_25 (O_25,N_49933,N_49976);
xor UO_26 (O_26,N_49969,N_49899);
and UO_27 (O_27,N_49752,N_49967);
nand UO_28 (O_28,N_49896,N_49882);
xnor UO_29 (O_29,N_49780,N_49953);
nand UO_30 (O_30,N_49827,N_49947);
nor UO_31 (O_31,N_49992,N_49926);
nand UO_32 (O_32,N_49903,N_49855);
nand UO_33 (O_33,N_49767,N_49887);
nor UO_34 (O_34,N_49817,N_49893);
nor UO_35 (O_35,N_49766,N_49911);
and UO_36 (O_36,N_49946,N_49812);
or UO_37 (O_37,N_49810,N_49831);
nand UO_38 (O_38,N_49828,N_49854);
and UO_39 (O_39,N_49814,N_49997);
xnor UO_40 (O_40,N_49936,N_49930);
nand UO_41 (O_41,N_49822,N_49870);
or UO_42 (O_42,N_49986,N_49783);
and UO_43 (O_43,N_49800,N_49863);
nand UO_44 (O_44,N_49994,N_49765);
or UO_45 (O_45,N_49784,N_49923);
nor UO_46 (O_46,N_49815,N_49821);
and UO_47 (O_47,N_49900,N_49981);
and UO_48 (O_48,N_49888,N_49908);
or UO_49 (O_49,N_49949,N_49850);
or UO_50 (O_50,N_49788,N_49771);
and UO_51 (O_51,N_49974,N_49818);
xnor UO_52 (O_52,N_49977,N_49836);
nor UO_53 (O_53,N_49790,N_49915);
nor UO_54 (O_54,N_49901,N_49928);
nor UO_55 (O_55,N_49914,N_49813);
and UO_56 (O_56,N_49996,N_49945);
or UO_57 (O_57,N_49823,N_49802);
or UO_58 (O_58,N_49940,N_49789);
nand UO_59 (O_59,N_49846,N_49751);
xor UO_60 (O_60,N_49868,N_49966);
nand UO_61 (O_61,N_49935,N_49889);
or UO_62 (O_62,N_49934,N_49830);
and UO_63 (O_63,N_49847,N_49978);
or UO_64 (O_64,N_49857,N_49761);
and UO_65 (O_65,N_49964,N_49991);
or UO_66 (O_66,N_49762,N_49941);
nor UO_67 (O_67,N_49797,N_49808);
xnor UO_68 (O_68,N_49839,N_49798);
and UO_69 (O_69,N_49902,N_49921);
or UO_70 (O_70,N_49999,N_49913);
or UO_71 (O_71,N_49984,N_49759);
nor UO_72 (O_72,N_49849,N_49998);
nor UO_73 (O_73,N_49993,N_49816);
and UO_74 (O_74,N_49905,N_49804);
and UO_75 (O_75,N_49881,N_49763);
xor UO_76 (O_76,N_49890,N_49809);
xor UO_77 (O_77,N_49811,N_49975);
nand UO_78 (O_78,N_49910,N_49968);
nor UO_79 (O_79,N_49867,N_49886);
or UO_80 (O_80,N_49922,N_49785);
nand UO_81 (O_81,N_49774,N_49972);
and UO_82 (O_82,N_49859,N_49956);
and UO_83 (O_83,N_49962,N_49760);
or UO_84 (O_84,N_49989,N_49856);
nor UO_85 (O_85,N_49965,N_49796);
and UO_86 (O_86,N_49758,N_49880);
or UO_87 (O_87,N_49885,N_49750);
nand UO_88 (O_88,N_49861,N_49753);
nand UO_89 (O_89,N_49779,N_49959);
or UO_90 (O_90,N_49958,N_49840);
nor UO_91 (O_91,N_49782,N_49837);
and UO_92 (O_92,N_49909,N_49919);
nand UO_93 (O_93,N_49793,N_49825);
or UO_94 (O_94,N_49851,N_49897);
xor UO_95 (O_95,N_49904,N_49980);
or UO_96 (O_96,N_49769,N_49898);
nand UO_97 (O_97,N_49925,N_49757);
nand UO_98 (O_98,N_49918,N_49787);
nor UO_99 (O_99,N_49990,N_49799);
nor UO_100 (O_100,N_49942,N_49848);
nand UO_101 (O_101,N_49944,N_49819);
xnor UO_102 (O_102,N_49920,N_49895);
nor UO_103 (O_103,N_49971,N_49775);
or UO_104 (O_104,N_49865,N_49872);
nand UO_105 (O_105,N_49792,N_49801);
or UO_106 (O_106,N_49891,N_49960);
and UO_107 (O_107,N_49892,N_49858);
and UO_108 (O_108,N_49807,N_49842);
and UO_109 (O_109,N_49754,N_49871);
or UO_110 (O_110,N_49970,N_49829);
xnor UO_111 (O_111,N_49937,N_49988);
and UO_112 (O_112,N_49894,N_49778);
xor UO_113 (O_113,N_49877,N_49907);
and UO_114 (O_114,N_49884,N_49841);
nand UO_115 (O_115,N_49875,N_49773);
or UO_116 (O_116,N_49806,N_49955);
nor UO_117 (O_117,N_49948,N_49770);
xor UO_118 (O_118,N_49776,N_49939);
nand UO_119 (O_119,N_49852,N_49963);
nand UO_120 (O_120,N_49781,N_49951);
or UO_121 (O_121,N_49791,N_49906);
nand UO_122 (O_122,N_49917,N_49916);
or UO_123 (O_123,N_49869,N_49835);
or UO_124 (O_124,N_49755,N_49878);
nor UO_125 (O_125,N_49966,N_49873);
and UO_126 (O_126,N_49782,N_49932);
or UO_127 (O_127,N_49966,N_49900);
or UO_128 (O_128,N_49892,N_49968);
nand UO_129 (O_129,N_49905,N_49812);
or UO_130 (O_130,N_49770,N_49791);
xor UO_131 (O_131,N_49771,N_49964);
xnor UO_132 (O_132,N_49782,N_49973);
and UO_133 (O_133,N_49981,N_49957);
nor UO_134 (O_134,N_49981,N_49842);
xnor UO_135 (O_135,N_49840,N_49997);
nand UO_136 (O_136,N_49793,N_49843);
or UO_137 (O_137,N_49884,N_49831);
or UO_138 (O_138,N_49759,N_49919);
xor UO_139 (O_139,N_49837,N_49902);
xor UO_140 (O_140,N_49843,N_49833);
or UO_141 (O_141,N_49916,N_49831);
and UO_142 (O_142,N_49828,N_49888);
xor UO_143 (O_143,N_49922,N_49940);
and UO_144 (O_144,N_49952,N_49863);
nand UO_145 (O_145,N_49958,N_49846);
or UO_146 (O_146,N_49903,N_49952);
xor UO_147 (O_147,N_49756,N_49951);
or UO_148 (O_148,N_49979,N_49933);
and UO_149 (O_149,N_49865,N_49916);
nor UO_150 (O_150,N_49891,N_49836);
nand UO_151 (O_151,N_49923,N_49981);
or UO_152 (O_152,N_49804,N_49836);
nand UO_153 (O_153,N_49800,N_49973);
and UO_154 (O_154,N_49893,N_49940);
nand UO_155 (O_155,N_49830,N_49845);
xor UO_156 (O_156,N_49845,N_49812);
and UO_157 (O_157,N_49780,N_49852);
and UO_158 (O_158,N_49868,N_49848);
or UO_159 (O_159,N_49798,N_49940);
or UO_160 (O_160,N_49886,N_49854);
xnor UO_161 (O_161,N_49935,N_49900);
or UO_162 (O_162,N_49845,N_49999);
nand UO_163 (O_163,N_49987,N_49991);
nand UO_164 (O_164,N_49830,N_49980);
nor UO_165 (O_165,N_49794,N_49776);
or UO_166 (O_166,N_49824,N_49821);
nor UO_167 (O_167,N_49946,N_49874);
xnor UO_168 (O_168,N_49960,N_49931);
or UO_169 (O_169,N_49998,N_49839);
nand UO_170 (O_170,N_49882,N_49755);
xor UO_171 (O_171,N_49943,N_49882);
xor UO_172 (O_172,N_49834,N_49822);
and UO_173 (O_173,N_49974,N_49856);
and UO_174 (O_174,N_49772,N_49986);
or UO_175 (O_175,N_49810,N_49833);
nor UO_176 (O_176,N_49957,N_49915);
nand UO_177 (O_177,N_49786,N_49876);
xor UO_178 (O_178,N_49826,N_49885);
xor UO_179 (O_179,N_49867,N_49901);
nand UO_180 (O_180,N_49964,N_49758);
xnor UO_181 (O_181,N_49841,N_49828);
and UO_182 (O_182,N_49889,N_49820);
nor UO_183 (O_183,N_49937,N_49757);
nand UO_184 (O_184,N_49802,N_49989);
and UO_185 (O_185,N_49985,N_49965);
xor UO_186 (O_186,N_49771,N_49847);
and UO_187 (O_187,N_49910,N_49866);
or UO_188 (O_188,N_49811,N_49964);
xor UO_189 (O_189,N_49754,N_49792);
nand UO_190 (O_190,N_49993,N_49916);
nand UO_191 (O_191,N_49780,N_49806);
nor UO_192 (O_192,N_49845,N_49908);
nand UO_193 (O_193,N_49924,N_49866);
nand UO_194 (O_194,N_49833,N_49760);
xor UO_195 (O_195,N_49795,N_49947);
xor UO_196 (O_196,N_49946,N_49872);
nand UO_197 (O_197,N_49894,N_49985);
or UO_198 (O_198,N_49928,N_49809);
or UO_199 (O_199,N_49948,N_49871);
or UO_200 (O_200,N_49933,N_49940);
nor UO_201 (O_201,N_49967,N_49814);
xor UO_202 (O_202,N_49770,N_49928);
and UO_203 (O_203,N_49779,N_49826);
and UO_204 (O_204,N_49962,N_49791);
and UO_205 (O_205,N_49991,N_49801);
nor UO_206 (O_206,N_49770,N_49924);
nand UO_207 (O_207,N_49977,N_49965);
and UO_208 (O_208,N_49753,N_49982);
and UO_209 (O_209,N_49851,N_49861);
xnor UO_210 (O_210,N_49935,N_49866);
xor UO_211 (O_211,N_49900,N_49891);
or UO_212 (O_212,N_49995,N_49932);
nor UO_213 (O_213,N_49850,N_49830);
nor UO_214 (O_214,N_49938,N_49943);
xnor UO_215 (O_215,N_49875,N_49981);
and UO_216 (O_216,N_49859,N_49795);
or UO_217 (O_217,N_49925,N_49861);
xnor UO_218 (O_218,N_49945,N_49836);
or UO_219 (O_219,N_49810,N_49794);
nand UO_220 (O_220,N_49845,N_49776);
and UO_221 (O_221,N_49872,N_49858);
xor UO_222 (O_222,N_49845,N_49753);
nor UO_223 (O_223,N_49921,N_49849);
nor UO_224 (O_224,N_49925,N_49956);
nand UO_225 (O_225,N_49860,N_49963);
nor UO_226 (O_226,N_49815,N_49854);
xor UO_227 (O_227,N_49786,N_49873);
nor UO_228 (O_228,N_49916,N_49947);
xnor UO_229 (O_229,N_49910,N_49750);
nand UO_230 (O_230,N_49842,N_49866);
xor UO_231 (O_231,N_49878,N_49775);
and UO_232 (O_232,N_49909,N_49878);
or UO_233 (O_233,N_49896,N_49849);
nand UO_234 (O_234,N_49910,N_49964);
and UO_235 (O_235,N_49943,N_49759);
nand UO_236 (O_236,N_49750,N_49894);
or UO_237 (O_237,N_49812,N_49997);
nor UO_238 (O_238,N_49831,N_49976);
or UO_239 (O_239,N_49899,N_49788);
nand UO_240 (O_240,N_49776,N_49754);
and UO_241 (O_241,N_49860,N_49901);
xor UO_242 (O_242,N_49938,N_49883);
and UO_243 (O_243,N_49810,N_49963);
and UO_244 (O_244,N_49773,N_49863);
nor UO_245 (O_245,N_49793,N_49924);
nor UO_246 (O_246,N_49869,N_49788);
nor UO_247 (O_247,N_49967,N_49872);
and UO_248 (O_248,N_49928,N_49957);
nand UO_249 (O_249,N_49818,N_49936);
or UO_250 (O_250,N_49929,N_49774);
or UO_251 (O_251,N_49779,N_49979);
nor UO_252 (O_252,N_49901,N_49777);
and UO_253 (O_253,N_49940,N_49811);
and UO_254 (O_254,N_49782,N_49917);
and UO_255 (O_255,N_49882,N_49875);
nand UO_256 (O_256,N_49807,N_49915);
nor UO_257 (O_257,N_49925,N_49881);
nand UO_258 (O_258,N_49928,N_49979);
or UO_259 (O_259,N_49765,N_49962);
nor UO_260 (O_260,N_49864,N_49990);
xnor UO_261 (O_261,N_49931,N_49911);
nand UO_262 (O_262,N_49954,N_49844);
and UO_263 (O_263,N_49868,N_49962);
or UO_264 (O_264,N_49958,N_49897);
or UO_265 (O_265,N_49784,N_49974);
nor UO_266 (O_266,N_49787,N_49887);
nand UO_267 (O_267,N_49970,N_49973);
nor UO_268 (O_268,N_49778,N_49756);
nor UO_269 (O_269,N_49911,N_49923);
and UO_270 (O_270,N_49889,N_49825);
or UO_271 (O_271,N_49889,N_49852);
nor UO_272 (O_272,N_49892,N_49761);
or UO_273 (O_273,N_49942,N_49886);
nand UO_274 (O_274,N_49940,N_49979);
or UO_275 (O_275,N_49872,N_49961);
xor UO_276 (O_276,N_49880,N_49784);
xor UO_277 (O_277,N_49890,N_49922);
nor UO_278 (O_278,N_49915,N_49921);
and UO_279 (O_279,N_49967,N_49899);
or UO_280 (O_280,N_49872,N_49857);
nor UO_281 (O_281,N_49891,N_49945);
and UO_282 (O_282,N_49987,N_49996);
and UO_283 (O_283,N_49873,N_49761);
nand UO_284 (O_284,N_49841,N_49932);
and UO_285 (O_285,N_49918,N_49779);
nand UO_286 (O_286,N_49798,N_49915);
nor UO_287 (O_287,N_49985,N_49932);
and UO_288 (O_288,N_49887,N_49774);
xnor UO_289 (O_289,N_49838,N_49957);
xnor UO_290 (O_290,N_49835,N_49970);
or UO_291 (O_291,N_49844,N_49923);
nand UO_292 (O_292,N_49821,N_49843);
and UO_293 (O_293,N_49769,N_49781);
xor UO_294 (O_294,N_49936,N_49793);
or UO_295 (O_295,N_49770,N_49885);
xor UO_296 (O_296,N_49966,N_49904);
nor UO_297 (O_297,N_49956,N_49890);
nor UO_298 (O_298,N_49811,N_49831);
or UO_299 (O_299,N_49872,N_49817);
or UO_300 (O_300,N_49953,N_49982);
and UO_301 (O_301,N_49885,N_49850);
or UO_302 (O_302,N_49831,N_49812);
or UO_303 (O_303,N_49793,N_49833);
and UO_304 (O_304,N_49948,N_49805);
xor UO_305 (O_305,N_49815,N_49751);
nor UO_306 (O_306,N_49765,N_49998);
nand UO_307 (O_307,N_49792,N_49771);
and UO_308 (O_308,N_49903,N_49986);
or UO_309 (O_309,N_49816,N_49805);
xor UO_310 (O_310,N_49974,N_49925);
and UO_311 (O_311,N_49882,N_49988);
nor UO_312 (O_312,N_49962,N_49853);
and UO_313 (O_313,N_49783,N_49892);
and UO_314 (O_314,N_49880,N_49999);
nand UO_315 (O_315,N_49946,N_49800);
nor UO_316 (O_316,N_49891,N_49877);
nor UO_317 (O_317,N_49841,N_49916);
or UO_318 (O_318,N_49909,N_49892);
nor UO_319 (O_319,N_49823,N_49861);
nand UO_320 (O_320,N_49765,N_49946);
nor UO_321 (O_321,N_49796,N_49975);
nand UO_322 (O_322,N_49993,N_49865);
xnor UO_323 (O_323,N_49844,N_49806);
or UO_324 (O_324,N_49859,N_49825);
or UO_325 (O_325,N_49813,N_49910);
and UO_326 (O_326,N_49878,N_49786);
nor UO_327 (O_327,N_49786,N_49991);
xor UO_328 (O_328,N_49984,N_49997);
nor UO_329 (O_329,N_49804,N_49946);
or UO_330 (O_330,N_49844,N_49760);
and UO_331 (O_331,N_49753,N_49785);
xnor UO_332 (O_332,N_49772,N_49999);
nand UO_333 (O_333,N_49976,N_49918);
xor UO_334 (O_334,N_49939,N_49927);
xnor UO_335 (O_335,N_49813,N_49856);
and UO_336 (O_336,N_49866,N_49890);
xnor UO_337 (O_337,N_49836,N_49801);
or UO_338 (O_338,N_49807,N_49852);
xnor UO_339 (O_339,N_49931,N_49863);
nor UO_340 (O_340,N_49769,N_49884);
or UO_341 (O_341,N_49763,N_49858);
nand UO_342 (O_342,N_49995,N_49934);
and UO_343 (O_343,N_49793,N_49998);
nand UO_344 (O_344,N_49998,N_49870);
nand UO_345 (O_345,N_49917,N_49826);
xnor UO_346 (O_346,N_49824,N_49978);
nand UO_347 (O_347,N_49881,N_49764);
and UO_348 (O_348,N_49883,N_49880);
xor UO_349 (O_349,N_49911,N_49771);
and UO_350 (O_350,N_49857,N_49816);
and UO_351 (O_351,N_49888,N_49844);
nor UO_352 (O_352,N_49899,N_49906);
or UO_353 (O_353,N_49797,N_49867);
or UO_354 (O_354,N_49841,N_49820);
and UO_355 (O_355,N_49778,N_49855);
xor UO_356 (O_356,N_49852,N_49916);
or UO_357 (O_357,N_49832,N_49884);
and UO_358 (O_358,N_49782,N_49957);
nor UO_359 (O_359,N_49975,N_49895);
or UO_360 (O_360,N_49819,N_49942);
or UO_361 (O_361,N_49950,N_49804);
xnor UO_362 (O_362,N_49915,N_49975);
and UO_363 (O_363,N_49964,N_49887);
xor UO_364 (O_364,N_49891,N_49778);
and UO_365 (O_365,N_49937,N_49786);
xnor UO_366 (O_366,N_49920,N_49880);
or UO_367 (O_367,N_49763,N_49924);
xnor UO_368 (O_368,N_49821,N_49999);
xnor UO_369 (O_369,N_49765,N_49857);
nor UO_370 (O_370,N_49800,N_49960);
nor UO_371 (O_371,N_49764,N_49805);
nand UO_372 (O_372,N_49872,N_49804);
xnor UO_373 (O_373,N_49996,N_49761);
and UO_374 (O_374,N_49968,N_49832);
nand UO_375 (O_375,N_49773,N_49860);
or UO_376 (O_376,N_49897,N_49954);
and UO_377 (O_377,N_49798,N_49832);
or UO_378 (O_378,N_49832,N_49929);
xor UO_379 (O_379,N_49966,N_49880);
and UO_380 (O_380,N_49840,N_49993);
nand UO_381 (O_381,N_49839,N_49804);
and UO_382 (O_382,N_49968,N_49988);
or UO_383 (O_383,N_49959,N_49785);
or UO_384 (O_384,N_49988,N_49944);
xnor UO_385 (O_385,N_49888,N_49981);
xor UO_386 (O_386,N_49839,N_49891);
xnor UO_387 (O_387,N_49884,N_49941);
nand UO_388 (O_388,N_49943,N_49884);
or UO_389 (O_389,N_49866,N_49959);
nor UO_390 (O_390,N_49818,N_49903);
nor UO_391 (O_391,N_49768,N_49940);
and UO_392 (O_392,N_49796,N_49979);
xor UO_393 (O_393,N_49829,N_49861);
nand UO_394 (O_394,N_49862,N_49995);
nor UO_395 (O_395,N_49888,N_49800);
or UO_396 (O_396,N_49981,N_49935);
nand UO_397 (O_397,N_49969,N_49974);
and UO_398 (O_398,N_49911,N_49980);
xnor UO_399 (O_399,N_49890,N_49767);
and UO_400 (O_400,N_49797,N_49776);
nor UO_401 (O_401,N_49852,N_49837);
xor UO_402 (O_402,N_49927,N_49942);
xor UO_403 (O_403,N_49963,N_49851);
xor UO_404 (O_404,N_49972,N_49959);
nand UO_405 (O_405,N_49950,N_49772);
nor UO_406 (O_406,N_49974,N_49789);
nor UO_407 (O_407,N_49918,N_49932);
nor UO_408 (O_408,N_49968,N_49955);
xor UO_409 (O_409,N_49764,N_49844);
and UO_410 (O_410,N_49873,N_49911);
nor UO_411 (O_411,N_49840,N_49861);
or UO_412 (O_412,N_49884,N_49838);
xnor UO_413 (O_413,N_49955,N_49946);
nand UO_414 (O_414,N_49883,N_49992);
and UO_415 (O_415,N_49871,N_49771);
or UO_416 (O_416,N_49951,N_49875);
and UO_417 (O_417,N_49761,N_49768);
or UO_418 (O_418,N_49922,N_49891);
xnor UO_419 (O_419,N_49853,N_49773);
or UO_420 (O_420,N_49815,N_49993);
xor UO_421 (O_421,N_49864,N_49775);
and UO_422 (O_422,N_49928,N_49985);
and UO_423 (O_423,N_49980,N_49861);
and UO_424 (O_424,N_49957,N_49998);
or UO_425 (O_425,N_49964,N_49953);
xor UO_426 (O_426,N_49757,N_49865);
nand UO_427 (O_427,N_49958,N_49797);
and UO_428 (O_428,N_49829,N_49852);
and UO_429 (O_429,N_49820,N_49842);
and UO_430 (O_430,N_49760,N_49803);
nor UO_431 (O_431,N_49940,N_49876);
xor UO_432 (O_432,N_49773,N_49777);
nand UO_433 (O_433,N_49978,N_49821);
nand UO_434 (O_434,N_49856,N_49903);
xnor UO_435 (O_435,N_49824,N_49896);
nand UO_436 (O_436,N_49987,N_49895);
nand UO_437 (O_437,N_49882,N_49888);
xor UO_438 (O_438,N_49859,N_49896);
or UO_439 (O_439,N_49945,N_49942);
and UO_440 (O_440,N_49997,N_49860);
and UO_441 (O_441,N_49941,N_49863);
nor UO_442 (O_442,N_49788,N_49850);
nor UO_443 (O_443,N_49895,N_49943);
xor UO_444 (O_444,N_49901,N_49765);
or UO_445 (O_445,N_49897,N_49756);
nand UO_446 (O_446,N_49790,N_49804);
nor UO_447 (O_447,N_49868,N_49886);
xnor UO_448 (O_448,N_49882,N_49751);
nor UO_449 (O_449,N_49989,N_49756);
xnor UO_450 (O_450,N_49867,N_49784);
xnor UO_451 (O_451,N_49869,N_49755);
xnor UO_452 (O_452,N_49945,N_49854);
nor UO_453 (O_453,N_49943,N_49822);
xor UO_454 (O_454,N_49915,N_49967);
nand UO_455 (O_455,N_49829,N_49803);
nor UO_456 (O_456,N_49779,N_49816);
and UO_457 (O_457,N_49883,N_49907);
xnor UO_458 (O_458,N_49901,N_49863);
nand UO_459 (O_459,N_49823,N_49785);
nand UO_460 (O_460,N_49893,N_49939);
and UO_461 (O_461,N_49784,N_49833);
xnor UO_462 (O_462,N_49822,N_49775);
nand UO_463 (O_463,N_49992,N_49805);
or UO_464 (O_464,N_49913,N_49909);
xor UO_465 (O_465,N_49864,N_49875);
xor UO_466 (O_466,N_49895,N_49988);
xnor UO_467 (O_467,N_49755,N_49773);
and UO_468 (O_468,N_49861,N_49872);
nor UO_469 (O_469,N_49824,N_49900);
nand UO_470 (O_470,N_49998,N_49995);
nor UO_471 (O_471,N_49831,N_49996);
nand UO_472 (O_472,N_49756,N_49767);
nor UO_473 (O_473,N_49817,N_49943);
xor UO_474 (O_474,N_49863,N_49987);
nor UO_475 (O_475,N_49988,N_49775);
nor UO_476 (O_476,N_49978,N_49937);
or UO_477 (O_477,N_49888,N_49924);
and UO_478 (O_478,N_49854,N_49833);
nand UO_479 (O_479,N_49876,N_49753);
or UO_480 (O_480,N_49929,N_49962);
xnor UO_481 (O_481,N_49898,N_49930);
nor UO_482 (O_482,N_49775,N_49916);
and UO_483 (O_483,N_49911,N_49851);
nand UO_484 (O_484,N_49935,N_49902);
nor UO_485 (O_485,N_49864,N_49886);
nand UO_486 (O_486,N_49935,N_49808);
xnor UO_487 (O_487,N_49872,N_49853);
xor UO_488 (O_488,N_49965,N_49874);
nor UO_489 (O_489,N_49977,N_49983);
nand UO_490 (O_490,N_49954,N_49884);
and UO_491 (O_491,N_49912,N_49974);
nand UO_492 (O_492,N_49808,N_49893);
xnor UO_493 (O_493,N_49856,N_49956);
nand UO_494 (O_494,N_49764,N_49787);
or UO_495 (O_495,N_49773,N_49936);
nor UO_496 (O_496,N_49937,N_49830);
nand UO_497 (O_497,N_49983,N_49860);
xor UO_498 (O_498,N_49790,N_49818);
nand UO_499 (O_499,N_49878,N_49923);
or UO_500 (O_500,N_49868,N_49927);
xnor UO_501 (O_501,N_49790,N_49874);
and UO_502 (O_502,N_49917,N_49829);
nor UO_503 (O_503,N_49875,N_49778);
nand UO_504 (O_504,N_49765,N_49799);
nand UO_505 (O_505,N_49774,N_49838);
nor UO_506 (O_506,N_49907,N_49765);
or UO_507 (O_507,N_49982,N_49865);
nor UO_508 (O_508,N_49774,N_49788);
nand UO_509 (O_509,N_49835,N_49920);
nor UO_510 (O_510,N_49786,N_49821);
nor UO_511 (O_511,N_49812,N_49853);
nand UO_512 (O_512,N_49924,N_49752);
or UO_513 (O_513,N_49772,N_49798);
or UO_514 (O_514,N_49825,N_49808);
or UO_515 (O_515,N_49896,N_49856);
nor UO_516 (O_516,N_49758,N_49764);
nor UO_517 (O_517,N_49886,N_49953);
nor UO_518 (O_518,N_49849,N_49868);
and UO_519 (O_519,N_49893,N_49904);
nor UO_520 (O_520,N_49892,N_49914);
nor UO_521 (O_521,N_49881,N_49863);
nor UO_522 (O_522,N_49812,N_49773);
and UO_523 (O_523,N_49859,N_49811);
and UO_524 (O_524,N_49888,N_49933);
xor UO_525 (O_525,N_49999,N_49939);
nor UO_526 (O_526,N_49854,N_49770);
or UO_527 (O_527,N_49969,N_49901);
nand UO_528 (O_528,N_49925,N_49872);
or UO_529 (O_529,N_49782,N_49888);
or UO_530 (O_530,N_49940,N_49914);
nand UO_531 (O_531,N_49767,N_49938);
or UO_532 (O_532,N_49786,N_49973);
nand UO_533 (O_533,N_49908,N_49918);
xnor UO_534 (O_534,N_49855,N_49876);
nand UO_535 (O_535,N_49976,N_49884);
and UO_536 (O_536,N_49880,N_49817);
xnor UO_537 (O_537,N_49885,N_49872);
or UO_538 (O_538,N_49928,N_49755);
nand UO_539 (O_539,N_49776,N_49854);
nor UO_540 (O_540,N_49761,N_49850);
or UO_541 (O_541,N_49758,N_49984);
nand UO_542 (O_542,N_49779,N_49961);
and UO_543 (O_543,N_49852,N_49982);
and UO_544 (O_544,N_49814,N_49939);
xnor UO_545 (O_545,N_49905,N_49777);
and UO_546 (O_546,N_49987,N_49876);
nand UO_547 (O_547,N_49970,N_49960);
and UO_548 (O_548,N_49969,N_49845);
and UO_549 (O_549,N_49965,N_49929);
and UO_550 (O_550,N_49764,N_49937);
and UO_551 (O_551,N_49951,N_49877);
or UO_552 (O_552,N_49786,N_49918);
or UO_553 (O_553,N_49845,N_49921);
nor UO_554 (O_554,N_49769,N_49902);
and UO_555 (O_555,N_49864,N_49757);
xor UO_556 (O_556,N_49873,N_49796);
and UO_557 (O_557,N_49867,N_49939);
or UO_558 (O_558,N_49945,N_49785);
xor UO_559 (O_559,N_49835,N_49888);
nor UO_560 (O_560,N_49940,N_49853);
nand UO_561 (O_561,N_49793,N_49983);
nand UO_562 (O_562,N_49885,N_49793);
or UO_563 (O_563,N_49961,N_49934);
or UO_564 (O_564,N_49775,N_49979);
xor UO_565 (O_565,N_49954,N_49860);
xnor UO_566 (O_566,N_49992,N_49868);
xnor UO_567 (O_567,N_49992,N_49963);
xnor UO_568 (O_568,N_49871,N_49770);
nand UO_569 (O_569,N_49912,N_49910);
and UO_570 (O_570,N_49766,N_49885);
xnor UO_571 (O_571,N_49924,N_49881);
and UO_572 (O_572,N_49977,N_49963);
nor UO_573 (O_573,N_49847,N_49881);
xor UO_574 (O_574,N_49957,N_49798);
or UO_575 (O_575,N_49791,N_49976);
nor UO_576 (O_576,N_49782,N_49874);
nor UO_577 (O_577,N_49783,N_49944);
and UO_578 (O_578,N_49850,N_49781);
or UO_579 (O_579,N_49844,N_49797);
and UO_580 (O_580,N_49999,N_49969);
and UO_581 (O_581,N_49821,N_49875);
and UO_582 (O_582,N_49935,N_49825);
nand UO_583 (O_583,N_49899,N_49859);
or UO_584 (O_584,N_49788,N_49805);
or UO_585 (O_585,N_49801,N_49876);
and UO_586 (O_586,N_49796,N_49821);
nor UO_587 (O_587,N_49869,N_49860);
nand UO_588 (O_588,N_49916,N_49951);
nor UO_589 (O_589,N_49758,N_49974);
nor UO_590 (O_590,N_49877,N_49760);
or UO_591 (O_591,N_49991,N_49944);
and UO_592 (O_592,N_49763,N_49823);
and UO_593 (O_593,N_49939,N_49933);
and UO_594 (O_594,N_49761,N_49781);
and UO_595 (O_595,N_49816,N_49945);
and UO_596 (O_596,N_49836,N_49852);
and UO_597 (O_597,N_49882,N_49949);
nand UO_598 (O_598,N_49912,N_49965);
nor UO_599 (O_599,N_49916,N_49776);
or UO_600 (O_600,N_49969,N_49822);
or UO_601 (O_601,N_49895,N_49867);
nor UO_602 (O_602,N_49922,N_49765);
nor UO_603 (O_603,N_49825,N_49924);
xnor UO_604 (O_604,N_49754,N_49997);
or UO_605 (O_605,N_49995,N_49793);
xor UO_606 (O_606,N_49758,N_49934);
nand UO_607 (O_607,N_49894,N_49920);
or UO_608 (O_608,N_49783,N_49925);
xnor UO_609 (O_609,N_49911,N_49945);
nor UO_610 (O_610,N_49773,N_49790);
and UO_611 (O_611,N_49957,N_49871);
nand UO_612 (O_612,N_49751,N_49992);
nand UO_613 (O_613,N_49848,N_49941);
or UO_614 (O_614,N_49950,N_49917);
or UO_615 (O_615,N_49939,N_49891);
nand UO_616 (O_616,N_49962,N_49935);
xnor UO_617 (O_617,N_49916,N_49949);
nand UO_618 (O_618,N_49887,N_49818);
nand UO_619 (O_619,N_49908,N_49941);
and UO_620 (O_620,N_49971,N_49770);
nand UO_621 (O_621,N_49775,N_49932);
nor UO_622 (O_622,N_49881,N_49920);
xnor UO_623 (O_623,N_49808,N_49930);
or UO_624 (O_624,N_49979,N_49830);
xor UO_625 (O_625,N_49821,N_49884);
or UO_626 (O_626,N_49981,N_49789);
xnor UO_627 (O_627,N_49912,N_49848);
or UO_628 (O_628,N_49985,N_49863);
nor UO_629 (O_629,N_49883,N_49890);
nor UO_630 (O_630,N_49811,N_49789);
and UO_631 (O_631,N_49954,N_49776);
nand UO_632 (O_632,N_49901,N_49835);
nand UO_633 (O_633,N_49994,N_49792);
and UO_634 (O_634,N_49889,N_49903);
nand UO_635 (O_635,N_49841,N_49816);
xnor UO_636 (O_636,N_49908,N_49976);
nand UO_637 (O_637,N_49840,N_49807);
xnor UO_638 (O_638,N_49762,N_49978);
or UO_639 (O_639,N_49947,N_49872);
and UO_640 (O_640,N_49811,N_49989);
nor UO_641 (O_641,N_49887,N_49884);
nor UO_642 (O_642,N_49962,N_49941);
nor UO_643 (O_643,N_49879,N_49774);
nor UO_644 (O_644,N_49899,N_49849);
nand UO_645 (O_645,N_49936,N_49896);
nand UO_646 (O_646,N_49963,N_49871);
xor UO_647 (O_647,N_49986,N_49753);
and UO_648 (O_648,N_49993,N_49924);
xor UO_649 (O_649,N_49918,N_49981);
nand UO_650 (O_650,N_49773,N_49959);
xnor UO_651 (O_651,N_49917,N_49779);
nand UO_652 (O_652,N_49956,N_49838);
nor UO_653 (O_653,N_49980,N_49883);
xor UO_654 (O_654,N_49775,N_49814);
nor UO_655 (O_655,N_49815,N_49927);
xnor UO_656 (O_656,N_49759,N_49921);
nand UO_657 (O_657,N_49802,N_49895);
nand UO_658 (O_658,N_49844,N_49774);
and UO_659 (O_659,N_49777,N_49973);
nand UO_660 (O_660,N_49850,N_49925);
nor UO_661 (O_661,N_49948,N_49783);
nor UO_662 (O_662,N_49959,N_49761);
nand UO_663 (O_663,N_49815,N_49909);
or UO_664 (O_664,N_49936,N_49888);
nand UO_665 (O_665,N_49835,N_49797);
nand UO_666 (O_666,N_49878,N_49964);
and UO_667 (O_667,N_49928,N_49829);
nor UO_668 (O_668,N_49835,N_49981);
or UO_669 (O_669,N_49875,N_49937);
nor UO_670 (O_670,N_49998,N_49981);
nand UO_671 (O_671,N_49753,N_49808);
nand UO_672 (O_672,N_49985,N_49872);
or UO_673 (O_673,N_49774,N_49994);
nor UO_674 (O_674,N_49832,N_49852);
or UO_675 (O_675,N_49979,N_49834);
nand UO_676 (O_676,N_49852,N_49850);
nand UO_677 (O_677,N_49780,N_49938);
nand UO_678 (O_678,N_49848,N_49772);
and UO_679 (O_679,N_49868,N_49876);
nand UO_680 (O_680,N_49793,N_49854);
nor UO_681 (O_681,N_49936,N_49825);
and UO_682 (O_682,N_49949,N_49907);
nand UO_683 (O_683,N_49984,N_49780);
xor UO_684 (O_684,N_49956,N_49930);
nor UO_685 (O_685,N_49761,N_49815);
nand UO_686 (O_686,N_49753,N_49931);
xnor UO_687 (O_687,N_49756,N_49777);
nand UO_688 (O_688,N_49766,N_49855);
and UO_689 (O_689,N_49788,N_49943);
xnor UO_690 (O_690,N_49750,N_49888);
xnor UO_691 (O_691,N_49817,N_49847);
and UO_692 (O_692,N_49811,N_49839);
and UO_693 (O_693,N_49956,N_49992);
xnor UO_694 (O_694,N_49851,N_49868);
xnor UO_695 (O_695,N_49774,N_49841);
nand UO_696 (O_696,N_49750,N_49804);
or UO_697 (O_697,N_49781,N_49867);
and UO_698 (O_698,N_49829,N_49869);
nand UO_699 (O_699,N_49970,N_49882);
nor UO_700 (O_700,N_49835,N_49998);
and UO_701 (O_701,N_49837,N_49893);
nand UO_702 (O_702,N_49857,N_49846);
xor UO_703 (O_703,N_49819,N_49947);
xnor UO_704 (O_704,N_49857,N_49876);
xnor UO_705 (O_705,N_49954,N_49889);
nand UO_706 (O_706,N_49933,N_49910);
or UO_707 (O_707,N_49933,N_49835);
nand UO_708 (O_708,N_49886,N_49993);
and UO_709 (O_709,N_49808,N_49995);
nand UO_710 (O_710,N_49972,N_49971);
or UO_711 (O_711,N_49912,N_49811);
and UO_712 (O_712,N_49890,N_49900);
and UO_713 (O_713,N_49769,N_49754);
or UO_714 (O_714,N_49831,N_49754);
nand UO_715 (O_715,N_49885,N_49870);
or UO_716 (O_716,N_49996,N_49913);
nor UO_717 (O_717,N_49992,N_49787);
nor UO_718 (O_718,N_49761,N_49852);
xnor UO_719 (O_719,N_49805,N_49894);
nand UO_720 (O_720,N_49913,N_49750);
and UO_721 (O_721,N_49834,N_49890);
or UO_722 (O_722,N_49873,N_49758);
nor UO_723 (O_723,N_49852,N_49863);
nand UO_724 (O_724,N_49855,N_49825);
or UO_725 (O_725,N_49901,N_49931);
nand UO_726 (O_726,N_49948,N_49983);
xor UO_727 (O_727,N_49895,N_49804);
xnor UO_728 (O_728,N_49835,N_49927);
xnor UO_729 (O_729,N_49773,N_49912);
and UO_730 (O_730,N_49786,N_49955);
nand UO_731 (O_731,N_49997,N_49837);
nor UO_732 (O_732,N_49813,N_49962);
nand UO_733 (O_733,N_49999,N_49903);
and UO_734 (O_734,N_49760,N_49757);
and UO_735 (O_735,N_49948,N_49845);
nand UO_736 (O_736,N_49764,N_49837);
nand UO_737 (O_737,N_49956,N_49954);
nor UO_738 (O_738,N_49873,N_49853);
or UO_739 (O_739,N_49756,N_49870);
xor UO_740 (O_740,N_49941,N_49894);
nor UO_741 (O_741,N_49868,N_49921);
nand UO_742 (O_742,N_49776,N_49752);
nand UO_743 (O_743,N_49930,N_49814);
or UO_744 (O_744,N_49944,N_49953);
and UO_745 (O_745,N_49797,N_49964);
or UO_746 (O_746,N_49968,N_49890);
xnor UO_747 (O_747,N_49977,N_49810);
and UO_748 (O_748,N_49861,N_49932);
or UO_749 (O_749,N_49797,N_49965);
nor UO_750 (O_750,N_49769,N_49823);
or UO_751 (O_751,N_49894,N_49858);
xnor UO_752 (O_752,N_49991,N_49998);
or UO_753 (O_753,N_49841,N_49989);
nor UO_754 (O_754,N_49895,N_49773);
or UO_755 (O_755,N_49803,N_49987);
nor UO_756 (O_756,N_49790,N_49933);
xnor UO_757 (O_757,N_49831,N_49966);
nand UO_758 (O_758,N_49901,N_49945);
nor UO_759 (O_759,N_49789,N_49791);
or UO_760 (O_760,N_49752,N_49798);
nor UO_761 (O_761,N_49942,N_49904);
nor UO_762 (O_762,N_49890,N_49937);
xor UO_763 (O_763,N_49952,N_49772);
nor UO_764 (O_764,N_49944,N_49945);
nand UO_765 (O_765,N_49912,N_49758);
nor UO_766 (O_766,N_49795,N_49754);
nor UO_767 (O_767,N_49755,N_49787);
and UO_768 (O_768,N_49785,N_49963);
xnor UO_769 (O_769,N_49791,N_49772);
nor UO_770 (O_770,N_49944,N_49912);
nor UO_771 (O_771,N_49874,N_49972);
or UO_772 (O_772,N_49880,N_49995);
and UO_773 (O_773,N_49992,N_49764);
nor UO_774 (O_774,N_49894,N_49804);
nor UO_775 (O_775,N_49812,N_49979);
nand UO_776 (O_776,N_49930,N_49875);
nor UO_777 (O_777,N_49915,N_49801);
and UO_778 (O_778,N_49898,N_49916);
or UO_779 (O_779,N_49764,N_49955);
nand UO_780 (O_780,N_49842,N_49960);
nand UO_781 (O_781,N_49775,N_49819);
nor UO_782 (O_782,N_49868,N_49836);
nand UO_783 (O_783,N_49845,N_49766);
nor UO_784 (O_784,N_49993,N_49880);
nor UO_785 (O_785,N_49945,N_49780);
xor UO_786 (O_786,N_49793,N_49751);
and UO_787 (O_787,N_49936,N_49977);
and UO_788 (O_788,N_49938,N_49956);
and UO_789 (O_789,N_49890,N_49771);
nand UO_790 (O_790,N_49851,N_49923);
or UO_791 (O_791,N_49932,N_49854);
nor UO_792 (O_792,N_49921,N_49776);
or UO_793 (O_793,N_49784,N_49828);
nand UO_794 (O_794,N_49768,N_49947);
and UO_795 (O_795,N_49803,N_49892);
xor UO_796 (O_796,N_49781,N_49817);
nor UO_797 (O_797,N_49915,N_49919);
nor UO_798 (O_798,N_49813,N_49995);
or UO_799 (O_799,N_49754,N_49759);
and UO_800 (O_800,N_49802,N_49836);
nand UO_801 (O_801,N_49845,N_49893);
and UO_802 (O_802,N_49772,N_49817);
nor UO_803 (O_803,N_49855,N_49863);
and UO_804 (O_804,N_49926,N_49923);
or UO_805 (O_805,N_49777,N_49833);
and UO_806 (O_806,N_49915,N_49796);
nor UO_807 (O_807,N_49976,N_49794);
nand UO_808 (O_808,N_49852,N_49849);
nor UO_809 (O_809,N_49811,N_49865);
xor UO_810 (O_810,N_49882,N_49756);
nor UO_811 (O_811,N_49961,N_49952);
nor UO_812 (O_812,N_49800,N_49953);
nor UO_813 (O_813,N_49769,N_49802);
nor UO_814 (O_814,N_49945,N_49865);
xor UO_815 (O_815,N_49759,N_49867);
nand UO_816 (O_816,N_49807,N_49943);
or UO_817 (O_817,N_49978,N_49834);
nor UO_818 (O_818,N_49784,N_49829);
and UO_819 (O_819,N_49990,N_49984);
or UO_820 (O_820,N_49887,N_49989);
nand UO_821 (O_821,N_49768,N_49885);
or UO_822 (O_822,N_49907,N_49971);
or UO_823 (O_823,N_49905,N_49820);
xor UO_824 (O_824,N_49884,N_49765);
or UO_825 (O_825,N_49939,N_49819);
nand UO_826 (O_826,N_49756,N_49871);
and UO_827 (O_827,N_49796,N_49901);
and UO_828 (O_828,N_49864,N_49972);
xnor UO_829 (O_829,N_49990,N_49873);
nand UO_830 (O_830,N_49899,N_49959);
or UO_831 (O_831,N_49839,N_49954);
or UO_832 (O_832,N_49855,N_49819);
nand UO_833 (O_833,N_49991,N_49767);
xor UO_834 (O_834,N_49759,N_49945);
and UO_835 (O_835,N_49927,N_49832);
nand UO_836 (O_836,N_49775,N_49915);
nand UO_837 (O_837,N_49814,N_49983);
and UO_838 (O_838,N_49786,N_49783);
xnor UO_839 (O_839,N_49808,N_49807);
and UO_840 (O_840,N_49950,N_49944);
or UO_841 (O_841,N_49952,N_49808);
xnor UO_842 (O_842,N_49985,N_49851);
nor UO_843 (O_843,N_49762,N_49794);
nand UO_844 (O_844,N_49847,N_49808);
xnor UO_845 (O_845,N_49813,N_49998);
and UO_846 (O_846,N_49850,N_49990);
nand UO_847 (O_847,N_49912,N_49989);
and UO_848 (O_848,N_49870,N_49957);
xnor UO_849 (O_849,N_49929,N_49838);
and UO_850 (O_850,N_49931,N_49944);
xnor UO_851 (O_851,N_49984,N_49841);
nor UO_852 (O_852,N_49772,N_49978);
nor UO_853 (O_853,N_49804,N_49918);
or UO_854 (O_854,N_49796,N_49993);
nor UO_855 (O_855,N_49852,N_49886);
or UO_856 (O_856,N_49847,N_49897);
or UO_857 (O_857,N_49860,N_49864);
and UO_858 (O_858,N_49889,N_49888);
and UO_859 (O_859,N_49782,N_49982);
and UO_860 (O_860,N_49859,N_49955);
and UO_861 (O_861,N_49849,N_49940);
or UO_862 (O_862,N_49785,N_49762);
nor UO_863 (O_863,N_49771,N_49938);
xor UO_864 (O_864,N_49979,N_49839);
or UO_865 (O_865,N_49992,N_49824);
and UO_866 (O_866,N_49757,N_49877);
nor UO_867 (O_867,N_49873,N_49863);
and UO_868 (O_868,N_49875,N_49927);
nand UO_869 (O_869,N_49852,N_49877);
xor UO_870 (O_870,N_49911,N_49809);
or UO_871 (O_871,N_49859,N_49960);
or UO_872 (O_872,N_49914,N_49844);
nand UO_873 (O_873,N_49884,N_49844);
xnor UO_874 (O_874,N_49882,N_49857);
or UO_875 (O_875,N_49792,N_49762);
and UO_876 (O_876,N_49755,N_49768);
nand UO_877 (O_877,N_49835,N_49924);
xor UO_878 (O_878,N_49898,N_49838);
and UO_879 (O_879,N_49936,N_49917);
nor UO_880 (O_880,N_49946,N_49801);
nand UO_881 (O_881,N_49803,N_49906);
and UO_882 (O_882,N_49846,N_49902);
nor UO_883 (O_883,N_49776,N_49960);
xor UO_884 (O_884,N_49904,N_49752);
nor UO_885 (O_885,N_49755,N_49987);
nand UO_886 (O_886,N_49898,N_49784);
nor UO_887 (O_887,N_49761,N_49962);
and UO_888 (O_888,N_49847,N_49880);
and UO_889 (O_889,N_49996,N_49823);
or UO_890 (O_890,N_49865,N_49765);
nor UO_891 (O_891,N_49839,N_49763);
xnor UO_892 (O_892,N_49804,N_49976);
nand UO_893 (O_893,N_49841,N_49751);
and UO_894 (O_894,N_49959,N_49827);
and UO_895 (O_895,N_49855,N_49988);
and UO_896 (O_896,N_49937,N_49925);
or UO_897 (O_897,N_49947,N_49875);
xor UO_898 (O_898,N_49921,N_49830);
or UO_899 (O_899,N_49824,N_49807);
and UO_900 (O_900,N_49909,N_49916);
and UO_901 (O_901,N_49767,N_49818);
nand UO_902 (O_902,N_49891,N_49782);
or UO_903 (O_903,N_49914,N_49785);
nand UO_904 (O_904,N_49994,N_49979);
and UO_905 (O_905,N_49904,N_49911);
nor UO_906 (O_906,N_49903,N_49907);
nor UO_907 (O_907,N_49901,N_49839);
xor UO_908 (O_908,N_49810,N_49924);
nor UO_909 (O_909,N_49852,N_49759);
xnor UO_910 (O_910,N_49754,N_49996);
nand UO_911 (O_911,N_49949,N_49978);
or UO_912 (O_912,N_49756,N_49928);
nand UO_913 (O_913,N_49823,N_49902);
or UO_914 (O_914,N_49979,N_49836);
nor UO_915 (O_915,N_49781,N_49844);
xnor UO_916 (O_916,N_49815,N_49998);
nor UO_917 (O_917,N_49891,N_49813);
nor UO_918 (O_918,N_49799,N_49814);
nand UO_919 (O_919,N_49807,N_49858);
nor UO_920 (O_920,N_49793,N_49993);
nand UO_921 (O_921,N_49834,N_49846);
nor UO_922 (O_922,N_49916,N_49812);
nor UO_923 (O_923,N_49830,N_49888);
or UO_924 (O_924,N_49863,N_49937);
or UO_925 (O_925,N_49963,N_49892);
nand UO_926 (O_926,N_49818,N_49753);
and UO_927 (O_927,N_49776,N_49992);
nor UO_928 (O_928,N_49866,N_49843);
nor UO_929 (O_929,N_49864,N_49770);
or UO_930 (O_930,N_49878,N_49872);
nor UO_931 (O_931,N_49751,N_49770);
nand UO_932 (O_932,N_49859,N_49769);
nor UO_933 (O_933,N_49833,N_49753);
and UO_934 (O_934,N_49949,N_49950);
xor UO_935 (O_935,N_49859,N_49936);
nor UO_936 (O_936,N_49988,N_49956);
nor UO_937 (O_937,N_49958,N_49971);
or UO_938 (O_938,N_49978,N_49815);
nor UO_939 (O_939,N_49792,N_49955);
nand UO_940 (O_940,N_49818,N_49979);
and UO_941 (O_941,N_49814,N_49991);
and UO_942 (O_942,N_49993,N_49763);
nor UO_943 (O_943,N_49888,N_49969);
nor UO_944 (O_944,N_49834,N_49958);
nor UO_945 (O_945,N_49844,N_49991);
nand UO_946 (O_946,N_49960,N_49813);
and UO_947 (O_947,N_49913,N_49882);
or UO_948 (O_948,N_49854,N_49860);
or UO_949 (O_949,N_49856,N_49770);
or UO_950 (O_950,N_49798,N_49775);
nand UO_951 (O_951,N_49961,N_49827);
xnor UO_952 (O_952,N_49996,N_49846);
or UO_953 (O_953,N_49920,N_49757);
xor UO_954 (O_954,N_49953,N_49926);
and UO_955 (O_955,N_49773,N_49838);
and UO_956 (O_956,N_49987,N_49905);
nor UO_957 (O_957,N_49766,N_49839);
xnor UO_958 (O_958,N_49794,N_49788);
and UO_959 (O_959,N_49811,N_49949);
or UO_960 (O_960,N_49844,N_49917);
and UO_961 (O_961,N_49899,N_49907);
or UO_962 (O_962,N_49821,N_49956);
nand UO_963 (O_963,N_49761,N_49788);
nor UO_964 (O_964,N_49809,N_49947);
nor UO_965 (O_965,N_49868,N_49759);
or UO_966 (O_966,N_49793,N_49933);
nand UO_967 (O_967,N_49957,N_49948);
nand UO_968 (O_968,N_49821,N_49787);
nand UO_969 (O_969,N_49838,N_49982);
nor UO_970 (O_970,N_49953,N_49906);
xnor UO_971 (O_971,N_49802,N_49956);
nand UO_972 (O_972,N_49910,N_49751);
nand UO_973 (O_973,N_49875,N_49819);
xnor UO_974 (O_974,N_49770,N_49792);
nor UO_975 (O_975,N_49925,N_49906);
nor UO_976 (O_976,N_49796,N_49943);
and UO_977 (O_977,N_49955,N_49800);
nor UO_978 (O_978,N_49784,N_49947);
nand UO_979 (O_979,N_49892,N_49989);
and UO_980 (O_980,N_49873,N_49810);
nand UO_981 (O_981,N_49910,N_49906);
nor UO_982 (O_982,N_49841,N_49959);
or UO_983 (O_983,N_49969,N_49778);
xnor UO_984 (O_984,N_49934,N_49861);
and UO_985 (O_985,N_49941,N_49841);
nor UO_986 (O_986,N_49950,N_49953);
and UO_987 (O_987,N_49761,N_49928);
nand UO_988 (O_988,N_49782,N_49996);
and UO_989 (O_989,N_49966,N_49950);
or UO_990 (O_990,N_49887,N_49794);
and UO_991 (O_991,N_49865,N_49887);
xor UO_992 (O_992,N_49814,N_49861);
or UO_993 (O_993,N_49826,N_49830);
xor UO_994 (O_994,N_49938,N_49759);
xnor UO_995 (O_995,N_49946,N_49974);
or UO_996 (O_996,N_49751,N_49952);
nor UO_997 (O_997,N_49785,N_49770);
nor UO_998 (O_998,N_49951,N_49976);
xor UO_999 (O_999,N_49840,N_49913);
nand UO_1000 (O_1000,N_49915,N_49888);
xor UO_1001 (O_1001,N_49813,N_49763);
and UO_1002 (O_1002,N_49825,N_49921);
and UO_1003 (O_1003,N_49755,N_49775);
and UO_1004 (O_1004,N_49930,N_49759);
nand UO_1005 (O_1005,N_49866,N_49786);
or UO_1006 (O_1006,N_49969,N_49886);
or UO_1007 (O_1007,N_49822,N_49899);
nand UO_1008 (O_1008,N_49774,N_49955);
and UO_1009 (O_1009,N_49992,N_49978);
and UO_1010 (O_1010,N_49843,N_49910);
nor UO_1011 (O_1011,N_49948,N_49765);
nor UO_1012 (O_1012,N_49953,N_49995);
or UO_1013 (O_1013,N_49831,N_49994);
or UO_1014 (O_1014,N_49820,N_49825);
and UO_1015 (O_1015,N_49940,N_49846);
or UO_1016 (O_1016,N_49913,N_49983);
nor UO_1017 (O_1017,N_49765,N_49766);
nor UO_1018 (O_1018,N_49868,N_49956);
or UO_1019 (O_1019,N_49838,N_49865);
or UO_1020 (O_1020,N_49948,N_49930);
or UO_1021 (O_1021,N_49885,N_49973);
nor UO_1022 (O_1022,N_49868,N_49817);
and UO_1023 (O_1023,N_49821,N_49908);
or UO_1024 (O_1024,N_49780,N_49935);
nor UO_1025 (O_1025,N_49792,N_49863);
xnor UO_1026 (O_1026,N_49755,N_49952);
or UO_1027 (O_1027,N_49766,N_49913);
and UO_1028 (O_1028,N_49793,N_49797);
xor UO_1029 (O_1029,N_49838,N_49802);
xor UO_1030 (O_1030,N_49854,N_49753);
and UO_1031 (O_1031,N_49772,N_49850);
nand UO_1032 (O_1032,N_49925,N_49973);
nor UO_1033 (O_1033,N_49919,N_49961);
nand UO_1034 (O_1034,N_49949,N_49960);
nand UO_1035 (O_1035,N_49912,N_49772);
nand UO_1036 (O_1036,N_49872,N_49840);
nor UO_1037 (O_1037,N_49974,N_49866);
nor UO_1038 (O_1038,N_49911,N_49799);
nand UO_1039 (O_1039,N_49758,N_49767);
or UO_1040 (O_1040,N_49802,N_49967);
or UO_1041 (O_1041,N_49864,N_49913);
nor UO_1042 (O_1042,N_49961,N_49796);
nand UO_1043 (O_1043,N_49764,N_49828);
nor UO_1044 (O_1044,N_49924,N_49846);
and UO_1045 (O_1045,N_49987,N_49758);
or UO_1046 (O_1046,N_49974,N_49828);
and UO_1047 (O_1047,N_49894,N_49843);
or UO_1048 (O_1048,N_49913,N_49969);
nor UO_1049 (O_1049,N_49872,N_49956);
nand UO_1050 (O_1050,N_49843,N_49893);
xnor UO_1051 (O_1051,N_49962,N_49968);
nand UO_1052 (O_1052,N_49982,N_49929);
xnor UO_1053 (O_1053,N_49992,N_49904);
nand UO_1054 (O_1054,N_49968,N_49800);
and UO_1055 (O_1055,N_49807,N_49976);
and UO_1056 (O_1056,N_49765,N_49826);
and UO_1057 (O_1057,N_49989,N_49945);
nor UO_1058 (O_1058,N_49977,N_49770);
nor UO_1059 (O_1059,N_49922,N_49775);
xor UO_1060 (O_1060,N_49795,N_49815);
nor UO_1061 (O_1061,N_49861,N_49941);
nand UO_1062 (O_1062,N_49934,N_49798);
nand UO_1063 (O_1063,N_49783,N_49814);
nor UO_1064 (O_1064,N_49790,N_49907);
xnor UO_1065 (O_1065,N_49778,N_49913);
and UO_1066 (O_1066,N_49777,N_49926);
and UO_1067 (O_1067,N_49918,N_49781);
xnor UO_1068 (O_1068,N_49799,N_49775);
nand UO_1069 (O_1069,N_49963,N_49873);
xor UO_1070 (O_1070,N_49916,N_49826);
or UO_1071 (O_1071,N_49817,N_49879);
nand UO_1072 (O_1072,N_49764,N_49963);
xor UO_1073 (O_1073,N_49934,N_49897);
xnor UO_1074 (O_1074,N_49771,N_49784);
or UO_1075 (O_1075,N_49974,N_49774);
and UO_1076 (O_1076,N_49996,N_49861);
or UO_1077 (O_1077,N_49786,N_49879);
xor UO_1078 (O_1078,N_49955,N_49908);
xnor UO_1079 (O_1079,N_49762,N_49996);
and UO_1080 (O_1080,N_49961,N_49891);
nor UO_1081 (O_1081,N_49918,N_49992);
nand UO_1082 (O_1082,N_49825,N_49764);
or UO_1083 (O_1083,N_49906,N_49807);
nor UO_1084 (O_1084,N_49889,N_49964);
xnor UO_1085 (O_1085,N_49923,N_49804);
and UO_1086 (O_1086,N_49833,N_49894);
nor UO_1087 (O_1087,N_49974,N_49878);
and UO_1088 (O_1088,N_49980,N_49916);
nand UO_1089 (O_1089,N_49910,N_49868);
and UO_1090 (O_1090,N_49847,N_49751);
and UO_1091 (O_1091,N_49809,N_49872);
xor UO_1092 (O_1092,N_49821,N_49762);
xor UO_1093 (O_1093,N_49980,N_49804);
xnor UO_1094 (O_1094,N_49756,N_49997);
nand UO_1095 (O_1095,N_49825,N_49890);
or UO_1096 (O_1096,N_49922,N_49754);
xnor UO_1097 (O_1097,N_49810,N_49993);
xnor UO_1098 (O_1098,N_49754,N_49798);
or UO_1099 (O_1099,N_49817,N_49910);
xnor UO_1100 (O_1100,N_49884,N_49879);
xnor UO_1101 (O_1101,N_49787,N_49822);
xor UO_1102 (O_1102,N_49801,N_49796);
nand UO_1103 (O_1103,N_49975,N_49815);
and UO_1104 (O_1104,N_49862,N_49922);
nor UO_1105 (O_1105,N_49830,N_49990);
and UO_1106 (O_1106,N_49794,N_49954);
nand UO_1107 (O_1107,N_49760,N_49961);
nand UO_1108 (O_1108,N_49836,N_49792);
or UO_1109 (O_1109,N_49819,N_49831);
nand UO_1110 (O_1110,N_49945,N_49824);
and UO_1111 (O_1111,N_49987,N_49913);
nand UO_1112 (O_1112,N_49751,N_49972);
nor UO_1113 (O_1113,N_49991,N_49755);
xor UO_1114 (O_1114,N_49769,N_49822);
or UO_1115 (O_1115,N_49833,N_49752);
nand UO_1116 (O_1116,N_49963,N_49984);
nor UO_1117 (O_1117,N_49831,N_49971);
and UO_1118 (O_1118,N_49945,N_49760);
xor UO_1119 (O_1119,N_49770,N_49973);
nand UO_1120 (O_1120,N_49821,N_49954);
nor UO_1121 (O_1121,N_49997,N_49874);
and UO_1122 (O_1122,N_49989,N_49953);
xnor UO_1123 (O_1123,N_49799,N_49896);
nor UO_1124 (O_1124,N_49795,N_49827);
or UO_1125 (O_1125,N_49916,N_49768);
and UO_1126 (O_1126,N_49765,N_49915);
or UO_1127 (O_1127,N_49888,N_49883);
or UO_1128 (O_1128,N_49884,N_49930);
or UO_1129 (O_1129,N_49818,N_49911);
and UO_1130 (O_1130,N_49768,N_49846);
nor UO_1131 (O_1131,N_49857,N_49771);
nor UO_1132 (O_1132,N_49777,N_49959);
nand UO_1133 (O_1133,N_49862,N_49896);
nor UO_1134 (O_1134,N_49762,N_49802);
and UO_1135 (O_1135,N_49937,N_49855);
and UO_1136 (O_1136,N_49840,N_49924);
nor UO_1137 (O_1137,N_49846,N_49864);
or UO_1138 (O_1138,N_49828,N_49818);
xnor UO_1139 (O_1139,N_49962,N_49885);
xnor UO_1140 (O_1140,N_49896,N_49917);
nor UO_1141 (O_1141,N_49761,N_49865);
nor UO_1142 (O_1142,N_49925,N_49938);
nand UO_1143 (O_1143,N_49931,N_49980);
nand UO_1144 (O_1144,N_49847,N_49850);
nor UO_1145 (O_1145,N_49804,N_49917);
nor UO_1146 (O_1146,N_49946,N_49925);
nand UO_1147 (O_1147,N_49960,N_49973);
or UO_1148 (O_1148,N_49842,N_49964);
nand UO_1149 (O_1149,N_49968,N_49860);
nand UO_1150 (O_1150,N_49829,N_49992);
nor UO_1151 (O_1151,N_49875,N_49914);
or UO_1152 (O_1152,N_49897,N_49985);
or UO_1153 (O_1153,N_49907,N_49813);
or UO_1154 (O_1154,N_49925,N_49891);
nor UO_1155 (O_1155,N_49786,N_49931);
xor UO_1156 (O_1156,N_49904,N_49837);
nor UO_1157 (O_1157,N_49997,N_49830);
nand UO_1158 (O_1158,N_49929,N_49848);
and UO_1159 (O_1159,N_49770,N_49960);
or UO_1160 (O_1160,N_49814,N_49864);
or UO_1161 (O_1161,N_49908,N_49790);
and UO_1162 (O_1162,N_49962,N_49769);
nor UO_1163 (O_1163,N_49897,N_49803);
xor UO_1164 (O_1164,N_49753,N_49787);
xnor UO_1165 (O_1165,N_49754,N_49990);
xor UO_1166 (O_1166,N_49786,N_49788);
nand UO_1167 (O_1167,N_49982,N_49761);
nor UO_1168 (O_1168,N_49936,N_49961);
and UO_1169 (O_1169,N_49950,N_49842);
and UO_1170 (O_1170,N_49784,N_49961);
or UO_1171 (O_1171,N_49837,N_49943);
xor UO_1172 (O_1172,N_49759,N_49964);
nand UO_1173 (O_1173,N_49884,N_49889);
nor UO_1174 (O_1174,N_49936,N_49794);
xnor UO_1175 (O_1175,N_49791,N_49905);
or UO_1176 (O_1176,N_49992,N_49779);
xnor UO_1177 (O_1177,N_49895,N_49771);
or UO_1178 (O_1178,N_49851,N_49778);
and UO_1179 (O_1179,N_49890,N_49850);
and UO_1180 (O_1180,N_49820,N_49881);
or UO_1181 (O_1181,N_49872,N_49849);
xnor UO_1182 (O_1182,N_49957,N_49954);
and UO_1183 (O_1183,N_49954,N_49870);
and UO_1184 (O_1184,N_49926,N_49892);
nor UO_1185 (O_1185,N_49968,N_49908);
nand UO_1186 (O_1186,N_49999,N_49979);
nand UO_1187 (O_1187,N_49791,N_49920);
nand UO_1188 (O_1188,N_49916,N_49878);
and UO_1189 (O_1189,N_49815,N_49793);
nand UO_1190 (O_1190,N_49770,N_49999);
nor UO_1191 (O_1191,N_49850,N_49954);
xnor UO_1192 (O_1192,N_49759,N_49807);
nor UO_1193 (O_1193,N_49848,N_49915);
nor UO_1194 (O_1194,N_49956,N_49971);
and UO_1195 (O_1195,N_49774,N_49897);
nor UO_1196 (O_1196,N_49856,N_49897);
nor UO_1197 (O_1197,N_49900,N_49870);
nand UO_1198 (O_1198,N_49830,N_49849);
xor UO_1199 (O_1199,N_49866,N_49851);
nor UO_1200 (O_1200,N_49845,N_49971);
or UO_1201 (O_1201,N_49799,N_49867);
nand UO_1202 (O_1202,N_49938,N_49856);
nor UO_1203 (O_1203,N_49759,N_49941);
or UO_1204 (O_1204,N_49886,N_49905);
nand UO_1205 (O_1205,N_49890,N_49943);
or UO_1206 (O_1206,N_49906,N_49999);
or UO_1207 (O_1207,N_49955,N_49916);
xnor UO_1208 (O_1208,N_49836,N_49992);
xor UO_1209 (O_1209,N_49798,N_49777);
xnor UO_1210 (O_1210,N_49754,N_49779);
or UO_1211 (O_1211,N_49901,N_49781);
and UO_1212 (O_1212,N_49935,N_49817);
or UO_1213 (O_1213,N_49838,N_49786);
or UO_1214 (O_1214,N_49829,N_49934);
xnor UO_1215 (O_1215,N_49877,N_49929);
nor UO_1216 (O_1216,N_49856,N_49952);
nand UO_1217 (O_1217,N_49767,N_49873);
nor UO_1218 (O_1218,N_49799,N_49806);
and UO_1219 (O_1219,N_49950,N_49865);
nand UO_1220 (O_1220,N_49817,N_49864);
xor UO_1221 (O_1221,N_49992,N_49837);
xnor UO_1222 (O_1222,N_49856,N_49916);
xnor UO_1223 (O_1223,N_49812,N_49791);
nand UO_1224 (O_1224,N_49871,N_49946);
nand UO_1225 (O_1225,N_49802,N_49941);
nand UO_1226 (O_1226,N_49939,N_49910);
or UO_1227 (O_1227,N_49888,N_49788);
and UO_1228 (O_1228,N_49831,N_49931);
nand UO_1229 (O_1229,N_49976,N_49894);
xor UO_1230 (O_1230,N_49862,N_49848);
or UO_1231 (O_1231,N_49793,N_49979);
or UO_1232 (O_1232,N_49860,N_49989);
xor UO_1233 (O_1233,N_49881,N_49824);
or UO_1234 (O_1234,N_49901,N_49988);
nor UO_1235 (O_1235,N_49832,N_49910);
nand UO_1236 (O_1236,N_49954,N_49938);
and UO_1237 (O_1237,N_49987,N_49951);
nor UO_1238 (O_1238,N_49895,N_49750);
nand UO_1239 (O_1239,N_49789,N_49800);
nand UO_1240 (O_1240,N_49842,N_49983);
or UO_1241 (O_1241,N_49823,N_49993);
or UO_1242 (O_1242,N_49964,N_49821);
and UO_1243 (O_1243,N_49909,N_49772);
and UO_1244 (O_1244,N_49900,N_49867);
or UO_1245 (O_1245,N_49983,N_49756);
nand UO_1246 (O_1246,N_49921,N_49946);
or UO_1247 (O_1247,N_49951,N_49989);
and UO_1248 (O_1248,N_49762,N_49895);
nor UO_1249 (O_1249,N_49915,N_49834);
nor UO_1250 (O_1250,N_49787,N_49812);
and UO_1251 (O_1251,N_49882,N_49764);
nand UO_1252 (O_1252,N_49803,N_49985);
xnor UO_1253 (O_1253,N_49799,N_49986);
nand UO_1254 (O_1254,N_49905,N_49770);
and UO_1255 (O_1255,N_49829,N_49765);
nor UO_1256 (O_1256,N_49979,N_49785);
or UO_1257 (O_1257,N_49989,N_49932);
or UO_1258 (O_1258,N_49930,N_49955);
nand UO_1259 (O_1259,N_49865,N_49933);
xor UO_1260 (O_1260,N_49873,N_49936);
nor UO_1261 (O_1261,N_49930,N_49813);
nor UO_1262 (O_1262,N_49902,N_49892);
nand UO_1263 (O_1263,N_49753,N_49910);
nand UO_1264 (O_1264,N_49794,N_49952);
or UO_1265 (O_1265,N_49861,N_49820);
nor UO_1266 (O_1266,N_49855,N_49769);
xor UO_1267 (O_1267,N_49927,N_49870);
nand UO_1268 (O_1268,N_49833,N_49975);
nand UO_1269 (O_1269,N_49853,N_49765);
and UO_1270 (O_1270,N_49770,N_49901);
or UO_1271 (O_1271,N_49837,N_49922);
or UO_1272 (O_1272,N_49917,N_49847);
or UO_1273 (O_1273,N_49888,N_49971);
nand UO_1274 (O_1274,N_49809,N_49828);
or UO_1275 (O_1275,N_49861,N_49923);
xor UO_1276 (O_1276,N_49882,N_49798);
nor UO_1277 (O_1277,N_49822,N_49842);
or UO_1278 (O_1278,N_49955,N_49892);
and UO_1279 (O_1279,N_49828,N_49822);
and UO_1280 (O_1280,N_49896,N_49930);
or UO_1281 (O_1281,N_49978,N_49893);
nor UO_1282 (O_1282,N_49942,N_49964);
xor UO_1283 (O_1283,N_49818,N_49797);
and UO_1284 (O_1284,N_49790,N_49803);
nand UO_1285 (O_1285,N_49885,N_49963);
nor UO_1286 (O_1286,N_49873,N_49893);
xnor UO_1287 (O_1287,N_49853,N_49982);
or UO_1288 (O_1288,N_49958,N_49983);
nor UO_1289 (O_1289,N_49758,N_49893);
and UO_1290 (O_1290,N_49858,N_49802);
and UO_1291 (O_1291,N_49899,N_49909);
or UO_1292 (O_1292,N_49871,N_49856);
or UO_1293 (O_1293,N_49901,N_49766);
xor UO_1294 (O_1294,N_49907,N_49885);
and UO_1295 (O_1295,N_49894,N_49781);
and UO_1296 (O_1296,N_49910,N_49886);
and UO_1297 (O_1297,N_49853,N_49956);
nor UO_1298 (O_1298,N_49830,N_49954);
or UO_1299 (O_1299,N_49765,N_49880);
nand UO_1300 (O_1300,N_49770,N_49753);
or UO_1301 (O_1301,N_49898,N_49751);
nor UO_1302 (O_1302,N_49963,N_49919);
or UO_1303 (O_1303,N_49957,N_49969);
and UO_1304 (O_1304,N_49818,N_49859);
and UO_1305 (O_1305,N_49817,N_49900);
and UO_1306 (O_1306,N_49853,N_49939);
nor UO_1307 (O_1307,N_49762,N_49994);
and UO_1308 (O_1308,N_49841,N_49970);
nor UO_1309 (O_1309,N_49958,N_49976);
and UO_1310 (O_1310,N_49756,N_49802);
nor UO_1311 (O_1311,N_49997,N_49947);
nand UO_1312 (O_1312,N_49866,N_49886);
nor UO_1313 (O_1313,N_49767,N_49863);
or UO_1314 (O_1314,N_49902,N_49760);
or UO_1315 (O_1315,N_49875,N_49892);
nand UO_1316 (O_1316,N_49917,N_49817);
or UO_1317 (O_1317,N_49771,N_49845);
xor UO_1318 (O_1318,N_49911,N_49842);
xor UO_1319 (O_1319,N_49799,N_49897);
nor UO_1320 (O_1320,N_49886,N_49954);
nor UO_1321 (O_1321,N_49806,N_49791);
or UO_1322 (O_1322,N_49874,N_49986);
nand UO_1323 (O_1323,N_49899,N_49895);
nor UO_1324 (O_1324,N_49804,N_49822);
nor UO_1325 (O_1325,N_49953,N_49976);
or UO_1326 (O_1326,N_49855,N_49857);
nor UO_1327 (O_1327,N_49813,N_49889);
and UO_1328 (O_1328,N_49785,N_49918);
nand UO_1329 (O_1329,N_49757,N_49968);
nand UO_1330 (O_1330,N_49852,N_49830);
nor UO_1331 (O_1331,N_49772,N_49939);
nor UO_1332 (O_1332,N_49769,N_49856);
and UO_1333 (O_1333,N_49865,N_49944);
and UO_1334 (O_1334,N_49984,N_49910);
and UO_1335 (O_1335,N_49760,N_49963);
and UO_1336 (O_1336,N_49936,N_49854);
nand UO_1337 (O_1337,N_49904,N_49825);
nand UO_1338 (O_1338,N_49872,N_49835);
nor UO_1339 (O_1339,N_49948,N_49884);
nor UO_1340 (O_1340,N_49878,N_49912);
or UO_1341 (O_1341,N_49921,N_49952);
and UO_1342 (O_1342,N_49937,N_49800);
xor UO_1343 (O_1343,N_49873,N_49847);
xnor UO_1344 (O_1344,N_49859,N_49895);
xor UO_1345 (O_1345,N_49816,N_49943);
or UO_1346 (O_1346,N_49854,N_49983);
or UO_1347 (O_1347,N_49932,N_49933);
nand UO_1348 (O_1348,N_49963,N_49912);
xor UO_1349 (O_1349,N_49988,N_49905);
nor UO_1350 (O_1350,N_49854,N_49759);
nor UO_1351 (O_1351,N_49768,N_49881);
xor UO_1352 (O_1352,N_49788,N_49959);
and UO_1353 (O_1353,N_49905,N_49873);
xor UO_1354 (O_1354,N_49995,N_49922);
or UO_1355 (O_1355,N_49868,N_49933);
xnor UO_1356 (O_1356,N_49936,N_49893);
nor UO_1357 (O_1357,N_49767,N_49785);
or UO_1358 (O_1358,N_49782,N_49875);
or UO_1359 (O_1359,N_49975,N_49807);
or UO_1360 (O_1360,N_49958,N_49855);
or UO_1361 (O_1361,N_49929,N_49926);
nand UO_1362 (O_1362,N_49759,N_49900);
and UO_1363 (O_1363,N_49854,N_49976);
nand UO_1364 (O_1364,N_49827,N_49823);
or UO_1365 (O_1365,N_49954,N_49790);
nand UO_1366 (O_1366,N_49955,N_49881);
nor UO_1367 (O_1367,N_49843,N_49945);
or UO_1368 (O_1368,N_49998,N_49945);
or UO_1369 (O_1369,N_49778,N_49878);
xnor UO_1370 (O_1370,N_49788,N_49798);
xnor UO_1371 (O_1371,N_49879,N_49923);
and UO_1372 (O_1372,N_49791,N_49895);
and UO_1373 (O_1373,N_49957,N_49939);
nor UO_1374 (O_1374,N_49951,N_49871);
or UO_1375 (O_1375,N_49954,N_49862);
xor UO_1376 (O_1376,N_49782,N_49861);
and UO_1377 (O_1377,N_49903,N_49976);
xnor UO_1378 (O_1378,N_49845,N_49892);
and UO_1379 (O_1379,N_49790,N_49923);
or UO_1380 (O_1380,N_49766,N_49904);
nand UO_1381 (O_1381,N_49949,N_49803);
or UO_1382 (O_1382,N_49806,N_49771);
nor UO_1383 (O_1383,N_49999,N_49978);
xor UO_1384 (O_1384,N_49858,N_49859);
nand UO_1385 (O_1385,N_49760,N_49787);
and UO_1386 (O_1386,N_49832,N_49947);
nor UO_1387 (O_1387,N_49990,N_49958);
xnor UO_1388 (O_1388,N_49969,N_49754);
xor UO_1389 (O_1389,N_49829,N_49836);
and UO_1390 (O_1390,N_49915,N_49899);
and UO_1391 (O_1391,N_49932,N_49849);
and UO_1392 (O_1392,N_49926,N_49903);
nand UO_1393 (O_1393,N_49794,N_49999);
and UO_1394 (O_1394,N_49772,N_49775);
xor UO_1395 (O_1395,N_49822,N_49774);
xnor UO_1396 (O_1396,N_49984,N_49843);
nand UO_1397 (O_1397,N_49799,N_49957);
xnor UO_1398 (O_1398,N_49883,N_49781);
or UO_1399 (O_1399,N_49766,N_49873);
xor UO_1400 (O_1400,N_49810,N_49916);
xor UO_1401 (O_1401,N_49843,N_49880);
nor UO_1402 (O_1402,N_49973,N_49979);
or UO_1403 (O_1403,N_49851,N_49926);
nor UO_1404 (O_1404,N_49980,N_49872);
and UO_1405 (O_1405,N_49798,N_49817);
or UO_1406 (O_1406,N_49931,N_49985);
nor UO_1407 (O_1407,N_49861,N_49868);
nand UO_1408 (O_1408,N_49872,N_49944);
xnor UO_1409 (O_1409,N_49790,N_49851);
nand UO_1410 (O_1410,N_49760,N_49912);
and UO_1411 (O_1411,N_49839,N_49933);
or UO_1412 (O_1412,N_49830,N_49858);
or UO_1413 (O_1413,N_49902,N_49896);
xor UO_1414 (O_1414,N_49919,N_49952);
nand UO_1415 (O_1415,N_49837,N_49972);
and UO_1416 (O_1416,N_49823,N_49901);
or UO_1417 (O_1417,N_49959,N_49912);
nor UO_1418 (O_1418,N_49793,N_49762);
nor UO_1419 (O_1419,N_49929,N_49843);
and UO_1420 (O_1420,N_49861,N_49830);
or UO_1421 (O_1421,N_49990,N_49863);
nand UO_1422 (O_1422,N_49907,N_49781);
or UO_1423 (O_1423,N_49871,N_49860);
and UO_1424 (O_1424,N_49872,N_49868);
nor UO_1425 (O_1425,N_49917,N_49971);
nand UO_1426 (O_1426,N_49928,N_49927);
xor UO_1427 (O_1427,N_49910,N_49838);
xor UO_1428 (O_1428,N_49923,N_49769);
xnor UO_1429 (O_1429,N_49939,N_49898);
nand UO_1430 (O_1430,N_49876,N_49933);
xor UO_1431 (O_1431,N_49822,N_49912);
and UO_1432 (O_1432,N_49894,N_49854);
and UO_1433 (O_1433,N_49795,N_49861);
xnor UO_1434 (O_1434,N_49923,N_49768);
or UO_1435 (O_1435,N_49895,N_49925);
xnor UO_1436 (O_1436,N_49978,N_49759);
nand UO_1437 (O_1437,N_49829,N_49899);
or UO_1438 (O_1438,N_49959,N_49888);
xnor UO_1439 (O_1439,N_49809,N_49999);
nand UO_1440 (O_1440,N_49875,N_49841);
or UO_1441 (O_1441,N_49941,N_49751);
or UO_1442 (O_1442,N_49773,N_49930);
and UO_1443 (O_1443,N_49781,N_49871);
or UO_1444 (O_1444,N_49862,N_49813);
or UO_1445 (O_1445,N_49836,N_49815);
or UO_1446 (O_1446,N_49951,N_49825);
nand UO_1447 (O_1447,N_49829,N_49959);
or UO_1448 (O_1448,N_49776,N_49919);
or UO_1449 (O_1449,N_49817,N_49905);
or UO_1450 (O_1450,N_49994,N_49914);
nor UO_1451 (O_1451,N_49756,N_49783);
xnor UO_1452 (O_1452,N_49877,N_49966);
nand UO_1453 (O_1453,N_49759,N_49813);
nor UO_1454 (O_1454,N_49981,N_49967);
xor UO_1455 (O_1455,N_49790,N_49868);
nand UO_1456 (O_1456,N_49883,N_49771);
xnor UO_1457 (O_1457,N_49791,N_49981);
and UO_1458 (O_1458,N_49818,N_49833);
nand UO_1459 (O_1459,N_49797,N_49975);
nor UO_1460 (O_1460,N_49851,N_49757);
xnor UO_1461 (O_1461,N_49943,N_49958);
xnor UO_1462 (O_1462,N_49888,N_49774);
xnor UO_1463 (O_1463,N_49783,N_49886);
nand UO_1464 (O_1464,N_49911,N_49813);
and UO_1465 (O_1465,N_49763,N_49805);
and UO_1466 (O_1466,N_49759,N_49927);
and UO_1467 (O_1467,N_49751,N_49960);
nor UO_1468 (O_1468,N_49979,N_49989);
or UO_1469 (O_1469,N_49930,N_49783);
or UO_1470 (O_1470,N_49778,N_49957);
and UO_1471 (O_1471,N_49862,N_49855);
xnor UO_1472 (O_1472,N_49879,N_49934);
nor UO_1473 (O_1473,N_49850,N_49860);
xor UO_1474 (O_1474,N_49900,N_49779);
or UO_1475 (O_1475,N_49909,N_49895);
and UO_1476 (O_1476,N_49925,N_49980);
or UO_1477 (O_1477,N_49812,N_49898);
and UO_1478 (O_1478,N_49901,N_49882);
and UO_1479 (O_1479,N_49860,N_49862);
or UO_1480 (O_1480,N_49772,N_49801);
nand UO_1481 (O_1481,N_49960,N_49942);
nand UO_1482 (O_1482,N_49829,N_49809);
and UO_1483 (O_1483,N_49925,N_49820);
xor UO_1484 (O_1484,N_49970,N_49803);
nor UO_1485 (O_1485,N_49983,N_49835);
nand UO_1486 (O_1486,N_49790,N_49811);
xnor UO_1487 (O_1487,N_49827,N_49778);
or UO_1488 (O_1488,N_49902,N_49873);
xor UO_1489 (O_1489,N_49842,N_49782);
xor UO_1490 (O_1490,N_49873,N_49992);
xor UO_1491 (O_1491,N_49857,N_49773);
xor UO_1492 (O_1492,N_49873,N_49819);
xor UO_1493 (O_1493,N_49968,N_49778);
nand UO_1494 (O_1494,N_49985,N_49883);
nand UO_1495 (O_1495,N_49962,N_49940);
nor UO_1496 (O_1496,N_49750,N_49945);
and UO_1497 (O_1497,N_49801,N_49957);
and UO_1498 (O_1498,N_49928,N_49911);
xor UO_1499 (O_1499,N_49819,N_49867);
xnor UO_1500 (O_1500,N_49925,N_49827);
or UO_1501 (O_1501,N_49964,N_49830);
or UO_1502 (O_1502,N_49969,N_49837);
nor UO_1503 (O_1503,N_49905,N_49792);
or UO_1504 (O_1504,N_49938,N_49806);
xnor UO_1505 (O_1505,N_49800,N_49859);
nand UO_1506 (O_1506,N_49909,N_49809);
and UO_1507 (O_1507,N_49963,N_49895);
xnor UO_1508 (O_1508,N_49964,N_49817);
xor UO_1509 (O_1509,N_49796,N_49810);
or UO_1510 (O_1510,N_49826,N_49825);
nor UO_1511 (O_1511,N_49766,N_49926);
xor UO_1512 (O_1512,N_49985,N_49852);
nand UO_1513 (O_1513,N_49808,N_49853);
xor UO_1514 (O_1514,N_49853,N_49847);
nor UO_1515 (O_1515,N_49890,N_49941);
or UO_1516 (O_1516,N_49758,N_49935);
and UO_1517 (O_1517,N_49946,N_49767);
nand UO_1518 (O_1518,N_49845,N_49923);
nand UO_1519 (O_1519,N_49949,N_49995);
nor UO_1520 (O_1520,N_49837,N_49910);
and UO_1521 (O_1521,N_49770,N_49858);
nor UO_1522 (O_1522,N_49954,N_49852);
nand UO_1523 (O_1523,N_49863,N_49968);
and UO_1524 (O_1524,N_49967,N_49956);
xor UO_1525 (O_1525,N_49924,N_49833);
and UO_1526 (O_1526,N_49903,N_49918);
nor UO_1527 (O_1527,N_49980,N_49876);
nand UO_1528 (O_1528,N_49799,N_49838);
or UO_1529 (O_1529,N_49782,N_49852);
nand UO_1530 (O_1530,N_49785,N_49765);
and UO_1531 (O_1531,N_49865,N_49837);
xnor UO_1532 (O_1532,N_49840,N_49931);
and UO_1533 (O_1533,N_49799,N_49829);
and UO_1534 (O_1534,N_49897,N_49852);
or UO_1535 (O_1535,N_49945,N_49761);
nand UO_1536 (O_1536,N_49785,N_49813);
xor UO_1537 (O_1537,N_49919,N_49840);
xnor UO_1538 (O_1538,N_49970,N_49943);
and UO_1539 (O_1539,N_49995,N_49896);
and UO_1540 (O_1540,N_49839,N_49816);
nor UO_1541 (O_1541,N_49817,N_49898);
nor UO_1542 (O_1542,N_49956,N_49989);
xor UO_1543 (O_1543,N_49801,N_49933);
nand UO_1544 (O_1544,N_49789,N_49962);
xnor UO_1545 (O_1545,N_49823,N_49961);
nand UO_1546 (O_1546,N_49770,N_49893);
xor UO_1547 (O_1547,N_49951,N_49923);
nor UO_1548 (O_1548,N_49925,N_49889);
nor UO_1549 (O_1549,N_49881,N_49949);
and UO_1550 (O_1550,N_49841,N_49982);
xor UO_1551 (O_1551,N_49814,N_49751);
and UO_1552 (O_1552,N_49991,N_49764);
and UO_1553 (O_1553,N_49889,N_49907);
xnor UO_1554 (O_1554,N_49789,N_49953);
xnor UO_1555 (O_1555,N_49900,N_49784);
and UO_1556 (O_1556,N_49928,N_49910);
nand UO_1557 (O_1557,N_49947,N_49879);
or UO_1558 (O_1558,N_49989,N_49754);
and UO_1559 (O_1559,N_49781,N_49806);
or UO_1560 (O_1560,N_49927,N_49794);
nor UO_1561 (O_1561,N_49993,N_49851);
xnor UO_1562 (O_1562,N_49990,N_49997);
nor UO_1563 (O_1563,N_49786,N_49971);
nor UO_1564 (O_1564,N_49997,N_49946);
and UO_1565 (O_1565,N_49819,N_49810);
or UO_1566 (O_1566,N_49763,N_49753);
and UO_1567 (O_1567,N_49933,N_49789);
xnor UO_1568 (O_1568,N_49953,N_49952);
or UO_1569 (O_1569,N_49751,N_49943);
nor UO_1570 (O_1570,N_49946,N_49885);
and UO_1571 (O_1571,N_49888,N_49965);
xor UO_1572 (O_1572,N_49964,N_49810);
or UO_1573 (O_1573,N_49787,N_49829);
or UO_1574 (O_1574,N_49972,N_49826);
nand UO_1575 (O_1575,N_49887,N_49924);
nor UO_1576 (O_1576,N_49937,N_49885);
or UO_1577 (O_1577,N_49917,N_49828);
nor UO_1578 (O_1578,N_49837,N_49875);
xor UO_1579 (O_1579,N_49753,N_49996);
and UO_1580 (O_1580,N_49814,N_49829);
nor UO_1581 (O_1581,N_49763,N_49957);
nor UO_1582 (O_1582,N_49942,N_49755);
xnor UO_1583 (O_1583,N_49752,N_49842);
nor UO_1584 (O_1584,N_49849,N_49835);
or UO_1585 (O_1585,N_49913,N_49867);
nand UO_1586 (O_1586,N_49892,N_49777);
xor UO_1587 (O_1587,N_49848,N_49963);
xnor UO_1588 (O_1588,N_49877,N_49815);
xor UO_1589 (O_1589,N_49907,N_49843);
nand UO_1590 (O_1590,N_49936,N_49972);
xnor UO_1591 (O_1591,N_49789,N_49938);
nor UO_1592 (O_1592,N_49850,N_49952);
and UO_1593 (O_1593,N_49990,N_49885);
nand UO_1594 (O_1594,N_49754,N_49941);
and UO_1595 (O_1595,N_49937,N_49870);
nor UO_1596 (O_1596,N_49805,N_49806);
xor UO_1597 (O_1597,N_49842,N_49916);
nor UO_1598 (O_1598,N_49750,N_49826);
nand UO_1599 (O_1599,N_49828,N_49855);
or UO_1600 (O_1600,N_49873,N_49930);
nand UO_1601 (O_1601,N_49936,N_49982);
nor UO_1602 (O_1602,N_49842,N_49851);
or UO_1603 (O_1603,N_49976,N_49869);
nand UO_1604 (O_1604,N_49834,N_49900);
xor UO_1605 (O_1605,N_49908,N_49869);
or UO_1606 (O_1606,N_49919,N_49779);
nor UO_1607 (O_1607,N_49988,N_49904);
and UO_1608 (O_1608,N_49937,N_49804);
or UO_1609 (O_1609,N_49790,N_49949);
nor UO_1610 (O_1610,N_49891,N_49890);
nor UO_1611 (O_1611,N_49884,N_49963);
xor UO_1612 (O_1612,N_49894,N_49842);
nor UO_1613 (O_1613,N_49790,N_49802);
and UO_1614 (O_1614,N_49837,N_49790);
xor UO_1615 (O_1615,N_49989,N_49935);
nand UO_1616 (O_1616,N_49788,N_49814);
and UO_1617 (O_1617,N_49774,N_49998);
nor UO_1618 (O_1618,N_49879,N_49773);
xor UO_1619 (O_1619,N_49950,N_49816);
nor UO_1620 (O_1620,N_49791,N_49932);
nor UO_1621 (O_1621,N_49936,N_49929);
or UO_1622 (O_1622,N_49779,N_49810);
nor UO_1623 (O_1623,N_49864,N_49927);
nor UO_1624 (O_1624,N_49994,N_49750);
xor UO_1625 (O_1625,N_49771,N_49866);
xnor UO_1626 (O_1626,N_49775,N_49993);
and UO_1627 (O_1627,N_49909,N_49750);
or UO_1628 (O_1628,N_49837,N_49938);
nor UO_1629 (O_1629,N_49750,N_49836);
xnor UO_1630 (O_1630,N_49757,N_49777);
and UO_1631 (O_1631,N_49982,N_49995);
nor UO_1632 (O_1632,N_49773,N_49922);
nor UO_1633 (O_1633,N_49799,N_49864);
nor UO_1634 (O_1634,N_49983,N_49916);
nand UO_1635 (O_1635,N_49949,N_49823);
nand UO_1636 (O_1636,N_49926,N_49813);
nor UO_1637 (O_1637,N_49821,N_49795);
or UO_1638 (O_1638,N_49968,N_49817);
nor UO_1639 (O_1639,N_49888,N_49786);
nor UO_1640 (O_1640,N_49801,N_49854);
nand UO_1641 (O_1641,N_49885,N_49951);
xnor UO_1642 (O_1642,N_49913,N_49830);
or UO_1643 (O_1643,N_49815,N_49835);
nand UO_1644 (O_1644,N_49842,N_49791);
nand UO_1645 (O_1645,N_49947,N_49889);
nand UO_1646 (O_1646,N_49960,N_49975);
nand UO_1647 (O_1647,N_49810,N_49965);
xor UO_1648 (O_1648,N_49983,N_49795);
nand UO_1649 (O_1649,N_49836,N_49803);
or UO_1650 (O_1650,N_49797,N_49894);
nor UO_1651 (O_1651,N_49858,N_49984);
nor UO_1652 (O_1652,N_49979,N_49889);
xor UO_1653 (O_1653,N_49803,N_49764);
xor UO_1654 (O_1654,N_49975,N_49931);
and UO_1655 (O_1655,N_49916,N_49756);
nand UO_1656 (O_1656,N_49954,N_49949);
nand UO_1657 (O_1657,N_49974,N_49803);
or UO_1658 (O_1658,N_49822,N_49770);
or UO_1659 (O_1659,N_49813,N_49938);
or UO_1660 (O_1660,N_49950,N_49873);
nor UO_1661 (O_1661,N_49898,N_49858);
and UO_1662 (O_1662,N_49989,N_49954);
and UO_1663 (O_1663,N_49815,N_49781);
and UO_1664 (O_1664,N_49988,N_49935);
nor UO_1665 (O_1665,N_49816,N_49815);
nor UO_1666 (O_1666,N_49909,N_49902);
and UO_1667 (O_1667,N_49891,N_49985);
xnor UO_1668 (O_1668,N_49931,N_49838);
and UO_1669 (O_1669,N_49776,N_49831);
xnor UO_1670 (O_1670,N_49965,N_49920);
nor UO_1671 (O_1671,N_49810,N_49906);
or UO_1672 (O_1672,N_49893,N_49928);
nor UO_1673 (O_1673,N_49879,N_49875);
and UO_1674 (O_1674,N_49966,N_49979);
or UO_1675 (O_1675,N_49751,N_49977);
or UO_1676 (O_1676,N_49942,N_49982);
and UO_1677 (O_1677,N_49935,N_49753);
nand UO_1678 (O_1678,N_49987,N_49979);
nor UO_1679 (O_1679,N_49768,N_49924);
or UO_1680 (O_1680,N_49817,N_49981);
nand UO_1681 (O_1681,N_49875,N_49787);
nor UO_1682 (O_1682,N_49991,N_49938);
nor UO_1683 (O_1683,N_49820,N_49953);
nor UO_1684 (O_1684,N_49924,N_49926);
nor UO_1685 (O_1685,N_49837,N_49964);
nand UO_1686 (O_1686,N_49787,N_49801);
and UO_1687 (O_1687,N_49763,N_49785);
or UO_1688 (O_1688,N_49975,N_49830);
or UO_1689 (O_1689,N_49993,N_49876);
nor UO_1690 (O_1690,N_49918,N_49880);
xor UO_1691 (O_1691,N_49873,N_49964);
nor UO_1692 (O_1692,N_49884,N_49798);
and UO_1693 (O_1693,N_49898,N_49792);
xor UO_1694 (O_1694,N_49912,N_49836);
nand UO_1695 (O_1695,N_49995,N_49888);
nand UO_1696 (O_1696,N_49998,N_49788);
xor UO_1697 (O_1697,N_49757,N_49837);
or UO_1698 (O_1698,N_49765,N_49832);
xor UO_1699 (O_1699,N_49791,N_49891);
and UO_1700 (O_1700,N_49956,N_49771);
or UO_1701 (O_1701,N_49951,N_49981);
or UO_1702 (O_1702,N_49857,N_49770);
nor UO_1703 (O_1703,N_49914,N_49907);
or UO_1704 (O_1704,N_49994,N_49913);
xor UO_1705 (O_1705,N_49849,N_49846);
and UO_1706 (O_1706,N_49972,N_49750);
and UO_1707 (O_1707,N_49952,N_49889);
nand UO_1708 (O_1708,N_49904,N_49789);
nand UO_1709 (O_1709,N_49801,N_49972);
or UO_1710 (O_1710,N_49908,N_49983);
nor UO_1711 (O_1711,N_49811,N_49957);
xor UO_1712 (O_1712,N_49835,N_49794);
nor UO_1713 (O_1713,N_49782,N_49969);
xnor UO_1714 (O_1714,N_49882,N_49817);
xor UO_1715 (O_1715,N_49859,N_49891);
xnor UO_1716 (O_1716,N_49941,N_49831);
or UO_1717 (O_1717,N_49986,N_49801);
and UO_1718 (O_1718,N_49759,N_49962);
and UO_1719 (O_1719,N_49967,N_49789);
nor UO_1720 (O_1720,N_49888,N_49966);
or UO_1721 (O_1721,N_49968,N_49866);
xor UO_1722 (O_1722,N_49907,N_49987);
or UO_1723 (O_1723,N_49961,N_49943);
and UO_1724 (O_1724,N_49780,N_49869);
and UO_1725 (O_1725,N_49792,N_49883);
xnor UO_1726 (O_1726,N_49972,N_49992);
xor UO_1727 (O_1727,N_49860,N_49970);
and UO_1728 (O_1728,N_49901,N_49846);
xor UO_1729 (O_1729,N_49964,N_49831);
and UO_1730 (O_1730,N_49899,N_49996);
xnor UO_1731 (O_1731,N_49912,N_49894);
xor UO_1732 (O_1732,N_49964,N_49909);
xnor UO_1733 (O_1733,N_49768,N_49932);
and UO_1734 (O_1734,N_49770,N_49888);
or UO_1735 (O_1735,N_49756,N_49877);
xnor UO_1736 (O_1736,N_49798,N_49878);
and UO_1737 (O_1737,N_49801,N_49752);
nor UO_1738 (O_1738,N_49941,N_49776);
nor UO_1739 (O_1739,N_49914,N_49962);
nor UO_1740 (O_1740,N_49918,N_49782);
xnor UO_1741 (O_1741,N_49979,N_49794);
xnor UO_1742 (O_1742,N_49787,N_49795);
nor UO_1743 (O_1743,N_49812,N_49918);
nand UO_1744 (O_1744,N_49750,N_49823);
nand UO_1745 (O_1745,N_49866,N_49837);
nand UO_1746 (O_1746,N_49780,N_49907);
and UO_1747 (O_1747,N_49774,N_49757);
and UO_1748 (O_1748,N_49853,N_49948);
xnor UO_1749 (O_1749,N_49943,N_49865);
nor UO_1750 (O_1750,N_49920,N_49925);
nand UO_1751 (O_1751,N_49812,N_49785);
xnor UO_1752 (O_1752,N_49889,N_49912);
nor UO_1753 (O_1753,N_49780,N_49992);
xnor UO_1754 (O_1754,N_49903,N_49792);
and UO_1755 (O_1755,N_49855,N_49822);
xor UO_1756 (O_1756,N_49840,N_49854);
nor UO_1757 (O_1757,N_49871,N_49768);
xnor UO_1758 (O_1758,N_49854,N_49934);
nor UO_1759 (O_1759,N_49846,N_49976);
and UO_1760 (O_1760,N_49773,N_49872);
xnor UO_1761 (O_1761,N_49893,N_49856);
or UO_1762 (O_1762,N_49950,N_49916);
and UO_1763 (O_1763,N_49860,N_49845);
nand UO_1764 (O_1764,N_49942,N_49857);
nor UO_1765 (O_1765,N_49813,N_49951);
and UO_1766 (O_1766,N_49994,N_49884);
nand UO_1767 (O_1767,N_49948,N_49833);
and UO_1768 (O_1768,N_49866,N_49914);
xor UO_1769 (O_1769,N_49756,N_49923);
and UO_1770 (O_1770,N_49974,N_49891);
or UO_1771 (O_1771,N_49975,N_49988);
nor UO_1772 (O_1772,N_49771,N_49927);
and UO_1773 (O_1773,N_49945,N_49925);
or UO_1774 (O_1774,N_49875,N_49956);
xor UO_1775 (O_1775,N_49866,N_49796);
and UO_1776 (O_1776,N_49802,N_49916);
nand UO_1777 (O_1777,N_49798,N_49954);
xnor UO_1778 (O_1778,N_49923,N_49860);
nor UO_1779 (O_1779,N_49966,N_49908);
and UO_1780 (O_1780,N_49975,N_49801);
nand UO_1781 (O_1781,N_49869,N_49953);
nand UO_1782 (O_1782,N_49752,N_49870);
and UO_1783 (O_1783,N_49960,N_49881);
and UO_1784 (O_1784,N_49751,N_49763);
xor UO_1785 (O_1785,N_49889,N_49761);
and UO_1786 (O_1786,N_49777,N_49890);
and UO_1787 (O_1787,N_49890,N_49892);
xor UO_1788 (O_1788,N_49977,N_49917);
or UO_1789 (O_1789,N_49961,N_49917);
nand UO_1790 (O_1790,N_49991,N_49915);
and UO_1791 (O_1791,N_49851,N_49815);
xnor UO_1792 (O_1792,N_49759,N_49800);
nand UO_1793 (O_1793,N_49932,N_49801);
nand UO_1794 (O_1794,N_49790,N_49951);
nor UO_1795 (O_1795,N_49834,N_49988);
and UO_1796 (O_1796,N_49764,N_49975);
nor UO_1797 (O_1797,N_49952,N_49795);
xor UO_1798 (O_1798,N_49804,N_49974);
or UO_1799 (O_1799,N_49940,N_49804);
or UO_1800 (O_1800,N_49939,N_49808);
nor UO_1801 (O_1801,N_49839,N_49787);
or UO_1802 (O_1802,N_49889,N_49966);
nand UO_1803 (O_1803,N_49903,N_49781);
and UO_1804 (O_1804,N_49768,N_49845);
nor UO_1805 (O_1805,N_49967,N_49775);
xor UO_1806 (O_1806,N_49813,N_49913);
xor UO_1807 (O_1807,N_49986,N_49814);
nor UO_1808 (O_1808,N_49850,N_49794);
nand UO_1809 (O_1809,N_49842,N_49857);
or UO_1810 (O_1810,N_49844,N_49828);
or UO_1811 (O_1811,N_49822,N_49782);
and UO_1812 (O_1812,N_49902,N_49971);
xor UO_1813 (O_1813,N_49825,N_49874);
and UO_1814 (O_1814,N_49974,N_49845);
nor UO_1815 (O_1815,N_49815,N_49754);
or UO_1816 (O_1816,N_49895,N_49933);
nor UO_1817 (O_1817,N_49882,N_49845);
or UO_1818 (O_1818,N_49930,N_49949);
nand UO_1819 (O_1819,N_49924,N_49858);
or UO_1820 (O_1820,N_49936,N_49769);
nor UO_1821 (O_1821,N_49914,N_49996);
xor UO_1822 (O_1822,N_49900,N_49925);
or UO_1823 (O_1823,N_49918,N_49813);
or UO_1824 (O_1824,N_49763,N_49760);
xor UO_1825 (O_1825,N_49939,N_49771);
and UO_1826 (O_1826,N_49864,N_49964);
nor UO_1827 (O_1827,N_49777,N_49831);
xnor UO_1828 (O_1828,N_49777,N_49962);
nand UO_1829 (O_1829,N_49888,N_49794);
xnor UO_1830 (O_1830,N_49845,N_49929);
nor UO_1831 (O_1831,N_49901,N_49907);
and UO_1832 (O_1832,N_49985,N_49972);
and UO_1833 (O_1833,N_49824,N_49939);
or UO_1834 (O_1834,N_49889,N_49828);
nor UO_1835 (O_1835,N_49985,N_49943);
nand UO_1836 (O_1836,N_49986,N_49933);
or UO_1837 (O_1837,N_49937,N_49769);
nand UO_1838 (O_1838,N_49859,N_49790);
xnor UO_1839 (O_1839,N_49926,N_49951);
nand UO_1840 (O_1840,N_49860,N_49815);
nor UO_1841 (O_1841,N_49852,N_49874);
xor UO_1842 (O_1842,N_49902,N_49822);
xor UO_1843 (O_1843,N_49873,N_49996);
nor UO_1844 (O_1844,N_49959,N_49878);
or UO_1845 (O_1845,N_49873,N_49949);
nor UO_1846 (O_1846,N_49864,N_49906);
nand UO_1847 (O_1847,N_49941,N_49871);
and UO_1848 (O_1848,N_49876,N_49869);
and UO_1849 (O_1849,N_49862,N_49968);
and UO_1850 (O_1850,N_49954,N_49961);
xnor UO_1851 (O_1851,N_49930,N_49836);
or UO_1852 (O_1852,N_49857,N_49837);
xnor UO_1853 (O_1853,N_49965,N_49938);
or UO_1854 (O_1854,N_49887,N_49853);
nand UO_1855 (O_1855,N_49981,N_49751);
or UO_1856 (O_1856,N_49905,N_49855);
or UO_1857 (O_1857,N_49902,N_49753);
nor UO_1858 (O_1858,N_49896,N_49986);
nand UO_1859 (O_1859,N_49893,N_49788);
nor UO_1860 (O_1860,N_49886,N_49779);
nor UO_1861 (O_1861,N_49877,N_49851);
nor UO_1862 (O_1862,N_49779,N_49860);
nor UO_1863 (O_1863,N_49819,N_49836);
nand UO_1864 (O_1864,N_49808,N_49945);
nor UO_1865 (O_1865,N_49825,N_49944);
nor UO_1866 (O_1866,N_49940,N_49946);
and UO_1867 (O_1867,N_49842,N_49847);
and UO_1868 (O_1868,N_49862,N_49934);
or UO_1869 (O_1869,N_49950,N_49886);
nor UO_1870 (O_1870,N_49987,N_49789);
xor UO_1871 (O_1871,N_49805,N_49901);
nor UO_1872 (O_1872,N_49835,N_49854);
nor UO_1873 (O_1873,N_49874,N_49812);
nor UO_1874 (O_1874,N_49979,N_49998);
and UO_1875 (O_1875,N_49855,N_49885);
or UO_1876 (O_1876,N_49858,N_49906);
or UO_1877 (O_1877,N_49943,N_49976);
nand UO_1878 (O_1878,N_49986,N_49927);
or UO_1879 (O_1879,N_49787,N_49830);
xnor UO_1880 (O_1880,N_49766,N_49945);
nor UO_1881 (O_1881,N_49984,N_49894);
and UO_1882 (O_1882,N_49843,N_49753);
and UO_1883 (O_1883,N_49938,N_49916);
or UO_1884 (O_1884,N_49866,N_49971);
nand UO_1885 (O_1885,N_49930,N_49882);
or UO_1886 (O_1886,N_49873,N_49952);
nor UO_1887 (O_1887,N_49818,N_49841);
or UO_1888 (O_1888,N_49837,N_49780);
xor UO_1889 (O_1889,N_49774,N_49926);
nand UO_1890 (O_1890,N_49760,N_49818);
nor UO_1891 (O_1891,N_49882,N_49869);
and UO_1892 (O_1892,N_49932,N_49922);
nand UO_1893 (O_1893,N_49970,N_49950);
nor UO_1894 (O_1894,N_49862,N_49986);
and UO_1895 (O_1895,N_49960,N_49807);
nor UO_1896 (O_1896,N_49884,N_49939);
xnor UO_1897 (O_1897,N_49771,N_49759);
nor UO_1898 (O_1898,N_49775,N_49790);
and UO_1899 (O_1899,N_49963,N_49888);
nor UO_1900 (O_1900,N_49882,N_49906);
xnor UO_1901 (O_1901,N_49858,N_49965);
xnor UO_1902 (O_1902,N_49809,N_49923);
nand UO_1903 (O_1903,N_49829,N_49838);
xor UO_1904 (O_1904,N_49886,N_49945);
or UO_1905 (O_1905,N_49787,N_49967);
xnor UO_1906 (O_1906,N_49837,N_49941);
and UO_1907 (O_1907,N_49758,N_49849);
nor UO_1908 (O_1908,N_49771,N_49754);
nor UO_1909 (O_1909,N_49922,N_49780);
nor UO_1910 (O_1910,N_49756,N_49993);
and UO_1911 (O_1911,N_49947,N_49825);
or UO_1912 (O_1912,N_49804,N_49874);
xor UO_1913 (O_1913,N_49916,N_49990);
and UO_1914 (O_1914,N_49998,N_49963);
or UO_1915 (O_1915,N_49830,N_49873);
nand UO_1916 (O_1916,N_49808,N_49941);
xnor UO_1917 (O_1917,N_49751,N_49937);
xor UO_1918 (O_1918,N_49960,N_49879);
or UO_1919 (O_1919,N_49932,N_49994);
or UO_1920 (O_1920,N_49949,N_49852);
nand UO_1921 (O_1921,N_49983,N_49978);
nand UO_1922 (O_1922,N_49930,N_49867);
and UO_1923 (O_1923,N_49880,N_49815);
nor UO_1924 (O_1924,N_49979,N_49828);
or UO_1925 (O_1925,N_49929,N_49986);
and UO_1926 (O_1926,N_49926,N_49960);
nor UO_1927 (O_1927,N_49888,N_49953);
nor UO_1928 (O_1928,N_49777,N_49878);
and UO_1929 (O_1929,N_49769,N_49814);
nor UO_1930 (O_1930,N_49986,N_49773);
nor UO_1931 (O_1931,N_49757,N_49946);
nand UO_1932 (O_1932,N_49854,N_49933);
xor UO_1933 (O_1933,N_49927,N_49850);
xnor UO_1934 (O_1934,N_49758,N_49803);
or UO_1935 (O_1935,N_49964,N_49787);
xor UO_1936 (O_1936,N_49891,N_49937);
nor UO_1937 (O_1937,N_49822,N_49766);
and UO_1938 (O_1938,N_49811,N_49878);
nand UO_1939 (O_1939,N_49861,N_49975);
and UO_1940 (O_1940,N_49894,N_49857);
and UO_1941 (O_1941,N_49911,N_49958);
or UO_1942 (O_1942,N_49866,N_49836);
and UO_1943 (O_1943,N_49939,N_49997);
and UO_1944 (O_1944,N_49956,N_49974);
and UO_1945 (O_1945,N_49925,N_49884);
nand UO_1946 (O_1946,N_49893,N_49829);
nand UO_1947 (O_1947,N_49885,N_49879);
and UO_1948 (O_1948,N_49755,N_49885);
and UO_1949 (O_1949,N_49963,N_49782);
or UO_1950 (O_1950,N_49910,N_49877);
nand UO_1951 (O_1951,N_49762,N_49989);
nand UO_1952 (O_1952,N_49766,N_49983);
and UO_1953 (O_1953,N_49813,N_49796);
nand UO_1954 (O_1954,N_49752,N_49841);
or UO_1955 (O_1955,N_49775,N_49764);
or UO_1956 (O_1956,N_49944,N_49924);
nor UO_1957 (O_1957,N_49779,N_49793);
nand UO_1958 (O_1958,N_49976,N_49798);
or UO_1959 (O_1959,N_49836,N_49987);
xor UO_1960 (O_1960,N_49854,N_49942);
xor UO_1961 (O_1961,N_49992,N_49970);
or UO_1962 (O_1962,N_49905,N_49771);
and UO_1963 (O_1963,N_49920,N_49802);
nor UO_1964 (O_1964,N_49764,N_49834);
and UO_1965 (O_1965,N_49830,N_49788);
xor UO_1966 (O_1966,N_49759,N_49810);
xnor UO_1967 (O_1967,N_49855,N_49925);
and UO_1968 (O_1968,N_49916,N_49822);
xor UO_1969 (O_1969,N_49833,N_49885);
nand UO_1970 (O_1970,N_49764,N_49790);
xor UO_1971 (O_1971,N_49831,N_49772);
or UO_1972 (O_1972,N_49923,N_49849);
and UO_1973 (O_1973,N_49839,N_49894);
and UO_1974 (O_1974,N_49924,N_49879);
nor UO_1975 (O_1975,N_49847,N_49858);
or UO_1976 (O_1976,N_49804,N_49814);
and UO_1977 (O_1977,N_49951,N_49986);
and UO_1978 (O_1978,N_49865,N_49769);
and UO_1979 (O_1979,N_49916,N_49960);
nand UO_1980 (O_1980,N_49755,N_49904);
or UO_1981 (O_1981,N_49754,N_49885);
nor UO_1982 (O_1982,N_49897,N_49931);
or UO_1983 (O_1983,N_49983,N_49970);
nand UO_1984 (O_1984,N_49773,N_49766);
or UO_1985 (O_1985,N_49864,N_49845);
xor UO_1986 (O_1986,N_49813,N_49764);
or UO_1987 (O_1987,N_49924,N_49960);
nor UO_1988 (O_1988,N_49934,N_49783);
nand UO_1989 (O_1989,N_49935,N_49922);
xor UO_1990 (O_1990,N_49829,N_49938);
xor UO_1991 (O_1991,N_49952,N_49972);
xor UO_1992 (O_1992,N_49882,N_49989);
or UO_1993 (O_1993,N_49998,N_49935);
nand UO_1994 (O_1994,N_49926,N_49866);
or UO_1995 (O_1995,N_49826,N_49780);
or UO_1996 (O_1996,N_49793,N_49968);
nand UO_1997 (O_1997,N_49955,N_49897);
nor UO_1998 (O_1998,N_49944,N_49834);
and UO_1999 (O_1999,N_49921,N_49953);
nor UO_2000 (O_2000,N_49821,N_49919);
xor UO_2001 (O_2001,N_49859,N_49911);
nand UO_2002 (O_2002,N_49814,N_49873);
and UO_2003 (O_2003,N_49996,N_49882);
nor UO_2004 (O_2004,N_49758,N_49896);
or UO_2005 (O_2005,N_49944,N_49804);
nor UO_2006 (O_2006,N_49896,N_49803);
and UO_2007 (O_2007,N_49872,N_49839);
nand UO_2008 (O_2008,N_49848,N_49878);
nand UO_2009 (O_2009,N_49938,N_49887);
or UO_2010 (O_2010,N_49882,N_49841);
or UO_2011 (O_2011,N_49859,N_49906);
xor UO_2012 (O_2012,N_49885,N_49842);
or UO_2013 (O_2013,N_49913,N_49925);
nand UO_2014 (O_2014,N_49783,N_49770);
and UO_2015 (O_2015,N_49897,N_49904);
xnor UO_2016 (O_2016,N_49958,N_49791);
nor UO_2017 (O_2017,N_49956,N_49750);
nand UO_2018 (O_2018,N_49988,N_49811);
xnor UO_2019 (O_2019,N_49792,N_49900);
nor UO_2020 (O_2020,N_49867,N_49852);
and UO_2021 (O_2021,N_49974,N_49935);
xnor UO_2022 (O_2022,N_49951,N_49991);
xnor UO_2023 (O_2023,N_49833,N_49923);
nand UO_2024 (O_2024,N_49760,N_49766);
or UO_2025 (O_2025,N_49972,N_49945);
nand UO_2026 (O_2026,N_49812,N_49844);
xnor UO_2027 (O_2027,N_49827,N_49880);
and UO_2028 (O_2028,N_49974,N_49963);
nor UO_2029 (O_2029,N_49886,N_49834);
and UO_2030 (O_2030,N_49771,N_49948);
xnor UO_2031 (O_2031,N_49863,N_49899);
nand UO_2032 (O_2032,N_49981,N_49996);
nor UO_2033 (O_2033,N_49916,N_49895);
and UO_2034 (O_2034,N_49836,N_49899);
nand UO_2035 (O_2035,N_49970,N_49957);
and UO_2036 (O_2036,N_49765,N_49759);
nor UO_2037 (O_2037,N_49814,N_49892);
or UO_2038 (O_2038,N_49808,N_49898);
nor UO_2039 (O_2039,N_49969,N_49859);
nand UO_2040 (O_2040,N_49986,N_49967);
or UO_2041 (O_2041,N_49931,N_49996);
nor UO_2042 (O_2042,N_49977,N_49866);
or UO_2043 (O_2043,N_49823,N_49964);
nand UO_2044 (O_2044,N_49867,N_49963);
nand UO_2045 (O_2045,N_49808,N_49999);
nor UO_2046 (O_2046,N_49884,N_49962);
nand UO_2047 (O_2047,N_49775,N_49975);
nor UO_2048 (O_2048,N_49820,N_49848);
and UO_2049 (O_2049,N_49756,N_49902);
and UO_2050 (O_2050,N_49972,N_49999);
xor UO_2051 (O_2051,N_49829,N_49800);
or UO_2052 (O_2052,N_49833,N_49889);
nand UO_2053 (O_2053,N_49976,N_49829);
nand UO_2054 (O_2054,N_49897,N_49917);
xnor UO_2055 (O_2055,N_49880,N_49938);
nor UO_2056 (O_2056,N_49868,N_49754);
or UO_2057 (O_2057,N_49792,N_49941);
and UO_2058 (O_2058,N_49846,N_49770);
and UO_2059 (O_2059,N_49762,N_49801);
or UO_2060 (O_2060,N_49897,N_49760);
xor UO_2061 (O_2061,N_49823,N_49814);
or UO_2062 (O_2062,N_49770,N_49920);
nor UO_2063 (O_2063,N_49941,N_49761);
or UO_2064 (O_2064,N_49848,N_49795);
and UO_2065 (O_2065,N_49914,N_49850);
and UO_2066 (O_2066,N_49835,N_49841);
xor UO_2067 (O_2067,N_49970,N_49842);
or UO_2068 (O_2068,N_49783,N_49872);
nand UO_2069 (O_2069,N_49942,N_49956);
or UO_2070 (O_2070,N_49988,N_49767);
nand UO_2071 (O_2071,N_49919,N_49918);
nor UO_2072 (O_2072,N_49795,N_49959);
xor UO_2073 (O_2073,N_49965,N_49903);
nor UO_2074 (O_2074,N_49899,N_49988);
or UO_2075 (O_2075,N_49765,N_49960);
nor UO_2076 (O_2076,N_49789,N_49922);
or UO_2077 (O_2077,N_49840,N_49975);
nand UO_2078 (O_2078,N_49903,N_49801);
xnor UO_2079 (O_2079,N_49958,N_49805);
nor UO_2080 (O_2080,N_49811,N_49887);
or UO_2081 (O_2081,N_49794,N_49861);
xnor UO_2082 (O_2082,N_49864,N_49935);
nand UO_2083 (O_2083,N_49787,N_49868);
nand UO_2084 (O_2084,N_49971,N_49949);
nand UO_2085 (O_2085,N_49807,N_49980);
xor UO_2086 (O_2086,N_49996,N_49778);
nand UO_2087 (O_2087,N_49898,N_49997);
nand UO_2088 (O_2088,N_49994,N_49875);
and UO_2089 (O_2089,N_49841,N_49874);
nor UO_2090 (O_2090,N_49825,N_49869);
xor UO_2091 (O_2091,N_49868,N_49839);
xor UO_2092 (O_2092,N_49808,N_49990);
nor UO_2093 (O_2093,N_49970,N_49966);
or UO_2094 (O_2094,N_49797,N_49812);
nand UO_2095 (O_2095,N_49955,N_49888);
xnor UO_2096 (O_2096,N_49815,N_49939);
and UO_2097 (O_2097,N_49901,N_49884);
or UO_2098 (O_2098,N_49839,N_49802);
and UO_2099 (O_2099,N_49785,N_49876);
nand UO_2100 (O_2100,N_49906,N_49784);
nor UO_2101 (O_2101,N_49850,N_49796);
or UO_2102 (O_2102,N_49909,N_49866);
and UO_2103 (O_2103,N_49847,N_49783);
and UO_2104 (O_2104,N_49948,N_49826);
or UO_2105 (O_2105,N_49930,N_49857);
nor UO_2106 (O_2106,N_49899,N_49834);
nand UO_2107 (O_2107,N_49906,N_49924);
and UO_2108 (O_2108,N_49861,N_49781);
xor UO_2109 (O_2109,N_49987,N_49810);
and UO_2110 (O_2110,N_49750,N_49993);
and UO_2111 (O_2111,N_49899,N_49997);
nand UO_2112 (O_2112,N_49942,N_49770);
or UO_2113 (O_2113,N_49795,N_49860);
nand UO_2114 (O_2114,N_49893,N_49775);
xnor UO_2115 (O_2115,N_49908,N_49876);
nand UO_2116 (O_2116,N_49776,N_49761);
xnor UO_2117 (O_2117,N_49949,N_49994);
and UO_2118 (O_2118,N_49755,N_49993);
or UO_2119 (O_2119,N_49794,N_49884);
nor UO_2120 (O_2120,N_49911,N_49780);
or UO_2121 (O_2121,N_49808,N_49915);
or UO_2122 (O_2122,N_49878,N_49960);
and UO_2123 (O_2123,N_49871,N_49978);
xnor UO_2124 (O_2124,N_49985,N_49988);
or UO_2125 (O_2125,N_49984,N_49848);
and UO_2126 (O_2126,N_49763,N_49821);
and UO_2127 (O_2127,N_49901,N_49780);
or UO_2128 (O_2128,N_49910,N_49907);
nand UO_2129 (O_2129,N_49960,N_49849);
nor UO_2130 (O_2130,N_49898,N_49980);
nor UO_2131 (O_2131,N_49758,N_49937);
or UO_2132 (O_2132,N_49983,N_49783);
nand UO_2133 (O_2133,N_49894,N_49775);
xnor UO_2134 (O_2134,N_49826,N_49911);
nor UO_2135 (O_2135,N_49989,N_49926);
nand UO_2136 (O_2136,N_49859,N_49931);
xor UO_2137 (O_2137,N_49862,N_49767);
and UO_2138 (O_2138,N_49758,N_49752);
xor UO_2139 (O_2139,N_49894,N_49763);
and UO_2140 (O_2140,N_49822,N_49783);
or UO_2141 (O_2141,N_49969,N_49847);
and UO_2142 (O_2142,N_49886,N_49853);
or UO_2143 (O_2143,N_49913,N_49803);
xor UO_2144 (O_2144,N_49865,N_49926);
or UO_2145 (O_2145,N_49964,N_49951);
xor UO_2146 (O_2146,N_49869,N_49906);
xor UO_2147 (O_2147,N_49875,N_49833);
xnor UO_2148 (O_2148,N_49820,N_49821);
or UO_2149 (O_2149,N_49894,N_49808);
nand UO_2150 (O_2150,N_49768,N_49779);
xor UO_2151 (O_2151,N_49991,N_49792);
or UO_2152 (O_2152,N_49760,N_49970);
or UO_2153 (O_2153,N_49930,N_49878);
nand UO_2154 (O_2154,N_49876,N_49983);
nor UO_2155 (O_2155,N_49980,N_49797);
or UO_2156 (O_2156,N_49971,N_49926);
nand UO_2157 (O_2157,N_49850,N_49763);
nor UO_2158 (O_2158,N_49994,N_49899);
or UO_2159 (O_2159,N_49995,N_49819);
nand UO_2160 (O_2160,N_49958,N_49777);
xnor UO_2161 (O_2161,N_49773,N_49951);
nand UO_2162 (O_2162,N_49947,N_49775);
or UO_2163 (O_2163,N_49975,N_49821);
and UO_2164 (O_2164,N_49925,N_49909);
nor UO_2165 (O_2165,N_49926,N_49823);
or UO_2166 (O_2166,N_49979,N_49902);
or UO_2167 (O_2167,N_49824,N_49960);
nor UO_2168 (O_2168,N_49778,N_49869);
and UO_2169 (O_2169,N_49827,N_49915);
xnor UO_2170 (O_2170,N_49979,N_49900);
and UO_2171 (O_2171,N_49797,N_49801);
and UO_2172 (O_2172,N_49816,N_49979);
or UO_2173 (O_2173,N_49790,N_49812);
nor UO_2174 (O_2174,N_49750,N_49788);
nor UO_2175 (O_2175,N_49910,N_49985);
nand UO_2176 (O_2176,N_49791,N_49892);
nor UO_2177 (O_2177,N_49893,N_49995);
or UO_2178 (O_2178,N_49811,N_49870);
or UO_2179 (O_2179,N_49779,N_49844);
or UO_2180 (O_2180,N_49879,N_49911);
or UO_2181 (O_2181,N_49848,N_49960);
and UO_2182 (O_2182,N_49762,N_49820);
and UO_2183 (O_2183,N_49917,N_49981);
nand UO_2184 (O_2184,N_49938,N_49996);
nand UO_2185 (O_2185,N_49880,N_49787);
and UO_2186 (O_2186,N_49929,N_49890);
nor UO_2187 (O_2187,N_49846,N_49917);
nand UO_2188 (O_2188,N_49752,N_49826);
and UO_2189 (O_2189,N_49871,N_49991);
xor UO_2190 (O_2190,N_49899,N_49797);
nand UO_2191 (O_2191,N_49921,N_49905);
nand UO_2192 (O_2192,N_49900,N_49955);
or UO_2193 (O_2193,N_49794,N_49763);
and UO_2194 (O_2194,N_49751,N_49957);
and UO_2195 (O_2195,N_49960,N_49794);
xor UO_2196 (O_2196,N_49762,N_49925);
nand UO_2197 (O_2197,N_49932,N_49975);
nand UO_2198 (O_2198,N_49970,N_49872);
xor UO_2199 (O_2199,N_49895,N_49795);
xor UO_2200 (O_2200,N_49763,N_49920);
or UO_2201 (O_2201,N_49783,N_49821);
or UO_2202 (O_2202,N_49912,N_49920);
and UO_2203 (O_2203,N_49878,N_49973);
nor UO_2204 (O_2204,N_49875,N_49786);
xnor UO_2205 (O_2205,N_49905,N_49839);
xnor UO_2206 (O_2206,N_49759,N_49988);
and UO_2207 (O_2207,N_49806,N_49974);
nor UO_2208 (O_2208,N_49873,N_49956);
or UO_2209 (O_2209,N_49972,N_49762);
xor UO_2210 (O_2210,N_49992,N_49964);
nor UO_2211 (O_2211,N_49862,N_49992);
nand UO_2212 (O_2212,N_49855,N_49973);
or UO_2213 (O_2213,N_49977,N_49859);
and UO_2214 (O_2214,N_49817,N_49903);
and UO_2215 (O_2215,N_49837,N_49800);
nand UO_2216 (O_2216,N_49981,N_49851);
and UO_2217 (O_2217,N_49909,N_49886);
xor UO_2218 (O_2218,N_49907,N_49769);
nor UO_2219 (O_2219,N_49884,N_49824);
and UO_2220 (O_2220,N_49974,N_49795);
and UO_2221 (O_2221,N_49826,N_49899);
nor UO_2222 (O_2222,N_49861,N_49987);
xnor UO_2223 (O_2223,N_49959,N_49750);
xor UO_2224 (O_2224,N_49838,N_49952);
nor UO_2225 (O_2225,N_49998,N_49975);
nand UO_2226 (O_2226,N_49754,N_49829);
nor UO_2227 (O_2227,N_49787,N_49900);
nand UO_2228 (O_2228,N_49876,N_49944);
xor UO_2229 (O_2229,N_49764,N_49962);
nand UO_2230 (O_2230,N_49940,N_49884);
and UO_2231 (O_2231,N_49959,N_49843);
nor UO_2232 (O_2232,N_49793,N_49809);
and UO_2233 (O_2233,N_49780,N_49766);
or UO_2234 (O_2234,N_49788,N_49822);
nand UO_2235 (O_2235,N_49826,N_49802);
and UO_2236 (O_2236,N_49814,N_49899);
xor UO_2237 (O_2237,N_49867,N_49857);
nor UO_2238 (O_2238,N_49989,N_49964);
xor UO_2239 (O_2239,N_49868,N_49867);
and UO_2240 (O_2240,N_49860,N_49817);
nor UO_2241 (O_2241,N_49773,N_49931);
and UO_2242 (O_2242,N_49874,N_49996);
nand UO_2243 (O_2243,N_49961,N_49984);
xnor UO_2244 (O_2244,N_49877,N_49784);
xnor UO_2245 (O_2245,N_49833,N_49921);
nand UO_2246 (O_2246,N_49901,N_49877);
or UO_2247 (O_2247,N_49764,N_49860);
and UO_2248 (O_2248,N_49850,N_49926);
xor UO_2249 (O_2249,N_49848,N_49858);
or UO_2250 (O_2250,N_49899,N_49808);
or UO_2251 (O_2251,N_49875,N_49922);
and UO_2252 (O_2252,N_49971,N_49878);
xnor UO_2253 (O_2253,N_49943,N_49915);
and UO_2254 (O_2254,N_49877,N_49985);
nand UO_2255 (O_2255,N_49824,N_49942);
or UO_2256 (O_2256,N_49895,N_49758);
and UO_2257 (O_2257,N_49920,N_49762);
or UO_2258 (O_2258,N_49981,N_49871);
nand UO_2259 (O_2259,N_49988,N_49770);
nand UO_2260 (O_2260,N_49896,N_49829);
nand UO_2261 (O_2261,N_49763,N_49880);
xnor UO_2262 (O_2262,N_49782,N_49946);
xor UO_2263 (O_2263,N_49816,N_49755);
nand UO_2264 (O_2264,N_49898,N_49761);
nor UO_2265 (O_2265,N_49890,N_49859);
or UO_2266 (O_2266,N_49823,N_49781);
or UO_2267 (O_2267,N_49773,N_49792);
nand UO_2268 (O_2268,N_49968,N_49864);
xnor UO_2269 (O_2269,N_49992,N_49979);
xnor UO_2270 (O_2270,N_49853,N_49803);
nor UO_2271 (O_2271,N_49871,N_49810);
nor UO_2272 (O_2272,N_49853,N_49906);
nor UO_2273 (O_2273,N_49959,N_49852);
or UO_2274 (O_2274,N_49906,N_49814);
xnor UO_2275 (O_2275,N_49890,N_49842);
nor UO_2276 (O_2276,N_49859,N_49958);
nor UO_2277 (O_2277,N_49970,N_49769);
nand UO_2278 (O_2278,N_49897,N_49977);
or UO_2279 (O_2279,N_49937,N_49967);
xor UO_2280 (O_2280,N_49976,N_49892);
nand UO_2281 (O_2281,N_49987,N_49869);
and UO_2282 (O_2282,N_49875,N_49847);
nand UO_2283 (O_2283,N_49957,N_49849);
xnor UO_2284 (O_2284,N_49769,N_49784);
nor UO_2285 (O_2285,N_49810,N_49932);
or UO_2286 (O_2286,N_49821,N_49930);
xnor UO_2287 (O_2287,N_49826,N_49996);
or UO_2288 (O_2288,N_49903,N_49882);
and UO_2289 (O_2289,N_49791,N_49827);
and UO_2290 (O_2290,N_49774,N_49799);
and UO_2291 (O_2291,N_49872,N_49851);
nor UO_2292 (O_2292,N_49801,N_49976);
xnor UO_2293 (O_2293,N_49864,N_49816);
nor UO_2294 (O_2294,N_49929,N_49808);
nor UO_2295 (O_2295,N_49984,N_49896);
and UO_2296 (O_2296,N_49920,N_49766);
xnor UO_2297 (O_2297,N_49914,N_49752);
xnor UO_2298 (O_2298,N_49857,N_49784);
and UO_2299 (O_2299,N_49823,N_49928);
xor UO_2300 (O_2300,N_49956,N_49998);
nand UO_2301 (O_2301,N_49868,N_49908);
xnor UO_2302 (O_2302,N_49857,N_49840);
or UO_2303 (O_2303,N_49832,N_49954);
nor UO_2304 (O_2304,N_49997,N_49942);
nor UO_2305 (O_2305,N_49843,N_49813);
nor UO_2306 (O_2306,N_49883,N_49937);
and UO_2307 (O_2307,N_49903,N_49779);
and UO_2308 (O_2308,N_49960,N_49768);
nand UO_2309 (O_2309,N_49828,N_49806);
xnor UO_2310 (O_2310,N_49755,N_49780);
xnor UO_2311 (O_2311,N_49806,N_49964);
or UO_2312 (O_2312,N_49786,N_49865);
nand UO_2313 (O_2313,N_49796,N_49894);
and UO_2314 (O_2314,N_49926,N_49849);
nand UO_2315 (O_2315,N_49761,N_49895);
xor UO_2316 (O_2316,N_49756,N_49773);
and UO_2317 (O_2317,N_49803,N_49937);
and UO_2318 (O_2318,N_49798,N_49905);
or UO_2319 (O_2319,N_49785,N_49794);
or UO_2320 (O_2320,N_49959,N_49765);
nor UO_2321 (O_2321,N_49893,N_49805);
nor UO_2322 (O_2322,N_49820,N_49892);
or UO_2323 (O_2323,N_49853,N_49907);
nor UO_2324 (O_2324,N_49759,N_49968);
xnor UO_2325 (O_2325,N_49752,N_49966);
nand UO_2326 (O_2326,N_49941,N_49810);
xor UO_2327 (O_2327,N_49830,N_49940);
xor UO_2328 (O_2328,N_49921,N_49892);
nand UO_2329 (O_2329,N_49924,N_49930);
or UO_2330 (O_2330,N_49837,N_49772);
nor UO_2331 (O_2331,N_49895,N_49811);
or UO_2332 (O_2332,N_49864,N_49811);
nor UO_2333 (O_2333,N_49870,N_49960);
nand UO_2334 (O_2334,N_49750,N_49818);
and UO_2335 (O_2335,N_49907,N_49776);
xor UO_2336 (O_2336,N_49777,N_49953);
nand UO_2337 (O_2337,N_49821,N_49937);
and UO_2338 (O_2338,N_49793,N_49761);
xor UO_2339 (O_2339,N_49823,N_49761);
nor UO_2340 (O_2340,N_49890,N_49754);
and UO_2341 (O_2341,N_49947,N_49801);
and UO_2342 (O_2342,N_49806,N_49779);
and UO_2343 (O_2343,N_49997,N_49750);
and UO_2344 (O_2344,N_49777,N_49944);
xnor UO_2345 (O_2345,N_49800,N_49824);
and UO_2346 (O_2346,N_49992,N_49886);
xnor UO_2347 (O_2347,N_49874,N_49894);
nand UO_2348 (O_2348,N_49828,N_49994);
or UO_2349 (O_2349,N_49915,N_49828);
or UO_2350 (O_2350,N_49785,N_49977);
and UO_2351 (O_2351,N_49948,N_49919);
and UO_2352 (O_2352,N_49939,N_49970);
and UO_2353 (O_2353,N_49848,N_49970);
nand UO_2354 (O_2354,N_49760,N_49921);
nor UO_2355 (O_2355,N_49785,N_49831);
xor UO_2356 (O_2356,N_49955,N_49824);
and UO_2357 (O_2357,N_49950,N_49802);
nand UO_2358 (O_2358,N_49939,N_49823);
nand UO_2359 (O_2359,N_49922,N_49860);
nor UO_2360 (O_2360,N_49835,N_49829);
or UO_2361 (O_2361,N_49893,N_49858);
or UO_2362 (O_2362,N_49920,N_49939);
or UO_2363 (O_2363,N_49847,N_49862);
nand UO_2364 (O_2364,N_49962,N_49822);
nand UO_2365 (O_2365,N_49781,N_49908);
xor UO_2366 (O_2366,N_49957,N_49999);
nand UO_2367 (O_2367,N_49765,N_49881);
nor UO_2368 (O_2368,N_49756,N_49973);
or UO_2369 (O_2369,N_49856,N_49857);
and UO_2370 (O_2370,N_49848,N_49824);
or UO_2371 (O_2371,N_49846,N_49835);
nor UO_2372 (O_2372,N_49926,N_49984);
and UO_2373 (O_2373,N_49777,N_49767);
nand UO_2374 (O_2374,N_49970,N_49800);
or UO_2375 (O_2375,N_49837,N_49820);
nor UO_2376 (O_2376,N_49931,N_49776);
xor UO_2377 (O_2377,N_49842,N_49881);
xor UO_2378 (O_2378,N_49866,N_49867);
nand UO_2379 (O_2379,N_49933,N_49960);
and UO_2380 (O_2380,N_49756,N_49801);
nor UO_2381 (O_2381,N_49925,N_49753);
and UO_2382 (O_2382,N_49770,N_49865);
or UO_2383 (O_2383,N_49811,N_49803);
and UO_2384 (O_2384,N_49794,N_49993);
xor UO_2385 (O_2385,N_49827,N_49916);
or UO_2386 (O_2386,N_49968,N_49897);
and UO_2387 (O_2387,N_49991,N_49837);
or UO_2388 (O_2388,N_49973,N_49943);
xor UO_2389 (O_2389,N_49996,N_49847);
and UO_2390 (O_2390,N_49799,N_49950);
xnor UO_2391 (O_2391,N_49766,N_49776);
or UO_2392 (O_2392,N_49776,N_49997);
or UO_2393 (O_2393,N_49810,N_49908);
or UO_2394 (O_2394,N_49909,N_49806);
nand UO_2395 (O_2395,N_49762,N_49917);
nor UO_2396 (O_2396,N_49860,N_49820);
and UO_2397 (O_2397,N_49904,N_49930);
or UO_2398 (O_2398,N_49831,N_49834);
or UO_2399 (O_2399,N_49926,N_49977);
xor UO_2400 (O_2400,N_49905,N_49755);
xnor UO_2401 (O_2401,N_49886,N_49822);
nand UO_2402 (O_2402,N_49868,N_49804);
xnor UO_2403 (O_2403,N_49962,N_49826);
xnor UO_2404 (O_2404,N_49873,N_49860);
or UO_2405 (O_2405,N_49844,N_49952);
xor UO_2406 (O_2406,N_49858,N_49930);
nand UO_2407 (O_2407,N_49977,N_49881);
nor UO_2408 (O_2408,N_49846,N_49910);
xor UO_2409 (O_2409,N_49885,N_49979);
and UO_2410 (O_2410,N_49819,N_49764);
xnor UO_2411 (O_2411,N_49756,N_49751);
nand UO_2412 (O_2412,N_49786,N_49900);
and UO_2413 (O_2413,N_49862,N_49955);
nand UO_2414 (O_2414,N_49967,N_49882);
xor UO_2415 (O_2415,N_49925,N_49885);
and UO_2416 (O_2416,N_49930,N_49838);
nand UO_2417 (O_2417,N_49828,N_49954);
nand UO_2418 (O_2418,N_49967,N_49828);
and UO_2419 (O_2419,N_49960,N_49755);
nand UO_2420 (O_2420,N_49840,N_49806);
or UO_2421 (O_2421,N_49813,N_49957);
nand UO_2422 (O_2422,N_49985,N_49848);
xor UO_2423 (O_2423,N_49950,N_49855);
or UO_2424 (O_2424,N_49795,N_49993);
or UO_2425 (O_2425,N_49772,N_49926);
and UO_2426 (O_2426,N_49861,N_49819);
xor UO_2427 (O_2427,N_49837,N_49920);
and UO_2428 (O_2428,N_49782,N_49987);
nor UO_2429 (O_2429,N_49853,N_49938);
xor UO_2430 (O_2430,N_49888,N_49864);
xnor UO_2431 (O_2431,N_49778,N_49799);
nor UO_2432 (O_2432,N_49987,N_49882);
xor UO_2433 (O_2433,N_49845,N_49885);
nor UO_2434 (O_2434,N_49846,N_49812);
nand UO_2435 (O_2435,N_49996,N_49853);
and UO_2436 (O_2436,N_49912,N_49933);
xnor UO_2437 (O_2437,N_49870,N_49894);
xor UO_2438 (O_2438,N_49790,N_49887);
or UO_2439 (O_2439,N_49894,N_49968);
xnor UO_2440 (O_2440,N_49785,N_49868);
xnor UO_2441 (O_2441,N_49995,N_49935);
xor UO_2442 (O_2442,N_49848,N_49996);
nand UO_2443 (O_2443,N_49892,N_49975);
or UO_2444 (O_2444,N_49953,N_49931);
nor UO_2445 (O_2445,N_49952,N_49775);
xnor UO_2446 (O_2446,N_49915,N_49982);
nand UO_2447 (O_2447,N_49966,N_49856);
xor UO_2448 (O_2448,N_49939,N_49886);
nor UO_2449 (O_2449,N_49759,N_49951);
nand UO_2450 (O_2450,N_49900,N_49902);
and UO_2451 (O_2451,N_49797,N_49946);
xnor UO_2452 (O_2452,N_49863,N_49914);
and UO_2453 (O_2453,N_49765,N_49862);
or UO_2454 (O_2454,N_49763,N_49840);
xor UO_2455 (O_2455,N_49761,N_49821);
nand UO_2456 (O_2456,N_49795,N_49940);
nand UO_2457 (O_2457,N_49975,N_49976);
and UO_2458 (O_2458,N_49754,N_49767);
nor UO_2459 (O_2459,N_49990,N_49943);
xor UO_2460 (O_2460,N_49913,N_49954);
nand UO_2461 (O_2461,N_49933,N_49798);
and UO_2462 (O_2462,N_49939,N_49954);
and UO_2463 (O_2463,N_49857,N_49887);
xnor UO_2464 (O_2464,N_49921,N_49924);
or UO_2465 (O_2465,N_49846,N_49822);
xor UO_2466 (O_2466,N_49897,N_49841);
nor UO_2467 (O_2467,N_49987,N_49780);
nor UO_2468 (O_2468,N_49933,N_49773);
xor UO_2469 (O_2469,N_49784,N_49796);
nor UO_2470 (O_2470,N_49848,N_49811);
nand UO_2471 (O_2471,N_49860,N_49834);
nor UO_2472 (O_2472,N_49792,N_49983);
or UO_2473 (O_2473,N_49799,N_49966);
nor UO_2474 (O_2474,N_49988,N_49880);
xnor UO_2475 (O_2475,N_49924,N_49925);
xor UO_2476 (O_2476,N_49868,N_49801);
and UO_2477 (O_2477,N_49783,N_49883);
xor UO_2478 (O_2478,N_49881,N_49887);
nor UO_2479 (O_2479,N_49750,N_49806);
xor UO_2480 (O_2480,N_49813,N_49854);
nand UO_2481 (O_2481,N_49864,N_49809);
and UO_2482 (O_2482,N_49779,N_49833);
nand UO_2483 (O_2483,N_49987,N_49866);
and UO_2484 (O_2484,N_49879,N_49781);
nand UO_2485 (O_2485,N_49791,N_49753);
or UO_2486 (O_2486,N_49829,N_49949);
xnor UO_2487 (O_2487,N_49855,N_49886);
or UO_2488 (O_2488,N_49964,N_49894);
nand UO_2489 (O_2489,N_49889,N_49992);
and UO_2490 (O_2490,N_49830,N_49972);
nand UO_2491 (O_2491,N_49991,N_49830);
xor UO_2492 (O_2492,N_49952,N_49924);
nand UO_2493 (O_2493,N_49954,N_49983);
or UO_2494 (O_2494,N_49995,N_49850);
xnor UO_2495 (O_2495,N_49844,N_49876);
nor UO_2496 (O_2496,N_49862,N_49874);
and UO_2497 (O_2497,N_49767,N_49752);
nor UO_2498 (O_2498,N_49834,N_49924);
and UO_2499 (O_2499,N_49986,N_49796);
and UO_2500 (O_2500,N_49859,N_49905);
or UO_2501 (O_2501,N_49910,N_49929);
nor UO_2502 (O_2502,N_49835,N_49928);
xor UO_2503 (O_2503,N_49921,N_49910);
or UO_2504 (O_2504,N_49761,N_49867);
or UO_2505 (O_2505,N_49966,N_49800);
nand UO_2506 (O_2506,N_49977,N_49874);
nor UO_2507 (O_2507,N_49914,N_49839);
nor UO_2508 (O_2508,N_49774,N_49958);
xnor UO_2509 (O_2509,N_49842,N_49793);
nand UO_2510 (O_2510,N_49781,N_49933);
nor UO_2511 (O_2511,N_49834,N_49947);
xor UO_2512 (O_2512,N_49890,N_49889);
and UO_2513 (O_2513,N_49869,N_49881);
and UO_2514 (O_2514,N_49804,N_49992);
and UO_2515 (O_2515,N_49812,N_49850);
and UO_2516 (O_2516,N_49807,N_49887);
or UO_2517 (O_2517,N_49825,N_49880);
and UO_2518 (O_2518,N_49797,N_49850);
nor UO_2519 (O_2519,N_49954,N_49856);
or UO_2520 (O_2520,N_49976,N_49820);
and UO_2521 (O_2521,N_49895,N_49847);
nor UO_2522 (O_2522,N_49914,N_49925);
xnor UO_2523 (O_2523,N_49779,N_49778);
nand UO_2524 (O_2524,N_49878,N_49993);
nand UO_2525 (O_2525,N_49903,N_49885);
or UO_2526 (O_2526,N_49765,N_49784);
nor UO_2527 (O_2527,N_49863,N_49778);
xor UO_2528 (O_2528,N_49815,N_49772);
and UO_2529 (O_2529,N_49810,N_49828);
nand UO_2530 (O_2530,N_49798,N_49938);
nor UO_2531 (O_2531,N_49982,N_49764);
nor UO_2532 (O_2532,N_49859,N_49998);
nor UO_2533 (O_2533,N_49833,N_49956);
nand UO_2534 (O_2534,N_49975,N_49786);
or UO_2535 (O_2535,N_49906,N_49804);
and UO_2536 (O_2536,N_49773,N_49784);
or UO_2537 (O_2537,N_49971,N_49957);
nor UO_2538 (O_2538,N_49868,N_49915);
nor UO_2539 (O_2539,N_49792,N_49920);
nand UO_2540 (O_2540,N_49934,N_49806);
or UO_2541 (O_2541,N_49866,N_49826);
and UO_2542 (O_2542,N_49943,N_49933);
nor UO_2543 (O_2543,N_49858,N_49958);
nor UO_2544 (O_2544,N_49850,N_49947);
nor UO_2545 (O_2545,N_49883,N_49852);
xnor UO_2546 (O_2546,N_49990,N_49962);
and UO_2547 (O_2547,N_49909,N_49762);
or UO_2548 (O_2548,N_49802,N_49909);
nand UO_2549 (O_2549,N_49966,N_49943);
xnor UO_2550 (O_2550,N_49995,N_49752);
nor UO_2551 (O_2551,N_49794,N_49898);
or UO_2552 (O_2552,N_49958,N_49944);
xor UO_2553 (O_2553,N_49772,N_49812);
xnor UO_2554 (O_2554,N_49779,N_49788);
xor UO_2555 (O_2555,N_49775,N_49911);
xor UO_2556 (O_2556,N_49784,N_49851);
xor UO_2557 (O_2557,N_49841,N_49986);
nand UO_2558 (O_2558,N_49915,N_49831);
and UO_2559 (O_2559,N_49927,N_49776);
or UO_2560 (O_2560,N_49986,N_49884);
and UO_2561 (O_2561,N_49915,N_49939);
nor UO_2562 (O_2562,N_49961,N_49910);
nand UO_2563 (O_2563,N_49777,N_49812);
nand UO_2564 (O_2564,N_49834,N_49993);
or UO_2565 (O_2565,N_49959,N_49803);
xor UO_2566 (O_2566,N_49927,N_49819);
xnor UO_2567 (O_2567,N_49761,N_49861);
nand UO_2568 (O_2568,N_49828,N_49874);
nor UO_2569 (O_2569,N_49767,N_49804);
and UO_2570 (O_2570,N_49992,N_49932);
nand UO_2571 (O_2571,N_49815,N_49916);
and UO_2572 (O_2572,N_49945,N_49976);
nand UO_2573 (O_2573,N_49832,N_49817);
or UO_2574 (O_2574,N_49867,N_49752);
xnor UO_2575 (O_2575,N_49895,N_49991);
and UO_2576 (O_2576,N_49980,N_49772);
and UO_2577 (O_2577,N_49926,N_49869);
xnor UO_2578 (O_2578,N_49884,N_49823);
nor UO_2579 (O_2579,N_49863,N_49989);
and UO_2580 (O_2580,N_49887,N_49956);
nor UO_2581 (O_2581,N_49934,N_49914);
and UO_2582 (O_2582,N_49843,N_49791);
and UO_2583 (O_2583,N_49817,N_49844);
and UO_2584 (O_2584,N_49887,N_49886);
xnor UO_2585 (O_2585,N_49921,N_49793);
or UO_2586 (O_2586,N_49767,N_49909);
or UO_2587 (O_2587,N_49830,N_49796);
nor UO_2588 (O_2588,N_49924,N_49843);
xnor UO_2589 (O_2589,N_49893,N_49819);
nand UO_2590 (O_2590,N_49767,N_49808);
and UO_2591 (O_2591,N_49767,N_49817);
and UO_2592 (O_2592,N_49949,N_49945);
nor UO_2593 (O_2593,N_49927,N_49787);
and UO_2594 (O_2594,N_49911,N_49908);
nand UO_2595 (O_2595,N_49922,N_49929);
nand UO_2596 (O_2596,N_49815,N_49881);
or UO_2597 (O_2597,N_49992,N_49819);
and UO_2598 (O_2598,N_49899,N_49916);
xor UO_2599 (O_2599,N_49986,N_49790);
or UO_2600 (O_2600,N_49998,N_49831);
xnor UO_2601 (O_2601,N_49806,N_49939);
xor UO_2602 (O_2602,N_49837,N_49830);
nor UO_2603 (O_2603,N_49853,N_49814);
nor UO_2604 (O_2604,N_49759,N_49887);
or UO_2605 (O_2605,N_49966,N_49905);
nor UO_2606 (O_2606,N_49791,N_49802);
nand UO_2607 (O_2607,N_49857,N_49820);
nor UO_2608 (O_2608,N_49958,N_49809);
xor UO_2609 (O_2609,N_49929,N_49953);
or UO_2610 (O_2610,N_49849,N_49969);
nor UO_2611 (O_2611,N_49871,N_49853);
and UO_2612 (O_2612,N_49936,N_49791);
nor UO_2613 (O_2613,N_49862,N_49991);
nand UO_2614 (O_2614,N_49798,N_49980);
nor UO_2615 (O_2615,N_49879,N_49941);
xor UO_2616 (O_2616,N_49807,N_49826);
xor UO_2617 (O_2617,N_49945,N_49846);
or UO_2618 (O_2618,N_49880,N_49973);
or UO_2619 (O_2619,N_49772,N_49996);
xor UO_2620 (O_2620,N_49822,N_49913);
xnor UO_2621 (O_2621,N_49957,N_49973);
nor UO_2622 (O_2622,N_49793,N_49892);
and UO_2623 (O_2623,N_49806,N_49778);
xnor UO_2624 (O_2624,N_49761,N_49870);
and UO_2625 (O_2625,N_49973,N_49932);
nor UO_2626 (O_2626,N_49891,N_49797);
and UO_2627 (O_2627,N_49841,N_49994);
or UO_2628 (O_2628,N_49959,N_49927);
and UO_2629 (O_2629,N_49879,N_49909);
nand UO_2630 (O_2630,N_49837,N_49822);
and UO_2631 (O_2631,N_49914,N_49842);
xnor UO_2632 (O_2632,N_49918,N_49985);
nor UO_2633 (O_2633,N_49752,N_49897);
or UO_2634 (O_2634,N_49791,N_49792);
xnor UO_2635 (O_2635,N_49974,N_49936);
nor UO_2636 (O_2636,N_49837,N_49926);
nand UO_2637 (O_2637,N_49878,N_49797);
and UO_2638 (O_2638,N_49968,N_49853);
or UO_2639 (O_2639,N_49965,N_49988);
and UO_2640 (O_2640,N_49837,N_49841);
and UO_2641 (O_2641,N_49858,N_49758);
and UO_2642 (O_2642,N_49790,N_49841);
and UO_2643 (O_2643,N_49795,N_49924);
and UO_2644 (O_2644,N_49764,N_49761);
nor UO_2645 (O_2645,N_49880,N_49891);
and UO_2646 (O_2646,N_49891,N_49874);
nor UO_2647 (O_2647,N_49967,N_49795);
and UO_2648 (O_2648,N_49895,N_49938);
or UO_2649 (O_2649,N_49816,N_49939);
nor UO_2650 (O_2650,N_49992,N_49980);
and UO_2651 (O_2651,N_49769,N_49863);
or UO_2652 (O_2652,N_49814,N_49771);
and UO_2653 (O_2653,N_49786,N_49760);
nor UO_2654 (O_2654,N_49946,N_49807);
xnor UO_2655 (O_2655,N_49904,N_49923);
nand UO_2656 (O_2656,N_49771,N_49909);
xor UO_2657 (O_2657,N_49778,N_49922);
or UO_2658 (O_2658,N_49793,N_49967);
xor UO_2659 (O_2659,N_49792,N_49839);
nor UO_2660 (O_2660,N_49759,N_49954);
xnor UO_2661 (O_2661,N_49901,N_49973);
nor UO_2662 (O_2662,N_49929,N_49802);
and UO_2663 (O_2663,N_49774,N_49991);
nor UO_2664 (O_2664,N_49751,N_49917);
or UO_2665 (O_2665,N_49795,N_49760);
xor UO_2666 (O_2666,N_49975,N_49850);
xnor UO_2667 (O_2667,N_49774,N_49808);
or UO_2668 (O_2668,N_49767,N_49973);
or UO_2669 (O_2669,N_49936,N_49855);
nand UO_2670 (O_2670,N_49956,N_49761);
nor UO_2671 (O_2671,N_49817,N_49873);
nand UO_2672 (O_2672,N_49929,N_49899);
and UO_2673 (O_2673,N_49920,N_49822);
nand UO_2674 (O_2674,N_49921,N_49918);
nand UO_2675 (O_2675,N_49851,N_49819);
nor UO_2676 (O_2676,N_49842,N_49792);
nor UO_2677 (O_2677,N_49862,N_49914);
nand UO_2678 (O_2678,N_49993,N_49902);
nand UO_2679 (O_2679,N_49859,N_49897);
and UO_2680 (O_2680,N_49922,N_49930);
nand UO_2681 (O_2681,N_49998,N_49948);
and UO_2682 (O_2682,N_49856,N_49753);
xnor UO_2683 (O_2683,N_49816,N_49947);
nand UO_2684 (O_2684,N_49797,N_49773);
nor UO_2685 (O_2685,N_49828,N_49895);
xnor UO_2686 (O_2686,N_49858,N_49792);
nand UO_2687 (O_2687,N_49996,N_49813);
nor UO_2688 (O_2688,N_49765,N_49867);
nor UO_2689 (O_2689,N_49977,N_49752);
and UO_2690 (O_2690,N_49790,N_49852);
xnor UO_2691 (O_2691,N_49928,N_49995);
and UO_2692 (O_2692,N_49923,N_49952);
or UO_2693 (O_2693,N_49869,N_49971);
nor UO_2694 (O_2694,N_49893,N_49915);
and UO_2695 (O_2695,N_49972,N_49765);
xnor UO_2696 (O_2696,N_49805,N_49944);
and UO_2697 (O_2697,N_49903,N_49956);
and UO_2698 (O_2698,N_49905,N_49849);
and UO_2699 (O_2699,N_49930,N_49946);
xor UO_2700 (O_2700,N_49784,N_49787);
nor UO_2701 (O_2701,N_49833,N_49995);
or UO_2702 (O_2702,N_49916,N_49820);
or UO_2703 (O_2703,N_49757,N_49921);
nand UO_2704 (O_2704,N_49882,N_49977);
xnor UO_2705 (O_2705,N_49870,N_49760);
nand UO_2706 (O_2706,N_49810,N_49856);
xor UO_2707 (O_2707,N_49966,N_49842);
xnor UO_2708 (O_2708,N_49792,N_49778);
xnor UO_2709 (O_2709,N_49965,N_49780);
and UO_2710 (O_2710,N_49968,N_49851);
xnor UO_2711 (O_2711,N_49859,N_49807);
nor UO_2712 (O_2712,N_49914,N_49834);
and UO_2713 (O_2713,N_49873,N_49780);
nand UO_2714 (O_2714,N_49908,N_49838);
nand UO_2715 (O_2715,N_49872,N_49958);
nand UO_2716 (O_2716,N_49992,N_49753);
nor UO_2717 (O_2717,N_49918,N_49774);
or UO_2718 (O_2718,N_49893,N_49822);
xnor UO_2719 (O_2719,N_49945,N_49851);
xnor UO_2720 (O_2720,N_49787,N_49827);
and UO_2721 (O_2721,N_49856,N_49874);
xnor UO_2722 (O_2722,N_49889,N_49814);
nand UO_2723 (O_2723,N_49802,N_49884);
nor UO_2724 (O_2724,N_49802,N_49984);
or UO_2725 (O_2725,N_49827,N_49797);
or UO_2726 (O_2726,N_49912,N_49774);
or UO_2727 (O_2727,N_49753,N_49784);
xor UO_2728 (O_2728,N_49937,N_49807);
nand UO_2729 (O_2729,N_49912,N_49823);
and UO_2730 (O_2730,N_49795,N_49884);
and UO_2731 (O_2731,N_49840,N_49891);
and UO_2732 (O_2732,N_49752,N_49956);
xnor UO_2733 (O_2733,N_49874,N_49913);
nand UO_2734 (O_2734,N_49933,N_49761);
nand UO_2735 (O_2735,N_49770,N_49956);
and UO_2736 (O_2736,N_49834,N_49850);
and UO_2737 (O_2737,N_49971,N_49803);
nand UO_2738 (O_2738,N_49852,N_49903);
and UO_2739 (O_2739,N_49878,N_49939);
nand UO_2740 (O_2740,N_49923,N_49943);
nor UO_2741 (O_2741,N_49896,N_49880);
nand UO_2742 (O_2742,N_49910,N_49867);
or UO_2743 (O_2743,N_49887,N_49993);
and UO_2744 (O_2744,N_49775,N_49777);
xnor UO_2745 (O_2745,N_49750,N_49751);
or UO_2746 (O_2746,N_49977,N_49922);
or UO_2747 (O_2747,N_49902,N_49847);
xnor UO_2748 (O_2748,N_49766,N_49890);
xor UO_2749 (O_2749,N_49910,N_49922);
nor UO_2750 (O_2750,N_49810,N_49872);
or UO_2751 (O_2751,N_49952,N_49888);
nand UO_2752 (O_2752,N_49948,N_49869);
and UO_2753 (O_2753,N_49757,N_49859);
xor UO_2754 (O_2754,N_49889,N_49838);
nor UO_2755 (O_2755,N_49970,N_49771);
nand UO_2756 (O_2756,N_49803,N_49849);
and UO_2757 (O_2757,N_49902,N_49918);
or UO_2758 (O_2758,N_49887,N_49948);
and UO_2759 (O_2759,N_49803,N_49864);
nand UO_2760 (O_2760,N_49791,N_49815);
nor UO_2761 (O_2761,N_49902,N_49754);
xnor UO_2762 (O_2762,N_49871,N_49787);
xnor UO_2763 (O_2763,N_49963,N_49981);
nand UO_2764 (O_2764,N_49763,N_49826);
or UO_2765 (O_2765,N_49909,N_49847);
or UO_2766 (O_2766,N_49972,N_49836);
or UO_2767 (O_2767,N_49904,N_49883);
nand UO_2768 (O_2768,N_49976,N_49778);
xnor UO_2769 (O_2769,N_49882,N_49919);
nand UO_2770 (O_2770,N_49949,N_49996);
nor UO_2771 (O_2771,N_49891,N_49931);
or UO_2772 (O_2772,N_49940,N_49814);
nand UO_2773 (O_2773,N_49797,N_49772);
nor UO_2774 (O_2774,N_49766,N_49948);
or UO_2775 (O_2775,N_49893,N_49968);
nand UO_2776 (O_2776,N_49931,N_49849);
nor UO_2777 (O_2777,N_49857,N_49923);
or UO_2778 (O_2778,N_49818,N_49918);
nor UO_2779 (O_2779,N_49942,N_49955);
and UO_2780 (O_2780,N_49963,N_49886);
xnor UO_2781 (O_2781,N_49954,N_49982);
and UO_2782 (O_2782,N_49949,N_49856);
and UO_2783 (O_2783,N_49835,N_49812);
and UO_2784 (O_2784,N_49984,N_49982);
nor UO_2785 (O_2785,N_49920,N_49932);
or UO_2786 (O_2786,N_49811,N_49757);
and UO_2787 (O_2787,N_49758,N_49885);
nor UO_2788 (O_2788,N_49987,N_49984);
or UO_2789 (O_2789,N_49914,N_49888);
xnor UO_2790 (O_2790,N_49843,N_49897);
nor UO_2791 (O_2791,N_49944,N_49995);
nor UO_2792 (O_2792,N_49810,N_49950);
xor UO_2793 (O_2793,N_49819,N_49870);
or UO_2794 (O_2794,N_49843,N_49879);
nor UO_2795 (O_2795,N_49916,N_49888);
nor UO_2796 (O_2796,N_49835,N_49905);
xnor UO_2797 (O_2797,N_49786,N_49983);
xor UO_2798 (O_2798,N_49837,N_49765);
xor UO_2799 (O_2799,N_49893,N_49921);
or UO_2800 (O_2800,N_49829,N_49868);
and UO_2801 (O_2801,N_49964,N_49832);
nand UO_2802 (O_2802,N_49980,N_49908);
or UO_2803 (O_2803,N_49821,N_49780);
or UO_2804 (O_2804,N_49771,N_49772);
xor UO_2805 (O_2805,N_49815,N_49979);
or UO_2806 (O_2806,N_49898,N_49854);
xnor UO_2807 (O_2807,N_49824,N_49873);
nand UO_2808 (O_2808,N_49965,N_49846);
and UO_2809 (O_2809,N_49807,N_49875);
or UO_2810 (O_2810,N_49786,N_49906);
xnor UO_2811 (O_2811,N_49765,N_49830);
nor UO_2812 (O_2812,N_49916,N_49963);
nand UO_2813 (O_2813,N_49918,N_49987);
xor UO_2814 (O_2814,N_49816,N_49886);
and UO_2815 (O_2815,N_49885,N_49866);
or UO_2816 (O_2816,N_49882,N_49859);
and UO_2817 (O_2817,N_49797,N_49986);
and UO_2818 (O_2818,N_49961,N_49893);
nor UO_2819 (O_2819,N_49832,N_49942);
xor UO_2820 (O_2820,N_49789,N_49998);
xor UO_2821 (O_2821,N_49750,N_49922);
and UO_2822 (O_2822,N_49908,N_49999);
nand UO_2823 (O_2823,N_49810,N_49843);
nand UO_2824 (O_2824,N_49992,N_49923);
xor UO_2825 (O_2825,N_49882,N_49945);
xnor UO_2826 (O_2826,N_49797,N_49988);
xor UO_2827 (O_2827,N_49797,N_49884);
nor UO_2828 (O_2828,N_49988,N_49850);
xnor UO_2829 (O_2829,N_49788,N_49978);
nand UO_2830 (O_2830,N_49844,N_49910);
nor UO_2831 (O_2831,N_49792,N_49975);
nor UO_2832 (O_2832,N_49880,N_49981);
nand UO_2833 (O_2833,N_49857,N_49824);
or UO_2834 (O_2834,N_49976,N_49862);
nand UO_2835 (O_2835,N_49811,N_49918);
xor UO_2836 (O_2836,N_49893,N_49841);
and UO_2837 (O_2837,N_49945,N_49930);
xor UO_2838 (O_2838,N_49770,N_49929);
nor UO_2839 (O_2839,N_49954,N_49857);
and UO_2840 (O_2840,N_49911,N_49887);
or UO_2841 (O_2841,N_49819,N_49929);
or UO_2842 (O_2842,N_49991,N_49958);
and UO_2843 (O_2843,N_49859,N_49819);
xnor UO_2844 (O_2844,N_49779,N_49976);
and UO_2845 (O_2845,N_49785,N_49793);
or UO_2846 (O_2846,N_49999,N_49829);
nor UO_2847 (O_2847,N_49847,N_49944);
nand UO_2848 (O_2848,N_49894,N_49970);
and UO_2849 (O_2849,N_49848,N_49888);
xor UO_2850 (O_2850,N_49842,N_49925);
nand UO_2851 (O_2851,N_49897,N_49781);
nand UO_2852 (O_2852,N_49758,N_49756);
or UO_2853 (O_2853,N_49804,N_49975);
or UO_2854 (O_2854,N_49923,N_49838);
nor UO_2855 (O_2855,N_49986,N_49995);
xor UO_2856 (O_2856,N_49870,N_49754);
nor UO_2857 (O_2857,N_49820,N_49815);
nor UO_2858 (O_2858,N_49950,N_49767);
and UO_2859 (O_2859,N_49777,N_49935);
or UO_2860 (O_2860,N_49820,N_49949);
or UO_2861 (O_2861,N_49800,N_49994);
and UO_2862 (O_2862,N_49992,N_49828);
xor UO_2863 (O_2863,N_49971,N_49764);
nor UO_2864 (O_2864,N_49833,N_49790);
nor UO_2865 (O_2865,N_49836,N_49822);
or UO_2866 (O_2866,N_49783,N_49908);
nor UO_2867 (O_2867,N_49826,N_49843);
nor UO_2868 (O_2868,N_49761,N_49842);
nor UO_2869 (O_2869,N_49848,N_49932);
xnor UO_2870 (O_2870,N_49831,N_49775);
and UO_2871 (O_2871,N_49945,N_49794);
nand UO_2872 (O_2872,N_49853,N_49916);
and UO_2873 (O_2873,N_49793,N_49817);
and UO_2874 (O_2874,N_49967,N_49883);
and UO_2875 (O_2875,N_49931,N_49905);
or UO_2876 (O_2876,N_49915,N_49978);
and UO_2877 (O_2877,N_49845,N_49927);
nand UO_2878 (O_2878,N_49815,N_49830);
and UO_2879 (O_2879,N_49753,N_49884);
nand UO_2880 (O_2880,N_49938,N_49983);
or UO_2881 (O_2881,N_49889,N_49986);
xnor UO_2882 (O_2882,N_49931,N_49758);
xor UO_2883 (O_2883,N_49883,N_49918);
and UO_2884 (O_2884,N_49833,N_49837);
or UO_2885 (O_2885,N_49757,N_49965);
xnor UO_2886 (O_2886,N_49789,N_49841);
and UO_2887 (O_2887,N_49855,N_49759);
nand UO_2888 (O_2888,N_49914,N_49906);
and UO_2889 (O_2889,N_49871,N_49976);
or UO_2890 (O_2890,N_49963,N_49752);
nand UO_2891 (O_2891,N_49898,N_49818);
nand UO_2892 (O_2892,N_49912,N_49956);
nand UO_2893 (O_2893,N_49892,N_49788);
or UO_2894 (O_2894,N_49786,N_49851);
xnor UO_2895 (O_2895,N_49946,N_49771);
nor UO_2896 (O_2896,N_49965,N_49754);
xor UO_2897 (O_2897,N_49983,N_49859);
nor UO_2898 (O_2898,N_49867,N_49794);
and UO_2899 (O_2899,N_49884,N_49826);
nand UO_2900 (O_2900,N_49782,N_49860);
xnor UO_2901 (O_2901,N_49905,N_49919);
or UO_2902 (O_2902,N_49961,N_49770);
nand UO_2903 (O_2903,N_49774,N_49780);
and UO_2904 (O_2904,N_49954,N_49772);
or UO_2905 (O_2905,N_49851,N_49752);
nor UO_2906 (O_2906,N_49817,N_49899);
and UO_2907 (O_2907,N_49903,N_49921);
or UO_2908 (O_2908,N_49755,N_49826);
nand UO_2909 (O_2909,N_49801,N_49753);
nand UO_2910 (O_2910,N_49919,N_49880);
or UO_2911 (O_2911,N_49780,N_49800);
xor UO_2912 (O_2912,N_49830,N_49981);
or UO_2913 (O_2913,N_49940,N_49838);
nor UO_2914 (O_2914,N_49883,N_49814);
nor UO_2915 (O_2915,N_49769,N_49917);
and UO_2916 (O_2916,N_49901,N_49755);
xor UO_2917 (O_2917,N_49828,N_49840);
nand UO_2918 (O_2918,N_49821,N_49859);
xor UO_2919 (O_2919,N_49905,N_49945);
nand UO_2920 (O_2920,N_49812,N_49838);
xor UO_2921 (O_2921,N_49980,N_49837);
and UO_2922 (O_2922,N_49995,N_49857);
or UO_2923 (O_2923,N_49978,N_49840);
nor UO_2924 (O_2924,N_49842,N_49996);
and UO_2925 (O_2925,N_49801,N_49804);
or UO_2926 (O_2926,N_49826,N_49995);
or UO_2927 (O_2927,N_49952,N_49991);
nor UO_2928 (O_2928,N_49792,N_49990);
xnor UO_2929 (O_2929,N_49802,N_49961);
and UO_2930 (O_2930,N_49879,N_49847);
nand UO_2931 (O_2931,N_49813,N_49788);
and UO_2932 (O_2932,N_49758,N_49850);
and UO_2933 (O_2933,N_49966,N_49985);
or UO_2934 (O_2934,N_49861,N_49966);
nand UO_2935 (O_2935,N_49860,N_49750);
nor UO_2936 (O_2936,N_49854,N_49915);
xnor UO_2937 (O_2937,N_49902,N_49991);
nand UO_2938 (O_2938,N_49879,N_49830);
and UO_2939 (O_2939,N_49958,N_49781);
and UO_2940 (O_2940,N_49811,N_49857);
nand UO_2941 (O_2941,N_49854,N_49922);
or UO_2942 (O_2942,N_49962,N_49821);
or UO_2943 (O_2943,N_49911,N_49779);
and UO_2944 (O_2944,N_49899,N_49801);
xor UO_2945 (O_2945,N_49762,N_49845);
xor UO_2946 (O_2946,N_49833,N_49896);
or UO_2947 (O_2947,N_49930,N_49937);
nor UO_2948 (O_2948,N_49861,N_49971);
and UO_2949 (O_2949,N_49862,N_49926);
nand UO_2950 (O_2950,N_49785,N_49964);
nor UO_2951 (O_2951,N_49924,N_49933);
nor UO_2952 (O_2952,N_49765,N_49931);
nand UO_2953 (O_2953,N_49795,N_49819);
nand UO_2954 (O_2954,N_49997,N_49968);
and UO_2955 (O_2955,N_49900,N_49850);
nor UO_2956 (O_2956,N_49948,N_49994);
nor UO_2957 (O_2957,N_49976,N_49793);
nor UO_2958 (O_2958,N_49987,N_49952);
nor UO_2959 (O_2959,N_49779,N_49908);
nand UO_2960 (O_2960,N_49996,N_49883);
nand UO_2961 (O_2961,N_49772,N_49814);
nor UO_2962 (O_2962,N_49766,N_49896);
and UO_2963 (O_2963,N_49765,N_49910);
and UO_2964 (O_2964,N_49756,N_49836);
nand UO_2965 (O_2965,N_49999,N_49837);
xor UO_2966 (O_2966,N_49904,N_49836);
and UO_2967 (O_2967,N_49984,N_49762);
nand UO_2968 (O_2968,N_49814,N_49886);
xnor UO_2969 (O_2969,N_49761,N_49968);
nand UO_2970 (O_2970,N_49941,N_49875);
or UO_2971 (O_2971,N_49922,N_49957);
nor UO_2972 (O_2972,N_49798,N_49920);
xor UO_2973 (O_2973,N_49911,N_49895);
and UO_2974 (O_2974,N_49905,N_49781);
nand UO_2975 (O_2975,N_49771,N_49982);
and UO_2976 (O_2976,N_49941,N_49793);
xor UO_2977 (O_2977,N_49815,N_49765);
and UO_2978 (O_2978,N_49752,N_49971);
nor UO_2979 (O_2979,N_49974,N_49943);
nand UO_2980 (O_2980,N_49900,N_49807);
nor UO_2981 (O_2981,N_49968,N_49953);
xnor UO_2982 (O_2982,N_49939,N_49821);
nor UO_2983 (O_2983,N_49805,N_49818);
nor UO_2984 (O_2984,N_49807,N_49966);
xnor UO_2985 (O_2985,N_49864,N_49892);
and UO_2986 (O_2986,N_49863,N_49954);
nand UO_2987 (O_2987,N_49826,N_49891);
xnor UO_2988 (O_2988,N_49859,N_49750);
nand UO_2989 (O_2989,N_49924,N_49865);
nand UO_2990 (O_2990,N_49974,N_49825);
nand UO_2991 (O_2991,N_49867,N_49839);
nor UO_2992 (O_2992,N_49763,N_49903);
xnor UO_2993 (O_2993,N_49830,N_49836);
nand UO_2994 (O_2994,N_49905,N_49939);
and UO_2995 (O_2995,N_49832,N_49762);
or UO_2996 (O_2996,N_49970,N_49805);
nor UO_2997 (O_2997,N_49837,N_49978);
and UO_2998 (O_2998,N_49756,N_49771);
xor UO_2999 (O_2999,N_49931,N_49818);
and UO_3000 (O_3000,N_49946,N_49873);
or UO_3001 (O_3001,N_49776,N_49789);
or UO_3002 (O_3002,N_49913,N_49993);
xnor UO_3003 (O_3003,N_49994,N_49856);
xor UO_3004 (O_3004,N_49885,N_49847);
nand UO_3005 (O_3005,N_49953,N_49811);
nand UO_3006 (O_3006,N_49959,N_49816);
nor UO_3007 (O_3007,N_49851,N_49979);
nand UO_3008 (O_3008,N_49933,N_49828);
or UO_3009 (O_3009,N_49986,N_49907);
nor UO_3010 (O_3010,N_49980,N_49775);
nor UO_3011 (O_3011,N_49913,N_49895);
and UO_3012 (O_3012,N_49823,N_49858);
or UO_3013 (O_3013,N_49752,N_49880);
nand UO_3014 (O_3014,N_49843,N_49859);
nand UO_3015 (O_3015,N_49945,N_49983);
and UO_3016 (O_3016,N_49809,N_49946);
nand UO_3017 (O_3017,N_49945,N_49932);
xnor UO_3018 (O_3018,N_49967,N_49980);
xor UO_3019 (O_3019,N_49821,N_49805);
and UO_3020 (O_3020,N_49861,N_49877);
nor UO_3021 (O_3021,N_49818,N_49846);
nor UO_3022 (O_3022,N_49862,N_49821);
or UO_3023 (O_3023,N_49909,N_49953);
or UO_3024 (O_3024,N_49766,N_49888);
and UO_3025 (O_3025,N_49925,N_49853);
or UO_3026 (O_3026,N_49813,N_49921);
or UO_3027 (O_3027,N_49828,N_49750);
nor UO_3028 (O_3028,N_49980,N_49929);
or UO_3029 (O_3029,N_49883,N_49906);
xor UO_3030 (O_3030,N_49829,N_49924);
nor UO_3031 (O_3031,N_49753,N_49842);
and UO_3032 (O_3032,N_49853,N_49946);
nor UO_3033 (O_3033,N_49886,N_49997);
or UO_3034 (O_3034,N_49863,N_49891);
xnor UO_3035 (O_3035,N_49865,N_49925);
and UO_3036 (O_3036,N_49874,N_49780);
nand UO_3037 (O_3037,N_49915,N_49935);
nor UO_3038 (O_3038,N_49892,N_49980);
nand UO_3039 (O_3039,N_49938,N_49795);
nand UO_3040 (O_3040,N_49853,N_49941);
or UO_3041 (O_3041,N_49820,N_49919);
or UO_3042 (O_3042,N_49884,N_49905);
or UO_3043 (O_3043,N_49832,N_49950);
and UO_3044 (O_3044,N_49795,N_49856);
nor UO_3045 (O_3045,N_49899,N_49917);
and UO_3046 (O_3046,N_49944,N_49955);
nand UO_3047 (O_3047,N_49859,N_49962);
and UO_3048 (O_3048,N_49829,N_49915);
or UO_3049 (O_3049,N_49758,N_49936);
and UO_3050 (O_3050,N_49858,N_49798);
or UO_3051 (O_3051,N_49773,N_49908);
and UO_3052 (O_3052,N_49807,N_49882);
xor UO_3053 (O_3053,N_49811,N_49932);
and UO_3054 (O_3054,N_49818,N_49836);
nor UO_3055 (O_3055,N_49792,N_49862);
nand UO_3056 (O_3056,N_49750,N_49944);
nor UO_3057 (O_3057,N_49946,N_49827);
nor UO_3058 (O_3058,N_49885,N_49821);
or UO_3059 (O_3059,N_49859,N_49827);
and UO_3060 (O_3060,N_49857,N_49879);
or UO_3061 (O_3061,N_49928,N_49898);
or UO_3062 (O_3062,N_49970,N_49881);
nor UO_3063 (O_3063,N_49983,N_49957);
nand UO_3064 (O_3064,N_49975,N_49970);
nand UO_3065 (O_3065,N_49852,N_49809);
nand UO_3066 (O_3066,N_49802,N_49755);
nand UO_3067 (O_3067,N_49870,N_49896);
nand UO_3068 (O_3068,N_49927,N_49923);
nand UO_3069 (O_3069,N_49793,N_49929);
xor UO_3070 (O_3070,N_49946,N_49927);
xor UO_3071 (O_3071,N_49864,N_49804);
and UO_3072 (O_3072,N_49992,N_49782);
and UO_3073 (O_3073,N_49967,N_49973);
xor UO_3074 (O_3074,N_49957,N_49873);
nor UO_3075 (O_3075,N_49826,N_49873);
nand UO_3076 (O_3076,N_49830,N_49846);
or UO_3077 (O_3077,N_49876,N_49901);
xor UO_3078 (O_3078,N_49757,N_49806);
and UO_3079 (O_3079,N_49809,N_49756);
or UO_3080 (O_3080,N_49897,N_49789);
and UO_3081 (O_3081,N_49841,N_49954);
and UO_3082 (O_3082,N_49793,N_49989);
nor UO_3083 (O_3083,N_49750,N_49905);
nand UO_3084 (O_3084,N_49788,N_49961);
xor UO_3085 (O_3085,N_49969,N_49788);
xnor UO_3086 (O_3086,N_49788,N_49858);
nor UO_3087 (O_3087,N_49947,N_49788);
and UO_3088 (O_3088,N_49964,N_49865);
nand UO_3089 (O_3089,N_49975,N_49989);
or UO_3090 (O_3090,N_49927,N_49954);
and UO_3091 (O_3091,N_49944,N_49897);
nand UO_3092 (O_3092,N_49792,N_49915);
xnor UO_3093 (O_3093,N_49839,N_49779);
nor UO_3094 (O_3094,N_49956,N_49918);
nor UO_3095 (O_3095,N_49857,N_49758);
nor UO_3096 (O_3096,N_49932,N_49919);
or UO_3097 (O_3097,N_49932,N_49873);
or UO_3098 (O_3098,N_49922,N_49808);
nand UO_3099 (O_3099,N_49791,N_49942);
or UO_3100 (O_3100,N_49972,N_49785);
xnor UO_3101 (O_3101,N_49958,N_49762);
nor UO_3102 (O_3102,N_49983,N_49772);
and UO_3103 (O_3103,N_49758,N_49908);
and UO_3104 (O_3104,N_49771,N_49987);
xor UO_3105 (O_3105,N_49948,N_49967);
and UO_3106 (O_3106,N_49867,N_49760);
xnor UO_3107 (O_3107,N_49793,N_49804);
nand UO_3108 (O_3108,N_49879,N_49778);
and UO_3109 (O_3109,N_49995,N_49865);
or UO_3110 (O_3110,N_49861,N_49995);
nand UO_3111 (O_3111,N_49940,N_49783);
or UO_3112 (O_3112,N_49884,N_49772);
and UO_3113 (O_3113,N_49904,N_49933);
or UO_3114 (O_3114,N_49976,N_49825);
and UO_3115 (O_3115,N_49963,N_49936);
and UO_3116 (O_3116,N_49863,N_49948);
or UO_3117 (O_3117,N_49794,N_49905);
nor UO_3118 (O_3118,N_49803,N_49902);
nand UO_3119 (O_3119,N_49797,N_49889);
nor UO_3120 (O_3120,N_49916,N_49766);
and UO_3121 (O_3121,N_49752,N_49789);
xor UO_3122 (O_3122,N_49820,N_49987);
or UO_3123 (O_3123,N_49767,N_49933);
nand UO_3124 (O_3124,N_49859,N_49857);
nand UO_3125 (O_3125,N_49900,N_49796);
and UO_3126 (O_3126,N_49895,N_49950);
or UO_3127 (O_3127,N_49974,N_49996);
nor UO_3128 (O_3128,N_49980,N_49863);
nand UO_3129 (O_3129,N_49774,N_49874);
xnor UO_3130 (O_3130,N_49925,N_49791);
or UO_3131 (O_3131,N_49854,N_49963);
xnor UO_3132 (O_3132,N_49894,N_49955);
nand UO_3133 (O_3133,N_49814,N_49942);
and UO_3134 (O_3134,N_49956,N_49762);
nor UO_3135 (O_3135,N_49751,N_49909);
xor UO_3136 (O_3136,N_49990,N_49912);
nor UO_3137 (O_3137,N_49904,N_49866);
nor UO_3138 (O_3138,N_49855,N_49915);
or UO_3139 (O_3139,N_49855,N_49750);
or UO_3140 (O_3140,N_49896,N_49941);
xor UO_3141 (O_3141,N_49932,N_49803);
nor UO_3142 (O_3142,N_49965,N_49897);
xor UO_3143 (O_3143,N_49765,N_49801);
or UO_3144 (O_3144,N_49790,N_49840);
nand UO_3145 (O_3145,N_49981,N_49891);
or UO_3146 (O_3146,N_49898,N_49984);
xor UO_3147 (O_3147,N_49785,N_49841);
and UO_3148 (O_3148,N_49937,N_49850);
xor UO_3149 (O_3149,N_49850,N_49977);
nand UO_3150 (O_3150,N_49766,N_49814);
xor UO_3151 (O_3151,N_49885,N_49817);
and UO_3152 (O_3152,N_49860,N_49935);
and UO_3153 (O_3153,N_49963,N_49969);
nor UO_3154 (O_3154,N_49760,N_49756);
and UO_3155 (O_3155,N_49948,N_49896);
or UO_3156 (O_3156,N_49757,N_49770);
nand UO_3157 (O_3157,N_49774,N_49765);
nor UO_3158 (O_3158,N_49771,N_49826);
or UO_3159 (O_3159,N_49755,N_49947);
and UO_3160 (O_3160,N_49857,N_49955);
xnor UO_3161 (O_3161,N_49811,N_49844);
nor UO_3162 (O_3162,N_49986,N_49861);
xnor UO_3163 (O_3163,N_49813,N_49751);
nor UO_3164 (O_3164,N_49844,N_49881);
xnor UO_3165 (O_3165,N_49796,N_49917);
nand UO_3166 (O_3166,N_49839,N_49834);
or UO_3167 (O_3167,N_49869,N_49855);
and UO_3168 (O_3168,N_49866,N_49945);
or UO_3169 (O_3169,N_49772,N_49881);
xnor UO_3170 (O_3170,N_49921,N_49998);
nor UO_3171 (O_3171,N_49956,N_49965);
or UO_3172 (O_3172,N_49956,N_49941);
nand UO_3173 (O_3173,N_49968,N_49899);
nand UO_3174 (O_3174,N_49888,N_49984);
or UO_3175 (O_3175,N_49806,N_49789);
xor UO_3176 (O_3176,N_49878,N_49781);
nor UO_3177 (O_3177,N_49808,N_49884);
nor UO_3178 (O_3178,N_49918,N_49817);
nor UO_3179 (O_3179,N_49786,N_49817);
and UO_3180 (O_3180,N_49917,N_49794);
xor UO_3181 (O_3181,N_49835,N_49911);
or UO_3182 (O_3182,N_49993,N_49969);
or UO_3183 (O_3183,N_49873,N_49884);
nor UO_3184 (O_3184,N_49957,N_49966);
nand UO_3185 (O_3185,N_49988,N_49751);
and UO_3186 (O_3186,N_49944,N_49833);
and UO_3187 (O_3187,N_49867,N_49935);
nand UO_3188 (O_3188,N_49825,N_49785);
or UO_3189 (O_3189,N_49896,N_49904);
xnor UO_3190 (O_3190,N_49977,N_49933);
or UO_3191 (O_3191,N_49850,N_49784);
or UO_3192 (O_3192,N_49871,N_49959);
and UO_3193 (O_3193,N_49840,N_49867);
nand UO_3194 (O_3194,N_49925,N_49978);
nand UO_3195 (O_3195,N_49875,N_49766);
nand UO_3196 (O_3196,N_49938,N_49750);
nand UO_3197 (O_3197,N_49941,N_49904);
and UO_3198 (O_3198,N_49893,N_49905);
nand UO_3199 (O_3199,N_49904,N_49956);
nor UO_3200 (O_3200,N_49980,N_49960);
xor UO_3201 (O_3201,N_49875,N_49912);
or UO_3202 (O_3202,N_49872,N_49913);
or UO_3203 (O_3203,N_49819,N_49954);
nor UO_3204 (O_3204,N_49970,N_49979);
or UO_3205 (O_3205,N_49822,N_49768);
or UO_3206 (O_3206,N_49879,N_49998);
nor UO_3207 (O_3207,N_49884,N_49852);
or UO_3208 (O_3208,N_49994,N_49804);
or UO_3209 (O_3209,N_49752,N_49888);
xnor UO_3210 (O_3210,N_49868,N_49820);
or UO_3211 (O_3211,N_49821,N_49936);
nor UO_3212 (O_3212,N_49888,N_49873);
or UO_3213 (O_3213,N_49848,N_49886);
nand UO_3214 (O_3214,N_49802,N_49998);
nor UO_3215 (O_3215,N_49947,N_49914);
or UO_3216 (O_3216,N_49822,N_49933);
or UO_3217 (O_3217,N_49850,N_49936);
or UO_3218 (O_3218,N_49915,N_49955);
nand UO_3219 (O_3219,N_49952,N_49995);
nor UO_3220 (O_3220,N_49902,N_49950);
xnor UO_3221 (O_3221,N_49951,N_49906);
nand UO_3222 (O_3222,N_49787,N_49929);
nand UO_3223 (O_3223,N_49927,N_49834);
nor UO_3224 (O_3224,N_49948,N_49976);
nand UO_3225 (O_3225,N_49954,N_49796);
nor UO_3226 (O_3226,N_49872,N_49798);
xnor UO_3227 (O_3227,N_49933,N_49995);
or UO_3228 (O_3228,N_49753,N_49755);
nand UO_3229 (O_3229,N_49890,N_49788);
nor UO_3230 (O_3230,N_49868,N_49814);
xnor UO_3231 (O_3231,N_49936,N_49839);
or UO_3232 (O_3232,N_49958,N_49940);
or UO_3233 (O_3233,N_49825,N_49842);
nor UO_3234 (O_3234,N_49985,N_49795);
nor UO_3235 (O_3235,N_49757,N_49763);
xor UO_3236 (O_3236,N_49924,N_49997);
xnor UO_3237 (O_3237,N_49940,N_49788);
nand UO_3238 (O_3238,N_49914,N_49896);
nor UO_3239 (O_3239,N_49983,N_49858);
nor UO_3240 (O_3240,N_49929,N_49948);
nor UO_3241 (O_3241,N_49909,N_49976);
xnor UO_3242 (O_3242,N_49973,N_49991);
nand UO_3243 (O_3243,N_49896,N_49935);
nor UO_3244 (O_3244,N_49775,N_49767);
nand UO_3245 (O_3245,N_49870,N_49795);
or UO_3246 (O_3246,N_49952,N_49940);
nor UO_3247 (O_3247,N_49807,N_49876);
xor UO_3248 (O_3248,N_49858,N_49922);
nor UO_3249 (O_3249,N_49836,N_49823);
nand UO_3250 (O_3250,N_49823,N_49990);
xnor UO_3251 (O_3251,N_49772,N_49882);
xnor UO_3252 (O_3252,N_49947,N_49899);
or UO_3253 (O_3253,N_49767,N_49883);
or UO_3254 (O_3254,N_49890,N_49962);
xor UO_3255 (O_3255,N_49856,N_49760);
nand UO_3256 (O_3256,N_49849,N_49763);
xor UO_3257 (O_3257,N_49970,N_49989);
nand UO_3258 (O_3258,N_49837,N_49895);
and UO_3259 (O_3259,N_49863,N_49766);
and UO_3260 (O_3260,N_49778,N_49887);
or UO_3261 (O_3261,N_49904,N_49870);
nand UO_3262 (O_3262,N_49906,N_49790);
xor UO_3263 (O_3263,N_49997,N_49883);
nand UO_3264 (O_3264,N_49859,N_49938);
nand UO_3265 (O_3265,N_49990,N_49758);
nor UO_3266 (O_3266,N_49922,N_49752);
and UO_3267 (O_3267,N_49922,N_49802);
xnor UO_3268 (O_3268,N_49872,N_49750);
nand UO_3269 (O_3269,N_49793,N_49982);
and UO_3270 (O_3270,N_49998,N_49895);
nand UO_3271 (O_3271,N_49982,N_49983);
xor UO_3272 (O_3272,N_49941,N_49967);
or UO_3273 (O_3273,N_49826,N_49776);
and UO_3274 (O_3274,N_49844,N_49893);
or UO_3275 (O_3275,N_49977,N_49790);
nand UO_3276 (O_3276,N_49773,N_49990);
nand UO_3277 (O_3277,N_49931,N_49782);
xnor UO_3278 (O_3278,N_49972,N_49777);
nand UO_3279 (O_3279,N_49977,N_49878);
and UO_3280 (O_3280,N_49835,N_49937);
and UO_3281 (O_3281,N_49793,N_49944);
nor UO_3282 (O_3282,N_49914,N_49879);
nand UO_3283 (O_3283,N_49972,N_49940);
nor UO_3284 (O_3284,N_49864,N_49918);
and UO_3285 (O_3285,N_49857,N_49996);
and UO_3286 (O_3286,N_49865,N_49947);
nor UO_3287 (O_3287,N_49996,N_49876);
xor UO_3288 (O_3288,N_49912,N_49819);
or UO_3289 (O_3289,N_49754,N_49838);
nor UO_3290 (O_3290,N_49773,N_49764);
nand UO_3291 (O_3291,N_49940,N_49840);
xnor UO_3292 (O_3292,N_49887,N_49859);
and UO_3293 (O_3293,N_49828,N_49849);
xor UO_3294 (O_3294,N_49927,N_49782);
nor UO_3295 (O_3295,N_49874,N_49967);
or UO_3296 (O_3296,N_49981,N_49761);
xor UO_3297 (O_3297,N_49807,N_49833);
nor UO_3298 (O_3298,N_49896,N_49790);
and UO_3299 (O_3299,N_49968,N_49868);
xnor UO_3300 (O_3300,N_49869,N_49783);
xor UO_3301 (O_3301,N_49809,N_49866);
nand UO_3302 (O_3302,N_49767,N_49761);
nand UO_3303 (O_3303,N_49976,N_49960);
nor UO_3304 (O_3304,N_49837,N_49887);
and UO_3305 (O_3305,N_49856,N_49840);
or UO_3306 (O_3306,N_49868,N_49832);
nor UO_3307 (O_3307,N_49962,N_49942);
nand UO_3308 (O_3308,N_49775,N_49888);
nor UO_3309 (O_3309,N_49997,N_49952);
xnor UO_3310 (O_3310,N_49932,N_49758);
or UO_3311 (O_3311,N_49958,N_49795);
nand UO_3312 (O_3312,N_49961,N_49980);
nor UO_3313 (O_3313,N_49841,N_49788);
nor UO_3314 (O_3314,N_49839,N_49971);
or UO_3315 (O_3315,N_49836,N_49759);
nor UO_3316 (O_3316,N_49955,N_49980);
or UO_3317 (O_3317,N_49898,N_49903);
nor UO_3318 (O_3318,N_49770,N_49902);
nor UO_3319 (O_3319,N_49879,N_49782);
nand UO_3320 (O_3320,N_49798,N_49894);
and UO_3321 (O_3321,N_49951,N_49954);
xor UO_3322 (O_3322,N_49874,N_49861);
nand UO_3323 (O_3323,N_49980,N_49880);
nand UO_3324 (O_3324,N_49791,N_49752);
and UO_3325 (O_3325,N_49816,N_49855);
or UO_3326 (O_3326,N_49957,N_49960);
xor UO_3327 (O_3327,N_49757,N_49766);
xor UO_3328 (O_3328,N_49762,N_49944);
and UO_3329 (O_3329,N_49936,N_49750);
xnor UO_3330 (O_3330,N_49883,N_49884);
or UO_3331 (O_3331,N_49766,N_49790);
xnor UO_3332 (O_3332,N_49917,N_49822);
nand UO_3333 (O_3333,N_49872,N_49796);
nor UO_3334 (O_3334,N_49780,N_49997);
nor UO_3335 (O_3335,N_49986,N_49998);
or UO_3336 (O_3336,N_49751,N_49934);
xor UO_3337 (O_3337,N_49965,N_49841);
and UO_3338 (O_3338,N_49886,N_49750);
nand UO_3339 (O_3339,N_49876,N_49961);
or UO_3340 (O_3340,N_49942,N_49976);
nor UO_3341 (O_3341,N_49807,N_49880);
and UO_3342 (O_3342,N_49784,N_49789);
nand UO_3343 (O_3343,N_49759,N_49917);
and UO_3344 (O_3344,N_49809,N_49865);
nand UO_3345 (O_3345,N_49870,N_49785);
xor UO_3346 (O_3346,N_49777,N_49938);
nor UO_3347 (O_3347,N_49891,N_49788);
or UO_3348 (O_3348,N_49795,N_49935);
and UO_3349 (O_3349,N_49976,N_49767);
and UO_3350 (O_3350,N_49939,N_49906);
or UO_3351 (O_3351,N_49829,N_49772);
and UO_3352 (O_3352,N_49782,N_49955);
and UO_3353 (O_3353,N_49947,N_49993);
and UO_3354 (O_3354,N_49876,N_49843);
or UO_3355 (O_3355,N_49814,N_49760);
and UO_3356 (O_3356,N_49915,N_49764);
and UO_3357 (O_3357,N_49808,N_49881);
xor UO_3358 (O_3358,N_49808,N_49956);
or UO_3359 (O_3359,N_49960,N_49795);
xor UO_3360 (O_3360,N_49842,N_49789);
nor UO_3361 (O_3361,N_49787,N_49911);
and UO_3362 (O_3362,N_49873,N_49960);
nand UO_3363 (O_3363,N_49847,N_49934);
or UO_3364 (O_3364,N_49933,N_49811);
and UO_3365 (O_3365,N_49865,N_49885);
nor UO_3366 (O_3366,N_49839,N_49908);
or UO_3367 (O_3367,N_49802,N_49997);
or UO_3368 (O_3368,N_49758,N_49947);
xnor UO_3369 (O_3369,N_49857,N_49960);
and UO_3370 (O_3370,N_49868,N_49859);
or UO_3371 (O_3371,N_49828,N_49870);
and UO_3372 (O_3372,N_49821,N_49968);
nor UO_3373 (O_3373,N_49912,N_49763);
xnor UO_3374 (O_3374,N_49911,N_49983);
or UO_3375 (O_3375,N_49969,N_49948);
and UO_3376 (O_3376,N_49911,N_49962);
or UO_3377 (O_3377,N_49836,N_49890);
nor UO_3378 (O_3378,N_49894,N_49897);
nor UO_3379 (O_3379,N_49938,N_49870);
xnor UO_3380 (O_3380,N_49905,N_49879);
nand UO_3381 (O_3381,N_49931,N_49873);
xnor UO_3382 (O_3382,N_49872,N_49799);
xnor UO_3383 (O_3383,N_49870,N_49884);
xnor UO_3384 (O_3384,N_49909,N_49839);
nor UO_3385 (O_3385,N_49818,N_49944);
nor UO_3386 (O_3386,N_49948,N_49907);
or UO_3387 (O_3387,N_49966,N_49872);
nand UO_3388 (O_3388,N_49806,N_49972);
nand UO_3389 (O_3389,N_49950,N_49812);
nor UO_3390 (O_3390,N_49929,N_49903);
or UO_3391 (O_3391,N_49951,N_49901);
xor UO_3392 (O_3392,N_49752,N_49919);
xor UO_3393 (O_3393,N_49808,N_49856);
xnor UO_3394 (O_3394,N_49955,N_49868);
or UO_3395 (O_3395,N_49832,N_49900);
and UO_3396 (O_3396,N_49896,N_49958);
and UO_3397 (O_3397,N_49899,N_49928);
nor UO_3398 (O_3398,N_49842,N_49871);
or UO_3399 (O_3399,N_49815,N_49893);
and UO_3400 (O_3400,N_49986,N_49838);
or UO_3401 (O_3401,N_49831,N_49855);
or UO_3402 (O_3402,N_49866,N_49950);
or UO_3403 (O_3403,N_49947,N_49855);
or UO_3404 (O_3404,N_49872,N_49850);
nor UO_3405 (O_3405,N_49949,N_49862);
nor UO_3406 (O_3406,N_49990,N_49789);
xnor UO_3407 (O_3407,N_49809,N_49995);
and UO_3408 (O_3408,N_49986,N_49769);
xnor UO_3409 (O_3409,N_49856,N_49870);
nand UO_3410 (O_3410,N_49899,N_49783);
nor UO_3411 (O_3411,N_49889,N_49823);
nor UO_3412 (O_3412,N_49966,N_49826);
or UO_3413 (O_3413,N_49988,N_49867);
or UO_3414 (O_3414,N_49849,N_49965);
nor UO_3415 (O_3415,N_49827,N_49837);
nor UO_3416 (O_3416,N_49824,N_49885);
nand UO_3417 (O_3417,N_49778,N_49946);
or UO_3418 (O_3418,N_49792,N_49947);
nor UO_3419 (O_3419,N_49814,N_49884);
nand UO_3420 (O_3420,N_49995,N_49926);
and UO_3421 (O_3421,N_49992,N_49949);
and UO_3422 (O_3422,N_49811,N_49783);
nand UO_3423 (O_3423,N_49804,N_49849);
or UO_3424 (O_3424,N_49790,N_49890);
or UO_3425 (O_3425,N_49898,N_49797);
or UO_3426 (O_3426,N_49911,N_49938);
xnor UO_3427 (O_3427,N_49931,N_49910);
and UO_3428 (O_3428,N_49863,N_49973);
nor UO_3429 (O_3429,N_49984,N_49889);
and UO_3430 (O_3430,N_49960,N_49947);
or UO_3431 (O_3431,N_49956,N_49766);
nor UO_3432 (O_3432,N_49775,N_49849);
nand UO_3433 (O_3433,N_49886,N_49882);
and UO_3434 (O_3434,N_49856,N_49805);
nor UO_3435 (O_3435,N_49866,N_49777);
xor UO_3436 (O_3436,N_49920,N_49761);
nor UO_3437 (O_3437,N_49900,N_49771);
xnor UO_3438 (O_3438,N_49773,N_49956);
xnor UO_3439 (O_3439,N_49996,N_49911);
xor UO_3440 (O_3440,N_49862,N_49981);
or UO_3441 (O_3441,N_49866,N_49850);
nor UO_3442 (O_3442,N_49841,N_49848);
xor UO_3443 (O_3443,N_49945,N_49839);
xor UO_3444 (O_3444,N_49950,N_49988);
nand UO_3445 (O_3445,N_49761,N_49967);
and UO_3446 (O_3446,N_49929,N_49873);
and UO_3447 (O_3447,N_49797,N_49840);
xnor UO_3448 (O_3448,N_49854,N_49797);
nor UO_3449 (O_3449,N_49762,N_49757);
xor UO_3450 (O_3450,N_49923,N_49826);
xor UO_3451 (O_3451,N_49968,N_49993);
nor UO_3452 (O_3452,N_49776,N_49902);
nor UO_3453 (O_3453,N_49853,N_49957);
or UO_3454 (O_3454,N_49855,N_49921);
and UO_3455 (O_3455,N_49911,N_49941);
xor UO_3456 (O_3456,N_49993,N_49827);
nand UO_3457 (O_3457,N_49794,N_49837);
nor UO_3458 (O_3458,N_49825,N_49799);
and UO_3459 (O_3459,N_49942,N_49775);
nand UO_3460 (O_3460,N_49983,N_49823);
nor UO_3461 (O_3461,N_49883,N_49829);
or UO_3462 (O_3462,N_49866,N_49849);
nand UO_3463 (O_3463,N_49773,N_49837);
xor UO_3464 (O_3464,N_49917,N_49856);
and UO_3465 (O_3465,N_49931,N_49915);
nand UO_3466 (O_3466,N_49819,N_49982);
nor UO_3467 (O_3467,N_49951,N_49774);
nor UO_3468 (O_3468,N_49865,N_49768);
or UO_3469 (O_3469,N_49945,N_49965);
nor UO_3470 (O_3470,N_49754,N_49873);
or UO_3471 (O_3471,N_49806,N_49927);
and UO_3472 (O_3472,N_49865,N_49823);
or UO_3473 (O_3473,N_49753,N_49835);
or UO_3474 (O_3474,N_49835,N_49938);
or UO_3475 (O_3475,N_49796,N_49863);
xnor UO_3476 (O_3476,N_49929,N_49863);
nor UO_3477 (O_3477,N_49964,N_49935);
or UO_3478 (O_3478,N_49782,N_49866);
or UO_3479 (O_3479,N_49766,N_49752);
or UO_3480 (O_3480,N_49758,N_49925);
nor UO_3481 (O_3481,N_49989,N_49752);
or UO_3482 (O_3482,N_49934,N_49919);
xnor UO_3483 (O_3483,N_49805,N_49853);
nand UO_3484 (O_3484,N_49937,N_49939);
xnor UO_3485 (O_3485,N_49948,N_49984);
and UO_3486 (O_3486,N_49913,N_49837);
nand UO_3487 (O_3487,N_49879,N_49878);
nor UO_3488 (O_3488,N_49894,N_49773);
and UO_3489 (O_3489,N_49957,N_49956);
nand UO_3490 (O_3490,N_49981,N_49945);
and UO_3491 (O_3491,N_49935,N_49967);
or UO_3492 (O_3492,N_49778,N_49817);
nand UO_3493 (O_3493,N_49826,N_49893);
xnor UO_3494 (O_3494,N_49983,N_49953);
or UO_3495 (O_3495,N_49773,N_49948);
nand UO_3496 (O_3496,N_49782,N_49778);
or UO_3497 (O_3497,N_49855,N_49960);
xnor UO_3498 (O_3498,N_49949,N_49801);
xnor UO_3499 (O_3499,N_49866,N_49934);
and UO_3500 (O_3500,N_49856,N_49875);
nand UO_3501 (O_3501,N_49796,N_49805);
or UO_3502 (O_3502,N_49948,N_49946);
xnor UO_3503 (O_3503,N_49954,N_49861);
nor UO_3504 (O_3504,N_49974,N_49885);
nor UO_3505 (O_3505,N_49976,N_49935);
xnor UO_3506 (O_3506,N_49985,N_49994);
or UO_3507 (O_3507,N_49945,N_49964);
nor UO_3508 (O_3508,N_49793,N_49857);
nor UO_3509 (O_3509,N_49753,N_49812);
xnor UO_3510 (O_3510,N_49886,N_49971);
nor UO_3511 (O_3511,N_49829,N_49819);
and UO_3512 (O_3512,N_49937,N_49953);
nand UO_3513 (O_3513,N_49811,N_49868);
nor UO_3514 (O_3514,N_49860,N_49894);
xor UO_3515 (O_3515,N_49816,N_49818);
or UO_3516 (O_3516,N_49760,N_49940);
or UO_3517 (O_3517,N_49912,N_49935);
or UO_3518 (O_3518,N_49841,N_49960);
nand UO_3519 (O_3519,N_49846,N_49867);
nor UO_3520 (O_3520,N_49875,N_49878);
nand UO_3521 (O_3521,N_49783,N_49922);
nor UO_3522 (O_3522,N_49846,N_49938);
and UO_3523 (O_3523,N_49782,N_49862);
nor UO_3524 (O_3524,N_49983,N_49988);
nand UO_3525 (O_3525,N_49872,N_49778);
nand UO_3526 (O_3526,N_49903,N_49933);
or UO_3527 (O_3527,N_49850,N_49814);
and UO_3528 (O_3528,N_49928,N_49914);
or UO_3529 (O_3529,N_49774,N_49970);
nor UO_3530 (O_3530,N_49861,N_49850);
nor UO_3531 (O_3531,N_49958,N_49864);
or UO_3532 (O_3532,N_49936,N_49808);
nand UO_3533 (O_3533,N_49909,N_49974);
nand UO_3534 (O_3534,N_49848,N_49760);
xor UO_3535 (O_3535,N_49774,N_49775);
xnor UO_3536 (O_3536,N_49836,N_49978);
xnor UO_3537 (O_3537,N_49972,N_49902);
nand UO_3538 (O_3538,N_49874,N_49951);
and UO_3539 (O_3539,N_49819,N_49868);
nand UO_3540 (O_3540,N_49909,N_49842);
xor UO_3541 (O_3541,N_49946,N_49984);
xor UO_3542 (O_3542,N_49979,N_49934);
xnor UO_3543 (O_3543,N_49935,N_49997);
nand UO_3544 (O_3544,N_49952,N_49800);
xor UO_3545 (O_3545,N_49877,N_49750);
nand UO_3546 (O_3546,N_49889,N_49830);
nand UO_3547 (O_3547,N_49902,N_49771);
xor UO_3548 (O_3548,N_49812,N_49754);
or UO_3549 (O_3549,N_49798,N_49926);
and UO_3550 (O_3550,N_49980,N_49859);
or UO_3551 (O_3551,N_49970,N_49875);
or UO_3552 (O_3552,N_49916,N_49908);
nor UO_3553 (O_3553,N_49908,N_49771);
nor UO_3554 (O_3554,N_49890,N_49761);
xor UO_3555 (O_3555,N_49863,N_49874);
and UO_3556 (O_3556,N_49969,N_49961);
xor UO_3557 (O_3557,N_49907,N_49872);
and UO_3558 (O_3558,N_49869,N_49817);
and UO_3559 (O_3559,N_49772,N_49841);
nor UO_3560 (O_3560,N_49896,N_49903);
or UO_3561 (O_3561,N_49779,N_49835);
or UO_3562 (O_3562,N_49873,N_49981);
nand UO_3563 (O_3563,N_49807,N_49951);
and UO_3564 (O_3564,N_49774,N_49987);
or UO_3565 (O_3565,N_49776,N_49778);
and UO_3566 (O_3566,N_49962,N_49788);
nor UO_3567 (O_3567,N_49862,N_49798);
and UO_3568 (O_3568,N_49778,N_49842);
and UO_3569 (O_3569,N_49902,N_49966);
nor UO_3570 (O_3570,N_49788,N_49948);
and UO_3571 (O_3571,N_49915,N_49869);
nor UO_3572 (O_3572,N_49811,N_49904);
xor UO_3573 (O_3573,N_49854,N_49862);
and UO_3574 (O_3574,N_49980,N_49995);
nor UO_3575 (O_3575,N_49869,N_49820);
and UO_3576 (O_3576,N_49890,N_49940);
or UO_3577 (O_3577,N_49875,N_49978);
nand UO_3578 (O_3578,N_49832,N_49935);
or UO_3579 (O_3579,N_49838,N_49796);
nand UO_3580 (O_3580,N_49766,N_49949);
and UO_3581 (O_3581,N_49862,N_49757);
or UO_3582 (O_3582,N_49950,N_49852);
xor UO_3583 (O_3583,N_49887,N_49888);
nor UO_3584 (O_3584,N_49982,N_49928);
and UO_3585 (O_3585,N_49889,N_49965);
and UO_3586 (O_3586,N_49926,N_49890);
and UO_3587 (O_3587,N_49995,N_49763);
xor UO_3588 (O_3588,N_49989,N_49999);
and UO_3589 (O_3589,N_49877,N_49819);
and UO_3590 (O_3590,N_49929,N_49891);
nor UO_3591 (O_3591,N_49760,N_49933);
xor UO_3592 (O_3592,N_49805,N_49920);
nor UO_3593 (O_3593,N_49884,N_49875);
nor UO_3594 (O_3594,N_49936,N_49996);
and UO_3595 (O_3595,N_49887,N_49895);
and UO_3596 (O_3596,N_49981,N_49812);
nand UO_3597 (O_3597,N_49826,N_49849);
xnor UO_3598 (O_3598,N_49773,N_49877);
nand UO_3599 (O_3599,N_49826,N_49903);
nor UO_3600 (O_3600,N_49823,N_49765);
nand UO_3601 (O_3601,N_49897,N_49777);
nor UO_3602 (O_3602,N_49767,N_49865);
xor UO_3603 (O_3603,N_49823,N_49830);
nor UO_3604 (O_3604,N_49861,N_49799);
or UO_3605 (O_3605,N_49983,N_49974);
nor UO_3606 (O_3606,N_49854,N_49938);
nor UO_3607 (O_3607,N_49989,N_49866);
nand UO_3608 (O_3608,N_49886,N_49775);
or UO_3609 (O_3609,N_49814,N_49856);
and UO_3610 (O_3610,N_49969,N_49976);
or UO_3611 (O_3611,N_49950,N_49900);
and UO_3612 (O_3612,N_49979,N_49752);
or UO_3613 (O_3613,N_49861,N_49931);
nand UO_3614 (O_3614,N_49932,N_49983);
or UO_3615 (O_3615,N_49940,N_49906);
or UO_3616 (O_3616,N_49948,N_49975);
xor UO_3617 (O_3617,N_49865,N_49906);
or UO_3618 (O_3618,N_49943,N_49798);
nand UO_3619 (O_3619,N_49835,N_49941);
nor UO_3620 (O_3620,N_49915,N_49923);
xor UO_3621 (O_3621,N_49788,N_49824);
nand UO_3622 (O_3622,N_49769,N_49968);
nand UO_3623 (O_3623,N_49801,N_49791);
or UO_3624 (O_3624,N_49818,N_49792);
xnor UO_3625 (O_3625,N_49878,N_49877);
xor UO_3626 (O_3626,N_49825,N_49922);
and UO_3627 (O_3627,N_49820,N_49936);
or UO_3628 (O_3628,N_49987,N_49877);
and UO_3629 (O_3629,N_49810,N_49868);
and UO_3630 (O_3630,N_49936,N_49900);
nor UO_3631 (O_3631,N_49988,N_49931);
or UO_3632 (O_3632,N_49897,N_49815);
nand UO_3633 (O_3633,N_49781,N_49965);
nand UO_3634 (O_3634,N_49765,N_49795);
or UO_3635 (O_3635,N_49852,N_49932);
or UO_3636 (O_3636,N_49846,N_49891);
nor UO_3637 (O_3637,N_49788,N_49823);
or UO_3638 (O_3638,N_49908,N_49887);
and UO_3639 (O_3639,N_49792,N_49760);
and UO_3640 (O_3640,N_49769,N_49819);
xnor UO_3641 (O_3641,N_49998,N_49854);
or UO_3642 (O_3642,N_49923,N_49895);
or UO_3643 (O_3643,N_49894,N_49824);
and UO_3644 (O_3644,N_49860,N_49982);
nand UO_3645 (O_3645,N_49995,N_49869);
or UO_3646 (O_3646,N_49777,N_49872);
xnor UO_3647 (O_3647,N_49973,N_49775);
and UO_3648 (O_3648,N_49786,N_49939);
nor UO_3649 (O_3649,N_49981,N_49952);
and UO_3650 (O_3650,N_49930,N_49958);
and UO_3651 (O_3651,N_49958,N_49932);
and UO_3652 (O_3652,N_49802,N_49973);
or UO_3653 (O_3653,N_49805,N_49768);
and UO_3654 (O_3654,N_49970,N_49762);
xor UO_3655 (O_3655,N_49943,N_49811);
and UO_3656 (O_3656,N_49789,N_49854);
or UO_3657 (O_3657,N_49753,N_49968);
or UO_3658 (O_3658,N_49907,N_49805);
nand UO_3659 (O_3659,N_49764,N_49931);
and UO_3660 (O_3660,N_49769,N_49830);
or UO_3661 (O_3661,N_49819,N_49891);
xnor UO_3662 (O_3662,N_49951,N_49927);
xor UO_3663 (O_3663,N_49963,N_49863);
xnor UO_3664 (O_3664,N_49975,N_49752);
nor UO_3665 (O_3665,N_49967,N_49994);
nor UO_3666 (O_3666,N_49908,N_49772);
nand UO_3667 (O_3667,N_49996,N_49977);
nor UO_3668 (O_3668,N_49873,N_49882);
nand UO_3669 (O_3669,N_49941,N_49752);
xnor UO_3670 (O_3670,N_49821,N_49990);
nand UO_3671 (O_3671,N_49978,N_49971);
xor UO_3672 (O_3672,N_49917,N_49991);
nor UO_3673 (O_3673,N_49960,N_49953);
xnor UO_3674 (O_3674,N_49939,N_49944);
nand UO_3675 (O_3675,N_49856,N_49926);
xnor UO_3676 (O_3676,N_49992,N_49933);
xnor UO_3677 (O_3677,N_49886,N_49865);
xor UO_3678 (O_3678,N_49951,N_49840);
xnor UO_3679 (O_3679,N_49864,N_49767);
nand UO_3680 (O_3680,N_49872,N_49759);
xor UO_3681 (O_3681,N_49803,N_49768);
nor UO_3682 (O_3682,N_49978,N_49970);
xor UO_3683 (O_3683,N_49940,N_49919);
nand UO_3684 (O_3684,N_49998,N_49900);
nand UO_3685 (O_3685,N_49750,N_49791);
nor UO_3686 (O_3686,N_49988,N_49881);
or UO_3687 (O_3687,N_49939,N_49998);
nand UO_3688 (O_3688,N_49932,N_49858);
nand UO_3689 (O_3689,N_49974,N_49770);
nor UO_3690 (O_3690,N_49765,N_49878);
and UO_3691 (O_3691,N_49907,N_49767);
or UO_3692 (O_3692,N_49965,N_49917);
xor UO_3693 (O_3693,N_49914,N_49965);
nand UO_3694 (O_3694,N_49843,N_49892);
nor UO_3695 (O_3695,N_49834,N_49816);
xor UO_3696 (O_3696,N_49781,N_49854);
nand UO_3697 (O_3697,N_49777,N_49877);
and UO_3698 (O_3698,N_49779,N_49950);
nand UO_3699 (O_3699,N_49872,N_49912);
nor UO_3700 (O_3700,N_49934,N_49923);
nand UO_3701 (O_3701,N_49915,N_49956);
nand UO_3702 (O_3702,N_49810,N_49887);
or UO_3703 (O_3703,N_49933,N_49873);
or UO_3704 (O_3704,N_49942,N_49974);
or UO_3705 (O_3705,N_49895,N_49796);
xor UO_3706 (O_3706,N_49835,N_49919);
nor UO_3707 (O_3707,N_49994,N_49757);
and UO_3708 (O_3708,N_49757,N_49884);
or UO_3709 (O_3709,N_49853,N_49959);
and UO_3710 (O_3710,N_49829,N_49902);
and UO_3711 (O_3711,N_49870,N_49984);
nor UO_3712 (O_3712,N_49930,N_49792);
and UO_3713 (O_3713,N_49975,N_49799);
nand UO_3714 (O_3714,N_49972,N_49840);
xor UO_3715 (O_3715,N_49768,N_49831);
xor UO_3716 (O_3716,N_49756,N_49823);
nand UO_3717 (O_3717,N_49852,N_49900);
and UO_3718 (O_3718,N_49900,N_49881);
xor UO_3719 (O_3719,N_49804,N_49934);
xnor UO_3720 (O_3720,N_49850,N_49958);
xor UO_3721 (O_3721,N_49846,N_49993);
xnor UO_3722 (O_3722,N_49954,N_49758);
or UO_3723 (O_3723,N_49927,N_49852);
xnor UO_3724 (O_3724,N_49912,N_49756);
nor UO_3725 (O_3725,N_49845,N_49765);
xor UO_3726 (O_3726,N_49934,N_49909);
or UO_3727 (O_3727,N_49965,N_49787);
or UO_3728 (O_3728,N_49995,N_49895);
xnor UO_3729 (O_3729,N_49797,N_49961);
xor UO_3730 (O_3730,N_49864,N_49790);
nor UO_3731 (O_3731,N_49866,N_49792);
xor UO_3732 (O_3732,N_49826,N_49774);
nor UO_3733 (O_3733,N_49997,N_49994);
nor UO_3734 (O_3734,N_49751,N_49783);
nand UO_3735 (O_3735,N_49938,N_49799);
or UO_3736 (O_3736,N_49865,N_49948);
or UO_3737 (O_3737,N_49757,N_49986);
and UO_3738 (O_3738,N_49763,N_49822);
or UO_3739 (O_3739,N_49952,N_49938);
nor UO_3740 (O_3740,N_49753,N_49820);
and UO_3741 (O_3741,N_49901,N_49963);
or UO_3742 (O_3742,N_49762,N_49932);
or UO_3743 (O_3743,N_49813,N_49967);
nor UO_3744 (O_3744,N_49803,N_49868);
xor UO_3745 (O_3745,N_49809,N_49920);
or UO_3746 (O_3746,N_49796,N_49840);
and UO_3747 (O_3747,N_49821,N_49767);
or UO_3748 (O_3748,N_49817,N_49814);
or UO_3749 (O_3749,N_49995,N_49874);
nand UO_3750 (O_3750,N_49896,N_49778);
nand UO_3751 (O_3751,N_49938,N_49980);
nand UO_3752 (O_3752,N_49951,N_49886);
nand UO_3753 (O_3753,N_49916,N_49761);
nand UO_3754 (O_3754,N_49802,N_49925);
or UO_3755 (O_3755,N_49834,N_49974);
nor UO_3756 (O_3756,N_49849,N_49877);
or UO_3757 (O_3757,N_49819,N_49852);
nand UO_3758 (O_3758,N_49981,N_49855);
or UO_3759 (O_3759,N_49754,N_49840);
and UO_3760 (O_3760,N_49789,N_49792);
and UO_3761 (O_3761,N_49812,N_49952);
nor UO_3762 (O_3762,N_49907,N_49915);
and UO_3763 (O_3763,N_49847,N_49957);
nand UO_3764 (O_3764,N_49973,N_49950);
or UO_3765 (O_3765,N_49762,N_49848);
or UO_3766 (O_3766,N_49910,N_49967);
nor UO_3767 (O_3767,N_49849,N_49754);
xnor UO_3768 (O_3768,N_49955,N_49970);
and UO_3769 (O_3769,N_49947,N_49770);
nand UO_3770 (O_3770,N_49760,N_49770);
and UO_3771 (O_3771,N_49905,N_49811);
and UO_3772 (O_3772,N_49818,N_49773);
nor UO_3773 (O_3773,N_49898,N_49868);
nor UO_3774 (O_3774,N_49874,N_49823);
nor UO_3775 (O_3775,N_49884,N_49877);
nor UO_3776 (O_3776,N_49985,N_49825);
nand UO_3777 (O_3777,N_49854,N_49940);
nor UO_3778 (O_3778,N_49916,N_49795);
and UO_3779 (O_3779,N_49794,N_49795);
or UO_3780 (O_3780,N_49778,N_49821);
nand UO_3781 (O_3781,N_49931,N_49834);
and UO_3782 (O_3782,N_49806,N_49904);
or UO_3783 (O_3783,N_49788,N_49778);
and UO_3784 (O_3784,N_49869,N_49782);
and UO_3785 (O_3785,N_49900,N_49968);
xor UO_3786 (O_3786,N_49784,N_49905);
or UO_3787 (O_3787,N_49811,N_49824);
nand UO_3788 (O_3788,N_49823,N_49835);
xnor UO_3789 (O_3789,N_49773,N_49776);
xor UO_3790 (O_3790,N_49756,N_49994);
nor UO_3791 (O_3791,N_49972,N_49846);
xnor UO_3792 (O_3792,N_49820,N_49922);
and UO_3793 (O_3793,N_49915,N_49833);
or UO_3794 (O_3794,N_49890,N_49820);
nand UO_3795 (O_3795,N_49822,N_49909);
nor UO_3796 (O_3796,N_49913,N_49948);
and UO_3797 (O_3797,N_49822,N_49895);
and UO_3798 (O_3798,N_49935,N_49794);
xor UO_3799 (O_3799,N_49976,N_49929);
nand UO_3800 (O_3800,N_49844,N_49846);
nand UO_3801 (O_3801,N_49792,N_49895);
xnor UO_3802 (O_3802,N_49846,N_49918);
and UO_3803 (O_3803,N_49947,N_49866);
and UO_3804 (O_3804,N_49874,N_49953);
nor UO_3805 (O_3805,N_49772,N_49886);
or UO_3806 (O_3806,N_49823,N_49775);
nor UO_3807 (O_3807,N_49893,N_49953);
nand UO_3808 (O_3808,N_49821,N_49920);
nand UO_3809 (O_3809,N_49910,N_49946);
nand UO_3810 (O_3810,N_49936,N_49983);
xnor UO_3811 (O_3811,N_49897,N_49846);
nand UO_3812 (O_3812,N_49989,N_49821);
or UO_3813 (O_3813,N_49992,N_49875);
and UO_3814 (O_3814,N_49927,N_49831);
or UO_3815 (O_3815,N_49895,N_49892);
nor UO_3816 (O_3816,N_49956,N_49784);
xnor UO_3817 (O_3817,N_49915,N_49815);
or UO_3818 (O_3818,N_49883,N_49916);
xor UO_3819 (O_3819,N_49802,N_49761);
nor UO_3820 (O_3820,N_49820,N_49931);
nand UO_3821 (O_3821,N_49957,N_49920);
nor UO_3822 (O_3822,N_49973,N_49791);
and UO_3823 (O_3823,N_49982,N_49850);
nor UO_3824 (O_3824,N_49878,N_49900);
nand UO_3825 (O_3825,N_49864,N_49962);
xor UO_3826 (O_3826,N_49844,N_49848);
nor UO_3827 (O_3827,N_49777,N_49931);
xnor UO_3828 (O_3828,N_49905,N_49751);
and UO_3829 (O_3829,N_49982,N_49784);
and UO_3830 (O_3830,N_49952,N_49861);
nand UO_3831 (O_3831,N_49936,N_49909);
nor UO_3832 (O_3832,N_49929,N_49800);
nand UO_3833 (O_3833,N_49976,N_49876);
xnor UO_3834 (O_3834,N_49986,N_49909);
or UO_3835 (O_3835,N_49819,N_49924);
or UO_3836 (O_3836,N_49901,N_49894);
and UO_3837 (O_3837,N_49855,N_49770);
and UO_3838 (O_3838,N_49962,N_49946);
xnor UO_3839 (O_3839,N_49872,N_49816);
nand UO_3840 (O_3840,N_49867,N_49942);
and UO_3841 (O_3841,N_49817,N_49887);
xnor UO_3842 (O_3842,N_49798,N_49889);
nor UO_3843 (O_3843,N_49902,N_49864);
nand UO_3844 (O_3844,N_49983,N_49811);
nor UO_3845 (O_3845,N_49962,N_49758);
and UO_3846 (O_3846,N_49994,N_49938);
nand UO_3847 (O_3847,N_49874,N_49973);
and UO_3848 (O_3848,N_49900,N_49967);
xnor UO_3849 (O_3849,N_49981,N_49861);
or UO_3850 (O_3850,N_49877,N_49937);
or UO_3851 (O_3851,N_49830,N_49911);
nor UO_3852 (O_3852,N_49911,N_49763);
or UO_3853 (O_3853,N_49937,N_49922);
nor UO_3854 (O_3854,N_49885,N_49915);
and UO_3855 (O_3855,N_49977,N_49938);
and UO_3856 (O_3856,N_49858,N_49825);
or UO_3857 (O_3857,N_49947,N_49952);
nand UO_3858 (O_3858,N_49824,N_49997);
xnor UO_3859 (O_3859,N_49790,N_49967);
xnor UO_3860 (O_3860,N_49813,N_49973);
and UO_3861 (O_3861,N_49829,N_49871);
nand UO_3862 (O_3862,N_49816,N_49918);
xor UO_3863 (O_3863,N_49927,N_49931);
nand UO_3864 (O_3864,N_49798,N_49808);
and UO_3865 (O_3865,N_49863,N_49808);
xor UO_3866 (O_3866,N_49914,N_49915);
or UO_3867 (O_3867,N_49941,N_49842);
or UO_3868 (O_3868,N_49892,N_49936);
and UO_3869 (O_3869,N_49865,N_49942);
and UO_3870 (O_3870,N_49968,N_49772);
xnor UO_3871 (O_3871,N_49798,N_49928);
xor UO_3872 (O_3872,N_49911,N_49772);
nand UO_3873 (O_3873,N_49790,N_49857);
xnor UO_3874 (O_3874,N_49861,N_49893);
and UO_3875 (O_3875,N_49845,N_49993);
xor UO_3876 (O_3876,N_49763,N_49907);
and UO_3877 (O_3877,N_49988,N_49982);
and UO_3878 (O_3878,N_49895,N_49972);
or UO_3879 (O_3879,N_49824,N_49866);
xor UO_3880 (O_3880,N_49869,N_49961);
and UO_3881 (O_3881,N_49932,N_49913);
xor UO_3882 (O_3882,N_49863,N_49825);
or UO_3883 (O_3883,N_49840,N_49936);
xor UO_3884 (O_3884,N_49961,N_49912);
nor UO_3885 (O_3885,N_49908,N_49936);
and UO_3886 (O_3886,N_49986,N_49904);
or UO_3887 (O_3887,N_49776,N_49825);
nand UO_3888 (O_3888,N_49849,N_49993);
nand UO_3889 (O_3889,N_49982,N_49950);
and UO_3890 (O_3890,N_49943,N_49952);
nand UO_3891 (O_3891,N_49900,N_49997);
nor UO_3892 (O_3892,N_49787,N_49811);
and UO_3893 (O_3893,N_49929,N_49842);
and UO_3894 (O_3894,N_49917,N_49924);
or UO_3895 (O_3895,N_49763,N_49974);
xor UO_3896 (O_3896,N_49773,N_49822);
xor UO_3897 (O_3897,N_49892,N_49894);
xnor UO_3898 (O_3898,N_49949,N_49997);
or UO_3899 (O_3899,N_49812,N_49996);
and UO_3900 (O_3900,N_49960,N_49899);
nand UO_3901 (O_3901,N_49972,N_49829);
nor UO_3902 (O_3902,N_49814,N_49785);
and UO_3903 (O_3903,N_49767,N_49959);
and UO_3904 (O_3904,N_49898,N_49803);
and UO_3905 (O_3905,N_49805,N_49773);
nand UO_3906 (O_3906,N_49885,N_49935);
xnor UO_3907 (O_3907,N_49809,N_49751);
nor UO_3908 (O_3908,N_49977,N_49811);
nand UO_3909 (O_3909,N_49999,N_49864);
nor UO_3910 (O_3910,N_49771,N_49751);
or UO_3911 (O_3911,N_49795,N_49858);
or UO_3912 (O_3912,N_49913,N_49851);
or UO_3913 (O_3913,N_49960,N_49909);
and UO_3914 (O_3914,N_49882,N_49895);
xor UO_3915 (O_3915,N_49837,N_49845);
nand UO_3916 (O_3916,N_49809,N_49932);
nand UO_3917 (O_3917,N_49871,N_49930);
xnor UO_3918 (O_3918,N_49989,N_49937);
or UO_3919 (O_3919,N_49800,N_49822);
nand UO_3920 (O_3920,N_49973,N_49939);
and UO_3921 (O_3921,N_49810,N_49859);
nor UO_3922 (O_3922,N_49990,N_49815);
and UO_3923 (O_3923,N_49907,N_49792);
and UO_3924 (O_3924,N_49762,N_49828);
nand UO_3925 (O_3925,N_49974,N_49953);
xor UO_3926 (O_3926,N_49906,N_49936);
nor UO_3927 (O_3927,N_49906,N_49760);
xnor UO_3928 (O_3928,N_49946,N_49911);
and UO_3929 (O_3929,N_49911,N_49883);
xnor UO_3930 (O_3930,N_49920,N_49875);
or UO_3931 (O_3931,N_49838,N_49868);
xor UO_3932 (O_3932,N_49941,N_49981);
or UO_3933 (O_3933,N_49916,N_49911);
and UO_3934 (O_3934,N_49993,N_49856);
xnor UO_3935 (O_3935,N_49967,N_49876);
and UO_3936 (O_3936,N_49832,N_49830);
and UO_3937 (O_3937,N_49976,N_49999);
nor UO_3938 (O_3938,N_49881,N_49893);
or UO_3939 (O_3939,N_49864,N_49976);
and UO_3940 (O_3940,N_49979,N_49880);
and UO_3941 (O_3941,N_49948,N_49813);
xnor UO_3942 (O_3942,N_49840,N_49994);
nor UO_3943 (O_3943,N_49834,N_49884);
nor UO_3944 (O_3944,N_49797,N_49833);
or UO_3945 (O_3945,N_49857,N_49787);
nand UO_3946 (O_3946,N_49802,N_49902);
or UO_3947 (O_3947,N_49841,N_49854);
nor UO_3948 (O_3948,N_49801,N_49914);
and UO_3949 (O_3949,N_49769,N_49807);
or UO_3950 (O_3950,N_49910,N_49857);
xnor UO_3951 (O_3951,N_49797,N_49869);
or UO_3952 (O_3952,N_49780,N_49866);
nand UO_3953 (O_3953,N_49973,N_49779);
nor UO_3954 (O_3954,N_49929,N_49777);
or UO_3955 (O_3955,N_49940,N_49860);
or UO_3956 (O_3956,N_49917,N_49755);
and UO_3957 (O_3957,N_49916,N_49877);
nor UO_3958 (O_3958,N_49844,N_49992);
and UO_3959 (O_3959,N_49916,N_49798);
or UO_3960 (O_3960,N_49809,N_49972);
nand UO_3961 (O_3961,N_49798,N_49999);
or UO_3962 (O_3962,N_49883,N_49843);
xor UO_3963 (O_3963,N_49885,N_49989);
nand UO_3964 (O_3964,N_49870,N_49963);
or UO_3965 (O_3965,N_49792,N_49970);
or UO_3966 (O_3966,N_49897,N_49855);
xnor UO_3967 (O_3967,N_49974,N_49959);
xnor UO_3968 (O_3968,N_49914,N_49910);
xor UO_3969 (O_3969,N_49919,N_49998);
or UO_3970 (O_3970,N_49956,N_49843);
or UO_3971 (O_3971,N_49971,N_49848);
nor UO_3972 (O_3972,N_49801,N_49759);
and UO_3973 (O_3973,N_49794,N_49857);
xnor UO_3974 (O_3974,N_49880,N_49877);
xor UO_3975 (O_3975,N_49860,N_49938);
nand UO_3976 (O_3976,N_49781,N_49882);
nor UO_3977 (O_3977,N_49997,N_49872);
nor UO_3978 (O_3978,N_49980,N_49758);
xnor UO_3979 (O_3979,N_49969,N_49807);
nand UO_3980 (O_3980,N_49916,N_49913);
xnor UO_3981 (O_3981,N_49806,N_49911);
nor UO_3982 (O_3982,N_49844,N_49877);
nand UO_3983 (O_3983,N_49972,N_49960);
xnor UO_3984 (O_3984,N_49867,N_49959);
nand UO_3985 (O_3985,N_49797,N_49876);
xor UO_3986 (O_3986,N_49830,N_49953);
nand UO_3987 (O_3987,N_49954,N_49975);
nor UO_3988 (O_3988,N_49828,N_49878);
xnor UO_3989 (O_3989,N_49830,N_49848);
nor UO_3990 (O_3990,N_49859,N_49855);
and UO_3991 (O_3991,N_49820,N_49967);
or UO_3992 (O_3992,N_49825,N_49805);
xnor UO_3993 (O_3993,N_49762,N_49829);
and UO_3994 (O_3994,N_49990,N_49906);
nor UO_3995 (O_3995,N_49758,N_49762);
nand UO_3996 (O_3996,N_49826,N_49790);
or UO_3997 (O_3997,N_49977,N_49907);
nor UO_3998 (O_3998,N_49924,N_49877);
xnor UO_3999 (O_3999,N_49842,N_49965);
or UO_4000 (O_4000,N_49914,N_49918);
nand UO_4001 (O_4001,N_49794,N_49875);
xnor UO_4002 (O_4002,N_49784,N_49995);
nand UO_4003 (O_4003,N_49878,N_49779);
or UO_4004 (O_4004,N_49766,N_49941);
nand UO_4005 (O_4005,N_49838,N_49856);
or UO_4006 (O_4006,N_49977,N_49774);
nand UO_4007 (O_4007,N_49952,N_49756);
nand UO_4008 (O_4008,N_49901,N_49752);
nor UO_4009 (O_4009,N_49769,N_49864);
or UO_4010 (O_4010,N_49881,N_49789);
nand UO_4011 (O_4011,N_49829,N_49947);
and UO_4012 (O_4012,N_49909,N_49777);
nand UO_4013 (O_4013,N_49782,N_49983);
nand UO_4014 (O_4014,N_49988,N_49938);
xnor UO_4015 (O_4015,N_49790,N_49973);
nor UO_4016 (O_4016,N_49862,N_49999);
xor UO_4017 (O_4017,N_49932,N_49820);
or UO_4018 (O_4018,N_49757,N_49960);
nand UO_4019 (O_4019,N_49856,N_49986);
or UO_4020 (O_4020,N_49987,N_49850);
and UO_4021 (O_4021,N_49845,N_49820);
and UO_4022 (O_4022,N_49999,N_49952);
xnor UO_4023 (O_4023,N_49847,N_49799);
nor UO_4024 (O_4024,N_49996,N_49991);
or UO_4025 (O_4025,N_49980,N_49973);
nand UO_4026 (O_4026,N_49897,N_49858);
nor UO_4027 (O_4027,N_49929,N_49918);
or UO_4028 (O_4028,N_49925,N_49755);
and UO_4029 (O_4029,N_49915,N_49794);
xnor UO_4030 (O_4030,N_49827,N_49960);
nand UO_4031 (O_4031,N_49890,N_49897);
xor UO_4032 (O_4032,N_49923,N_49866);
nand UO_4033 (O_4033,N_49935,N_49788);
nand UO_4034 (O_4034,N_49776,N_49917);
xor UO_4035 (O_4035,N_49757,N_49892);
xnor UO_4036 (O_4036,N_49961,N_49828);
or UO_4037 (O_4037,N_49847,N_49933);
nand UO_4038 (O_4038,N_49872,N_49780);
or UO_4039 (O_4039,N_49764,N_49868);
and UO_4040 (O_4040,N_49830,N_49882);
nand UO_4041 (O_4041,N_49810,N_49775);
or UO_4042 (O_4042,N_49875,N_49836);
nand UO_4043 (O_4043,N_49869,N_49925);
nand UO_4044 (O_4044,N_49774,N_49853);
xor UO_4045 (O_4045,N_49994,N_49992);
and UO_4046 (O_4046,N_49901,N_49759);
xnor UO_4047 (O_4047,N_49956,N_49780);
or UO_4048 (O_4048,N_49932,N_49955);
xnor UO_4049 (O_4049,N_49818,N_49947);
nor UO_4050 (O_4050,N_49863,N_49966);
and UO_4051 (O_4051,N_49857,N_49967);
and UO_4052 (O_4052,N_49769,N_49880);
or UO_4053 (O_4053,N_49813,N_49905);
and UO_4054 (O_4054,N_49758,N_49972);
nand UO_4055 (O_4055,N_49764,N_49877);
nand UO_4056 (O_4056,N_49918,N_49973);
or UO_4057 (O_4057,N_49943,N_49853);
or UO_4058 (O_4058,N_49796,N_49951);
xnor UO_4059 (O_4059,N_49900,N_49946);
nand UO_4060 (O_4060,N_49911,N_49917);
and UO_4061 (O_4061,N_49821,N_49800);
nor UO_4062 (O_4062,N_49774,N_49949);
or UO_4063 (O_4063,N_49891,N_49783);
and UO_4064 (O_4064,N_49987,N_49784);
nand UO_4065 (O_4065,N_49774,N_49821);
xnor UO_4066 (O_4066,N_49867,N_49946);
or UO_4067 (O_4067,N_49814,N_49958);
xnor UO_4068 (O_4068,N_49873,N_49844);
or UO_4069 (O_4069,N_49857,N_49926);
or UO_4070 (O_4070,N_49785,N_49875);
xnor UO_4071 (O_4071,N_49753,N_49895);
xor UO_4072 (O_4072,N_49914,N_49782);
xnor UO_4073 (O_4073,N_49802,N_49947);
xor UO_4074 (O_4074,N_49773,N_49750);
and UO_4075 (O_4075,N_49750,N_49977);
xor UO_4076 (O_4076,N_49866,N_49922);
and UO_4077 (O_4077,N_49790,N_49965);
nand UO_4078 (O_4078,N_49875,N_49995);
nand UO_4079 (O_4079,N_49930,N_49818);
and UO_4080 (O_4080,N_49941,N_49959);
nand UO_4081 (O_4081,N_49788,N_49780);
and UO_4082 (O_4082,N_49914,N_49939);
xnor UO_4083 (O_4083,N_49753,N_49837);
nand UO_4084 (O_4084,N_49886,N_49863);
and UO_4085 (O_4085,N_49838,N_49917);
nor UO_4086 (O_4086,N_49832,N_49981);
nand UO_4087 (O_4087,N_49980,N_49951);
nand UO_4088 (O_4088,N_49964,N_49751);
nor UO_4089 (O_4089,N_49822,N_49935);
or UO_4090 (O_4090,N_49982,N_49961);
xnor UO_4091 (O_4091,N_49932,N_49806);
xor UO_4092 (O_4092,N_49977,N_49856);
nand UO_4093 (O_4093,N_49872,N_49789);
nand UO_4094 (O_4094,N_49800,N_49814);
nor UO_4095 (O_4095,N_49810,N_49984);
nand UO_4096 (O_4096,N_49927,N_49855);
nor UO_4097 (O_4097,N_49999,N_49936);
or UO_4098 (O_4098,N_49906,N_49933);
nor UO_4099 (O_4099,N_49761,N_49860);
or UO_4100 (O_4100,N_49882,N_49890);
nand UO_4101 (O_4101,N_49754,N_49832);
nor UO_4102 (O_4102,N_49790,N_49878);
nand UO_4103 (O_4103,N_49794,N_49755);
or UO_4104 (O_4104,N_49842,N_49811);
nor UO_4105 (O_4105,N_49900,N_49842);
nor UO_4106 (O_4106,N_49774,N_49944);
and UO_4107 (O_4107,N_49800,N_49903);
nor UO_4108 (O_4108,N_49891,N_49842);
nand UO_4109 (O_4109,N_49758,N_49790);
xnor UO_4110 (O_4110,N_49898,N_49958);
and UO_4111 (O_4111,N_49990,N_49989);
nand UO_4112 (O_4112,N_49943,N_49980);
and UO_4113 (O_4113,N_49769,N_49794);
xnor UO_4114 (O_4114,N_49838,N_49772);
xnor UO_4115 (O_4115,N_49830,N_49870);
xor UO_4116 (O_4116,N_49908,N_49917);
and UO_4117 (O_4117,N_49937,N_49991);
and UO_4118 (O_4118,N_49832,N_49766);
nor UO_4119 (O_4119,N_49924,N_49860);
or UO_4120 (O_4120,N_49997,N_49820);
nor UO_4121 (O_4121,N_49822,N_49930);
nand UO_4122 (O_4122,N_49961,N_49884);
nor UO_4123 (O_4123,N_49979,N_49925);
nor UO_4124 (O_4124,N_49944,N_49796);
and UO_4125 (O_4125,N_49921,N_49831);
and UO_4126 (O_4126,N_49877,N_49817);
xor UO_4127 (O_4127,N_49834,N_49752);
and UO_4128 (O_4128,N_49987,N_49823);
xnor UO_4129 (O_4129,N_49827,N_49865);
xnor UO_4130 (O_4130,N_49860,N_49772);
nand UO_4131 (O_4131,N_49947,N_49963);
nor UO_4132 (O_4132,N_49922,N_49887);
or UO_4133 (O_4133,N_49884,N_49953);
or UO_4134 (O_4134,N_49855,N_49963);
nor UO_4135 (O_4135,N_49872,N_49766);
nand UO_4136 (O_4136,N_49818,N_49862);
nor UO_4137 (O_4137,N_49909,N_49800);
nor UO_4138 (O_4138,N_49753,N_49948);
nor UO_4139 (O_4139,N_49847,N_49884);
nor UO_4140 (O_4140,N_49945,N_49773);
xor UO_4141 (O_4141,N_49913,N_49968);
nand UO_4142 (O_4142,N_49969,N_49933);
xnor UO_4143 (O_4143,N_49992,N_49895);
nor UO_4144 (O_4144,N_49993,N_49806);
nand UO_4145 (O_4145,N_49862,N_49756);
nor UO_4146 (O_4146,N_49921,N_49880);
xnor UO_4147 (O_4147,N_49987,N_49940);
xor UO_4148 (O_4148,N_49954,N_49981);
or UO_4149 (O_4149,N_49974,N_49970);
and UO_4150 (O_4150,N_49780,N_49982);
and UO_4151 (O_4151,N_49984,N_49942);
nand UO_4152 (O_4152,N_49887,N_49963);
or UO_4153 (O_4153,N_49876,N_49885);
nand UO_4154 (O_4154,N_49972,N_49892);
or UO_4155 (O_4155,N_49956,N_49979);
xor UO_4156 (O_4156,N_49945,N_49779);
nor UO_4157 (O_4157,N_49962,N_49966);
nand UO_4158 (O_4158,N_49927,N_49811);
and UO_4159 (O_4159,N_49868,N_49960);
nand UO_4160 (O_4160,N_49942,N_49954);
and UO_4161 (O_4161,N_49980,N_49755);
or UO_4162 (O_4162,N_49966,N_49884);
nor UO_4163 (O_4163,N_49784,N_49843);
nand UO_4164 (O_4164,N_49955,N_49929);
and UO_4165 (O_4165,N_49763,N_49994);
nor UO_4166 (O_4166,N_49818,N_49759);
nand UO_4167 (O_4167,N_49982,N_49818);
nor UO_4168 (O_4168,N_49829,N_49791);
nor UO_4169 (O_4169,N_49844,N_49988);
nor UO_4170 (O_4170,N_49979,N_49908);
and UO_4171 (O_4171,N_49813,N_49925);
xor UO_4172 (O_4172,N_49987,N_49829);
nor UO_4173 (O_4173,N_49808,N_49954);
nor UO_4174 (O_4174,N_49813,N_49823);
nor UO_4175 (O_4175,N_49772,N_49976);
xnor UO_4176 (O_4176,N_49962,N_49948);
nor UO_4177 (O_4177,N_49883,N_49974);
xor UO_4178 (O_4178,N_49813,N_49964);
xor UO_4179 (O_4179,N_49830,N_49843);
nor UO_4180 (O_4180,N_49805,N_49859);
and UO_4181 (O_4181,N_49838,N_49758);
xor UO_4182 (O_4182,N_49802,N_49863);
xor UO_4183 (O_4183,N_49774,N_49868);
nand UO_4184 (O_4184,N_49776,N_49920);
or UO_4185 (O_4185,N_49904,N_49918);
and UO_4186 (O_4186,N_49880,N_49761);
and UO_4187 (O_4187,N_49794,N_49765);
and UO_4188 (O_4188,N_49920,N_49902);
nand UO_4189 (O_4189,N_49820,N_49979);
and UO_4190 (O_4190,N_49961,N_49890);
and UO_4191 (O_4191,N_49820,N_49982);
nor UO_4192 (O_4192,N_49804,N_49938);
nor UO_4193 (O_4193,N_49846,N_49862);
and UO_4194 (O_4194,N_49917,N_49912);
or UO_4195 (O_4195,N_49961,N_49758);
xor UO_4196 (O_4196,N_49924,N_49867);
nand UO_4197 (O_4197,N_49896,N_49916);
xor UO_4198 (O_4198,N_49809,N_49998);
nor UO_4199 (O_4199,N_49818,N_49946);
and UO_4200 (O_4200,N_49950,N_49910);
and UO_4201 (O_4201,N_49903,N_49945);
or UO_4202 (O_4202,N_49961,N_49889);
nand UO_4203 (O_4203,N_49971,N_49916);
nand UO_4204 (O_4204,N_49764,N_49861);
and UO_4205 (O_4205,N_49812,N_49971);
or UO_4206 (O_4206,N_49974,N_49906);
or UO_4207 (O_4207,N_49972,N_49821);
xnor UO_4208 (O_4208,N_49902,N_49957);
xor UO_4209 (O_4209,N_49816,N_49811);
or UO_4210 (O_4210,N_49915,N_49846);
or UO_4211 (O_4211,N_49932,N_49780);
or UO_4212 (O_4212,N_49941,N_49803);
nand UO_4213 (O_4213,N_49782,N_49828);
or UO_4214 (O_4214,N_49827,N_49792);
nor UO_4215 (O_4215,N_49972,N_49878);
nor UO_4216 (O_4216,N_49888,N_49857);
or UO_4217 (O_4217,N_49817,N_49788);
and UO_4218 (O_4218,N_49868,N_49935);
nand UO_4219 (O_4219,N_49910,N_49911);
and UO_4220 (O_4220,N_49859,N_49786);
xor UO_4221 (O_4221,N_49755,N_49930);
or UO_4222 (O_4222,N_49779,N_49948);
and UO_4223 (O_4223,N_49962,N_49874);
nand UO_4224 (O_4224,N_49967,N_49817);
and UO_4225 (O_4225,N_49886,N_49769);
nand UO_4226 (O_4226,N_49839,N_49828);
and UO_4227 (O_4227,N_49914,N_49819);
nand UO_4228 (O_4228,N_49865,N_49864);
and UO_4229 (O_4229,N_49967,N_49990);
nand UO_4230 (O_4230,N_49865,N_49968);
xnor UO_4231 (O_4231,N_49931,N_49990);
xnor UO_4232 (O_4232,N_49766,N_49887);
xor UO_4233 (O_4233,N_49752,N_49997);
nor UO_4234 (O_4234,N_49880,N_49963);
or UO_4235 (O_4235,N_49886,N_49787);
or UO_4236 (O_4236,N_49822,N_49925);
and UO_4237 (O_4237,N_49778,N_49789);
or UO_4238 (O_4238,N_49969,N_49816);
and UO_4239 (O_4239,N_49888,N_49803);
or UO_4240 (O_4240,N_49959,N_49920);
and UO_4241 (O_4241,N_49937,N_49752);
xnor UO_4242 (O_4242,N_49937,N_49943);
or UO_4243 (O_4243,N_49875,N_49943);
or UO_4244 (O_4244,N_49856,N_49887);
nor UO_4245 (O_4245,N_49979,N_49784);
nand UO_4246 (O_4246,N_49956,N_49803);
nand UO_4247 (O_4247,N_49933,N_49806);
nor UO_4248 (O_4248,N_49892,N_49945);
and UO_4249 (O_4249,N_49900,N_49964);
or UO_4250 (O_4250,N_49836,N_49771);
or UO_4251 (O_4251,N_49968,N_49858);
xnor UO_4252 (O_4252,N_49779,N_49901);
nand UO_4253 (O_4253,N_49766,N_49966);
xor UO_4254 (O_4254,N_49989,N_49850);
or UO_4255 (O_4255,N_49871,N_49878);
xnor UO_4256 (O_4256,N_49857,N_49911);
xor UO_4257 (O_4257,N_49951,N_49911);
and UO_4258 (O_4258,N_49832,N_49763);
nor UO_4259 (O_4259,N_49831,N_49890);
and UO_4260 (O_4260,N_49832,N_49865);
xnor UO_4261 (O_4261,N_49831,N_49760);
xor UO_4262 (O_4262,N_49808,N_49950);
and UO_4263 (O_4263,N_49875,N_49756);
nand UO_4264 (O_4264,N_49900,N_49875);
xnor UO_4265 (O_4265,N_49804,N_49903);
xnor UO_4266 (O_4266,N_49980,N_49856);
nand UO_4267 (O_4267,N_49881,N_49878);
and UO_4268 (O_4268,N_49880,N_49852);
nand UO_4269 (O_4269,N_49762,N_49751);
nor UO_4270 (O_4270,N_49886,N_49917);
nor UO_4271 (O_4271,N_49792,N_49852);
nor UO_4272 (O_4272,N_49760,N_49830);
nand UO_4273 (O_4273,N_49973,N_49976);
xor UO_4274 (O_4274,N_49912,N_49948);
or UO_4275 (O_4275,N_49914,N_49807);
nand UO_4276 (O_4276,N_49866,N_49846);
nand UO_4277 (O_4277,N_49952,N_49752);
and UO_4278 (O_4278,N_49934,N_49791);
and UO_4279 (O_4279,N_49787,N_49988);
or UO_4280 (O_4280,N_49891,N_49762);
nor UO_4281 (O_4281,N_49787,N_49934);
and UO_4282 (O_4282,N_49760,N_49964);
xnor UO_4283 (O_4283,N_49912,N_49971);
nor UO_4284 (O_4284,N_49911,N_49773);
and UO_4285 (O_4285,N_49989,N_49910);
nor UO_4286 (O_4286,N_49915,N_49928);
nand UO_4287 (O_4287,N_49994,N_49986);
nand UO_4288 (O_4288,N_49765,N_49988);
nand UO_4289 (O_4289,N_49905,N_49834);
nor UO_4290 (O_4290,N_49895,N_49846);
xor UO_4291 (O_4291,N_49810,N_49850);
xnor UO_4292 (O_4292,N_49772,N_49805);
and UO_4293 (O_4293,N_49780,N_49991);
nand UO_4294 (O_4294,N_49925,N_49921);
nor UO_4295 (O_4295,N_49821,N_49806);
xnor UO_4296 (O_4296,N_49800,N_49915);
or UO_4297 (O_4297,N_49914,N_49927);
xnor UO_4298 (O_4298,N_49782,N_49941);
or UO_4299 (O_4299,N_49874,N_49757);
xor UO_4300 (O_4300,N_49824,N_49820);
nor UO_4301 (O_4301,N_49884,N_49896);
xor UO_4302 (O_4302,N_49903,N_49866);
and UO_4303 (O_4303,N_49799,N_49967);
or UO_4304 (O_4304,N_49801,N_49802);
and UO_4305 (O_4305,N_49823,N_49931);
or UO_4306 (O_4306,N_49821,N_49904);
nor UO_4307 (O_4307,N_49826,N_49758);
xor UO_4308 (O_4308,N_49786,N_49942);
xnor UO_4309 (O_4309,N_49885,N_49836);
nand UO_4310 (O_4310,N_49864,N_49956);
nor UO_4311 (O_4311,N_49815,N_49947);
or UO_4312 (O_4312,N_49895,N_49826);
nor UO_4313 (O_4313,N_49847,N_49952);
and UO_4314 (O_4314,N_49908,N_49856);
xor UO_4315 (O_4315,N_49829,N_49993);
nand UO_4316 (O_4316,N_49982,N_49789);
xor UO_4317 (O_4317,N_49921,N_49841);
nand UO_4318 (O_4318,N_49974,N_49917);
xnor UO_4319 (O_4319,N_49802,N_49966);
nand UO_4320 (O_4320,N_49989,N_49801);
nor UO_4321 (O_4321,N_49754,N_49850);
xor UO_4322 (O_4322,N_49981,N_49810);
or UO_4323 (O_4323,N_49949,N_49781);
and UO_4324 (O_4324,N_49846,N_49790);
or UO_4325 (O_4325,N_49802,N_49852);
and UO_4326 (O_4326,N_49858,N_49943);
nor UO_4327 (O_4327,N_49772,N_49823);
or UO_4328 (O_4328,N_49825,N_49856);
nor UO_4329 (O_4329,N_49810,N_49883);
nand UO_4330 (O_4330,N_49854,N_49928);
xnor UO_4331 (O_4331,N_49793,N_49953);
xnor UO_4332 (O_4332,N_49905,N_49788);
or UO_4333 (O_4333,N_49975,N_49999);
nand UO_4334 (O_4334,N_49992,N_49900);
and UO_4335 (O_4335,N_49795,N_49782);
or UO_4336 (O_4336,N_49781,N_49961);
nand UO_4337 (O_4337,N_49952,N_49892);
xor UO_4338 (O_4338,N_49994,N_49946);
nand UO_4339 (O_4339,N_49962,N_49816);
nor UO_4340 (O_4340,N_49808,N_49835);
nand UO_4341 (O_4341,N_49810,N_49846);
nor UO_4342 (O_4342,N_49832,N_49980);
or UO_4343 (O_4343,N_49938,N_49762);
or UO_4344 (O_4344,N_49795,N_49937);
or UO_4345 (O_4345,N_49876,N_49891);
or UO_4346 (O_4346,N_49877,N_49805);
or UO_4347 (O_4347,N_49883,N_49768);
nor UO_4348 (O_4348,N_49822,N_49926);
and UO_4349 (O_4349,N_49946,N_49852);
nor UO_4350 (O_4350,N_49981,N_49752);
nor UO_4351 (O_4351,N_49793,N_49905);
nand UO_4352 (O_4352,N_49818,N_49882);
nand UO_4353 (O_4353,N_49995,N_49835);
and UO_4354 (O_4354,N_49827,N_49839);
or UO_4355 (O_4355,N_49966,N_49915);
nand UO_4356 (O_4356,N_49908,N_49849);
xnor UO_4357 (O_4357,N_49854,N_49777);
xor UO_4358 (O_4358,N_49777,N_49946);
nand UO_4359 (O_4359,N_49905,N_49874);
nor UO_4360 (O_4360,N_49857,N_49985);
nand UO_4361 (O_4361,N_49765,N_49889);
nor UO_4362 (O_4362,N_49800,N_49834);
nand UO_4363 (O_4363,N_49839,N_49948);
or UO_4364 (O_4364,N_49959,N_49893);
xnor UO_4365 (O_4365,N_49901,N_49763);
nand UO_4366 (O_4366,N_49961,N_49908);
nor UO_4367 (O_4367,N_49939,N_49988);
or UO_4368 (O_4368,N_49794,N_49774);
xnor UO_4369 (O_4369,N_49934,N_49762);
nand UO_4370 (O_4370,N_49869,N_49851);
xor UO_4371 (O_4371,N_49990,N_49963);
xor UO_4372 (O_4372,N_49820,N_49770);
nor UO_4373 (O_4373,N_49778,N_49777);
xnor UO_4374 (O_4374,N_49786,N_49836);
and UO_4375 (O_4375,N_49780,N_49846);
nand UO_4376 (O_4376,N_49984,N_49927);
xor UO_4377 (O_4377,N_49824,N_49818);
and UO_4378 (O_4378,N_49990,N_49975);
and UO_4379 (O_4379,N_49811,N_49973);
xor UO_4380 (O_4380,N_49928,N_49848);
and UO_4381 (O_4381,N_49872,N_49752);
and UO_4382 (O_4382,N_49985,N_49957);
and UO_4383 (O_4383,N_49771,N_49937);
nand UO_4384 (O_4384,N_49960,N_49968);
nor UO_4385 (O_4385,N_49859,N_49893);
nor UO_4386 (O_4386,N_49857,N_49938);
and UO_4387 (O_4387,N_49766,N_49984);
nor UO_4388 (O_4388,N_49943,N_49839);
xnor UO_4389 (O_4389,N_49876,N_49923);
nor UO_4390 (O_4390,N_49906,N_49836);
or UO_4391 (O_4391,N_49756,N_49828);
xnor UO_4392 (O_4392,N_49923,N_49948);
xnor UO_4393 (O_4393,N_49880,N_49970);
and UO_4394 (O_4394,N_49834,N_49791);
or UO_4395 (O_4395,N_49986,N_49855);
xnor UO_4396 (O_4396,N_49860,N_49900);
nand UO_4397 (O_4397,N_49858,N_49805);
and UO_4398 (O_4398,N_49954,N_49915);
xor UO_4399 (O_4399,N_49859,N_49803);
xor UO_4400 (O_4400,N_49800,N_49901);
xor UO_4401 (O_4401,N_49959,N_49971);
xor UO_4402 (O_4402,N_49821,N_49808);
nand UO_4403 (O_4403,N_49808,N_49873);
nor UO_4404 (O_4404,N_49871,N_49779);
xnor UO_4405 (O_4405,N_49957,N_49803);
nor UO_4406 (O_4406,N_49863,N_49857);
and UO_4407 (O_4407,N_49915,N_49999);
and UO_4408 (O_4408,N_49877,N_49828);
and UO_4409 (O_4409,N_49751,N_49958);
or UO_4410 (O_4410,N_49879,N_49935);
and UO_4411 (O_4411,N_49796,N_49897);
xnor UO_4412 (O_4412,N_49821,N_49836);
and UO_4413 (O_4413,N_49804,N_49916);
or UO_4414 (O_4414,N_49942,N_49792);
xnor UO_4415 (O_4415,N_49930,N_49776);
and UO_4416 (O_4416,N_49775,N_49868);
xnor UO_4417 (O_4417,N_49840,N_49812);
and UO_4418 (O_4418,N_49943,N_49983);
nand UO_4419 (O_4419,N_49862,N_49913);
nand UO_4420 (O_4420,N_49812,N_49813);
nand UO_4421 (O_4421,N_49946,N_49836);
and UO_4422 (O_4422,N_49842,N_49808);
or UO_4423 (O_4423,N_49791,N_49819);
nand UO_4424 (O_4424,N_49898,N_49811);
nand UO_4425 (O_4425,N_49872,N_49793);
xnor UO_4426 (O_4426,N_49970,N_49913);
xnor UO_4427 (O_4427,N_49790,N_49911);
and UO_4428 (O_4428,N_49913,N_49878);
or UO_4429 (O_4429,N_49876,N_49906);
and UO_4430 (O_4430,N_49971,N_49862);
nand UO_4431 (O_4431,N_49867,N_49768);
nor UO_4432 (O_4432,N_49867,N_49980);
xnor UO_4433 (O_4433,N_49871,N_49911);
and UO_4434 (O_4434,N_49784,N_49925);
nor UO_4435 (O_4435,N_49870,N_49827);
or UO_4436 (O_4436,N_49822,N_49900);
and UO_4437 (O_4437,N_49960,N_49783);
xor UO_4438 (O_4438,N_49919,N_49771);
xor UO_4439 (O_4439,N_49839,N_49799);
and UO_4440 (O_4440,N_49895,N_49829);
nor UO_4441 (O_4441,N_49854,N_49969);
nor UO_4442 (O_4442,N_49982,N_49857);
or UO_4443 (O_4443,N_49841,N_49849);
or UO_4444 (O_4444,N_49851,N_49967);
and UO_4445 (O_4445,N_49913,N_49918);
nor UO_4446 (O_4446,N_49775,N_49853);
and UO_4447 (O_4447,N_49952,N_49964);
nor UO_4448 (O_4448,N_49949,N_49768);
and UO_4449 (O_4449,N_49767,N_49983);
nand UO_4450 (O_4450,N_49792,N_49810);
or UO_4451 (O_4451,N_49900,N_49754);
xor UO_4452 (O_4452,N_49835,N_49942);
nand UO_4453 (O_4453,N_49857,N_49776);
and UO_4454 (O_4454,N_49882,N_49850);
and UO_4455 (O_4455,N_49978,N_49793);
xor UO_4456 (O_4456,N_49758,N_49904);
nand UO_4457 (O_4457,N_49806,N_49793);
or UO_4458 (O_4458,N_49774,N_49889);
nand UO_4459 (O_4459,N_49804,N_49919);
or UO_4460 (O_4460,N_49901,N_49764);
nand UO_4461 (O_4461,N_49797,N_49967);
xor UO_4462 (O_4462,N_49848,N_49797);
and UO_4463 (O_4463,N_49927,N_49885);
nand UO_4464 (O_4464,N_49858,N_49941);
nand UO_4465 (O_4465,N_49936,N_49783);
or UO_4466 (O_4466,N_49807,N_49866);
xor UO_4467 (O_4467,N_49773,N_49823);
nand UO_4468 (O_4468,N_49935,N_49855);
and UO_4469 (O_4469,N_49872,N_49906);
nand UO_4470 (O_4470,N_49867,N_49999);
xor UO_4471 (O_4471,N_49760,N_49949);
nand UO_4472 (O_4472,N_49891,N_49965);
nor UO_4473 (O_4473,N_49957,N_49759);
or UO_4474 (O_4474,N_49758,N_49863);
and UO_4475 (O_4475,N_49819,N_49949);
xor UO_4476 (O_4476,N_49958,N_49980);
and UO_4477 (O_4477,N_49878,N_49771);
or UO_4478 (O_4478,N_49873,N_49945);
xnor UO_4479 (O_4479,N_49793,N_49928);
and UO_4480 (O_4480,N_49818,N_49984);
or UO_4481 (O_4481,N_49858,N_49925);
or UO_4482 (O_4482,N_49861,N_49815);
nor UO_4483 (O_4483,N_49760,N_49832);
or UO_4484 (O_4484,N_49776,N_49955);
nor UO_4485 (O_4485,N_49773,N_49934);
nor UO_4486 (O_4486,N_49919,N_49897);
nor UO_4487 (O_4487,N_49756,N_49833);
nand UO_4488 (O_4488,N_49754,N_49948);
nor UO_4489 (O_4489,N_49784,N_49819);
nor UO_4490 (O_4490,N_49784,N_49921);
nor UO_4491 (O_4491,N_49890,N_49801);
or UO_4492 (O_4492,N_49900,N_49789);
xnor UO_4493 (O_4493,N_49804,N_49820);
xor UO_4494 (O_4494,N_49939,N_49945);
xnor UO_4495 (O_4495,N_49888,N_49797);
nor UO_4496 (O_4496,N_49807,N_49857);
and UO_4497 (O_4497,N_49970,N_49824);
xnor UO_4498 (O_4498,N_49848,N_49847);
and UO_4499 (O_4499,N_49806,N_49857);
or UO_4500 (O_4500,N_49799,N_49979);
nand UO_4501 (O_4501,N_49769,N_49850);
nand UO_4502 (O_4502,N_49826,N_49890);
nor UO_4503 (O_4503,N_49938,N_49773);
nor UO_4504 (O_4504,N_49811,N_49971);
or UO_4505 (O_4505,N_49782,N_49780);
xor UO_4506 (O_4506,N_49964,N_49866);
and UO_4507 (O_4507,N_49874,N_49845);
nor UO_4508 (O_4508,N_49988,N_49757);
nor UO_4509 (O_4509,N_49873,N_49865);
and UO_4510 (O_4510,N_49887,N_49831);
or UO_4511 (O_4511,N_49983,N_49995);
or UO_4512 (O_4512,N_49957,N_49924);
nor UO_4513 (O_4513,N_49932,N_49842);
and UO_4514 (O_4514,N_49759,N_49965);
xnor UO_4515 (O_4515,N_49759,N_49897);
or UO_4516 (O_4516,N_49902,N_49861);
nand UO_4517 (O_4517,N_49988,N_49892);
or UO_4518 (O_4518,N_49791,N_49950);
or UO_4519 (O_4519,N_49810,N_49762);
xor UO_4520 (O_4520,N_49802,N_49930);
and UO_4521 (O_4521,N_49945,N_49801);
xnor UO_4522 (O_4522,N_49914,N_49764);
xnor UO_4523 (O_4523,N_49923,N_49893);
nor UO_4524 (O_4524,N_49880,N_49833);
nor UO_4525 (O_4525,N_49989,N_49911);
or UO_4526 (O_4526,N_49930,N_49856);
xnor UO_4527 (O_4527,N_49789,N_49828);
nor UO_4528 (O_4528,N_49758,N_49750);
or UO_4529 (O_4529,N_49882,N_49934);
xnor UO_4530 (O_4530,N_49923,N_49922);
and UO_4531 (O_4531,N_49973,N_49871);
and UO_4532 (O_4532,N_49838,N_49869);
xor UO_4533 (O_4533,N_49838,N_49880);
nand UO_4534 (O_4534,N_49781,N_49845);
nand UO_4535 (O_4535,N_49808,N_49828);
xnor UO_4536 (O_4536,N_49809,N_49853);
and UO_4537 (O_4537,N_49916,N_49927);
or UO_4538 (O_4538,N_49944,N_49908);
or UO_4539 (O_4539,N_49865,N_49978);
nand UO_4540 (O_4540,N_49853,N_49879);
nor UO_4541 (O_4541,N_49863,N_49861);
nand UO_4542 (O_4542,N_49898,N_49841);
xor UO_4543 (O_4543,N_49957,N_49779);
nor UO_4544 (O_4544,N_49805,N_49921);
and UO_4545 (O_4545,N_49872,N_49864);
nand UO_4546 (O_4546,N_49933,N_49896);
or UO_4547 (O_4547,N_49754,N_49970);
xor UO_4548 (O_4548,N_49856,N_49780);
nand UO_4549 (O_4549,N_49842,N_49821);
xnor UO_4550 (O_4550,N_49957,N_49986);
and UO_4551 (O_4551,N_49761,N_49974);
nor UO_4552 (O_4552,N_49818,N_49870);
xnor UO_4553 (O_4553,N_49977,N_49817);
xnor UO_4554 (O_4554,N_49902,N_49810);
and UO_4555 (O_4555,N_49870,N_49955);
nand UO_4556 (O_4556,N_49849,N_49792);
and UO_4557 (O_4557,N_49811,N_49765);
nand UO_4558 (O_4558,N_49817,N_49866);
nand UO_4559 (O_4559,N_49944,N_49926);
and UO_4560 (O_4560,N_49924,N_49973);
and UO_4561 (O_4561,N_49820,N_49759);
nand UO_4562 (O_4562,N_49858,N_49824);
nand UO_4563 (O_4563,N_49918,N_49831);
nand UO_4564 (O_4564,N_49940,N_49938);
xnor UO_4565 (O_4565,N_49778,N_49791);
nor UO_4566 (O_4566,N_49919,N_49766);
nand UO_4567 (O_4567,N_49892,N_49865);
nand UO_4568 (O_4568,N_49949,N_49787);
and UO_4569 (O_4569,N_49798,N_49959);
xor UO_4570 (O_4570,N_49997,N_49843);
nor UO_4571 (O_4571,N_49954,N_49947);
and UO_4572 (O_4572,N_49819,N_49889);
nor UO_4573 (O_4573,N_49929,N_49815);
or UO_4574 (O_4574,N_49817,N_49992);
xor UO_4575 (O_4575,N_49834,N_49928);
xnor UO_4576 (O_4576,N_49966,N_49982);
xor UO_4577 (O_4577,N_49763,N_49977);
nor UO_4578 (O_4578,N_49971,N_49882);
xnor UO_4579 (O_4579,N_49974,N_49881);
nand UO_4580 (O_4580,N_49927,N_49792);
and UO_4581 (O_4581,N_49829,N_49793);
nor UO_4582 (O_4582,N_49849,N_49855);
or UO_4583 (O_4583,N_49812,N_49975);
nand UO_4584 (O_4584,N_49777,N_49994);
nor UO_4585 (O_4585,N_49799,N_49972);
nand UO_4586 (O_4586,N_49910,N_49974);
xor UO_4587 (O_4587,N_49777,N_49995);
nand UO_4588 (O_4588,N_49857,N_49827);
nor UO_4589 (O_4589,N_49986,N_49791);
nor UO_4590 (O_4590,N_49804,N_49936);
xnor UO_4591 (O_4591,N_49969,N_49985);
and UO_4592 (O_4592,N_49802,N_49882);
and UO_4593 (O_4593,N_49870,N_49950);
xor UO_4594 (O_4594,N_49950,N_49814);
or UO_4595 (O_4595,N_49915,N_49835);
nand UO_4596 (O_4596,N_49840,N_49768);
or UO_4597 (O_4597,N_49901,N_49874);
nand UO_4598 (O_4598,N_49892,N_49801);
or UO_4599 (O_4599,N_49862,N_49911);
and UO_4600 (O_4600,N_49824,N_49850);
and UO_4601 (O_4601,N_49861,N_49864);
or UO_4602 (O_4602,N_49797,N_49851);
xnor UO_4603 (O_4603,N_49875,N_49849);
xnor UO_4604 (O_4604,N_49756,N_49906);
nor UO_4605 (O_4605,N_49831,N_49847);
nand UO_4606 (O_4606,N_49815,N_49750);
and UO_4607 (O_4607,N_49752,N_49790);
xnor UO_4608 (O_4608,N_49808,N_49925);
and UO_4609 (O_4609,N_49966,N_49956);
and UO_4610 (O_4610,N_49864,N_49949);
and UO_4611 (O_4611,N_49903,N_49902);
nor UO_4612 (O_4612,N_49979,N_49997);
xor UO_4613 (O_4613,N_49764,N_49980);
nand UO_4614 (O_4614,N_49963,N_49775);
nor UO_4615 (O_4615,N_49904,N_49935);
nor UO_4616 (O_4616,N_49943,N_49934);
and UO_4617 (O_4617,N_49938,N_49904);
nor UO_4618 (O_4618,N_49946,N_49783);
or UO_4619 (O_4619,N_49828,N_49848);
and UO_4620 (O_4620,N_49862,N_49839);
nand UO_4621 (O_4621,N_49777,N_49950);
and UO_4622 (O_4622,N_49831,N_49765);
or UO_4623 (O_4623,N_49783,N_49990);
nand UO_4624 (O_4624,N_49800,N_49979);
or UO_4625 (O_4625,N_49848,N_49887);
and UO_4626 (O_4626,N_49893,N_49983);
xor UO_4627 (O_4627,N_49908,N_49988);
or UO_4628 (O_4628,N_49930,N_49974);
nand UO_4629 (O_4629,N_49886,N_49875);
nand UO_4630 (O_4630,N_49972,N_49773);
or UO_4631 (O_4631,N_49925,N_49954);
and UO_4632 (O_4632,N_49766,N_49796);
nor UO_4633 (O_4633,N_49947,N_49967);
or UO_4634 (O_4634,N_49830,N_49797);
xor UO_4635 (O_4635,N_49890,N_49912);
and UO_4636 (O_4636,N_49987,N_49750);
xor UO_4637 (O_4637,N_49825,N_49787);
nand UO_4638 (O_4638,N_49945,N_49904);
and UO_4639 (O_4639,N_49895,N_49842);
xnor UO_4640 (O_4640,N_49843,N_49824);
and UO_4641 (O_4641,N_49983,N_49896);
nor UO_4642 (O_4642,N_49765,N_49952);
xor UO_4643 (O_4643,N_49893,N_49790);
or UO_4644 (O_4644,N_49752,N_49822);
and UO_4645 (O_4645,N_49835,N_49978);
or UO_4646 (O_4646,N_49751,N_49989);
nor UO_4647 (O_4647,N_49993,N_49838);
nor UO_4648 (O_4648,N_49752,N_49898);
xnor UO_4649 (O_4649,N_49962,N_49969);
or UO_4650 (O_4650,N_49853,N_49966);
xor UO_4651 (O_4651,N_49802,N_49994);
xor UO_4652 (O_4652,N_49982,N_49939);
xnor UO_4653 (O_4653,N_49762,N_49797);
and UO_4654 (O_4654,N_49828,N_49986);
xnor UO_4655 (O_4655,N_49891,N_49841);
xnor UO_4656 (O_4656,N_49887,N_49826);
xnor UO_4657 (O_4657,N_49918,N_49916);
nor UO_4658 (O_4658,N_49768,N_49771);
or UO_4659 (O_4659,N_49898,N_49883);
xnor UO_4660 (O_4660,N_49785,N_49973);
nor UO_4661 (O_4661,N_49962,N_49881);
xor UO_4662 (O_4662,N_49983,N_49944);
and UO_4663 (O_4663,N_49888,N_49951);
nor UO_4664 (O_4664,N_49806,N_49819);
and UO_4665 (O_4665,N_49985,N_49782);
nand UO_4666 (O_4666,N_49836,N_49959);
and UO_4667 (O_4667,N_49899,N_49877);
nand UO_4668 (O_4668,N_49887,N_49966);
or UO_4669 (O_4669,N_49810,N_49959);
xor UO_4670 (O_4670,N_49850,N_49981);
or UO_4671 (O_4671,N_49932,N_49929);
nand UO_4672 (O_4672,N_49988,N_49890);
nor UO_4673 (O_4673,N_49969,N_49955);
nor UO_4674 (O_4674,N_49814,N_49859);
or UO_4675 (O_4675,N_49932,N_49864);
xor UO_4676 (O_4676,N_49963,N_49801);
xor UO_4677 (O_4677,N_49809,N_49844);
and UO_4678 (O_4678,N_49790,N_49921);
nor UO_4679 (O_4679,N_49863,N_49822);
and UO_4680 (O_4680,N_49850,N_49777);
nor UO_4681 (O_4681,N_49946,N_49838);
xnor UO_4682 (O_4682,N_49816,N_49952);
nor UO_4683 (O_4683,N_49889,N_49904);
or UO_4684 (O_4684,N_49782,N_49826);
xnor UO_4685 (O_4685,N_49997,N_49962);
or UO_4686 (O_4686,N_49849,N_49778);
nor UO_4687 (O_4687,N_49987,N_49932);
and UO_4688 (O_4688,N_49931,N_49870);
or UO_4689 (O_4689,N_49924,N_49937);
or UO_4690 (O_4690,N_49778,N_49767);
or UO_4691 (O_4691,N_49894,N_49958);
nand UO_4692 (O_4692,N_49778,N_49900);
nor UO_4693 (O_4693,N_49794,N_49882);
nor UO_4694 (O_4694,N_49845,N_49750);
nand UO_4695 (O_4695,N_49881,N_49959);
nor UO_4696 (O_4696,N_49842,N_49794);
and UO_4697 (O_4697,N_49935,N_49802);
and UO_4698 (O_4698,N_49839,N_49973);
or UO_4699 (O_4699,N_49832,N_49847);
nand UO_4700 (O_4700,N_49900,N_49884);
or UO_4701 (O_4701,N_49986,N_49775);
xnor UO_4702 (O_4702,N_49756,N_49797);
nand UO_4703 (O_4703,N_49985,N_49934);
nand UO_4704 (O_4704,N_49946,N_49796);
nand UO_4705 (O_4705,N_49967,N_49859);
nor UO_4706 (O_4706,N_49833,N_49809);
or UO_4707 (O_4707,N_49935,N_49881);
or UO_4708 (O_4708,N_49896,N_49898);
xor UO_4709 (O_4709,N_49832,N_49888);
xnor UO_4710 (O_4710,N_49790,N_49776);
and UO_4711 (O_4711,N_49869,N_49984);
or UO_4712 (O_4712,N_49831,N_49804);
nand UO_4713 (O_4713,N_49933,N_49770);
or UO_4714 (O_4714,N_49911,N_49866);
or UO_4715 (O_4715,N_49864,N_49793);
xnor UO_4716 (O_4716,N_49772,N_49904);
nand UO_4717 (O_4717,N_49992,N_49903);
nand UO_4718 (O_4718,N_49880,N_49754);
xor UO_4719 (O_4719,N_49968,N_49980);
and UO_4720 (O_4720,N_49773,N_49917);
or UO_4721 (O_4721,N_49840,N_49822);
and UO_4722 (O_4722,N_49972,N_49957);
and UO_4723 (O_4723,N_49880,N_49941);
nand UO_4724 (O_4724,N_49891,N_49883);
nor UO_4725 (O_4725,N_49844,N_49866);
and UO_4726 (O_4726,N_49853,N_49841);
or UO_4727 (O_4727,N_49970,N_49988);
nor UO_4728 (O_4728,N_49955,N_49798);
or UO_4729 (O_4729,N_49838,N_49897);
or UO_4730 (O_4730,N_49933,N_49985);
or UO_4731 (O_4731,N_49790,N_49800);
nand UO_4732 (O_4732,N_49750,N_49898);
nand UO_4733 (O_4733,N_49876,N_49986);
nand UO_4734 (O_4734,N_49757,N_49891);
xor UO_4735 (O_4735,N_49916,N_49817);
and UO_4736 (O_4736,N_49915,N_49945);
nor UO_4737 (O_4737,N_49885,N_49816);
or UO_4738 (O_4738,N_49988,N_49885);
xnor UO_4739 (O_4739,N_49972,N_49963);
nand UO_4740 (O_4740,N_49778,N_49750);
or UO_4741 (O_4741,N_49901,N_49983);
xnor UO_4742 (O_4742,N_49915,N_49847);
nand UO_4743 (O_4743,N_49871,N_49924);
or UO_4744 (O_4744,N_49850,N_49983);
and UO_4745 (O_4745,N_49836,N_49982);
and UO_4746 (O_4746,N_49791,N_49899);
xnor UO_4747 (O_4747,N_49865,N_49784);
xnor UO_4748 (O_4748,N_49943,N_49880);
xnor UO_4749 (O_4749,N_49923,N_49884);
and UO_4750 (O_4750,N_49990,N_49827);
and UO_4751 (O_4751,N_49925,N_49918);
and UO_4752 (O_4752,N_49917,N_49757);
or UO_4753 (O_4753,N_49978,N_49822);
nand UO_4754 (O_4754,N_49890,N_49970);
xnor UO_4755 (O_4755,N_49991,N_49990);
and UO_4756 (O_4756,N_49965,N_49828);
nor UO_4757 (O_4757,N_49823,N_49905);
xor UO_4758 (O_4758,N_49780,N_49758);
nand UO_4759 (O_4759,N_49789,N_49823);
xnor UO_4760 (O_4760,N_49763,N_49799);
or UO_4761 (O_4761,N_49844,N_49820);
nor UO_4762 (O_4762,N_49873,N_49765);
or UO_4763 (O_4763,N_49953,N_49838);
xor UO_4764 (O_4764,N_49804,N_49848);
xor UO_4765 (O_4765,N_49814,N_49852);
xnor UO_4766 (O_4766,N_49923,N_49750);
nand UO_4767 (O_4767,N_49922,N_49945);
nand UO_4768 (O_4768,N_49926,N_49945);
or UO_4769 (O_4769,N_49876,N_49955);
and UO_4770 (O_4770,N_49974,N_49955);
nor UO_4771 (O_4771,N_49834,N_49828);
nor UO_4772 (O_4772,N_49921,N_49858);
and UO_4773 (O_4773,N_49821,N_49855);
and UO_4774 (O_4774,N_49947,N_49905);
nand UO_4775 (O_4775,N_49789,N_49798);
nor UO_4776 (O_4776,N_49834,N_49841);
and UO_4777 (O_4777,N_49805,N_49922);
or UO_4778 (O_4778,N_49966,N_49765);
nand UO_4779 (O_4779,N_49931,N_49883);
nand UO_4780 (O_4780,N_49777,N_49970);
xnor UO_4781 (O_4781,N_49971,N_49773);
xnor UO_4782 (O_4782,N_49859,N_49767);
nand UO_4783 (O_4783,N_49994,N_49766);
and UO_4784 (O_4784,N_49865,N_49970);
xnor UO_4785 (O_4785,N_49927,N_49846);
and UO_4786 (O_4786,N_49938,N_49885);
nor UO_4787 (O_4787,N_49833,N_49947);
and UO_4788 (O_4788,N_49817,N_49902);
xor UO_4789 (O_4789,N_49881,N_49965);
nand UO_4790 (O_4790,N_49926,N_49974);
xor UO_4791 (O_4791,N_49890,N_49854);
nand UO_4792 (O_4792,N_49867,N_49955);
nand UO_4793 (O_4793,N_49786,N_49770);
nand UO_4794 (O_4794,N_49983,N_49952);
and UO_4795 (O_4795,N_49968,N_49874);
xor UO_4796 (O_4796,N_49974,N_49852);
nor UO_4797 (O_4797,N_49814,N_49960);
nor UO_4798 (O_4798,N_49992,N_49977);
xnor UO_4799 (O_4799,N_49812,N_49806);
nor UO_4800 (O_4800,N_49876,N_49758);
nor UO_4801 (O_4801,N_49913,N_49826);
or UO_4802 (O_4802,N_49882,N_49871);
and UO_4803 (O_4803,N_49981,N_49958);
and UO_4804 (O_4804,N_49858,N_49957);
nand UO_4805 (O_4805,N_49947,N_49951);
and UO_4806 (O_4806,N_49857,N_49812);
and UO_4807 (O_4807,N_49957,N_49909);
xnor UO_4808 (O_4808,N_49903,N_49837);
and UO_4809 (O_4809,N_49996,N_49951);
and UO_4810 (O_4810,N_49780,N_49796);
and UO_4811 (O_4811,N_49799,N_49868);
and UO_4812 (O_4812,N_49874,N_49919);
nand UO_4813 (O_4813,N_49944,N_49879);
and UO_4814 (O_4814,N_49977,N_49930);
xor UO_4815 (O_4815,N_49927,N_49958);
or UO_4816 (O_4816,N_49940,N_49791);
nand UO_4817 (O_4817,N_49984,N_49906);
xnor UO_4818 (O_4818,N_49891,N_49989);
xor UO_4819 (O_4819,N_49942,N_49938);
or UO_4820 (O_4820,N_49930,N_49984);
or UO_4821 (O_4821,N_49863,N_49793);
or UO_4822 (O_4822,N_49898,N_49948);
xor UO_4823 (O_4823,N_49758,N_49909);
xor UO_4824 (O_4824,N_49877,N_49814);
and UO_4825 (O_4825,N_49938,N_49825);
nor UO_4826 (O_4826,N_49915,N_49753);
nand UO_4827 (O_4827,N_49901,N_49896);
nor UO_4828 (O_4828,N_49951,N_49786);
nor UO_4829 (O_4829,N_49987,N_49822);
and UO_4830 (O_4830,N_49843,N_49852);
nor UO_4831 (O_4831,N_49898,N_49819);
or UO_4832 (O_4832,N_49808,N_49782);
and UO_4833 (O_4833,N_49915,N_49937);
and UO_4834 (O_4834,N_49778,N_49841);
and UO_4835 (O_4835,N_49903,N_49816);
or UO_4836 (O_4836,N_49964,N_49800);
and UO_4837 (O_4837,N_49826,N_49947);
and UO_4838 (O_4838,N_49792,N_49787);
xor UO_4839 (O_4839,N_49879,N_49807);
or UO_4840 (O_4840,N_49844,N_49771);
nor UO_4841 (O_4841,N_49899,N_49978);
and UO_4842 (O_4842,N_49912,N_49840);
nand UO_4843 (O_4843,N_49904,N_49817);
or UO_4844 (O_4844,N_49991,N_49904);
nand UO_4845 (O_4845,N_49842,N_49844);
nor UO_4846 (O_4846,N_49919,N_49843);
nand UO_4847 (O_4847,N_49989,N_49969);
xor UO_4848 (O_4848,N_49850,N_49858);
and UO_4849 (O_4849,N_49815,N_49833);
and UO_4850 (O_4850,N_49880,N_49889);
nand UO_4851 (O_4851,N_49797,N_49763);
nor UO_4852 (O_4852,N_49899,N_49855);
nor UO_4853 (O_4853,N_49905,N_49797);
nor UO_4854 (O_4854,N_49831,N_49758);
or UO_4855 (O_4855,N_49889,N_49906);
xnor UO_4856 (O_4856,N_49978,N_49866);
xor UO_4857 (O_4857,N_49976,N_49896);
or UO_4858 (O_4858,N_49924,N_49958);
xor UO_4859 (O_4859,N_49797,N_49755);
and UO_4860 (O_4860,N_49971,N_49754);
and UO_4861 (O_4861,N_49764,N_49977);
and UO_4862 (O_4862,N_49968,N_49969);
nand UO_4863 (O_4863,N_49942,N_49878);
nand UO_4864 (O_4864,N_49763,N_49844);
nor UO_4865 (O_4865,N_49831,N_49993);
or UO_4866 (O_4866,N_49945,N_49867);
nor UO_4867 (O_4867,N_49823,N_49793);
and UO_4868 (O_4868,N_49782,N_49800);
and UO_4869 (O_4869,N_49988,N_49783);
and UO_4870 (O_4870,N_49855,N_49760);
or UO_4871 (O_4871,N_49876,N_49979);
and UO_4872 (O_4872,N_49899,N_49821);
nand UO_4873 (O_4873,N_49946,N_49760);
nor UO_4874 (O_4874,N_49889,N_49882);
and UO_4875 (O_4875,N_49781,N_49796);
nor UO_4876 (O_4876,N_49852,N_49996);
nor UO_4877 (O_4877,N_49901,N_49756);
and UO_4878 (O_4878,N_49776,N_49886);
or UO_4879 (O_4879,N_49767,N_49920);
and UO_4880 (O_4880,N_49791,N_49794);
nor UO_4881 (O_4881,N_49984,N_49970);
and UO_4882 (O_4882,N_49852,N_49777);
nand UO_4883 (O_4883,N_49966,N_49815);
and UO_4884 (O_4884,N_49755,N_49958);
or UO_4885 (O_4885,N_49834,N_49997);
nor UO_4886 (O_4886,N_49918,N_49862);
nand UO_4887 (O_4887,N_49801,N_49778);
and UO_4888 (O_4888,N_49822,N_49765);
or UO_4889 (O_4889,N_49937,N_49811);
nor UO_4890 (O_4890,N_49839,N_49805);
and UO_4891 (O_4891,N_49811,N_49974);
nor UO_4892 (O_4892,N_49977,N_49787);
and UO_4893 (O_4893,N_49786,N_49800);
and UO_4894 (O_4894,N_49821,N_49888);
and UO_4895 (O_4895,N_49936,N_49827);
nand UO_4896 (O_4896,N_49938,N_49923);
nor UO_4897 (O_4897,N_49879,N_49963);
xnor UO_4898 (O_4898,N_49799,N_49902);
nand UO_4899 (O_4899,N_49861,N_49845);
and UO_4900 (O_4900,N_49801,N_49790);
and UO_4901 (O_4901,N_49951,N_49757);
or UO_4902 (O_4902,N_49949,N_49977);
or UO_4903 (O_4903,N_49755,N_49807);
or UO_4904 (O_4904,N_49936,N_49915);
nor UO_4905 (O_4905,N_49997,N_49989);
or UO_4906 (O_4906,N_49874,N_49974);
nand UO_4907 (O_4907,N_49774,N_49941);
or UO_4908 (O_4908,N_49933,N_49921);
or UO_4909 (O_4909,N_49777,N_49982);
nor UO_4910 (O_4910,N_49796,N_49779);
xnor UO_4911 (O_4911,N_49783,N_49943);
and UO_4912 (O_4912,N_49767,N_49931);
or UO_4913 (O_4913,N_49786,N_49929);
and UO_4914 (O_4914,N_49767,N_49835);
xor UO_4915 (O_4915,N_49934,N_49833);
nand UO_4916 (O_4916,N_49846,N_49926);
nor UO_4917 (O_4917,N_49948,N_49798);
and UO_4918 (O_4918,N_49945,N_49884);
nand UO_4919 (O_4919,N_49927,N_49780);
nand UO_4920 (O_4920,N_49763,N_49956);
nor UO_4921 (O_4921,N_49852,N_49913);
or UO_4922 (O_4922,N_49829,N_49851);
nor UO_4923 (O_4923,N_49750,N_49864);
xnor UO_4924 (O_4924,N_49877,N_49762);
nor UO_4925 (O_4925,N_49832,N_49801);
nor UO_4926 (O_4926,N_49829,N_49920);
and UO_4927 (O_4927,N_49781,N_49926);
or UO_4928 (O_4928,N_49969,N_49949);
and UO_4929 (O_4929,N_49827,N_49850);
nand UO_4930 (O_4930,N_49927,N_49960);
or UO_4931 (O_4931,N_49853,N_49960);
or UO_4932 (O_4932,N_49868,N_49862);
nand UO_4933 (O_4933,N_49906,N_49915);
xnor UO_4934 (O_4934,N_49788,N_49837);
nor UO_4935 (O_4935,N_49993,N_49946);
or UO_4936 (O_4936,N_49897,N_49806);
or UO_4937 (O_4937,N_49835,N_49967);
nand UO_4938 (O_4938,N_49970,N_49962);
and UO_4939 (O_4939,N_49943,N_49881);
and UO_4940 (O_4940,N_49824,N_49827);
or UO_4941 (O_4941,N_49826,N_49959);
nor UO_4942 (O_4942,N_49888,N_49825);
or UO_4943 (O_4943,N_49982,N_49881);
xor UO_4944 (O_4944,N_49763,N_49831);
and UO_4945 (O_4945,N_49914,N_49780);
nand UO_4946 (O_4946,N_49932,N_49845);
nand UO_4947 (O_4947,N_49997,N_49893);
nand UO_4948 (O_4948,N_49771,N_49841);
or UO_4949 (O_4949,N_49807,N_49921);
or UO_4950 (O_4950,N_49922,N_49811);
nand UO_4951 (O_4951,N_49795,N_49911);
and UO_4952 (O_4952,N_49763,N_49771);
xor UO_4953 (O_4953,N_49825,N_49827);
and UO_4954 (O_4954,N_49971,N_49955);
or UO_4955 (O_4955,N_49942,N_49879);
nor UO_4956 (O_4956,N_49983,N_49891);
and UO_4957 (O_4957,N_49884,N_49817);
nand UO_4958 (O_4958,N_49814,N_49995);
nor UO_4959 (O_4959,N_49803,N_49845);
xnor UO_4960 (O_4960,N_49864,N_49973);
and UO_4961 (O_4961,N_49752,N_49896);
nand UO_4962 (O_4962,N_49932,N_49997);
nand UO_4963 (O_4963,N_49783,N_49796);
xor UO_4964 (O_4964,N_49977,N_49789);
nand UO_4965 (O_4965,N_49951,N_49839);
nand UO_4966 (O_4966,N_49791,N_49960);
nand UO_4967 (O_4967,N_49967,N_49821);
and UO_4968 (O_4968,N_49828,N_49942);
xnor UO_4969 (O_4969,N_49999,N_49797);
nor UO_4970 (O_4970,N_49940,N_49777);
and UO_4971 (O_4971,N_49988,N_49964);
and UO_4972 (O_4972,N_49869,N_49913);
or UO_4973 (O_4973,N_49917,N_49874);
nor UO_4974 (O_4974,N_49840,N_49782);
nor UO_4975 (O_4975,N_49843,N_49799);
xor UO_4976 (O_4976,N_49880,N_49791);
or UO_4977 (O_4977,N_49958,N_49987);
and UO_4978 (O_4978,N_49977,N_49771);
nor UO_4979 (O_4979,N_49936,N_49801);
nor UO_4980 (O_4980,N_49979,N_49845);
or UO_4981 (O_4981,N_49974,N_49990);
nor UO_4982 (O_4982,N_49798,N_49942);
nand UO_4983 (O_4983,N_49770,N_49895);
nand UO_4984 (O_4984,N_49792,N_49753);
and UO_4985 (O_4985,N_49996,N_49792);
or UO_4986 (O_4986,N_49793,N_49870);
and UO_4987 (O_4987,N_49959,N_49787);
nor UO_4988 (O_4988,N_49909,N_49947);
nand UO_4989 (O_4989,N_49954,N_49764);
nand UO_4990 (O_4990,N_49882,N_49763);
xnor UO_4991 (O_4991,N_49847,N_49896);
nor UO_4992 (O_4992,N_49808,N_49993);
and UO_4993 (O_4993,N_49980,N_49954);
and UO_4994 (O_4994,N_49999,N_49816);
or UO_4995 (O_4995,N_49791,N_49822);
nand UO_4996 (O_4996,N_49942,N_49872);
xor UO_4997 (O_4997,N_49892,N_49755);
or UO_4998 (O_4998,N_49778,N_49989);
nand UO_4999 (O_4999,N_49786,N_49915);
endmodule