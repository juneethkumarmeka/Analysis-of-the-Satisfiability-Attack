module basic_500_3000_500_5_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_408,In_332);
and U1 (N_1,In_240,In_255);
and U2 (N_2,In_125,In_476);
or U3 (N_3,In_177,In_15);
xnor U4 (N_4,In_368,In_374);
nand U5 (N_5,In_217,In_95);
nand U6 (N_6,In_78,In_309);
nor U7 (N_7,In_353,In_461);
and U8 (N_8,In_93,In_124);
nand U9 (N_9,In_43,In_170);
xor U10 (N_10,In_399,In_320);
nand U11 (N_11,In_107,In_335);
nand U12 (N_12,In_284,In_406);
nor U13 (N_13,In_263,In_135);
or U14 (N_14,In_387,In_407);
xnor U15 (N_15,In_236,In_56);
or U16 (N_16,In_178,In_106);
nand U17 (N_17,In_73,In_375);
or U18 (N_18,In_94,In_244);
nand U19 (N_19,In_46,In_120);
nor U20 (N_20,In_79,In_467);
or U21 (N_21,In_328,In_62);
or U22 (N_22,In_163,In_299);
and U23 (N_23,In_355,In_341);
nand U24 (N_24,In_475,In_168);
nor U25 (N_25,In_455,In_482);
and U26 (N_26,In_26,In_12);
nor U27 (N_27,In_42,In_491);
nand U28 (N_28,In_342,In_462);
or U29 (N_29,In_452,In_227);
or U30 (N_30,In_267,In_164);
nand U31 (N_31,In_154,In_54);
and U32 (N_32,In_212,In_82);
and U33 (N_33,In_5,In_325);
or U34 (N_34,In_45,In_354);
nand U35 (N_35,In_444,In_105);
or U36 (N_36,In_490,In_9);
nor U37 (N_37,In_349,In_428);
or U38 (N_38,In_142,In_228);
or U39 (N_39,In_216,In_454);
and U40 (N_40,In_189,In_239);
or U41 (N_41,In_259,In_118);
and U42 (N_42,In_226,In_38);
or U43 (N_43,In_283,In_485);
and U44 (N_44,In_439,In_415);
and U45 (N_45,In_99,In_384);
and U46 (N_46,In_235,In_151);
and U47 (N_47,In_278,In_186);
nand U48 (N_48,In_366,In_130);
or U49 (N_49,In_197,In_331);
or U50 (N_50,In_131,In_139);
nor U51 (N_51,In_53,In_250);
and U52 (N_52,In_191,In_393);
or U53 (N_53,In_49,In_345);
nor U54 (N_54,In_499,In_385);
nand U55 (N_55,In_29,In_13);
and U56 (N_56,In_58,In_258);
or U57 (N_57,In_60,In_100);
and U58 (N_58,In_460,In_492);
and U59 (N_59,In_322,In_3);
nor U60 (N_60,In_27,In_184);
nand U61 (N_61,In_425,In_363);
or U62 (N_62,In_33,In_223);
or U63 (N_63,In_442,In_487);
nor U64 (N_64,In_8,In_372);
nor U65 (N_65,In_419,In_338);
nand U66 (N_66,In_55,In_149);
or U67 (N_67,In_451,In_463);
and U68 (N_68,In_378,In_296);
and U69 (N_69,In_376,In_411);
and U70 (N_70,In_39,In_126);
nor U71 (N_71,In_167,In_72);
or U72 (N_72,In_192,In_31);
nor U73 (N_73,In_185,In_478);
or U74 (N_74,In_420,In_351);
nor U75 (N_75,In_306,In_447);
nor U76 (N_76,In_104,In_183);
nand U77 (N_77,In_249,In_219);
nand U78 (N_78,In_300,In_290);
and U79 (N_79,In_64,In_22);
or U80 (N_80,In_254,In_247);
nor U81 (N_81,In_358,In_129);
nor U82 (N_82,In_238,In_352);
nor U83 (N_83,In_230,In_148);
nand U84 (N_84,In_484,In_357);
and U85 (N_85,In_251,In_295);
and U86 (N_86,In_233,In_396);
and U87 (N_87,In_280,In_279);
and U88 (N_88,In_222,In_336);
or U89 (N_89,In_18,In_37);
or U90 (N_90,In_285,In_339);
and U91 (N_91,In_133,In_398);
nand U92 (N_92,In_416,In_426);
or U93 (N_93,In_289,In_234);
nor U94 (N_94,In_413,In_66);
nor U95 (N_95,In_272,In_44);
and U96 (N_96,In_496,In_147);
nand U97 (N_97,In_369,In_114);
or U98 (N_98,In_174,In_75);
and U99 (N_99,In_266,In_382);
nor U100 (N_100,In_268,In_248);
and U101 (N_101,In_483,In_152);
nor U102 (N_102,In_294,In_136);
and U103 (N_103,In_179,In_346);
or U104 (N_104,In_434,In_456);
nor U105 (N_105,In_457,In_450);
and U106 (N_106,In_314,In_344);
and U107 (N_107,In_221,In_122);
or U108 (N_108,In_220,In_246);
nor U109 (N_109,In_313,In_423);
nor U110 (N_110,In_340,In_310);
nand U111 (N_111,In_421,In_394);
and U112 (N_112,In_422,In_440);
nor U113 (N_113,In_291,In_229);
nand U114 (N_114,In_176,In_480);
nor U115 (N_115,In_337,In_318);
and U116 (N_116,In_424,In_269);
nand U117 (N_117,In_157,In_101);
or U118 (N_118,In_397,In_199);
and U119 (N_119,In_202,In_145);
nor U120 (N_120,In_270,In_165);
and U121 (N_121,In_11,In_326);
or U122 (N_122,In_281,In_321);
nor U123 (N_123,In_333,In_103);
and U124 (N_124,In_86,In_276);
and U125 (N_125,In_453,In_111);
nor U126 (N_126,In_19,In_493);
and U127 (N_127,In_465,In_418);
and U128 (N_128,In_97,In_243);
nor U129 (N_129,In_21,In_256);
or U130 (N_130,In_65,In_57);
nand U131 (N_131,In_260,In_274);
nand U132 (N_132,In_116,In_377);
nand U133 (N_133,In_262,In_14);
or U134 (N_134,In_265,In_412);
or U135 (N_135,In_445,In_200);
nand U136 (N_136,In_297,In_92);
nand U137 (N_137,In_30,In_10);
and U138 (N_138,In_359,In_261);
nand U139 (N_139,In_273,In_298);
and U140 (N_140,In_213,In_446);
nand U141 (N_141,In_218,In_305);
nor U142 (N_142,In_315,In_67);
nor U143 (N_143,In_96,In_41);
and U144 (N_144,In_311,In_119);
and U145 (N_145,In_121,In_312);
and U146 (N_146,In_373,In_171);
nor U147 (N_147,In_379,In_90);
nor U148 (N_148,In_25,In_209);
nand U149 (N_149,In_401,In_390);
nand U150 (N_150,In_253,In_205);
nor U151 (N_151,In_464,In_370);
and U152 (N_152,In_159,In_417);
nand U153 (N_153,In_391,In_409);
or U154 (N_154,In_365,In_431);
or U155 (N_155,In_51,In_190);
nor U156 (N_156,In_257,In_201);
nand U157 (N_157,In_360,In_180);
or U158 (N_158,In_316,In_83);
and U159 (N_159,In_308,In_195);
or U160 (N_160,In_182,In_252);
nand U161 (N_161,In_225,In_395);
nand U162 (N_162,In_172,In_34);
nor U163 (N_163,In_347,In_128);
nand U164 (N_164,In_286,In_486);
nand U165 (N_165,In_132,In_59);
and U166 (N_166,In_323,In_329);
nand U167 (N_167,In_473,In_245);
and U168 (N_168,In_113,In_211);
nand U169 (N_169,In_292,In_98);
nand U170 (N_170,In_293,In_466);
and U171 (N_171,In_459,In_361);
and U172 (N_172,In_153,In_74);
nor U173 (N_173,In_140,In_63);
and U174 (N_174,In_348,In_224);
or U175 (N_175,In_437,In_489);
nand U176 (N_176,In_61,In_88);
or U177 (N_177,In_242,In_410);
nor U178 (N_178,In_343,In_498);
nor U179 (N_179,In_32,In_468);
nor U180 (N_180,In_123,In_48);
nand U181 (N_181,In_141,In_441);
or U182 (N_182,In_364,In_169);
and U183 (N_183,In_414,In_134);
and U184 (N_184,In_317,In_303);
and U185 (N_185,In_334,In_85);
nand U186 (N_186,In_231,In_77);
nand U187 (N_187,In_495,In_68);
nand U188 (N_188,In_443,In_367);
and U189 (N_189,In_2,In_472);
and U190 (N_190,In_458,In_324);
and U191 (N_191,In_356,In_20);
or U192 (N_192,In_102,In_181);
nor U193 (N_193,In_319,In_108);
nor U194 (N_194,In_112,In_282);
and U195 (N_195,In_388,In_194);
nor U196 (N_196,In_403,In_16);
and U197 (N_197,In_166,In_214);
and U198 (N_198,In_50,In_474);
nor U199 (N_199,In_156,In_430);
nor U200 (N_200,In_481,In_84);
or U201 (N_201,In_138,In_362);
nor U202 (N_202,In_173,In_404);
and U203 (N_203,In_302,In_47);
and U204 (N_204,In_386,In_160);
and U205 (N_205,In_69,In_40);
and U206 (N_206,In_232,In_203);
nor U207 (N_207,In_400,In_448);
and U208 (N_208,In_381,In_155);
nor U209 (N_209,In_237,In_469);
and U210 (N_210,In_198,In_497);
or U211 (N_211,In_1,In_80);
nor U212 (N_212,In_71,In_188);
nand U213 (N_213,In_162,In_193);
or U214 (N_214,In_241,In_402);
nand U215 (N_215,In_0,In_161);
nor U216 (N_216,In_115,In_350);
or U217 (N_217,In_158,In_36);
nand U218 (N_218,In_210,In_277);
nand U219 (N_219,In_81,In_144);
nor U220 (N_220,In_429,In_432);
or U221 (N_221,In_494,In_206);
nor U222 (N_222,In_204,In_470);
nor U223 (N_223,In_150,In_208);
nor U224 (N_224,In_6,In_389);
or U225 (N_225,In_383,In_264);
and U226 (N_226,In_477,In_91);
nor U227 (N_227,In_110,In_392);
nand U228 (N_228,In_23,In_187);
nor U229 (N_229,In_196,In_438);
or U230 (N_230,In_127,In_330);
nand U231 (N_231,In_109,In_287);
and U232 (N_232,In_405,In_479);
nor U233 (N_233,In_89,In_288);
or U234 (N_234,In_488,In_146);
nand U235 (N_235,In_436,In_327);
nor U236 (N_236,In_35,In_435);
and U237 (N_237,In_207,In_87);
nor U238 (N_238,In_70,In_17);
or U239 (N_239,In_117,In_215);
and U240 (N_240,In_28,In_307);
nor U241 (N_241,In_143,In_175);
or U242 (N_242,In_427,In_380);
or U243 (N_243,In_271,In_7);
or U244 (N_244,In_433,In_76);
or U245 (N_245,In_24,In_137);
or U246 (N_246,In_371,In_52);
nor U247 (N_247,In_275,In_449);
nor U248 (N_248,In_304,In_471);
or U249 (N_249,In_301,In_4);
or U250 (N_250,In_256,In_287);
nand U251 (N_251,In_335,In_286);
or U252 (N_252,In_139,In_430);
or U253 (N_253,In_441,In_269);
or U254 (N_254,In_180,In_364);
nor U255 (N_255,In_35,In_473);
nor U256 (N_256,In_332,In_262);
or U257 (N_257,In_154,In_52);
or U258 (N_258,In_124,In_34);
nor U259 (N_259,In_152,In_115);
nand U260 (N_260,In_74,In_135);
and U261 (N_261,In_429,In_334);
nand U262 (N_262,In_259,In_412);
nor U263 (N_263,In_299,In_78);
or U264 (N_264,In_253,In_51);
nand U265 (N_265,In_428,In_151);
or U266 (N_266,In_454,In_260);
or U267 (N_267,In_71,In_445);
or U268 (N_268,In_179,In_47);
and U269 (N_269,In_47,In_361);
and U270 (N_270,In_430,In_4);
nor U271 (N_271,In_19,In_382);
and U272 (N_272,In_242,In_164);
nand U273 (N_273,In_376,In_35);
nor U274 (N_274,In_440,In_428);
and U275 (N_275,In_408,In_280);
nand U276 (N_276,In_147,In_358);
and U277 (N_277,In_42,In_382);
nand U278 (N_278,In_339,In_147);
nor U279 (N_279,In_422,In_323);
nand U280 (N_280,In_147,In_371);
and U281 (N_281,In_143,In_381);
nor U282 (N_282,In_462,In_302);
nand U283 (N_283,In_28,In_300);
nand U284 (N_284,In_227,In_136);
nor U285 (N_285,In_134,In_218);
and U286 (N_286,In_498,In_360);
or U287 (N_287,In_251,In_60);
or U288 (N_288,In_343,In_389);
nand U289 (N_289,In_7,In_390);
nor U290 (N_290,In_233,In_129);
and U291 (N_291,In_323,In_343);
nand U292 (N_292,In_196,In_233);
or U293 (N_293,In_232,In_377);
or U294 (N_294,In_458,In_133);
or U295 (N_295,In_13,In_111);
and U296 (N_296,In_170,In_473);
and U297 (N_297,In_215,In_246);
nor U298 (N_298,In_134,In_301);
or U299 (N_299,In_176,In_400);
or U300 (N_300,In_251,In_74);
nand U301 (N_301,In_357,In_455);
or U302 (N_302,In_159,In_426);
nand U303 (N_303,In_146,In_249);
or U304 (N_304,In_92,In_111);
nand U305 (N_305,In_198,In_343);
nor U306 (N_306,In_382,In_25);
nor U307 (N_307,In_204,In_400);
nor U308 (N_308,In_414,In_319);
nand U309 (N_309,In_379,In_254);
nor U310 (N_310,In_225,In_381);
nor U311 (N_311,In_227,In_9);
nor U312 (N_312,In_331,In_173);
nand U313 (N_313,In_123,In_377);
nor U314 (N_314,In_65,In_168);
nand U315 (N_315,In_226,In_356);
nand U316 (N_316,In_240,In_459);
nor U317 (N_317,In_433,In_117);
and U318 (N_318,In_497,In_252);
nand U319 (N_319,In_135,In_99);
and U320 (N_320,In_493,In_165);
nor U321 (N_321,In_55,In_484);
nand U322 (N_322,In_101,In_131);
or U323 (N_323,In_51,In_465);
or U324 (N_324,In_470,In_377);
nor U325 (N_325,In_280,In_427);
nor U326 (N_326,In_227,In_427);
nor U327 (N_327,In_77,In_456);
nand U328 (N_328,In_260,In_497);
or U329 (N_329,In_180,In_340);
or U330 (N_330,In_450,In_363);
and U331 (N_331,In_135,In_56);
or U332 (N_332,In_265,In_376);
nor U333 (N_333,In_182,In_38);
nor U334 (N_334,In_395,In_330);
nor U335 (N_335,In_317,In_335);
nor U336 (N_336,In_222,In_81);
and U337 (N_337,In_426,In_74);
and U338 (N_338,In_105,In_156);
and U339 (N_339,In_139,In_225);
or U340 (N_340,In_96,In_51);
nor U341 (N_341,In_352,In_249);
nand U342 (N_342,In_407,In_246);
nor U343 (N_343,In_450,In_73);
nor U344 (N_344,In_325,In_460);
nand U345 (N_345,In_427,In_248);
and U346 (N_346,In_5,In_328);
nand U347 (N_347,In_269,In_407);
and U348 (N_348,In_196,In_288);
nand U349 (N_349,In_401,In_416);
and U350 (N_350,In_207,In_302);
or U351 (N_351,In_235,In_293);
or U352 (N_352,In_1,In_275);
nor U353 (N_353,In_107,In_165);
nand U354 (N_354,In_232,In_487);
nor U355 (N_355,In_405,In_194);
or U356 (N_356,In_262,In_341);
and U357 (N_357,In_450,In_425);
nor U358 (N_358,In_132,In_143);
nor U359 (N_359,In_188,In_235);
nor U360 (N_360,In_377,In_69);
nand U361 (N_361,In_22,In_258);
nor U362 (N_362,In_328,In_38);
nor U363 (N_363,In_262,In_368);
or U364 (N_364,In_24,In_245);
or U365 (N_365,In_178,In_270);
or U366 (N_366,In_265,In_435);
and U367 (N_367,In_64,In_2);
and U368 (N_368,In_76,In_342);
nor U369 (N_369,In_469,In_371);
or U370 (N_370,In_237,In_131);
nand U371 (N_371,In_405,In_74);
nor U372 (N_372,In_259,In_74);
and U373 (N_373,In_333,In_468);
nand U374 (N_374,In_467,In_205);
and U375 (N_375,In_91,In_195);
or U376 (N_376,In_240,In_93);
nor U377 (N_377,In_5,In_210);
or U378 (N_378,In_261,In_471);
nor U379 (N_379,In_282,In_68);
or U380 (N_380,In_66,In_273);
or U381 (N_381,In_96,In_470);
xor U382 (N_382,In_93,In_336);
and U383 (N_383,In_39,In_233);
nand U384 (N_384,In_325,In_388);
or U385 (N_385,In_2,In_57);
and U386 (N_386,In_190,In_321);
nor U387 (N_387,In_379,In_46);
or U388 (N_388,In_369,In_4);
nor U389 (N_389,In_263,In_120);
nand U390 (N_390,In_249,In_412);
nor U391 (N_391,In_132,In_136);
nand U392 (N_392,In_286,In_211);
or U393 (N_393,In_280,In_174);
or U394 (N_394,In_57,In_401);
nand U395 (N_395,In_306,In_249);
and U396 (N_396,In_316,In_131);
nor U397 (N_397,In_344,In_173);
or U398 (N_398,In_417,In_234);
nand U399 (N_399,In_171,In_446);
nor U400 (N_400,In_430,In_54);
nand U401 (N_401,In_446,In_460);
or U402 (N_402,In_175,In_112);
nand U403 (N_403,In_237,In_365);
nand U404 (N_404,In_312,In_188);
nor U405 (N_405,In_64,In_257);
and U406 (N_406,In_123,In_256);
or U407 (N_407,In_486,In_451);
and U408 (N_408,In_95,In_291);
nor U409 (N_409,In_426,In_398);
and U410 (N_410,In_431,In_201);
nand U411 (N_411,In_243,In_269);
nor U412 (N_412,In_149,In_233);
and U413 (N_413,In_96,In_122);
and U414 (N_414,In_312,In_323);
nor U415 (N_415,In_276,In_180);
or U416 (N_416,In_189,In_206);
and U417 (N_417,In_306,In_245);
and U418 (N_418,In_479,In_367);
or U419 (N_419,In_9,In_379);
and U420 (N_420,In_239,In_475);
or U421 (N_421,In_171,In_124);
nor U422 (N_422,In_35,In_180);
nor U423 (N_423,In_162,In_276);
or U424 (N_424,In_2,In_249);
nand U425 (N_425,In_237,In_184);
and U426 (N_426,In_287,In_96);
nor U427 (N_427,In_341,In_128);
nor U428 (N_428,In_350,In_292);
nor U429 (N_429,In_159,In_398);
nor U430 (N_430,In_282,In_123);
and U431 (N_431,In_257,In_213);
nor U432 (N_432,In_301,In_16);
and U433 (N_433,In_304,In_414);
and U434 (N_434,In_338,In_95);
nand U435 (N_435,In_91,In_416);
and U436 (N_436,In_90,In_485);
nor U437 (N_437,In_238,In_202);
nand U438 (N_438,In_304,In_486);
nor U439 (N_439,In_400,In_20);
nor U440 (N_440,In_186,In_487);
nand U441 (N_441,In_332,In_325);
nand U442 (N_442,In_425,In_491);
nand U443 (N_443,In_223,In_236);
or U444 (N_444,In_183,In_76);
nor U445 (N_445,In_240,In_409);
nor U446 (N_446,In_215,In_253);
nand U447 (N_447,In_104,In_318);
xor U448 (N_448,In_196,In_395);
or U449 (N_449,In_288,In_116);
nor U450 (N_450,In_167,In_93);
nand U451 (N_451,In_402,In_363);
and U452 (N_452,In_233,In_165);
nor U453 (N_453,In_5,In_346);
and U454 (N_454,In_437,In_227);
nand U455 (N_455,In_355,In_316);
or U456 (N_456,In_186,In_43);
nor U457 (N_457,In_205,In_412);
or U458 (N_458,In_189,In_405);
nor U459 (N_459,In_335,In_297);
or U460 (N_460,In_170,In_433);
or U461 (N_461,In_257,In_106);
or U462 (N_462,In_317,In_346);
or U463 (N_463,In_28,In_309);
nor U464 (N_464,In_390,In_457);
nand U465 (N_465,In_467,In_64);
and U466 (N_466,In_214,In_70);
and U467 (N_467,In_497,In_142);
and U468 (N_468,In_45,In_397);
nor U469 (N_469,In_85,In_357);
or U470 (N_470,In_395,In_406);
nand U471 (N_471,In_237,In_112);
or U472 (N_472,In_496,In_459);
nor U473 (N_473,In_225,In_472);
nand U474 (N_474,In_329,In_10);
nor U475 (N_475,In_386,In_476);
nor U476 (N_476,In_263,In_237);
xor U477 (N_477,In_86,In_96);
nand U478 (N_478,In_412,In_256);
nand U479 (N_479,In_57,In_489);
nand U480 (N_480,In_484,In_393);
and U481 (N_481,In_467,In_169);
nand U482 (N_482,In_301,In_2);
and U483 (N_483,In_357,In_72);
nand U484 (N_484,In_392,In_444);
and U485 (N_485,In_441,In_391);
or U486 (N_486,In_207,In_265);
nor U487 (N_487,In_447,In_378);
nor U488 (N_488,In_182,In_451);
nor U489 (N_489,In_337,In_203);
or U490 (N_490,In_461,In_167);
or U491 (N_491,In_197,In_163);
and U492 (N_492,In_481,In_402);
and U493 (N_493,In_255,In_102);
nor U494 (N_494,In_189,In_253);
nand U495 (N_495,In_228,In_441);
and U496 (N_496,In_108,In_34);
nand U497 (N_497,In_77,In_125);
and U498 (N_498,In_51,In_217);
nand U499 (N_499,In_447,In_241);
xnor U500 (N_500,In_104,In_57);
nor U501 (N_501,In_27,In_373);
and U502 (N_502,In_73,In_381);
or U503 (N_503,In_60,In_7);
nand U504 (N_504,In_436,In_226);
nor U505 (N_505,In_157,In_326);
and U506 (N_506,In_342,In_346);
nor U507 (N_507,In_260,In_217);
nor U508 (N_508,In_383,In_378);
and U509 (N_509,In_387,In_152);
and U510 (N_510,In_199,In_333);
and U511 (N_511,In_316,In_39);
or U512 (N_512,In_193,In_43);
nor U513 (N_513,In_374,In_296);
and U514 (N_514,In_488,In_212);
and U515 (N_515,In_456,In_283);
nand U516 (N_516,In_357,In_125);
or U517 (N_517,In_12,In_64);
nand U518 (N_518,In_145,In_9);
nand U519 (N_519,In_230,In_284);
or U520 (N_520,In_33,In_194);
and U521 (N_521,In_419,In_173);
or U522 (N_522,In_127,In_441);
nor U523 (N_523,In_36,In_253);
or U524 (N_524,In_407,In_235);
nand U525 (N_525,In_471,In_70);
and U526 (N_526,In_375,In_456);
nand U527 (N_527,In_37,In_131);
nand U528 (N_528,In_366,In_185);
nand U529 (N_529,In_177,In_186);
nand U530 (N_530,In_281,In_357);
nor U531 (N_531,In_255,In_325);
and U532 (N_532,In_87,In_100);
nor U533 (N_533,In_287,In_295);
nand U534 (N_534,In_196,In_261);
and U535 (N_535,In_235,In_144);
or U536 (N_536,In_431,In_181);
nand U537 (N_537,In_427,In_26);
nor U538 (N_538,In_245,In_388);
and U539 (N_539,In_420,In_209);
nor U540 (N_540,In_115,In_240);
nor U541 (N_541,In_5,In_383);
nand U542 (N_542,In_126,In_181);
xnor U543 (N_543,In_456,In_426);
or U544 (N_544,In_113,In_120);
nand U545 (N_545,In_13,In_100);
nor U546 (N_546,In_436,In_473);
nor U547 (N_547,In_454,In_484);
and U548 (N_548,In_482,In_38);
and U549 (N_549,In_236,In_182);
nand U550 (N_550,In_339,In_305);
nor U551 (N_551,In_69,In_122);
nand U552 (N_552,In_326,In_404);
nor U553 (N_553,In_129,In_147);
and U554 (N_554,In_128,In_230);
and U555 (N_555,In_346,In_181);
nand U556 (N_556,In_249,In_98);
or U557 (N_557,In_221,In_424);
nor U558 (N_558,In_66,In_303);
and U559 (N_559,In_261,In_159);
and U560 (N_560,In_34,In_206);
and U561 (N_561,In_469,In_349);
and U562 (N_562,In_254,In_426);
or U563 (N_563,In_194,In_377);
nor U564 (N_564,In_433,In_144);
nand U565 (N_565,In_12,In_192);
and U566 (N_566,In_211,In_3);
xnor U567 (N_567,In_312,In_325);
or U568 (N_568,In_184,In_462);
nand U569 (N_569,In_109,In_383);
or U570 (N_570,In_357,In_353);
or U571 (N_571,In_9,In_231);
nand U572 (N_572,In_405,In_165);
nand U573 (N_573,In_113,In_202);
and U574 (N_574,In_377,In_214);
nand U575 (N_575,In_71,In_337);
nor U576 (N_576,In_335,In_482);
or U577 (N_577,In_30,In_256);
and U578 (N_578,In_467,In_395);
or U579 (N_579,In_233,In_409);
and U580 (N_580,In_209,In_138);
and U581 (N_581,In_157,In_224);
nand U582 (N_582,In_493,In_54);
nand U583 (N_583,In_107,In_464);
and U584 (N_584,In_436,In_479);
nor U585 (N_585,In_474,In_93);
or U586 (N_586,In_245,In_186);
and U587 (N_587,In_173,In_99);
or U588 (N_588,In_26,In_97);
and U589 (N_589,In_91,In_420);
or U590 (N_590,In_228,In_363);
nand U591 (N_591,In_22,In_227);
and U592 (N_592,In_47,In_120);
nor U593 (N_593,In_276,In_434);
nor U594 (N_594,In_460,In_135);
nor U595 (N_595,In_204,In_330);
nor U596 (N_596,In_24,In_368);
nand U597 (N_597,In_457,In_312);
nand U598 (N_598,In_351,In_250);
and U599 (N_599,In_134,In_158);
or U600 (N_600,N_395,N_590);
nand U601 (N_601,N_476,N_57);
and U602 (N_602,N_62,N_322);
and U603 (N_603,N_261,N_9);
nor U604 (N_604,N_508,N_377);
nand U605 (N_605,N_234,N_162);
or U606 (N_606,N_315,N_132);
nor U607 (N_607,N_169,N_477);
and U608 (N_608,N_595,N_555);
nand U609 (N_609,N_482,N_328);
xnor U610 (N_610,N_63,N_324);
nor U611 (N_611,N_164,N_306);
nor U612 (N_612,N_405,N_274);
nor U613 (N_613,N_280,N_188);
nor U614 (N_614,N_128,N_20);
and U615 (N_615,N_537,N_354);
nand U616 (N_616,N_446,N_109);
nand U617 (N_617,N_309,N_499);
or U618 (N_618,N_97,N_443);
nand U619 (N_619,N_168,N_526);
and U620 (N_620,N_409,N_282);
and U621 (N_621,N_198,N_331);
xor U622 (N_622,N_372,N_156);
nand U623 (N_623,N_58,N_213);
nand U624 (N_624,N_359,N_289);
or U625 (N_625,N_146,N_390);
or U626 (N_626,N_424,N_119);
or U627 (N_627,N_468,N_226);
and U628 (N_628,N_129,N_279);
nor U629 (N_629,N_28,N_91);
or U630 (N_630,N_158,N_16);
nor U631 (N_631,N_136,N_380);
nor U632 (N_632,N_458,N_336);
and U633 (N_633,N_467,N_243);
nand U634 (N_634,N_242,N_364);
or U635 (N_635,N_233,N_301);
nor U636 (N_636,N_286,N_6);
nor U637 (N_637,N_398,N_50);
xnor U638 (N_638,N_216,N_444);
nor U639 (N_639,N_370,N_399);
nand U640 (N_640,N_149,N_13);
and U641 (N_641,N_59,N_358);
and U642 (N_642,N_277,N_452);
xor U643 (N_643,N_382,N_278);
and U644 (N_644,N_108,N_22);
and U645 (N_645,N_423,N_394);
nor U646 (N_646,N_171,N_321);
nor U647 (N_647,N_159,N_337);
nand U648 (N_648,N_250,N_193);
and U649 (N_649,N_173,N_522);
nor U650 (N_650,N_362,N_412);
or U651 (N_651,N_256,N_589);
nor U652 (N_652,N_167,N_204);
or U653 (N_653,N_512,N_130);
and U654 (N_654,N_392,N_435);
nor U655 (N_655,N_562,N_599);
or U656 (N_656,N_383,N_96);
and U657 (N_657,N_471,N_77);
nor U658 (N_658,N_304,N_148);
and U659 (N_659,N_459,N_384);
nand U660 (N_660,N_554,N_369);
or U661 (N_661,N_411,N_70);
and U662 (N_662,N_191,N_560);
nand U663 (N_663,N_347,N_527);
nor U664 (N_664,N_351,N_115);
and U665 (N_665,N_549,N_426);
nand U666 (N_666,N_201,N_397);
or U667 (N_667,N_273,N_150);
and U668 (N_668,N_564,N_469);
or U669 (N_669,N_550,N_567);
or U670 (N_670,N_186,N_406);
nand U671 (N_671,N_539,N_401);
nand U672 (N_672,N_75,N_525);
or U673 (N_673,N_12,N_245);
nand U674 (N_674,N_396,N_393);
nand U675 (N_675,N_429,N_160);
nand U676 (N_676,N_323,N_232);
or U677 (N_677,N_574,N_83);
and U678 (N_678,N_532,N_504);
nand U679 (N_679,N_34,N_78);
and U680 (N_680,N_586,N_182);
nor U681 (N_681,N_592,N_408);
or U682 (N_682,N_440,N_219);
and U683 (N_683,N_436,N_457);
nor U684 (N_684,N_90,N_583);
nor U685 (N_685,N_536,N_214);
nand U686 (N_686,N_461,N_338);
nor U687 (N_687,N_262,N_177);
and U688 (N_688,N_531,N_137);
nand U689 (N_689,N_30,N_462);
or U690 (N_690,N_495,N_346);
or U691 (N_691,N_47,N_41);
and U692 (N_692,N_546,N_183);
nor U693 (N_693,N_294,N_76);
or U694 (N_694,N_51,N_366);
nand U695 (N_695,N_378,N_4);
or U696 (N_696,N_500,N_180);
nor U697 (N_697,N_195,N_179);
nand U698 (N_698,N_221,N_343);
nand U699 (N_699,N_127,N_237);
nand U700 (N_700,N_283,N_120);
and U701 (N_701,N_478,N_84);
and U702 (N_702,N_253,N_285);
or U703 (N_703,N_433,N_535);
and U704 (N_704,N_33,N_502);
and U705 (N_705,N_140,N_0);
or U706 (N_706,N_441,N_86);
nand U707 (N_707,N_481,N_208);
nor U708 (N_708,N_207,N_229);
and U709 (N_709,N_507,N_327);
and U710 (N_710,N_330,N_202);
nand U711 (N_711,N_316,N_473);
nand U712 (N_712,N_260,N_295);
or U713 (N_713,N_225,N_192);
and U714 (N_714,N_485,N_329);
nor U715 (N_715,N_552,N_530);
nor U716 (N_716,N_326,N_422);
nand U717 (N_717,N_486,N_463);
or U718 (N_718,N_506,N_587);
nand U719 (N_719,N_116,N_52);
and U720 (N_720,N_534,N_439);
nor U721 (N_721,N_565,N_8);
and U722 (N_722,N_15,N_352);
and U723 (N_723,N_480,N_453);
nor U724 (N_724,N_573,N_529);
and U725 (N_725,N_310,N_494);
and U726 (N_726,N_227,N_342);
and U727 (N_727,N_118,N_81);
and U728 (N_728,N_498,N_542);
and U729 (N_729,N_135,N_110);
nor U730 (N_730,N_489,N_17);
and U731 (N_731,N_428,N_79);
nand U732 (N_732,N_111,N_284);
nand U733 (N_733,N_217,N_1);
nand U734 (N_734,N_187,N_7);
nor U735 (N_735,N_38,N_355);
nor U736 (N_736,N_484,N_367);
nand U737 (N_737,N_60,N_246);
nor U738 (N_738,N_123,N_153);
nand U739 (N_739,N_302,N_548);
nand U740 (N_740,N_54,N_487);
nand U741 (N_741,N_212,N_174);
nand U742 (N_742,N_319,N_597);
nand U743 (N_743,N_298,N_2);
nand U744 (N_744,N_449,N_505);
and U745 (N_745,N_416,N_563);
or U746 (N_746,N_48,N_27);
nor U747 (N_747,N_68,N_223);
or U748 (N_748,N_185,N_345);
and U749 (N_749,N_475,N_568);
and U750 (N_750,N_228,N_559);
nor U751 (N_751,N_511,N_403);
nor U752 (N_752,N_584,N_385);
nor U753 (N_753,N_272,N_579);
nor U754 (N_754,N_203,N_538);
nor U755 (N_755,N_196,N_107);
and U756 (N_756,N_23,N_49);
or U757 (N_757,N_124,N_572);
nand U758 (N_758,N_210,N_145);
nand U759 (N_759,N_308,N_190);
nand U760 (N_760,N_281,N_155);
nand U761 (N_761,N_556,N_543);
nor U762 (N_762,N_430,N_222);
nor U763 (N_763,N_438,N_236);
or U764 (N_764,N_305,N_26);
and U765 (N_765,N_239,N_455);
nand U766 (N_766,N_580,N_102);
and U767 (N_767,N_402,N_501);
and U768 (N_768,N_252,N_161);
nor U769 (N_769,N_66,N_348);
nor U770 (N_770,N_126,N_561);
nor U771 (N_771,N_11,N_540);
nand U772 (N_772,N_19,N_518);
or U773 (N_773,N_288,N_10);
or U774 (N_774,N_425,N_447);
or U775 (N_775,N_307,N_332);
or U776 (N_776,N_39,N_200);
or U777 (N_777,N_244,N_492);
nor U778 (N_778,N_205,N_259);
or U779 (N_779,N_264,N_598);
nor U780 (N_780,N_206,N_588);
and U781 (N_781,N_464,N_176);
nand U782 (N_782,N_303,N_296);
nor U783 (N_783,N_254,N_379);
and U784 (N_784,N_42,N_69);
or U785 (N_785,N_163,N_551);
or U786 (N_786,N_299,N_88);
or U787 (N_787,N_133,N_29);
and U788 (N_788,N_85,N_98);
and U789 (N_789,N_404,N_381);
or U790 (N_790,N_341,N_40);
or U791 (N_791,N_553,N_516);
nor U792 (N_792,N_357,N_215);
nand U793 (N_793,N_44,N_139);
nor U794 (N_794,N_271,N_94);
and U795 (N_795,N_391,N_99);
and U796 (N_796,N_544,N_350);
or U797 (N_797,N_576,N_419);
and U798 (N_798,N_65,N_18);
and U799 (N_799,N_292,N_21);
nor U800 (N_800,N_270,N_172);
nor U801 (N_801,N_56,N_312);
nor U802 (N_802,N_365,N_87);
or U803 (N_803,N_231,N_194);
nand U804 (N_804,N_479,N_593);
and U805 (N_805,N_71,N_434);
and U806 (N_806,N_368,N_258);
nor U807 (N_807,N_14,N_491);
nand U808 (N_808,N_141,N_493);
nand U809 (N_809,N_165,N_442);
nor U810 (N_810,N_175,N_437);
nand U811 (N_811,N_389,N_325);
or U812 (N_812,N_519,N_121);
nor U813 (N_813,N_5,N_386);
nand U814 (N_814,N_95,N_503);
nor U815 (N_815,N_445,N_67);
and U816 (N_816,N_374,N_266);
and U817 (N_817,N_427,N_334);
or U818 (N_818,N_344,N_74);
nand U819 (N_819,N_515,N_72);
or U820 (N_820,N_300,N_496);
nand U821 (N_821,N_240,N_199);
and U822 (N_822,N_353,N_104);
and U823 (N_823,N_117,N_569);
nor U824 (N_824,N_418,N_35);
xnor U825 (N_825,N_275,N_361);
nor U826 (N_826,N_454,N_147);
or U827 (N_827,N_388,N_36);
or U828 (N_828,N_510,N_349);
and U829 (N_829,N_43,N_46);
and U830 (N_830,N_170,N_73);
and U831 (N_831,N_520,N_356);
nor U832 (N_832,N_460,N_92);
nand U833 (N_833,N_166,N_513);
nor U834 (N_834,N_276,N_410);
and U835 (N_835,N_267,N_112);
or U836 (N_836,N_230,N_297);
or U837 (N_837,N_456,N_413);
nand U838 (N_838,N_255,N_157);
nand U839 (N_839,N_363,N_218);
and U840 (N_840,N_596,N_93);
nor U841 (N_841,N_541,N_293);
or U842 (N_842,N_415,N_82);
and U843 (N_843,N_64,N_474);
or U844 (N_844,N_263,N_220);
or U845 (N_845,N_497,N_318);
nor U846 (N_846,N_448,N_178);
or U847 (N_847,N_470,N_247);
or U848 (N_848,N_31,N_578);
nor U849 (N_849,N_483,N_545);
nor U850 (N_850,N_523,N_122);
or U851 (N_851,N_407,N_131);
nor U852 (N_852,N_450,N_209);
nand U853 (N_853,N_557,N_431);
nand U854 (N_854,N_333,N_80);
or U855 (N_855,N_101,N_524);
or U856 (N_856,N_594,N_181);
nor U857 (N_857,N_375,N_61);
nor U858 (N_858,N_314,N_142);
or U859 (N_859,N_3,N_241);
or U860 (N_860,N_340,N_514);
nand U861 (N_861,N_373,N_224);
nand U862 (N_862,N_189,N_238);
and U863 (N_863,N_211,N_290);
nand U864 (N_864,N_197,N_184);
nand U865 (N_865,N_151,N_339);
nor U866 (N_866,N_25,N_582);
nand U867 (N_867,N_591,N_103);
and U868 (N_868,N_32,N_420);
and U869 (N_869,N_414,N_387);
and U870 (N_870,N_488,N_53);
nand U871 (N_871,N_509,N_417);
or U872 (N_872,N_235,N_360);
nand U873 (N_873,N_251,N_24);
or U874 (N_874,N_269,N_558);
or U875 (N_875,N_581,N_287);
or U876 (N_876,N_376,N_517);
nand U877 (N_877,N_313,N_45);
nand U878 (N_878,N_55,N_268);
or U879 (N_879,N_465,N_106);
nand U880 (N_880,N_490,N_114);
or U881 (N_881,N_89,N_154);
and U882 (N_882,N_143,N_317);
nor U883 (N_883,N_421,N_575);
nor U884 (N_884,N_432,N_585);
nor U885 (N_885,N_533,N_138);
nand U886 (N_886,N_570,N_144);
or U887 (N_887,N_37,N_320);
nor U888 (N_888,N_100,N_547);
and U889 (N_889,N_249,N_257);
nor U890 (N_890,N_265,N_134);
nand U891 (N_891,N_571,N_577);
nor U892 (N_892,N_113,N_105);
or U893 (N_893,N_335,N_311);
nand U894 (N_894,N_291,N_152);
or U895 (N_895,N_248,N_466);
or U896 (N_896,N_125,N_400);
or U897 (N_897,N_521,N_528);
nand U898 (N_898,N_371,N_451);
or U899 (N_899,N_472,N_566);
nand U900 (N_900,N_313,N_386);
and U901 (N_901,N_313,N_542);
or U902 (N_902,N_385,N_564);
nor U903 (N_903,N_553,N_459);
nand U904 (N_904,N_303,N_170);
or U905 (N_905,N_282,N_89);
or U906 (N_906,N_271,N_566);
and U907 (N_907,N_293,N_118);
and U908 (N_908,N_295,N_405);
nand U909 (N_909,N_263,N_231);
or U910 (N_910,N_320,N_53);
nand U911 (N_911,N_92,N_154);
and U912 (N_912,N_169,N_512);
and U913 (N_913,N_471,N_85);
nand U914 (N_914,N_125,N_306);
nor U915 (N_915,N_145,N_528);
or U916 (N_916,N_340,N_213);
nor U917 (N_917,N_28,N_221);
or U918 (N_918,N_412,N_396);
nor U919 (N_919,N_96,N_10);
nand U920 (N_920,N_449,N_426);
or U921 (N_921,N_119,N_157);
and U922 (N_922,N_396,N_69);
nand U923 (N_923,N_333,N_546);
and U924 (N_924,N_257,N_20);
nand U925 (N_925,N_346,N_80);
nor U926 (N_926,N_567,N_288);
or U927 (N_927,N_186,N_407);
or U928 (N_928,N_518,N_136);
nand U929 (N_929,N_154,N_571);
or U930 (N_930,N_227,N_440);
and U931 (N_931,N_482,N_368);
or U932 (N_932,N_586,N_186);
and U933 (N_933,N_338,N_280);
nor U934 (N_934,N_202,N_297);
and U935 (N_935,N_151,N_104);
nor U936 (N_936,N_377,N_463);
and U937 (N_937,N_597,N_596);
nor U938 (N_938,N_230,N_288);
and U939 (N_939,N_441,N_237);
nand U940 (N_940,N_311,N_200);
and U941 (N_941,N_581,N_69);
and U942 (N_942,N_236,N_106);
and U943 (N_943,N_428,N_372);
nor U944 (N_944,N_287,N_275);
or U945 (N_945,N_276,N_109);
nor U946 (N_946,N_50,N_469);
and U947 (N_947,N_311,N_495);
nand U948 (N_948,N_427,N_162);
and U949 (N_949,N_481,N_54);
or U950 (N_950,N_47,N_596);
nand U951 (N_951,N_149,N_285);
and U952 (N_952,N_505,N_245);
nand U953 (N_953,N_170,N_110);
and U954 (N_954,N_140,N_528);
nand U955 (N_955,N_269,N_70);
or U956 (N_956,N_238,N_104);
nand U957 (N_957,N_94,N_319);
and U958 (N_958,N_293,N_504);
and U959 (N_959,N_557,N_247);
nor U960 (N_960,N_453,N_348);
nand U961 (N_961,N_59,N_189);
and U962 (N_962,N_320,N_55);
and U963 (N_963,N_460,N_408);
or U964 (N_964,N_498,N_518);
nand U965 (N_965,N_33,N_477);
nor U966 (N_966,N_288,N_99);
nor U967 (N_967,N_179,N_154);
or U968 (N_968,N_352,N_461);
or U969 (N_969,N_429,N_273);
and U970 (N_970,N_120,N_417);
and U971 (N_971,N_111,N_485);
nand U972 (N_972,N_150,N_15);
nand U973 (N_973,N_47,N_526);
nor U974 (N_974,N_582,N_545);
and U975 (N_975,N_551,N_295);
nand U976 (N_976,N_282,N_283);
nand U977 (N_977,N_555,N_2);
nor U978 (N_978,N_508,N_164);
or U979 (N_979,N_19,N_436);
nor U980 (N_980,N_396,N_516);
or U981 (N_981,N_276,N_131);
nor U982 (N_982,N_543,N_537);
or U983 (N_983,N_493,N_371);
nor U984 (N_984,N_463,N_506);
nor U985 (N_985,N_263,N_270);
xor U986 (N_986,N_452,N_72);
and U987 (N_987,N_22,N_305);
xnor U988 (N_988,N_473,N_555);
and U989 (N_989,N_139,N_267);
and U990 (N_990,N_483,N_98);
nor U991 (N_991,N_256,N_226);
nand U992 (N_992,N_7,N_305);
and U993 (N_993,N_213,N_337);
and U994 (N_994,N_456,N_262);
nand U995 (N_995,N_487,N_525);
or U996 (N_996,N_477,N_32);
nor U997 (N_997,N_198,N_296);
nand U998 (N_998,N_446,N_209);
or U999 (N_999,N_404,N_372);
nand U1000 (N_1000,N_114,N_250);
nand U1001 (N_1001,N_156,N_101);
or U1002 (N_1002,N_561,N_64);
nand U1003 (N_1003,N_225,N_443);
and U1004 (N_1004,N_460,N_175);
and U1005 (N_1005,N_33,N_490);
and U1006 (N_1006,N_552,N_284);
or U1007 (N_1007,N_417,N_441);
nand U1008 (N_1008,N_452,N_156);
nor U1009 (N_1009,N_344,N_393);
or U1010 (N_1010,N_360,N_595);
xnor U1011 (N_1011,N_120,N_463);
or U1012 (N_1012,N_94,N_260);
or U1013 (N_1013,N_183,N_426);
nand U1014 (N_1014,N_450,N_401);
nor U1015 (N_1015,N_441,N_61);
or U1016 (N_1016,N_542,N_254);
xor U1017 (N_1017,N_574,N_599);
and U1018 (N_1018,N_403,N_10);
or U1019 (N_1019,N_313,N_61);
nor U1020 (N_1020,N_593,N_106);
nand U1021 (N_1021,N_313,N_105);
nor U1022 (N_1022,N_95,N_545);
and U1023 (N_1023,N_263,N_219);
nand U1024 (N_1024,N_192,N_268);
nor U1025 (N_1025,N_194,N_80);
nand U1026 (N_1026,N_213,N_470);
or U1027 (N_1027,N_294,N_564);
and U1028 (N_1028,N_214,N_113);
or U1029 (N_1029,N_504,N_102);
or U1030 (N_1030,N_324,N_555);
nor U1031 (N_1031,N_179,N_248);
and U1032 (N_1032,N_71,N_98);
nand U1033 (N_1033,N_236,N_192);
or U1034 (N_1034,N_195,N_518);
or U1035 (N_1035,N_12,N_540);
nand U1036 (N_1036,N_425,N_241);
or U1037 (N_1037,N_381,N_472);
nor U1038 (N_1038,N_357,N_534);
or U1039 (N_1039,N_65,N_576);
or U1040 (N_1040,N_123,N_132);
and U1041 (N_1041,N_146,N_169);
xor U1042 (N_1042,N_243,N_90);
nor U1043 (N_1043,N_486,N_478);
nand U1044 (N_1044,N_190,N_82);
nor U1045 (N_1045,N_57,N_166);
nor U1046 (N_1046,N_527,N_29);
or U1047 (N_1047,N_539,N_550);
or U1048 (N_1048,N_458,N_548);
nand U1049 (N_1049,N_24,N_187);
nor U1050 (N_1050,N_200,N_568);
nand U1051 (N_1051,N_221,N_179);
and U1052 (N_1052,N_461,N_551);
or U1053 (N_1053,N_98,N_104);
nand U1054 (N_1054,N_284,N_37);
or U1055 (N_1055,N_323,N_512);
nand U1056 (N_1056,N_237,N_275);
and U1057 (N_1057,N_481,N_256);
nor U1058 (N_1058,N_429,N_286);
and U1059 (N_1059,N_154,N_597);
or U1060 (N_1060,N_235,N_346);
and U1061 (N_1061,N_0,N_26);
and U1062 (N_1062,N_216,N_381);
and U1063 (N_1063,N_308,N_126);
nor U1064 (N_1064,N_468,N_514);
or U1065 (N_1065,N_455,N_382);
or U1066 (N_1066,N_265,N_333);
and U1067 (N_1067,N_331,N_281);
nor U1068 (N_1068,N_493,N_445);
nor U1069 (N_1069,N_364,N_211);
nand U1070 (N_1070,N_126,N_263);
and U1071 (N_1071,N_226,N_291);
and U1072 (N_1072,N_464,N_509);
or U1073 (N_1073,N_443,N_384);
nand U1074 (N_1074,N_217,N_476);
nor U1075 (N_1075,N_371,N_116);
nor U1076 (N_1076,N_179,N_3);
nor U1077 (N_1077,N_33,N_29);
nor U1078 (N_1078,N_392,N_63);
nor U1079 (N_1079,N_100,N_348);
nor U1080 (N_1080,N_578,N_502);
nor U1081 (N_1081,N_36,N_514);
nor U1082 (N_1082,N_427,N_413);
or U1083 (N_1083,N_98,N_204);
or U1084 (N_1084,N_366,N_287);
or U1085 (N_1085,N_561,N_114);
and U1086 (N_1086,N_402,N_535);
or U1087 (N_1087,N_444,N_505);
and U1088 (N_1088,N_482,N_227);
nand U1089 (N_1089,N_440,N_267);
nor U1090 (N_1090,N_139,N_215);
and U1091 (N_1091,N_120,N_450);
or U1092 (N_1092,N_269,N_402);
nand U1093 (N_1093,N_313,N_152);
or U1094 (N_1094,N_456,N_540);
nand U1095 (N_1095,N_339,N_550);
and U1096 (N_1096,N_493,N_590);
nor U1097 (N_1097,N_454,N_7);
and U1098 (N_1098,N_388,N_502);
or U1099 (N_1099,N_57,N_486);
or U1100 (N_1100,N_464,N_189);
nor U1101 (N_1101,N_543,N_334);
nand U1102 (N_1102,N_98,N_377);
and U1103 (N_1103,N_119,N_537);
or U1104 (N_1104,N_344,N_58);
nand U1105 (N_1105,N_324,N_438);
nand U1106 (N_1106,N_227,N_358);
nand U1107 (N_1107,N_40,N_5);
or U1108 (N_1108,N_569,N_173);
nand U1109 (N_1109,N_9,N_378);
nor U1110 (N_1110,N_16,N_92);
nor U1111 (N_1111,N_18,N_259);
or U1112 (N_1112,N_109,N_561);
nor U1113 (N_1113,N_412,N_289);
or U1114 (N_1114,N_550,N_464);
and U1115 (N_1115,N_496,N_449);
nor U1116 (N_1116,N_561,N_212);
and U1117 (N_1117,N_230,N_55);
or U1118 (N_1118,N_78,N_378);
nor U1119 (N_1119,N_138,N_206);
nand U1120 (N_1120,N_518,N_334);
or U1121 (N_1121,N_599,N_142);
nor U1122 (N_1122,N_113,N_182);
and U1123 (N_1123,N_237,N_163);
nor U1124 (N_1124,N_399,N_395);
or U1125 (N_1125,N_224,N_382);
and U1126 (N_1126,N_426,N_372);
and U1127 (N_1127,N_29,N_187);
or U1128 (N_1128,N_28,N_476);
and U1129 (N_1129,N_331,N_443);
nand U1130 (N_1130,N_529,N_321);
nand U1131 (N_1131,N_413,N_583);
or U1132 (N_1132,N_480,N_525);
nand U1133 (N_1133,N_167,N_300);
and U1134 (N_1134,N_103,N_527);
nor U1135 (N_1135,N_369,N_349);
or U1136 (N_1136,N_2,N_271);
nand U1137 (N_1137,N_596,N_534);
nor U1138 (N_1138,N_430,N_28);
and U1139 (N_1139,N_102,N_314);
and U1140 (N_1140,N_61,N_28);
nand U1141 (N_1141,N_592,N_350);
or U1142 (N_1142,N_424,N_510);
or U1143 (N_1143,N_262,N_72);
nor U1144 (N_1144,N_362,N_394);
nor U1145 (N_1145,N_535,N_99);
nor U1146 (N_1146,N_538,N_137);
nand U1147 (N_1147,N_92,N_311);
nor U1148 (N_1148,N_563,N_425);
nand U1149 (N_1149,N_84,N_115);
nand U1150 (N_1150,N_291,N_279);
nor U1151 (N_1151,N_501,N_526);
nor U1152 (N_1152,N_272,N_414);
or U1153 (N_1153,N_228,N_269);
nor U1154 (N_1154,N_447,N_583);
nor U1155 (N_1155,N_288,N_576);
or U1156 (N_1156,N_173,N_493);
nand U1157 (N_1157,N_219,N_157);
and U1158 (N_1158,N_504,N_166);
or U1159 (N_1159,N_462,N_26);
nor U1160 (N_1160,N_249,N_324);
or U1161 (N_1161,N_123,N_259);
nor U1162 (N_1162,N_15,N_79);
nor U1163 (N_1163,N_85,N_597);
nand U1164 (N_1164,N_138,N_335);
or U1165 (N_1165,N_508,N_557);
nor U1166 (N_1166,N_88,N_93);
or U1167 (N_1167,N_200,N_399);
and U1168 (N_1168,N_140,N_453);
and U1169 (N_1169,N_462,N_586);
and U1170 (N_1170,N_359,N_164);
nor U1171 (N_1171,N_154,N_517);
or U1172 (N_1172,N_343,N_441);
nand U1173 (N_1173,N_264,N_311);
and U1174 (N_1174,N_195,N_440);
or U1175 (N_1175,N_244,N_510);
and U1176 (N_1176,N_343,N_3);
or U1177 (N_1177,N_591,N_113);
or U1178 (N_1178,N_359,N_541);
nor U1179 (N_1179,N_561,N_160);
nand U1180 (N_1180,N_98,N_525);
nand U1181 (N_1181,N_353,N_283);
nor U1182 (N_1182,N_14,N_390);
nor U1183 (N_1183,N_574,N_316);
or U1184 (N_1184,N_132,N_542);
and U1185 (N_1185,N_217,N_420);
or U1186 (N_1186,N_128,N_240);
or U1187 (N_1187,N_450,N_94);
or U1188 (N_1188,N_121,N_303);
nand U1189 (N_1189,N_227,N_510);
or U1190 (N_1190,N_596,N_429);
or U1191 (N_1191,N_301,N_327);
nor U1192 (N_1192,N_2,N_111);
and U1193 (N_1193,N_31,N_527);
nor U1194 (N_1194,N_49,N_533);
and U1195 (N_1195,N_151,N_180);
nand U1196 (N_1196,N_16,N_292);
nor U1197 (N_1197,N_49,N_399);
nor U1198 (N_1198,N_316,N_511);
and U1199 (N_1199,N_144,N_320);
nand U1200 (N_1200,N_955,N_761);
nand U1201 (N_1201,N_953,N_1096);
nand U1202 (N_1202,N_1183,N_1196);
or U1203 (N_1203,N_898,N_1065);
and U1204 (N_1204,N_695,N_704);
and U1205 (N_1205,N_1166,N_684);
and U1206 (N_1206,N_832,N_1095);
nand U1207 (N_1207,N_1146,N_874);
nand U1208 (N_1208,N_852,N_1014);
or U1209 (N_1209,N_778,N_970);
nor U1210 (N_1210,N_998,N_893);
nor U1211 (N_1211,N_933,N_733);
nand U1212 (N_1212,N_697,N_908);
or U1213 (N_1213,N_653,N_1160);
and U1214 (N_1214,N_828,N_1163);
and U1215 (N_1215,N_948,N_1091);
nor U1216 (N_1216,N_631,N_782);
or U1217 (N_1217,N_865,N_1104);
and U1218 (N_1218,N_1083,N_706);
nor U1219 (N_1219,N_714,N_1126);
or U1220 (N_1220,N_651,N_1124);
and U1221 (N_1221,N_1022,N_793);
nand U1222 (N_1222,N_637,N_1165);
or U1223 (N_1223,N_947,N_765);
nor U1224 (N_1224,N_996,N_649);
and U1225 (N_1225,N_1050,N_1079);
nor U1226 (N_1226,N_785,N_1120);
or U1227 (N_1227,N_875,N_892);
or U1228 (N_1228,N_1142,N_784);
nor U1229 (N_1229,N_731,N_963);
nor U1230 (N_1230,N_1094,N_889);
and U1231 (N_1231,N_909,N_1038);
or U1232 (N_1232,N_1167,N_1198);
or U1233 (N_1233,N_1059,N_1036);
nand U1234 (N_1234,N_879,N_999);
nand U1235 (N_1235,N_757,N_853);
nand U1236 (N_1236,N_610,N_701);
or U1237 (N_1237,N_717,N_827);
or U1238 (N_1238,N_788,N_972);
or U1239 (N_1239,N_973,N_1074);
nand U1240 (N_1240,N_762,N_1180);
nor U1241 (N_1241,N_1129,N_635);
and U1242 (N_1242,N_1153,N_1128);
or U1243 (N_1243,N_664,N_661);
and U1244 (N_1244,N_862,N_692);
or U1245 (N_1245,N_900,N_927);
or U1246 (N_1246,N_1093,N_1009);
nor U1247 (N_1247,N_801,N_691);
and U1248 (N_1248,N_1181,N_1134);
or U1249 (N_1249,N_1087,N_794);
nand U1250 (N_1250,N_698,N_677);
nand U1251 (N_1251,N_1067,N_759);
nand U1252 (N_1252,N_1112,N_887);
nor U1253 (N_1253,N_650,N_858);
nand U1254 (N_1254,N_670,N_622);
nor U1255 (N_1255,N_1184,N_1194);
and U1256 (N_1256,N_643,N_819);
nand U1257 (N_1257,N_781,N_1044);
or U1258 (N_1258,N_660,N_825);
nor U1259 (N_1259,N_768,N_730);
nor U1260 (N_1260,N_659,N_620);
and U1261 (N_1261,N_1043,N_1188);
nor U1262 (N_1262,N_837,N_954);
and U1263 (N_1263,N_1187,N_876);
and U1264 (N_1264,N_810,N_1136);
nand U1265 (N_1265,N_872,N_1131);
xor U1266 (N_1266,N_1052,N_713);
nand U1267 (N_1267,N_1192,N_878);
or U1268 (N_1268,N_811,N_974);
nand U1269 (N_1269,N_814,N_1001);
nor U1270 (N_1270,N_686,N_1016);
or U1271 (N_1271,N_743,N_1049);
xnor U1272 (N_1272,N_1057,N_772);
and U1273 (N_1273,N_997,N_803);
nand U1274 (N_1274,N_940,N_1173);
nand U1275 (N_1275,N_729,N_756);
or U1276 (N_1276,N_1199,N_1042);
nand U1277 (N_1277,N_1141,N_726);
nand U1278 (N_1278,N_978,N_669);
or U1279 (N_1279,N_930,N_735);
or U1280 (N_1280,N_616,N_849);
and U1281 (N_1281,N_1062,N_1070);
nand U1282 (N_1282,N_682,N_945);
or U1283 (N_1283,N_942,N_1168);
nand U1284 (N_1284,N_877,N_894);
nor U1285 (N_1285,N_831,N_617);
nor U1286 (N_1286,N_979,N_964);
and U1287 (N_1287,N_1013,N_612);
or U1288 (N_1288,N_817,N_1021);
nor U1289 (N_1289,N_615,N_1040);
nor U1290 (N_1290,N_621,N_609);
nand U1291 (N_1291,N_962,N_1089);
nor U1292 (N_1292,N_1018,N_640);
nand U1293 (N_1293,N_1078,N_1086);
or U1294 (N_1294,N_1024,N_604);
nand U1295 (N_1295,N_806,N_611);
xor U1296 (N_1296,N_1159,N_1020);
nor U1297 (N_1297,N_1154,N_952);
or U1298 (N_1298,N_987,N_624);
and U1299 (N_1299,N_1017,N_843);
and U1300 (N_1300,N_995,N_917);
xor U1301 (N_1301,N_606,N_1008);
and U1302 (N_1302,N_1101,N_671);
nand U1303 (N_1303,N_1063,N_1152);
nand U1304 (N_1304,N_712,N_725);
nor U1305 (N_1305,N_993,N_656);
or U1306 (N_1306,N_923,N_925);
and U1307 (N_1307,N_949,N_1138);
or U1308 (N_1308,N_738,N_1125);
nor U1309 (N_1309,N_1190,N_668);
nor U1310 (N_1310,N_657,N_935);
nand U1311 (N_1311,N_1097,N_944);
and U1312 (N_1312,N_899,N_773);
nor U1313 (N_1313,N_746,N_914);
nand U1314 (N_1314,N_626,N_1121);
and U1315 (N_1315,N_1133,N_1143);
nand U1316 (N_1316,N_859,N_1003);
or U1317 (N_1317,N_1130,N_1127);
nor U1318 (N_1318,N_797,N_848);
or U1319 (N_1319,N_745,N_702);
and U1320 (N_1320,N_834,N_981);
or U1321 (N_1321,N_1108,N_1045);
and U1322 (N_1322,N_946,N_603);
or U1323 (N_1323,N_1041,N_928);
nand U1324 (N_1324,N_913,N_992);
xnor U1325 (N_1325,N_957,N_646);
nor U1326 (N_1326,N_1118,N_775);
or U1327 (N_1327,N_1186,N_880);
or U1328 (N_1328,N_911,N_699);
and U1329 (N_1329,N_1178,N_1034);
and U1330 (N_1330,N_783,N_690);
nand U1331 (N_1331,N_1002,N_1117);
or U1332 (N_1332,N_990,N_847);
and U1333 (N_1333,N_984,N_627);
nand U1334 (N_1334,N_904,N_685);
nand U1335 (N_1335,N_939,N_1077);
or U1336 (N_1336,N_618,N_1053);
nor U1337 (N_1337,N_1195,N_1135);
nand U1338 (N_1338,N_816,N_798);
nand U1339 (N_1339,N_753,N_679);
or U1340 (N_1340,N_766,N_1072);
nor U1341 (N_1341,N_951,N_840);
and U1342 (N_1342,N_857,N_1028);
and U1343 (N_1343,N_1122,N_958);
nor U1344 (N_1344,N_829,N_1076);
and U1345 (N_1345,N_718,N_683);
and U1346 (N_1346,N_655,N_960);
nor U1347 (N_1347,N_632,N_1189);
nand U1348 (N_1348,N_749,N_719);
nor U1349 (N_1349,N_915,N_737);
or U1350 (N_1350,N_771,N_804);
nand U1351 (N_1351,N_1106,N_823);
and U1352 (N_1352,N_1007,N_1177);
nand U1353 (N_1353,N_1137,N_774);
nor U1354 (N_1354,N_967,N_1000);
and U1355 (N_1355,N_634,N_977);
or U1356 (N_1356,N_918,N_1010);
nor U1357 (N_1357,N_807,N_689);
and U1358 (N_1358,N_1157,N_1026);
xor U1359 (N_1359,N_851,N_1098);
and U1360 (N_1360,N_906,N_1164);
nor U1361 (N_1361,N_675,N_826);
or U1362 (N_1362,N_1169,N_868);
nand U1363 (N_1363,N_1100,N_1033);
and U1364 (N_1364,N_739,N_786);
and U1365 (N_1365,N_813,N_1035);
nand U1366 (N_1366,N_1174,N_763);
nor U1367 (N_1367,N_716,N_922);
nor U1368 (N_1368,N_934,N_777);
or U1369 (N_1369,N_959,N_787);
nand U1370 (N_1370,N_924,N_792);
or U1371 (N_1371,N_854,N_869);
or U1372 (N_1372,N_950,N_1139);
and U1373 (N_1373,N_1051,N_976);
and U1374 (N_1374,N_1176,N_790);
and U1375 (N_1375,N_600,N_883);
nand U1376 (N_1376,N_1155,N_1030);
nand U1377 (N_1377,N_750,N_1114);
nor U1378 (N_1378,N_938,N_932);
nor U1379 (N_1379,N_1069,N_985);
nor U1380 (N_1380,N_644,N_921);
and U1381 (N_1381,N_1175,N_916);
nor U1382 (N_1382,N_1032,N_665);
and U1383 (N_1383,N_890,N_715);
and U1384 (N_1384,N_1088,N_795);
or U1385 (N_1385,N_855,N_1081);
xnor U1386 (N_1386,N_989,N_838);
nand U1387 (N_1387,N_1193,N_667);
nor U1388 (N_1388,N_870,N_1172);
nand U1389 (N_1389,N_1113,N_645);
nand U1390 (N_1390,N_796,N_666);
or U1391 (N_1391,N_920,N_866);
nor U1392 (N_1392,N_1099,N_639);
nand U1393 (N_1393,N_986,N_1054);
nor U1394 (N_1394,N_1185,N_727);
and U1395 (N_1395,N_732,N_882);
and U1396 (N_1396,N_791,N_1151);
nand U1397 (N_1397,N_888,N_1111);
nand U1398 (N_1398,N_780,N_802);
or U1399 (N_1399,N_647,N_605);
and U1400 (N_1400,N_980,N_710);
or U1401 (N_1401,N_1132,N_630);
xnor U1402 (N_1402,N_1068,N_754);
nand U1403 (N_1403,N_864,N_1055);
nor U1404 (N_1404,N_1197,N_895);
nand U1405 (N_1405,N_601,N_1161);
nand U1406 (N_1406,N_1075,N_943);
and U1407 (N_1407,N_681,N_789);
nand U1408 (N_1408,N_672,N_742);
nor U1409 (N_1409,N_613,N_1092);
or U1410 (N_1410,N_720,N_1046);
nand U1411 (N_1411,N_1056,N_1023);
or U1412 (N_1412,N_805,N_641);
nor U1413 (N_1413,N_711,N_1148);
or U1414 (N_1414,N_770,N_931);
nand U1415 (N_1415,N_1012,N_994);
nand U1416 (N_1416,N_619,N_891);
or U1417 (N_1417,N_901,N_1039);
and U1418 (N_1418,N_723,N_736);
nor U1419 (N_1419,N_968,N_969);
nor U1420 (N_1420,N_982,N_636);
and U1421 (N_1421,N_856,N_815);
nor U1422 (N_1422,N_863,N_1085);
and U1423 (N_1423,N_760,N_693);
nand U1424 (N_1424,N_747,N_991);
and U1425 (N_1425,N_1029,N_642);
and U1426 (N_1426,N_841,N_734);
and U1427 (N_1427,N_965,N_799);
and U1428 (N_1428,N_873,N_809);
and U1429 (N_1429,N_1162,N_1109);
and U1430 (N_1430,N_721,N_897);
nand U1431 (N_1431,N_673,N_839);
or U1432 (N_1432,N_929,N_678);
or U1433 (N_1433,N_842,N_755);
and U1434 (N_1434,N_680,N_1082);
and U1435 (N_1435,N_674,N_1058);
or U1436 (N_1436,N_1080,N_936);
nand U1437 (N_1437,N_687,N_1060);
or U1438 (N_1438,N_1144,N_836);
or U1439 (N_1439,N_662,N_971);
or U1440 (N_1440,N_941,N_1156);
and U1441 (N_1441,N_709,N_1084);
nand U1442 (N_1442,N_966,N_676);
nor U1443 (N_1443,N_1171,N_845);
nor U1444 (N_1444,N_744,N_818);
nor U1445 (N_1445,N_1047,N_975);
and U1446 (N_1446,N_1145,N_912);
nor U1447 (N_1447,N_1090,N_1147);
nand U1448 (N_1448,N_722,N_779);
nand U1449 (N_1449,N_752,N_625);
and U1450 (N_1450,N_767,N_1191);
nand U1451 (N_1451,N_886,N_1011);
nand U1452 (N_1452,N_688,N_1179);
and U1453 (N_1453,N_919,N_1105);
nor U1454 (N_1454,N_820,N_1027);
nand U1455 (N_1455,N_902,N_764);
nor U1456 (N_1456,N_821,N_881);
nand U1457 (N_1457,N_700,N_1005);
or U1458 (N_1458,N_769,N_988);
and U1459 (N_1459,N_758,N_741);
nor U1460 (N_1460,N_808,N_1158);
nor U1461 (N_1461,N_812,N_1066);
nor U1462 (N_1462,N_956,N_833);
nor U1463 (N_1463,N_696,N_844);
and U1464 (N_1464,N_1119,N_867);
nor U1465 (N_1465,N_652,N_623);
xor U1466 (N_1466,N_884,N_1103);
nand U1467 (N_1467,N_608,N_703);
nand U1468 (N_1468,N_1110,N_1071);
and U1469 (N_1469,N_707,N_1107);
nor U1470 (N_1470,N_860,N_1061);
or U1471 (N_1471,N_648,N_926);
or U1472 (N_1472,N_1015,N_830);
or U1473 (N_1473,N_1115,N_937);
and U1474 (N_1474,N_694,N_740);
and U1475 (N_1475,N_751,N_961);
or U1476 (N_1476,N_708,N_607);
nand U1477 (N_1477,N_1150,N_983);
nor U1478 (N_1478,N_776,N_896);
nor U1479 (N_1479,N_658,N_629);
nor U1480 (N_1480,N_903,N_822);
or U1481 (N_1481,N_910,N_1064);
nor U1482 (N_1482,N_905,N_835);
or U1483 (N_1483,N_1037,N_1006);
nor U1484 (N_1484,N_824,N_654);
xor U1485 (N_1485,N_628,N_885);
or U1486 (N_1486,N_1031,N_614);
nor U1487 (N_1487,N_1140,N_1019);
and U1488 (N_1488,N_1048,N_1073);
nand U1489 (N_1489,N_861,N_602);
nand U1490 (N_1490,N_1004,N_663);
nor U1491 (N_1491,N_871,N_1116);
or U1492 (N_1492,N_1182,N_1102);
nand U1493 (N_1493,N_1149,N_724);
nor U1494 (N_1494,N_907,N_846);
nor U1495 (N_1495,N_638,N_748);
or U1496 (N_1496,N_1123,N_850);
nand U1497 (N_1497,N_1025,N_705);
nand U1498 (N_1498,N_1170,N_728);
xnor U1499 (N_1499,N_633,N_800);
or U1500 (N_1500,N_620,N_1181);
nand U1501 (N_1501,N_867,N_874);
nand U1502 (N_1502,N_775,N_979);
nand U1503 (N_1503,N_613,N_1152);
xor U1504 (N_1504,N_974,N_655);
or U1505 (N_1505,N_604,N_1160);
or U1506 (N_1506,N_938,N_661);
xnor U1507 (N_1507,N_706,N_983);
nor U1508 (N_1508,N_1038,N_1196);
and U1509 (N_1509,N_839,N_640);
nand U1510 (N_1510,N_1077,N_1118);
and U1511 (N_1511,N_772,N_919);
nand U1512 (N_1512,N_1065,N_968);
or U1513 (N_1513,N_954,N_960);
and U1514 (N_1514,N_619,N_1072);
nor U1515 (N_1515,N_754,N_664);
nor U1516 (N_1516,N_715,N_708);
and U1517 (N_1517,N_1073,N_1134);
and U1518 (N_1518,N_788,N_1088);
nor U1519 (N_1519,N_671,N_913);
nor U1520 (N_1520,N_997,N_1065);
nand U1521 (N_1521,N_675,N_886);
nor U1522 (N_1522,N_1127,N_666);
nor U1523 (N_1523,N_643,N_650);
nand U1524 (N_1524,N_646,N_912);
and U1525 (N_1525,N_697,N_1135);
nand U1526 (N_1526,N_1075,N_845);
and U1527 (N_1527,N_635,N_831);
nor U1528 (N_1528,N_1138,N_942);
nand U1529 (N_1529,N_690,N_923);
nor U1530 (N_1530,N_958,N_694);
nor U1531 (N_1531,N_1007,N_1154);
nand U1532 (N_1532,N_812,N_901);
and U1533 (N_1533,N_1167,N_944);
and U1534 (N_1534,N_872,N_1181);
nand U1535 (N_1535,N_756,N_712);
or U1536 (N_1536,N_919,N_671);
and U1537 (N_1537,N_987,N_628);
or U1538 (N_1538,N_963,N_763);
nand U1539 (N_1539,N_948,N_634);
nand U1540 (N_1540,N_794,N_715);
and U1541 (N_1541,N_965,N_1020);
nand U1542 (N_1542,N_1009,N_623);
or U1543 (N_1543,N_1107,N_1027);
and U1544 (N_1544,N_822,N_919);
or U1545 (N_1545,N_942,N_944);
nand U1546 (N_1546,N_820,N_950);
nand U1547 (N_1547,N_965,N_1118);
nand U1548 (N_1548,N_767,N_1163);
and U1549 (N_1549,N_947,N_966);
nor U1550 (N_1550,N_1133,N_655);
nor U1551 (N_1551,N_850,N_1035);
and U1552 (N_1552,N_831,N_1060);
nor U1553 (N_1553,N_1189,N_1080);
nand U1554 (N_1554,N_1151,N_800);
nor U1555 (N_1555,N_822,N_1094);
or U1556 (N_1556,N_990,N_673);
nand U1557 (N_1557,N_1043,N_1194);
and U1558 (N_1558,N_740,N_1088);
or U1559 (N_1559,N_1026,N_1110);
nand U1560 (N_1560,N_609,N_603);
and U1561 (N_1561,N_853,N_694);
or U1562 (N_1562,N_937,N_600);
or U1563 (N_1563,N_839,N_610);
or U1564 (N_1564,N_702,N_657);
and U1565 (N_1565,N_717,N_1177);
nor U1566 (N_1566,N_826,N_763);
or U1567 (N_1567,N_855,N_846);
nand U1568 (N_1568,N_1121,N_918);
nor U1569 (N_1569,N_693,N_858);
and U1570 (N_1570,N_1124,N_683);
and U1571 (N_1571,N_908,N_1018);
or U1572 (N_1572,N_1051,N_876);
and U1573 (N_1573,N_745,N_969);
nand U1574 (N_1574,N_964,N_1140);
xor U1575 (N_1575,N_1053,N_907);
xnor U1576 (N_1576,N_1004,N_684);
and U1577 (N_1577,N_983,N_918);
or U1578 (N_1578,N_611,N_864);
and U1579 (N_1579,N_983,N_887);
or U1580 (N_1580,N_975,N_842);
nor U1581 (N_1581,N_1035,N_899);
or U1582 (N_1582,N_694,N_663);
nand U1583 (N_1583,N_767,N_1028);
or U1584 (N_1584,N_900,N_835);
or U1585 (N_1585,N_1132,N_1073);
nand U1586 (N_1586,N_664,N_1176);
nor U1587 (N_1587,N_600,N_1014);
or U1588 (N_1588,N_947,N_1074);
nor U1589 (N_1589,N_628,N_823);
xor U1590 (N_1590,N_649,N_818);
nor U1591 (N_1591,N_813,N_752);
and U1592 (N_1592,N_992,N_880);
or U1593 (N_1593,N_807,N_978);
nor U1594 (N_1594,N_1163,N_943);
and U1595 (N_1595,N_1183,N_696);
nand U1596 (N_1596,N_770,N_1073);
nor U1597 (N_1597,N_850,N_799);
nor U1598 (N_1598,N_1099,N_1151);
nand U1599 (N_1599,N_1115,N_914);
nor U1600 (N_1600,N_1071,N_963);
and U1601 (N_1601,N_767,N_1175);
xnor U1602 (N_1602,N_1149,N_1095);
and U1603 (N_1603,N_729,N_1050);
or U1604 (N_1604,N_725,N_826);
and U1605 (N_1605,N_1160,N_839);
nor U1606 (N_1606,N_1106,N_744);
nor U1607 (N_1607,N_846,N_925);
nor U1608 (N_1608,N_767,N_732);
or U1609 (N_1609,N_737,N_856);
or U1610 (N_1610,N_630,N_798);
nor U1611 (N_1611,N_975,N_1137);
nand U1612 (N_1612,N_1047,N_953);
or U1613 (N_1613,N_609,N_684);
and U1614 (N_1614,N_1094,N_749);
and U1615 (N_1615,N_827,N_771);
nor U1616 (N_1616,N_965,N_1053);
nand U1617 (N_1617,N_603,N_652);
and U1618 (N_1618,N_997,N_1132);
and U1619 (N_1619,N_1080,N_1061);
and U1620 (N_1620,N_1053,N_1096);
or U1621 (N_1621,N_1125,N_754);
nand U1622 (N_1622,N_772,N_624);
or U1623 (N_1623,N_724,N_1142);
or U1624 (N_1624,N_917,N_632);
or U1625 (N_1625,N_624,N_1134);
nor U1626 (N_1626,N_613,N_925);
and U1627 (N_1627,N_1192,N_639);
and U1628 (N_1628,N_786,N_689);
nor U1629 (N_1629,N_752,N_884);
or U1630 (N_1630,N_965,N_817);
or U1631 (N_1631,N_642,N_1164);
nor U1632 (N_1632,N_812,N_1147);
nor U1633 (N_1633,N_1163,N_626);
xnor U1634 (N_1634,N_767,N_916);
and U1635 (N_1635,N_824,N_855);
or U1636 (N_1636,N_707,N_872);
nor U1637 (N_1637,N_817,N_809);
or U1638 (N_1638,N_942,N_1153);
or U1639 (N_1639,N_973,N_741);
and U1640 (N_1640,N_1058,N_879);
and U1641 (N_1641,N_732,N_1135);
or U1642 (N_1642,N_1199,N_1154);
nor U1643 (N_1643,N_1072,N_604);
or U1644 (N_1644,N_1140,N_1046);
nor U1645 (N_1645,N_922,N_906);
and U1646 (N_1646,N_1160,N_1083);
or U1647 (N_1647,N_797,N_760);
or U1648 (N_1648,N_713,N_845);
nor U1649 (N_1649,N_644,N_741);
and U1650 (N_1650,N_861,N_678);
nand U1651 (N_1651,N_974,N_653);
nand U1652 (N_1652,N_1115,N_652);
nand U1653 (N_1653,N_1156,N_1128);
and U1654 (N_1654,N_908,N_1115);
nor U1655 (N_1655,N_995,N_647);
or U1656 (N_1656,N_1136,N_1057);
or U1657 (N_1657,N_868,N_889);
nor U1658 (N_1658,N_644,N_1191);
and U1659 (N_1659,N_1129,N_754);
nand U1660 (N_1660,N_972,N_727);
nor U1661 (N_1661,N_818,N_1077);
and U1662 (N_1662,N_691,N_960);
or U1663 (N_1663,N_862,N_1101);
and U1664 (N_1664,N_858,N_918);
or U1665 (N_1665,N_909,N_876);
nor U1666 (N_1666,N_1162,N_636);
nand U1667 (N_1667,N_672,N_1188);
nand U1668 (N_1668,N_898,N_1106);
or U1669 (N_1669,N_958,N_1020);
or U1670 (N_1670,N_1066,N_712);
nand U1671 (N_1671,N_1065,N_863);
and U1672 (N_1672,N_881,N_827);
and U1673 (N_1673,N_672,N_767);
nand U1674 (N_1674,N_714,N_1119);
or U1675 (N_1675,N_932,N_1087);
nor U1676 (N_1676,N_608,N_1184);
nand U1677 (N_1677,N_869,N_798);
or U1678 (N_1678,N_921,N_1131);
or U1679 (N_1679,N_926,N_884);
and U1680 (N_1680,N_950,N_1137);
nand U1681 (N_1681,N_785,N_838);
nand U1682 (N_1682,N_750,N_625);
or U1683 (N_1683,N_1102,N_910);
and U1684 (N_1684,N_879,N_663);
and U1685 (N_1685,N_748,N_787);
nand U1686 (N_1686,N_695,N_850);
nand U1687 (N_1687,N_1053,N_1055);
nand U1688 (N_1688,N_877,N_1057);
nand U1689 (N_1689,N_674,N_1129);
nor U1690 (N_1690,N_1025,N_1076);
and U1691 (N_1691,N_804,N_698);
or U1692 (N_1692,N_946,N_887);
nor U1693 (N_1693,N_703,N_1072);
nand U1694 (N_1694,N_620,N_910);
nor U1695 (N_1695,N_790,N_747);
or U1696 (N_1696,N_1067,N_856);
and U1697 (N_1697,N_1070,N_1064);
nor U1698 (N_1698,N_1039,N_1158);
nor U1699 (N_1699,N_637,N_616);
nor U1700 (N_1700,N_1042,N_1038);
nand U1701 (N_1701,N_1035,N_775);
and U1702 (N_1702,N_1147,N_1125);
nor U1703 (N_1703,N_661,N_1109);
or U1704 (N_1704,N_954,N_1131);
or U1705 (N_1705,N_1015,N_817);
nand U1706 (N_1706,N_1002,N_867);
and U1707 (N_1707,N_820,N_873);
nand U1708 (N_1708,N_1148,N_997);
or U1709 (N_1709,N_1008,N_836);
nor U1710 (N_1710,N_1143,N_1104);
or U1711 (N_1711,N_739,N_690);
nand U1712 (N_1712,N_1005,N_1185);
nand U1713 (N_1713,N_1074,N_812);
nand U1714 (N_1714,N_1190,N_1030);
and U1715 (N_1715,N_1160,N_1037);
or U1716 (N_1716,N_618,N_880);
nor U1717 (N_1717,N_1107,N_652);
nor U1718 (N_1718,N_763,N_958);
nand U1719 (N_1719,N_893,N_634);
and U1720 (N_1720,N_685,N_858);
nor U1721 (N_1721,N_701,N_771);
and U1722 (N_1722,N_999,N_1158);
and U1723 (N_1723,N_848,N_1075);
and U1724 (N_1724,N_860,N_1065);
nor U1725 (N_1725,N_1050,N_1100);
and U1726 (N_1726,N_1039,N_769);
and U1727 (N_1727,N_693,N_802);
and U1728 (N_1728,N_742,N_804);
nand U1729 (N_1729,N_858,N_867);
nand U1730 (N_1730,N_987,N_672);
nand U1731 (N_1731,N_1154,N_842);
nor U1732 (N_1732,N_926,N_763);
or U1733 (N_1733,N_782,N_1159);
nand U1734 (N_1734,N_1131,N_1082);
and U1735 (N_1735,N_676,N_845);
and U1736 (N_1736,N_957,N_999);
nor U1737 (N_1737,N_800,N_859);
and U1738 (N_1738,N_1006,N_658);
nor U1739 (N_1739,N_1191,N_902);
or U1740 (N_1740,N_961,N_987);
xnor U1741 (N_1741,N_834,N_815);
and U1742 (N_1742,N_775,N_797);
and U1743 (N_1743,N_827,N_1091);
or U1744 (N_1744,N_753,N_736);
or U1745 (N_1745,N_783,N_808);
nand U1746 (N_1746,N_953,N_849);
nand U1747 (N_1747,N_1100,N_807);
or U1748 (N_1748,N_1103,N_1009);
and U1749 (N_1749,N_709,N_931);
nand U1750 (N_1750,N_878,N_843);
and U1751 (N_1751,N_858,N_957);
nand U1752 (N_1752,N_808,N_723);
nor U1753 (N_1753,N_1153,N_783);
or U1754 (N_1754,N_849,N_1117);
nand U1755 (N_1755,N_848,N_647);
or U1756 (N_1756,N_1125,N_1094);
and U1757 (N_1757,N_737,N_992);
nand U1758 (N_1758,N_784,N_968);
nor U1759 (N_1759,N_765,N_1153);
nand U1760 (N_1760,N_615,N_854);
or U1761 (N_1761,N_1126,N_757);
nor U1762 (N_1762,N_808,N_788);
nand U1763 (N_1763,N_957,N_886);
and U1764 (N_1764,N_1153,N_613);
and U1765 (N_1765,N_904,N_693);
or U1766 (N_1766,N_876,N_650);
nor U1767 (N_1767,N_876,N_974);
or U1768 (N_1768,N_654,N_642);
nand U1769 (N_1769,N_1141,N_727);
or U1770 (N_1770,N_1057,N_1133);
or U1771 (N_1771,N_967,N_623);
nor U1772 (N_1772,N_970,N_1039);
nor U1773 (N_1773,N_842,N_1037);
or U1774 (N_1774,N_1161,N_807);
and U1775 (N_1775,N_1138,N_832);
nor U1776 (N_1776,N_710,N_608);
nor U1777 (N_1777,N_686,N_903);
and U1778 (N_1778,N_873,N_1177);
and U1779 (N_1779,N_841,N_902);
nand U1780 (N_1780,N_899,N_864);
nand U1781 (N_1781,N_652,N_840);
nor U1782 (N_1782,N_733,N_621);
nor U1783 (N_1783,N_710,N_1122);
or U1784 (N_1784,N_1031,N_751);
nand U1785 (N_1785,N_1058,N_895);
nand U1786 (N_1786,N_720,N_1017);
nand U1787 (N_1787,N_984,N_1063);
nand U1788 (N_1788,N_620,N_830);
and U1789 (N_1789,N_1161,N_876);
nand U1790 (N_1790,N_751,N_795);
nand U1791 (N_1791,N_1029,N_836);
nand U1792 (N_1792,N_652,N_917);
nor U1793 (N_1793,N_1072,N_1144);
nor U1794 (N_1794,N_1139,N_627);
nor U1795 (N_1795,N_692,N_849);
and U1796 (N_1796,N_798,N_633);
nand U1797 (N_1797,N_803,N_956);
or U1798 (N_1798,N_754,N_1138);
and U1799 (N_1799,N_786,N_775);
nand U1800 (N_1800,N_1797,N_1303);
nor U1801 (N_1801,N_1446,N_1238);
nor U1802 (N_1802,N_1656,N_1706);
nor U1803 (N_1803,N_1421,N_1348);
and U1804 (N_1804,N_1464,N_1697);
nand U1805 (N_1805,N_1448,N_1372);
or U1806 (N_1806,N_1444,N_1544);
or U1807 (N_1807,N_1423,N_1213);
nor U1808 (N_1808,N_1300,N_1312);
or U1809 (N_1809,N_1595,N_1395);
and U1810 (N_1810,N_1385,N_1799);
nor U1811 (N_1811,N_1521,N_1618);
or U1812 (N_1812,N_1610,N_1251);
nor U1813 (N_1813,N_1513,N_1661);
nand U1814 (N_1814,N_1366,N_1653);
nand U1815 (N_1815,N_1319,N_1788);
nor U1816 (N_1816,N_1350,N_1465);
nor U1817 (N_1817,N_1655,N_1553);
nand U1818 (N_1818,N_1204,N_1639);
and U1819 (N_1819,N_1763,N_1267);
or U1820 (N_1820,N_1432,N_1714);
or U1821 (N_1821,N_1501,N_1232);
and U1822 (N_1822,N_1467,N_1662);
nand U1823 (N_1823,N_1449,N_1202);
nor U1824 (N_1824,N_1301,N_1256);
nor U1825 (N_1825,N_1684,N_1735);
nand U1826 (N_1826,N_1534,N_1364);
and U1827 (N_1827,N_1390,N_1623);
and U1828 (N_1828,N_1704,N_1396);
nand U1829 (N_1829,N_1636,N_1664);
nor U1830 (N_1830,N_1602,N_1537);
nand U1831 (N_1831,N_1792,N_1367);
and U1832 (N_1832,N_1777,N_1739);
nand U1833 (N_1833,N_1291,N_1292);
and U1834 (N_1834,N_1403,N_1708);
or U1835 (N_1835,N_1242,N_1563);
and U1836 (N_1836,N_1369,N_1517);
or U1837 (N_1837,N_1566,N_1480);
nor U1838 (N_1838,N_1712,N_1286);
nand U1839 (N_1839,N_1436,N_1689);
nand U1840 (N_1840,N_1453,N_1450);
nand U1841 (N_1841,N_1762,N_1798);
and U1842 (N_1842,N_1452,N_1404);
and U1843 (N_1843,N_1786,N_1568);
and U1844 (N_1844,N_1254,N_1383);
nor U1845 (N_1845,N_1783,N_1360);
and U1846 (N_1846,N_1670,N_1295);
and U1847 (N_1847,N_1339,N_1514);
or U1848 (N_1848,N_1278,N_1665);
nand U1849 (N_1849,N_1525,N_1549);
or U1850 (N_1850,N_1299,N_1379);
or U1851 (N_1851,N_1541,N_1754);
nor U1852 (N_1852,N_1377,N_1418);
or U1853 (N_1853,N_1523,N_1635);
nor U1854 (N_1854,N_1229,N_1615);
or U1855 (N_1855,N_1311,N_1620);
nor U1856 (N_1856,N_1764,N_1674);
and U1857 (N_1857,N_1780,N_1410);
and U1858 (N_1858,N_1782,N_1614);
and U1859 (N_1859,N_1422,N_1234);
nand U1860 (N_1860,N_1499,N_1428);
nand U1861 (N_1861,N_1732,N_1381);
and U1862 (N_1862,N_1268,N_1645);
and U1863 (N_1863,N_1356,N_1679);
nor U1864 (N_1864,N_1622,N_1616);
and U1865 (N_1865,N_1641,N_1472);
and U1866 (N_1866,N_1203,N_1208);
nand U1867 (N_1867,N_1424,N_1279);
nor U1868 (N_1868,N_1680,N_1555);
nand U1869 (N_1869,N_1584,N_1742);
or U1870 (N_1870,N_1775,N_1470);
and U1871 (N_1871,N_1490,N_1439);
or U1872 (N_1872,N_1649,N_1334);
nand U1873 (N_1873,N_1337,N_1559);
nand U1874 (N_1874,N_1768,N_1711);
or U1875 (N_1875,N_1543,N_1216);
or U1876 (N_1876,N_1500,N_1416);
nor U1877 (N_1877,N_1625,N_1591);
nor U1878 (N_1878,N_1374,N_1382);
nor U1879 (N_1879,N_1743,N_1407);
and U1880 (N_1880,N_1315,N_1210);
and U1881 (N_1881,N_1321,N_1699);
and U1882 (N_1882,N_1435,N_1351);
or U1883 (N_1883,N_1494,N_1533);
xor U1884 (N_1884,N_1495,N_1668);
nand U1885 (N_1885,N_1751,N_1605);
and U1886 (N_1886,N_1389,N_1252);
or U1887 (N_1887,N_1522,N_1545);
nor U1888 (N_1888,N_1236,N_1427);
and U1889 (N_1889,N_1406,N_1235);
or U1890 (N_1890,N_1658,N_1222);
and U1891 (N_1891,N_1681,N_1542);
nor U1892 (N_1892,N_1642,N_1491);
and U1893 (N_1893,N_1617,N_1225);
and U1894 (N_1894,N_1758,N_1727);
nand U1895 (N_1895,N_1486,N_1437);
or U1896 (N_1896,N_1509,N_1333);
nand U1897 (N_1897,N_1506,N_1323);
nand U1898 (N_1898,N_1289,N_1710);
and U1899 (N_1899,N_1508,N_1765);
and U1900 (N_1900,N_1536,N_1206);
or U1901 (N_1901,N_1590,N_1211);
and U1902 (N_1902,N_1717,N_1487);
or U1903 (N_1903,N_1707,N_1497);
nand U1904 (N_1904,N_1217,N_1769);
or U1905 (N_1905,N_1705,N_1774);
and U1906 (N_1906,N_1475,N_1718);
or U1907 (N_1907,N_1535,N_1572);
or U1908 (N_1908,N_1220,N_1551);
nand U1909 (N_1909,N_1200,N_1269);
xnor U1910 (N_1910,N_1785,N_1488);
nand U1911 (N_1911,N_1247,N_1586);
or U1912 (N_1912,N_1729,N_1532);
nand U1913 (N_1913,N_1474,N_1651);
nor U1914 (N_1914,N_1611,N_1515);
or U1915 (N_1915,N_1271,N_1405);
or U1916 (N_1916,N_1752,N_1737);
or U1917 (N_1917,N_1414,N_1657);
nor U1918 (N_1918,N_1631,N_1720);
and U1919 (N_1919,N_1524,N_1736);
nand U1920 (N_1920,N_1565,N_1368);
nor U1921 (N_1921,N_1519,N_1596);
or U1922 (N_1922,N_1275,N_1233);
and U1923 (N_1923,N_1361,N_1546);
nand U1924 (N_1924,N_1626,N_1294);
and U1925 (N_1925,N_1527,N_1398);
and U1926 (N_1926,N_1692,N_1759);
nor U1927 (N_1927,N_1454,N_1322);
nor U1928 (N_1928,N_1671,N_1702);
nand U1929 (N_1929,N_1346,N_1634);
nor U1930 (N_1930,N_1358,N_1660);
or U1931 (N_1931,N_1592,N_1621);
nand U1932 (N_1932,N_1290,N_1362);
nand U1933 (N_1933,N_1391,N_1633);
and U1934 (N_1934,N_1325,N_1304);
nor U1935 (N_1935,N_1434,N_1579);
nor U1936 (N_1936,N_1518,N_1409);
or U1937 (N_1937,N_1261,N_1462);
nand U1938 (N_1938,N_1250,N_1726);
nor U1939 (N_1939,N_1274,N_1673);
or U1940 (N_1940,N_1746,N_1505);
nor U1941 (N_1941,N_1237,N_1309);
nor U1942 (N_1942,N_1260,N_1531);
or U1943 (N_1943,N_1357,N_1608);
nand U1944 (N_1944,N_1516,N_1770);
or U1945 (N_1945,N_1226,N_1701);
and U1946 (N_1946,N_1687,N_1569);
or U1947 (N_1947,N_1700,N_1393);
nand U1948 (N_1948,N_1588,N_1589);
nor U1949 (N_1949,N_1246,N_1547);
nor U1950 (N_1950,N_1779,N_1789);
and U1951 (N_1951,N_1760,N_1438);
nand U1952 (N_1952,N_1354,N_1576);
or U1953 (N_1953,N_1709,N_1277);
nor U1954 (N_1954,N_1288,N_1682);
nor U1955 (N_1955,N_1540,N_1666);
nor U1956 (N_1956,N_1593,N_1442);
and U1957 (N_1957,N_1329,N_1265);
nand U1958 (N_1958,N_1400,N_1643);
or U1959 (N_1959,N_1308,N_1628);
and U1960 (N_1960,N_1761,N_1570);
or U1961 (N_1961,N_1577,N_1772);
nand U1962 (N_1962,N_1793,N_1280);
and U1963 (N_1963,N_1561,N_1359);
nand U1964 (N_1964,N_1646,N_1599);
nor U1965 (N_1965,N_1338,N_1629);
nand U1966 (N_1966,N_1728,N_1207);
and U1967 (N_1967,N_1753,N_1460);
nand U1968 (N_1968,N_1266,N_1511);
nand U1969 (N_1969,N_1723,N_1459);
or U1970 (N_1970,N_1219,N_1734);
and U1971 (N_1971,N_1552,N_1744);
nor U1972 (N_1972,N_1458,N_1371);
and U1973 (N_1973,N_1581,N_1557);
and U1974 (N_1974,N_1594,N_1784);
nor U1975 (N_1975,N_1310,N_1669);
or U1976 (N_1976,N_1417,N_1672);
or U1977 (N_1977,N_1526,N_1392);
nand U1978 (N_1978,N_1270,N_1420);
and U1979 (N_1979,N_1489,N_1415);
and U1980 (N_1980,N_1571,N_1205);
or U1981 (N_1981,N_1675,N_1328);
and U1982 (N_1982,N_1724,N_1693);
nand U1983 (N_1983,N_1214,N_1688);
and U1984 (N_1984,N_1209,N_1259);
nor U1985 (N_1985,N_1476,N_1324);
nor U1986 (N_1986,N_1567,N_1482);
or U1987 (N_1987,N_1694,N_1335);
nor U1988 (N_1988,N_1388,N_1663);
or U1989 (N_1989,N_1493,N_1484);
nand U1990 (N_1990,N_1483,N_1326);
nand U1991 (N_1991,N_1451,N_1791);
and U1992 (N_1992,N_1318,N_1347);
nor U1993 (N_1993,N_1223,N_1691);
or U1994 (N_1994,N_1587,N_1554);
or U1995 (N_1995,N_1650,N_1573);
nor U1996 (N_1996,N_1678,N_1600);
nand U1997 (N_1997,N_1716,N_1425);
and U1998 (N_1998,N_1747,N_1239);
nand U1999 (N_1999,N_1738,N_1426);
or U2000 (N_2000,N_1469,N_1212);
nand U2001 (N_2001,N_1609,N_1457);
nor U2002 (N_2002,N_1394,N_1245);
or U2003 (N_2003,N_1598,N_1507);
nor U2004 (N_2004,N_1479,N_1273);
or U2005 (N_2005,N_1740,N_1296);
and U2006 (N_2006,N_1638,N_1698);
or U2007 (N_2007,N_1471,N_1637);
and U2008 (N_2008,N_1750,N_1307);
nand U2009 (N_2009,N_1316,N_1456);
nand U2010 (N_2010,N_1647,N_1272);
nand U2011 (N_2011,N_1276,N_1455);
nor U2012 (N_2012,N_1243,N_1336);
and U2013 (N_2013,N_1257,N_1604);
nor U2014 (N_2014,N_1380,N_1560);
or U2015 (N_2015,N_1607,N_1677);
or U2016 (N_2016,N_1477,N_1504);
nor U2017 (N_2017,N_1468,N_1375);
nand U2018 (N_2018,N_1648,N_1630);
nor U2019 (N_2019,N_1227,N_1498);
nor U2020 (N_2020,N_1613,N_1384);
nand U2021 (N_2021,N_1492,N_1757);
nand U2022 (N_2022,N_1787,N_1461);
nor U2023 (N_2023,N_1244,N_1287);
and U2024 (N_2024,N_1249,N_1281);
and U2025 (N_2025,N_1731,N_1745);
and U2026 (N_2026,N_1686,N_1433);
and U2027 (N_2027,N_1332,N_1703);
or U2028 (N_2028,N_1248,N_1305);
nor U2029 (N_2029,N_1285,N_1264);
or U2030 (N_2030,N_1370,N_1578);
or U2031 (N_2031,N_1640,N_1725);
or U2032 (N_2032,N_1564,N_1741);
nor U2033 (N_2033,N_1431,N_1376);
nand U2034 (N_2034,N_1463,N_1255);
and U2035 (N_2035,N_1466,N_1696);
nand U2036 (N_2036,N_1582,N_1715);
and U2037 (N_2037,N_1363,N_1503);
xor U2038 (N_2038,N_1685,N_1345);
nand U2039 (N_2039,N_1297,N_1317);
or U2040 (N_2040,N_1512,N_1221);
or U2041 (N_2041,N_1749,N_1550);
or U2042 (N_2042,N_1408,N_1654);
nor U2043 (N_2043,N_1413,N_1228);
nand U2044 (N_2044,N_1201,N_1539);
and U2045 (N_2045,N_1313,N_1302);
and U2046 (N_2046,N_1342,N_1481);
nand U2047 (N_2047,N_1218,N_1676);
nand U2048 (N_2048,N_1430,N_1721);
nor U2049 (N_2049,N_1722,N_1538);
or U2050 (N_2050,N_1314,N_1766);
or U2051 (N_2051,N_1473,N_1652);
and U2052 (N_2052,N_1343,N_1349);
nor U2053 (N_2053,N_1373,N_1767);
xnor U2054 (N_2054,N_1529,N_1253);
nand U2055 (N_2055,N_1478,N_1585);
and U2056 (N_2056,N_1619,N_1352);
or U2057 (N_2057,N_1293,N_1298);
and U2058 (N_2058,N_1224,N_1580);
nor U2059 (N_2059,N_1306,N_1773);
nand U2060 (N_2060,N_1776,N_1445);
or U2061 (N_2061,N_1282,N_1355);
nand U2062 (N_2062,N_1558,N_1231);
and U2063 (N_2063,N_1713,N_1440);
or U2064 (N_2064,N_1344,N_1790);
nor U2065 (N_2065,N_1719,N_1443);
xnor U2066 (N_2066,N_1378,N_1262);
xor U2067 (N_2067,N_1730,N_1331);
or U2068 (N_2068,N_1612,N_1411);
or U2069 (N_2069,N_1556,N_1624);
or U2070 (N_2070,N_1695,N_1429);
nor U2071 (N_2071,N_1530,N_1606);
nand U2072 (N_2072,N_1283,N_1485);
and U2073 (N_2073,N_1632,N_1601);
nand U2074 (N_2074,N_1365,N_1230);
or U2075 (N_2075,N_1402,N_1447);
or U2076 (N_2076,N_1387,N_1690);
nor U2077 (N_2077,N_1627,N_1240);
nor U2078 (N_2078,N_1755,N_1778);
or U2079 (N_2079,N_1353,N_1284);
and U2080 (N_2080,N_1320,N_1756);
nor U2081 (N_2081,N_1397,N_1330);
nand U2082 (N_2082,N_1795,N_1340);
nand U2083 (N_2083,N_1510,N_1667);
nor U2084 (N_2084,N_1327,N_1644);
nand U2085 (N_2085,N_1258,N_1419);
or U2086 (N_2086,N_1771,N_1520);
and U2087 (N_2087,N_1341,N_1575);
and U2088 (N_2088,N_1796,N_1781);
and U2089 (N_2089,N_1603,N_1401);
nand U2090 (N_2090,N_1597,N_1528);
or U2091 (N_2091,N_1502,N_1733);
nor U2092 (N_2092,N_1562,N_1399);
and U2093 (N_2093,N_1412,N_1683);
nand U2094 (N_2094,N_1215,N_1583);
nand U2095 (N_2095,N_1794,N_1263);
and U2096 (N_2096,N_1548,N_1659);
nor U2097 (N_2097,N_1441,N_1748);
nand U2098 (N_2098,N_1241,N_1574);
nand U2099 (N_2099,N_1496,N_1386);
nand U2100 (N_2100,N_1452,N_1346);
and U2101 (N_2101,N_1253,N_1434);
nand U2102 (N_2102,N_1768,N_1483);
nand U2103 (N_2103,N_1462,N_1513);
nor U2104 (N_2104,N_1299,N_1277);
and U2105 (N_2105,N_1466,N_1242);
nor U2106 (N_2106,N_1264,N_1788);
and U2107 (N_2107,N_1453,N_1216);
nor U2108 (N_2108,N_1642,N_1769);
or U2109 (N_2109,N_1415,N_1222);
or U2110 (N_2110,N_1393,N_1243);
nor U2111 (N_2111,N_1545,N_1354);
nand U2112 (N_2112,N_1574,N_1495);
or U2113 (N_2113,N_1543,N_1496);
and U2114 (N_2114,N_1403,N_1307);
or U2115 (N_2115,N_1773,N_1514);
or U2116 (N_2116,N_1762,N_1389);
or U2117 (N_2117,N_1577,N_1331);
or U2118 (N_2118,N_1641,N_1475);
nor U2119 (N_2119,N_1422,N_1640);
and U2120 (N_2120,N_1791,N_1553);
nor U2121 (N_2121,N_1525,N_1604);
nor U2122 (N_2122,N_1548,N_1751);
nor U2123 (N_2123,N_1253,N_1698);
nor U2124 (N_2124,N_1527,N_1730);
xnor U2125 (N_2125,N_1682,N_1320);
nor U2126 (N_2126,N_1313,N_1370);
or U2127 (N_2127,N_1545,N_1532);
and U2128 (N_2128,N_1467,N_1685);
and U2129 (N_2129,N_1664,N_1365);
or U2130 (N_2130,N_1672,N_1455);
and U2131 (N_2131,N_1628,N_1629);
nor U2132 (N_2132,N_1622,N_1466);
nor U2133 (N_2133,N_1326,N_1699);
nand U2134 (N_2134,N_1315,N_1213);
nand U2135 (N_2135,N_1724,N_1295);
nor U2136 (N_2136,N_1327,N_1575);
and U2137 (N_2137,N_1535,N_1740);
nor U2138 (N_2138,N_1645,N_1488);
and U2139 (N_2139,N_1758,N_1262);
or U2140 (N_2140,N_1712,N_1251);
nor U2141 (N_2141,N_1572,N_1621);
or U2142 (N_2142,N_1505,N_1382);
and U2143 (N_2143,N_1531,N_1673);
or U2144 (N_2144,N_1422,N_1618);
xor U2145 (N_2145,N_1711,N_1305);
or U2146 (N_2146,N_1707,N_1681);
nand U2147 (N_2147,N_1218,N_1436);
nor U2148 (N_2148,N_1573,N_1632);
and U2149 (N_2149,N_1460,N_1540);
nor U2150 (N_2150,N_1722,N_1570);
or U2151 (N_2151,N_1691,N_1313);
or U2152 (N_2152,N_1690,N_1393);
or U2153 (N_2153,N_1648,N_1308);
nand U2154 (N_2154,N_1324,N_1506);
or U2155 (N_2155,N_1710,N_1268);
or U2156 (N_2156,N_1494,N_1327);
or U2157 (N_2157,N_1799,N_1749);
and U2158 (N_2158,N_1435,N_1560);
and U2159 (N_2159,N_1252,N_1690);
and U2160 (N_2160,N_1787,N_1725);
nand U2161 (N_2161,N_1356,N_1489);
nand U2162 (N_2162,N_1564,N_1228);
nand U2163 (N_2163,N_1727,N_1652);
nand U2164 (N_2164,N_1482,N_1744);
nor U2165 (N_2165,N_1664,N_1783);
xor U2166 (N_2166,N_1452,N_1632);
and U2167 (N_2167,N_1546,N_1424);
or U2168 (N_2168,N_1699,N_1742);
nand U2169 (N_2169,N_1657,N_1717);
nand U2170 (N_2170,N_1203,N_1358);
and U2171 (N_2171,N_1229,N_1379);
nor U2172 (N_2172,N_1319,N_1657);
and U2173 (N_2173,N_1719,N_1489);
or U2174 (N_2174,N_1738,N_1658);
nor U2175 (N_2175,N_1432,N_1399);
or U2176 (N_2176,N_1319,N_1627);
nand U2177 (N_2177,N_1428,N_1286);
nor U2178 (N_2178,N_1213,N_1728);
and U2179 (N_2179,N_1563,N_1414);
nand U2180 (N_2180,N_1427,N_1391);
or U2181 (N_2181,N_1690,N_1665);
or U2182 (N_2182,N_1337,N_1771);
nor U2183 (N_2183,N_1525,N_1782);
nor U2184 (N_2184,N_1216,N_1425);
or U2185 (N_2185,N_1466,N_1516);
or U2186 (N_2186,N_1614,N_1201);
and U2187 (N_2187,N_1382,N_1510);
nor U2188 (N_2188,N_1367,N_1247);
nand U2189 (N_2189,N_1325,N_1415);
and U2190 (N_2190,N_1645,N_1568);
and U2191 (N_2191,N_1637,N_1486);
nand U2192 (N_2192,N_1232,N_1361);
and U2193 (N_2193,N_1654,N_1575);
nand U2194 (N_2194,N_1669,N_1258);
or U2195 (N_2195,N_1452,N_1716);
nand U2196 (N_2196,N_1250,N_1424);
nor U2197 (N_2197,N_1592,N_1649);
nand U2198 (N_2198,N_1444,N_1622);
nor U2199 (N_2199,N_1760,N_1414);
nand U2200 (N_2200,N_1377,N_1791);
or U2201 (N_2201,N_1625,N_1561);
and U2202 (N_2202,N_1284,N_1739);
nand U2203 (N_2203,N_1736,N_1635);
nand U2204 (N_2204,N_1503,N_1530);
nor U2205 (N_2205,N_1252,N_1473);
nand U2206 (N_2206,N_1482,N_1339);
and U2207 (N_2207,N_1226,N_1224);
or U2208 (N_2208,N_1692,N_1350);
nor U2209 (N_2209,N_1304,N_1758);
nand U2210 (N_2210,N_1416,N_1545);
and U2211 (N_2211,N_1340,N_1579);
or U2212 (N_2212,N_1636,N_1793);
and U2213 (N_2213,N_1328,N_1529);
nand U2214 (N_2214,N_1332,N_1654);
nand U2215 (N_2215,N_1701,N_1678);
and U2216 (N_2216,N_1470,N_1268);
or U2217 (N_2217,N_1260,N_1701);
nand U2218 (N_2218,N_1287,N_1424);
nand U2219 (N_2219,N_1594,N_1418);
and U2220 (N_2220,N_1343,N_1316);
and U2221 (N_2221,N_1619,N_1473);
nor U2222 (N_2222,N_1559,N_1571);
and U2223 (N_2223,N_1303,N_1521);
nand U2224 (N_2224,N_1534,N_1450);
nand U2225 (N_2225,N_1377,N_1784);
nor U2226 (N_2226,N_1655,N_1639);
or U2227 (N_2227,N_1670,N_1488);
nand U2228 (N_2228,N_1731,N_1554);
nor U2229 (N_2229,N_1490,N_1442);
nand U2230 (N_2230,N_1749,N_1714);
or U2231 (N_2231,N_1226,N_1361);
and U2232 (N_2232,N_1773,N_1333);
and U2233 (N_2233,N_1386,N_1489);
nand U2234 (N_2234,N_1687,N_1425);
nor U2235 (N_2235,N_1364,N_1231);
nand U2236 (N_2236,N_1768,N_1769);
and U2237 (N_2237,N_1766,N_1487);
and U2238 (N_2238,N_1225,N_1342);
nor U2239 (N_2239,N_1456,N_1638);
and U2240 (N_2240,N_1445,N_1293);
nand U2241 (N_2241,N_1726,N_1436);
nand U2242 (N_2242,N_1299,N_1348);
or U2243 (N_2243,N_1313,N_1637);
and U2244 (N_2244,N_1289,N_1429);
and U2245 (N_2245,N_1299,N_1709);
nand U2246 (N_2246,N_1584,N_1461);
nand U2247 (N_2247,N_1605,N_1438);
nor U2248 (N_2248,N_1268,N_1225);
nor U2249 (N_2249,N_1298,N_1315);
or U2250 (N_2250,N_1668,N_1731);
nand U2251 (N_2251,N_1605,N_1645);
and U2252 (N_2252,N_1258,N_1783);
nor U2253 (N_2253,N_1386,N_1722);
xnor U2254 (N_2254,N_1705,N_1263);
nor U2255 (N_2255,N_1331,N_1490);
and U2256 (N_2256,N_1584,N_1266);
nand U2257 (N_2257,N_1711,N_1526);
or U2258 (N_2258,N_1663,N_1632);
nor U2259 (N_2259,N_1365,N_1707);
nor U2260 (N_2260,N_1238,N_1763);
and U2261 (N_2261,N_1578,N_1366);
and U2262 (N_2262,N_1390,N_1309);
and U2263 (N_2263,N_1682,N_1794);
nor U2264 (N_2264,N_1240,N_1726);
and U2265 (N_2265,N_1691,N_1426);
and U2266 (N_2266,N_1509,N_1770);
nand U2267 (N_2267,N_1297,N_1637);
or U2268 (N_2268,N_1791,N_1349);
or U2269 (N_2269,N_1766,N_1264);
or U2270 (N_2270,N_1756,N_1364);
nand U2271 (N_2271,N_1696,N_1431);
nand U2272 (N_2272,N_1580,N_1759);
and U2273 (N_2273,N_1756,N_1681);
xor U2274 (N_2274,N_1501,N_1248);
nand U2275 (N_2275,N_1583,N_1603);
and U2276 (N_2276,N_1787,N_1754);
nor U2277 (N_2277,N_1549,N_1709);
and U2278 (N_2278,N_1776,N_1334);
and U2279 (N_2279,N_1399,N_1571);
or U2280 (N_2280,N_1675,N_1355);
and U2281 (N_2281,N_1618,N_1372);
nand U2282 (N_2282,N_1662,N_1210);
and U2283 (N_2283,N_1229,N_1653);
and U2284 (N_2284,N_1264,N_1270);
nand U2285 (N_2285,N_1320,N_1387);
nand U2286 (N_2286,N_1204,N_1368);
or U2287 (N_2287,N_1363,N_1704);
and U2288 (N_2288,N_1279,N_1352);
and U2289 (N_2289,N_1215,N_1728);
or U2290 (N_2290,N_1318,N_1712);
or U2291 (N_2291,N_1487,N_1604);
and U2292 (N_2292,N_1742,N_1319);
or U2293 (N_2293,N_1653,N_1455);
nor U2294 (N_2294,N_1486,N_1549);
nor U2295 (N_2295,N_1633,N_1275);
or U2296 (N_2296,N_1527,N_1450);
nor U2297 (N_2297,N_1274,N_1646);
nor U2298 (N_2298,N_1337,N_1429);
nand U2299 (N_2299,N_1442,N_1536);
and U2300 (N_2300,N_1446,N_1650);
nor U2301 (N_2301,N_1567,N_1782);
nor U2302 (N_2302,N_1796,N_1707);
nand U2303 (N_2303,N_1730,N_1647);
and U2304 (N_2304,N_1680,N_1571);
and U2305 (N_2305,N_1469,N_1363);
or U2306 (N_2306,N_1513,N_1694);
and U2307 (N_2307,N_1511,N_1653);
nor U2308 (N_2308,N_1767,N_1238);
nor U2309 (N_2309,N_1243,N_1200);
and U2310 (N_2310,N_1293,N_1501);
and U2311 (N_2311,N_1439,N_1280);
nand U2312 (N_2312,N_1698,N_1286);
nand U2313 (N_2313,N_1400,N_1595);
and U2314 (N_2314,N_1708,N_1367);
and U2315 (N_2315,N_1337,N_1514);
nand U2316 (N_2316,N_1690,N_1786);
nand U2317 (N_2317,N_1599,N_1285);
nand U2318 (N_2318,N_1603,N_1472);
or U2319 (N_2319,N_1296,N_1703);
or U2320 (N_2320,N_1267,N_1568);
and U2321 (N_2321,N_1403,N_1417);
and U2322 (N_2322,N_1485,N_1740);
nand U2323 (N_2323,N_1443,N_1448);
xnor U2324 (N_2324,N_1698,N_1470);
and U2325 (N_2325,N_1345,N_1330);
or U2326 (N_2326,N_1465,N_1421);
nor U2327 (N_2327,N_1311,N_1369);
or U2328 (N_2328,N_1435,N_1758);
or U2329 (N_2329,N_1402,N_1733);
and U2330 (N_2330,N_1287,N_1735);
and U2331 (N_2331,N_1645,N_1211);
nand U2332 (N_2332,N_1588,N_1636);
nor U2333 (N_2333,N_1650,N_1243);
nand U2334 (N_2334,N_1342,N_1430);
and U2335 (N_2335,N_1431,N_1526);
or U2336 (N_2336,N_1752,N_1310);
or U2337 (N_2337,N_1222,N_1734);
nor U2338 (N_2338,N_1657,N_1392);
and U2339 (N_2339,N_1323,N_1790);
nand U2340 (N_2340,N_1315,N_1478);
or U2341 (N_2341,N_1635,N_1374);
or U2342 (N_2342,N_1311,N_1256);
and U2343 (N_2343,N_1233,N_1472);
and U2344 (N_2344,N_1262,N_1258);
or U2345 (N_2345,N_1530,N_1511);
nand U2346 (N_2346,N_1614,N_1549);
and U2347 (N_2347,N_1310,N_1352);
and U2348 (N_2348,N_1399,N_1729);
nand U2349 (N_2349,N_1686,N_1202);
and U2350 (N_2350,N_1254,N_1774);
and U2351 (N_2351,N_1665,N_1216);
and U2352 (N_2352,N_1218,N_1319);
nand U2353 (N_2353,N_1517,N_1377);
and U2354 (N_2354,N_1776,N_1404);
or U2355 (N_2355,N_1514,N_1481);
nor U2356 (N_2356,N_1723,N_1508);
and U2357 (N_2357,N_1449,N_1514);
nor U2358 (N_2358,N_1738,N_1708);
nor U2359 (N_2359,N_1737,N_1544);
nor U2360 (N_2360,N_1230,N_1447);
and U2361 (N_2361,N_1297,N_1599);
and U2362 (N_2362,N_1606,N_1316);
nand U2363 (N_2363,N_1465,N_1219);
or U2364 (N_2364,N_1486,N_1571);
nor U2365 (N_2365,N_1220,N_1571);
and U2366 (N_2366,N_1751,N_1537);
nand U2367 (N_2367,N_1266,N_1252);
or U2368 (N_2368,N_1535,N_1451);
nor U2369 (N_2369,N_1500,N_1257);
and U2370 (N_2370,N_1240,N_1686);
nor U2371 (N_2371,N_1732,N_1517);
and U2372 (N_2372,N_1677,N_1618);
nand U2373 (N_2373,N_1532,N_1354);
nor U2374 (N_2374,N_1350,N_1708);
nand U2375 (N_2375,N_1401,N_1411);
nand U2376 (N_2376,N_1675,N_1751);
nand U2377 (N_2377,N_1464,N_1292);
and U2378 (N_2378,N_1578,N_1698);
and U2379 (N_2379,N_1725,N_1408);
and U2380 (N_2380,N_1787,N_1767);
or U2381 (N_2381,N_1615,N_1410);
and U2382 (N_2382,N_1527,N_1633);
and U2383 (N_2383,N_1522,N_1294);
or U2384 (N_2384,N_1423,N_1242);
or U2385 (N_2385,N_1304,N_1550);
or U2386 (N_2386,N_1754,N_1422);
and U2387 (N_2387,N_1592,N_1435);
and U2388 (N_2388,N_1682,N_1498);
or U2389 (N_2389,N_1394,N_1296);
nand U2390 (N_2390,N_1302,N_1369);
nor U2391 (N_2391,N_1308,N_1799);
and U2392 (N_2392,N_1400,N_1619);
and U2393 (N_2393,N_1597,N_1499);
nand U2394 (N_2394,N_1790,N_1727);
or U2395 (N_2395,N_1416,N_1426);
nand U2396 (N_2396,N_1311,N_1755);
or U2397 (N_2397,N_1247,N_1429);
or U2398 (N_2398,N_1701,N_1559);
nor U2399 (N_2399,N_1606,N_1772);
and U2400 (N_2400,N_2084,N_2335);
nor U2401 (N_2401,N_2353,N_2271);
or U2402 (N_2402,N_2075,N_1970);
nor U2403 (N_2403,N_2056,N_2113);
nand U2404 (N_2404,N_2085,N_2312);
and U2405 (N_2405,N_1863,N_2374);
nor U2406 (N_2406,N_2384,N_1969);
nor U2407 (N_2407,N_2072,N_2106);
and U2408 (N_2408,N_1848,N_2235);
nand U2409 (N_2409,N_2135,N_2361);
or U2410 (N_2410,N_1880,N_2129);
nor U2411 (N_2411,N_1869,N_1883);
or U2412 (N_2412,N_2303,N_2371);
and U2413 (N_2413,N_2150,N_2051);
or U2414 (N_2414,N_2182,N_2111);
nor U2415 (N_2415,N_1908,N_1836);
nand U2416 (N_2416,N_2260,N_2004);
and U2417 (N_2417,N_2318,N_2214);
or U2418 (N_2418,N_2146,N_1844);
nand U2419 (N_2419,N_2267,N_2003);
and U2420 (N_2420,N_2366,N_2045);
nand U2421 (N_2421,N_1859,N_2245);
or U2422 (N_2422,N_2376,N_1973);
or U2423 (N_2423,N_1841,N_1989);
and U2424 (N_2424,N_2096,N_2383);
nand U2425 (N_2425,N_2041,N_2259);
nand U2426 (N_2426,N_2270,N_2205);
nor U2427 (N_2427,N_2298,N_1920);
and U2428 (N_2428,N_1937,N_2121);
nor U2429 (N_2429,N_2310,N_1926);
nor U2430 (N_2430,N_2037,N_2350);
and U2431 (N_2431,N_2141,N_2388);
and U2432 (N_2432,N_2014,N_2108);
nand U2433 (N_2433,N_2345,N_1906);
or U2434 (N_2434,N_2151,N_2273);
or U2435 (N_2435,N_2367,N_2039);
or U2436 (N_2436,N_2391,N_2282);
and U2437 (N_2437,N_2149,N_1837);
or U2438 (N_2438,N_2170,N_2394);
nand U2439 (N_2439,N_2128,N_1825);
or U2440 (N_2440,N_1853,N_2065);
and U2441 (N_2441,N_2015,N_2148);
nor U2442 (N_2442,N_1835,N_2239);
nand U2443 (N_2443,N_2049,N_2192);
or U2444 (N_2444,N_2197,N_2082);
nand U2445 (N_2445,N_2287,N_1830);
nand U2446 (N_2446,N_1999,N_2316);
or U2447 (N_2447,N_2342,N_2329);
and U2448 (N_2448,N_1854,N_2105);
nand U2449 (N_2449,N_2138,N_1925);
and U2450 (N_2450,N_2324,N_1953);
nand U2451 (N_2451,N_2132,N_2022);
nor U2452 (N_2452,N_1885,N_1914);
nor U2453 (N_2453,N_2363,N_2044);
nor U2454 (N_2454,N_2089,N_2248);
nand U2455 (N_2455,N_1949,N_2175);
nor U2456 (N_2456,N_2078,N_2364);
nor U2457 (N_2457,N_1899,N_2166);
nor U2458 (N_2458,N_2274,N_1918);
and U2459 (N_2459,N_1988,N_2092);
nand U2460 (N_2460,N_2055,N_1803);
nor U2461 (N_2461,N_2086,N_1986);
and U2462 (N_2462,N_2352,N_2358);
or U2463 (N_2463,N_2008,N_2220);
and U2464 (N_2464,N_2378,N_1807);
nor U2465 (N_2465,N_2326,N_2024);
nor U2466 (N_2466,N_1958,N_2377);
nor U2467 (N_2467,N_2144,N_1978);
nor U2468 (N_2468,N_1829,N_2227);
nor U2469 (N_2469,N_2261,N_1931);
nand U2470 (N_2470,N_1947,N_1942);
or U2471 (N_2471,N_2201,N_2278);
and U2472 (N_2472,N_1802,N_2140);
nor U2473 (N_2473,N_2397,N_2334);
nand U2474 (N_2474,N_2372,N_2018);
and U2475 (N_2475,N_2059,N_2308);
nor U2476 (N_2476,N_1913,N_1984);
and U2477 (N_2477,N_2076,N_2338);
nand U2478 (N_2478,N_2188,N_2153);
nor U2479 (N_2479,N_2299,N_2203);
or U2480 (N_2480,N_2221,N_1983);
and U2481 (N_2481,N_1816,N_1946);
or U2482 (N_2482,N_2002,N_2233);
nand U2483 (N_2483,N_2266,N_1977);
nand U2484 (N_2484,N_2207,N_1855);
or U2485 (N_2485,N_2293,N_2213);
nand U2486 (N_2486,N_2053,N_2143);
and U2487 (N_2487,N_2191,N_2000);
or U2488 (N_2488,N_1887,N_1974);
or U2489 (N_2489,N_1871,N_1804);
nor U2490 (N_2490,N_2011,N_1826);
or U2491 (N_2491,N_1993,N_1957);
nor U2492 (N_2492,N_1858,N_2058);
nor U2493 (N_2493,N_2385,N_2167);
and U2494 (N_2494,N_1895,N_1875);
nand U2495 (N_2495,N_1805,N_2124);
nor U2496 (N_2496,N_2046,N_2171);
and U2497 (N_2497,N_2160,N_1818);
and U2498 (N_2498,N_2328,N_2262);
nand U2499 (N_2499,N_2231,N_2225);
nand U2500 (N_2500,N_1929,N_2375);
nand U2501 (N_2501,N_1877,N_2208);
or U2502 (N_2502,N_1847,N_1801);
and U2503 (N_2503,N_2200,N_2063);
or U2504 (N_2504,N_1922,N_1980);
nor U2505 (N_2505,N_2288,N_1945);
or U2506 (N_2506,N_2064,N_2365);
nand U2507 (N_2507,N_2336,N_2032);
and U2508 (N_2508,N_2280,N_1924);
and U2509 (N_2509,N_2038,N_2252);
or U2510 (N_2510,N_2211,N_2222);
and U2511 (N_2511,N_1898,N_2346);
and U2512 (N_2512,N_2165,N_1897);
or U2513 (N_2513,N_2322,N_1891);
or U2514 (N_2514,N_1971,N_1867);
or U2515 (N_2515,N_1907,N_2209);
nor U2516 (N_2516,N_2136,N_2370);
or U2517 (N_2517,N_1972,N_2180);
nand U2518 (N_2518,N_2110,N_2242);
nand U2519 (N_2519,N_2118,N_2265);
or U2520 (N_2520,N_2253,N_1903);
nand U2521 (N_2521,N_2283,N_1811);
nand U2522 (N_2522,N_2284,N_1991);
nand U2523 (N_2523,N_2119,N_2176);
and U2524 (N_2524,N_2177,N_1919);
nand U2525 (N_2525,N_2134,N_2381);
nand U2526 (N_2526,N_2195,N_2054);
or U2527 (N_2527,N_1956,N_1881);
nand U2528 (N_2528,N_1938,N_2306);
and U2529 (N_2529,N_2154,N_2027);
or U2530 (N_2530,N_2157,N_1806);
nand U2531 (N_2531,N_2190,N_2216);
nand U2532 (N_2532,N_1936,N_1981);
nor U2533 (N_2533,N_1954,N_2099);
or U2534 (N_2534,N_2295,N_2393);
and U2535 (N_2535,N_2343,N_2204);
and U2536 (N_2536,N_1962,N_2043);
or U2537 (N_2537,N_1966,N_2247);
nor U2538 (N_2538,N_2382,N_1889);
and U2539 (N_2539,N_2301,N_2183);
and U2540 (N_2540,N_2268,N_2198);
or U2541 (N_2541,N_2010,N_1948);
nand U2542 (N_2542,N_1862,N_2093);
nand U2543 (N_2543,N_2351,N_1992);
nor U2544 (N_2544,N_2215,N_2300);
and U2545 (N_2545,N_1896,N_2071);
or U2546 (N_2546,N_2229,N_1968);
or U2547 (N_2547,N_2088,N_2289);
nand U2548 (N_2548,N_2291,N_1856);
nand U2549 (N_2549,N_2158,N_2147);
or U2550 (N_2550,N_2142,N_2103);
and U2551 (N_2551,N_2159,N_1876);
nor U2552 (N_2552,N_1813,N_2276);
or U2553 (N_2553,N_1838,N_1912);
and U2554 (N_2554,N_2028,N_2073);
nor U2555 (N_2555,N_2025,N_2285);
or U2556 (N_2556,N_1870,N_2035);
xor U2557 (N_2557,N_1932,N_1845);
nor U2558 (N_2558,N_2033,N_2369);
and U2559 (N_2559,N_2001,N_2311);
or U2560 (N_2560,N_1990,N_2390);
nor U2561 (N_2561,N_1901,N_2052);
nor U2562 (N_2562,N_2019,N_2320);
nor U2563 (N_2563,N_1843,N_1902);
nand U2564 (N_2564,N_2309,N_1996);
nor U2565 (N_2565,N_2185,N_2199);
nand U2566 (N_2566,N_1861,N_1995);
and U2567 (N_2567,N_2281,N_1900);
nand U2568 (N_2568,N_2137,N_2187);
nor U2569 (N_2569,N_1888,N_1943);
and U2570 (N_2570,N_2067,N_2258);
nor U2571 (N_2571,N_2169,N_2243);
and U2572 (N_2572,N_1909,N_1874);
and U2573 (N_2573,N_2272,N_2087);
nand U2574 (N_2574,N_2079,N_2083);
or U2575 (N_2575,N_2050,N_2164);
or U2576 (N_2576,N_2319,N_1911);
or U2577 (N_2577,N_2219,N_1828);
nor U2578 (N_2578,N_2396,N_1927);
or U2579 (N_2579,N_1873,N_1872);
and U2580 (N_2580,N_2029,N_2189);
and U2581 (N_2581,N_1808,N_2355);
nand U2582 (N_2582,N_2179,N_2020);
nand U2583 (N_2583,N_2057,N_2254);
and U2584 (N_2584,N_2330,N_1821);
and U2585 (N_2585,N_2347,N_2237);
nor U2586 (N_2586,N_2292,N_1851);
or U2587 (N_2587,N_2206,N_2104);
or U2588 (N_2588,N_2304,N_1951);
and U2589 (N_2589,N_1985,N_1941);
or U2590 (N_2590,N_2095,N_2249);
nor U2591 (N_2591,N_2339,N_2307);
or U2592 (N_2592,N_1979,N_1967);
or U2593 (N_2593,N_2202,N_2122);
nand U2594 (N_2594,N_2362,N_2314);
nor U2595 (N_2595,N_2256,N_2332);
nor U2596 (N_2596,N_2244,N_2115);
or U2597 (N_2597,N_1930,N_1917);
nor U2598 (N_2598,N_2062,N_2098);
or U2599 (N_2599,N_2255,N_2163);
and U2600 (N_2600,N_1950,N_2047);
nor U2601 (N_2601,N_1886,N_2226);
and U2602 (N_2602,N_1849,N_1923);
and U2603 (N_2603,N_1976,N_1833);
or U2604 (N_2604,N_2349,N_1940);
or U2605 (N_2605,N_2090,N_2246);
nand U2606 (N_2606,N_2109,N_2181);
nor U2607 (N_2607,N_2107,N_1893);
nand U2608 (N_2608,N_1834,N_2210);
nand U2609 (N_2609,N_2005,N_2184);
or U2610 (N_2610,N_2036,N_1832);
nor U2611 (N_2611,N_1846,N_1960);
and U2612 (N_2612,N_1842,N_1878);
or U2613 (N_2613,N_2392,N_2102);
nor U2614 (N_2614,N_2114,N_2130);
nand U2615 (N_2615,N_2241,N_2077);
nand U2616 (N_2616,N_2100,N_1975);
and U2617 (N_2617,N_2359,N_2126);
or U2618 (N_2618,N_1819,N_2123);
and U2619 (N_2619,N_2368,N_2277);
nor U2620 (N_2620,N_2315,N_1904);
nor U2621 (N_2621,N_2162,N_1916);
and U2622 (N_2622,N_2238,N_2145);
nor U2623 (N_2623,N_2091,N_2275);
and U2624 (N_2624,N_2264,N_2186);
nor U2625 (N_2625,N_2380,N_1852);
nand U2626 (N_2626,N_2070,N_2156);
or U2627 (N_2627,N_2340,N_1952);
nand U2628 (N_2628,N_2399,N_2069);
nand U2629 (N_2629,N_1961,N_2006);
nor U2630 (N_2630,N_2168,N_1910);
nand U2631 (N_2631,N_1884,N_2257);
and U2632 (N_2632,N_1860,N_2373);
nand U2633 (N_2633,N_2196,N_1892);
and U2634 (N_2634,N_1894,N_2223);
or U2635 (N_2635,N_2269,N_2060);
nor U2636 (N_2636,N_2357,N_1823);
nand U2637 (N_2637,N_2080,N_2236);
nand U2638 (N_2638,N_2012,N_2302);
nor U2639 (N_2639,N_2026,N_2290);
and U2640 (N_2640,N_2341,N_2354);
or U2641 (N_2641,N_2356,N_2133);
nand U2642 (N_2642,N_1879,N_2230);
nand U2643 (N_2643,N_1865,N_2331);
and U2644 (N_2644,N_2021,N_1965);
and U2645 (N_2645,N_1994,N_2321);
or U2646 (N_2646,N_1982,N_1822);
nor U2647 (N_2647,N_2017,N_1840);
or U2648 (N_2648,N_2074,N_2240);
or U2649 (N_2649,N_2296,N_1815);
nor U2650 (N_2650,N_1882,N_2161);
or U2651 (N_2651,N_2117,N_1814);
nor U2652 (N_2652,N_2323,N_2066);
or U2653 (N_2653,N_2386,N_2034);
and U2654 (N_2654,N_1928,N_1817);
and U2655 (N_2655,N_1831,N_1866);
nor U2656 (N_2656,N_1850,N_1935);
or U2657 (N_2657,N_2048,N_2007);
nand U2658 (N_2658,N_2305,N_2313);
or U2659 (N_2659,N_2379,N_2031);
and U2660 (N_2660,N_2061,N_2218);
and U2661 (N_2661,N_2232,N_1905);
and U2662 (N_2662,N_2294,N_2337);
and U2663 (N_2663,N_1890,N_1939);
nor U2664 (N_2664,N_1987,N_1820);
nand U2665 (N_2665,N_2172,N_2116);
and U2666 (N_2666,N_1959,N_2217);
and U2667 (N_2667,N_2398,N_2228);
and U2668 (N_2668,N_2234,N_2327);
nand U2669 (N_2669,N_2224,N_1827);
or U2670 (N_2670,N_2317,N_2094);
or U2671 (N_2671,N_2125,N_1800);
nand U2672 (N_2672,N_2040,N_1944);
nor U2673 (N_2673,N_2030,N_2286);
and U2674 (N_2674,N_2131,N_1921);
or U2675 (N_2675,N_1934,N_1868);
nor U2676 (N_2676,N_2178,N_2120);
or U2677 (N_2677,N_1809,N_2279);
or U2678 (N_2678,N_2251,N_2081);
nor U2679 (N_2679,N_1857,N_2297);
or U2680 (N_2680,N_2139,N_2155);
nor U2681 (N_2681,N_2023,N_2193);
nand U2682 (N_2682,N_2127,N_1915);
nor U2683 (N_2683,N_1964,N_2068);
and U2684 (N_2684,N_2112,N_1824);
or U2685 (N_2685,N_2348,N_2042);
or U2686 (N_2686,N_2389,N_2333);
nor U2687 (N_2687,N_2387,N_2360);
and U2688 (N_2688,N_2013,N_2174);
and U2689 (N_2689,N_2250,N_2325);
or U2690 (N_2690,N_2395,N_2173);
nor U2691 (N_2691,N_2009,N_2212);
and U2692 (N_2692,N_1998,N_1963);
or U2693 (N_2693,N_1955,N_2263);
nor U2694 (N_2694,N_1810,N_1997);
and U2695 (N_2695,N_2016,N_2152);
and U2696 (N_2696,N_2194,N_2344);
nand U2697 (N_2697,N_2097,N_1933);
and U2698 (N_2698,N_1839,N_1812);
nand U2699 (N_2699,N_2101,N_1864);
nand U2700 (N_2700,N_1930,N_2382);
and U2701 (N_2701,N_2010,N_1884);
nor U2702 (N_2702,N_2196,N_2193);
or U2703 (N_2703,N_1827,N_2295);
nor U2704 (N_2704,N_1982,N_1926);
nand U2705 (N_2705,N_1986,N_1850);
or U2706 (N_2706,N_2361,N_1827);
or U2707 (N_2707,N_1959,N_2184);
or U2708 (N_2708,N_2257,N_2256);
and U2709 (N_2709,N_2040,N_2295);
nor U2710 (N_2710,N_1843,N_2309);
nand U2711 (N_2711,N_1836,N_1942);
or U2712 (N_2712,N_2377,N_2179);
and U2713 (N_2713,N_2108,N_2306);
xor U2714 (N_2714,N_1807,N_1846);
and U2715 (N_2715,N_2296,N_2062);
or U2716 (N_2716,N_2360,N_2219);
nand U2717 (N_2717,N_2217,N_2084);
nor U2718 (N_2718,N_2368,N_2372);
or U2719 (N_2719,N_1977,N_2146);
and U2720 (N_2720,N_2085,N_1908);
or U2721 (N_2721,N_1920,N_2054);
or U2722 (N_2722,N_2361,N_2391);
and U2723 (N_2723,N_1857,N_2111);
nor U2724 (N_2724,N_1806,N_2136);
nor U2725 (N_2725,N_1828,N_2230);
nand U2726 (N_2726,N_2016,N_2025);
nand U2727 (N_2727,N_1938,N_2234);
and U2728 (N_2728,N_1896,N_2325);
and U2729 (N_2729,N_2379,N_1973);
or U2730 (N_2730,N_2121,N_2298);
or U2731 (N_2731,N_1852,N_2344);
or U2732 (N_2732,N_2228,N_2264);
nor U2733 (N_2733,N_1809,N_1948);
and U2734 (N_2734,N_1988,N_1999);
and U2735 (N_2735,N_2030,N_2332);
or U2736 (N_2736,N_1864,N_2201);
xor U2737 (N_2737,N_2355,N_2224);
and U2738 (N_2738,N_2064,N_1849);
nand U2739 (N_2739,N_2181,N_1948);
nor U2740 (N_2740,N_1845,N_1902);
or U2741 (N_2741,N_2035,N_1854);
nand U2742 (N_2742,N_2056,N_1992);
nor U2743 (N_2743,N_2102,N_2161);
nor U2744 (N_2744,N_2131,N_2249);
or U2745 (N_2745,N_2144,N_1997);
and U2746 (N_2746,N_2204,N_2197);
nor U2747 (N_2747,N_2158,N_1919);
nor U2748 (N_2748,N_2371,N_2171);
nor U2749 (N_2749,N_1892,N_2168);
nor U2750 (N_2750,N_2330,N_2303);
nand U2751 (N_2751,N_2151,N_2030);
or U2752 (N_2752,N_2119,N_2353);
and U2753 (N_2753,N_1910,N_1871);
or U2754 (N_2754,N_2237,N_1827);
nand U2755 (N_2755,N_1928,N_1956);
or U2756 (N_2756,N_2220,N_1843);
nand U2757 (N_2757,N_1802,N_2135);
and U2758 (N_2758,N_2252,N_2395);
nand U2759 (N_2759,N_2151,N_1928);
or U2760 (N_2760,N_1867,N_2284);
nor U2761 (N_2761,N_2250,N_2202);
or U2762 (N_2762,N_1903,N_1840);
or U2763 (N_2763,N_2051,N_2040);
and U2764 (N_2764,N_1993,N_1964);
nand U2765 (N_2765,N_2121,N_2044);
nand U2766 (N_2766,N_1823,N_2136);
nand U2767 (N_2767,N_2239,N_1891);
and U2768 (N_2768,N_1958,N_2076);
or U2769 (N_2769,N_2368,N_2041);
or U2770 (N_2770,N_2109,N_1971);
nor U2771 (N_2771,N_2071,N_1800);
nor U2772 (N_2772,N_2272,N_2120);
or U2773 (N_2773,N_2161,N_2068);
and U2774 (N_2774,N_2056,N_1905);
nor U2775 (N_2775,N_2203,N_2266);
nand U2776 (N_2776,N_2240,N_1881);
nand U2777 (N_2777,N_1874,N_2163);
and U2778 (N_2778,N_1903,N_1895);
nand U2779 (N_2779,N_2138,N_1982);
nor U2780 (N_2780,N_2244,N_1823);
and U2781 (N_2781,N_2303,N_2070);
or U2782 (N_2782,N_1984,N_2211);
and U2783 (N_2783,N_2339,N_2230);
and U2784 (N_2784,N_2294,N_2147);
or U2785 (N_2785,N_1899,N_2314);
and U2786 (N_2786,N_1829,N_1987);
nor U2787 (N_2787,N_2027,N_2100);
nand U2788 (N_2788,N_1977,N_1826);
nor U2789 (N_2789,N_2292,N_2128);
or U2790 (N_2790,N_1848,N_2388);
nand U2791 (N_2791,N_1896,N_2371);
and U2792 (N_2792,N_1982,N_2379);
or U2793 (N_2793,N_1800,N_1899);
and U2794 (N_2794,N_1952,N_2287);
or U2795 (N_2795,N_1973,N_2314);
nand U2796 (N_2796,N_1800,N_2180);
nor U2797 (N_2797,N_2048,N_2171);
nand U2798 (N_2798,N_1906,N_2155);
and U2799 (N_2799,N_1881,N_2023);
nor U2800 (N_2800,N_2166,N_2032);
and U2801 (N_2801,N_2344,N_1990);
and U2802 (N_2802,N_2097,N_2176);
or U2803 (N_2803,N_2382,N_1979);
nand U2804 (N_2804,N_2048,N_1926);
nor U2805 (N_2805,N_2259,N_2018);
and U2806 (N_2806,N_2110,N_2090);
and U2807 (N_2807,N_2049,N_1976);
and U2808 (N_2808,N_2214,N_1978);
nand U2809 (N_2809,N_2285,N_1856);
and U2810 (N_2810,N_2307,N_1988);
and U2811 (N_2811,N_2054,N_1918);
nand U2812 (N_2812,N_2273,N_1944);
nand U2813 (N_2813,N_2159,N_2098);
or U2814 (N_2814,N_2315,N_2243);
xnor U2815 (N_2815,N_1937,N_1849);
or U2816 (N_2816,N_2190,N_1993);
and U2817 (N_2817,N_1955,N_2313);
and U2818 (N_2818,N_2224,N_2218);
and U2819 (N_2819,N_2334,N_2289);
nor U2820 (N_2820,N_2065,N_2387);
nor U2821 (N_2821,N_2014,N_2186);
nand U2822 (N_2822,N_2199,N_2348);
nand U2823 (N_2823,N_2207,N_1898);
and U2824 (N_2824,N_2220,N_2044);
nand U2825 (N_2825,N_2218,N_2323);
nor U2826 (N_2826,N_1987,N_2085);
or U2827 (N_2827,N_2249,N_2219);
and U2828 (N_2828,N_2138,N_1979);
nand U2829 (N_2829,N_2334,N_2006);
nand U2830 (N_2830,N_1900,N_2244);
nor U2831 (N_2831,N_2312,N_2006);
nand U2832 (N_2832,N_2108,N_1947);
and U2833 (N_2833,N_1950,N_1898);
and U2834 (N_2834,N_1968,N_1943);
or U2835 (N_2835,N_2328,N_1937);
nand U2836 (N_2836,N_1949,N_2343);
nor U2837 (N_2837,N_2050,N_1899);
or U2838 (N_2838,N_2011,N_1871);
or U2839 (N_2839,N_2125,N_2145);
nand U2840 (N_2840,N_2162,N_1942);
nand U2841 (N_2841,N_1968,N_2337);
nor U2842 (N_2842,N_2127,N_1855);
nand U2843 (N_2843,N_2093,N_1974);
or U2844 (N_2844,N_2386,N_2321);
and U2845 (N_2845,N_1819,N_1817);
nor U2846 (N_2846,N_2248,N_2086);
nand U2847 (N_2847,N_1908,N_2225);
and U2848 (N_2848,N_2397,N_2313);
nand U2849 (N_2849,N_2092,N_1934);
or U2850 (N_2850,N_2086,N_2234);
and U2851 (N_2851,N_2266,N_1827);
nand U2852 (N_2852,N_2240,N_1963);
and U2853 (N_2853,N_2091,N_2002);
and U2854 (N_2854,N_1863,N_2009);
and U2855 (N_2855,N_2256,N_1872);
nor U2856 (N_2856,N_2321,N_2239);
or U2857 (N_2857,N_2351,N_1983);
or U2858 (N_2858,N_2166,N_2228);
or U2859 (N_2859,N_1892,N_2345);
and U2860 (N_2860,N_2194,N_2121);
nor U2861 (N_2861,N_2269,N_1961);
nor U2862 (N_2862,N_2282,N_1856);
and U2863 (N_2863,N_1803,N_1831);
nor U2864 (N_2864,N_1898,N_2126);
or U2865 (N_2865,N_1869,N_2290);
and U2866 (N_2866,N_2200,N_2107);
and U2867 (N_2867,N_2235,N_2272);
nor U2868 (N_2868,N_1942,N_2251);
or U2869 (N_2869,N_1991,N_1864);
nand U2870 (N_2870,N_2321,N_2246);
or U2871 (N_2871,N_2130,N_1989);
or U2872 (N_2872,N_2364,N_2003);
nand U2873 (N_2873,N_2008,N_1952);
nand U2874 (N_2874,N_2153,N_2209);
nor U2875 (N_2875,N_2111,N_2369);
or U2876 (N_2876,N_1960,N_1919);
nor U2877 (N_2877,N_1919,N_2006);
nor U2878 (N_2878,N_2304,N_2278);
and U2879 (N_2879,N_2036,N_2244);
nand U2880 (N_2880,N_2333,N_1929);
and U2881 (N_2881,N_1955,N_1911);
and U2882 (N_2882,N_1984,N_2027);
and U2883 (N_2883,N_1944,N_1892);
and U2884 (N_2884,N_1817,N_2057);
nor U2885 (N_2885,N_1827,N_2061);
nor U2886 (N_2886,N_1848,N_2140);
or U2887 (N_2887,N_2172,N_2151);
nor U2888 (N_2888,N_1938,N_2354);
nand U2889 (N_2889,N_2035,N_2331);
and U2890 (N_2890,N_2129,N_2165);
nand U2891 (N_2891,N_2202,N_1959);
nor U2892 (N_2892,N_2083,N_2322);
nand U2893 (N_2893,N_1816,N_1993);
and U2894 (N_2894,N_1818,N_2221);
and U2895 (N_2895,N_2221,N_2257);
and U2896 (N_2896,N_2354,N_2000);
or U2897 (N_2897,N_1809,N_2149);
nand U2898 (N_2898,N_1944,N_2048);
or U2899 (N_2899,N_1980,N_2183);
and U2900 (N_2900,N_2012,N_2378);
or U2901 (N_2901,N_2015,N_1931);
nand U2902 (N_2902,N_1999,N_2301);
or U2903 (N_2903,N_2343,N_2151);
or U2904 (N_2904,N_2338,N_1807);
xor U2905 (N_2905,N_2085,N_1914);
and U2906 (N_2906,N_1991,N_1973);
and U2907 (N_2907,N_2010,N_2008);
or U2908 (N_2908,N_1928,N_2368);
or U2909 (N_2909,N_1938,N_1942);
nor U2910 (N_2910,N_1847,N_2067);
or U2911 (N_2911,N_2254,N_2145);
or U2912 (N_2912,N_2166,N_1999);
or U2913 (N_2913,N_1834,N_2138);
and U2914 (N_2914,N_2298,N_1898);
or U2915 (N_2915,N_1858,N_2208);
and U2916 (N_2916,N_1835,N_2290);
xor U2917 (N_2917,N_2215,N_1971);
nor U2918 (N_2918,N_1920,N_2157);
nor U2919 (N_2919,N_2011,N_2374);
and U2920 (N_2920,N_2282,N_2289);
nand U2921 (N_2921,N_2138,N_2014);
and U2922 (N_2922,N_2376,N_2265);
nand U2923 (N_2923,N_2129,N_2221);
or U2924 (N_2924,N_2367,N_1970);
or U2925 (N_2925,N_2384,N_1893);
nor U2926 (N_2926,N_2048,N_1925);
nand U2927 (N_2927,N_2233,N_2217);
nor U2928 (N_2928,N_2149,N_2230);
and U2929 (N_2929,N_2069,N_2242);
nor U2930 (N_2930,N_1833,N_2234);
nor U2931 (N_2931,N_2043,N_2044);
or U2932 (N_2932,N_2163,N_2133);
or U2933 (N_2933,N_1973,N_2137);
and U2934 (N_2934,N_1898,N_2217);
nor U2935 (N_2935,N_2130,N_2009);
nand U2936 (N_2936,N_2068,N_2330);
nand U2937 (N_2937,N_1966,N_1803);
or U2938 (N_2938,N_2225,N_2052);
nand U2939 (N_2939,N_1914,N_1979);
or U2940 (N_2940,N_2108,N_2274);
or U2941 (N_2941,N_2249,N_2308);
and U2942 (N_2942,N_2133,N_1866);
or U2943 (N_2943,N_2274,N_1876);
nor U2944 (N_2944,N_1816,N_1885);
or U2945 (N_2945,N_2133,N_2311);
nand U2946 (N_2946,N_1839,N_1828);
or U2947 (N_2947,N_2015,N_1840);
and U2948 (N_2948,N_2379,N_2293);
nor U2949 (N_2949,N_2226,N_1988);
nand U2950 (N_2950,N_2055,N_2147);
nor U2951 (N_2951,N_2165,N_2192);
and U2952 (N_2952,N_2376,N_2092);
nand U2953 (N_2953,N_1872,N_2075);
nor U2954 (N_2954,N_2084,N_2281);
and U2955 (N_2955,N_2012,N_2293);
nor U2956 (N_2956,N_2074,N_2042);
nand U2957 (N_2957,N_1963,N_2046);
and U2958 (N_2958,N_1812,N_1914);
or U2959 (N_2959,N_1864,N_1857);
or U2960 (N_2960,N_2033,N_2048);
or U2961 (N_2961,N_2170,N_2174);
or U2962 (N_2962,N_2357,N_2362);
xor U2963 (N_2963,N_1819,N_2131);
or U2964 (N_2964,N_1864,N_2297);
nand U2965 (N_2965,N_2042,N_1859);
or U2966 (N_2966,N_1826,N_2158);
xor U2967 (N_2967,N_2129,N_2345);
or U2968 (N_2968,N_1812,N_1962);
nor U2969 (N_2969,N_2133,N_1926);
and U2970 (N_2970,N_1815,N_2248);
nor U2971 (N_2971,N_1980,N_2002);
nand U2972 (N_2972,N_2353,N_1893);
nand U2973 (N_2973,N_1948,N_2197);
nand U2974 (N_2974,N_2369,N_2281);
and U2975 (N_2975,N_2259,N_1808);
and U2976 (N_2976,N_2128,N_2133);
or U2977 (N_2977,N_2297,N_2213);
and U2978 (N_2978,N_2068,N_2116);
nand U2979 (N_2979,N_2292,N_1802);
nor U2980 (N_2980,N_1826,N_2196);
and U2981 (N_2981,N_1814,N_2340);
nand U2982 (N_2982,N_2100,N_1838);
and U2983 (N_2983,N_1937,N_2249);
and U2984 (N_2984,N_2309,N_2193);
or U2985 (N_2985,N_2027,N_2040);
nor U2986 (N_2986,N_2286,N_2011);
nor U2987 (N_2987,N_1911,N_2316);
and U2988 (N_2988,N_2325,N_2003);
nor U2989 (N_2989,N_1859,N_2383);
nor U2990 (N_2990,N_2028,N_2284);
nand U2991 (N_2991,N_1938,N_1918);
nor U2992 (N_2992,N_2109,N_1896);
or U2993 (N_2993,N_2370,N_2225);
or U2994 (N_2994,N_1953,N_2230);
nand U2995 (N_2995,N_2196,N_2270);
nor U2996 (N_2996,N_1922,N_1918);
and U2997 (N_2997,N_2043,N_2169);
and U2998 (N_2998,N_2354,N_2100);
nor U2999 (N_2999,N_2186,N_2312);
and UO_0 (O_0,N_2483,N_2806);
nor UO_1 (O_1,N_2992,N_2593);
and UO_2 (O_2,N_2762,N_2929);
and UO_3 (O_3,N_2881,N_2428);
or UO_4 (O_4,N_2606,N_2818);
or UO_5 (O_5,N_2678,N_2566);
nor UO_6 (O_6,N_2877,N_2713);
nor UO_7 (O_7,N_2452,N_2447);
and UO_8 (O_8,N_2586,N_2807);
nor UO_9 (O_9,N_2965,N_2982);
or UO_10 (O_10,N_2578,N_2697);
nor UO_11 (O_11,N_2621,N_2766);
nand UO_12 (O_12,N_2505,N_2928);
nor UO_13 (O_13,N_2625,N_2976);
or UO_14 (O_14,N_2668,N_2801);
and UO_15 (O_15,N_2522,N_2635);
and UO_16 (O_16,N_2579,N_2799);
or UO_17 (O_17,N_2478,N_2465);
or UO_18 (O_18,N_2661,N_2845);
nor UO_19 (O_19,N_2690,N_2736);
or UO_20 (O_20,N_2826,N_2617);
and UO_21 (O_21,N_2676,N_2922);
nor UO_22 (O_22,N_2981,N_2842);
and UO_23 (O_23,N_2620,N_2864);
nand UO_24 (O_24,N_2879,N_2726);
or UO_25 (O_25,N_2665,N_2449);
nor UO_26 (O_26,N_2888,N_2411);
nor UO_27 (O_27,N_2567,N_2724);
and UO_28 (O_28,N_2471,N_2921);
nand UO_29 (O_29,N_2454,N_2918);
nor UO_30 (O_30,N_2557,N_2910);
and UO_31 (O_31,N_2605,N_2562);
or UO_32 (O_32,N_2413,N_2927);
and UO_33 (O_33,N_2470,N_2570);
nor UO_34 (O_34,N_2901,N_2462);
nand UO_35 (O_35,N_2775,N_2531);
and UO_36 (O_36,N_2804,N_2843);
or UO_37 (O_37,N_2402,N_2925);
or UO_38 (O_38,N_2651,N_2791);
nor UO_39 (O_39,N_2935,N_2916);
and UO_40 (O_40,N_2481,N_2688);
or UO_41 (O_41,N_2498,N_2718);
nor UO_42 (O_42,N_2978,N_2815);
nand UO_43 (O_43,N_2829,N_2455);
and UO_44 (O_44,N_2512,N_2953);
nand UO_45 (O_45,N_2565,N_2971);
or UO_46 (O_46,N_2754,N_2519);
nand UO_47 (O_47,N_2752,N_2735);
nor UO_48 (O_48,N_2527,N_2418);
and UO_49 (O_49,N_2896,N_2938);
nor UO_50 (O_50,N_2614,N_2407);
nor UO_51 (O_51,N_2420,N_2467);
and UO_52 (O_52,N_2995,N_2924);
and UO_53 (O_53,N_2627,N_2692);
nor UO_54 (O_54,N_2583,N_2933);
or UO_55 (O_55,N_2847,N_2488);
nand UO_56 (O_56,N_2573,N_2577);
nor UO_57 (O_57,N_2765,N_2968);
or UO_58 (O_58,N_2819,N_2850);
nand UO_59 (O_59,N_2874,N_2648);
nand UO_60 (O_60,N_2550,N_2542);
nand UO_61 (O_61,N_2739,N_2619);
or UO_62 (O_62,N_2670,N_2764);
nand UO_63 (O_63,N_2628,N_2997);
nand UO_64 (O_64,N_2825,N_2482);
or UO_65 (O_65,N_2949,N_2437);
nor UO_66 (O_66,N_2950,N_2930);
and UO_67 (O_67,N_2569,N_2689);
nand UO_68 (O_68,N_2464,N_2860);
or UO_69 (O_69,N_2975,N_2987);
nand UO_70 (O_70,N_2994,N_2841);
and UO_71 (O_71,N_2683,N_2876);
nand UO_72 (O_72,N_2400,N_2789);
or UO_73 (O_73,N_2497,N_2989);
nand UO_74 (O_74,N_2969,N_2908);
nand UO_75 (O_75,N_2664,N_2636);
or UO_76 (O_76,N_2787,N_2761);
and UO_77 (O_77,N_2687,N_2607);
or UO_78 (O_78,N_2778,N_2824);
and UO_79 (O_79,N_2433,N_2990);
nor UO_80 (O_80,N_2812,N_2538);
nor UO_81 (O_81,N_2532,N_2656);
nor UO_82 (O_82,N_2592,N_2721);
nand UO_83 (O_83,N_2962,N_2551);
nand UO_84 (O_84,N_2673,N_2750);
and UO_85 (O_85,N_2900,N_2536);
and UO_86 (O_86,N_2895,N_2558);
and UO_87 (O_87,N_2448,N_2897);
and UO_88 (O_88,N_2608,N_2612);
nand UO_89 (O_89,N_2491,N_2838);
nand UO_90 (O_90,N_2693,N_2459);
nor UO_91 (O_91,N_2514,N_2633);
or UO_92 (O_92,N_2823,N_2996);
nand UO_93 (O_93,N_2817,N_2554);
nor UO_94 (O_94,N_2870,N_2698);
and UO_95 (O_95,N_2469,N_2474);
nand UO_96 (O_96,N_2979,N_2759);
nand UO_97 (O_97,N_2903,N_2999);
nor UO_98 (O_98,N_2944,N_2832);
nand UO_99 (O_99,N_2463,N_2486);
and UO_100 (O_100,N_2731,N_2744);
nor UO_101 (O_101,N_2964,N_2575);
xor UO_102 (O_102,N_2917,N_2590);
nand UO_103 (O_103,N_2604,N_2827);
or UO_104 (O_104,N_2571,N_2779);
or UO_105 (O_105,N_2507,N_2476);
nand UO_106 (O_106,N_2539,N_2889);
nand UO_107 (O_107,N_2510,N_2568);
nor UO_108 (O_108,N_2553,N_2913);
nand UO_109 (O_109,N_2410,N_2423);
or UO_110 (O_110,N_2453,N_2403);
and UO_111 (O_111,N_2704,N_2937);
or UO_112 (O_112,N_2967,N_2501);
and UO_113 (O_113,N_2760,N_2591);
and UO_114 (O_114,N_2757,N_2525);
nand UO_115 (O_115,N_2408,N_2772);
or UO_116 (O_116,N_2416,N_2776);
nor UO_117 (O_117,N_2502,N_2645);
nor UO_118 (O_118,N_2419,N_2540);
or UO_119 (O_119,N_2667,N_2626);
nor UO_120 (O_120,N_2638,N_2641);
and UO_121 (O_121,N_2973,N_2631);
nor UO_122 (O_122,N_2868,N_2809);
nor UO_123 (O_123,N_2485,N_2686);
and UO_124 (O_124,N_2831,N_2743);
and UO_125 (O_125,N_2839,N_2887);
nand UO_126 (O_126,N_2785,N_2492);
nor UO_127 (O_127,N_2833,N_2884);
nand UO_128 (O_128,N_2909,N_2820);
nand UO_129 (O_129,N_2977,N_2873);
nand UO_130 (O_130,N_2438,N_2948);
or UO_131 (O_131,N_2882,N_2442);
or UO_132 (O_132,N_2797,N_2646);
nor UO_133 (O_133,N_2998,N_2706);
and UO_134 (O_134,N_2985,N_2931);
or UO_135 (O_135,N_2669,N_2986);
nand UO_136 (O_136,N_2563,N_2749);
nand UO_137 (O_137,N_2640,N_2781);
or UO_138 (O_138,N_2970,N_2880);
and UO_139 (O_139,N_2600,N_2770);
and UO_140 (O_140,N_2663,N_2537);
nand UO_141 (O_141,N_2649,N_2814);
and UO_142 (O_142,N_2729,N_2763);
and UO_143 (O_143,N_2677,N_2701);
or UO_144 (O_144,N_2616,N_2461);
nor UO_145 (O_145,N_2800,N_2601);
nor UO_146 (O_146,N_2871,N_2533);
nand UO_147 (O_147,N_2867,N_2862);
and UO_148 (O_148,N_2598,N_2431);
nor UO_149 (O_149,N_2782,N_2658);
nand UO_150 (O_150,N_2587,N_2624);
and UO_151 (O_151,N_2803,N_2836);
nor UO_152 (O_152,N_2556,N_2458);
nand UO_153 (O_153,N_2585,N_2639);
nor UO_154 (O_154,N_2541,N_2523);
nand UO_155 (O_155,N_2849,N_2786);
and UO_156 (O_156,N_2712,N_2615);
nor UO_157 (O_157,N_2495,N_2682);
and UO_158 (O_158,N_2572,N_2508);
and UO_159 (O_159,N_2517,N_2883);
or UO_160 (O_160,N_2430,N_2574);
and UO_161 (O_161,N_2655,N_2866);
or UO_162 (O_162,N_2552,N_2777);
nand UO_163 (O_163,N_2709,N_2936);
nand UO_164 (O_164,N_2952,N_2675);
or UO_165 (O_165,N_2886,N_2424);
nor UO_166 (O_166,N_2629,N_2773);
or UO_167 (O_167,N_2544,N_2691);
or UO_168 (O_168,N_2429,N_2644);
nor UO_169 (O_169,N_2548,N_2679);
and UO_170 (O_170,N_2671,N_2623);
and UO_171 (O_171,N_2802,N_2466);
and UO_172 (O_172,N_2526,N_2984);
and UO_173 (O_173,N_2659,N_2769);
or UO_174 (O_174,N_2489,N_2504);
or UO_175 (O_175,N_2810,N_2611);
or UO_176 (O_176,N_2564,N_2852);
or UO_177 (O_177,N_2496,N_2549);
or UO_178 (O_178,N_2920,N_2932);
and UO_179 (O_179,N_2945,N_2710);
nand UO_180 (O_180,N_2946,N_2794);
and UO_181 (O_181,N_2436,N_2748);
nand UO_182 (O_182,N_2939,N_2840);
nor UO_183 (O_183,N_2457,N_2740);
or UO_184 (O_184,N_2584,N_2830);
nor UO_185 (O_185,N_2811,N_2609);
nand UO_186 (O_186,N_2595,N_2406);
and UO_187 (O_187,N_2923,N_2943);
nand UO_188 (O_188,N_2518,N_2561);
nor UO_189 (O_189,N_2893,N_2798);
and UO_190 (O_190,N_2894,N_2737);
and UO_191 (O_191,N_2503,N_2892);
nor UO_192 (O_192,N_2869,N_2912);
nor UO_193 (O_193,N_2974,N_2741);
nor UO_194 (O_194,N_2711,N_2906);
and UO_195 (O_195,N_2947,N_2404);
nand UO_196 (O_196,N_2813,N_2528);
nand UO_197 (O_197,N_2911,N_2926);
nand UO_198 (O_198,N_2432,N_2768);
or UO_199 (O_199,N_2699,N_2632);
nor UO_200 (O_200,N_2630,N_2755);
or UO_201 (O_201,N_2942,N_2914);
and UO_202 (O_202,N_2951,N_2865);
nor UO_203 (O_203,N_2854,N_2547);
and UO_204 (O_204,N_2828,N_2720);
nor UO_205 (O_205,N_2618,N_2705);
and UO_206 (O_206,N_2837,N_2793);
or UO_207 (O_207,N_2796,N_2746);
or UO_208 (O_208,N_2473,N_2515);
or UO_209 (O_209,N_2634,N_2719);
or UO_210 (O_210,N_2784,N_2652);
or UO_211 (O_211,N_2780,N_2961);
and UO_212 (O_212,N_2956,N_2477);
or UO_213 (O_213,N_2674,N_2885);
nor UO_214 (O_214,N_2816,N_2940);
and UO_215 (O_215,N_2622,N_2941);
and UO_216 (O_216,N_2958,N_2957);
nand UO_217 (O_217,N_2702,N_2460);
and UO_218 (O_218,N_2808,N_2468);
nor UO_219 (O_219,N_2848,N_2555);
and UO_220 (O_220,N_2963,N_2899);
or UO_221 (O_221,N_2439,N_2855);
or UO_222 (O_222,N_2694,N_2955);
nand UO_223 (O_223,N_2657,N_2907);
and UO_224 (O_224,N_2890,N_2530);
or UO_225 (O_225,N_2560,N_2988);
nand UO_226 (O_226,N_2723,N_2753);
xnor UO_227 (O_227,N_2576,N_2446);
nand UO_228 (O_228,N_2412,N_2602);
nand UO_229 (O_229,N_2653,N_2422);
nand UO_230 (O_230,N_2822,N_2745);
and UO_231 (O_231,N_2851,N_2844);
nand UO_232 (O_232,N_2756,N_2805);
nor UO_233 (O_233,N_2733,N_2445);
and UO_234 (O_234,N_2500,N_2863);
nor UO_235 (O_235,N_2654,N_2613);
and UO_236 (O_236,N_2487,N_2513);
and UO_237 (O_237,N_2858,N_2727);
nor UO_238 (O_238,N_2660,N_2685);
or UO_239 (O_239,N_2767,N_2856);
nor UO_240 (O_240,N_2788,N_2915);
nand UO_241 (O_241,N_2730,N_2680);
nand UO_242 (O_242,N_2742,N_2588);
or UO_243 (O_243,N_2905,N_2747);
nand UO_244 (O_244,N_2993,N_2472);
xor UO_245 (O_245,N_2405,N_2603);
or UO_246 (O_246,N_2451,N_2891);
and UO_247 (O_247,N_2425,N_2716);
nor UO_248 (O_248,N_2734,N_2738);
or UO_249 (O_249,N_2700,N_2919);
and UO_250 (O_250,N_2696,N_2427);
nand UO_251 (O_251,N_2494,N_2972);
nor UO_252 (O_252,N_2511,N_2835);
nand UO_253 (O_253,N_2898,N_2516);
nor UO_254 (O_254,N_2834,N_2792);
nor UO_255 (O_255,N_2934,N_2846);
and UO_256 (O_256,N_2875,N_2417);
nand UO_257 (O_257,N_2904,N_2681);
nor UO_258 (O_258,N_2450,N_2695);
or UO_259 (O_259,N_2581,N_2758);
or UO_260 (O_260,N_2966,N_2751);
and UO_261 (O_261,N_2524,N_2983);
and UO_262 (O_262,N_2703,N_2857);
xnor UO_263 (O_263,N_2443,N_2859);
or UO_264 (O_264,N_2545,N_2534);
nor UO_265 (O_265,N_2401,N_2421);
nor UO_266 (O_266,N_2684,N_2980);
nand UO_267 (O_267,N_2434,N_2959);
and UO_268 (O_268,N_2861,N_2774);
nand UO_269 (O_269,N_2444,N_2415);
nor UO_270 (O_270,N_2441,N_2662);
nand UO_271 (O_271,N_2509,N_2535);
or UO_272 (O_272,N_2506,N_2484);
nand UO_273 (O_273,N_2580,N_2546);
nor UO_274 (O_274,N_2732,N_2435);
nand UO_275 (O_275,N_2414,N_2960);
and UO_276 (O_276,N_2821,N_2582);
and UO_277 (O_277,N_2878,N_2795);
or UO_278 (O_278,N_2650,N_2479);
nand UO_279 (O_279,N_2493,N_2637);
nor UO_280 (O_280,N_2475,N_2599);
nand UO_281 (O_281,N_2643,N_2783);
or UO_282 (O_282,N_2589,N_2672);
and UO_283 (O_283,N_2728,N_2642);
nand UO_284 (O_284,N_2771,N_2543);
nor UO_285 (O_285,N_2440,N_2717);
and UO_286 (O_286,N_2499,N_2872);
or UO_287 (O_287,N_2559,N_2666);
nand UO_288 (O_288,N_2521,N_2902);
and UO_289 (O_289,N_2596,N_2954);
nor UO_290 (O_290,N_2456,N_2722);
nand UO_291 (O_291,N_2991,N_2490);
or UO_292 (O_292,N_2715,N_2520);
and UO_293 (O_293,N_2708,N_2597);
and UO_294 (O_294,N_2714,N_2853);
nor UO_295 (O_295,N_2426,N_2790);
nor UO_296 (O_296,N_2480,N_2647);
and UO_297 (O_297,N_2725,N_2707);
nand UO_298 (O_298,N_2409,N_2594);
nor UO_299 (O_299,N_2610,N_2529);
or UO_300 (O_300,N_2629,N_2641);
nand UO_301 (O_301,N_2755,N_2876);
and UO_302 (O_302,N_2960,N_2910);
or UO_303 (O_303,N_2429,N_2451);
nor UO_304 (O_304,N_2829,N_2673);
or UO_305 (O_305,N_2804,N_2484);
nand UO_306 (O_306,N_2945,N_2837);
or UO_307 (O_307,N_2723,N_2937);
nand UO_308 (O_308,N_2654,N_2500);
and UO_309 (O_309,N_2877,N_2875);
and UO_310 (O_310,N_2698,N_2644);
nand UO_311 (O_311,N_2892,N_2735);
and UO_312 (O_312,N_2590,N_2677);
nand UO_313 (O_313,N_2835,N_2425);
or UO_314 (O_314,N_2650,N_2469);
and UO_315 (O_315,N_2920,N_2419);
xnor UO_316 (O_316,N_2523,N_2712);
nand UO_317 (O_317,N_2540,N_2405);
and UO_318 (O_318,N_2683,N_2544);
or UO_319 (O_319,N_2626,N_2579);
or UO_320 (O_320,N_2461,N_2854);
nand UO_321 (O_321,N_2688,N_2792);
or UO_322 (O_322,N_2614,N_2942);
nor UO_323 (O_323,N_2857,N_2890);
nor UO_324 (O_324,N_2807,N_2976);
nor UO_325 (O_325,N_2658,N_2743);
nand UO_326 (O_326,N_2990,N_2437);
or UO_327 (O_327,N_2751,N_2627);
nand UO_328 (O_328,N_2660,N_2722);
nor UO_329 (O_329,N_2721,N_2919);
nor UO_330 (O_330,N_2575,N_2736);
or UO_331 (O_331,N_2993,N_2892);
or UO_332 (O_332,N_2800,N_2732);
and UO_333 (O_333,N_2923,N_2478);
or UO_334 (O_334,N_2500,N_2669);
nand UO_335 (O_335,N_2613,N_2525);
and UO_336 (O_336,N_2655,N_2565);
nand UO_337 (O_337,N_2528,N_2426);
nand UO_338 (O_338,N_2973,N_2796);
and UO_339 (O_339,N_2599,N_2946);
nor UO_340 (O_340,N_2778,N_2471);
nor UO_341 (O_341,N_2482,N_2472);
nor UO_342 (O_342,N_2414,N_2431);
or UO_343 (O_343,N_2559,N_2718);
and UO_344 (O_344,N_2525,N_2431);
nor UO_345 (O_345,N_2916,N_2992);
or UO_346 (O_346,N_2808,N_2761);
or UO_347 (O_347,N_2840,N_2827);
or UO_348 (O_348,N_2483,N_2847);
nand UO_349 (O_349,N_2559,N_2480);
nor UO_350 (O_350,N_2625,N_2488);
or UO_351 (O_351,N_2554,N_2429);
nand UO_352 (O_352,N_2426,N_2463);
nor UO_353 (O_353,N_2807,N_2997);
nand UO_354 (O_354,N_2669,N_2933);
nor UO_355 (O_355,N_2460,N_2602);
nand UO_356 (O_356,N_2868,N_2735);
or UO_357 (O_357,N_2662,N_2912);
nand UO_358 (O_358,N_2535,N_2781);
or UO_359 (O_359,N_2818,N_2584);
and UO_360 (O_360,N_2466,N_2656);
and UO_361 (O_361,N_2650,N_2531);
and UO_362 (O_362,N_2587,N_2901);
nand UO_363 (O_363,N_2899,N_2483);
nand UO_364 (O_364,N_2498,N_2517);
xnor UO_365 (O_365,N_2436,N_2552);
nor UO_366 (O_366,N_2892,N_2531);
or UO_367 (O_367,N_2560,N_2496);
and UO_368 (O_368,N_2753,N_2968);
or UO_369 (O_369,N_2475,N_2697);
nand UO_370 (O_370,N_2636,N_2467);
nand UO_371 (O_371,N_2703,N_2713);
nor UO_372 (O_372,N_2440,N_2926);
nand UO_373 (O_373,N_2631,N_2412);
and UO_374 (O_374,N_2594,N_2505);
and UO_375 (O_375,N_2627,N_2982);
or UO_376 (O_376,N_2540,N_2764);
nand UO_377 (O_377,N_2514,N_2731);
and UO_378 (O_378,N_2994,N_2918);
nand UO_379 (O_379,N_2713,N_2553);
nand UO_380 (O_380,N_2785,N_2548);
nand UO_381 (O_381,N_2426,N_2682);
or UO_382 (O_382,N_2824,N_2524);
nand UO_383 (O_383,N_2720,N_2987);
nand UO_384 (O_384,N_2870,N_2496);
nor UO_385 (O_385,N_2663,N_2776);
nor UO_386 (O_386,N_2763,N_2476);
and UO_387 (O_387,N_2669,N_2433);
nand UO_388 (O_388,N_2719,N_2995);
or UO_389 (O_389,N_2910,N_2829);
nor UO_390 (O_390,N_2577,N_2659);
or UO_391 (O_391,N_2742,N_2569);
nand UO_392 (O_392,N_2707,N_2710);
nor UO_393 (O_393,N_2556,N_2530);
and UO_394 (O_394,N_2775,N_2883);
nand UO_395 (O_395,N_2633,N_2976);
or UO_396 (O_396,N_2747,N_2924);
nor UO_397 (O_397,N_2932,N_2565);
nand UO_398 (O_398,N_2521,N_2626);
and UO_399 (O_399,N_2485,N_2885);
nand UO_400 (O_400,N_2725,N_2537);
and UO_401 (O_401,N_2595,N_2977);
and UO_402 (O_402,N_2550,N_2468);
and UO_403 (O_403,N_2544,N_2706);
nand UO_404 (O_404,N_2478,N_2627);
and UO_405 (O_405,N_2893,N_2653);
nor UO_406 (O_406,N_2697,N_2720);
nand UO_407 (O_407,N_2543,N_2566);
nor UO_408 (O_408,N_2449,N_2688);
and UO_409 (O_409,N_2449,N_2553);
and UO_410 (O_410,N_2783,N_2960);
nor UO_411 (O_411,N_2990,N_2425);
and UO_412 (O_412,N_2840,N_2584);
and UO_413 (O_413,N_2949,N_2516);
nand UO_414 (O_414,N_2696,N_2730);
nor UO_415 (O_415,N_2967,N_2436);
nand UO_416 (O_416,N_2822,N_2508);
nand UO_417 (O_417,N_2821,N_2972);
and UO_418 (O_418,N_2564,N_2769);
nand UO_419 (O_419,N_2714,N_2640);
or UO_420 (O_420,N_2903,N_2666);
or UO_421 (O_421,N_2893,N_2764);
and UO_422 (O_422,N_2933,N_2475);
or UO_423 (O_423,N_2884,N_2999);
nand UO_424 (O_424,N_2755,N_2641);
and UO_425 (O_425,N_2800,N_2653);
nor UO_426 (O_426,N_2943,N_2973);
nand UO_427 (O_427,N_2644,N_2712);
nand UO_428 (O_428,N_2622,N_2647);
nand UO_429 (O_429,N_2540,N_2859);
nor UO_430 (O_430,N_2943,N_2466);
and UO_431 (O_431,N_2416,N_2792);
nand UO_432 (O_432,N_2575,N_2804);
and UO_433 (O_433,N_2946,N_2400);
xnor UO_434 (O_434,N_2555,N_2781);
or UO_435 (O_435,N_2695,N_2879);
nand UO_436 (O_436,N_2856,N_2606);
nor UO_437 (O_437,N_2984,N_2913);
and UO_438 (O_438,N_2707,N_2949);
nand UO_439 (O_439,N_2995,N_2548);
or UO_440 (O_440,N_2603,N_2577);
xor UO_441 (O_441,N_2897,N_2760);
or UO_442 (O_442,N_2440,N_2561);
nor UO_443 (O_443,N_2471,N_2701);
and UO_444 (O_444,N_2823,N_2868);
nand UO_445 (O_445,N_2573,N_2605);
and UO_446 (O_446,N_2505,N_2556);
nand UO_447 (O_447,N_2506,N_2643);
or UO_448 (O_448,N_2813,N_2506);
and UO_449 (O_449,N_2656,N_2936);
or UO_450 (O_450,N_2404,N_2967);
nor UO_451 (O_451,N_2785,N_2504);
nor UO_452 (O_452,N_2907,N_2557);
nor UO_453 (O_453,N_2633,N_2464);
and UO_454 (O_454,N_2486,N_2714);
nor UO_455 (O_455,N_2990,N_2529);
nor UO_456 (O_456,N_2471,N_2565);
nand UO_457 (O_457,N_2709,N_2954);
and UO_458 (O_458,N_2698,N_2919);
and UO_459 (O_459,N_2648,N_2407);
nor UO_460 (O_460,N_2910,N_2612);
nand UO_461 (O_461,N_2646,N_2804);
or UO_462 (O_462,N_2800,N_2585);
nor UO_463 (O_463,N_2669,N_2882);
or UO_464 (O_464,N_2685,N_2407);
nor UO_465 (O_465,N_2674,N_2657);
or UO_466 (O_466,N_2893,N_2805);
and UO_467 (O_467,N_2768,N_2435);
or UO_468 (O_468,N_2880,N_2954);
nand UO_469 (O_469,N_2481,N_2659);
and UO_470 (O_470,N_2997,N_2939);
and UO_471 (O_471,N_2883,N_2926);
and UO_472 (O_472,N_2789,N_2566);
nand UO_473 (O_473,N_2405,N_2658);
nand UO_474 (O_474,N_2871,N_2780);
nor UO_475 (O_475,N_2783,N_2466);
nor UO_476 (O_476,N_2414,N_2583);
and UO_477 (O_477,N_2770,N_2717);
nor UO_478 (O_478,N_2878,N_2606);
and UO_479 (O_479,N_2823,N_2611);
nand UO_480 (O_480,N_2510,N_2923);
and UO_481 (O_481,N_2715,N_2993);
or UO_482 (O_482,N_2899,N_2420);
nand UO_483 (O_483,N_2850,N_2535);
nor UO_484 (O_484,N_2903,N_2610);
nor UO_485 (O_485,N_2668,N_2434);
nand UO_486 (O_486,N_2655,N_2727);
and UO_487 (O_487,N_2723,N_2466);
or UO_488 (O_488,N_2676,N_2578);
and UO_489 (O_489,N_2629,N_2964);
and UO_490 (O_490,N_2744,N_2974);
nand UO_491 (O_491,N_2818,N_2547);
and UO_492 (O_492,N_2475,N_2559);
and UO_493 (O_493,N_2465,N_2574);
nand UO_494 (O_494,N_2532,N_2899);
or UO_495 (O_495,N_2915,N_2824);
nand UO_496 (O_496,N_2569,N_2771);
or UO_497 (O_497,N_2971,N_2935);
or UO_498 (O_498,N_2874,N_2947);
nor UO_499 (O_499,N_2908,N_2763);
endmodule