module basic_750_5000_1000_25_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_387,In_596);
nor U1 (N_1,In_498,In_367);
xor U2 (N_2,In_46,In_144);
nor U3 (N_3,In_126,In_523);
nand U4 (N_4,In_518,In_339);
nor U5 (N_5,In_43,In_592);
nor U6 (N_6,In_431,In_478);
and U7 (N_7,In_652,In_270);
and U8 (N_8,In_469,In_665);
nor U9 (N_9,In_409,In_308);
nor U10 (N_10,In_325,In_109);
or U11 (N_11,In_334,In_646);
nor U12 (N_12,In_280,In_193);
xnor U13 (N_13,In_50,In_128);
and U14 (N_14,In_602,In_224);
nor U15 (N_15,In_163,In_636);
xnor U16 (N_16,In_98,In_371);
xnor U17 (N_17,In_1,In_623);
nor U18 (N_18,In_451,In_385);
nand U19 (N_19,In_117,In_737);
nor U20 (N_20,In_169,In_287);
or U21 (N_21,In_439,In_87);
nor U22 (N_22,In_324,In_356);
or U23 (N_23,In_400,In_353);
or U24 (N_24,In_668,In_233);
or U25 (N_25,In_634,In_45);
nand U26 (N_26,In_4,In_140);
nand U27 (N_27,In_440,In_532);
nand U28 (N_28,In_467,In_729);
nand U29 (N_29,In_115,In_395);
and U30 (N_30,In_514,In_305);
and U31 (N_31,In_146,In_41);
nand U32 (N_32,In_640,In_338);
or U33 (N_33,In_494,In_554);
nor U34 (N_34,In_534,In_249);
xnor U35 (N_35,In_205,In_165);
and U36 (N_36,In_706,In_317);
or U37 (N_37,In_717,In_629);
and U38 (N_38,In_113,In_522);
nor U39 (N_39,In_340,In_747);
nor U40 (N_40,In_226,In_227);
or U41 (N_41,In_282,In_502);
nand U42 (N_42,In_506,In_656);
nor U43 (N_43,In_734,In_242);
nand U44 (N_44,In_357,In_670);
xnor U45 (N_45,In_120,In_8);
nor U46 (N_46,In_61,In_276);
nor U47 (N_47,In_574,In_66);
nand U48 (N_48,In_289,In_172);
nor U49 (N_49,In_582,In_157);
or U50 (N_50,In_654,In_265);
xor U51 (N_51,In_175,In_277);
nor U52 (N_52,In_295,In_208);
nand U53 (N_53,In_296,In_151);
nor U54 (N_54,In_560,In_192);
or U55 (N_55,In_7,In_627);
nor U56 (N_56,In_472,In_487);
nand U57 (N_57,In_744,In_139);
nand U58 (N_58,In_229,In_369);
nand U59 (N_59,In_373,In_630);
nor U60 (N_60,In_633,In_631);
nor U61 (N_61,In_632,In_490);
nor U62 (N_62,In_118,In_228);
and U63 (N_63,In_189,In_283);
nor U64 (N_64,In_86,In_37);
nand U65 (N_65,In_692,In_589);
or U66 (N_66,In_417,In_9);
nand U67 (N_67,In_444,In_588);
xnor U68 (N_68,In_424,In_569);
or U69 (N_69,In_655,In_218);
nor U70 (N_70,In_606,In_637);
nand U71 (N_71,In_314,In_438);
nand U72 (N_72,In_136,In_465);
nor U73 (N_73,In_191,In_455);
or U74 (N_74,In_694,In_161);
or U75 (N_75,In_206,In_272);
xor U76 (N_76,In_69,In_20);
and U77 (N_77,In_111,In_515);
and U78 (N_78,In_285,In_59);
or U79 (N_79,In_448,In_557);
nor U80 (N_80,In_368,In_407);
nand U81 (N_81,In_209,In_6);
or U82 (N_82,In_56,In_318);
and U83 (N_83,In_330,In_129);
nand U84 (N_84,In_311,In_306);
nor U85 (N_85,In_708,In_57);
xor U86 (N_86,In_695,In_466);
and U87 (N_87,In_432,In_540);
nand U88 (N_88,In_718,In_32);
xor U89 (N_89,In_132,In_658);
or U90 (N_90,In_99,In_29);
and U91 (N_91,In_122,In_578);
and U92 (N_92,In_573,In_667);
and U93 (N_93,In_164,In_275);
nor U94 (N_94,In_689,In_457);
or U95 (N_95,In_571,In_619);
nor U96 (N_96,In_89,In_664);
nor U97 (N_97,In_396,In_178);
and U98 (N_98,In_669,In_649);
nand U99 (N_99,In_92,In_549);
nand U100 (N_100,In_564,In_452);
and U101 (N_101,In_47,In_732);
and U102 (N_102,In_555,In_435);
or U103 (N_103,In_67,In_60);
and U104 (N_104,In_595,In_131);
and U105 (N_105,In_547,In_240);
and U106 (N_106,In_468,In_323);
nand U107 (N_107,In_359,In_261);
nor U108 (N_108,In_418,In_587);
nor U109 (N_109,In_450,In_106);
and U110 (N_110,In_74,In_464);
and U111 (N_111,In_121,In_603);
or U112 (N_112,In_470,In_214);
and U113 (N_113,In_365,In_590);
and U114 (N_114,In_671,In_13);
or U115 (N_115,In_543,In_95);
and U116 (N_116,In_181,In_358);
or U117 (N_117,In_347,In_421);
nor U118 (N_118,In_625,In_71);
nand U119 (N_119,In_23,In_516);
or U120 (N_120,In_705,In_363);
and U121 (N_121,In_138,In_576);
nand U122 (N_122,In_538,In_458);
or U123 (N_123,In_196,In_412);
nor U124 (N_124,In_133,In_537);
nor U125 (N_125,In_608,In_666);
and U126 (N_126,In_374,In_195);
and U127 (N_127,In_350,In_408);
nand U128 (N_128,In_610,In_416);
nor U129 (N_129,In_645,In_93);
and U130 (N_130,In_94,In_333);
or U131 (N_131,In_217,In_279);
nor U132 (N_132,In_362,In_425);
and U133 (N_133,In_220,In_551);
and U134 (N_134,In_171,In_28);
or U135 (N_135,In_449,In_507);
nand U136 (N_136,In_264,In_294);
and U137 (N_137,In_79,In_326);
and U138 (N_138,In_320,In_179);
nor U139 (N_139,In_379,In_236);
nand U140 (N_140,In_263,In_488);
or U141 (N_141,In_696,In_268);
and U142 (N_142,In_745,In_319);
nand U143 (N_143,In_251,In_186);
nor U144 (N_144,In_419,In_401);
xor U145 (N_145,In_716,In_476);
nor U146 (N_146,In_485,In_75);
or U147 (N_147,In_710,In_552);
and U148 (N_148,In_513,In_415);
or U149 (N_149,In_39,In_651);
nand U150 (N_150,In_512,In_255);
and U151 (N_151,In_199,In_130);
nor U152 (N_152,In_230,In_693);
or U153 (N_153,In_124,In_313);
and U154 (N_154,In_386,In_200);
nand U155 (N_155,In_360,In_125);
and U156 (N_156,In_536,In_245);
nor U157 (N_157,In_674,In_375);
xnor U158 (N_158,In_723,In_720);
nand U159 (N_159,In_486,In_650);
and U160 (N_160,In_341,In_137);
nand U161 (N_161,In_127,In_351);
nor U162 (N_162,In_613,In_10);
and U163 (N_163,In_624,In_70);
nand U164 (N_164,In_489,In_315);
nor U165 (N_165,In_594,In_198);
and U166 (N_166,In_604,In_119);
nand U167 (N_167,In_90,In_447);
nor U168 (N_168,In_626,In_382);
nor U169 (N_169,In_31,In_662);
nor U170 (N_170,In_687,In_539);
and U171 (N_171,In_611,In_302);
or U172 (N_172,In_65,In_724);
and U173 (N_173,In_390,In_202);
and U174 (N_174,In_85,In_167);
xnor U175 (N_175,In_445,In_474);
and U176 (N_176,In_591,In_568);
or U177 (N_177,In_252,In_82);
nor U178 (N_178,In_135,In_453);
nor U179 (N_179,In_101,In_410);
nand U180 (N_180,In_150,In_316);
xor U181 (N_181,In_584,In_701);
and U182 (N_182,In_511,In_484);
or U183 (N_183,In_677,In_258);
xor U184 (N_184,In_617,In_566);
nor U185 (N_185,In_53,In_598);
nand U186 (N_186,In_682,In_612);
or U187 (N_187,In_739,In_54);
and U188 (N_188,In_309,In_620);
and U189 (N_189,In_746,In_149);
nor U190 (N_190,In_736,In_562);
or U191 (N_191,In_232,In_535);
and U192 (N_192,In_436,In_203);
and U193 (N_193,In_81,In_530);
or U194 (N_194,In_712,In_225);
or U195 (N_195,In_68,In_256);
or U196 (N_196,In_212,In_491);
xnor U197 (N_197,In_678,In_621);
or U198 (N_198,In_709,In_288);
or U199 (N_199,In_681,In_103);
and U200 (N_200,N_28,In_471);
or U201 (N_201,N_54,In_703);
and U202 (N_202,In_370,In_123);
or U203 (N_203,In_607,N_47);
nand U204 (N_204,In_411,In_749);
nand U205 (N_205,In_312,N_98);
nand U206 (N_206,In_394,In_194);
nor U207 (N_207,N_86,In_567);
xnor U208 (N_208,N_129,N_51);
nand U209 (N_209,In_583,In_173);
nor U210 (N_210,N_104,In_40);
nor U211 (N_211,In_461,In_727);
and U212 (N_212,In_672,In_17);
and U213 (N_213,N_30,In_248);
nor U214 (N_214,In_542,N_7);
and U215 (N_215,In_231,In_235);
nor U216 (N_216,In_699,In_241);
or U217 (N_217,In_378,In_273);
or U218 (N_218,N_46,In_345);
nor U219 (N_219,In_433,N_151);
xor U220 (N_220,In_473,In_211);
nor U221 (N_221,N_146,In_177);
nor U222 (N_222,In_354,In_336);
nor U223 (N_223,N_65,N_69);
nand U224 (N_224,N_153,In_180);
nor U225 (N_225,N_147,N_44);
or U226 (N_226,N_143,In_600);
or U227 (N_227,N_87,N_63);
or U228 (N_228,In_643,N_29);
nor U229 (N_229,N_128,N_97);
xor U230 (N_230,In_748,In_11);
nand U231 (N_231,N_174,In_735);
nand U232 (N_232,In_266,N_183);
or U233 (N_233,In_24,N_64);
nand U234 (N_234,In_2,In_274);
or U235 (N_235,In_381,In_77);
or U236 (N_236,In_648,In_361);
xnor U237 (N_237,In_237,N_42);
nor U238 (N_238,In_586,In_286);
or U239 (N_239,In_391,N_50);
nor U240 (N_240,In_114,In_52);
or U241 (N_241,In_337,In_559);
xor U242 (N_242,N_74,In_254);
nor U243 (N_243,In_215,N_32);
and U244 (N_244,In_392,In_281);
nor U245 (N_245,In_257,In_174);
nand U246 (N_246,In_344,In_153);
and U247 (N_247,N_145,In_501);
and U248 (N_248,N_23,N_77);
or U249 (N_249,In_335,In_247);
and U250 (N_250,N_31,In_221);
nor U251 (N_251,N_173,In_580);
nor U252 (N_252,N_114,In_141);
or U253 (N_253,In_524,In_558);
or U254 (N_254,In_572,In_622);
nor U255 (N_255,In_207,In_609);
and U256 (N_256,In_721,N_17);
or U257 (N_257,N_1,In_553);
or U258 (N_258,In_366,N_101);
nand U259 (N_259,In_0,N_112);
and U260 (N_260,N_109,In_188);
or U261 (N_261,In_154,N_21);
nor U262 (N_262,In_22,In_742);
nand U263 (N_263,In_73,In_176);
nor U264 (N_264,In_641,N_144);
or U265 (N_265,N_24,N_89);
nor U266 (N_266,In_342,N_190);
nor U267 (N_267,In_644,In_147);
nand U268 (N_268,In_38,In_104);
nand U269 (N_269,N_139,N_177);
xnor U270 (N_270,N_90,In_628);
nand U271 (N_271,In_480,In_499);
nand U272 (N_272,In_26,In_690);
nor U273 (N_273,In_18,In_372);
xnor U274 (N_274,In_639,In_715);
or U275 (N_275,In_5,In_300);
nand U276 (N_276,In_441,N_166);
and U277 (N_277,N_93,In_505);
nor U278 (N_278,N_12,In_204);
or U279 (N_279,In_322,In_91);
xor U280 (N_280,In_223,In_76);
and U281 (N_281,In_327,In_49);
xnor U282 (N_282,In_349,In_346);
xor U283 (N_283,In_533,In_714);
or U284 (N_284,In_399,N_102);
or U285 (N_285,In_548,In_243);
or U286 (N_286,In_679,In_145);
or U287 (N_287,In_635,In_605);
nand U288 (N_288,In_546,In_166);
and U289 (N_289,N_136,In_529);
nand U290 (N_290,In_234,In_743);
and U291 (N_291,N_71,N_161);
xor U292 (N_292,In_437,In_201);
nand U293 (N_293,N_25,N_194);
nand U294 (N_294,In_544,In_48);
nand U295 (N_295,N_176,In_72);
or U296 (N_296,In_577,N_178);
nand U297 (N_297,N_8,In_383);
xnor U298 (N_298,In_526,N_111);
or U299 (N_299,N_19,N_66);
and U300 (N_300,In_663,In_238);
nand U301 (N_301,In_707,In_301);
or U302 (N_302,N_164,In_269);
nand U303 (N_303,In_618,In_397);
or U304 (N_304,In_393,In_58);
and U305 (N_305,In_152,N_4);
or U306 (N_306,In_25,In_427);
and U307 (N_307,In_730,N_2);
nand U308 (N_308,N_148,N_160);
xor U309 (N_309,N_76,In_642);
or U310 (N_310,In_293,N_192);
and U311 (N_311,N_172,In_691);
xor U312 (N_312,In_570,In_414);
nand U313 (N_313,In_297,In_443);
xnor U314 (N_314,N_13,In_291);
or U315 (N_315,In_3,In_481);
nor U316 (N_316,In_298,In_83);
nor U317 (N_317,N_67,In_680);
nand U318 (N_318,N_105,In_384);
and U319 (N_319,In_100,In_290);
and U320 (N_320,In_422,N_122);
nor U321 (N_321,In_711,N_180);
and U322 (N_322,N_167,In_517);
nor U323 (N_323,N_198,N_33);
and U324 (N_324,N_41,N_20);
or U325 (N_325,N_120,In_700);
nand U326 (N_326,In_599,In_62);
and U327 (N_327,In_244,In_376);
or U328 (N_328,N_57,N_40);
nand U329 (N_329,In_246,N_11);
nand U330 (N_330,N_94,N_156);
and U331 (N_331,In_685,In_426);
or U332 (N_332,In_44,N_186);
nand U333 (N_333,In_686,In_134);
nor U334 (N_334,In_96,In_565);
nor U335 (N_335,N_140,In_497);
nand U336 (N_336,In_84,N_61);
and U337 (N_337,In_329,In_477);
nor U338 (N_338,N_85,In_16);
and U339 (N_339,In_492,In_697);
or U340 (N_340,N_119,N_159);
nor U341 (N_341,In_657,N_187);
or U342 (N_342,N_191,In_462);
nand U343 (N_343,N_59,N_127);
or U344 (N_344,N_132,In_148);
and U345 (N_345,N_75,In_110);
and U346 (N_346,N_35,N_110);
and U347 (N_347,In_331,In_504);
nand U348 (N_348,In_525,N_83);
and U349 (N_349,In_182,In_404);
xor U350 (N_350,In_740,In_500);
or U351 (N_351,In_88,In_262);
nand U352 (N_352,N_48,N_125);
nand U353 (N_353,N_137,N_189);
nand U354 (N_354,N_26,In_423);
nand U355 (N_355,In_728,In_731);
or U356 (N_356,In_398,In_63);
and U357 (N_357,In_460,In_213);
nand U358 (N_358,In_284,In_42);
nand U359 (N_359,N_169,N_18);
nor U360 (N_360,In_267,In_185);
nand U361 (N_361,N_168,N_22);
xnor U362 (N_362,In_475,In_556);
xor U363 (N_363,In_653,In_521);
nor U364 (N_364,N_108,In_343);
or U365 (N_365,In_15,In_14);
and U366 (N_366,N_107,In_733);
and U367 (N_367,In_105,In_509);
and U368 (N_368,In_698,N_60);
and U369 (N_369,N_16,In_429);
nand U370 (N_370,N_130,In_299);
or U371 (N_371,In_510,N_188);
and U372 (N_372,In_479,N_68);
and U373 (N_373,N_73,In_51);
nor U374 (N_374,In_434,In_702);
nor U375 (N_375,In_321,In_36);
and U376 (N_376,N_175,N_126);
xnor U377 (N_377,In_80,N_79);
or U378 (N_378,N_34,N_113);
and U379 (N_379,In_638,N_196);
nand U380 (N_380,In_676,N_92);
nor U381 (N_381,In_442,N_197);
or U382 (N_382,In_725,N_78);
and U383 (N_383,In_688,In_33);
nand U384 (N_384,In_722,In_456);
nor U385 (N_385,In_719,In_210);
or U386 (N_386,N_5,In_12);
nand U387 (N_387,In_550,N_116);
nand U388 (N_388,N_95,In_260);
xnor U389 (N_389,N_55,In_495);
and U390 (N_390,N_72,N_37);
nand U391 (N_391,In_459,In_520);
nor U392 (N_392,In_683,In_107);
and U393 (N_393,In_483,N_36);
xor U394 (N_394,N_115,In_541);
nor U395 (N_395,N_117,N_58);
nand U396 (N_396,N_103,In_405);
xor U397 (N_397,N_84,In_303);
nor U398 (N_398,In_328,In_519);
or U399 (N_399,In_168,In_585);
nor U400 (N_400,N_170,In_527);
nor U401 (N_401,N_231,N_350);
nor U402 (N_402,N_277,N_269);
or U403 (N_403,N_287,In_116);
nand U404 (N_404,N_236,N_38);
and U405 (N_405,N_265,In_112);
nor U406 (N_406,N_238,N_100);
nor U407 (N_407,N_138,In_304);
nand U408 (N_408,In_183,N_49);
and U409 (N_409,N_232,In_593);
xor U410 (N_410,In_184,N_165);
and U411 (N_411,N_264,N_181);
nor U412 (N_412,N_227,N_157);
or U413 (N_413,N_27,N_339);
nor U414 (N_414,N_202,In_352);
nor U415 (N_415,In_575,In_239);
and U416 (N_416,N_272,N_267);
nor U417 (N_417,N_361,In_482);
nand U418 (N_418,In_219,In_250);
xnor U419 (N_419,N_389,N_305);
nand U420 (N_420,N_133,N_282);
nor U421 (N_421,In_159,N_289);
nand U422 (N_422,In_222,In_271);
nor U423 (N_423,N_256,N_141);
nand U424 (N_424,N_301,In_216);
and U425 (N_425,N_9,N_193);
nand U426 (N_426,N_155,N_281);
nor U427 (N_427,N_14,N_296);
xor U428 (N_428,N_241,N_106);
xnor U429 (N_429,N_134,N_373);
nor U430 (N_430,N_248,N_351);
and U431 (N_431,N_366,N_369);
and U432 (N_432,N_229,In_713);
and U433 (N_433,N_200,N_304);
or U434 (N_434,In_190,In_413);
or U435 (N_435,In_463,N_362);
or U436 (N_436,N_221,N_397);
nor U437 (N_437,N_328,N_162);
nand U438 (N_438,In_78,N_284);
and U439 (N_439,N_0,N_230);
or U440 (N_440,N_210,In_97);
and U441 (N_441,N_355,In_348);
or U442 (N_442,In_143,N_324);
nor U443 (N_443,N_317,N_99);
nor U444 (N_444,N_294,N_368);
and U445 (N_445,N_358,In_446);
or U446 (N_446,N_244,N_270);
xnor U447 (N_447,N_285,N_246);
nand U448 (N_448,N_390,N_247);
and U449 (N_449,N_380,N_52);
nand U450 (N_450,N_332,N_303);
and U451 (N_451,N_399,N_288);
and U452 (N_452,N_53,N_152);
or U453 (N_453,N_179,N_204);
and U454 (N_454,N_216,In_108);
nor U455 (N_455,N_331,N_70);
or U456 (N_456,N_314,N_81);
or U457 (N_457,In_563,N_245);
nor U458 (N_458,N_290,N_365);
or U459 (N_459,In_684,N_336);
nand U460 (N_460,In_614,N_131);
or U461 (N_461,N_279,N_249);
nand U462 (N_462,N_320,N_222);
and U463 (N_463,N_88,N_10);
and U464 (N_464,N_201,N_185);
nor U465 (N_465,N_171,N_310);
nand U466 (N_466,In_428,N_217);
or U467 (N_467,N_292,In_155);
nand U468 (N_468,N_302,N_370);
nand U469 (N_469,N_309,In_310);
nor U470 (N_470,In_19,N_359);
nor U471 (N_471,N_376,N_184);
and U472 (N_472,N_315,N_383);
or U473 (N_473,N_253,N_118);
nor U474 (N_474,In_253,N_271);
nand U475 (N_475,In_581,N_291);
nor U476 (N_476,N_298,N_391);
or U477 (N_477,N_352,N_307);
nand U478 (N_478,In_661,N_6);
nand U479 (N_479,In_27,N_224);
xnor U480 (N_480,N_276,In_402);
and U481 (N_481,N_308,N_39);
and U482 (N_482,In_615,N_325);
nor U483 (N_483,N_283,N_357);
or U484 (N_484,In_454,N_318);
xnor U485 (N_485,N_327,In_726);
xnor U486 (N_486,In_528,N_257);
and U487 (N_487,In_158,N_237);
nor U488 (N_488,N_158,In_102);
nand U489 (N_489,In_332,N_393);
and U490 (N_490,In_64,N_82);
nand U491 (N_491,N_396,N_394);
nor U492 (N_492,N_223,N_385);
and U493 (N_493,N_258,N_225);
or U494 (N_494,N_3,N_323);
and U495 (N_495,In_738,In_389);
nand U496 (N_496,N_382,N_395);
or U497 (N_497,N_199,N_345);
or U498 (N_498,N_326,N_316);
and U499 (N_499,N_56,In_741);
and U500 (N_500,In_160,In_377);
xor U501 (N_501,In_30,N_206);
or U502 (N_502,N_295,N_252);
and U503 (N_503,N_228,N_377);
nor U504 (N_504,N_340,N_163);
xor U505 (N_505,In_493,N_347);
nor U506 (N_506,N_242,N_299);
and U507 (N_507,N_205,N_226);
xor U508 (N_508,In_531,In_579);
xor U509 (N_509,N_208,N_263);
nor U510 (N_510,N_251,N_378);
and U511 (N_511,N_313,In_430);
or U512 (N_512,N_214,In_420);
xnor U513 (N_513,N_322,In_545);
or U514 (N_514,N_135,In_616);
nor U515 (N_515,N_330,N_334);
nand U516 (N_516,N_363,N_374);
or U517 (N_517,In_503,N_312);
nor U518 (N_518,N_346,N_342);
nor U519 (N_519,In_170,N_311);
xnor U520 (N_520,N_234,N_356);
nand U521 (N_521,N_275,In_34);
nand U522 (N_522,N_379,N_371);
or U523 (N_523,N_297,In_659);
and U524 (N_524,N_235,N_364);
nand U525 (N_525,N_212,In_21);
nand U526 (N_526,In_142,N_349);
or U527 (N_527,In_673,N_381);
nor U528 (N_528,In_162,N_286);
nand U529 (N_529,N_62,N_384);
nor U530 (N_530,N_333,In_496);
nand U531 (N_531,N_149,N_195);
and U532 (N_532,N_337,N_211);
nand U533 (N_533,N_343,N_259);
xor U534 (N_534,N_15,N_91);
nand U535 (N_535,N_280,In_660);
nor U536 (N_536,In_35,N_239);
or U537 (N_537,N_338,N_250);
nor U538 (N_538,N_335,In_55);
nand U539 (N_539,N_80,N_388);
or U540 (N_540,In_561,In_364);
or U541 (N_541,In_197,N_240);
nand U542 (N_542,In_355,N_348);
and U543 (N_543,N_367,N_306);
nor U544 (N_544,N_121,In_601);
or U545 (N_545,In_597,N_142);
nand U546 (N_546,N_154,In_187);
nand U547 (N_547,N_341,N_124);
nand U548 (N_548,In_675,In_704);
xnor U549 (N_549,In_647,N_255);
xor U550 (N_550,N_344,In_380);
nor U551 (N_551,N_43,N_207);
and U552 (N_552,N_213,N_266);
or U553 (N_553,N_273,N_392);
or U554 (N_554,In_307,N_375);
nand U555 (N_555,N_372,N_96);
nand U556 (N_556,N_254,In_292);
nand U557 (N_557,N_360,N_243);
xnor U558 (N_558,N_274,In_156);
or U559 (N_559,N_268,N_150);
nor U560 (N_560,N_220,N_209);
xor U561 (N_561,N_398,N_203);
nor U562 (N_562,N_45,In_508);
nand U563 (N_563,N_261,N_123);
or U564 (N_564,N_215,N_293);
nor U565 (N_565,N_262,In_259);
nand U566 (N_566,N_233,In_403);
and U567 (N_567,In_388,N_182);
xor U568 (N_568,N_278,N_353);
nor U569 (N_569,In_406,N_319);
and U570 (N_570,In_278,N_321);
nor U571 (N_571,N_218,N_386);
or U572 (N_572,N_300,N_219);
or U573 (N_573,N_260,N_387);
nor U574 (N_574,N_329,N_354);
or U575 (N_575,N_252,In_304);
nor U576 (N_576,N_371,N_99);
nand U577 (N_577,N_396,In_659);
nor U578 (N_578,N_329,In_307);
xnor U579 (N_579,N_390,N_208);
or U580 (N_580,N_9,N_15);
nor U581 (N_581,N_208,In_332);
xnor U582 (N_582,In_420,In_34);
nand U583 (N_583,In_675,N_287);
nor U584 (N_584,N_171,N_138);
nand U585 (N_585,N_277,In_143);
and U586 (N_586,N_346,N_154);
nor U587 (N_587,In_454,N_121);
nand U588 (N_588,In_713,N_296);
and U589 (N_589,N_135,N_358);
and U590 (N_590,N_121,N_96);
xnor U591 (N_591,N_313,N_391);
nor U592 (N_592,In_659,N_361);
or U593 (N_593,N_284,N_385);
or U594 (N_594,N_15,N_70);
or U595 (N_595,In_332,N_38);
nand U596 (N_596,N_300,N_389);
nand U597 (N_597,N_307,In_190);
nand U598 (N_598,N_226,N_39);
xor U599 (N_599,N_217,N_70);
nand U600 (N_600,N_468,N_471);
or U601 (N_601,N_569,N_497);
xnor U602 (N_602,N_402,N_546);
and U603 (N_603,N_582,N_484);
nand U604 (N_604,N_407,N_430);
nor U605 (N_605,N_577,N_405);
and U606 (N_606,N_505,N_429);
nand U607 (N_607,N_481,N_476);
and U608 (N_608,N_451,N_529);
nor U609 (N_609,N_444,N_564);
nor U610 (N_610,N_563,N_473);
nand U611 (N_611,N_499,N_493);
and U612 (N_612,N_470,N_524);
nand U613 (N_613,N_480,N_597);
nor U614 (N_614,N_513,N_442);
nand U615 (N_615,N_464,N_543);
nor U616 (N_616,N_446,N_447);
and U617 (N_617,N_594,N_580);
xnor U618 (N_618,N_579,N_590);
nor U619 (N_619,N_408,N_454);
nand U620 (N_620,N_581,N_552);
and U621 (N_621,N_475,N_437);
nor U622 (N_622,N_494,N_438);
nor U623 (N_623,N_414,N_586);
or U624 (N_624,N_521,N_401);
xnor U625 (N_625,N_489,N_547);
nor U626 (N_626,N_424,N_558);
and U627 (N_627,N_436,N_504);
nand U628 (N_628,N_526,N_434);
nand U629 (N_629,N_512,N_465);
and U630 (N_630,N_488,N_453);
nand U631 (N_631,N_435,N_461);
and U632 (N_632,N_531,N_587);
nand U633 (N_633,N_583,N_425);
nor U634 (N_634,N_472,N_517);
nor U635 (N_635,N_568,N_427);
nor U636 (N_636,N_432,N_518);
and U637 (N_637,N_422,N_466);
nand U638 (N_638,N_503,N_538);
xor U639 (N_639,N_522,N_441);
nand U640 (N_640,N_527,N_445);
nand U641 (N_641,N_485,N_553);
and U642 (N_642,N_539,N_423);
nand U643 (N_643,N_421,N_491);
and U644 (N_644,N_544,N_535);
xor U645 (N_645,N_428,N_506);
nand U646 (N_646,N_495,N_534);
nand U647 (N_647,N_567,N_431);
nand U648 (N_648,N_554,N_459);
nor U649 (N_649,N_456,N_508);
or U650 (N_650,N_572,N_448);
or U651 (N_651,N_565,N_440);
xnor U652 (N_652,N_460,N_509);
nand U653 (N_653,N_498,N_542);
or U654 (N_654,N_500,N_496);
nand U655 (N_655,N_528,N_467);
or U656 (N_656,N_479,N_541);
nor U657 (N_657,N_549,N_417);
xnor U658 (N_658,N_410,N_449);
and U659 (N_659,N_566,N_426);
or U660 (N_660,N_536,N_557);
nor U661 (N_661,N_501,N_584);
or U662 (N_662,N_462,N_502);
or U663 (N_663,N_574,N_575);
nor U664 (N_664,N_540,N_562);
nand U665 (N_665,N_477,N_550);
nand U666 (N_666,N_433,N_419);
xor U667 (N_667,N_515,N_571);
nand U668 (N_668,N_516,N_415);
nand U669 (N_669,N_457,N_537);
or U670 (N_670,N_598,N_450);
xor U671 (N_671,N_548,N_570);
or U672 (N_672,N_585,N_403);
nand U673 (N_673,N_591,N_592);
and U674 (N_674,N_555,N_593);
and U675 (N_675,N_439,N_523);
nand U676 (N_676,N_474,N_576);
or U677 (N_677,N_455,N_469);
or U678 (N_678,N_595,N_533);
and U679 (N_679,N_409,N_483);
nand U680 (N_680,N_482,N_404);
nand U681 (N_681,N_599,N_452);
nor U682 (N_682,N_463,N_406);
or U683 (N_683,N_458,N_507);
and U684 (N_684,N_532,N_400);
and U685 (N_685,N_588,N_411);
nor U686 (N_686,N_520,N_596);
or U687 (N_687,N_525,N_556);
nor U688 (N_688,N_416,N_514);
or U689 (N_689,N_559,N_412);
nor U690 (N_690,N_418,N_490);
and U691 (N_691,N_560,N_561);
and U692 (N_692,N_511,N_420);
or U693 (N_693,N_413,N_487);
nand U694 (N_694,N_486,N_492);
nand U695 (N_695,N_530,N_573);
or U696 (N_696,N_519,N_478);
nor U697 (N_697,N_510,N_551);
xnor U698 (N_698,N_589,N_578);
xnor U699 (N_699,N_443,N_545);
and U700 (N_700,N_424,N_582);
or U701 (N_701,N_402,N_522);
or U702 (N_702,N_522,N_512);
nor U703 (N_703,N_578,N_447);
nand U704 (N_704,N_563,N_487);
nor U705 (N_705,N_565,N_413);
or U706 (N_706,N_434,N_408);
and U707 (N_707,N_422,N_476);
nor U708 (N_708,N_430,N_534);
nand U709 (N_709,N_593,N_581);
nand U710 (N_710,N_583,N_406);
xor U711 (N_711,N_471,N_485);
nand U712 (N_712,N_487,N_431);
and U713 (N_713,N_592,N_547);
and U714 (N_714,N_452,N_511);
nor U715 (N_715,N_514,N_446);
nor U716 (N_716,N_485,N_517);
and U717 (N_717,N_449,N_525);
and U718 (N_718,N_452,N_460);
nor U719 (N_719,N_583,N_556);
or U720 (N_720,N_509,N_548);
nand U721 (N_721,N_504,N_564);
and U722 (N_722,N_454,N_442);
or U723 (N_723,N_417,N_447);
or U724 (N_724,N_433,N_475);
nor U725 (N_725,N_440,N_406);
xnor U726 (N_726,N_442,N_517);
nand U727 (N_727,N_492,N_590);
nand U728 (N_728,N_565,N_546);
and U729 (N_729,N_583,N_561);
and U730 (N_730,N_503,N_583);
xnor U731 (N_731,N_445,N_524);
nand U732 (N_732,N_480,N_491);
and U733 (N_733,N_444,N_591);
nand U734 (N_734,N_491,N_540);
nor U735 (N_735,N_493,N_473);
nand U736 (N_736,N_486,N_414);
or U737 (N_737,N_400,N_520);
or U738 (N_738,N_405,N_545);
xnor U739 (N_739,N_497,N_514);
xor U740 (N_740,N_468,N_432);
and U741 (N_741,N_469,N_556);
and U742 (N_742,N_484,N_546);
or U743 (N_743,N_508,N_553);
or U744 (N_744,N_501,N_474);
nor U745 (N_745,N_549,N_416);
or U746 (N_746,N_403,N_410);
xnor U747 (N_747,N_485,N_492);
and U748 (N_748,N_544,N_537);
nand U749 (N_749,N_514,N_418);
nor U750 (N_750,N_495,N_473);
xor U751 (N_751,N_465,N_548);
nand U752 (N_752,N_551,N_572);
nor U753 (N_753,N_454,N_494);
and U754 (N_754,N_446,N_569);
nand U755 (N_755,N_444,N_451);
nand U756 (N_756,N_533,N_559);
or U757 (N_757,N_583,N_569);
or U758 (N_758,N_563,N_474);
xor U759 (N_759,N_537,N_490);
xnor U760 (N_760,N_501,N_489);
nor U761 (N_761,N_519,N_412);
nor U762 (N_762,N_581,N_491);
xnor U763 (N_763,N_442,N_522);
or U764 (N_764,N_432,N_509);
and U765 (N_765,N_419,N_534);
and U766 (N_766,N_484,N_424);
nor U767 (N_767,N_432,N_496);
and U768 (N_768,N_556,N_566);
xor U769 (N_769,N_513,N_476);
or U770 (N_770,N_428,N_577);
or U771 (N_771,N_467,N_429);
and U772 (N_772,N_577,N_586);
nor U773 (N_773,N_578,N_527);
nor U774 (N_774,N_482,N_412);
nand U775 (N_775,N_455,N_539);
nor U776 (N_776,N_507,N_565);
or U777 (N_777,N_433,N_474);
xor U778 (N_778,N_536,N_459);
nor U779 (N_779,N_531,N_545);
or U780 (N_780,N_506,N_558);
nand U781 (N_781,N_410,N_557);
xnor U782 (N_782,N_471,N_575);
xor U783 (N_783,N_525,N_437);
xor U784 (N_784,N_430,N_449);
nand U785 (N_785,N_514,N_456);
nor U786 (N_786,N_513,N_552);
nor U787 (N_787,N_476,N_503);
xnor U788 (N_788,N_423,N_493);
nand U789 (N_789,N_401,N_488);
and U790 (N_790,N_521,N_551);
and U791 (N_791,N_443,N_527);
or U792 (N_792,N_511,N_462);
or U793 (N_793,N_458,N_540);
and U794 (N_794,N_404,N_524);
xnor U795 (N_795,N_563,N_564);
or U796 (N_796,N_409,N_587);
and U797 (N_797,N_586,N_556);
and U798 (N_798,N_556,N_567);
nand U799 (N_799,N_597,N_591);
nor U800 (N_800,N_611,N_694);
nand U801 (N_801,N_794,N_702);
nand U802 (N_802,N_766,N_604);
or U803 (N_803,N_771,N_684);
and U804 (N_804,N_600,N_745);
nand U805 (N_805,N_797,N_648);
xnor U806 (N_806,N_635,N_751);
or U807 (N_807,N_731,N_720);
and U808 (N_808,N_748,N_718);
nor U809 (N_809,N_746,N_735);
nor U810 (N_810,N_743,N_703);
nand U811 (N_811,N_693,N_753);
and U812 (N_812,N_659,N_668);
nand U813 (N_813,N_613,N_630);
and U814 (N_814,N_642,N_717);
or U815 (N_815,N_618,N_780);
and U816 (N_816,N_793,N_632);
nor U817 (N_817,N_733,N_616);
nor U818 (N_818,N_678,N_624);
nor U819 (N_819,N_602,N_614);
xor U820 (N_820,N_747,N_656);
or U821 (N_821,N_760,N_645);
and U822 (N_822,N_629,N_625);
nand U823 (N_823,N_687,N_701);
nor U824 (N_824,N_615,N_640);
xor U825 (N_825,N_691,N_665);
nor U826 (N_826,N_727,N_763);
nand U827 (N_827,N_709,N_700);
nor U828 (N_828,N_790,N_627);
and U829 (N_829,N_698,N_667);
xnor U830 (N_830,N_696,N_758);
nor U831 (N_831,N_712,N_690);
nand U832 (N_832,N_719,N_734);
or U833 (N_833,N_791,N_744);
nand U834 (N_834,N_786,N_750);
nor U835 (N_835,N_787,N_776);
or U836 (N_836,N_646,N_664);
and U837 (N_837,N_673,N_626);
nand U838 (N_838,N_738,N_666);
nor U839 (N_839,N_644,N_796);
or U840 (N_840,N_772,N_730);
nand U841 (N_841,N_637,N_603);
nor U842 (N_842,N_674,N_695);
and U843 (N_843,N_728,N_605);
nor U844 (N_844,N_610,N_788);
nor U845 (N_845,N_639,N_708);
and U846 (N_846,N_774,N_707);
or U847 (N_847,N_762,N_683);
and U848 (N_848,N_619,N_757);
nor U849 (N_849,N_620,N_677);
nor U850 (N_850,N_737,N_653);
xor U851 (N_851,N_652,N_699);
xor U852 (N_852,N_617,N_785);
nand U853 (N_853,N_658,N_792);
and U854 (N_854,N_641,N_779);
or U855 (N_855,N_675,N_752);
nor U856 (N_856,N_732,N_676);
or U857 (N_857,N_713,N_756);
or U858 (N_858,N_606,N_633);
or U859 (N_859,N_649,N_775);
and U860 (N_860,N_672,N_657);
nand U861 (N_861,N_777,N_782);
or U862 (N_862,N_685,N_716);
or U863 (N_863,N_773,N_679);
and U864 (N_864,N_768,N_755);
nand U865 (N_865,N_722,N_634);
or U866 (N_866,N_705,N_706);
nor U867 (N_867,N_724,N_628);
and U868 (N_868,N_654,N_741);
or U869 (N_869,N_669,N_798);
nor U870 (N_870,N_608,N_789);
or U871 (N_871,N_650,N_764);
nand U872 (N_872,N_686,N_609);
nor U873 (N_873,N_670,N_710);
or U874 (N_874,N_697,N_795);
nor U875 (N_875,N_740,N_621);
nor U876 (N_876,N_799,N_759);
and U877 (N_877,N_784,N_754);
nor U878 (N_878,N_761,N_682);
nor U879 (N_879,N_715,N_636);
or U880 (N_880,N_729,N_783);
xor U881 (N_881,N_736,N_623);
nor U882 (N_882,N_767,N_688);
nor U883 (N_883,N_631,N_781);
nor U884 (N_884,N_726,N_770);
nor U885 (N_885,N_663,N_704);
and U886 (N_886,N_638,N_661);
and U887 (N_887,N_739,N_671);
nand U888 (N_888,N_660,N_643);
or U889 (N_889,N_680,N_769);
nor U890 (N_890,N_607,N_622);
and U891 (N_891,N_749,N_692);
nor U892 (N_892,N_714,N_778);
xnor U893 (N_893,N_742,N_647);
or U894 (N_894,N_711,N_655);
nor U895 (N_895,N_601,N_765);
or U896 (N_896,N_725,N_651);
nand U897 (N_897,N_662,N_689);
nor U898 (N_898,N_612,N_681);
nor U899 (N_899,N_723,N_721);
nand U900 (N_900,N_691,N_655);
and U901 (N_901,N_774,N_713);
or U902 (N_902,N_602,N_651);
or U903 (N_903,N_664,N_644);
nor U904 (N_904,N_761,N_608);
xnor U905 (N_905,N_617,N_760);
and U906 (N_906,N_603,N_602);
and U907 (N_907,N_630,N_794);
or U908 (N_908,N_671,N_683);
and U909 (N_909,N_694,N_721);
or U910 (N_910,N_633,N_794);
or U911 (N_911,N_645,N_673);
xor U912 (N_912,N_767,N_709);
and U913 (N_913,N_711,N_729);
nand U914 (N_914,N_771,N_672);
nand U915 (N_915,N_715,N_708);
or U916 (N_916,N_602,N_623);
or U917 (N_917,N_699,N_613);
nand U918 (N_918,N_657,N_728);
nor U919 (N_919,N_615,N_614);
nor U920 (N_920,N_684,N_680);
xor U921 (N_921,N_682,N_668);
nand U922 (N_922,N_648,N_732);
or U923 (N_923,N_707,N_797);
and U924 (N_924,N_779,N_742);
nor U925 (N_925,N_630,N_791);
nand U926 (N_926,N_741,N_636);
nor U927 (N_927,N_687,N_620);
nand U928 (N_928,N_669,N_760);
and U929 (N_929,N_617,N_601);
nand U930 (N_930,N_631,N_611);
and U931 (N_931,N_777,N_652);
or U932 (N_932,N_703,N_694);
or U933 (N_933,N_774,N_749);
nor U934 (N_934,N_724,N_657);
nor U935 (N_935,N_737,N_788);
or U936 (N_936,N_640,N_778);
nand U937 (N_937,N_720,N_773);
or U938 (N_938,N_782,N_609);
and U939 (N_939,N_718,N_770);
nand U940 (N_940,N_703,N_620);
nor U941 (N_941,N_684,N_667);
nand U942 (N_942,N_690,N_683);
or U943 (N_943,N_736,N_633);
and U944 (N_944,N_656,N_658);
nand U945 (N_945,N_720,N_793);
and U946 (N_946,N_795,N_691);
nor U947 (N_947,N_675,N_715);
nand U948 (N_948,N_659,N_749);
nand U949 (N_949,N_785,N_699);
nand U950 (N_950,N_743,N_612);
or U951 (N_951,N_644,N_646);
nand U952 (N_952,N_627,N_678);
nand U953 (N_953,N_751,N_626);
or U954 (N_954,N_658,N_682);
and U955 (N_955,N_720,N_659);
nand U956 (N_956,N_747,N_743);
and U957 (N_957,N_643,N_622);
and U958 (N_958,N_712,N_797);
and U959 (N_959,N_661,N_697);
or U960 (N_960,N_729,N_657);
nor U961 (N_961,N_789,N_778);
xor U962 (N_962,N_661,N_682);
and U963 (N_963,N_735,N_612);
nand U964 (N_964,N_741,N_730);
or U965 (N_965,N_607,N_731);
or U966 (N_966,N_623,N_605);
and U967 (N_967,N_671,N_686);
and U968 (N_968,N_725,N_697);
xor U969 (N_969,N_718,N_699);
and U970 (N_970,N_739,N_632);
nor U971 (N_971,N_666,N_730);
nor U972 (N_972,N_640,N_774);
xnor U973 (N_973,N_732,N_649);
nor U974 (N_974,N_791,N_618);
nor U975 (N_975,N_689,N_747);
xnor U976 (N_976,N_619,N_686);
nor U977 (N_977,N_636,N_776);
or U978 (N_978,N_663,N_722);
or U979 (N_979,N_696,N_630);
nor U980 (N_980,N_760,N_611);
nand U981 (N_981,N_603,N_620);
and U982 (N_982,N_706,N_730);
or U983 (N_983,N_751,N_738);
nand U984 (N_984,N_742,N_663);
nor U985 (N_985,N_797,N_695);
nand U986 (N_986,N_683,N_720);
or U987 (N_987,N_780,N_708);
and U988 (N_988,N_624,N_760);
and U989 (N_989,N_694,N_786);
or U990 (N_990,N_616,N_776);
nand U991 (N_991,N_774,N_751);
nand U992 (N_992,N_647,N_681);
nand U993 (N_993,N_743,N_653);
nand U994 (N_994,N_789,N_618);
nand U995 (N_995,N_791,N_687);
and U996 (N_996,N_784,N_785);
nand U997 (N_997,N_663,N_640);
and U998 (N_998,N_733,N_710);
nor U999 (N_999,N_704,N_646);
or U1000 (N_1000,N_848,N_997);
nor U1001 (N_1001,N_937,N_901);
nor U1002 (N_1002,N_841,N_895);
nand U1003 (N_1003,N_993,N_900);
and U1004 (N_1004,N_885,N_941);
and U1005 (N_1005,N_827,N_852);
nand U1006 (N_1006,N_909,N_850);
xor U1007 (N_1007,N_843,N_920);
and U1008 (N_1008,N_971,N_931);
nand U1009 (N_1009,N_950,N_991);
nor U1010 (N_1010,N_805,N_803);
and U1011 (N_1011,N_954,N_844);
or U1012 (N_1012,N_932,N_964);
or U1013 (N_1013,N_983,N_921);
and U1014 (N_1014,N_908,N_888);
or U1015 (N_1015,N_966,N_936);
nor U1016 (N_1016,N_818,N_802);
xnor U1017 (N_1017,N_899,N_872);
nand U1018 (N_1018,N_861,N_834);
or U1019 (N_1019,N_855,N_912);
or U1020 (N_1020,N_978,N_825);
nand U1021 (N_1021,N_836,N_924);
or U1022 (N_1022,N_985,N_892);
nand U1023 (N_1023,N_819,N_878);
nand U1024 (N_1024,N_907,N_846);
and U1025 (N_1025,N_961,N_915);
nor U1026 (N_1026,N_994,N_972);
nand U1027 (N_1027,N_820,N_982);
or U1028 (N_1028,N_979,N_829);
nand U1029 (N_1029,N_943,N_989);
nor U1030 (N_1030,N_815,N_823);
nand U1031 (N_1031,N_864,N_999);
and U1032 (N_1032,N_877,N_956);
nor U1033 (N_1033,N_927,N_988);
nand U1034 (N_1034,N_976,N_811);
nor U1035 (N_1035,N_859,N_830);
nand U1036 (N_1036,N_889,N_824);
nand U1037 (N_1037,N_886,N_874);
xnor U1038 (N_1038,N_948,N_856);
nor U1039 (N_1039,N_832,N_807);
and U1040 (N_1040,N_902,N_887);
and U1041 (N_1041,N_868,N_928);
and U1042 (N_1042,N_817,N_967);
nand U1043 (N_1043,N_810,N_970);
nor U1044 (N_1044,N_934,N_821);
or U1045 (N_1045,N_858,N_867);
or U1046 (N_1046,N_980,N_905);
and U1047 (N_1047,N_857,N_891);
and U1048 (N_1048,N_959,N_847);
nor U1049 (N_1049,N_840,N_945);
nand U1050 (N_1050,N_849,N_952);
nand U1051 (N_1051,N_863,N_801);
or U1052 (N_1052,N_914,N_873);
or U1053 (N_1053,N_963,N_944);
and U1054 (N_1054,N_884,N_879);
nor U1055 (N_1055,N_860,N_837);
or U1056 (N_1056,N_939,N_923);
nor U1057 (N_1057,N_975,N_922);
nor U1058 (N_1058,N_953,N_929);
or U1059 (N_1059,N_942,N_808);
nor U1060 (N_1060,N_933,N_987);
xnor U1061 (N_1061,N_965,N_813);
and U1062 (N_1062,N_947,N_842);
and U1063 (N_1063,N_853,N_903);
nor U1064 (N_1064,N_940,N_804);
xnor U1065 (N_1065,N_870,N_938);
nand U1066 (N_1066,N_866,N_816);
nor U1067 (N_1067,N_962,N_833);
nand U1068 (N_1068,N_916,N_995);
nand U1069 (N_1069,N_919,N_973);
and U1070 (N_1070,N_875,N_838);
and U1071 (N_1071,N_960,N_935);
nand U1072 (N_1072,N_930,N_896);
and U1073 (N_1073,N_809,N_835);
xor U1074 (N_1074,N_906,N_998);
and U1075 (N_1075,N_862,N_992);
or U1076 (N_1076,N_969,N_831);
nand U1077 (N_1077,N_865,N_883);
xnor U1078 (N_1078,N_996,N_845);
or U1079 (N_1079,N_926,N_910);
or U1080 (N_1080,N_917,N_957);
nand U1081 (N_1081,N_977,N_918);
nor U1082 (N_1082,N_814,N_881);
or U1083 (N_1083,N_981,N_949);
nand U1084 (N_1084,N_913,N_876);
or U1085 (N_1085,N_826,N_822);
and U1086 (N_1086,N_951,N_968);
or U1087 (N_1087,N_974,N_904);
nor U1088 (N_1088,N_894,N_946);
xnor U1089 (N_1089,N_871,N_806);
or U1090 (N_1090,N_925,N_893);
xnor U1091 (N_1091,N_880,N_986);
nor U1092 (N_1092,N_898,N_955);
and U1093 (N_1093,N_839,N_984);
and U1094 (N_1094,N_990,N_812);
and U1095 (N_1095,N_897,N_958);
and U1096 (N_1096,N_890,N_828);
nor U1097 (N_1097,N_869,N_911);
and U1098 (N_1098,N_854,N_851);
or U1099 (N_1099,N_882,N_800);
nand U1100 (N_1100,N_876,N_817);
nor U1101 (N_1101,N_814,N_964);
xnor U1102 (N_1102,N_987,N_926);
and U1103 (N_1103,N_907,N_994);
or U1104 (N_1104,N_857,N_916);
nand U1105 (N_1105,N_800,N_817);
nand U1106 (N_1106,N_900,N_920);
and U1107 (N_1107,N_997,N_953);
nor U1108 (N_1108,N_827,N_874);
nand U1109 (N_1109,N_927,N_844);
and U1110 (N_1110,N_892,N_845);
xor U1111 (N_1111,N_933,N_873);
or U1112 (N_1112,N_897,N_937);
nand U1113 (N_1113,N_888,N_830);
or U1114 (N_1114,N_869,N_985);
and U1115 (N_1115,N_980,N_919);
nand U1116 (N_1116,N_973,N_905);
xor U1117 (N_1117,N_818,N_898);
or U1118 (N_1118,N_824,N_899);
and U1119 (N_1119,N_884,N_849);
and U1120 (N_1120,N_935,N_823);
xor U1121 (N_1121,N_932,N_999);
nand U1122 (N_1122,N_854,N_889);
or U1123 (N_1123,N_971,N_984);
nor U1124 (N_1124,N_834,N_803);
nand U1125 (N_1125,N_845,N_847);
nand U1126 (N_1126,N_980,N_909);
nand U1127 (N_1127,N_895,N_868);
or U1128 (N_1128,N_969,N_912);
or U1129 (N_1129,N_942,N_921);
or U1130 (N_1130,N_807,N_960);
or U1131 (N_1131,N_858,N_856);
nand U1132 (N_1132,N_957,N_808);
or U1133 (N_1133,N_941,N_884);
or U1134 (N_1134,N_827,N_887);
and U1135 (N_1135,N_874,N_877);
or U1136 (N_1136,N_907,N_826);
and U1137 (N_1137,N_854,N_875);
nor U1138 (N_1138,N_942,N_805);
nor U1139 (N_1139,N_926,N_886);
xnor U1140 (N_1140,N_860,N_852);
or U1141 (N_1141,N_878,N_836);
nand U1142 (N_1142,N_941,N_845);
or U1143 (N_1143,N_968,N_845);
and U1144 (N_1144,N_947,N_821);
xor U1145 (N_1145,N_916,N_913);
xor U1146 (N_1146,N_817,N_838);
nand U1147 (N_1147,N_982,N_992);
xor U1148 (N_1148,N_870,N_871);
or U1149 (N_1149,N_810,N_849);
and U1150 (N_1150,N_932,N_865);
nand U1151 (N_1151,N_945,N_842);
or U1152 (N_1152,N_914,N_931);
nand U1153 (N_1153,N_930,N_853);
and U1154 (N_1154,N_812,N_971);
nand U1155 (N_1155,N_814,N_808);
or U1156 (N_1156,N_905,N_916);
or U1157 (N_1157,N_821,N_905);
nand U1158 (N_1158,N_965,N_930);
xnor U1159 (N_1159,N_951,N_938);
nand U1160 (N_1160,N_839,N_845);
nand U1161 (N_1161,N_929,N_942);
nor U1162 (N_1162,N_973,N_944);
and U1163 (N_1163,N_814,N_825);
xnor U1164 (N_1164,N_967,N_955);
nand U1165 (N_1165,N_946,N_826);
or U1166 (N_1166,N_992,N_879);
nor U1167 (N_1167,N_862,N_902);
or U1168 (N_1168,N_979,N_902);
nand U1169 (N_1169,N_873,N_863);
xnor U1170 (N_1170,N_985,N_999);
nor U1171 (N_1171,N_873,N_862);
and U1172 (N_1172,N_843,N_881);
and U1173 (N_1173,N_870,N_809);
or U1174 (N_1174,N_846,N_822);
and U1175 (N_1175,N_824,N_930);
nor U1176 (N_1176,N_886,N_879);
nand U1177 (N_1177,N_949,N_845);
nand U1178 (N_1178,N_933,N_947);
xor U1179 (N_1179,N_871,N_895);
nor U1180 (N_1180,N_964,N_963);
nor U1181 (N_1181,N_984,N_832);
or U1182 (N_1182,N_930,N_820);
nand U1183 (N_1183,N_970,N_879);
or U1184 (N_1184,N_874,N_851);
nand U1185 (N_1185,N_998,N_977);
nor U1186 (N_1186,N_995,N_918);
or U1187 (N_1187,N_853,N_890);
or U1188 (N_1188,N_868,N_894);
and U1189 (N_1189,N_934,N_901);
nand U1190 (N_1190,N_934,N_816);
and U1191 (N_1191,N_925,N_869);
and U1192 (N_1192,N_895,N_970);
nand U1193 (N_1193,N_861,N_979);
xor U1194 (N_1194,N_862,N_878);
nor U1195 (N_1195,N_930,N_848);
and U1196 (N_1196,N_999,N_899);
nor U1197 (N_1197,N_986,N_815);
and U1198 (N_1198,N_933,N_918);
nor U1199 (N_1199,N_953,N_962);
or U1200 (N_1200,N_1042,N_1009);
or U1201 (N_1201,N_1121,N_1017);
nor U1202 (N_1202,N_1118,N_1189);
nand U1203 (N_1203,N_1123,N_1081);
nand U1204 (N_1204,N_1111,N_1178);
and U1205 (N_1205,N_1059,N_1045);
nand U1206 (N_1206,N_1099,N_1164);
and U1207 (N_1207,N_1133,N_1030);
xor U1208 (N_1208,N_1135,N_1144);
and U1209 (N_1209,N_1061,N_1028);
nor U1210 (N_1210,N_1103,N_1003);
or U1211 (N_1211,N_1177,N_1181);
and U1212 (N_1212,N_1152,N_1086);
or U1213 (N_1213,N_1070,N_1127);
and U1214 (N_1214,N_1018,N_1014);
and U1215 (N_1215,N_1026,N_1155);
nand U1216 (N_1216,N_1115,N_1038);
nor U1217 (N_1217,N_1027,N_1004);
and U1218 (N_1218,N_1168,N_1142);
and U1219 (N_1219,N_1074,N_1107);
or U1220 (N_1220,N_1058,N_1062);
and U1221 (N_1221,N_1194,N_1160);
or U1222 (N_1222,N_1049,N_1110);
or U1223 (N_1223,N_1101,N_1015);
or U1224 (N_1224,N_1088,N_1041);
nand U1225 (N_1225,N_1102,N_1165);
and U1226 (N_1226,N_1093,N_1040);
nand U1227 (N_1227,N_1117,N_1192);
and U1228 (N_1228,N_1098,N_1173);
nor U1229 (N_1229,N_1166,N_1188);
xor U1230 (N_1230,N_1193,N_1186);
xor U1231 (N_1231,N_1159,N_1037);
nor U1232 (N_1232,N_1172,N_1196);
and U1233 (N_1233,N_1079,N_1089);
nand U1234 (N_1234,N_1151,N_1000);
or U1235 (N_1235,N_1112,N_1180);
nor U1236 (N_1236,N_1091,N_1134);
or U1237 (N_1237,N_1119,N_1199);
nand U1238 (N_1238,N_1161,N_1002);
nand U1239 (N_1239,N_1106,N_1136);
and U1240 (N_1240,N_1043,N_1185);
nor U1241 (N_1241,N_1031,N_1109);
and U1242 (N_1242,N_1016,N_1174);
nor U1243 (N_1243,N_1184,N_1073);
or U1244 (N_1244,N_1021,N_1146);
nand U1245 (N_1245,N_1092,N_1060);
and U1246 (N_1246,N_1063,N_1046);
and U1247 (N_1247,N_1154,N_1039);
nor U1248 (N_1248,N_1057,N_1066);
or U1249 (N_1249,N_1150,N_1048);
or U1250 (N_1250,N_1095,N_1055);
nand U1251 (N_1251,N_1100,N_1076);
nand U1252 (N_1252,N_1024,N_1094);
nand U1253 (N_1253,N_1114,N_1011);
nand U1254 (N_1254,N_1108,N_1120);
and U1255 (N_1255,N_1047,N_1010);
or U1256 (N_1256,N_1087,N_1001);
nor U1257 (N_1257,N_1141,N_1113);
nand U1258 (N_1258,N_1068,N_1147);
nor U1259 (N_1259,N_1128,N_1122);
nand U1260 (N_1260,N_1025,N_1191);
nor U1261 (N_1261,N_1158,N_1163);
nor U1262 (N_1262,N_1175,N_1105);
nand U1263 (N_1263,N_1097,N_1006);
or U1264 (N_1264,N_1149,N_1138);
nand U1265 (N_1265,N_1032,N_1036);
or U1266 (N_1266,N_1082,N_1080);
nand U1267 (N_1267,N_1183,N_1019);
and U1268 (N_1268,N_1020,N_1145);
or U1269 (N_1269,N_1033,N_1069);
nor U1270 (N_1270,N_1129,N_1085);
nor U1271 (N_1271,N_1169,N_1077);
nor U1272 (N_1272,N_1052,N_1187);
and U1273 (N_1273,N_1007,N_1124);
or U1274 (N_1274,N_1053,N_1198);
nor U1275 (N_1275,N_1195,N_1131);
nand U1276 (N_1276,N_1075,N_1176);
or U1277 (N_1277,N_1179,N_1035);
nor U1278 (N_1278,N_1054,N_1072);
xnor U1279 (N_1279,N_1125,N_1023);
nor U1280 (N_1280,N_1140,N_1167);
nand U1281 (N_1281,N_1005,N_1170);
nand U1282 (N_1282,N_1050,N_1156);
or U1283 (N_1283,N_1116,N_1126);
or U1284 (N_1284,N_1153,N_1143);
xor U1285 (N_1285,N_1190,N_1130);
nand U1286 (N_1286,N_1051,N_1182);
or U1287 (N_1287,N_1139,N_1148);
nor U1288 (N_1288,N_1197,N_1071);
or U1289 (N_1289,N_1078,N_1132);
nand U1290 (N_1290,N_1029,N_1067);
nand U1291 (N_1291,N_1162,N_1022);
nand U1292 (N_1292,N_1084,N_1044);
xnor U1293 (N_1293,N_1064,N_1137);
and U1294 (N_1294,N_1083,N_1096);
nand U1295 (N_1295,N_1012,N_1104);
xnor U1296 (N_1296,N_1013,N_1090);
or U1297 (N_1297,N_1034,N_1171);
xor U1298 (N_1298,N_1157,N_1056);
or U1299 (N_1299,N_1008,N_1065);
or U1300 (N_1300,N_1158,N_1064);
and U1301 (N_1301,N_1163,N_1198);
or U1302 (N_1302,N_1193,N_1150);
or U1303 (N_1303,N_1076,N_1111);
nand U1304 (N_1304,N_1011,N_1048);
or U1305 (N_1305,N_1019,N_1091);
and U1306 (N_1306,N_1102,N_1156);
xor U1307 (N_1307,N_1051,N_1116);
or U1308 (N_1308,N_1018,N_1019);
or U1309 (N_1309,N_1154,N_1051);
or U1310 (N_1310,N_1035,N_1138);
nand U1311 (N_1311,N_1016,N_1149);
nand U1312 (N_1312,N_1022,N_1130);
and U1313 (N_1313,N_1096,N_1177);
nand U1314 (N_1314,N_1016,N_1064);
or U1315 (N_1315,N_1088,N_1179);
nand U1316 (N_1316,N_1157,N_1007);
nand U1317 (N_1317,N_1190,N_1168);
and U1318 (N_1318,N_1004,N_1015);
or U1319 (N_1319,N_1084,N_1188);
or U1320 (N_1320,N_1082,N_1009);
nand U1321 (N_1321,N_1175,N_1148);
and U1322 (N_1322,N_1078,N_1099);
and U1323 (N_1323,N_1181,N_1194);
nand U1324 (N_1324,N_1188,N_1004);
and U1325 (N_1325,N_1084,N_1077);
xor U1326 (N_1326,N_1136,N_1168);
or U1327 (N_1327,N_1038,N_1001);
nor U1328 (N_1328,N_1107,N_1062);
nand U1329 (N_1329,N_1001,N_1134);
nand U1330 (N_1330,N_1155,N_1183);
and U1331 (N_1331,N_1097,N_1042);
xor U1332 (N_1332,N_1031,N_1171);
xnor U1333 (N_1333,N_1022,N_1031);
xnor U1334 (N_1334,N_1122,N_1022);
nor U1335 (N_1335,N_1067,N_1186);
or U1336 (N_1336,N_1183,N_1149);
and U1337 (N_1337,N_1166,N_1081);
nor U1338 (N_1338,N_1188,N_1100);
and U1339 (N_1339,N_1131,N_1017);
nor U1340 (N_1340,N_1067,N_1080);
nand U1341 (N_1341,N_1143,N_1075);
or U1342 (N_1342,N_1150,N_1176);
nand U1343 (N_1343,N_1048,N_1028);
or U1344 (N_1344,N_1030,N_1169);
nand U1345 (N_1345,N_1072,N_1001);
or U1346 (N_1346,N_1004,N_1071);
nand U1347 (N_1347,N_1032,N_1021);
or U1348 (N_1348,N_1098,N_1184);
nor U1349 (N_1349,N_1095,N_1066);
nor U1350 (N_1350,N_1012,N_1009);
or U1351 (N_1351,N_1152,N_1008);
and U1352 (N_1352,N_1003,N_1162);
or U1353 (N_1353,N_1163,N_1039);
or U1354 (N_1354,N_1054,N_1124);
nor U1355 (N_1355,N_1193,N_1016);
and U1356 (N_1356,N_1123,N_1131);
xor U1357 (N_1357,N_1155,N_1192);
or U1358 (N_1358,N_1186,N_1155);
and U1359 (N_1359,N_1031,N_1137);
nand U1360 (N_1360,N_1136,N_1130);
nand U1361 (N_1361,N_1056,N_1188);
nand U1362 (N_1362,N_1090,N_1132);
nor U1363 (N_1363,N_1112,N_1163);
nand U1364 (N_1364,N_1041,N_1199);
nand U1365 (N_1365,N_1123,N_1021);
xor U1366 (N_1366,N_1098,N_1034);
nor U1367 (N_1367,N_1051,N_1181);
nor U1368 (N_1368,N_1177,N_1193);
xor U1369 (N_1369,N_1155,N_1128);
nand U1370 (N_1370,N_1137,N_1075);
or U1371 (N_1371,N_1127,N_1069);
xor U1372 (N_1372,N_1001,N_1115);
nand U1373 (N_1373,N_1030,N_1182);
nand U1374 (N_1374,N_1028,N_1164);
or U1375 (N_1375,N_1108,N_1110);
nand U1376 (N_1376,N_1144,N_1049);
nand U1377 (N_1377,N_1123,N_1020);
xnor U1378 (N_1378,N_1189,N_1072);
nor U1379 (N_1379,N_1098,N_1099);
nand U1380 (N_1380,N_1043,N_1010);
or U1381 (N_1381,N_1008,N_1088);
nor U1382 (N_1382,N_1054,N_1185);
nand U1383 (N_1383,N_1103,N_1184);
or U1384 (N_1384,N_1192,N_1007);
nor U1385 (N_1385,N_1002,N_1005);
xor U1386 (N_1386,N_1006,N_1058);
nor U1387 (N_1387,N_1027,N_1191);
nand U1388 (N_1388,N_1084,N_1194);
nor U1389 (N_1389,N_1196,N_1029);
or U1390 (N_1390,N_1146,N_1077);
or U1391 (N_1391,N_1174,N_1081);
xnor U1392 (N_1392,N_1063,N_1015);
xor U1393 (N_1393,N_1092,N_1155);
xnor U1394 (N_1394,N_1108,N_1136);
or U1395 (N_1395,N_1034,N_1176);
nor U1396 (N_1396,N_1054,N_1078);
or U1397 (N_1397,N_1050,N_1190);
nor U1398 (N_1398,N_1101,N_1130);
and U1399 (N_1399,N_1181,N_1144);
or U1400 (N_1400,N_1377,N_1351);
and U1401 (N_1401,N_1236,N_1234);
nand U1402 (N_1402,N_1251,N_1244);
nor U1403 (N_1403,N_1393,N_1291);
nand U1404 (N_1404,N_1289,N_1370);
or U1405 (N_1405,N_1306,N_1305);
nor U1406 (N_1406,N_1241,N_1208);
or U1407 (N_1407,N_1249,N_1223);
nand U1408 (N_1408,N_1221,N_1255);
nor U1409 (N_1409,N_1358,N_1250);
or U1410 (N_1410,N_1385,N_1350);
and U1411 (N_1411,N_1212,N_1389);
nor U1412 (N_1412,N_1254,N_1313);
and U1413 (N_1413,N_1209,N_1292);
or U1414 (N_1414,N_1380,N_1323);
xor U1415 (N_1415,N_1359,N_1378);
nor U1416 (N_1416,N_1237,N_1398);
nor U1417 (N_1417,N_1344,N_1246);
and U1418 (N_1418,N_1384,N_1222);
nand U1419 (N_1419,N_1205,N_1258);
nor U1420 (N_1420,N_1207,N_1239);
xor U1421 (N_1421,N_1286,N_1215);
and U1422 (N_1422,N_1318,N_1211);
nand U1423 (N_1423,N_1352,N_1218);
and U1424 (N_1424,N_1354,N_1269);
nor U1425 (N_1425,N_1247,N_1217);
and U1426 (N_1426,N_1268,N_1348);
and U1427 (N_1427,N_1279,N_1369);
and U1428 (N_1428,N_1364,N_1259);
nand U1429 (N_1429,N_1395,N_1240);
nor U1430 (N_1430,N_1264,N_1252);
nor U1431 (N_1431,N_1256,N_1204);
nor U1432 (N_1432,N_1388,N_1299);
or U1433 (N_1433,N_1396,N_1266);
or U1434 (N_1434,N_1274,N_1338);
nand U1435 (N_1435,N_1276,N_1282);
xnor U1436 (N_1436,N_1257,N_1281);
nor U1437 (N_1437,N_1213,N_1301);
and U1438 (N_1438,N_1203,N_1300);
or U1439 (N_1439,N_1342,N_1332);
or U1440 (N_1440,N_1248,N_1227);
xor U1441 (N_1441,N_1297,N_1226);
nor U1442 (N_1442,N_1275,N_1220);
or U1443 (N_1443,N_1278,N_1345);
nor U1444 (N_1444,N_1312,N_1283);
nand U1445 (N_1445,N_1304,N_1273);
or U1446 (N_1446,N_1331,N_1375);
and U1447 (N_1447,N_1347,N_1231);
nand U1448 (N_1448,N_1309,N_1386);
nand U1449 (N_1449,N_1322,N_1319);
nand U1450 (N_1450,N_1262,N_1310);
nand U1451 (N_1451,N_1206,N_1360);
or U1452 (N_1452,N_1381,N_1260);
and U1453 (N_1453,N_1383,N_1397);
or U1454 (N_1454,N_1263,N_1242);
nand U1455 (N_1455,N_1390,N_1355);
or U1456 (N_1456,N_1376,N_1214);
nand U1457 (N_1457,N_1339,N_1361);
nand U1458 (N_1458,N_1210,N_1392);
nand U1459 (N_1459,N_1363,N_1349);
nor U1460 (N_1460,N_1325,N_1224);
nor U1461 (N_1461,N_1368,N_1357);
and U1462 (N_1462,N_1235,N_1294);
nand U1463 (N_1463,N_1394,N_1399);
or U1464 (N_1464,N_1253,N_1317);
and U1465 (N_1465,N_1298,N_1307);
xnor U1466 (N_1466,N_1277,N_1225);
xor U1467 (N_1467,N_1216,N_1233);
or U1468 (N_1468,N_1295,N_1232);
or U1469 (N_1469,N_1371,N_1314);
nand U1470 (N_1470,N_1328,N_1296);
and U1471 (N_1471,N_1336,N_1285);
nand U1472 (N_1472,N_1315,N_1372);
or U1473 (N_1473,N_1391,N_1270);
nor U1474 (N_1474,N_1238,N_1353);
nor U1475 (N_1475,N_1293,N_1302);
nor U1476 (N_1476,N_1201,N_1324);
nand U1477 (N_1477,N_1219,N_1265);
nand U1478 (N_1478,N_1316,N_1267);
nor U1479 (N_1479,N_1335,N_1303);
nor U1480 (N_1480,N_1374,N_1340);
or U1481 (N_1481,N_1280,N_1330);
nand U1482 (N_1482,N_1367,N_1382);
nand U1483 (N_1483,N_1365,N_1362);
nor U1484 (N_1484,N_1326,N_1230);
or U1485 (N_1485,N_1311,N_1346);
nor U1486 (N_1486,N_1272,N_1243);
nor U1487 (N_1487,N_1356,N_1287);
nand U1488 (N_1488,N_1229,N_1329);
and U1489 (N_1489,N_1202,N_1228);
xor U1490 (N_1490,N_1343,N_1288);
and U1491 (N_1491,N_1366,N_1261);
xor U1492 (N_1492,N_1308,N_1337);
and U1493 (N_1493,N_1333,N_1373);
or U1494 (N_1494,N_1320,N_1290);
nand U1495 (N_1495,N_1321,N_1271);
nor U1496 (N_1496,N_1200,N_1245);
xnor U1497 (N_1497,N_1341,N_1387);
or U1498 (N_1498,N_1327,N_1334);
or U1499 (N_1499,N_1379,N_1284);
and U1500 (N_1500,N_1321,N_1220);
or U1501 (N_1501,N_1243,N_1292);
or U1502 (N_1502,N_1345,N_1276);
and U1503 (N_1503,N_1232,N_1228);
nand U1504 (N_1504,N_1393,N_1281);
nand U1505 (N_1505,N_1244,N_1231);
or U1506 (N_1506,N_1394,N_1332);
nand U1507 (N_1507,N_1372,N_1264);
or U1508 (N_1508,N_1360,N_1349);
or U1509 (N_1509,N_1216,N_1211);
nand U1510 (N_1510,N_1381,N_1354);
or U1511 (N_1511,N_1281,N_1251);
xnor U1512 (N_1512,N_1212,N_1239);
and U1513 (N_1513,N_1264,N_1389);
and U1514 (N_1514,N_1211,N_1244);
and U1515 (N_1515,N_1344,N_1281);
or U1516 (N_1516,N_1300,N_1273);
nand U1517 (N_1517,N_1210,N_1314);
nand U1518 (N_1518,N_1343,N_1269);
nor U1519 (N_1519,N_1341,N_1333);
and U1520 (N_1520,N_1377,N_1324);
and U1521 (N_1521,N_1397,N_1352);
or U1522 (N_1522,N_1328,N_1204);
and U1523 (N_1523,N_1214,N_1291);
nand U1524 (N_1524,N_1223,N_1217);
and U1525 (N_1525,N_1361,N_1220);
nor U1526 (N_1526,N_1226,N_1370);
xor U1527 (N_1527,N_1302,N_1254);
and U1528 (N_1528,N_1260,N_1314);
nor U1529 (N_1529,N_1231,N_1353);
nand U1530 (N_1530,N_1224,N_1218);
and U1531 (N_1531,N_1286,N_1250);
nor U1532 (N_1532,N_1212,N_1282);
nand U1533 (N_1533,N_1251,N_1336);
or U1534 (N_1534,N_1279,N_1370);
nand U1535 (N_1535,N_1257,N_1331);
or U1536 (N_1536,N_1355,N_1389);
or U1537 (N_1537,N_1321,N_1229);
or U1538 (N_1538,N_1264,N_1382);
nor U1539 (N_1539,N_1247,N_1242);
nand U1540 (N_1540,N_1397,N_1338);
xnor U1541 (N_1541,N_1260,N_1227);
and U1542 (N_1542,N_1265,N_1326);
and U1543 (N_1543,N_1307,N_1253);
or U1544 (N_1544,N_1318,N_1257);
nor U1545 (N_1545,N_1256,N_1377);
nand U1546 (N_1546,N_1378,N_1346);
xnor U1547 (N_1547,N_1386,N_1290);
or U1548 (N_1548,N_1389,N_1273);
and U1549 (N_1549,N_1336,N_1346);
or U1550 (N_1550,N_1233,N_1255);
and U1551 (N_1551,N_1356,N_1298);
or U1552 (N_1552,N_1376,N_1341);
nand U1553 (N_1553,N_1292,N_1309);
nor U1554 (N_1554,N_1253,N_1282);
and U1555 (N_1555,N_1282,N_1338);
and U1556 (N_1556,N_1277,N_1228);
nand U1557 (N_1557,N_1372,N_1205);
nor U1558 (N_1558,N_1289,N_1371);
and U1559 (N_1559,N_1234,N_1215);
xor U1560 (N_1560,N_1303,N_1267);
or U1561 (N_1561,N_1301,N_1298);
and U1562 (N_1562,N_1244,N_1222);
nand U1563 (N_1563,N_1209,N_1349);
and U1564 (N_1564,N_1237,N_1295);
xor U1565 (N_1565,N_1306,N_1255);
xnor U1566 (N_1566,N_1272,N_1203);
xor U1567 (N_1567,N_1242,N_1386);
nor U1568 (N_1568,N_1330,N_1313);
and U1569 (N_1569,N_1395,N_1305);
nand U1570 (N_1570,N_1205,N_1249);
nor U1571 (N_1571,N_1247,N_1293);
nor U1572 (N_1572,N_1387,N_1321);
nand U1573 (N_1573,N_1215,N_1299);
nor U1574 (N_1574,N_1376,N_1230);
or U1575 (N_1575,N_1252,N_1319);
or U1576 (N_1576,N_1322,N_1398);
xnor U1577 (N_1577,N_1371,N_1300);
nor U1578 (N_1578,N_1333,N_1209);
or U1579 (N_1579,N_1380,N_1248);
and U1580 (N_1580,N_1205,N_1380);
and U1581 (N_1581,N_1259,N_1277);
xor U1582 (N_1582,N_1313,N_1363);
or U1583 (N_1583,N_1238,N_1215);
nor U1584 (N_1584,N_1323,N_1386);
nor U1585 (N_1585,N_1332,N_1311);
nor U1586 (N_1586,N_1280,N_1318);
nand U1587 (N_1587,N_1227,N_1210);
nor U1588 (N_1588,N_1246,N_1372);
xor U1589 (N_1589,N_1323,N_1212);
and U1590 (N_1590,N_1231,N_1213);
xor U1591 (N_1591,N_1335,N_1387);
and U1592 (N_1592,N_1279,N_1246);
xor U1593 (N_1593,N_1296,N_1283);
or U1594 (N_1594,N_1293,N_1284);
nand U1595 (N_1595,N_1349,N_1332);
or U1596 (N_1596,N_1340,N_1255);
or U1597 (N_1597,N_1341,N_1266);
or U1598 (N_1598,N_1302,N_1264);
and U1599 (N_1599,N_1245,N_1228);
or U1600 (N_1600,N_1439,N_1426);
and U1601 (N_1601,N_1511,N_1510);
and U1602 (N_1602,N_1573,N_1427);
or U1603 (N_1603,N_1412,N_1513);
or U1604 (N_1604,N_1588,N_1495);
nor U1605 (N_1605,N_1440,N_1536);
and U1606 (N_1606,N_1425,N_1544);
nor U1607 (N_1607,N_1416,N_1591);
or U1608 (N_1608,N_1414,N_1422);
or U1609 (N_1609,N_1443,N_1404);
or U1610 (N_1610,N_1571,N_1581);
or U1611 (N_1611,N_1428,N_1554);
nand U1612 (N_1612,N_1485,N_1491);
nand U1613 (N_1613,N_1456,N_1558);
or U1614 (N_1614,N_1441,N_1494);
or U1615 (N_1615,N_1519,N_1435);
or U1616 (N_1616,N_1538,N_1432);
or U1617 (N_1617,N_1560,N_1410);
and U1618 (N_1618,N_1406,N_1514);
xor U1619 (N_1619,N_1527,N_1534);
nand U1620 (N_1620,N_1447,N_1460);
or U1621 (N_1621,N_1545,N_1566);
nor U1622 (N_1622,N_1400,N_1457);
nand U1623 (N_1623,N_1501,N_1590);
and U1624 (N_1624,N_1521,N_1535);
nand U1625 (N_1625,N_1508,N_1458);
and U1626 (N_1626,N_1467,N_1587);
or U1627 (N_1627,N_1468,N_1476);
and U1628 (N_1628,N_1431,N_1595);
and U1629 (N_1629,N_1582,N_1503);
nor U1630 (N_1630,N_1483,N_1539);
xnor U1631 (N_1631,N_1482,N_1569);
and U1632 (N_1632,N_1528,N_1478);
and U1633 (N_1633,N_1499,N_1562);
or U1634 (N_1634,N_1515,N_1413);
nand U1635 (N_1635,N_1418,N_1448);
xnor U1636 (N_1636,N_1403,N_1533);
xnor U1637 (N_1637,N_1474,N_1472);
nor U1638 (N_1638,N_1437,N_1520);
nor U1639 (N_1639,N_1434,N_1529);
xnor U1640 (N_1640,N_1524,N_1549);
nand U1641 (N_1641,N_1548,N_1481);
nor U1642 (N_1642,N_1559,N_1461);
or U1643 (N_1643,N_1493,N_1540);
nor U1644 (N_1644,N_1570,N_1579);
nand U1645 (N_1645,N_1585,N_1598);
xor U1646 (N_1646,N_1480,N_1459);
nor U1647 (N_1647,N_1563,N_1543);
nor U1648 (N_1648,N_1522,N_1462);
or U1649 (N_1649,N_1445,N_1479);
and U1650 (N_1650,N_1407,N_1433);
xnor U1651 (N_1651,N_1504,N_1488);
nand U1652 (N_1652,N_1583,N_1594);
nand U1653 (N_1653,N_1596,N_1452);
xnor U1654 (N_1654,N_1575,N_1546);
nor U1655 (N_1655,N_1550,N_1597);
and U1656 (N_1656,N_1506,N_1576);
nand U1657 (N_1657,N_1430,N_1551);
and U1658 (N_1658,N_1516,N_1415);
nor U1659 (N_1659,N_1420,N_1568);
nand U1660 (N_1660,N_1487,N_1417);
and U1661 (N_1661,N_1592,N_1469);
and U1662 (N_1662,N_1401,N_1450);
or U1663 (N_1663,N_1453,N_1564);
nor U1664 (N_1664,N_1475,N_1466);
nand U1665 (N_1665,N_1567,N_1555);
nor U1666 (N_1666,N_1541,N_1486);
nand U1667 (N_1667,N_1577,N_1552);
and U1668 (N_1668,N_1542,N_1484);
and U1669 (N_1669,N_1423,N_1530);
and U1670 (N_1670,N_1537,N_1411);
and U1671 (N_1671,N_1455,N_1565);
nor U1672 (N_1672,N_1593,N_1557);
and U1673 (N_1673,N_1421,N_1589);
or U1674 (N_1674,N_1442,N_1429);
and U1675 (N_1675,N_1465,N_1553);
and U1676 (N_1676,N_1451,N_1502);
xor U1677 (N_1677,N_1578,N_1470);
or U1678 (N_1678,N_1505,N_1526);
nor U1679 (N_1679,N_1492,N_1497);
nor U1680 (N_1680,N_1517,N_1507);
xor U1681 (N_1681,N_1444,N_1556);
or U1682 (N_1682,N_1424,N_1402);
and U1683 (N_1683,N_1454,N_1409);
and U1684 (N_1684,N_1531,N_1496);
nand U1685 (N_1685,N_1580,N_1574);
or U1686 (N_1686,N_1561,N_1405);
nor U1687 (N_1687,N_1532,N_1471);
or U1688 (N_1688,N_1464,N_1489);
or U1689 (N_1689,N_1463,N_1586);
nor U1690 (N_1690,N_1584,N_1490);
nand U1691 (N_1691,N_1518,N_1547);
nor U1692 (N_1692,N_1449,N_1438);
and U1693 (N_1693,N_1572,N_1500);
nand U1694 (N_1694,N_1509,N_1477);
nor U1695 (N_1695,N_1446,N_1525);
nor U1696 (N_1696,N_1473,N_1498);
xor U1697 (N_1697,N_1408,N_1599);
nor U1698 (N_1698,N_1436,N_1523);
or U1699 (N_1699,N_1419,N_1512);
and U1700 (N_1700,N_1548,N_1457);
and U1701 (N_1701,N_1461,N_1579);
nor U1702 (N_1702,N_1509,N_1404);
nand U1703 (N_1703,N_1581,N_1517);
xnor U1704 (N_1704,N_1483,N_1419);
or U1705 (N_1705,N_1453,N_1443);
nor U1706 (N_1706,N_1526,N_1593);
and U1707 (N_1707,N_1447,N_1592);
and U1708 (N_1708,N_1473,N_1564);
or U1709 (N_1709,N_1469,N_1486);
or U1710 (N_1710,N_1491,N_1436);
nor U1711 (N_1711,N_1469,N_1436);
nor U1712 (N_1712,N_1408,N_1435);
nor U1713 (N_1713,N_1520,N_1489);
nor U1714 (N_1714,N_1485,N_1414);
and U1715 (N_1715,N_1535,N_1555);
and U1716 (N_1716,N_1419,N_1560);
and U1717 (N_1717,N_1576,N_1450);
or U1718 (N_1718,N_1591,N_1464);
or U1719 (N_1719,N_1417,N_1409);
nand U1720 (N_1720,N_1421,N_1559);
and U1721 (N_1721,N_1548,N_1441);
nand U1722 (N_1722,N_1467,N_1470);
nand U1723 (N_1723,N_1451,N_1550);
xnor U1724 (N_1724,N_1506,N_1566);
nand U1725 (N_1725,N_1410,N_1527);
nand U1726 (N_1726,N_1445,N_1495);
nand U1727 (N_1727,N_1554,N_1575);
or U1728 (N_1728,N_1407,N_1482);
and U1729 (N_1729,N_1580,N_1410);
nor U1730 (N_1730,N_1453,N_1565);
nor U1731 (N_1731,N_1433,N_1464);
nor U1732 (N_1732,N_1422,N_1502);
and U1733 (N_1733,N_1564,N_1495);
nand U1734 (N_1734,N_1478,N_1532);
or U1735 (N_1735,N_1597,N_1596);
or U1736 (N_1736,N_1407,N_1430);
and U1737 (N_1737,N_1422,N_1456);
xor U1738 (N_1738,N_1414,N_1503);
or U1739 (N_1739,N_1462,N_1434);
nand U1740 (N_1740,N_1426,N_1413);
or U1741 (N_1741,N_1536,N_1409);
nand U1742 (N_1742,N_1477,N_1415);
or U1743 (N_1743,N_1483,N_1502);
nor U1744 (N_1744,N_1458,N_1419);
or U1745 (N_1745,N_1405,N_1570);
or U1746 (N_1746,N_1525,N_1508);
xnor U1747 (N_1747,N_1585,N_1425);
and U1748 (N_1748,N_1552,N_1489);
and U1749 (N_1749,N_1452,N_1419);
xnor U1750 (N_1750,N_1595,N_1527);
and U1751 (N_1751,N_1577,N_1574);
nor U1752 (N_1752,N_1448,N_1581);
or U1753 (N_1753,N_1446,N_1468);
and U1754 (N_1754,N_1401,N_1492);
nor U1755 (N_1755,N_1428,N_1531);
nor U1756 (N_1756,N_1578,N_1475);
or U1757 (N_1757,N_1493,N_1474);
nand U1758 (N_1758,N_1587,N_1469);
nand U1759 (N_1759,N_1405,N_1585);
nand U1760 (N_1760,N_1478,N_1480);
and U1761 (N_1761,N_1445,N_1518);
nand U1762 (N_1762,N_1538,N_1514);
and U1763 (N_1763,N_1478,N_1456);
xnor U1764 (N_1764,N_1516,N_1536);
nor U1765 (N_1765,N_1506,N_1521);
nand U1766 (N_1766,N_1544,N_1462);
and U1767 (N_1767,N_1599,N_1482);
or U1768 (N_1768,N_1532,N_1539);
nor U1769 (N_1769,N_1461,N_1470);
or U1770 (N_1770,N_1457,N_1529);
nand U1771 (N_1771,N_1586,N_1483);
and U1772 (N_1772,N_1467,N_1490);
or U1773 (N_1773,N_1438,N_1545);
nor U1774 (N_1774,N_1453,N_1495);
nand U1775 (N_1775,N_1457,N_1517);
and U1776 (N_1776,N_1406,N_1503);
xnor U1777 (N_1777,N_1427,N_1588);
or U1778 (N_1778,N_1537,N_1538);
xor U1779 (N_1779,N_1548,N_1531);
nand U1780 (N_1780,N_1511,N_1543);
nor U1781 (N_1781,N_1578,N_1484);
or U1782 (N_1782,N_1542,N_1463);
nor U1783 (N_1783,N_1532,N_1480);
xor U1784 (N_1784,N_1510,N_1518);
and U1785 (N_1785,N_1579,N_1547);
nand U1786 (N_1786,N_1534,N_1452);
or U1787 (N_1787,N_1414,N_1440);
nor U1788 (N_1788,N_1576,N_1440);
and U1789 (N_1789,N_1475,N_1469);
nor U1790 (N_1790,N_1414,N_1558);
and U1791 (N_1791,N_1501,N_1553);
or U1792 (N_1792,N_1420,N_1540);
nand U1793 (N_1793,N_1450,N_1460);
nand U1794 (N_1794,N_1496,N_1555);
nand U1795 (N_1795,N_1589,N_1539);
and U1796 (N_1796,N_1559,N_1548);
or U1797 (N_1797,N_1566,N_1485);
nor U1798 (N_1798,N_1429,N_1517);
and U1799 (N_1799,N_1504,N_1425);
nor U1800 (N_1800,N_1654,N_1659);
nand U1801 (N_1801,N_1759,N_1601);
nor U1802 (N_1802,N_1729,N_1734);
and U1803 (N_1803,N_1674,N_1695);
xnor U1804 (N_1804,N_1693,N_1738);
xor U1805 (N_1805,N_1650,N_1651);
nor U1806 (N_1806,N_1747,N_1643);
or U1807 (N_1807,N_1764,N_1687);
and U1808 (N_1808,N_1779,N_1748);
or U1809 (N_1809,N_1602,N_1754);
nand U1810 (N_1810,N_1751,N_1706);
and U1811 (N_1811,N_1620,N_1635);
or U1812 (N_1812,N_1676,N_1797);
and U1813 (N_1813,N_1709,N_1788);
xor U1814 (N_1814,N_1786,N_1740);
nor U1815 (N_1815,N_1767,N_1636);
xnor U1816 (N_1816,N_1613,N_1616);
and U1817 (N_1817,N_1784,N_1609);
nor U1818 (N_1818,N_1691,N_1778);
and U1819 (N_1819,N_1648,N_1789);
nor U1820 (N_1820,N_1624,N_1663);
nor U1821 (N_1821,N_1652,N_1736);
or U1822 (N_1822,N_1628,N_1701);
and U1823 (N_1823,N_1666,N_1717);
nand U1824 (N_1824,N_1697,N_1753);
and U1825 (N_1825,N_1667,N_1684);
nor U1826 (N_1826,N_1661,N_1772);
nor U1827 (N_1827,N_1632,N_1669);
and U1828 (N_1828,N_1735,N_1644);
or U1829 (N_1829,N_1720,N_1639);
and U1830 (N_1830,N_1712,N_1622);
or U1831 (N_1831,N_1699,N_1749);
and U1832 (N_1832,N_1703,N_1606);
and U1833 (N_1833,N_1790,N_1782);
or U1834 (N_1834,N_1645,N_1721);
and U1835 (N_1835,N_1660,N_1785);
or U1836 (N_1836,N_1678,N_1728);
xnor U1837 (N_1837,N_1713,N_1617);
and U1838 (N_1838,N_1682,N_1675);
nand U1839 (N_1839,N_1756,N_1614);
nand U1840 (N_1840,N_1681,N_1683);
and U1841 (N_1841,N_1761,N_1627);
nand U1842 (N_1842,N_1664,N_1704);
xor U1843 (N_1843,N_1630,N_1714);
or U1844 (N_1844,N_1765,N_1696);
nor U1845 (N_1845,N_1724,N_1743);
or U1846 (N_1846,N_1710,N_1711);
or U1847 (N_1847,N_1791,N_1768);
nor U1848 (N_1848,N_1656,N_1780);
nand U1849 (N_1849,N_1757,N_1611);
nor U1850 (N_1850,N_1677,N_1688);
nand U1851 (N_1851,N_1625,N_1771);
and U1852 (N_1852,N_1731,N_1746);
nor U1853 (N_1853,N_1723,N_1774);
nor U1854 (N_1854,N_1670,N_1783);
or U1855 (N_1855,N_1726,N_1744);
nand U1856 (N_1856,N_1727,N_1621);
and U1857 (N_1857,N_1653,N_1618);
nand U1858 (N_1858,N_1775,N_1607);
nor U1859 (N_1859,N_1707,N_1662);
or U1860 (N_1860,N_1629,N_1750);
nand U1861 (N_1861,N_1657,N_1702);
and U1862 (N_1862,N_1686,N_1770);
xor U1863 (N_1863,N_1694,N_1692);
nor U1864 (N_1864,N_1649,N_1762);
and U1865 (N_1865,N_1673,N_1766);
or U1866 (N_1866,N_1631,N_1745);
nor U1867 (N_1867,N_1722,N_1798);
or U1868 (N_1868,N_1795,N_1742);
or U1869 (N_1869,N_1623,N_1741);
nor U1870 (N_1870,N_1689,N_1700);
and U1871 (N_1871,N_1626,N_1679);
or U1872 (N_1872,N_1604,N_1763);
nand U1873 (N_1873,N_1787,N_1752);
nor U1874 (N_1874,N_1793,N_1698);
or U1875 (N_1875,N_1610,N_1655);
nor U1876 (N_1876,N_1603,N_1758);
or U1877 (N_1877,N_1715,N_1605);
or U1878 (N_1878,N_1777,N_1725);
or U1879 (N_1879,N_1796,N_1612);
or U1880 (N_1880,N_1781,N_1640);
or U1881 (N_1881,N_1600,N_1776);
nor U1882 (N_1882,N_1646,N_1633);
and U1883 (N_1883,N_1794,N_1755);
nor U1884 (N_1884,N_1705,N_1619);
and U1885 (N_1885,N_1672,N_1665);
nor U1886 (N_1886,N_1792,N_1716);
or U1887 (N_1887,N_1773,N_1799);
and U1888 (N_1888,N_1769,N_1685);
and U1889 (N_1889,N_1638,N_1732);
and U1890 (N_1890,N_1641,N_1634);
nor U1891 (N_1891,N_1647,N_1637);
or U1892 (N_1892,N_1760,N_1719);
nand U1893 (N_1893,N_1608,N_1733);
nor U1894 (N_1894,N_1680,N_1668);
nand U1895 (N_1895,N_1658,N_1718);
nand U1896 (N_1896,N_1708,N_1615);
nand U1897 (N_1897,N_1671,N_1690);
or U1898 (N_1898,N_1642,N_1739);
xor U1899 (N_1899,N_1737,N_1730);
nand U1900 (N_1900,N_1660,N_1789);
nor U1901 (N_1901,N_1614,N_1678);
and U1902 (N_1902,N_1708,N_1681);
nand U1903 (N_1903,N_1794,N_1634);
or U1904 (N_1904,N_1786,N_1703);
nand U1905 (N_1905,N_1748,N_1793);
nor U1906 (N_1906,N_1710,N_1706);
nor U1907 (N_1907,N_1606,N_1660);
and U1908 (N_1908,N_1705,N_1665);
nand U1909 (N_1909,N_1744,N_1604);
nor U1910 (N_1910,N_1689,N_1610);
nand U1911 (N_1911,N_1711,N_1698);
nand U1912 (N_1912,N_1732,N_1789);
and U1913 (N_1913,N_1736,N_1796);
or U1914 (N_1914,N_1691,N_1612);
nand U1915 (N_1915,N_1618,N_1706);
or U1916 (N_1916,N_1740,N_1769);
xor U1917 (N_1917,N_1715,N_1771);
nand U1918 (N_1918,N_1707,N_1756);
or U1919 (N_1919,N_1753,N_1775);
nor U1920 (N_1920,N_1789,N_1610);
or U1921 (N_1921,N_1770,N_1708);
and U1922 (N_1922,N_1642,N_1789);
and U1923 (N_1923,N_1727,N_1642);
nor U1924 (N_1924,N_1716,N_1647);
or U1925 (N_1925,N_1624,N_1739);
nand U1926 (N_1926,N_1668,N_1713);
and U1927 (N_1927,N_1730,N_1686);
nand U1928 (N_1928,N_1750,N_1645);
and U1929 (N_1929,N_1742,N_1606);
nand U1930 (N_1930,N_1648,N_1702);
xnor U1931 (N_1931,N_1700,N_1748);
nor U1932 (N_1932,N_1769,N_1672);
or U1933 (N_1933,N_1798,N_1634);
nor U1934 (N_1934,N_1723,N_1688);
and U1935 (N_1935,N_1785,N_1721);
nor U1936 (N_1936,N_1648,N_1736);
nand U1937 (N_1937,N_1601,N_1667);
or U1938 (N_1938,N_1670,N_1775);
nand U1939 (N_1939,N_1651,N_1655);
and U1940 (N_1940,N_1641,N_1751);
xnor U1941 (N_1941,N_1782,N_1772);
nand U1942 (N_1942,N_1731,N_1730);
nor U1943 (N_1943,N_1634,N_1781);
nor U1944 (N_1944,N_1643,N_1730);
or U1945 (N_1945,N_1677,N_1794);
nor U1946 (N_1946,N_1658,N_1707);
nand U1947 (N_1947,N_1672,N_1632);
nand U1948 (N_1948,N_1769,N_1675);
or U1949 (N_1949,N_1797,N_1639);
and U1950 (N_1950,N_1782,N_1724);
nor U1951 (N_1951,N_1776,N_1717);
and U1952 (N_1952,N_1635,N_1671);
nor U1953 (N_1953,N_1791,N_1785);
or U1954 (N_1954,N_1611,N_1758);
or U1955 (N_1955,N_1745,N_1641);
nand U1956 (N_1956,N_1779,N_1753);
nor U1957 (N_1957,N_1600,N_1741);
or U1958 (N_1958,N_1641,N_1773);
or U1959 (N_1959,N_1659,N_1625);
or U1960 (N_1960,N_1773,N_1731);
or U1961 (N_1961,N_1712,N_1773);
nor U1962 (N_1962,N_1629,N_1675);
or U1963 (N_1963,N_1748,N_1708);
nand U1964 (N_1964,N_1750,N_1676);
and U1965 (N_1965,N_1791,N_1663);
and U1966 (N_1966,N_1755,N_1775);
nand U1967 (N_1967,N_1758,N_1607);
and U1968 (N_1968,N_1734,N_1606);
or U1969 (N_1969,N_1797,N_1723);
nor U1970 (N_1970,N_1763,N_1601);
xor U1971 (N_1971,N_1634,N_1691);
nor U1972 (N_1972,N_1672,N_1742);
or U1973 (N_1973,N_1693,N_1730);
and U1974 (N_1974,N_1770,N_1791);
nor U1975 (N_1975,N_1721,N_1750);
xnor U1976 (N_1976,N_1731,N_1675);
nor U1977 (N_1977,N_1614,N_1684);
or U1978 (N_1978,N_1624,N_1768);
xor U1979 (N_1979,N_1700,N_1660);
xnor U1980 (N_1980,N_1661,N_1768);
and U1981 (N_1981,N_1726,N_1618);
or U1982 (N_1982,N_1702,N_1780);
nand U1983 (N_1983,N_1612,N_1693);
nor U1984 (N_1984,N_1734,N_1625);
nor U1985 (N_1985,N_1749,N_1672);
or U1986 (N_1986,N_1622,N_1629);
xor U1987 (N_1987,N_1697,N_1743);
and U1988 (N_1988,N_1698,N_1749);
or U1989 (N_1989,N_1608,N_1686);
or U1990 (N_1990,N_1701,N_1650);
nand U1991 (N_1991,N_1657,N_1760);
and U1992 (N_1992,N_1629,N_1667);
or U1993 (N_1993,N_1718,N_1734);
and U1994 (N_1994,N_1603,N_1770);
and U1995 (N_1995,N_1720,N_1716);
or U1996 (N_1996,N_1739,N_1628);
or U1997 (N_1997,N_1715,N_1646);
xor U1998 (N_1998,N_1614,N_1720);
xor U1999 (N_1999,N_1736,N_1787);
or U2000 (N_2000,N_1886,N_1998);
nand U2001 (N_2001,N_1820,N_1822);
and U2002 (N_2002,N_1828,N_1959);
or U2003 (N_2003,N_1964,N_1970);
and U2004 (N_2004,N_1846,N_1803);
or U2005 (N_2005,N_1924,N_1962);
nor U2006 (N_2006,N_1901,N_1871);
nor U2007 (N_2007,N_1911,N_1995);
nand U2008 (N_2008,N_1832,N_1989);
or U2009 (N_2009,N_1807,N_1829);
nor U2010 (N_2010,N_1834,N_1870);
nand U2011 (N_2011,N_1931,N_1999);
and U2012 (N_2012,N_1902,N_1994);
xor U2013 (N_2013,N_1974,N_1900);
nand U2014 (N_2014,N_1950,N_1885);
and U2015 (N_2015,N_1876,N_1958);
nor U2016 (N_2016,N_1963,N_1907);
nor U2017 (N_2017,N_1819,N_1833);
nand U2018 (N_2018,N_1942,N_1977);
and U2019 (N_2019,N_1905,N_1938);
xnor U2020 (N_2020,N_1869,N_1985);
nand U2021 (N_2021,N_1939,N_1957);
nand U2022 (N_2022,N_1872,N_1918);
xnor U2023 (N_2023,N_1838,N_1862);
or U2024 (N_2024,N_1855,N_1866);
nand U2025 (N_2025,N_1880,N_1983);
nor U2026 (N_2026,N_1943,N_1926);
nand U2027 (N_2027,N_1920,N_1839);
nor U2028 (N_2028,N_1849,N_1837);
nand U2029 (N_2029,N_1863,N_1969);
and U2030 (N_2030,N_1945,N_1812);
nand U2031 (N_2031,N_1955,N_1823);
nand U2032 (N_2032,N_1996,N_1993);
or U2033 (N_2033,N_1952,N_1835);
nor U2034 (N_2034,N_1810,N_1878);
nand U2035 (N_2035,N_1818,N_1941);
and U2036 (N_2036,N_1842,N_1960);
or U2037 (N_2037,N_1843,N_1965);
and U2038 (N_2038,N_1917,N_1898);
or U2039 (N_2039,N_1847,N_1806);
xnor U2040 (N_2040,N_1895,N_1897);
and U2041 (N_2041,N_1936,N_1944);
or U2042 (N_2042,N_1916,N_1882);
or U2043 (N_2043,N_1976,N_1861);
or U2044 (N_2044,N_1913,N_1850);
and U2045 (N_2045,N_1830,N_1851);
nand U2046 (N_2046,N_1831,N_1968);
nor U2047 (N_2047,N_1910,N_1903);
nand U2048 (N_2048,N_1987,N_1986);
or U2049 (N_2049,N_1853,N_1802);
nand U2050 (N_2050,N_1899,N_1801);
nand U2051 (N_2051,N_1919,N_1845);
nand U2052 (N_2052,N_1951,N_1877);
nor U2053 (N_2053,N_1841,N_1865);
nand U2054 (N_2054,N_1844,N_1992);
nor U2055 (N_2055,N_1947,N_1981);
and U2056 (N_2056,N_1891,N_1815);
or U2057 (N_2057,N_1930,N_1809);
nand U2058 (N_2058,N_1932,N_1856);
and U2059 (N_2059,N_1873,N_1908);
and U2060 (N_2060,N_1933,N_1982);
or U2061 (N_2061,N_1867,N_1816);
and U2062 (N_2062,N_1953,N_1948);
nor U2063 (N_2063,N_1956,N_1997);
or U2064 (N_2064,N_1805,N_1935);
and U2065 (N_2065,N_1894,N_1949);
and U2066 (N_2066,N_1915,N_1811);
nor U2067 (N_2067,N_1961,N_1854);
nand U2068 (N_2068,N_1984,N_1858);
xnor U2069 (N_2069,N_1940,N_1884);
or U2070 (N_2070,N_1914,N_1966);
or U2071 (N_2071,N_1972,N_1860);
and U2072 (N_2072,N_1883,N_1859);
nor U2073 (N_2073,N_1973,N_1836);
or U2074 (N_2074,N_1922,N_1874);
or U2075 (N_2075,N_1875,N_1821);
nand U2076 (N_2076,N_1808,N_1813);
nand U2077 (N_2077,N_1889,N_1890);
or U2078 (N_2078,N_1909,N_1967);
and U2079 (N_2079,N_1923,N_1840);
or U2080 (N_2080,N_1824,N_1946);
and U2081 (N_2081,N_1925,N_1896);
or U2082 (N_2082,N_1825,N_1800);
and U2083 (N_2083,N_1857,N_1804);
nand U2084 (N_2084,N_1848,N_1881);
nor U2085 (N_2085,N_1827,N_1991);
and U2086 (N_2086,N_1927,N_1904);
and U2087 (N_2087,N_1864,N_1892);
nor U2088 (N_2088,N_1937,N_1906);
or U2089 (N_2089,N_1817,N_1912);
and U2090 (N_2090,N_1954,N_1921);
nor U2091 (N_2091,N_1980,N_1990);
and U2092 (N_2092,N_1928,N_1893);
nor U2093 (N_2093,N_1978,N_1887);
nor U2094 (N_2094,N_1971,N_1826);
and U2095 (N_2095,N_1868,N_1929);
or U2096 (N_2096,N_1879,N_1888);
nor U2097 (N_2097,N_1979,N_1814);
nand U2098 (N_2098,N_1852,N_1934);
and U2099 (N_2099,N_1988,N_1975);
or U2100 (N_2100,N_1855,N_1886);
nor U2101 (N_2101,N_1855,N_1972);
and U2102 (N_2102,N_1833,N_1905);
nand U2103 (N_2103,N_1953,N_1843);
nor U2104 (N_2104,N_1979,N_1878);
or U2105 (N_2105,N_1920,N_1898);
or U2106 (N_2106,N_1972,N_1951);
or U2107 (N_2107,N_1888,N_1944);
nor U2108 (N_2108,N_1914,N_1932);
and U2109 (N_2109,N_1973,N_1859);
nor U2110 (N_2110,N_1898,N_1947);
or U2111 (N_2111,N_1882,N_1981);
or U2112 (N_2112,N_1842,N_1869);
nand U2113 (N_2113,N_1809,N_1983);
nand U2114 (N_2114,N_1907,N_1872);
nand U2115 (N_2115,N_1992,N_1850);
or U2116 (N_2116,N_1916,N_1908);
or U2117 (N_2117,N_1878,N_1848);
nand U2118 (N_2118,N_1908,N_1992);
and U2119 (N_2119,N_1836,N_1932);
nand U2120 (N_2120,N_1849,N_1947);
nor U2121 (N_2121,N_1839,N_1834);
nand U2122 (N_2122,N_1866,N_1845);
or U2123 (N_2123,N_1917,N_1848);
or U2124 (N_2124,N_1921,N_1900);
nor U2125 (N_2125,N_1964,N_1987);
xor U2126 (N_2126,N_1869,N_1968);
nor U2127 (N_2127,N_1989,N_1948);
or U2128 (N_2128,N_1939,N_1960);
nor U2129 (N_2129,N_1910,N_1965);
and U2130 (N_2130,N_1903,N_1820);
or U2131 (N_2131,N_1988,N_1961);
or U2132 (N_2132,N_1999,N_1860);
nand U2133 (N_2133,N_1849,N_1949);
nand U2134 (N_2134,N_1883,N_1869);
nor U2135 (N_2135,N_1943,N_1909);
and U2136 (N_2136,N_1941,N_1974);
nor U2137 (N_2137,N_1891,N_1897);
or U2138 (N_2138,N_1873,N_1859);
xor U2139 (N_2139,N_1981,N_1895);
or U2140 (N_2140,N_1810,N_1835);
xor U2141 (N_2141,N_1852,N_1936);
or U2142 (N_2142,N_1841,N_1959);
nand U2143 (N_2143,N_1837,N_1893);
nor U2144 (N_2144,N_1960,N_1897);
or U2145 (N_2145,N_1967,N_1886);
and U2146 (N_2146,N_1869,N_1903);
and U2147 (N_2147,N_1998,N_1934);
and U2148 (N_2148,N_1805,N_1847);
nand U2149 (N_2149,N_1826,N_1961);
nor U2150 (N_2150,N_1880,N_1960);
nand U2151 (N_2151,N_1945,N_1842);
nand U2152 (N_2152,N_1869,N_1839);
and U2153 (N_2153,N_1892,N_1860);
nor U2154 (N_2154,N_1983,N_1891);
and U2155 (N_2155,N_1881,N_1841);
or U2156 (N_2156,N_1965,N_1959);
nand U2157 (N_2157,N_1818,N_1871);
nand U2158 (N_2158,N_1897,N_1811);
nor U2159 (N_2159,N_1884,N_1996);
nand U2160 (N_2160,N_1842,N_1903);
or U2161 (N_2161,N_1915,N_1911);
nor U2162 (N_2162,N_1942,N_1908);
xnor U2163 (N_2163,N_1891,N_1901);
or U2164 (N_2164,N_1853,N_1979);
nand U2165 (N_2165,N_1958,N_1932);
xor U2166 (N_2166,N_1925,N_1827);
and U2167 (N_2167,N_1824,N_1973);
nand U2168 (N_2168,N_1872,N_1843);
xor U2169 (N_2169,N_1841,N_1857);
and U2170 (N_2170,N_1869,N_1934);
or U2171 (N_2171,N_1818,N_1975);
and U2172 (N_2172,N_1988,N_1919);
nor U2173 (N_2173,N_1906,N_1908);
or U2174 (N_2174,N_1813,N_1824);
nor U2175 (N_2175,N_1901,N_1870);
xnor U2176 (N_2176,N_1950,N_1849);
and U2177 (N_2177,N_1868,N_1954);
nand U2178 (N_2178,N_1876,N_1909);
xor U2179 (N_2179,N_1938,N_1804);
or U2180 (N_2180,N_1988,N_1938);
nand U2181 (N_2181,N_1990,N_1913);
nor U2182 (N_2182,N_1938,N_1858);
nand U2183 (N_2183,N_1986,N_1910);
xnor U2184 (N_2184,N_1880,N_1873);
nand U2185 (N_2185,N_1992,N_1870);
or U2186 (N_2186,N_1822,N_1869);
nor U2187 (N_2187,N_1903,N_1813);
or U2188 (N_2188,N_1908,N_1854);
or U2189 (N_2189,N_1807,N_1835);
nor U2190 (N_2190,N_1827,N_1918);
nand U2191 (N_2191,N_1922,N_1968);
or U2192 (N_2192,N_1999,N_1974);
nor U2193 (N_2193,N_1979,N_1912);
nor U2194 (N_2194,N_1933,N_1804);
nor U2195 (N_2195,N_1997,N_1979);
or U2196 (N_2196,N_1838,N_1946);
nor U2197 (N_2197,N_1889,N_1852);
nand U2198 (N_2198,N_1872,N_1946);
and U2199 (N_2199,N_1993,N_1960);
and U2200 (N_2200,N_2082,N_2195);
or U2201 (N_2201,N_2060,N_2168);
or U2202 (N_2202,N_2027,N_2096);
nand U2203 (N_2203,N_2038,N_2137);
and U2204 (N_2204,N_2190,N_2171);
nand U2205 (N_2205,N_2126,N_2138);
or U2206 (N_2206,N_2173,N_2165);
or U2207 (N_2207,N_2024,N_2158);
nand U2208 (N_2208,N_2054,N_2150);
nand U2209 (N_2209,N_2066,N_2067);
nand U2210 (N_2210,N_2028,N_2118);
and U2211 (N_2211,N_2000,N_2035);
and U2212 (N_2212,N_2089,N_2070);
nand U2213 (N_2213,N_2104,N_2194);
nor U2214 (N_2214,N_2045,N_2065);
nor U2215 (N_2215,N_2021,N_2123);
and U2216 (N_2216,N_2134,N_2074);
nand U2217 (N_2217,N_2196,N_2088);
nand U2218 (N_2218,N_2050,N_2181);
nor U2219 (N_2219,N_2077,N_2078);
nor U2220 (N_2220,N_2106,N_2182);
nor U2221 (N_2221,N_2046,N_2175);
or U2222 (N_2222,N_2189,N_2115);
nor U2223 (N_2223,N_2052,N_2125);
nor U2224 (N_2224,N_2133,N_2107);
xnor U2225 (N_2225,N_2031,N_2009);
nand U2226 (N_2226,N_2049,N_2162);
nor U2227 (N_2227,N_2041,N_2176);
nand U2228 (N_2228,N_2006,N_2091);
and U2229 (N_2229,N_2018,N_2116);
xor U2230 (N_2230,N_2166,N_2111);
nor U2231 (N_2231,N_2174,N_2167);
or U2232 (N_2232,N_2026,N_2183);
nor U2233 (N_2233,N_2131,N_2101);
nand U2234 (N_2234,N_2136,N_2081);
and U2235 (N_2235,N_2037,N_2142);
nand U2236 (N_2236,N_2029,N_2177);
nand U2237 (N_2237,N_2008,N_2072);
and U2238 (N_2238,N_2170,N_2073);
nor U2239 (N_2239,N_2080,N_2120);
or U2240 (N_2240,N_2097,N_2003);
or U2241 (N_2241,N_2087,N_2098);
nand U2242 (N_2242,N_2139,N_2053);
and U2243 (N_2243,N_2076,N_2057);
nor U2244 (N_2244,N_2085,N_2005);
nor U2245 (N_2245,N_2105,N_2071);
nor U2246 (N_2246,N_2033,N_2148);
nor U2247 (N_2247,N_2153,N_2068);
nand U2248 (N_2248,N_2199,N_2132);
or U2249 (N_2249,N_2099,N_2164);
nor U2250 (N_2250,N_2193,N_2079);
and U2251 (N_2251,N_2093,N_2017);
and U2252 (N_2252,N_2198,N_2184);
or U2253 (N_2253,N_2015,N_2157);
and U2254 (N_2254,N_2064,N_2180);
nor U2255 (N_2255,N_2112,N_2151);
or U2256 (N_2256,N_2061,N_2141);
nor U2257 (N_2257,N_2127,N_2025);
and U2258 (N_2258,N_2178,N_2013);
and U2259 (N_2259,N_2149,N_2040);
xnor U2260 (N_2260,N_2179,N_2161);
xnor U2261 (N_2261,N_2192,N_2022);
nor U2262 (N_2262,N_2113,N_2187);
and U2263 (N_2263,N_2119,N_2083);
nor U2264 (N_2264,N_2020,N_2156);
nand U2265 (N_2265,N_2172,N_2152);
or U2266 (N_2266,N_2145,N_2154);
nor U2267 (N_2267,N_2129,N_2014);
nor U2268 (N_2268,N_2042,N_2100);
or U2269 (N_2269,N_2135,N_2095);
nor U2270 (N_2270,N_2011,N_2016);
nand U2271 (N_2271,N_2144,N_2147);
or U2272 (N_2272,N_2128,N_2036);
or U2273 (N_2273,N_2090,N_2086);
and U2274 (N_2274,N_2047,N_2103);
nor U2275 (N_2275,N_2058,N_2169);
nand U2276 (N_2276,N_2160,N_2124);
and U2277 (N_2277,N_2084,N_2117);
xor U2278 (N_2278,N_2102,N_2043);
nor U2279 (N_2279,N_2039,N_2010);
nor U2280 (N_2280,N_2002,N_2012);
or U2281 (N_2281,N_2030,N_2069);
nor U2282 (N_2282,N_2007,N_2122);
nor U2283 (N_2283,N_2109,N_2110);
nand U2284 (N_2284,N_2140,N_2019);
nor U2285 (N_2285,N_2004,N_2063);
and U2286 (N_2286,N_2055,N_2023);
nor U2287 (N_2287,N_2114,N_2001);
and U2288 (N_2288,N_2075,N_2059);
nand U2289 (N_2289,N_2188,N_2108);
or U2290 (N_2290,N_2186,N_2143);
and U2291 (N_2291,N_2034,N_2130);
and U2292 (N_2292,N_2032,N_2062);
or U2293 (N_2293,N_2163,N_2044);
xor U2294 (N_2294,N_2094,N_2092);
nand U2295 (N_2295,N_2121,N_2185);
or U2296 (N_2296,N_2048,N_2146);
nor U2297 (N_2297,N_2191,N_2197);
nor U2298 (N_2298,N_2155,N_2056);
and U2299 (N_2299,N_2051,N_2159);
or U2300 (N_2300,N_2137,N_2188);
and U2301 (N_2301,N_2072,N_2131);
and U2302 (N_2302,N_2080,N_2013);
nor U2303 (N_2303,N_2115,N_2051);
and U2304 (N_2304,N_2019,N_2076);
or U2305 (N_2305,N_2072,N_2023);
and U2306 (N_2306,N_2057,N_2027);
or U2307 (N_2307,N_2047,N_2118);
nand U2308 (N_2308,N_2004,N_2177);
and U2309 (N_2309,N_2046,N_2138);
xor U2310 (N_2310,N_2136,N_2061);
or U2311 (N_2311,N_2172,N_2146);
or U2312 (N_2312,N_2001,N_2103);
nand U2313 (N_2313,N_2069,N_2008);
and U2314 (N_2314,N_2195,N_2025);
nor U2315 (N_2315,N_2140,N_2146);
and U2316 (N_2316,N_2079,N_2065);
nor U2317 (N_2317,N_2150,N_2075);
nand U2318 (N_2318,N_2003,N_2001);
or U2319 (N_2319,N_2164,N_2118);
nor U2320 (N_2320,N_2066,N_2070);
or U2321 (N_2321,N_2056,N_2062);
or U2322 (N_2322,N_2185,N_2036);
and U2323 (N_2323,N_2102,N_2093);
or U2324 (N_2324,N_2142,N_2121);
and U2325 (N_2325,N_2053,N_2043);
and U2326 (N_2326,N_2012,N_2057);
or U2327 (N_2327,N_2093,N_2158);
nor U2328 (N_2328,N_2126,N_2023);
nand U2329 (N_2329,N_2192,N_2026);
or U2330 (N_2330,N_2087,N_2089);
nand U2331 (N_2331,N_2192,N_2111);
nand U2332 (N_2332,N_2144,N_2073);
nand U2333 (N_2333,N_2011,N_2181);
and U2334 (N_2334,N_2118,N_2183);
nand U2335 (N_2335,N_2123,N_2110);
or U2336 (N_2336,N_2103,N_2003);
nand U2337 (N_2337,N_2031,N_2004);
nor U2338 (N_2338,N_2132,N_2045);
nand U2339 (N_2339,N_2062,N_2175);
xnor U2340 (N_2340,N_2135,N_2048);
nand U2341 (N_2341,N_2120,N_2107);
and U2342 (N_2342,N_2107,N_2195);
nand U2343 (N_2343,N_2145,N_2196);
and U2344 (N_2344,N_2094,N_2085);
nor U2345 (N_2345,N_2044,N_2191);
and U2346 (N_2346,N_2166,N_2075);
and U2347 (N_2347,N_2007,N_2042);
nor U2348 (N_2348,N_2145,N_2108);
nand U2349 (N_2349,N_2147,N_2042);
nand U2350 (N_2350,N_2174,N_2018);
nor U2351 (N_2351,N_2063,N_2007);
nand U2352 (N_2352,N_2055,N_2138);
nor U2353 (N_2353,N_2183,N_2052);
nand U2354 (N_2354,N_2062,N_2053);
or U2355 (N_2355,N_2179,N_2083);
or U2356 (N_2356,N_2004,N_2108);
and U2357 (N_2357,N_2128,N_2154);
or U2358 (N_2358,N_2158,N_2103);
xnor U2359 (N_2359,N_2078,N_2182);
nand U2360 (N_2360,N_2068,N_2064);
nand U2361 (N_2361,N_2099,N_2142);
or U2362 (N_2362,N_2157,N_2192);
nand U2363 (N_2363,N_2178,N_2078);
or U2364 (N_2364,N_2165,N_2132);
and U2365 (N_2365,N_2150,N_2116);
and U2366 (N_2366,N_2147,N_2104);
nand U2367 (N_2367,N_2013,N_2193);
and U2368 (N_2368,N_2176,N_2183);
and U2369 (N_2369,N_2191,N_2136);
and U2370 (N_2370,N_2180,N_2031);
nor U2371 (N_2371,N_2184,N_2046);
nor U2372 (N_2372,N_2100,N_2168);
xnor U2373 (N_2373,N_2032,N_2002);
or U2374 (N_2374,N_2113,N_2061);
or U2375 (N_2375,N_2115,N_2098);
xnor U2376 (N_2376,N_2040,N_2094);
xnor U2377 (N_2377,N_2008,N_2042);
nor U2378 (N_2378,N_2189,N_2198);
nor U2379 (N_2379,N_2054,N_2091);
xor U2380 (N_2380,N_2173,N_2004);
nand U2381 (N_2381,N_2079,N_2162);
nand U2382 (N_2382,N_2086,N_2117);
or U2383 (N_2383,N_2077,N_2101);
and U2384 (N_2384,N_2079,N_2158);
and U2385 (N_2385,N_2022,N_2007);
nor U2386 (N_2386,N_2034,N_2041);
or U2387 (N_2387,N_2013,N_2139);
xnor U2388 (N_2388,N_2107,N_2198);
nand U2389 (N_2389,N_2199,N_2021);
nand U2390 (N_2390,N_2006,N_2070);
xnor U2391 (N_2391,N_2181,N_2165);
and U2392 (N_2392,N_2143,N_2069);
and U2393 (N_2393,N_2161,N_2101);
nor U2394 (N_2394,N_2100,N_2125);
and U2395 (N_2395,N_2069,N_2080);
xnor U2396 (N_2396,N_2145,N_2159);
nand U2397 (N_2397,N_2050,N_2149);
nor U2398 (N_2398,N_2162,N_2042);
nand U2399 (N_2399,N_2112,N_2094);
nand U2400 (N_2400,N_2227,N_2342);
xnor U2401 (N_2401,N_2250,N_2302);
nand U2402 (N_2402,N_2310,N_2350);
nand U2403 (N_2403,N_2271,N_2234);
nand U2404 (N_2404,N_2289,N_2371);
or U2405 (N_2405,N_2214,N_2359);
and U2406 (N_2406,N_2273,N_2333);
nand U2407 (N_2407,N_2389,N_2329);
or U2408 (N_2408,N_2279,N_2379);
nand U2409 (N_2409,N_2259,N_2318);
nand U2410 (N_2410,N_2395,N_2293);
or U2411 (N_2411,N_2363,N_2282);
nand U2412 (N_2412,N_2233,N_2303);
or U2413 (N_2413,N_2235,N_2205);
nand U2414 (N_2414,N_2320,N_2291);
or U2415 (N_2415,N_2284,N_2392);
xnor U2416 (N_2416,N_2307,N_2322);
and U2417 (N_2417,N_2203,N_2280);
nand U2418 (N_2418,N_2399,N_2351);
nor U2419 (N_2419,N_2255,N_2372);
xnor U2420 (N_2420,N_2297,N_2364);
and U2421 (N_2421,N_2335,N_2346);
nor U2422 (N_2422,N_2380,N_2308);
nand U2423 (N_2423,N_2296,N_2356);
or U2424 (N_2424,N_2301,N_2281);
xnor U2425 (N_2425,N_2261,N_2394);
and U2426 (N_2426,N_2200,N_2253);
and U2427 (N_2427,N_2258,N_2278);
or U2428 (N_2428,N_2388,N_2215);
or U2429 (N_2429,N_2304,N_2377);
nor U2430 (N_2430,N_2263,N_2332);
nand U2431 (N_2431,N_2376,N_2343);
or U2432 (N_2432,N_2353,N_2375);
nor U2433 (N_2433,N_2202,N_2286);
nand U2434 (N_2434,N_2244,N_2219);
xnor U2435 (N_2435,N_2225,N_2257);
and U2436 (N_2436,N_2306,N_2339);
nor U2437 (N_2437,N_2374,N_2313);
nand U2438 (N_2438,N_2347,N_2331);
or U2439 (N_2439,N_2209,N_2276);
or U2440 (N_2440,N_2290,N_2327);
xor U2441 (N_2441,N_2260,N_2230);
nand U2442 (N_2442,N_2217,N_2210);
nor U2443 (N_2443,N_2254,N_2393);
and U2444 (N_2444,N_2245,N_2362);
or U2445 (N_2445,N_2211,N_2323);
nor U2446 (N_2446,N_2358,N_2311);
nor U2447 (N_2447,N_2221,N_2229);
nor U2448 (N_2448,N_2352,N_2365);
and U2449 (N_2449,N_2228,N_2348);
nor U2450 (N_2450,N_2206,N_2237);
and U2451 (N_2451,N_2295,N_2357);
xnor U2452 (N_2452,N_2370,N_2220);
nor U2453 (N_2453,N_2288,N_2266);
nor U2454 (N_2454,N_2269,N_2275);
and U2455 (N_2455,N_2272,N_2345);
nor U2456 (N_2456,N_2251,N_2319);
or U2457 (N_2457,N_2246,N_2224);
nand U2458 (N_2458,N_2368,N_2277);
or U2459 (N_2459,N_2262,N_2315);
or U2460 (N_2460,N_2238,N_2354);
nand U2461 (N_2461,N_2326,N_2212);
and U2462 (N_2462,N_2330,N_2213);
or U2463 (N_2463,N_2385,N_2216);
xnor U2464 (N_2464,N_2242,N_2397);
and U2465 (N_2465,N_2270,N_2314);
or U2466 (N_2466,N_2325,N_2316);
nand U2467 (N_2467,N_2344,N_2373);
nor U2468 (N_2468,N_2252,N_2309);
nand U2469 (N_2469,N_2249,N_2384);
and U2470 (N_2470,N_2223,N_2240);
xnor U2471 (N_2471,N_2369,N_2265);
or U2472 (N_2472,N_2360,N_2232);
or U2473 (N_2473,N_2247,N_2267);
nand U2474 (N_2474,N_2366,N_2243);
nor U2475 (N_2475,N_2317,N_2248);
xnor U2476 (N_2476,N_2338,N_2231);
nor U2477 (N_2477,N_2387,N_2299);
and U2478 (N_2478,N_2341,N_2355);
or U2479 (N_2479,N_2298,N_2239);
and U2480 (N_2480,N_2305,N_2256);
xor U2481 (N_2481,N_2367,N_2336);
xor U2482 (N_2482,N_2340,N_2381);
or U2483 (N_2483,N_2398,N_2274);
and U2484 (N_2484,N_2218,N_2226);
nand U2485 (N_2485,N_2264,N_2321);
nor U2486 (N_2486,N_2312,N_2396);
or U2487 (N_2487,N_2241,N_2283);
nor U2488 (N_2488,N_2349,N_2300);
nor U2489 (N_2489,N_2208,N_2268);
nand U2490 (N_2490,N_2236,N_2383);
or U2491 (N_2491,N_2386,N_2390);
or U2492 (N_2492,N_2204,N_2337);
nand U2493 (N_2493,N_2222,N_2294);
and U2494 (N_2494,N_2382,N_2201);
nor U2495 (N_2495,N_2324,N_2287);
or U2496 (N_2496,N_2207,N_2334);
nand U2497 (N_2497,N_2328,N_2391);
and U2498 (N_2498,N_2285,N_2361);
and U2499 (N_2499,N_2292,N_2378);
and U2500 (N_2500,N_2338,N_2378);
and U2501 (N_2501,N_2203,N_2297);
xor U2502 (N_2502,N_2283,N_2351);
and U2503 (N_2503,N_2223,N_2315);
and U2504 (N_2504,N_2309,N_2225);
nor U2505 (N_2505,N_2247,N_2272);
nor U2506 (N_2506,N_2399,N_2305);
nor U2507 (N_2507,N_2221,N_2341);
xnor U2508 (N_2508,N_2226,N_2279);
nor U2509 (N_2509,N_2330,N_2283);
nor U2510 (N_2510,N_2295,N_2283);
and U2511 (N_2511,N_2217,N_2286);
nor U2512 (N_2512,N_2208,N_2275);
or U2513 (N_2513,N_2262,N_2287);
nor U2514 (N_2514,N_2342,N_2264);
or U2515 (N_2515,N_2220,N_2358);
xnor U2516 (N_2516,N_2369,N_2270);
nor U2517 (N_2517,N_2340,N_2237);
and U2518 (N_2518,N_2270,N_2376);
and U2519 (N_2519,N_2265,N_2347);
and U2520 (N_2520,N_2202,N_2231);
and U2521 (N_2521,N_2367,N_2294);
nor U2522 (N_2522,N_2210,N_2288);
or U2523 (N_2523,N_2316,N_2329);
nand U2524 (N_2524,N_2245,N_2285);
xor U2525 (N_2525,N_2372,N_2337);
or U2526 (N_2526,N_2290,N_2292);
and U2527 (N_2527,N_2219,N_2212);
nor U2528 (N_2528,N_2223,N_2254);
or U2529 (N_2529,N_2215,N_2335);
or U2530 (N_2530,N_2303,N_2336);
nor U2531 (N_2531,N_2331,N_2286);
nor U2532 (N_2532,N_2334,N_2339);
xor U2533 (N_2533,N_2286,N_2236);
or U2534 (N_2534,N_2202,N_2266);
nor U2535 (N_2535,N_2221,N_2231);
nor U2536 (N_2536,N_2394,N_2372);
or U2537 (N_2537,N_2374,N_2219);
and U2538 (N_2538,N_2323,N_2304);
xor U2539 (N_2539,N_2242,N_2382);
or U2540 (N_2540,N_2295,N_2392);
nand U2541 (N_2541,N_2241,N_2231);
or U2542 (N_2542,N_2397,N_2377);
nand U2543 (N_2543,N_2292,N_2256);
and U2544 (N_2544,N_2260,N_2280);
and U2545 (N_2545,N_2373,N_2380);
and U2546 (N_2546,N_2367,N_2342);
nand U2547 (N_2547,N_2239,N_2213);
nand U2548 (N_2548,N_2263,N_2210);
and U2549 (N_2549,N_2262,N_2239);
xnor U2550 (N_2550,N_2252,N_2232);
nor U2551 (N_2551,N_2278,N_2229);
and U2552 (N_2552,N_2286,N_2295);
nor U2553 (N_2553,N_2267,N_2234);
nand U2554 (N_2554,N_2221,N_2307);
and U2555 (N_2555,N_2359,N_2284);
or U2556 (N_2556,N_2298,N_2336);
nor U2557 (N_2557,N_2392,N_2288);
and U2558 (N_2558,N_2287,N_2383);
nand U2559 (N_2559,N_2357,N_2367);
or U2560 (N_2560,N_2242,N_2324);
nand U2561 (N_2561,N_2220,N_2331);
nor U2562 (N_2562,N_2372,N_2378);
nand U2563 (N_2563,N_2384,N_2345);
or U2564 (N_2564,N_2291,N_2363);
nand U2565 (N_2565,N_2298,N_2226);
nand U2566 (N_2566,N_2365,N_2368);
nand U2567 (N_2567,N_2200,N_2283);
and U2568 (N_2568,N_2392,N_2214);
nor U2569 (N_2569,N_2336,N_2347);
xnor U2570 (N_2570,N_2255,N_2257);
nor U2571 (N_2571,N_2370,N_2265);
or U2572 (N_2572,N_2239,N_2216);
nand U2573 (N_2573,N_2305,N_2279);
nor U2574 (N_2574,N_2363,N_2259);
or U2575 (N_2575,N_2389,N_2207);
nand U2576 (N_2576,N_2280,N_2307);
and U2577 (N_2577,N_2279,N_2388);
and U2578 (N_2578,N_2286,N_2279);
and U2579 (N_2579,N_2320,N_2376);
or U2580 (N_2580,N_2204,N_2393);
nor U2581 (N_2581,N_2209,N_2348);
or U2582 (N_2582,N_2397,N_2337);
nand U2583 (N_2583,N_2217,N_2271);
and U2584 (N_2584,N_2238,N_2233);
or U2585 (N_2585,N_2387,N_2221);
nor U2586 (N_2586,N_2207,N_2232);
nand U2587 (N_2587,N_2275,N_2200);
nand U2588 (N_2588,N_2334,N_2211);
nand U2589 (N_2589,N_2216,N_2272);
and U2590 (N_2590,N_2353,N_2380);
and U2591 (N_2591,N_2382,N_2359);
nor U2592 (N_2592,N_2338,N_2208);
and U2593 (N_2593,N_2222,N_2312);
nor U2594 (N_2594,N_2210,N_2214);
or U2595 (N_2595,N_2371,N_2257);
nor U2596 (N_2596,N_2396,N_2360);
and U2597 (N_2597,N_2272,N_2302);
and U2598 (N_2598,N_2345,N_2305);
or U2599 (N_2599,N_2380,N_2240);
nand U2600 (N_2600,N_2529,N_2464);
and U2601 (N_2601,N_2533,N_2522);
and U2602 (N_2602,N_2572,N_2558);
xor U2603 (N_2603,N_2591,N_2501);
xor U2604 (N_2604,N_2581,N_2478);
xnor U2605 (N_2605,N_2513,N_2553);
or U2606 (N_2606,N_2521,N_2406);
nand U2607 (N_2607,N_2476,N_2416);
nand U2608 (N_2608,N_2577,N_2466);
nand U2609 (N_2609,N_2550,N_2411);
xor U2610 (N_2610,N_2597,N_2505);
or U2611 (N_2611,N_2497,N_2530);
and U2612 (N_2612,N_2480,N_2507);
and U2613 (N_2613,N_2410,N_2515);
nor U2614 (N_2614,N_2576,N_2578);
and U2615 (N_2615,N_2523,N_2491);
nand U2616 (N_2616,N_2528,N_2459);
xor U2617 (N_2617,N_2428,N_2437);
nand U2618 (N_2618,N_2592,N_2451);
nor U2619 (N_2619,N_2403,N_2421);
nor U2620 (N_2620,N_2573,N_2435);
nor U2621 (N_2621,N_2520,N_2537);
or U2622 (N_2622,N_2482,N_2462);
xor U2623 (N_2623,N_2444,N_2594);
or U2624 (N_2624,N_2479,N_2542);
or U2625 (N_2625,N_2559,N_2524);
and U2626 (N_2626,N_2471,N_2575);
nand U2627 (N_2627,N_2568,N_2427);
and U2628 (N_2628,N_2450,N_2541);
or U2629 (N_2629,N_2493,N_2404);
xnor U2630 (N_2630,N_2409,N_2408);
xor U2631 (N_2631,N_2546,N_2475);
nand U2632 (N_2632,N_2543,N_2548);
or U2633 (N_2633,N_2489,N_2526);
nand U2634 (N_2634,N_2596,N_2422);
nand U2635 (N_2635,N_2414,N_2472);
xor U2636 (N_2636,N_2441,N_2419);
nor U2637 (N_2637,N_2487,N_2467);
and U2638 (N_2638,N_2498,N_2590);
or U2639 (N_2639,N_2585,N_2506);
or U2640 (N_2640,N_2504,N_2536);
and U2641 (N_2641,N_2439,N_2514);
xnor U2642 (N_2642,N_2458,N_2418);
and U2643 (N_2643,N_2447,N_2502);
or U2644 (N_2644,N_2474,N_2566);
and U2645 (N_2645,N_2547,N_2510);
and U2646 (N_2646,N_2534,N_2432);
nor U2647 (N_2647,N_2426,N_2595);
and U2648 (N_2648,N_2424,N_2454);
and U2649 (N_2649,N_2516,N_2519);
or U2650 (N_2650,N_2486,N_2512);
or U2651 (N_2651,N_2492,N_2425);
nand U2652 (N_2652,N_2582,N_2400);
and U2653 (N_2653,N_2586,N_2571);
and U2654 (N_2654,N_2412,N_2455);
nand U2655 (N_2655,N_2517,N_2552);
or U2656 (N_2656,N_2442,N_2511);
nor U2657 (N_2657,N_2490,N_2584);
nor U2658 (N_2658,N_2465,N_2405);
nand U2659 (N_2659,N_2461,N_2446);
nand U2660 (N_2660,N_2555,N_2463);
nor U2661 (N_2661,N_2440,N_2593);
or U2662 (N_2662,N_2433,N_2434);
and U2663 (N_2663,N_2532,N_2431);
nor U2664 (N_2664,N_2583,N_2495);
and U2665 (N_2665,N_2554,N_2560);
or U2666 (N_2666,N_2557,N_2415);
or U2667 (N_2667,N_2556,N_2470);
nor U2668 (N_2668,N_2598,N_2488);
and U2669 (N_2669,N_2564,N_2494);
xnor U2670 (N_2670,N_2587,N_2449);
nand U2671 (N_2671,N_2509,N_2599);
or U2672 (N_2672,N_2545,N_2429);
and U2673 (N_2673,N_2539,N_2473);
or U2674 (N_2674,N_2484,N_2570);
nor U2675 (N_2675,N_2496,N_2574);
nor U2676 (N_2676,N_2452,N_2540);
nor U2677 (N_2677,N_2469,N_2417);
and U2678 (N_2678,N_2535,N_2565);
and U2679 (N_2679,N_2485,N_2456);
nor U2680 (N_2680,N_2538,N_2460);
and U2681 (N_2681,N_2457,N_2567);
nor U2682 (N_2682,N_2436,N_2525);
or U2683 (N_2683,N_2551,N_2563);
nor U2684 (N_2684,N_2544,N_2561);
and U2685 (N_2685,N_2443,N_2468);
nand U2686 (N_2686,N_2562,N_2549);
or U2687 (N_2687,N_2481,N_2531);
and U2688 (N_2688,N_2518,N_2420);
and U2689 (N_2689,N_2477,N_2569);
and U2690 (N_2690,N_2503,N_2499);
xnor U2691 (N_2691,N_2453,N_2430);
or U2692 (N_2692,N_2407,N_2423);
and U2693 (N_2693,N_2579,N_2402);
or U2694 (N_2694,N_2580,N_2588);
nand U2695 (N_2695,N_2438,N_2445);
nand U2696 (N_2696,N_2500,N_2448);
or U2697 (N_2697,N_2508,N_2483);
nor U2698 (N_2698,N_2401,N_2413);
or U2699 (N_2699,N_2589,N_2527);
and U2700 (N_2700,N_2464,N_2545);
and U2701 (N_2701,N_2426,N_2518);
and U2702 (N_2702,N_2492,N_2435);
and U2703 (N_2703,N_2498,N_2400);
and U2704 (N_2704,N_2404,N_2578);
and U2705 (N_2705,N_2443,N_2440);
and U2706 (N_2706,N_2584,N_2469);
or U2707 (N_2707,N_2579,N_2599);
nor U2708 (N_2708,N_2501,N_2528);
or U2709 (N_2709,N_2544,N_2516);
and U2710 (N_2710,N_2573,N_2567);
nand U2711 (N_2711,N_2488,N_2538);
and U2712 (N_2712,N_2514,N_2522);
nand U2713 (N_2713,N_2584,N_2452);
or U2714 (N_2714,N_2516,N_2573);
nand U2715 (N_2715,N_2599,N_2431);
xor U2716 (N_2716,N_2497,N_2470);
and U2717 (N_2717,N_2517,N_2461);
and U2718 (N_2718,N_2549,N_2572);
and U2719 (N_2719,N_2450,N_2406);
and U2720 (N_2720,N_2473,N_2576);
and U2721 (N_2721,N_2534,N_2578);
and U2722 (N_2722,N_2531,N_2504);
or U2723 (N_2723,N_2452,N_2565);
nand U2724 (N_2724,N_2415,N_2451);
and U2725 (N_2725,N_2588,N_2521);
nor U2726 (N_2726,N_2513,N_2514);
xnor U2727 (N_2727,N_2420,N_2458);
nor U2728 (N_2728,N_2461,N_2578);
and U2729 (N_2729,N_2494,N_2539);
and U2730 (N_2730,N_2496,N_2499);
or U2731 (N_2731,N_2500,N_2590);
or U2732 (N_2732,N_2456,N_2557);
nand U2733 (N_2733,N_2468,N_2483);
and U2734 (N_2734,N_2547,N_2499);
nand U2735 (N_2735,N_2488,N_2458);
or U2736 (N_2736,N_2450,N_2512);
nand U2737 (N_2737,N_2410,N_2465);
or U2738 (N_2738,N_2438,N_2581);
nand U2739 (N_2739,N_2460,N_2524);
nor U2740 (N_2740,N_2506,N_2539);
and U2741 (N_2741,N_2492,N_2567);
or U2742 (N_2742,N_2443,N_2592);
and U2743 (N_2743,N_2578,N_2572);
and U2744 (N_2744,N_2569,N_2517);
and U2745 (N_2745,N_2449,N_2563);
xor U2746 (N_2746,N_2593,N_2495);
nor U2747 (N_2747,N_2565,N_2409);
nand U2748 (N_2748,N_2544,N_2548);
or U2749 (N_2749,N_2428,N_2561);
or U2750 (N_2750,N_2579,N_2524);
and U2751 (N_2751,N_2456,N_2495);
nor U2752 (N_2752,N_2512,N_2511);
or U2753 (N_2753,N_2524,N_2441);
or U2754 (N_2754,N_2462,N_2520);
or U2755 (N_2755,N_2486,N_2594);
xnor U2756 (N_2756,N_2595,N_2418);
nand U2757 (N_2757,N_2553,N_2554);
nor U2758 (N_2758,N_2412,N_2449);
nand U2759 (N_2759,N_2554,N_2484);
nand U2760 (N_2760,N_2468,N_2481);
and U2761 (N_2761,N_2509,N_2488);
nand U2762 (N_2762,N_2409,N_2550);
nand U2763 (N_2763,N_2513,N_2569);
xnor U2764 (N_2764,N_2536,N_2561);
xnor U2765 (N_2765,N_2593,N_2416);
or U2766 (N_2766,N_2566,N_2500);
or U2767 (N_2767,N_2478,N_2477);
xnor U2768 (N_2768,N_2572,N_2443);
and U2769 (N_2769,N_2521,N_2543);
and U2770 (N_2770,N_2476,N_2496);
nand U2771 (N_2771,N_2458,N_2550);
and U2772 (N_2772,N_2447,N_2554);
nor U2773 (N_2773,N_2543,N_2552);
and U2774 (N_2774,N_2456,N_2523);
nand U2775 (N_2775,N_2515,N_2489);
nand U2776 (N_2776,N_2418,N_2503);
or U2777 (N_2777,N_2443,N_2543);
nor U2778 (N_2778,N_2472,N_2592);
nor U2779 (N_2779,N_2406,N_2575);
xor U2780 (N_2780,N_2579,N_2466);
or U2781 (N_2781,N_2449,N_2551);
or U2782 (N_2782,N_2512,N_2402);
or U2783 (N_2783,N_2562,N_2413);
and U2784 (N_2784,N_2542,N_2585);
or U2785 (N_2785,N_2463,N_2585);
and U2786 (N_2786,N_2509,N_2534);
or U2787 (N_2787,N_2581,N_2418);
xor U2788 (N_2788,N_2498,N_2535);
nand U2789 (N_2789,N_2487,N_2577);
nor U2790 (N_2790,N_2494,N_2533);
nand U2791 (N_2791,N_2473,N_2408);
nand U2792 (N_2792,N_2547,N_2408);
and U2793 (N_2793,N_2400,N_2598);
xnor U2794 (N_2794,N_2447,N_2558);
or U2795 (N_2795,N_2441,N_2564);
and U2796 (N_2796,N_2465,N_2435);
and U2797 (N_2797,N_2437,N_2469);
nand U2798 (N_2798,N_2459,N_2481);
and U2799 (N_2799,N_2544,N_2453);
nand U2800 (N_2800,N_2672,N_2717);
or U2801 (N_2801,N_2784,N_2758);
or U2802 (N_2802,N_2696,N_2643);
nand U2803 (N_2803,N_2644,N_2660);
or U2804 (N_2804,N_2779,N_2687);
or U2805 (N_2805,N_2738,N_2653);
and U2806 (N_2806,N_2639,N_2716);
and U2807 (N_2807,N_2685,N_2769);
or U2808 (N_2808,N_2718,N_2621);
and U2809 (N_2809,N_2782,N_2787);
and U2810 (N_2810,N_2669,N_2745);
nand U2811 (N_2811,N_2775,N_2746);
or U2812 (N_2812,N_2663,N_2720);
xnor U2813 (N_2813,N_2659,N_2665);
or U2814 (N_2814,N_2645,N_2736);
nor U2815 (N_2815,N_2712,N_2654);
and U2816 (N_2816,N_2608,N_2630);
nand U2817 (N_2817,N_2636,N_2764);
nand U2818 (N_2818,N_2774,N_2631);
nand U2819 (N_2819,N_2789,N_2722);
or U2820 (N_2820,N_2701,N_2731);
or U2821 (N_2821,N_2661,N_2703);
or U2822 (N_2822,N_2686,N_2607);
nand U2823 (N_2823,N_2725,N_2617);
and U2824 (N_2824,N_2681,N_2773);
xor U2825 (N_2825,N_2757,N_2664);
nor U2826 (N_2826,N_2756,N_2702);
nor U2827 (N_2827,N_2605,N_2750);
nand U2828 (N_2828,N_2785,N_2695);
or U2829 (N_2829,N_2698,N_2693);
nand U2830 (N_2830,N_2791,N_2708);
and U2831 (N_2831,N_2793,N_2781);
or U2832 (N_2832,N_2700,N_2740);
and U2833 (N_2833,N_2632,N_2735);
nor U2834 (N_2834,N_2622,N_2710);
nor U2835 (N_2835,N_2620,N_2715);
nor U2836 (N_2836,N_2623,N_2797);
or U2837 (N_2837,N_2799,N_2603);
nor U2838 (N_2838,N_2743,N_2626);
and U2839 (N_2839,N_2638,N_2635);
xnor U2840 (N_2840,N_2737,N_2640);
nand U2841 (N_2841,N_2615,N_2684);
nor U2842 (N_2842,N_2748,N_2786);
nand U2843 (N_2843,N_2719,N_2762);
or U2844 (N_2844,N_2678,N_2657);
or U2845 (N_2845,N_2714,N_2723);
nand U2846 (N_2846,N_2747,N_2697);
nor U2847 (N_2847,N_2616,N_2790);
nand U2848 (N_2848,N_2755,N_2763);
nor U2849 (N_2849,N_2770,N_2674);
nor U2850 (N_2850,N_2772,N_2673);
nor U2851 (N_2851,N_2609,N_2727);
and U2852 (N_2852,N_2788,N_2732);
nor U2853 (N_2853,N_2689,N_2741);
xor U2854 (N_2854,N_2724,N_2628);
or U2855 (N_2855,N_2601,N_2726);
and U2856 (N_2856,N_2767,N_2706);
nor U2857 (N_2857,N_2766,N_2744);
or U2858 (N_2858,N_2705,N_2624);
nor U2859 (N_2859,N_2625,N_2713);
nand U2860 (N_2860,N_2780,N_2670);
or U2861 (N_2861,N_2629,N_2759);
or U2862 (N_2862,N_2652,N_2651);
or U2863 (N_2863,N_2733,N_2691);
xor U2864 (N_2864,N_2768,N_2682);
nand U2865 (N_2865,N_2679,N_2649);
nand U2866 (N_2866,N_2618,N_2760);
nand U2867 (N_2867,N_2683,N_2604);
or U2868 (N_2868,N_2734,N_2613);
nor U2869 (N_2869,N_2690,N_2730);
xor U2870 (N_2870,N_2761,N_2721);
and U2871 (N_2871,N_2602,N_2619);
and U2872 (N_2872,N_2704,N_2699);
and U2873 (N_2873,N_2610,N_2749);
nor U2874 (N_2874,N_2792,N_2655);
and U2875 (N_2875,N_2798,N_2666);
nand U2876 (N_2876,N_2688,N_2667);
nand U2877 (N_2877,N_2709,N_2728);
nand U2878 (N_2878,N_2739,N_2778);
and U2879 (N_2879,N_2742,N_2776);
and U2880 (N_2880,N_2633,N_2647);
nor U2881 (N_2881,N_2648,N_2765);
or U2882 (N_2882,N_2795,N_2777);
nor U2883 (N_2883,N_2796,N_2600);
or U2884 (N_2884,N_2675,N_2680);
nand U2885 (N_2885,N_2650,N_2692);
and U2886 (N_2886,N_2729,N_2753);
nor U2887 (N_2887,N_2606,N_2694);
nor U2888 (N_2888,N_2634,N_2646);
and U2889 (N_2889,N_2658,N_2794);
and U2890 (N_2890,N_2676,N_2614);
or U2891 (N_2891,N_2637,N_2612);
and U2892 (N_2892,N_2656,N_2711);
and U2893 (N_2893,N_2668,N_2754);
and U2894 (N_2894,N_2662,N_2783);
and U2895 (N_2895,N_2677,N_2627);
nand U2896 (N_2896,N_2641,N_2752);
and U2897 (N_2897,N_2751,N_2642);
or U2898 (N_2898,N_2671,N_2611);
or U2899 (N_2899,N_2707,N_2771);
nand U2900 (N_2900,N_2619,N_2621);
nor U2901 (N_2901,N_2721,N_2666);
or U2902 (N_2902,N_2684,N_2688);
or U2903 (N_2903,N_2752,N_2657);
nand U2904 (N_2904,N_2788,N_2770);
nor U2905 (N_2905,N_2687,N_2758);
nor U2906 (N_2906,N_2635,N_2622);
or U2907 (N_2907,N_2622,N_2604);
nor U2908 (N_2908,N_2772,N_2796);
nor U2909 (N_2909,N_2718,N_2784);
and U2910 (N_2910,N_2784,N_2749);
xnor U2911 (N_2911,N_2638,N_2778);
xor U2912 (N_2912,N_2606,N_2760);
or U2913 (N_2913,N_2684,N_2648);
nor U2914 (N_2914,N_2726,N_2633);
and U2915 (N_2915,N_2684,N_2639);
and U2916 (N_2916,N_2786,N_2645);
nand U2917 (N_2917,N_2644,N_2686);
nor U2918 (N_2918,N_2699,N_2614);
or U2919 (N_2919,N_2626,N_2781);
nand U2920 (N_2920,N_2776,N_2683);
and U2921 (N_2921,N_2631,N_2630);
nand U2922 (N_2922,N_2705,N_2625);
and U2923 (N_2923,N_2797,N_2715);
or U2924 (N_2924,N_2704,N_2625);
nor U2925 (N_2925,N_2742,N_2675);
nor U2926 (N_2926,N_2690,N_2724);
and U2927 (N_2927,N_2630,N_2678);
and U2928 (N_2928,N_2666,N_2606);
and U2929 (N_2929,N_2622,N_2642);
or U2930 (N_2930,N_2715,N_2628);
xor U2931 (N_2931,N_2614,N_2733);
nor U2932 (N_2932,N_2793,N_2711);
or U2933 (N_2933,N_2779,N_2617);
nor U2934 (N_2934,N_2640,N_2748);
nand U2935 (N_2935,N_2603,N_2774);
nor U2936 (N_2936,N_2776,N_2604);
and U2937 (N_2937,N_2624,N_2764);
and U2938 (N_2938,N_2753,N_2705);
and U2939 (N_2939,N_2765,N_2628);
and U2940 (N_2940,N_2749,N_2712);
or U2941 (N_2941,N_2680,N_2630);
nand U2942 (N_2942,N_2730,N_2611);
nand U2943 (N_2943,N_2658,N_2650);
nor U2944 (N_2944,N_2793,N_2749);
and U2945 (N_2945,N_2621,N_2633);
or U2946 (N_2946,N_2708,N_2727);
and U2947 (N_2947,N_2651,N_2603);
xor U2948 (N_2948,N_2751,N_2737);
and U2949 (N_2949,N_2692,N_2666);
nor U2950 (N_2950,N_2713,N_2783);
or U2951 (N_2951,N_2793,N_2774);
and U2952 (N_2952,N_2630,N_2703);
and U2953 (N_2953,N_2638,N_2779);
and U2954 (N_2954,N_2624,N_2655);
and U2955 (N_2955,N_2603,N_2657);
or U2956 (N_2956,N_2744,N_2756);
nand U2957 (N_2957,N_2784,N_2786);
or U2958 (N_2958,N_2724,N_2625);
xnor U2959 (N_2959,N_2667,N_2781);
nor U2960 (N_2960,N_2726,N_2644);
nor U2961 (N_2961,N_2659,N_2669);
and U2962 (N_2962,N_2687,N_2721);
nor U2963 (N_2963,N_2616,N_2649);
and U2964 (N_2964,N_2643,N_2648);
nand U2965 (N_2965,N_2655,N_2667);
nor U2966 (N_2966,N_2732,N_2695);
nor U2967 (N_2967,N_2721,N_2601);
nand U2968 (N_2968,N_2671,N_2706);
or U2969 (N_2969,N_2665,N_2601);
or U2970 (N_2970,N_2658,N_2689);
nor U2971 (N_2971,N_2712,N_2617);
or U2972 (N_2972,N_2779,N_2669);
xor U2973 (N_2973,N_2729,N_2603);
xnor U2974 (N_2974,N_2756,N_2758);
or U2975 (N_2975,N_2770,N_2695);
nor U2976 (N_2976,N_2717,N_2639);
nand U2977 (N_2977,N_2603,N_2749);
nor U2978 (N_2978,N_2771,N_2666);
or U2979 (N_2979,N_2697,N_2776);
and U2980 (N_2980,N_2680,N_2627);
xnor U2981 (N_2981,N_2671,N_2703);
or U2982 (N_2982,N_2694,N_2601);
nand U2983 (N_2983,N_2799,N_2699);
xnor U2984 (N_2984,N_2630,N_2611);
or U2985 (N_2985,N_2657,N_2715);
and U2986 (N_2986,N_2698,N_2653);
nand U2987 (N_2987,N_2798,N_2671);
and U2988 (N_2988,N_2633,N_2632);
xor U2989 (N_2989,N_2620,N_2658);
or U2990 (N_2990,N_2772,N_2798);
or U2991 (N_2991,N_2667,N_2643);
or U2992 (N_2992,N_2607,N_2606);
or U2993 (N_2993,N_2633,N_2669);
and U2994 (N_2994,N_2711,N_2686);
and U2995 (N_2995,N_2745,N_2758);
xnor U2996 (N_2996,N_2739,N_2685);
xnor U2997 (N_2997,N_2621,N_2615);
nor U2998 (N_2998,N_2751,N_2710);
nor U2999 (N_2999,N_2722,N_2625);
xor U3000 (N_3000,N_2925,N_2933);
nand U3001 (N_3001,N_2802,N_2865);
nand U3002 (N_3002,N_2854,N_2955);
nor U3003 (N_3003,N_2832,N_2860);
nand U3004 (N_3004,N_2801,N_2979);
and U3005 (N_3005,N_2842,N_2971);
nand U3006 (N_3006,N_2867,N_2815);
nand U3007 (N_3007,N_2841,N_2924);
nand U3008 (N_3008,N_2911,N_2866);
and U3009 (N_3009,N_2898,N_2923);
nand U3010 (N_3010,N_2847,N_2844);
or U3011 (N_3011,N_2883,N_2972);
nor U3012 (N_3012,N_2995,N_2856);
xnor U3013 (N_3013,N_2845,N_2896);
and U3014 (N_3014,N_2849,N_2919);
nand U3015 (N_3015,N_2948,N_2855);
and U3016 (N_3016,N_2994,N_2998);
and U3017 (N_3017,N_2997,N_2853);
xor U3018 (N_3018,N_2826,N_2804);
and U3019 (N_3019,N_2917,N_2813);
and U3020 (N_3020,N_2916,N_2862);
and U3021 (N_3021,N_2873,N_2934);
nor U3022 (N_3022,N_2991,N_2819);
nor U3023 (N_3023,N_2874,N_2899);
or U3024 (N_3024,N_2870,N_2810);
nand U3025 (N_3025,N_2953,N_2989);
and U3026 (N_3026,N_2894,N_2936);
or U3027 (N_3027,N_2820,N_2928);
nand U3028 (N_3028,N_2915,N_2885);
and U3029 (N_3029,N_2980,N_2960);
and U3030 (N_3030,N_2952,N_2942);
xnor U3031 (N_3031,N_2863,N_2852);
nor U3032 (N_3032,N_2950,N_2937);
or U3033 (N_3033,N_2939,N_2803);
or U3034 (N_3034,N_2886,N_2888);
and U3035 (N_3035,N_2914,N_2846);
nor U3036 (N_3036,N_2878,N_2800);
or U3037 (N_3037,N_2941,N_2814);
nand U3038 (N_3038,N_2977,N_2811);
and U3039 (N_3039,N_2918,N_2973);
and U3040 (N_3040,N_2943,N_2929);
or U3041 (N_3041,N_2876,N_2821);
nand U3042 (N_3042,N_2869,N_2981);
nand U3043 (N_3043,N_2965,N_2946);
nor U3044 (N_3044,N_2962,N_2868);
or U3045 (N_3045,N_2812,N_2909);
nand U3046 (N_3046,N_2831,N_2959);
xor U3047 (N_3047,N_2904,N_2891);
nor U3048 (N_3048,N_2947,N_2935);
and U3049 (N_3049,N_2949,N_2910);
and U3050 (N_3050,N_2875,N_2985);
and U3051 (N_3051,N_2912,N_2978);
nand U3052 (N_3052,N_2932,N_2835);
nor U3053 (N_3053,N_2822,N_2893);
nor U3054 (N_3054,N_2903,N_2839);
nand U3055 (N_3055,N_2818,N_2990);
and U3056 (N_3056,N_2882,N_2905);
nand U3057 (N_3057,N_2806,N_2834);
nand U3058 (N_3058,N_2817,N_2881);
nand U3059 (N_3059,N_2986,N_2906);
nor U3060 (N_3060,N_2830,N_2857);
nor U3061 (N_3061,N_2851,N_2879);
nand U3062 (N_3062,N_2807,N_2922);
nand U3063 (N_3063,N_2982,N_2956);
or U3064 (N_3064,N_2858,N_2833);
nand U3065 (N_3065,N_2996,N_2824);
and U3066 (N_3066,N_2827,N_2975);
and U3067 (N_3067,N_2816,N_2970);
and U3068 (N_3068,N_2829,N_2958);
nand U3069 (N_3069,N_2974,N_2907);
or U3070 (N_3070,N_2930,N_2961);
nand U3071 (N_3071,N_2871,N_2900);
and U3072 (N_3072,N_2902,N_2945);
nand U3073 (N_3073,N_2805,N_2987);
nand U3074 (N_3074,N_2843,N_2938);
or U3075 (N_3075,N_2966,N_2964);
nor U3076 (N_3076,N_2992,N_2957);
nor U3077 (N_3077,N_2895,N_2999);
nor U3078 (N_3078,N_2809,N_2861);
or U3079 (N_3079,N_2872,N_2892);
or U3080 (N_3080,N_2954,N_2983);
nand U3081 (N_3081,N_2920,N_2823);
and U3082 (N_3082,N_2963,N_2988);
nand U3083 (N_3083,N_2940,N_2969);
or U3084 (N_3084,N_2901,N_2859);
and U3085 (N_3085,N_2836,N_2968);
or U3086 (N_3086,N_2837,N_2877);
or U3087 (N_3087,N_2828,N_2840);
or U3088 (N_3088,N_2890,N_2887);
nand U3089 (N_3089,N_2921,N_2908);
or U3090 (N_3090,N_2984,N_2808);
nand U3091 (N_3091,N_2864,N_2976);
or U3092 (N_3092,N_2848,N_2913);
nor U3093 (N_3093,N_2880,N_2931);
nand U3094 (N_3094,N_2825,N_2951);
nor U3095 (N_3095,N_2993,N_2897);
and U3096 (N_3096,N_2838,N_2927);
nor U3097 (N_3097,N_2889,N_2926);
or U3098 (N_3098,N_2884,N_2944);
or U3099 (N_3099,N_2850,N_2967);
and U3100 (N_3100,N_2889,N_2821);
nor U3101 (N_3101,N_2987,N_2969);
nand U3102 (N_3102,N_2972,N_2948);
xor U3103 (N_3103,N_2981,N_2887);
and U3104 (N_3104,N_2879,N_2964);
nand U3105 (N_3105,N_2843,N_2967);
nand U3106 (N_3106,N_2803,N_2993);
nor U3107 (N_3107,N_2983,N_2808);
xor U3108 (N_3108,N_2866,N_2811);
or U3109 (N_3109,N_2978,N_2833);
or U3110 (N_3110,N_2810,N_2922);
and U3111 (N_3111,N_2901,N_2806);
nand U3112 (N_3112,N_2928,N_2822);
nor U3113 (N_3113,N_2848,N_2872);
nand U3114 (N_3114,N_2844,N_2944);
and U3115 (N_3115,N_2841,N_2901);
nand U3116 (N_3116,N_2995,N_2808);
nor U3117 (N_3117,N_2913,N_2831);
nand U3118 (N_3118,N_2924,N_2946);
nor U3119 (N_3119,N_2869,N_2884);
nor U3120 (N_3120,N_2819,N_2960);
nor U3121 (N_3121,N_2914,N_2982);
or U3122 (N_3122,N_2994,N_2917);
nor U3123 (N_3123,N_2826,N_2824);
nand U3124 (N_3124,N_2909,N_2895);
and U3125 (N_3125,N_2833,N_2912);
and U3126 (N_3126,N_2901,N_2863);
nor U3127 (N_3127,N_2824,N_2817);
nor U3128 (N_3128,N_2912,N_2905);
nor U3129 (N_3129,N_2810,N_2937);
nor U3130 (N_3130,N_2811,N_2890);
and U3131 (N_3131,N_2985,N_2890);
nor U3132 (N_3132,N_2938,N_2824);
or U3133 (N_3133,N_2858,N_2952);
and U3134 (N_3134,N_2875,N_2818);
or U3135 (N_3135,N_2907,N_2940);
or U3136 (N_3136,N_2882,N_2849);
nor U3137 (N_3137,N_2948,N_2822);
nand U3138 (N_3138,N_2934,N_2986);
nand U3139 (N_3139,N_2967,N_2999);
or U3140 (N_3140,N_2999,N_2804);
xor U3141 (N_3141,N_2923,N_2994);
and U3142 (N_3142,N_2875,N_2934);
or U3143 (N_3143,N_2893,N_2821);
nor U3144 (N_3144,N_2978,N_2819);
nand U3145 (N_3145,N_2891,N_2874);
nor U3146 (N_3146,N_2802,N_2932);
or U3147 (N_3147,N_2986,N_2970);
or U3148 (N_3148,N_2904,N_2946);
nor U3149 (N_3149,N_2964,N_2861);
and U3150 (N_3150,N_2805,N_2912);
and U3151 (N_3151,N_2931,N_2842);
and U3152 (N_3152,N_2968,N_2989);
xor U3153 (N_3153,N_2978,N_2972);
or U3154 (N_3154,N_2874,N_2909);
or U3155 (N_3155,N_2908,N_2900);
and U3156 (N_3156,N_2971,N_2844);
nand U3157 (N_3157,N_2903,N_2961);
or U3158 (N_3158,N_2921,N_2895);
and U3159 (N_3159,N_2969,N_2839);
nand U3160 (N_3160,N_2832,N_2876);
or U3161 (N_3161,N_2807,N_2814);
nand U3162 (N_3162,N_2969,N_2902);
nor U3163 (N_3163,N_2955,N_2805);
or U3164 (N_3164,N_2919,N_2810);
nor U3165 (N_3165,N_2940,N_2967);
and U3166 (N_3166,N_2858,N_2906);
nor U3167 (N_3167,N_2910,N_2995);
or U3168 (N_3168,N_2947,N_2978);
or U3169 (N_3169,N_2892,N_2888);
nand U3170 (N_3170,N_2960,N_2904);
or U3171 (N_3171,N_2944,N_2916);
xnor U3172 (N_3172,N_2910,N_2874);
or U3173 (N_3173,N_2808,N_2828);
or U3174 (N_3174,N_2803,N_2830);
xor U3175 (N_3175,N_2939,N_2860);
and U3176 (N_3176,N_2916,N_2861);
nand U3177 (N_3177,N_2804,N_2816);
and U3178 (N_3178,N_2850,N_2969);
and U3179 (N_3179,N_2934,N_2917);
xnor U3180 (N_3180,N_2890,N_2831);
or U3181 (N_3181,N_2915,N_2861);
nand U3182 (N_3182,N_2954,N_2844);
xnor U3183 (N_3183,N_2973,N_2970);
nor U3184 (N_3184,N_2928,N_2865);
and U3185 (N_3185,N_2902,N_2865);
or U3186 (N_3186,N_2905,N_2807);
nand U3187 (N_3187,N_2976,N_2863);
or U3188 (N_3188,N_2926,N_2803);
nor U3189 (N_3189,N_2993,N_2933);
nand U3190 (N_3190,N_2915,N_2833);
or U3191 (N_3191,N_2954,N_2962);
nor U3192 (N_3192,N_2897,N_2948);
xor U3193 (N_3193,N_2916,N_2959);
or U3194 (N_3194,N_2856,N_2969);
nand U3195 (N_3195,N_2919,N_2923);
nor U3196 (N_3196,N_2946,N_2841);
and U3197 (N_3197,N_2858,N_2925);
nand U3198 (N_3198,N_2870,N_2960);
nor U3199 (N_3199,N_2920,N_2910);
nand U3200 (N_3200,N_3003,N_3196);
and U3201 (N_3201,N_3034,N_3182);
nor U3202 (N_3202,N_3134,N_3090);
nand U3203 (N_3203,N_3190,N_3096);
or U3204 (N_3204,N_3011,N_3115);
nand U3205 (N_3205,N_3168,N_3112);
nor U3206 (N_3206,N_3147,N_3002);
nand U3207 (N_3207,N_3143,N_3169);
nand U3208 (N_3208,N_3083,N_3177);
and U3209 (N_3209,N_3114,N_3105);
nand U3210 (N_3210,N_3139,N_3015);
or U3211 (N_3211,N_3189,N_3078);
or U3212 (N_3212,N_3145,N_3038);
nand U3213 (N_3213,N_3197,N_3037);
nand U3214 (N_3214,N_3031,N_3164);
xnor U3215 (N_3215,N_3146,N_3106);
and U3216 (N_3216,N_3113,N_3155);
nand U3217 (N_3217,N_3174,N_3110);
or U3218 (N_3218,N_3148,N_3180);
and U3219 (N_3219,N_3127,N_3144);
nor U3220 (N_3220,N_3033,N_3188);
or U3221 (N_3221,N_3053,N_3157);
xor U3222 (N_3222,N_3131,N_3039);
nor U3223 (N_3223,N_3087,N_3023);
nand U3224 (N_3224,N_3156,N_3032);
nor U3225 (N_3225,N_3161,N_3019);
nand U3226 (N_3226,N_3176,N_3102);
nor U3227 (N_3227,N_3108,N_3130);
nor U3228 (N_3228,N_3116,N_3064);
and U3229 (N_3229,N_3178,N_3186);
or U3230 (N_3230,N_3104,N_3021);
and U3231 (N_3231,N_3119,N_3026);
or U3232 (N_3232,N_3158,N_3073);
or U3233 (N_3233,N_3010,N_3193);
or U3234 (N_3234,N_3137,N_3062);
nand U3235 (N_3235,N_3012,N_3018);
or U3236 (N_3236,N_3035,N_3092);
nand U3237 (N_3237,N_3198,N_3159);
and U3238 (N_3238,N_3132,N_3046);
or U3239 (N_3239,N_3063,N_3141);
and U3240 (N_3240,N_3009,N_3184);
nand U3241 (N_3241,N_3027,N_3067);
nand U3242 (N_3242,N_3179,N_3101);
nand U3243 (N_3243,N_3069,N_3070);
nor U3244 (N_3244,N_3000,N_3183);
or U3245 (N_3245,N_3066,N_3122);
xor U3246 (N_3246,N_3028,N_3054);
nor U3247 (N_3247,N_3040,N_3111);
or U3248 (N_3248,N_3138,N_3151);
nor U3249 (N_3249,N_3133,N_3160);
and U3250 (N_3250,N_3042,N_3055);
or U3251 (N_3251,N_3071,N_3172);
or U3252 (N_3252,N_3136,N_3056);
and U3253 (N_3253,N_3152,N_3058);
and U3254 (N_3254,N_3098,N_3175);
or U3255 (N_3255,N_3167,N_3068);
or U3256 (N_3256,N_3191,N_3125);
or U3257 (N_3257,N_3084,N_3118);
nor U3258 (N_3258,N_3006,N_3013);
nand U3259 (N_3259,N_3005,N_3004);
nand U3260 (N_3260,N_3060,N_3135);
nor U3261 (N_3261,N_3093,N_3045);
nor U3262 (N_3262,N_3036,N_3154);
nand U3263 (N_3263,N_3029,N_3050);
or U3264 (N_3264,N_3007,N_3030);
and U3265 (N_3265,N_3162,N_3149);
nand U3266 (N_3266,N_3049,N_3059);
xnor U3267 (N_3267,N_3089,N_3014);
nand U3268 (N_3268,N_3124,N_3001);
or U3269 (N_3269,N_3048,N_3041);
nor U3270 (N_3270,N_3128,N_3079);
nor U3271 (N_3271,N_3117,N_3044);
or U3272 (N_3272,N_3082,N_3187);
and U3273 (N_3273,N_3088,N_3153);
and U3274 (N_3274,N_3150,N_3194);
and U3275 (N_3275,N_3166,N_3076);
and U3276 (N_3276,N_3181,N_3192);
nor U3277 (N_3277,N_3121,N_3140);
and U3278 (N_3278,N_3099,N_3107);
nor U3279 (N_3279,N_3047,N_3074);
xnor U3280 (N_3280,N_3095,N_3185);
nand U3281 (N_3281,N_3022,N_3016);
nand U3282 (N_3282,N_3097,N_3165);
xnor U3283 (N_3283,N_3051,N_3072);
and U3284 (N_3284,N_3052,N_3142);
nand U3285 (N_3285,N_3024,N_3123);
or U3286 (N_3286,N_3086,N_3008);
nand U3287 (N_3287,N_3020,N_3109);
and U3288 (N_3288,N_3061,N_3043);
nor U3289 (N_3289,N_3077,N_3199);
and U3290 (N_3290,N_3171,N_3103);
nor U3291 (N_3291,N_3163,N_3080);
nor U3292 (N_3292,N_3094,N_3173);
nor U3293 (N_3293,N_3170,N_3091);
xnor U3294 (N_3294,N_3081,N_3075);
nand U3295 (N_3295,N_3100,N_3120);
and U3296 (N_3296,N_3057,N_3065);
and U3297 (N_3297,N_3126,N_3017);
or U3298 (N_3298,N_3025,N_3195);
and U3299 (N_3299,N_3085,N_3129);
nor U3300 (N_3300,N_3103,N_3057);
or U3301 (N_3301,N_3114,N_3185);
nand U3302 (N_3302,N_3012,N_3083);
and U3303 (N_3303,N_3019,N_3198);
xnor U3304 (N_3304,N_3134,N_3038);
and U3305 (N_3305,N_3037,N_3172);
nand U3306 (N_3306,N_3090,N_3144);
or U3307 (N_3307,N_3170,N_3019);
nand U3308 (N_3308,N_3186,N_3014);
nor U3309 (N_3309,N_3147,N_3005);
nand U3310 (N_3310,N_3110,N_3098);
nand U3311 (N_3311,N_3067,N_3048);
xnor U3312 (N_3312,N_3190,N_3097);
xnor U3313 (N_3313,N_3075,N_3131);
and U3314 (N_3314,N_3062,N_3059);
xor U3315 (N_3315,N_3168,N_3163);
and U3316 (N_3316,N_3137,N_3127);
nand U3317 (N_3317,N_3072,N_3133);
nor U3318 (N_3318,N_3066,N_3084);
xnor U3319 (N_3319,N_3055,N_3157);
nor U3320 (N_3320,N_3007,N_3115);
or U3321 (N_3321,N_3163,N_3033);
nand U3322 (N_3322,N_3102,N_3020);
nand U3323 (N_3323,N_3056,N_3166);
nor U3324 (N_3324,N_3040,N_3051);
nor U3325 (N_3325,N_3057,N_3185);
xnor U3326 (N_3326,N_3027,N_3007);
nand U3327 (N_3327,N_3086,N_3126);
nor U3328 (N_3328,N_3020,N_3124);
nor U3329 (N_3329,N_3083,N_3106);
nor U3330 (N_3330,N_3072,N_3087);
nand U3331 (N_3331,N_3116,N_3002);
nor U3332 (N_3332,N_3103,N_3173);
or U3333 (N_3333,N_3069,N_3155);
nor U3334 (N_3334,N_3077,N_3156);
nand U3335 (N_3335,N_3007,N_3187);
or U3336 (N_3336,N_3190,N_3192);
or U3337 (N_3337,N_3080,N_3117);
and U3338 (N_3338,N_3165,N_3033);
or U3339 (N_3339,N_3100,N_3013);
and U3340 (N_3340,N_3189,N_3018);
or U3341 (N_3341,N_3035,N_3192);
nand U3342 (N_3342,N_3144,N_3107);
xnor U3343 (N_3343,N_3182,N_3050);
or U3344 (N_3344,N_3144,N_3029);
or U3345 (N_3345,N_3044,N_3183);
and U3346 (N_3346,N_3121,N_3047);
nor U3347 (N_3347,N_3114,N_3099);
and U3348 (N_3348,N_3097,N_3043);
and U3349 (N_3349,N_3179,N_3123);
nand U3350 (N_3350,N_3141,N_3076);
nor U3351 (N_3351,N_3170,N_3177);
or U3352 (N_3352,N_3056,N_3187);
and U3353 (N_3353,N_3064,N_3189);
nand U3354 (N_3354,N_3058,N_3079);
xor U3355 (N_3355,N_3116,N_3192);
nand U3356 (N_3356,N_3043,N_3171);
nand U3357 (N_3357,N_3185,N_3176);
nand U3358 (N_3358,N_3121,N_3082);
xor U3359 (N_3359,N_3178,N_3188);
nand U3360 (N_3360,N_3004,N_3163);
nand U3361 (N_3361,N_3189,N_3030);
nor U3362 (N_3362,N_3083,N_3034);
or U3363 (N_3363,N_3118,N_3137);
xor U3364 (N_3364,N_3028,N_3181);
nor U3365 (N_3365,N_3198,N_3155);
or U3366 (N_3366,N_3133,N_3069);
nor U3367 (N_3367,N_3027,N_3033);
nor U3368 (N_3368,N_3037,N_3069);
or U3369 (N_3369,N_3050,N_3140);
and U3370 (N_3370,N_3080,N_3118);
nor U3371 (N_3371,N_3159,N_3111);
and U3372 (N_3372,N_3108,N_3067);
or U3373 (N_3373,N_3005,N_3122);
nor U3374 (N_3374,N_3082,N_3000);
nor U3375 (N_3375,N_3156,N_3069);
or U3376 (N_3376,N_3115,N_3037);
xnor U3377 (N_3377,N_3068,N_3096);
or U3378 (N_3378,N_3176,N_3146);
nor U3379 (N_3379,N_3190,N_3077);
nand U3380 (N_3380,N_3131,N_3100);
or U3381 (N_3381,N_3166,N_3190);
or U3382 (N_3382,N_3108,N_3079);
and U3383 (N_3383,N_3096,N_3154);
and U3384 (N_3384,N_3185,N_3168);
or U3385 (N_3385,N_3075,N_3084);
or U3386 (N_3386,N_3142,N_3140);
and U3387 (N_3387,N_3180,N_3173);
or U3388 (N_3388,N_3038,N_3151);
nor U3389 (N_3389,N_3128,N_3087);
nor U3390 (N_3390,N_3164,N_3022);
nor U3391 (N_3391,N_3117,N_3131);
nor U3392 (N_3392,N_3106,N_3038);
and U3393 (N_3393,N_3007,N_3118);
or U3394 (N_3394,N_3060,N_3004);
and U3395 (N_3395,N_3078,N_3075);
nand U3396 (N_3396,N_3162,N_3009);
or U3397 (N_3397,N_3012,N_3073);
nor U3398 (N_3398,N_3032,N_3101);
nand U3399 (N_3399,N_3190,N_3196);
and U3400 (N_3400,N_3370,N_3289);
or U3401 (N_3401,N_3356,N_3383);
nand U3402 (N_3402,N_3363,N_3320);
nand U3403 (N_3403,N_3206,N_3303);
nor U3404 (N_3404,N_3333,N_3244);
and U3405 (N_3405,N_3253,N_3255);
nand U3406 (N_3406,N_3212,N_3390);
and U3407 (N_3407,N_3224,N_3223);
nand U3408 (N_3408,N_3220,N_3273);
nor U3409 (N_3409,N_3314,N_3272);
or U3410 (N_3410,N_3330,N_3221);
xnor U3411 (N_3411,N_3319,N_3300);
and U3412 (N_3412,N_3386,N_3232);
nor U3413 (N_3413,N_3397,N_3277);
and U3414 (N_3414,N_3276,N_3343);
xnor U3415 (N_3415,N_3338,N_3382);
and U3416 (N_3416,N_3310,N_3268);
nand U3417 (N_3417,N_3213,N_3361);
xnor U3418 (N_3418,N_3252,N_3257);
and U3419 (N_3419,N_3282,N_3215);
nor U3420 (N_3420,N_3222,N_3379);
nand U3421 (N_3421,N_3207,N_3368);
and U3422 (N_3422,N_3243,N_3324);
or U3423 (N_3423,N_3201,N_3248);
and U3424 (N_3424,N_3348,N_3375);
xnor U3425 (N_3425,N_3246,N_3335);
nor U3426 (N_3426,N_3235,N_3360);
and U3427 (N_3427,N_3312,N_3290);
nor U3428 (N_3428,N_3292,N_3306);
nor U3429 (N_3429,N_3278,N_3214);
or U3430 (N_3430,N_3279,N_3229);
and U3431 (N_3431,N_3203,N_3263);
nor U3432 (N_3432,N_3316,N_3331);
and U3433 (N_3433,N_3259,N_3353);
or U3434 (N_3434,N_3346,N_3256);
xor U3435 (N_3435,N_3226,N_3281);
nor U3436 (N_3436,N_3274,N_3369);
and U3437 (N_3437,N_3339,N_3336);
or U3438 (N_3438,N_3315,N_3205);
or U3439 (N_3439,N_3250,N_3216);
and U3440 (N_3440,N_3371,N_3291);
nand U3441 (N_3441,N_3350,N_3347);
xnor U3442 (N_3442,N_3384,N_3210);
and U3443 (N_3443,N_3261,N_3366);
nand U3444 (N_3444,N_3355,N_3247);
nand U3445 (N_3445,N_3286,N_3349);
nand U3446 (N_3446,N_3385,N_3323);
or U3447 (N_3447,N_3301,N_3307);
nand U3448 (N_3448,N_3380,N_3337);
nor U3449 (N_3449,N_3254,N_3269);
nand U3450 (N_3450,N_3251,N_3398);
and U3451 (N_3451,N_3359,N_3395);
or U3452 (N_3452,N_3234,N_3230);
nor U3453 (N_3453,N_3364,N_3321);
xnor U3454 (N_3454,N_3211,N_3245);
nand U3455 (N_3455,N_3376,N_3202);
or U3456 (N_3456,N_3313,N_3354);
and U3457 (N_3457,N_3391,N_3294);
nand U3458 (N_3458,N_3372,N_3298);
nand U3459 (N_3459,N_3242,N_3342);
nand U3460 (N_3460,N_3362,N_3352);
xnor U3461 (N_3461,N_3233,N_3288);
nor U3462 (N_3462,N_3322,N_3326);
and U3463 (N_3463,N_3317,N_3284);
and U3464 (N_3464,N_3297,N_3208);
nand U3465 (N_3465,N_3332,N_3327);
nand U3466 (N_3466,N_3365,N_3329);
and U3467 (N_3467,N_3200,N_3374);
nand U3468 (N_3468,N_3396,N_3285);
or U3469 (N_3469,N_3225,N_3236);
nand U3470 (N_3470,N_3399,N_3377);
nor U3471 (N_3471,N_3340,N_3393);
or U3472 (N_3472,N_3344,N_3328);
and U3473 (N_3473,N_3238,N_3237);
or U3474 (N_3474,N_3296,N_3325);
or U3475 (N_3475,N_3345,N_3219);
and U3476 (N_3476,N_3381,N_3308);
nand U3477 (N_3477,N_3373,N_3387);
nand U3478 (N_3478,N_3388,N_3240);
and U3479 (N_3479,N_3204,N_3258);
nand U3480 (N_3480,N_3305,N_3394);
nor U3481 (N_3481,N_3239,N_3389);
or U3482 (N_3482,N_3264,N_3241);
and U3483 (N_3483,N_3351,N_3378);
nand U3484 (N_3484,N_3283,N_3265);
or U3485 (N_3485,N_3262,N_3275);
nand U3486 (N_3486,N_3280,N_3217);
xor U3487 (N_3487,N_3299,N_3302);
nor U3488 (N_3488,N_3227,N_3266);
nand U3489 (N_3489,N_3304,N_3231);
nand U3490 (N_3490,N_3218,N_3367);
and U3491 (N_3491,N_3270,N_3357);
and U3492 (N_3492,N_3271,N_3392);
nand U3493 (N_3493,N_3341,N_3358);
nor U3494 (N_3494,N_3293,N_3311);
or U3495 (N_3495,N_3287,N_3309);
nor U3496 (N_3496,N_3209,N_3260);
nor U3497 (N_3497,N_3295,N_3228);
and U3498 (N_3498,N_3318,N_3267);
or U3499 (N_3499,N_3334,N_3249);
xor U3500 (N_3500,N_3310,N_3360);
and U3501 (N_3501,N_3206,N_3333);
nand U3502 (N_3502,N_3280,N_3216);
nor U3503 (N_3503,N_3262,N_3244);
or U3504 (N_3504,N_3326,N_3221);
and U3505 (N_3505,N_3274,N_3295);
or U3506 (N_3506,N_3303,N_3298);
and U3507 (N_3507,N_3361,N_3359);
xor U3508 (N_3508,N_3347,N_3280);
nor U3509 (N_3509,N_3238,N_3261);
nand U3510 (N_3510,N_3314,N_3282);
nor U3511 (N_3511,N_3239,N_3221);
or U3512 (N_3512,N_3257,N_3360);
xor U3513 (N_3513,N_3396,N_3397);
nand U3514 (N_3514,N_3323,N_3294);
nand U3515 (N_3515,N_3324,N_3245);
nor U3516 (N_3516,N_3262,N_3248);
and U3517 (N_3517,N_3284,N_3333);
nand U3518 (N_3518,N_3293,N_3325);
nand U3519 (N_3519,N_3201,N_3257);
nand U3520 (N_3520,N_3248,N_3376);
nand U3521 (N_3521,N_3323,N_3225);
and U3522 (N_3522,N_3234,N_3255);
and U3523 (N_3523,N_3208,N_3357);
and U3524 (N_3524,N_3372,N_3378);
nand U3525 (N_3525,N_3266,N_3262);
or U3526 (N_3526,N_3203,N_3225);
and U3527 (N_3527,N_3337,N_3331);
nor U3528 (N_3528,N_3365,N_3333);
xnor U3529 (N_3529,N_3387,N_3348);
or U3530 (N_3530,N_3323,N_3311);
nand U3531 (N_3531,N_3271,N_3248);
and U3532 (N_3532,N_3298,N_3374);
nand U3533 (N_3533,N_3336,N_3278);
nand U3534 (N_3534,N_3268,N_3234);
or U3535 (N_3535,N_3358,N_3284);
xor U3536 (N_3536,N_3384,N_3361);
nand U3537 (N_3537,N_3283,N_3319);
and U3538 (N_3538,N_3254,N_3295);
nor U3539 (N_3539,N_3253,N_3313);
nand U3540 (N_3540,N_3314,N_3214);
nand U3541 (N_3541,N_3393,N_3289);
nand U3542 (N_3542,N_3360,N_3399);
and U3543 (N_3543,N_3316,N_3348);
nor U3544 (N_3544,N_3340,N_3367);
nand U3545 (N_3545,N_3390,N_3362);
or U3546 (N_3546,N_3246,N_3233);
nor U3547 (N_3547,N_3375,N_3379);
nand U3548 (N_3548,N_3296,N_3362);
or U3549 (N_3549,N_3354,N_3343);
and U3550 (N_3550,N_3279,N_3301);
and U3551 (N_3551,N_3295,N_3379);
or U3552 (N_3552,N_3375,N_3258);
xnor U3553 (N_3553,N_3395,N_3210);
and U3554 (N_3554,N_3356,N_3317);
or U3555 (N_3555,N_3309,N_3340);
xor U3556 (N_3556,N_3266,N_3310);
nand U3557 (N_3557,N_3300,N_3223);
nand U3558 (N_3558,N_3252,N_3359);
nor U3559 (N_3559,N_3326,N_3268);
nor U3560 (N_3560,N_3281,N_3286);
or U3561 (N_3561,N_3286,N_3305);
nand U3562 (N_3562,N_3227,N_3307);
and U3563 (N_3563,N_3326,N_3335);
nand U3564 (N_3564,N_3287,N_3316);
or U3565 (N_3565,N_3266,N_3211);
or U3566 (N_3566,N_3293,N_3233);
or U3567 (N_3567,N_3248,N_3359);
and U3568 (N_3568,N_3340,N_3289);
and U3569 (N_3569,N_3239,N_3379);
xnor U3570 (N_3570,N_3206,N_3398);
and U3571 (N_3571,N_3326,N_3384);
nand U3572 (N_3572,N_3251,N_3366);
nor U3573 (N_3573,N_3290,N_3282);
nor U3574 (N_3574,N_3391,N_3216);
or U3575 (N_3575,N_3274,N_3392);
nor U3576 (N_3576,N_3395,N_3328);
nor U3577 (N_3577,N_3202,N_3200);
nor U3578 (N_3578,N_3260,N_3296);
or U3579 (N_3579,N_3213,N_3209);
or U3580 (N_3580,N_3376,N_3209);
and U3581 (N_3581,N_3317,N_3232);
nor U3582 (N_3582,N_3313,N_3209);
nor U3583 (N_3583,N_3301,N_3223);
nor U3584 (N_3584,N_3393,N_3336);
and U3585 (N_3585,N_3265,N_3375);
nor U3586 (N_3586,N_3379,N_3289);
and U3587 (N_3587,N_3262,N_3253);
nor U3588 (N_3588,N_3272,N_3383);
nand U3589 (N_3589,N_3374,N_3328);
or U3590 (N_3590,N_3327,N_3263);
nand U3591 (N_3591,N_3238,N_3387);
and U3592 (N_3592,N_3246,N_3201);
and U3593 (N_3593,N_3256,N_3323);
nand U3594 (N_3594,N_3283,N_3259);
nand U3595 (N_3595,N_3212,N_3272);
and U3596 (N_3596,N_3225,N_3220);
nor U3597 (N_3597,N_3323,N_3341);
and U3598 (N_3598,N_3278,N_3298);
and U3599 (N_3599,N_3378,N_3336);
nor U3600 (N_3600,N_3456,N_3433);
or U3601 (N_3601,N_3560,N_3599);
nor U3602 (N_3602,N_3503,N_3478);
nand U3603 (N_3603,N_3512,N_3536);
and U3604 (N_3604,N_3515,N_3448);
nand U3605 (N_3605,N_3583,N_3501);
or U3606 (N_3606,N_3442,N_3513);
and U3607 (N_3607,N_3450,N_3443);
nand U3608 (N_3608,N_3577,N_3451);
nand U3609 (N_3609,N_3493,N_3487);
and U3610 (N_3610,N_3415,N_3570);
or U3611 (N_3611,N_3529,N_3564);
or U3612 (N_3612,N_3541,N_3550);
nor U3613 (N_3613,N_3518,N_3434);
or U3614 (N_3614,N_3579,N_3403);
and U3615 (N_3615,N_3426,N_3587);
xor U3616 (N_3616,N_3559,N_3427);
nor U3617 (N_3617,N_3429,N_3548);
nor U3618 (N_3618,N_3568,N_3527);
nor U3619 (N_3619,N_3432,N_3444);
or U3620 (N_3620,N_3406,N_3455);
nor U3621 (N_3621,N_3558,N_3537);
and U3622 (N_3622,N_3467,N_3555);
nor U3623 (N_3623,N_3596,N_3428);
and U3624 (N_3624,N_3419,N_3547);
and U3625 (N_3625,N_3422,N_3410);
and U3626 (N_3626,N_3592,N_3423);
nor U3627 (N_3627,N_3561,N_3458);
nand U3628 (N_3628,N_3418,N_3499);
nor U3629 (N_3629,N_3498,N_3543);
and U3630 (N_3630,N_3469,N_3552);
nand U3631 (N_3631,N_3597,N_3580);
and U3632 (N_3632,N_3439,N_3476);
nand U3633 (N_3633,N_3496,N_3472);
or U3634 (N_3634,N_3420,N_3486);
or U3635 (N_3635,N_3471,N_3437);
or U3636 (N_3636,N_3505,N_3562);
nor U3637 (N_3637,N_3495,N_3459);
or U3638 (N_3638,N_3573,N_3538);
or U3639 (N_3639,N_3400,N_3578);
xnor U3640 (N_3640,N_3470,N_3447);
and U3641 (N_3641,N_3526,N_3530);
nand U3642 (N_3642,N_3454,N_3521);
or U3643 (N_3643,N_3474,N_3457);
or U3644 (N_3644,N_3588,N_3522);
nor U3645 (N_3645,N_3563,N_3523);
and U3646 (N_3646,N_3424,N_3404);
or U3647 (N_3647,N_3453,N_3534);
xnor U3648 (N_3648,N_3413,N_3556);
nand U3649 (N_3649,N_3449,N_3566);
nor U3650 (N_3650,N_3576,N_3462);
nand U3651 (N_3651,N_3532,N_3551);
nand U3652 (N_3652,N_3594,N_3507);
nand U3653 (N_3653,N_3531,N_3553);
or U3654 (N_3654,N_3414,N_3539);
xor U3655 (N_3655,N_3520,N_3411);
nor U3656 (N_3656,N_3409,N_3416);
or U3657 (N_3657,N_3485,N_3595);
nor U3658 (N_3658,N_3510,N_3514);
nand U3659 (N_3659,N_3464,N_3517);
xnor U3660 (N_3660,N_3502,N_3598);
and U3661 (N_3661,N_3465,N_3504);
and U3662 (N_3662,N_3585,N_3519);
nand U3663 (N_3663,N_3571,N_3492);
nand U3664 (N_3664,N_3412,N_3490);
nor U3665 (N_3665,N_3491,N_3481);
nand U3666 (N_3666,N_3509,N_3483);
and U3667 (N_3667,N_3535,N_3452);
nand U3668 (N_3668,N_3431,N_3574);
and U3669 (N_3669,N_3525,N_3544);
or U3670 (N_3670,N_3497,N_3516);
nor U3671 (N_3671,N_3401,N_3549);
and U3672 (N_3672,N_3590,N_3473);
nor U3673 (N_3673,N_3435,N_3545);
or U3674 (N_3674,N_3479,N_3572);
and U3675 (N_3675,N_3557,N_3533);
and U3676 (N_3676,N_3528,N_3506);
or U3677 (N_3677,N_3584,N_3480);
nand U3678 (N_3678,N_3475,N_3575);
nand U3679 (N_3679,N_3546,N_3445);
or U3680 (N_3680,N_3582,N_3440);
nor U3681 (N_3681,N_3489,N_3569);
and U3682 (N_3682,N_3484,N_3436);
or U3683 (N_3683,N_3511,N_3463);
nand U3684 (N_3684,N_3554,N_3494);
and U3685 (N_3685,N_3460,N_3425);
and U3686 (N_3686,N_3482,N_3488);
nand U3687 (N_3687,N_3468,N_3461);
nor U3688 (N_3688,N_3586,N_3402);
nor U3689 (N_3689,N_3430,N_3567);
nor U3690 (N_3690,N_3438,N_3407);
nand U3691 (N_3691,N_3591,N_3565);
nand U3692 (N_3692,N_3524,N_3408);
or U3693 (N_3693,N_3500,N_3593);
nor U3694 (N_3694,N_3421,N_3441);
nand U3695 (N_3695,N_3477,N_3446);
and U3696 (N_3696,N_3508,N_3581);
nand U3697 (N_3697,N_3542,N_3589);
nand U3698 (N_3698,N_3466,N_3405);
or U3699 (N_3699,N_3417,N_3540);
nand U3700 (N_3700,N_3464,N_3510);
nand U3701 (N_3701,N_3466,N_3500);
and U3702 (N_3702,N_3485,N_3480);
nand U3703 (N_3703,N_3573,N_3455);
nand U3704 (N_3704,N_3548,N_3451);
and U3705 (N_3705,N_3592,N_3556);
nand U3706 (N_3706,N_3445,N_3420);
nor U3707 (N_3707,N_3519,N_3557);
nand U3708 (N_3708,N_3433,N_3468);
nand U3709 (N_3709,N_3447,N_3433);
nand U3710 (N_3710,N_3569,N_3577);
nor U3711 (N_3711,N_3567,N_3465);
nor U3712 (N_3712,N_3446,N_3552);
or U3713 (N_3713,N_3542,N_3487);
xor U3714 (N_3714,N_3502,N_3599);
or U3715 (N_3715,N_3475,N_3434);
nor U3716 (N_3716,N_3477,N_3448);
nor U3717 (N_3717,N_3454,N_3460);
or U3718 (N_3718,N_3435,N_3405);
nor U3719 (N_3719,N_3509,N_3458);
nand U3720 (N_3720,N_3462,N_3566);
nand U3721 (N_3721,N_3486,N_3409);
and U3722 (N_3722,N_3584,N_3566);
nand U3723 (N_3723,N_3411,N_3436);
nor U3724 (N_3724,N_3521,N_3511);
and U3725 (N_3725,N_3520,N_3499);
nand U3726 (N_3726,N_3481,N_3496);
nor U3727 (N_3727,N_3439,N_3536);
nand U3728 (N_3728,N_3507,N_3417);
xor U3729 (N_3729,N_3462,N_3474);
or U3730 (N_3730,N_3497,N_3550);
and U3731 (N_3731,N_3444,N_3526);
or U3732 (N_3732,N_3447,N_3411);
or U3733 (N_3733,N_3447,N_3415);
or U3734 (N_3734,N_3464,N_3411);
nand U3735 (N_3735,N_3532,N_3574);
nand U3736 (N_3736,N_3517,N_3505);
and U3737 (N_3737,N_3419,N_3594);
or U3738 (N_3738,N_3598,N_3491);
or U3739 (N_3739,N_3432,N_3562);
xnor U3740 (N_3740,N_3575,N_3545);
or U3741 (N_3741,N_3432,N_3470);
or U3742 (N_3742,N_3593,N_3403);
and U3743 (N_3743,N_3434,N_3436);
nand U3744 (N_3744,N_3469,N_3476);
nor U3745 (N_3745,N_3544,N_3510);
nor U3746 (N_3746,N_3449,N_3573);
xnor U3747 (N_3747,N_3500,N_3568);
and U3748 (N_3748,N_3494,N_3415);
and U3749 (N_3749,N_3440,N_3480);
nor U3750 (N_3750,N_3485,N_3557);
nor U3751 (N_3751,N_3499,N_3468);
xor U3752 (N_3752,N_3466,N_3593);
nand U3753 (N_3753,N_3571,N_3594);
nand U3754 (N_3754,N_3551,N_3445);
or U3755 (N_3755,N_3467,N_3568);
or U3756 (N_3756,N_3444,N_3561);
nand U3757 (N_3757,N_3488,N_3424);
or U3758 (N_3758,N_3423,N_3405);
nand U3759 (N_3759,N_3537,N_3420);
or U3760 (N_3760,N_3551,N_3472);
and U3761 (N_3761,N_3542,N_3534);
or U3762 (N_3762,N_3472,N_3412);
or U3763 (N_3763,N_3459,N_3546);
nand U3764 (N_3764,N_3575,N_3435);
nand U3765 (N_3765,N_3449,N_3539);
or U3766 (N_3766,N_3482,N_3567);
nor U3767 (N_3767,N_3452,N_3449);
nor U3768 (N_3768,N_3498,N_3522);
nor U3769 (N_3769,N_3469,N_3462);
nor U3770 (N_3770,N_3585,N_3529);
nand U3771 (N_3771,N_3406,N_3526);
xnor U3772 (N_3772,N_3425,N_3555);
or U3773 (N_3773,N_3554,N_3470);
or U3774 (N_3774,N_3546,N_3482);
nor U3775 (N_3775,N_3594,N_3514);
or U3776 (N_3776,N_3521,N_3481);
nand U3777 (N_3777,N_3422,N_3500);
and U3778 (N_3778,N_3403,N_3526);
and U3779 (N_3779,N_3520,N_3594);
nor U3780 (N_3780,N_3582,N_3598);
nand U3781 (N_3781,N_3424,N_3538);
and U3782 (N_3782,N_3477,N_3505);
or U3783 (N_3783,N_3530,N_3403);
nor U3784 (N_3784,N_3477,N_3474);
xor U3785 (N_3785,N_3422,N_3434);
or U3786 (N_3786,N_3546,N_3553);
nand U3787 (N_3787,N_3506,N_3559);
nand U3788 (N_3788,N_3555,N_3514);
nand U3789 (N_3789,N_3440,N_3552);
nor U3790 (N_3790,N_3596,N_3442);
nor U3791 (N_3791,N_3469,N_3598);
nor U3792 (N_3792,N_3473,N_3475);
nand U3793 (N_3793,N_3448,N_3463);
or U3794 (N_3794,N_3592,N_3470);
and U3795 (N_3795,N_3432,N_3408);
and U3796 (N_3796,N_3425,N_3482);
or U3797 (N_3797,N_3582,N_3523);
or U3798 (N_3798,N_3581,N_3599);
nor U3799 (N_3799,N_3405,N_3551);
or U3800 (N_3800,N_3742,N_3697);
nand U3801 (N_3801,N_3698,N_3774);
nor U3802 (N_3802,N_3750,N_3761);
or U3803 (N_3803,N_3605,N_3777);
nand U3804 (N_3804,N_3704,N_3794);
nor U3805 (N_3805,N_3642,N_3636);
and U3806 (N_3806,N_3647,N_3641);
or U3807 (N_3807,N_3771,N_3616);
and U3808 (N_3808,N_3671,N_3705);
and U3809 (N_3809,N_3633,N_3722);
and U3810 (N_3810,N_3619,N_3734);
nor U3811 (N_3811,N_3791,N_3747);
and U3812 (N_3812,N_3779,N_3731);
nand U3813 (N_3813,N_3737,N_3726);
nand U3814 (N_3814,N_3686,N_3606);
or U3815 (N_3815,N_3707,N_3732);
nor U3816 (N_3816,N_3646,N_3765);
or U3817 (N_3817,N_3643,N_3720);
or U3818 (N_3818,N_3645,N_3603);
or U3819 (N_3819,N_3628,N_3743);
and U3820 (N_3820,N_3692,N_3700);
xor U3821 (N_3821,N_3738,N_3718);
nor U3822 (N_3822,N_3710,N_3673);
nor U3823 (N_3823,N_3607,N_3650);
xnor U3824 (N_3824,N_3795,N_3683);
xnor U3825 (N_3825,N_3667,N_3712);
xor U3826 (N_3826,N_3784,N_3759);
nand U3827 (N_3827,N_3781,N_3776);
nand U3828 (N_3828,N_3680,N_3789);
nand U3829 (N_3829,N_3741,N_3608);
xor U3830 (N_3830,N_3798,N_3662);
or U3831 (N_3831,N_3681,N_3689);
or U3832 (N_3832,N_3748,N_3757);
and U3833 (N_3833,N_3649,N_3660);
or U3834 (N_3834,N_3752,N_3758);
and U3835 (N_3835,N_3753,N_3792);
nor U3836 (N_3836,N_3713,N_3620);
and U3837 (N_3837,N_3639,N_3631);
nor U3838 (N_3838,N_3688,N_3621);
xor U3839 (N_3839,N_3602,N_3721);
nor U3840 (N_3840,N_3701,N_3653);
nand U3841 (N_3841,N_3699,N_3624);
xnor U3842 (N_3842,N_3727,N_3678);
xnor U3843 (N_3843,N_3644,N_3687);
or U3844 (N_3844,N_3625,N_3638);
nand U3845 (N_3845,N_3714,N_3724);
nand U3846 (N_3846,N_3661,N_3780);
and U3847 (N_3847,N_3622,N_3790);
xor U3848 (N_3848,N_3610,N_3708);
nor U3849 (N_3849,N_3627,N_3711);
nand U3850 (N_3850,N_3611,N_3767);
nor U3851 (N_3851,N_3796,N_3666);
nand U3852 (N_3852,N_3773,N_3764);
nand U3853 (N_3853,N_3614,N_3623);
nor U3854 (N_3854,N_3648,N_3664);
nand U3855 (N_3855,N_3755,N_3740);
or U3856 (N_3856,N_3723,N_3655);
nand U3857 (N_3857,N_3744,N_3702);
nor U3858 (N_3858,N_3685,N_3768);
or U3859 (N_3859,N_3637,N_3677);
nor U3860 (N_3860,N_3690,N_3772);
and U3861 (N_3861,N_3668,N_3729);
nand U3862 (N_3862,N_3733,N_3600);
or U3863 (N_3863,N_3735,N_3775);
or U3864 (N_3864,N_3665,N_3736);
xnor U3865 (N_3865,N_3770,N_3635);
nor U3866 (N_3866,N_3651,N_3659);
nor U3867 (N_3867,N_3691,N_3760);
or U3868 (N_3868,N_3703,N_3717);
nand U3869 (N_3869,N_3745,N_3751);
and U3870 (N_3870,N_3684,N_3763);
nand U3871 (N_3871,N_3601,N_3618);
and U3872 (N_3872,N_3769,N_3694);
and U3873 (N_3873,N_3615,N_3675);
or U3874 (N_3874,N_3739,N_3785);
nor U3875 (N_3875,N_3746,N_3787);
or U3876 (N_3876,N_3682,N_3762);
and U3877 (N_3877,N_3630,N_3658);
or U3878 (N_3878,N_3696,N_3799);
and U3879 (N_3879,N_3797,N_3719);
nand U3880 (N_3880,N_3695,N_3728);
nor U3881 (N_3881,N_3730,N_3766);
and U3882 (N_3882,N_3632,N_3626);
nand U3883 (N_3883,N_3749,N_3634);
and U3884 (N_3884,N_3715,N_3674);
xor U3885 (N_3885,N_3693,N_3788);
or U3886 (N_3886,N_3640,N_3676);
nand U3887 (N_3887,N_3672,N_3756);
nand U3888 (N_3888,N_3778,N_3783);
xor U3889 (N_3889,N_3706,N_3617);
or U3890 (N_3890,N_3657,N_3604);
nand U3891 (N_3891,N_3679,N_3613);
and U3892 (N_3892,N_3609,N_3716);
or U3893 (N_3893,N_3670,N_3612);
or U3894 (N_3894,N_3793,N_3652);
or U3895 (N_3895,N_3754,N_3654);
and U3896 (N_3896,N_3725,N_3786);
and U3897 (N_3897,N_3629,N_3709);
nand U3898 (N_3898,N_3782,N_3656);
nand U3899 (N_3899,N_3663,N_3669);
nand U3900 (N_3900,N_3709,N_3645);
and U3901 (N_3901,N_3758,N_3613);
nor U3902 (N_3902,N_3666,N_3702);
xnor U3903 (N_3903,N_3695,N_3673);
and U3904 (N_3904,N_3776,N_3675);
and U3905 (N_3905,N_3634,N_3624);
and U3906 (N_3906,N_3669,N_3702);
and U3907 (N_3907,N_3721,N_3710);
nor U3908 (N_3908,N_3640,N_3691);
xor U3909 (N_3909,N_3612,N_3707);
or U3910 (N_3910,N_3788,N_3638);
nand U3911 (N_3911,N_3697,N_3798);
nor U3912 (N_3912,N_3663,N_3751);
and U3913 (N_3913,N_3726,N_3702);
and U3914 (N_3914,N_3788,N_3609);
or U3915 (N_3915,N_3643,N_3633);
nand U3916 (N_3916,N_3776,N_3626);
or U3917 (N_3917,N_3743,N_3754);
and U3918 (N_3918,N_3651,N_3674);
and U3919 (N_3919,N_3626,N_3634);
xor U3920 (N_3920,N_3689,N_3697);
nand U3921 (N_3921,N_3737,N_3723);
and U3922 (N_3922,N_3734,N_3724);
nor U3923 (N_3923,N_3605,N_3713);
and U3924 (N_3924,N_3619,N_3713);
nand U3925 (N_3925,N_3621,N_3713);
and U3926 (N_3926,N_3619,N_3636);
nand U3927 (N_3927,N_3767,N_3746);
xor U3928 (N_3928,N_3621,N_3774);
nand U3929 (N_3929,N_3602,N_3769);
or U3930 (N_3930,N_3668,N_3606);
or U3931 (N_3931,N_3686,N_3677);
nor U3932 (N_3932,N_3793,N_3677);
xor U3933 (N_3933,N_3638,N_3661);
nand U3934 (N_3934,N_3706,N_3791);
nor U3935 (N_3935,N_3638,N_3647);
nor U3936 (N_3936,N_3618,N_3672);
nor U3937 (N_3937,N_3722,N_3685);
nor U3938 (N_3938,N_3763,N_3709);
and U3939 (N_3939,N_3633,N_3701);
or U3940 (N_3940,N_3674,N_3664);
and U3941 (N_3941,N_3649,N_3641);
xor U3942 (N_3942,N_3748,N_3793);
nand U3943 (N_3943,N_3710,N_3645);
or U3944 (N_3944,N_3635,N_3659);
or U3945 (N_3945,N_3619,N_3609);
xor U3946 (N_3946,N_3716,N_3758);
or U3947 (N_3947,N_3614,N_3769);
or U3948 (N_3948,N_3605,N_3797);
nor U3949 (N_3949,N_3708,N_3629);
nor U3950 (N_3950,N_3748,N_3702);
nor U3951 (N_3951,N_3617,N_3753);
nor U3952 (N_3952,N_3700,N_3704);
nor U3953 (N_3953,N_3613,N_3602);
nor U3954 (N_3954,N_3777,N_3701);
nor U3955 (N_3955,N_3619,N_3632);
or U3956 (N_3956,N_3700,N_3787);
or U3957 (N_3957,N_3651,N_3708);
nand U3958 (N_3958,N_3619,N_3631);
nand U3959 (N_3959,N_3737,N_3667);
or U3960 (N_3960,N_3621,N_3639);
or U3961 (N_3961,N_3655,N_3767);
and U3962 (N_3962,N_3741,N_3612);
nor U3963 (N_3963,N_3696,N_3665);
or U3964 (N_3964,N_3664,N_3750);
nor U3965 (N_3965,N_3683,N_3671);
and U3966 (N_3966,N_3772,N_3791);
nor U3967 (N_3967,N_3766,N_3756);
nor U3968 (N_3968,N_3642,N_3755);
xnor U3969 (N_3969,N_3749,N_3671);
nor U3970 (N_3970,N_3620,N_3712);
nor U3971 (N_3971,N_3744,N_3755);
xor U3972 (N_3972,N_3788,N_3738);
and U3973 (N_3973,N_3689,N_3739);
nor U3974 (N_3974,N_3743,N_3770);
or U3975 (N_3975,N_3666,N_3618);
xnor U3976 (N_3976,N_3670,N_3641);
nor U3977 (N_3977,N_3603,N_3799);
nor U3978 (N_3978,N_3733,N_3646);
nor U3979 (N_3979,N_3791,N_3744);
nand U3980 (N_3980,N_3664,N_3716);
nand U3981 (N_3981,N_3657,N_3739);
nor U3982 (N_3982,N_3638,N_3797);
and U3983 (N_3983,N_3655,N_3783);
xor U3984 (N_3984,N_3786,N_3674);
and U3985 (N_3985,N_3659,N_3750);
nor U3986 (N_3986,N_3672,N_3611);
or U3987 (N_3987,N_3733,N_3679);
or U3988 (N_3988,N_3674,N_3788);
nand U3989 (N_3989,N_3654,N_3616);
nand U3990 (N_3990,N_3634,N_3701);
xnor U3991 (N_3991,N_3648,N_3630);
nor U3992 (N_3992,N_3742,N_3684);
nand U3993 (N_3993,N_3684,N_3746);
nor U3994 (N_3994,N_3748,N_3615);
nand U3995 (N_3995,N_3639,N_3756);
nand U3996 (N_3996,N_3632,N_3782);
nor U3997 (N_3997,N_3601,N_3644);
and U3998 (N_3998,N_3750,N_3771);
and U3999 (N_3999,N_3683,N_3698);
and U4000 (N_4000,N_3926,N_3971);
nand U4001 (N_4001,N_3851,N_3915);
and U4002 (N_4002,N_3939,N_3948);
nor U4003 (N_4003,N_3815,N_3959);
or U4004 (N_4004,N_3991,N_3924);
nor U4005 (N_4005,N_3841,N_3917);
nand U4006 (N_4006,N_3896,N_3942);
xnor U4007 (N_4007,N_3902,N_3923);
nor U4008 (N_4008,N_3919,N_3979);
nor U4009 (N_4009,N_3817,N_3863);
or U4010 (N_4010,N_3944,N_3989);
nor U4011 (N_4011,N_3850,N_3848);
and U4012 (N_4012,N_3930,N_3897);
nor U4013 (N_4013,N_3862,N_3999);
nor U4014 (N_4014,N_3810,N_3895);
xor U4015 (N_4015,N_3808,N_3833);
xnor U4016 (N_4016,N_3985,N_3866);
nand U4017 (N_4017,N_3882,N_3888);
or U4018 (N_4018,N_3945,N_3908);
or U4019 (N_4019,N_3837,N_3828);
and U4020 (N_4020,N_3932,N_3824);
nor U4021 (N_4021,N_3952,N_3860);
or U4022 (N_4022,N_3843,N_3921);
nand U4023 (N_4023,N_3885,N_3954);
nand U4024 (N_4024,N_3890,N_3823);
nor U4025 (N_4025,N_3835,N_3803);
nand U4026 (N_4026,N_3990,N_3820);
xor U4027 (N_4027,N_3859,N_3880);
and U4028 (N_4028,N_3879,N_3849);
and U4029 (N_4029,N_3805,N_3997);
nand U4030 (N_4030,N_3854,N_3929);
or U4031 (N_4031,N_3978,N_3918);
nor U4032 (N_4032,N_3844,N_3906);
xor U4033 (N_4033,N_3898,N_3927);
or U4034 (N_4034,N_3904,N_3818);
xnor U4035 (N_4035,N_3911,N_3840);
or U4036 (N_4036,N_3894,N_3813);
and U4037 (N_4037,N_3925,N_3940);
nand U4038 (N_4038,N_3861,N_3819);
nor U4039 (N_4039,N_3941,N_3877);
nand U4040 (N_4040,N_3827,N_3903);
or U4041 (N_4041,N_3907,N_3961);
and U4042 (N_4042,N_3936,N_3874);
xnor U4043 (N_4043,N_3992,N_3893);
and U4044 (N_4044,N_3957,N_3869);
nor U4045 (N_4045,N_3905,N_3809);
and U4046 (N_4046,N_3868,N_3900);
nor U4047 (N_4047,N_3949,N_3871);
xor U4048 (N_4048,N_3881,N_3857);
xor U4049 (N_4049,N_3987,N_3964);
nand U4050 (N_4050,N_3928,N_3858);
or U4051 (N_4051,N_3825,N_3811);
and U4052 (N_4052,N_3807,N_3922);
nand U4053 (N_4053,N_3878,N_3847);
or U4054 (N_4054,N_3812,N_3867);
or U4055 (N_4055,N_3875,N_3913);
nand U4056 (N_4056,N_3883,N_3886);
xnor U4057 (N_4057,N_3995,N_3855);
nand U4058 (N_4058,N_3884,N_3801);
xnor U4059 (N_4059,N_3994,N_3912);
nor U4060 (N_4060,N_3901,N_3951);
or U4061 (N_4061,N_3933,N_3977);
and U4062 (N_4062,N_3996,N_3832);
and U4063 (N_4063,N_3829,N_3943);
or U4064 (N_4064,N_3910,N_3983);
or U4065 (N_4065,N_3947,N_3974);
xor U4066 (N_4066,N_3950,N_3988);
nor U4067 (N_4067,N_3962,N_3852);
and U4068 (N_4068,N_3986,N_3980);
xnor U4069 (N_4069,N_3821,N_3814);
nand U4070 (N_4070,N_3842,N_3975);
or U4071 (N_4071,N_3804,N_3953);
nor U4072 (N_4072,N_3845,N_3838);
nor U4073 (N_4073,N_3806,N_3856);
nor U4074 (N_4074,N_3984,N_3876);
nand U4075 (N_4075,N_3937,N_3998);
nor U4076 (N_4076,N_3931,N_3872);
xnor U4077 (N_4077,N_3920,N_3899);
and U4078 (N_4078,N_3960,N_3834);
nand U4079 (N_4079,N_3969,N_3967);
nor U4080 (N_4080,N_3968,N_3830);
nor U4081 (N_4081,N_3836,N_3909);
and U4082 (N_4082,N_3955,N_3800);
nor U4083 (N_4083,N_3831,N_3914);
nor U4084 (N_4084,N_3935,N_3802);
nor U4085 (N_4085,N_3853,N_3873);
nor U4086 (N_4086,N_3839,N_3822);
or U4087 (N_4087,N_3958,N_3946);
nor U4088 (N_4088,N_3965,N_3816);
nor U4089 (N_4089,N_3956,N_3870);
and U4090 (N_4090,N_3993,N_3982);
nor U4091 (N_4091,N_3973,N_3889);
xor U4092 (N_4092,N_3966,N_3976);
xnor U4093 (N_4093,N_3963,N_3887);
nor U4094 (N_4094,N_3981,N_3865);
nor U4095 (N_4095,N_3916,N_3891);
nor U4096 (N_4096,N_3826,N_3972);
nor U4097 (N_4097,N_3846,N_3970);
nand U4098 (N_4098,N_3938,N_3892);
and U4099 (N_4099,N_3864,N_3934);
nor U4100 (N_4100,N_3913,N_3869);
nand U4101 (N_4101,N_3922,N_3913);
and U4102 (N_4102,N_3801,N_3842);
or U4103 (N_4103,N_3851,N_3821);
or U4104 (N_4104,N_3873,N_3836);
or U4105 (N_4105,N_3841,N_3851);
or U4106 (N_4106,N_3911,N_3875);
nand U4107 (N_4107,N_3978,N_3939);
xor U4108 (N_4108,N_3964,N_3919);
nor U4109 (N_4109,N_3897,N_3999);
and U4110 (N_4110,N_3941,N_3900);
or U4111 (N_4111,N_3814,N_3950);
xnor U4112 (N_4112,N_3953,N_3955);
nor U4113 (N_4113,N_3852,N_3971);
nand U4114 (N_4114,N_3961,N_3893);
xnor U4115 (N_4115,N_3953,N_3990);
nor U4116 (N_4116,N_3934,N_3985);
and U4117 (N_4117,N_3824,N_3885);
nand U4118 (N_4118,N_3999,N_3958);
or U4119 (N_4119,N_3973,N_3869);
and U4120 (N_4120,N_3838,N_3828);
nor U4121 (N_4121,N_3941,N_3873);
nand U4122 (N_4122,N_3905,N_3858);
or U4123 (N_4123,N_3980,N_3812);
nand U4124 (N_4124,N_3976,N_3855);
or U4125 (N_4125,N_3848,N_3970);
and U4126 (N_4126,N_3857,N_3924);
nor U4127 (N_4127,N_3929,N_3811);
xor U4128 (N_4128,N_3828,N_3884);
and U4129 (N_4129,N_3885,N_3864);
nand U4130 (N_4130,N_3970,N_3968);
or U4131 (N_4131,N_3902,N_3917);
and U4132 (N_4132,N_3875,N_3943);
and U4133 (N_4133,N_3848,N_3872);
nand U4134 (N_4134,N_3892,N_3880);
nor U4135 (N_4135,N_3925,N_3882);
or U4136 (N_4136,N_3919,N_3946);
nand U4137 (N_4137,N_3896,N_3880);
or U4138 (N_4138,N_3999,N_3933);
or U4139 (N_4139,N_3933,N_3961);
and U4140 (N_4140,N_3907,N_3934);
and U4141 (N_4141,N_3951,N_3964);
or U4142 (N_4142,N_3976,N_3804);
nand U4143 (N_4143,N_3972,N_3921);
nor U4144 (N_4144,N_3865,N_3898);
nor U4145 (N_4145,N_3823,N_3889);
and U4146 (N_4146,N_3869,N_3940);
or U4147 (N_4147,N_3869,N_3854);
and U4148 (N_4148,N_3978,N_3819);
xor U4149 (N_4149,N_3926,N_3882);
and U4150 (N_4150,N_3942,N_3955);
nand U4151 (N_4151,N_3859,N_3820);
nand U4152 (N_4152,N_3960,N_3945);
nor U4153 (N_4153,N_3805,N_3928);
or U4154 (N_4154,N_3851,N_3920);
nand U4155 (N_4155,N_3895,N_3893);
and U4156 (N_4156,N_3816,N_3970);
nor U4157 (N_4157,N_3834,N_3963);
or U4158 (N_4158,N_3824,N_3827);
and U4159 (N_4159,N_3987,N_3984);
nor U4160 (N_4160,N_3895,N_3872);
nand U4161 (N_4161,N_3935,N_3856);
and U4162 (N_4162,N_3878,N_3960);
nand U4163 (N_4163,N_3993,N_3912);
nor U4164 (N_4164,N_3906,N_3890);
and U4165 (N_4165,N_3888,N_3808);
xor U4166 (N_4166,N_3898,N_3802);
or U4167 (N_4167,N_3894,N_3860);
or U4168 (N_4168,N_3894,N_3871);
xnor U4169 (N_4169,N_3927,N_3880);
xnor U4170 (N_4170,N_3824,N_3843);
and U4171 (N_4171,N_3990,N_3950);
and U4172 (N_4172,N_3866,N_3970);
xor U4173 (N_4173,N_3982,N_3964);
and U4174 (N_4174,N_3838,N_3950);
nand U4175 (N_4175,N_3929,N_3850);
and U4176 (N_4176,N_3970,N_3987);
nor U4177 (N_4177,N_3993,N_3849);
nor U4178 (N_4178,N_3890,N_3944);
nand U4179 (N_4179,N_3987,N_3898);
and U4180 (N_4180,N_3937,N_3873);
nor U4181 (N_4181,N_3817,N_3824);
and U4182 (N_4182,N_3998,N_3904);
nand U4183 (N_4183,N_3995,N_3944);
and U4184 (N_4184,N_3939,N_3901);
nor U4185 (N_4185,N_3948,N_3968);
or U4186 (N_4186,N_3804,N_3901);
or U4187 (N_4187,N_3990,N_3943);
or U4188 (N_4188,N_3917,N_3819);
nor U4189 (N_4189,N_3885,N_3818);
and U4190 (N_4190,N_3897,N_3889);
or U4191 (N_4191,N_3852,N_3964);
or U4192 (N_4192,N_3825,N_3960);
and U4193 (N_4193,N_3906,N_3840);
or U4194 (N_4194,N_3993,N_3881);
and U4195 (N_4195,N_3865,N_3905);
nor U4196 (N_4196,N_3836,N_3996);
nand U4197 (N_4197,N_3877,N_3910);
nand U4198 (N_4198,N_3800,N_3839);
nor U4199 (N_4199,N_3855,N_3879);
and U4200 (N_4200,N_4181,N_4001);
xnor U4201 (N_4201,N_4092,N_4199);
and U4202 (N_4202,N_4071,N_4008);
nand U4203 (N_4203,N_4162,N_4119);
or U4204 (N_4204,N_4152,N_4195);
nor U4205 (N_4205,N_4073,N_4190);
or U4206 (N_4206,N_4034,N_4045);
and U4207 (N_4207,N_4136,N_4128);
and U4208 (N_4208,N_4068,N_4109);
or U4209 (N_4209,N_4060,N_4041);
nand U4210 (N_4210,N_4196,N_4006);
nor U4211 (N_4211,N_4043,N_4171);
and U4212 (N_4212,N_4053,N_4035);
nand U4213 (N_4213,N_4106,N_4098);
xor U4214 (N_4214,N_4062,N_4135);
or U4215 (N_4215,N_4069,N_4024);
nand U4216 (N_4216,N_4064,N_4016);
and U4217 (N_4217,N_4077,N_4058);
nor U4218 (N_4218,N_4185,N_4148);
nor U4219 (N_4219,N_4193,N_4030);
or U4220 (N_4220,N_4099,N_4141);
nor U4221 (N_4221,N_4054,N_4063);
nand U4222 (N_4222,N_4102,N_4118);
and U4223 (N_4223,N_4149,N_4015);
and U4224 (N_4224,N_4161,N_4114);
nor U4225 (N_4225,N_4066,N_4065);
or U4226 (N_4226,N_4166,N_4010);
nand U4227 (N_4227,N_4172,N_4078);
nor U4228 (N_4228,N_4103,N_4165);
nor U4229 (N_4229,N_4182,N_4127);
nor U4230 (N_4230,N_4133,N_4187);
and U4231 (N_4231,N_4059,N_4189);
nand U4232 (N_4232,N_4082,N_4140);
nor U4233 (N_4233,N_4186,N_4178);
and U4234 (N_4234,N_4017,N_4188);
and U4235 (N_4235,N_4067,N_4120);
nor U4236 (N_4236,N_4115,N_4046);
or U4237 (N_4237,N_4179,N_4101);
nor U4238 (N_4238,N_4139,N_4080);
and U4239 (N_4239,N_4021,N_4154);
nor U4240 (N_4240,N_4123,N_4143);
xor U4241 (N_4241,N_4198,N_4033);
and U4242 (N_4242,N_4048,N_4096);
nor U4243 (N_4243,N_4153,N_4144);
and U4244 (N_4244,N_4158,N_4022);
nor U4245 (N_4245,N_4192,N_4012);
and U4246 (N_4246,N_4029,N_4091);
xnor U4247 (N_4247,N_4094,N_4197);
xor U4248 (N_4248,N_4047,N_4163);
nand U4249 (N_4249,N_4168,N_4124);
and U4250 (N_4250,N_4121,N_4151);
nand U4251 (N_4251,N_4174,N_4145);
and U4252 (N_4252,N_4079,N_4037);
nand U4253 (N_4253,N_4134,N_4072);
nand U4254 (N_4254,N_4105,N_4052);
nand U4255 (N_4255,N_4100,N_4084);
or U4256 (N_4256,N_4019,N_4027);
and U4257 (N_4257,N_4057,N_4049);
and U4258 (N_4258,N_4113,N_4089);
or U4259 (N_4259,N_4093,N_4129);
and U4260 (N_4260,N_4110,N_4005);
and U4261 (N_4261,N_4117,N_4173);
and U4262 (N_4262,N_4097,N_4194);
nor U4263 (N_4263,N_4146,N_4050);
nor U4264 (N_4264,N_4164,N_4122);
xnor U4265 (N_4265,N_4061,N_4074);
nor U4266 (N_4266,N_4177,N_4051);
and U4267 (N_4267,N_4112,N_4031);
and U4268 (N_4268,N_4026,N_4036);
or U4269 (N_4269,N_4023,N_4085);
nand U4270 (N_4270,N_4137,N_4018);
nand U4271 (N_4271,N_4056,N_4183);
xor U4272 (N_4272,N_4087,N_4160);
or U4273 (N_4273,N_4108,N_4116);
and U4274 (N_4274,N_4000,N_4075);
xnor U4275 (N_4275,N_4167,N_4175);
or U4276 (N_4276,N_4011,N_4009);
or U4277 (N_4277,N_4138,N_4104);
nand U4278 (N_4278,N_4028,N_4020);
nor U4279 (N_4279,N_4088,N_4111);
and U4280 (N_4280,N_4142,N_4147);
or U4281 (N_4281,N_4076,N_4157);
and U4282 (N_4282,N_4083,N_4032);
nor U4283 (N_4283,N_4130,N_4014);
and U4284 (N_4284,N_4044,N_4191);
nand U4285 (N_4285,N_4180,N_4040);
xnor U4286 (N_4286,N_4013,N_4126);
or U4287 (N_4287,N_4055,N_4070);
xnor U4288 (N_4288,N_4184,N_4176);
or U4289 (N_4289,N_4007,N_4004);
xnor U4290 (N_4290,N_4156,N_4159);
and U4291 (N_4291,N_4170,N_4038);
nand U4292 (N_4292,N_4125,N_4107);
and U4293 (N_4293,N_4095,N_4042);
and U4294 (N_4294,N_4081,N_4086);
xor U4295 (N_4295,N_4155,N_4090);
or U4296 (N_4296,N_4002,N_4003);
nor U4297 (N_4297,N_4131,N_4132);
xor U4298 (N_4298,N_4150,N_4039);
nor U4299 (N_4299,N_4169,N_4025);
nand U4300 (N_4300,N_4043,N_4130);
and U4301 (N_4301,N_4167,N_4168);
nor U4302 (N_4302,N_4103,N_4104);
or U4303 (N_4303,N_4106,N_4096);
nor U4304 (N_4304,N_4106,N_4149);
nor U4305 (N_4305,N_4198,N_4009);
xor U4306 (N_4306,N_4175,N_4196);
and U4307 (N_4307,N_4045,N_4174);
and U4308 (N_4308,N_4041,N_4012);
nor U4309 (N_4309,N_4120,N_4108);
or U4310 (N_4310,N_4110,N_4007);
and U4311 (N_4311,N_4040,N_4128);
and U4312 (N_4312,N_4198,N_4064);
xnor U4313 (N_4313,N_4106,N_4145);
or U4314 (N_4314,N_4140,N_4191);
and U4315 (N_4315,N_4162,N_4071);
nor U4316 (N_4316,N_4023,N_4143);
nor U4317 (N_4317,N_4098,N_4093);
nor U4318 (N_4318,N_4160,N_4028);
xor U4319 (N_4319,N_4026,N_4092);
nand U4320 (N_4320,N_4123,N_4004);
and U4321 (N_4321,N_4048,N_4153);
or U4322 (N_4322,N_4049,N_4193);
nand U4323 (N_4323,N_4013,N_4122);
nor U4324 (N_4324,N_4187,N_4051);
or U4325 (N_4325,N_4143,N_4073);
or U4326 (N_4326,N_4156,N_4054);
nand U4327 (N_4327,N_4153,N_4046);
and U4328 (N_4328,N_4054,N_4144);
and U4329 (N_4329,N_4000,N_4001);
and U4330 (N_4330,N_4069,N_4035);
nor U4331 (N_4331,N_4131,N_4030);
nor U4332 (N_4332,N_4054,N_4060);
and U4333 (N_4333,N_4039,N_4184);
nand U4334 (N_4334,N_4194,N_4018);
nand U4335 (N_4335,N_4103,N_4096);
or U4336 (N_4336,N_4151,N_4186);
or U4337 (N_4337,N_4189,N_4179);
nand U4338 (N_4338,N_4099,N_4077);
nand U4339 (N_4339,N_4022,N_4159);
nand U4340 (N_4340,N_4061,N_4073);
or U4341 (N_4341,N_4049,N_4189);
xor U4342 (N_4342,N_4178,N_4053);
nand U4343 (N_4343,N_4070,N_4066);
nand U4344 (N_4344,N_4158,N_4129);
nand U4345 (N_4345,N_4155,N_4159);
nand U4346 (N_4346,N_4133,N_4147);
nand U4347 (N_4347,N_4110,N_4182);
and U4348 (N_4348,N_4173,N_4114);
nor U4349 (N_4349,N_4167,N_4128);
or U4350 (N_4350,N_4099,N_4175);
or U4351 (N_4351,N_4152,N_4071);
or U4352 (N_4352,N_4062,N_4108);
nand U4353 (N_4353,N_4105,N_4053);
and U4354 (N_4354,N_4142,N_4086);
xnor U4355 (N_4355,N_4147,N_4164);
nor U4356 (N_4356,N_4169,N_4102);
and U4357 (N_4357,N_4140,N_4112);
and U4358 (N_4358,N_4063,N_4143);
or U4359 (N_4359,N_4121,N_4138);
or U4360 (N_4360,N_4083,N_4165);
and U4361 (N_4361,N_4067,N_4074);
and U4362 (N_4362,N_4100,N_4013);
and U4363 (N_4363,N_4178,N_4005);
or U4364 (N_4364,N_4091,N_4063);
nor U4365 (N_4365,N_4049,N_4129);
nand U4366 (N_4366,N_4179,N_4083);
nor U4367 (N_4367,N_4080,N_4070);
nor U4368 (N_4368,N_4135,N_4169);
and U4369 (N_4369,N_4084,N_4116);
nand U4370 (N_4370,N_4032,N_4076);
nor U4371 (N_4371,N_4026,N_4148);
nand U4372 (N_4372,N_4044,N_4181);
and U4373 (N_4373,N_4067,N_4042);
or U4374 (N_4374,N_4181,N_4003);
or U4375 (N_4375,N_4087,N_4049);
nor U4376 (N_4376,N_4172,N_4179);
and U4377 (N_4377,N_4001,N_4125);
nor U4378 (N_4378,N_4085,N_4020);
nand U4379 (N_4379,N_4158,N_4159);
nand U4380 (N_4380,N_4143,N_4115);
and U4381 (N_4381,N_4188,N_4180);
or U4382 (N_4382,N_4044,N_4011);
nor U4383 (N_4383,N_4114,N_4121);
or U4384 (N_4384,N_4096,N_4094);
and U4385 (N_4385,N_4190,N_4025);
nand U4386 (N_4386,N_4167,N_4141);
nand U4387 (N_4387,N_4069,N_4037);
and U4388 (N_4388,N_4022,N_4086);
and U4389 (N_4389,N_4107,N_4108);
and U4390 (N_4390,N_4190,N_4106);
nand U4391 (N_4391,N_4028,N_4069);
nand U4392 (N_4392,N_4090,N_4145);
and U4393 (N_4393,N_4044,N_4154);
and U4394 (N_4394,N_4133,N_4030);
nor U4395 (N_4395,N_4120,N_4015);
or U4396 (N_4396,N_4197,N_4172);
and U4397 (N_4397,N_4167,N_4011);
nand U4398 (N_4398,N_4159,N_4090);
nand U4399 (N_4399,N_4160,N_4048);
nand U4400 (N_4400,N_4307,N_4225);
and U4401 (N_4401,N_4341,N_4357);
or U4402 (N_4402,N_4258,N_4284);
or U4403 (N_4403,N_4213,N_4324);
or U4404 (N_4404,N_4251,N_4244);
nand U4405 (N_4405,N_4374,N_4245);
and U4406 (N_4406,N_4385,N_4346);
or U4407 (N_4407,N_4369,N_4321);
xnor U4408 (N_4408,N_4399,N_4386);
or U4409 (N_4409,N_4351,N_4204);
nand U4410 (N_4410,N_4328,N_4260);
nand U4411 (N_4411,N_4222,N_4285);
and U4412 (N_4412,N_4206,N_4325);
nor U4413 (N_4413,N_4319,N_4326);
and U4414 (N_4414,N_4340,N_4229);
or U4415 (N_4415,N_4344,N_4203);
and U4416 (N_4416,N_4350,N_4280);
nand U4417 (N_4417,N_4202,N_4249);
or U4418 (N_4418,N_4308,N_4252);
xnor U4419 (N_4419,N_4335,N_4364);
xnor U4420 (N_4420,N_4309,N_4296);
or U4421 (N_4421,N_4283,N_4337);
or U4422 (N_4422,N_4233,N_4363);
nor U4423 (N_4423,N_4349,N_4231);
nand U4424 (N_4424,N_4247,N_4295);
nand U4425 (N_4425,N_4322,N_4312);
and U4426 (N_4426,N_4293,N_4348);
and U4427 (N_4427,N_4371,N_4359);
nand U4428 (N_4428,N_4212,N_4334);
nor U4429 (N_4429,N_4353,N_4393);
nor U4430 (N_4430,N_4299,N_4236);
or U4431 (N_4431,N_4288,N_4330);
nor U4432 (N_4432,N_4383,N_4224);
nand U4433 (N_4433,N_4230,N_4366);
nor U4434 (N_4434,N_4333,N_4388);
or U4435 (N_4435,N_4237,N_4358);
nor U4436 (N_4436,N_4235,N_4339);
nor U4437 (N_4437,N_4269,N_4368);
xnor U4438 (N_4438,N_4361,N_4292);
or U4439 (N_4439,N_4282,N_4271);
or U4440 (N_4440,N_4234,N_4226);
nor U4441 (N_4441,N_4318,N_4262);
or U4442 (N_4442,N_4354,N_4378);
nor U4443 (N_4443,N_4380,N_4327);
nor U4444 (N_4444,N_4273,N_4297);
and U4445 (N_4445,N_4360,N_4220);
and U4446 (N_4446,N_4270,N_4200);
xnor U4447 (N_4447,N_4395,N_4205);
or U4448 (N_4448,N_4384,N_4207);
and U4449 (N_4449,N_4215,N_4239);
xnor U4450 (N_4450,N_4209,N_4255);
xnor U4451 (N_4451,N_4331,N_4301);
nand U4452 (N_4452,N_4314,N_4355);
nor U4453 (N_4453,N_4281,N_4286);
xnor U4454 (N_4454,N_4390,N_4397);
nand U4455 (N_4455,N_4216,N_4365);
nand U4456 (N_4456,N_4242,N_4329);
or U4457 (N_4457,N_4310,N_4304);
nor U4458 (N_4458,N_4370,N_4243);
nor U4459 (N_4459,N_4223,N_4217);
xor U4460 (N_4460,N_4221,N_4256);
and U4461 (N_4461,N_4218,N_4317);
or U4462 (N_4462,N_4300,N_4291);
nor U4463 (N_4463,N_4267,N_4232);
xnor U4464 (N_4464,N_4208,N_4246);
or U4465 (N_4465,N_4290,N_4227);
or U4466 (N_4466,N_4392,N_4356);
nand U4467 (N_4467,N_4313,N_4382);
nor U4468 (N_4468,N_4289,N_4254);
or U4469 (N_4469,N_4277,N_4311);
and U4470 (N_4470,N_4373,N_4228);
xnor U4471 (N_4471,N_4320,N_4274);
and U4472 (N_4472,N_4265,N_4238);
or U4473 (N_4473,N_4323,N_4391);
nor U4474 (N_4474,N_4332,N_4315);
or U4475 (N_4475,N_4276,N_4347);
xnor U4476 (N_4476,N_4375,N_4303);
or U4477 (N_4477,N_4302,N_4261);
and U4478 (N_4478,N_4241,N_4367);
and U4479 (N_4479,N_4352,N_4305);
nand U4480 (N_4480,N_4372,N_4343);
and U4481 (N_4481,N_4272,N_4298);
nand U4482 (N_4482,N_4253,N_4396);
or U4483 (N_4483,N_4275,N_4259);
and U4484 (N_4484,N_4211,N_4381);
nor U4485 (N_4485,N_4263,N_4219);
or U4486 (N_4486,N_4387,N_4316);
and U4487 (N_4487,N_4345,N_4279);
nor U4488 (N_4488,N_4306,N_4240);
and U4489 (N_4489,N_4278,N_4268);
or U4490 (N_4490,N_4398,N_4214);
nor U4491 (N_4491,N_4336,N_4389);
nor U4492 (N_4492,N_4250,N_4377);
nand U4493 (N_4493,N_4264,N_4248);
and U4494 (N_4494,N_4210,N_4266);
nand U4495 (N_4495,N_4201,N_4287);
and U4496 (N_4496,N_4257,N_4362);
and U4497 (N_4497,N_4394,N_4342);
nor U4498 (N_4498,N_4338,N_4294);
nor U4499 (N_4499,N_4376,N_4379);
nor U4500 (N_4500,N_4243,N_4317);
and U4501 (N_4501,N_4213,N_4360);
or U4502 (N_4502,N_4235,N_4377);
or U4503 (N_4503,N_4339,N_4278);
xnor U4504 (N_4504,N_4258,N_4338);
or U4505 (N_4505,N_4366,N_4284);
nor U4506 (N_4506,N_4332,N_4263);
nand U4507 (N_4507,N_4328,N_4348);
or U4508 (N_4508,N_4309,N_4310);
nand U4509 (N_4509,N_4389,N_4207);
nand U4510 (N_4510,N_4371,N_4345);
or U4511 (N_4511,N_4270,N_4331);
or U4512 (N_4512,N_4251,N_4274);
nand U4513 (N_4513,N_4383,N_4390);
nand U4514 (N_4514,N_4223,N_4327);
and U4515 (N_4515,N_4225,N_4368);
and U4516 (N_4516,N_4246,N_4295);
nand U4517 (N_4517,N_4316,N_4276);
nand U4518 (N_4518,N_4242,N_4304);
nor U4519 (N_4519,N_4256,N_4243);
nor U4520 (N_4520,N_4360,N_4222);
nand U4521 (N_4521,N_4373,N_4202);
nand U4522 (N_4522,N_4337,N_4312);
nand U4523 (N_4523,N_4299,N_4273);
and U4524 (N_4524,N_4218,N_4262);
or U4525 (N_4525,N_4222,N_4367);
xor U4526 (N_4526,N_4360,N_4227);
and U4527 (N_4527,N_4362,N_4263);
and U4528 (N_4528,N_4243,N_4315);
xnor U4529 (N_4529,N_4390,N_4388);
and U4530 (N_4530,N_4394,N_4236);
nand U4531 (N_4531,N_4261,N_4283);
and U4532 (N_4532,N_4210,N_4392);
or U4533 (N_4533,N_4389,N_4273);
xnor U4534 (N_4534,N_4266,N_4311);
nor U4535 (N_4535,N_4264,N_4364);
xor U4536 (N_4536,N_4385,N_4225);
or U4537 (N_4537,N_4317,N_4399);
and U4538 (N_4538,N_4357,N_4329);
xnor U4539 (N_4539,N_4396,N_4350);
and U4540 (N_4540,N_4258,N_4310);
and U4541 (N_4541,N_4269,N_4369);
and U4542 (N_4542,N_4345,N_4218);
nand U4543 (N_4543,N_4308,N_4274);
nor U4544 (N_4544,N_4309,N_4339);
nor U4545 (N_4545,N_4321,N_4390);
nand U4546 (N_4546,N_4323,N_4252);
or U4547 (N_4547,N_4252,N_4313);
and U4548 (N_4548,N_4288,N_4367);
xnor U4549 (N_4549,N_4332,N_4326);
xnor U4550 (N_4550,N_4346,N_4295);
or U4551 (N_4551,N_4267,N_4374);
or U4552 (N_4552,N_4383,N_4247);
xor U4553 (N_4553,N_4386,N_4317);
nor U4554 (N_4554,N_4397,N_4234);
and U4555 (N_4555,N_4282,N_4243);
nand U4556 (N_4556,N_4309,N_4337);
or U4557 (N_4557,N_4225,N_4251);
or U4558 (N_4558,N_4319,N_4259);
and U4559 (N_4559,N_4325,N_4273);
nor U4560 (N_4560,N_4362,N_4205);
nor U4561 (N_4561,N_4384,N_4229);
nand U4562 (N_4562,N_4382,N_4217);
nand U4563 (N_4563,N_4283,N_4327);
or U4564 (N_4564,N_4331,N_4226);
or U4565 (N_4565,N_4233,N_4333);
nand U4566 (N_4566,N_4266,N_4259);
and U4567 (N_4567,N_4296,N_4390);
or U4568 (N_4568,N_4217,N_4224);
nor U4569 (N_4569,N_4358,N_4309);
nand U4570 (N_4570,N_4259,N_4315);
nand U4571 (N_4571,N_4266,N_4322);
xor U4572 (N_4572,N_4262,N_4339);
and U4573 (N_4573,N_4323,N_4201);
xor U4574 (N_4574,N_4253,N_4344);
nor U4575 (N_4575,N_4260,N_4388);
xor U4576 (N_4576,N_4320,N_4305);
xor U4577 (N_4577,N_4208,N_4289);
xor U4578 (N_4578,N_4380,N_4247);
and U4579 (N_4579,N_4221,N_4382);
or U4580 (N_4580,N_4393,N_4345);
and U4581 (N_4581,N_4347,N_4242);
xnor U4582 (N_4582,N_4255,N_4247);
xor U4583 (N_4583,N_4300,N_4385);
and U4584 (N_4584,N_4217,N_4280);
nand U4585 (N_4585,N_4363,N_4342);
xor U4586 (N_4586,N_4262,N_4263);
and U4587 (N_4587,N_4263,N_4273);
nor U4588 (N_4588,N_4246,N_4310);
nand U4589 (N_4589,N_4213,N_4205);
and U4590 (N_4590,N_4363,N_4207);
nor U4591 (N_4591,N_4214,N_4347);
nand U4592 (N_4592,N_4376,N_4352);
nand U4593 (N_4593,N_4328,N_4313);
nand U4594 (N_4594,N_4311,N_4238);
xor U4595 (N_4595,N_4340,N_4205);
or U4596 (N_4596,N_4328,N_4365);
and U4597 (N_4597,N_4359,N_4392);
nor U4598 (N_4598,N_4357,N_4363);
and U4599 (N_4599,N_4282,N_4203);
or U4600 (N_4600,N_4411,N_4487);
nand U4601 (N_4601,N_4583,N_4573);
nand U4602 (N_4602,N_4427,N_4428);
or U4603 (N_4603,N_4549,N_4563);
nor U4604 (N_4604,N_4524,N_4595);
nor U4605 (N_4605,N_4468,N_4537);
or U4606 (N_4606,N_4576,N_4435);
or U4607 (N_4607,N_4484,N_4580);
and U4608 (N_4608,N_4572,N_4598);
nor U4609 (N_4609,N_4492,N_4424);
nor U4610 (N_4610,N_4423,N_4494);
nand U4611 (N_4611,N_4543,N_4506);
nand U4612 (N_4612,N_4404,N_4504);
and U4613 (N_4613,N_4584,N_4593);
xnor U4614 (N_4614,N_4582,N_4432);
and U4615 (N_4615,N_4596,N_4415);
or U4616 (N_4616,N_4456,N_4564);
nand U4617 (N_4617,N_4536,N_4446);
nor U4618 (N_4618,N_4414,N_4416);
and U4619 (N_4619,N_4505,N_4457);
nand U4620 (N_4620,N_4480,N_4425);
and U4621 (N_4621,N_4526,N_4419);
nor U4622 (N_4622,N_4485,N_4471);
nor U4623 (N_4623,N_4532,N_4477);
or U4624 (N_4624,N_4525,N_4437);
nand U4625 (N_4625,N_4518,N_4516);
and U4626 (N_4626,N_4496,N_4531);
and U4627 (N_4627,N_4402,N_4553);
nand U4628 (N_4628,N_4412,N_4474);
or U4629 (N_4629,N_4426,N_4529);
nor U4630 (N_4630,N_4538,N_4491);
nor U4631 (N_4631,N_4574,N_4579);
or U4632 (N_4632,N_4567,N_4500);
and U4633 (N_4633,N_4522,N_4445);
and U4634 (N_4634,N_4489,N_4560);
nor U4635 (N_4635,N_4597,N_4565);
nor U4636 (N_4636,N_4463,N_4464);
nand U4637 (N_4637,N_4401,N_4586);
nor U4638 (N_4638,N_4542,N_4409);
nand U4639 (N_4639,N_4438,N_4420);
nor U4640 (N_4640,N_4514,N_4527);
nand U4641 (N_4641,N_4473,N_4444);
xnor U4642 (N_4642,N_4555,N_4433);
or U4643 (N_4643,N_4476,N_4509);
nand U4644 (N_4644,N_4460,N_4498);
and U4645 (N_4645,N_4588,N_4462);
xor U4646 (N_4646,N_4405,N_4515);
and U4647 (N_4647,N_4481,N_4510);
nand U4648 (N_4648,N_4407,N_4429);
nand U4649 (N_4649,N_4528,N_4413);
xor U4650 (N_4650,N_4459,N_4570);
or U4651 (N_4651,N_4478,N_4441);
nand U4652 (N_4652,N_4556,N_4517);
xnor U4653 (N_4653,N_4562,N_4447);
and U4654 (N_4654,N_4403,N_4568);
nand U4655 (N_4655,N_4502,N_4479);
nor U4656 (N_4656,N_4589,N_4451);
and U4657 (N_4657,N_4533,N_4512);
nor U4658 (N_4658,N_4503,N_4497);
and U4659 (N_4659,N_4535,N_4486);
or U4660 (N_4660,N_4470,N_4581);
nand U4661 (N_4661,N_4541,N_4440);
nor U4662 (N_4662,N_4434,N_4520);
nor U4663 (N_4663,N_4430,N_4507);
nor U4664 (N_4664,N_4467,N_4448);
nor U4665 (N_4665,N_4521,N_4530);
nand U4666 (N_4666,N_4453,N_4575);
nor U4667 (N_4667,N_4590,N_4548);
nor U4668 (N_4668,N_4594,N_4439);
and U4669 (N_4669,N_4569,N_4523);
or U4670 (N_4670,N_4483,N_4418);
xor U4671 (N_4671,N_4490,N_4436);
nor U4672 (N_4672,N_4550,N_4552);
or U4673 (N_4673,N_4469,N_4559);
nand U4674 (N_4674,N_4454,N_4511);
or U4675 (N_4675,N_4452,N_4475);
and U4676 (N_4676,N_4488,N_4539);
nand U4677 (N_4677,N_4466,N_4577);
nor U4678 (N_4678,N_4450,N_4431);
and U4679 (N_4679,N_4545,N_4461);
nand U4680 (N_4680,N_4482,N_4458);
and U4681 (N_4681,N_4442,N_4508);
nand U4682 (N_4682,N_4400,N_4410);
nand U4683 (N_4683,N_4546,N_4585);
nand U4684 (N_4684,N_4493,N_4587);
and U4685 (N_4685,N_4501,N_4557);
or U4686 (N_4686,N_4417,N_4561);
xnor U4687 (N_4687,N_4499,N_4421);
and U4688 (N_4688,N_4408,N_4472);
nor U4689 (N_4689,N_4551,N_4513);
nor U4690 (N_4690,N_4544,N_4465);
nand U4691 (N_4691,N_4455,N_4443);
nor U4692 (N_4692,N_4571,N_4406);
nand U4693 (N_4693,N_4495,N_4554);
nand U4694 (N_4694,N_4592,N_4547);
nand U4695 (N_4695,N_4566,N_4591);
and U4696 (N_4696,N_4519,N_4422);
or U4697 (N_4697,N_4578,N_4599);
xor U4698 (N_4698,N_4558,N_4540);
nand U4699 (N_4699,N_4449,N_4534);
and U4700 (N_4700,N_4449,N_4571);
xor U4701 (N_4701,N_4588,N_4448);
nand U4702 (N_4702,N_4412,N_4555);
xnor U4703 (N_4703,N_4495,N_4578);
xnor U4704 (N_4704,N_4506,N_4540);
nor U4705 (N_4705,N_4422,N_4538);
xor U4706 (N_4706,N_4456,N_4523);
nand U4707 (N_4707,N_4412,N_4569);
xor U4708 (N_4708,N_4407,N_4569);
and U4709 (N_4709,N_4444,N_4583);
or U4710 (N_4710,N_4486,N_4527);
nor U4711 (N_4711,N_4426,N_4551);
nor U4712 (N_4712,N_4410,N_4573);
or U4713 (N_4713,N_4485,N_4508);
and U4714 (N_4714,N_4476,N_4503);
or U4715 (N_4715,N_4411,N_4501);
nor U4716 (N_4716,N_4405,N_4592);
nor U4717 (N_4717,N_4592,N_4577);
nor U4718 (N_4718,N_4508,N_4513);
or U4719 (N_4719,N_4467,N_4435);
nand U4720 (N_4720,N_4423,N_4514);
nor U4721 (N_4721,N_4552,N_4584);
nor U4722 (N_4722,N_4492,N_4512);
or U4723 (N_4723,N_4451,N_4551);
and U4724 (N_4724,N_4506,N_4401);
nand U4725 (N_4725,N_4571,N_4506);
or U4726 (N_4726,N_4474,N_4591);
nor U4727 (N_4727,N_4455,N_4522);
nor U4728 (N_4728,N_4417,N_4407);
and U4729 (N_4729,N_4529,N_4487);
xnor U4730 (N_4730,N_4408,N_4455);
nand U4731 (N_4731,N_4581,N_4466);
nor U4732 (N_4732,N_4472,N_4568);
xor U4733 (N_4733,N_4472,N_4563);
nand U4734 (N_4734,N_4439,N_4417);
and U4735 (N_4735,N_4492,N_4586);
and U4736 (N_4736,N_4543,N_4570);
and U4737 (N_4737,N_4413,N_4495);
nor U4738 (N_4738,N_4596,N_4501);
nor U4739 (N_4739,N_4445,N_4591);
and U4740 (N_4740,N_4501,N_4443);
or U4741 (N_4741,N_4435,N_4481);
or U4742 (N_4742,N_4441,N_4448);
and U4743 (N_4743,N_4546,N_4588);
nand U4744 (N_4744,N_4517,N_4544);
or U4745 (N_4745,N_4487,N_4582);
nand U4746 (N_4746,N_4552,N_4490);
nand U4747 (N_4747,N_4557,N_4518);
or U4748 (N_4748,N_4543,N_4471);
and U4749 (N_4749,N_4482,N_4411);
nor U4750 (N_4750,N_4438,N_4472);
nand U4751 (N_4751,N_4547,N_4559);
or U4752 (N_4752,N_4445,N_4511);
xor U4753 (N_4753,N_4479,N_4498);
xnor U4754 (N_4754,N_4525,N_4433);
and U4755 (N_4755,N_4403,N_4586);
xnor U4756 (N_4756,N_4504,N_4571);
xnor U4757 (N_4757,N_4509,N_4590);
or U4758 (N_4758,N_4424,N_4522);
and U4759 (N_4759,N_4418,N_4570);
or U4760 (N_4760,N_4437,N_4501);
nand U4761 (N_4761,N_4489,N_4445);
and U4762 (N_4762,N_4416,N_4421);
nand U4763 (N_4763,N_4560,N_4427);
xor U4764 (N_4764,N_4585,N_4590);
xnor U4765 (N_4765,N_4507,N_4527);
or U4766 (N_4766,N_4457,N_4467);
or U4767 (N_4767,N_4570,N_4546);
and U4768 (N_4768,N_4425,N_4404);
nand U4769 (N_4769,N_4541,N_4460);
and U4770 (N_4770,N_4450,N_4438);
nand U4771 (N_4771,N_4522,N_4583);
nor U4772 (N_4772,N_4523,N_4572);
or U4773 (N_4773,N_4560,N_4488);
or U4774 (N_4774,N_4555,N_4546);
nor U4775 (N_4775,N_4434,N_4565);
nor U4776 (N_4776,N_4522,N_4557);
and U4777 (N_4777,N_4592,N_4440);
xor U4778 (N_4778,N_4504,N_4541);
nor U4779 (N_4779,N_4445,N_4527);
nor U4780 (N_4780,N_4419,N_4553);
nor U4781 (N_4781,N_4535,N_4507);
nor U4782 (N_4782,N_4496,N_4591);
and U4783 (N_4783,N_4440,N_4490);
or U4784 (N_4784,N_4594,N_4536);
and U4785 (N_4785,N_4493,N_4459);
or U4786 (N_4786,N_4468,N_4470);
or U4787 (N_4787,N_4516,N_4424);
nor U4788 (N_4788,N_4558,N_4463);
and U4789 (N_4789,N_4469,N_4575);
and U4790 (N_4790,N_4485,N_4584);
and U4791 (N_4791,N_4520,N_4508);
nand U4792 (N_4792,N_4518,N_4590);
nand U4793 (N_4793,N_4454,N_4473);
and U4794 (N_4794,N_4403,N_4459);
nor U4795 (N_4795,N_4589,N_4550);
and U4796 (N_4796,N_4433,N_4530);
nand U4797 (N_4797,N_4521,N_4490);
and U4798 (N_4798,N_4442,N_4417);
nor U4799 (N_4799,N_4470,N_4489);
nor U4800 (N_4800,N_4610,N_4795);
xor U4801 (N_4801,N_4701,N_4727);
and U4802 (N_4802,N_4758,N_4694);
nor U4803 (N_4803,N_4615,N_4789);
or U4804 (N_4804,N_4778,N_4638);
nand U4805 (N_4805,N_4613,N_4702);
and U4806 (N_4806,N_4611,N_4751);
or U4807 (N_4807,N_4743,N_4641);
or U4808 (N_4808,N_4606,N_4666);
nor U4809 (N_4809,N_4734,N_4756);
nor U4810 (N_4810,N_4621,N_4784);
nor U4811 (N_4811,N_4739,N_4726);
or U4812 (N_4812,N_4763,N_4632);
nor U4813 (N_4813,N_4740,N_4735);
or U4814 (N_4814,N_4768,N_4719);
nand U4815 (N_4815,N_4607,N_4733);
and U4816 (N_4816,N_4602,N_4648);
xor U4817 (N_4817,N_4637,N_4620);
and U4818 (N_4818,N_4672,N_4639);
and U4819 (N_4819,N_4731,N_4600);
nor U4820 (N_4820,N_4652,N_4781);
or U4821 (N_4821,N_4722,N_4640);
xnor U4822 (N_4822,N_4761,N_4715);
nor U4823 (N_4823,N_4757,N_4604);
nor U4824 (N_4824,N_4630,N_4732);
nand U4825 (N_4825,N_4646,N_4619);
and U4826 (N_4826,N_4780,N_4728);
and U4827 (N_4827,N_4710,N_4754);
nor U4828 (N_4828,N_4764,N_4762);
or U4829 (N_4829,N_4705,N_4643);
nor U4830 (N_4830,N_4696,N_4746);
or U4831 (N_4831,N_4624,N_4708);
nor U4832 (N_4832,N_4798,N_4683);
nor U4833 (N_4833,N_4797,N_4738);
nor U4834 (N_4834,N_4633,N_4603);
xnor U4835 (N_4835,N_4647,N_4659);
nor U4836 (N_4836,N_4662,N_4770);
nor U4837 (N_4837,N_4748,N_4676);
nor U4838 (N_4838,N_4622,N_4723);
or U4839 (N_4839,N_4707,N_4786);
nor U4840 (N_4840,N_4721,N_4777);
nand U4841 (N_4841,N_4767,N_4601);
xor U4842 (N_4842,N_4745,N_4670);
nand U4843 (N_4843,N_4725,N_4626);
or U4844 (N_4844,N_4799,N_4609);
nand U4845 (N_4845,N_4689,N_4627);
and U4846 (N_4846,N_4635,N_4629);
nor U4847 (N_4847,N_4703,N_4736);
nand U4848 (N_4848,N_4654,N_4680);
or U4849 (N_4849,N_4724,N_4644);
and U4850 (N_4850,N_4779,N_4753);
or U4851 (N_4851,N_4704,N_4608);
and U4852 (N_4852,N_4663,N_4712);
or U4853 (N_4853,N_4690,N_4782);
and U4854 (N_4854,N_4673,N_4628);
or U4855 (N_4855,N_4634,N_4636);
or U4856 (N_4856,N_4691,N_4656);
and U4857 (N_4857,N_4614,N_4776);
and U4858 (N_4858,N_4792,N_4669);
nor U4859 (N_4859,N_4688,N_4766);
nand U4860 (N_4860,N_4750,N_4625);
or U4861 (N_4861,N_4671,N_4759);
and U4862 (N_4862,N_4623,N_4700);
or U4863 (N_4863,N_4677,N_4665);
and U4864 (N_4864,N_4699,N_4649);
and U4865 (N_4865,N_4692,N_4791);
or U4866 (N_4866,N_4729,N_4769);
nand U4867 (N_4867,N_4749,N_4742);
and U4868 (N_4868,N_4657,N_4687);
and U4869 (N_4869,N_4771,N_4709);
nand U4870 (N_4870,N_4658,N_4716);
and U4871 (N_4871,N_4773,N_4655);
and U4872 (N_4872,N_4720,N_4775);
nand U4873 (N_4873,N_4681,N_4737);
nand U4874 (N_4874,N_4664,N_4772);
and U4875 (N_4875,N_4617,N_4645);
or U4876 (N_4876,N_4668,N_4783);
nor U4877 (N_4877,N_4741,N_4618);
nor U4878 (N_4878,N_4765,N_4612);
nor U4879 (N_4879,N_4711,N_4718);
nand U4880 (N_4880,N_4787,N_4674);
and U4881 (N_4881,N_4685,N_4679);
nor U4882 (N_4882,N_4744,N_4793);
nor U4883 (N_4883,N_4714,N_4695);
or U4884 (N_4884,N_4682,N_4774);
nand U4885 (N_4885,N_4686,N_4660);
nand U4886 (N_4886,N_4730,N_4693);
and U4887 (N_4887,N_4752,N_4706);
xor U4888 (N_4888,N_4631,N_4684);
or U4889 (N_4889,N_4760,N_4713);
and U4890 (N_4890,N_4788,N_4697);
nand U4891 (N_4891,N_4616,N_4675);
and U4892 (N_4892,N_4717,N_4796);
nand U4893 (N_4893,N_4661,N_4698);
nand U4894 (N_4894,N_4790,N_4605);
nor U4895 (N_4895,N_4667,N_4755);
and U4896 (N_4896,N_4650,N_4651);
xnor U4897 (N_4897,N_4642,N_4794);
and U4898 (N_4898,N_4747,N_4785);
or U4899 (N_4899,N_4678,N_4653);
nand U4900 (N_4900,N_4624,N_4715);
nor U4901 (N_4901,N_4759,N_4770);
or U4902 (N_4902,N_4779,N_4799);
xor U4903 (N_4903,N_4779,N_4692);
xor U4904 (N_4904,N_4607,N_4688);
and U4905 (N_4905,N_4648,N_4794);
nand U4906 (N_4906,N_4756,N_4646);
and U4907 (N_4907,N_4696,N_4688);
nand U4908 (N_4908,N_4618,N_4731);
nand U4909 (N_4909,N_4739,N_4755);
nor U4910 (N_4910,N_4740,N_4626);
or U4911 (N_4911,N_4660,N_4683);
xnor U4912 (N_4912,N_4785,N_4671);
nor U4913 (N_4913,N_4661,N_4658);
or U4914 (N_4914,N_4636,N_4773);
nand U4915 (N_4915,N_4603,N_4636);
nor U4916 (N_4916,N_4778,N_4768);
nand U4917 (N_4917,N_4708,N_4640);
nor U4918 (N_4918,N_4711,N_4674);
xnor U4919 (N_4919,N_4755,N_4798);
nor U4920 (N_4920,N_4718,N_4780);
and U4921 (N_4921,N_4711,N_4697);
and U4922 (N_4922,N_4657,N_4636);
or U4923 (N_4923,N_4743,N_4735);
nand U4924 (N_4924,N_4716,N_4797);
nand U4925 (N_4925,N_4654,N_4615);
nor U4926 (N_4926,N_4615,N_4798);
nand U4927 (N_4927,N_4680,N_4666);
nor U4928 (N_4928,N_4733,N_4693);
and U4929 (N_4929,N_4703,N_4739);
and U4930 (N_4930,N_4761,N_4695);
nand U4931 (N_4931,N_4745,N_4766);
or U4932 (N_4932,N_4655,N_4732);
nand U4933 (N_4933,N_4620,N_4755);
nand U4934 (N_4934,N_4694,N_4636);
nor U4935 (N_4935,N_4693,N_4783);
and U4936 (N_4936,N_4685,N_4600);
and U4937 (N_4937,N_4761,N_4738);
and U4938 (N_4938,N_4720,N_4756);
nand U4939 (N_4939,N_4718,N_4752);
or U4940 (N_4940,N_4693,N_4634);
nand U4941 (N_4941,N_4790,N_4776);
nor U4942 (N_4942,N_4775,N_4681);
nor U4943 (N_4943,N_4739,N_4756);
nand U4944 (N_4944,N_4717,N_4780);
nand U4945 (N_4945,N_4780,N_4733);
or U4946 (N_4946,N_4798,N_4629);
or U4947 (N_4947,N_4671,N_4657);
xnor U4948 (N_4948,N_4612,N_4615);
nand U4949 (N_4949,N_4724,N_4611);
nand U4950 (N_4950,N_4759,N_4665);
nor U4951 (N_4951,N_4633,N_4696);
and U4952 (N_4952,N_4751,N_4740);
or U4953 (N_4953,N_4782,N_4795);
xnor U4954 (N_4954,N_4790,N_4770);
nand U4955 (N_4955,N_4740,N_4768);
and U4956 (N_4956,N_4649,N_4635);
nor U4957 (N_4957,N_4747,N_4685);
or U4958 (N_4958,N_4660,N_4617);
and U4959 (N_4959,N_4610,N_4758);
nand U4960 (N_4960,N_4624,N_4760);
nand U4961 (N_4961,N_4637,N_4702);
nor U4962 (N_4962,N_4674,N_4719);
or U4963 (N_4963,N_4728,N_4671);
xor U4964 (N_4964,N_4600,N_4727);
nand U4965 (N_4965,N_4726,N_4797);
and U4966 (N_4966,N_4602,N_4781);
nor U4967 (N_4967,N_4678,N_4625);
nand U4968 (N_4968,N_4668,N_4798);
xnor U4969 (N_4969,N_4610,N_4751);
or U4970 (N_4970,N_4776,N_4747);
nor U4971 (N_4971,N_4723,N_4745);
nand U4972 (N_4972,N_4660,N_4640);
xnor U4973 (N_4973,N_4779,N_4683);
nand U4974 (N_4974,N_4758,N_4606);
xor U4975 (N_4975,N_4725,N_4610);
nand U4976 (N_4976,N_4652,N_4639);
or U4977 (N_4977,N_4739,N_4671);
nor U4978 (N_4978,N_4638,N_4767);
nor U4979 (N_4979,N_4767,N_4752);
nor U4980 (N_4980,N_4678,N_4672);
xnor U4981 (N_4981,N_4619,N_4718);
nand U4982 (N_4982,N_4642,N_4776);
nor U4983 (N_4983,N_4743,N_4695);
and U4984 (N_4984,N_4675,N_4660);
and U4985 (N_4985,N_4679,N_4640);
nand U4986 (N_4986,N_4718,N_4637);
nand U4987 (N_4987,N_4674,N_4701);
nor U4988 (N_4988,N_4748,N_4755);
or U4989 (N_4989,N_4638,N_4785);
and U4990 (N_4990,N_4603,N_4717);
nand U4991 (N_4991,N_4709,N_4658);
and U4992 (N_4992,N_4722,N_4797);
nor U4993 (N_4993,N_4687,N_4682);
or U4994 (N_4994,N_4627,N_4765);
or U4995 (N_4995,N_4739,N_4789);
or U4996 (N_4996,N_4633,N_4790);
and U4997 (N_4997,N_4715,N_4676);
nor U4998 (N_4998,N_4785,N_4607);
nand U4999 (N_4999,N_4642,N_4667);
and UO_0 (O_0,N_4997,N_4998);
nand UO_1 (O_1,N_4890,N_4937);
or UO_2 (O_2,N_4940,N_4802);
or UO_3 (O_3,N_4929,N_4949);
or UO_4 (O_4,N_4848,N_4861);
and UO_5 (O_5,N_4850,N_4892);
or UO_6 (O_6,N_4862,N_4962);
nand UO_7 (O_7,N_4883,N_4953);
nor UO_8 (O_8,N_4910,N_4809);
or UO_9 (O_9,N_4894,N_4915);
nand UO_10 (O_10,N_4877,N_4983);
nand UO_11 (O_11,N_4838,N_4907);
or UO_12 (O_12,N_4884,N_4930);
and UO_13 (O_13,N_4827,N_4934);
or UO_14 (O_14,N_4908,N_4987);
or UO_15 (O_15,N_4855,N_4904);
or UO_16 (O_16,N_4918,N_4852);
and UO_17 (O_17,N_4825,N_4868);
and UO_18 (O_18,N_4818,N_4831);
xnor UO_19 (O_19,N_4941,N_4836);
and UO_20 (O_20,N_4860,N_4970);
nor UO_21 (O_21,N_4826,N_4834);
nor UO_22 (O_22,N_4978,N_4810);
nor UO_23 (O_23,N_4963,N_4866);
xor UO_24 (O_24,N_4980,N_4916);
nand UO_25 (O_25,N_4820,N_4901);
xnor UO_26 (O_26,N_4927,N_4996);
nand UO_27 (O_27,N_4975,N_4951);
or UO_28 (O_28,N_4992,N_4812);
or UO_29 (O_29,N_4872,N_4986);
xnor UO_30 (O_30,N_4800,N_4909);
nor UO_31 (O_31,N_4804,N_4928);
and UO_32 (O_32,N_4981,N_4865);
and UO_33 (O_33,N_4973,N_4931);
nor UO_34 (O_34,N_4840,N_4921);
and UO_35 (O_35,N_4988,N_4943);
or UO_36 (O_36,N_4914,N_4801);
or UO_37 (O_37,N_4864,N_4858);
or UO_38 (O_38,N_4895,N_4964);
nand UO_39 (O_39,N_4869,N_4896);
nand UO_40 (O_40,N_4832,N_4830);
and UO_41 (O_41,N_4829,N_4935);
and UO_42 (O_42,N_4922,N_4936);
or UO_43 (O_43,N_4985,N_4903);
nor UO_44 (O_44,N_4821,N_4885);
or UO_45 (O_45,N_4873,N_4954);
and UO_46 (O_46,N_4841,N_4845);
nand UO_47 (O_47,N_4905,N_4969);
nor UO_48 (O_48,N_4984,N_4925);
nand UO_49 (O_49,N_4950,N_4815);
nand UO_50 (O_50,N_4991,N_4839);
and UO_51 (O_51,N_4944,N_4961);
nand UO_52 (O_52,N_4976,N_4814);
or UO_53 (O_53,N_4847,N_4882);
xnor UO_54 (O_54,N_4990,N_4870);
and UO_55 (O_55,N_4958,N_4971);
xor UO_56 (O_56,N_4968,N_4851);
or UO_57 (O_57,N_4875,N_4849);
nor UO_58 (O_58,N_4919,N_4822);
and UO_59 (O_59,N_4955,N_4967);
and UO_60 (O_60,N_4989,N_4833);
nor UO_61 (O_61,N_4876,N_4853);
and UO_62 (O_62,N_4911,N_4982);
xor UO_63 (O_63,N_4906,N_4899);
or UO_64 (O_64,N_4817,N_4898);
xor UO_65 (O_65,N_4867,N_4857);
or UO_66 (O_66,N_4881,N_4888);
nor UO_67 (O_67,N_4900,N_4965);
nor UO_68 (O_68,N_4854,N_4926);
xnor UO_69 (O_69,N_4917,N_4977);
or UO_70 (O_70,N_4924,N_4879);
or UO_71 (O_71,N_4979,N_4912);
nand UO_72 (O_72,N_4999,N_4803);
nor UO_73 (O_73,N_4939,N_4811);
xnor UO_74 (O_74,N_4956,N_4843);
nor UO_75 (O_75,N_4835,N_4871);
nor UO_76 (O_76,N_4807,N_4947);
nand UO_77 (O_77,N_4880,N_4932);
or UO_78 (O_78,N_4923,N_4946);
nor UO_79 (O_79,N_4886,N_4844);
nor UO_80 (O_80,N_4893,N_4957);
nor UO_81 (O_81,N_4952,N_4945);
xor UO_82 (O_82,N_4842,N_4995);
or UO_83 (O_83,N_4828,N_4994);
nand UO_84 (O_84,N_4805,N_4806);
nor UO_85 (O_85,N_4824,N_4813);
or UO_86 (O_86,N_4816,N_4846);
nand UO_87 (O_87,N_4913,N_4942);
and UO_88 (O_88,N_4808,N_4933);
xnor UO_89 (O_89,N_4897,N_4889);
xnor UO_90 (O_90,N_4887,N_4863);
and UO_91 (O_91,N_4959,N_4856);
or UO_92 (O_92,N_4823,N_4874);
xnor UO_93 (O_93,N_4920,N_4974);
or UO_94 (O_94,N_4902,N_4948);
nor UO_95 (O_95,N_4837,N_4819);
nand UO_96 (O_96,N_4972,N_4966);
nor UO_97 (O_97,N_4891,N_4938);
or UO_98 (O_98,N_4878,N_4993);
or UO_99 (O_99,N_4960,N_4859);
and UO_100 (O_100,N_4852,N_4943);
nand UO_101 (O_101,N_4854,N_4811);
nor UO_102 (O_102,N_4909,N_4849);
xor UO_103 (O_103,N_4970,N_4825);
or UO_104 (O_104,N_4835,N_4817);
or UO_105 (O_105,N_4872,N_4866);
or UO_106 (O_106,N_4816,N_4964);
and UO_107 (O_107,N_4945,N_4955);
and UO_108 (O_108,N_4866,N_4885);
nor UO_109 (O_109,N_4856,N_4839);
nand UO_110 (O_110,N_4828,N_4924);
nor UO_111 (O_111,N_4955,N_4900);
nand UO_112 (O_112,N_4886,N_4900);
nand UO_113 (O_113,N_4975,N_4878);
nor UO_114 (O_114,N_4975,N_4981);
or UO_115 (O_115,N_4944,N_4805);
nor UO_116 (O_116,N_4913,N_4958);
nor UO_117 (O_117,N_4978,N_4941);
nand UO_118 (O_118,N_4858,N_4810);
nor UO_119 (O_119,N_4821,N_4850);
and UO_120 (O_120,N_4806,N_4834);
xor UO_121 (O_121,N_4814,N_4804);
nand UO_122 (O_122,N_4836,N_4835);
nor UO_123 (O_123,N_4893,N_4903);
and UO_124 (O_124,N_4965,N_4806);
and UO_125 (O_125,N_4831,N_4868);
nand UO_126 (O_126,N_4917,N_4804);
nand UO_127 (O_127,N_4904,N_4827);
or UO_128 (O_128,N_4859,N_4812);
xnor UO_129 (O_129,N_4916,N_4879);
nor UO_130 (O_130,N_4837,N_4840);
nand UO_131 (O_131,N_4879,N_4994);
nand UO_132 (O_132,N_4907,N_4809);
or UO_133 (O_133,N_4926,N_4911);
and UO_134 (O_134,N_4889,N_4844);
and UO_135 (O_135,N_4898,N_4915);
nor UO_136 (O_136,N_4992,N_4839);
nand UO_137 (O_137,N_4857,N_4814);
nor UO_138 (O_138,N_4961,N_4829);
xor UO_139 (O_139,N_4811,N_4911);
and UO_140 (O_140,N_4904,N_4867);
or UO_141 (O_141,N_4873,N_4979);
nor UO_142 (O_142,N_4945,N_4839);
nand UO_143 (O_143,N_4802,N_4823);
nor UO_144 (O_144,N_4975,N_4976);
nand UO_145 (O_145,N_4803,N_4876);
and UO_146 (O_146,N_4920,N_4842);
nand UO_147 (O_147,N_4935,N_4840);
or UO_148 (O_148,N_4925,N_4825);
or UO_149 (O_149,N_4926,N_4820);
or UO_150 (O_150,N_4885,N_4850);
nand UO_151 (O_151,N_4967,N_4894);
or UO_152 (O_152,N_4974,N_4895);
nand UO_153 (O_153,N_4813,N_4984);
or UO_154 (O_154,N_4840,N_4942);
xnor UO_155 (O_155,N_4842,N_4898);
and UO_156 (O_156,N_4878,N_4856);
xor UO_157 (O_157,N_4856,N_4975);
and UO_158 (O_158,N_4944,N_4970);
and UO_159 (O_159,N_4994,N_4840);
xor UO_160 (O_160,N_4895,N_4878);
nor UO_161 (O_161,N_4837,N_4952);
xnor UO_162 (O_162,N_4857,N_4967);
and UO_163 (O_163,N_4991,N_4840);
or UO_164 (O_164,N_4972,N_4958);
and UO_165 (O_165,N_4800,N_4867);
xor UO_166 (O_166,N_4982,N_4974);
nand UO_167 (O_167,N_4973,N_4843);
xnor UO_168 (O_168,N_4916,N_4913);
and UO_169 (O_169,N_4896,N_4839);
nand UO_170 (O_170,N_4880,N_4937);
or UO_171 (O_171,N_4809,N_4949);
and UO_172 (O_172,N_4831,N_4890);
or UO_173 (O_173,N_4869,N_4859);
or UO_174 (O_174,N_4976,N_4872);
and UO_175 (O_175,N_4883,N_4900);
nor UO_176 (O_176,N_4839,N_4894);
or UO_177 (O_177,N_4973,N_4962);
nand UO_178 (O_178,N_4890,N_4842);
and UO_179 (O_179,N_4824,N_4942);
nand UO_180 (O_180,N_4953,N_4946);
or UO_181 (O_181,N_4978,N_4932);
nand UO_182 (O_182,N_4870,N_4911);
nor UO_183 (O_183,N_4991,N_4865);
nor UO_184 (O_184,N_4862,N_4966);
nand UO_185 (O_185,N_4890,N_4918);
nand UO_186 (O_186,N_4954,N_4842);
nand UO_187 (O_187,N_4976,N_4956);
or UO_188 (O_188,N_4864,N_4910);
and UO_189 (O_189,N_4913,N_4873);
nor UO_190 (O_190,N_4956,N_4907);
or UO_191 (O_191,N_4883,N_4877);
nor UO_192 (O_192,N_4838,N_4968);
nor UO_193 (O_193,N_4981,N_4894);
nand UO_194 (O_194,N_4936,N_4837);
nand UO_195 (O_195,N_4907,N_4938);
nand UO_196 (O_196,N_4875,N_4813);
nor UO_197 (O_197,N_4928,N_4974);
nand UO_198 (O_198,N_4806,N_4928);
or UO_199 (O_199,N_4883,N_4816);
nor UO_200 (O_200,N_4955,N_4848);
or UO_201 (O_201,N_4890,N_4830);
nor UO_202 (O_202,N_4863,N_4870);
and UO_203 (O_203,N_4899,N_4832);
xor UO_204 (O_204,N_4887,N_4813);
nor UO_205 (O_205,N_4910,N_4974);
or UO_206 (O_206,N_4941,N_4845);
and UO_207 (O_207,N_4946,N_4904);
nand UO_208 (O_208,N_4837,N_4971);
and UO_209 (O_209,N_4971,N_4887);
and UO_210 (O_210,N_4890,N_4803);
nor UO_211 (O_211,N_4957,N_4910);
xnor UO_212 (O_212,N_4812,N_4962);
nor UO_213 (O_213,N_4877,N_4814);
and UO_214 (O_214,N_4918,N_4900);
or UO_215 (O_215,N_4880,N_4814);
nand UO_216 (O_216,N_4931,N_4928);
or UO_217 (O_217,N_4816,N_4827);
xnor UO_218 (O_218,N_4921,N_4819);
nor UO_219 (O_219,N_4997,N_4815);
and UO_220 (O_220,N_4997,N_4890);
nor UO_221 (O_221,N_4950,N_4921);
and UO_222 (O_222,N_4962,N_4834);
nor UO_223 (O_223,N_4833,N_4932);
or UO_224 (O_224,N_4993,N_4930);
xnor UO_225 (O_225,N_4827,N_4896);
nand UO_226 (O_226,N_4978,N_4824);
or UO_227 (O_227,N_4990,N_4881);
or UO_228 (O_228,N_4911,N_4835);
nor UO_229 (O_229,N_4922,N_4964);
nand UO_230 (O_230,N_4833,N_4854);
and UO_231 (O_231,N_4957,N_4883);
xnor UO_232 (O_232,N_4977,N_4813);
nor UO_233 (O_233,N_4839,N_4980);
nor UO_234 (O_234,N_4825,N_4960);
nand UO_235 (O_235,N_4810,N_4975);
nor UO_236 (O_236,N_4889,N_4871);
and UO_237 (O_237,N_4825,N_4977);
or UO_238 (O_238,N_4902,N_4831);
and UO_239 (O_239,N_4894,N_4853);
or UO_240 (O_240,N_4801,N_4919);
nand UO_241 (O_241,N_4850,N_4886);
nor UO_242 (O_242,N_4961,N_4877);
nand UO_243 (O_243,N_4933,N_4927);
nand UO_244 (O_244,N_4854,N_4924);
xor UO_245 (O_245,N_4929,N_4996);
or UO_246 (O_246,N_4926,N_4881);
nor UO_247 (O_247,N_4979,N_4812);
and UO_248 (O_248,N_4839,N_4910);
xnor UO_249 (O_249,N_4964,N_4818);
or UO_250 (O_250,N_4913,N_4810);
xor UO_251 (O_251,N_4970,N_4968);
or UO_252 (O_252,N_4992,N_4961);
nand UO_253 (O_253,N_4881,N_4910);
nor UO_254 (O_254,N_4860,N_4918);
and UO_255 (O_255,N_4893,N_4856);
nor UO_256 (O_256,N_4979,N_4898);
and UO_257 (O_257,N_4887,N_4986);
or UO_258 (O_258,N_4949,N_4911);
xnor UO_259 (O_259,N_4984,N_4964);
nor UO_260 (O_260,N_4850,N_4987);
or UO_261 (O_261,N_4893,N_4896);
or UO_262 (O_262,N_4913,N_4816);
nand UO_263 (O_263,N_4811,N_4835);
or UO_264 (O_264,N_4857,N_4968);
and UO_265 (O_265,N_4998,N_4977);
and UO_266 (O_266,N_4913,N_4961);
nand UO_267 (O_267,N_4896,N_4945);
or UO_268 (O_268,N_4933,N_4892);
or UO_269 (O_269,N_4979,N_4961);
or UO_270 (O_270,N_4901,N_4873);
nand UO_271 (O_271,N_4965,N_4989);
and UO_272 (O_272,N_4948,N_4953);
nor UO_273 (O_273,N_4826,N_4838);
nand UO_274 (O_274,N_4998,N_4925);
and UO_275 (O_275,N_4804,N_4966);
nand UO_276 (O_276,N_4926,N_4839);
or UO_277 (O_277,N_4970,N_4962);
nor UO_278 (O_278,N_4938,N_4813);
nor UO_279 (O_279,N_4855,N_4948);
nand UO_280 (O_280,N_4982,N_4824);
xor UO_281 (O_281,N_4899,N_4990);
or UO_282 (O_282,N_4882,N_4887);
nand UO_283 (O_283,N_4939,N_4831);
nand UO_284 (O_284,N_4902,N_4809);
or UO_285 (O_285,N_4973,N_4835);
nand UO_286 (O_286,N_4937,N_4945);
and UO_287 (O_287,N_4839,N_4818);
nor UO_288 (O_288,N_4926,N_4912);
nor UO_289 (O_289,N_4911,N_4922);
nand UO_290 (O_290,N_4929,N_4843);
nand UO_291 (O_291,N_4943,N_4974);
and UO_292 (O_292,N_4909,N_4826);
or UO_293 (O_293,N_4853,N_4988);
nor UO_294 (O_294,N_4973,N_4965);
nor UO_295 (O_295,N_4912,N_4920);
and UO_296 (O_296,N_4830,N_4973);
nand UO_297 (O_297,N_4809,N_4891);
nand UO_298 (O_298,N_4800,N_4961);
nand UO_299 (O_299,N_4907,N_4922);
nor UO_300 (O_300,N_4962,N_4856);
nand UO_301 (O_301,N_4932,N_4908);
nand UO_302 (O_302,N_4987,N_4906);
nand UO_303 (O_303,N_4929,N_4818);
or UO_304 (O_304,N_4925,N_4869);
nor UO_305 (O_305,N_4937,N_4903);
or UO_306 (O_306,N_4950,N_4899);
and UO_307 (O_307,N_4981,N_4961);
nand UO_308 (O_308,N_4978,N_4811);
nor UO_309 (O_309,N_4851,N_4909);
nor UO_310 (O_310,N_4867,N_4932);
and UO_311 (O_311,N_4814,N_4979);
nor UO_312 (O_312,N_4908,N_4824);
and UO_313 (O_313,N_4816,N_4943);
nor UO_314 (O_314,N_4962,N_4938);
nor UO_315 (O_315,N_4939,N_4803);
nand UO_316 (O_316,N_4873,N_4941);
and UO_317 (O_317,N_4890,N_4893);
or UO_318 (O_318,N_4844,N_4946);
nor UO_319 (O_319,N_4812,N_4854);
nor UO_320 (O_320,N_4933,N_4894);
nand UO_321 (O_321,N_4914,N_4806);
or UO_322 (O_322,N_4979,N_4803);
nor UO_323 (O_323,N_4894,N_4931);
nand UO_324 (O_324,N_4853,N_4966);
and UO_325 (O_325,N_4919,N_4873);
and UO_326 (O_326,N_4803,N_4870);
and UO_327 (O_327,N_4912,N_4944);
xor UO_328 (O_328,N_4859,N_4815);
nor UO_329 (O_329,N_4987,N_4868);
and UO_330 (O_330,N_4866,N_4847);
nor UO_331 (O_331,N_4907,N_4972);
nor UO_332 (O_332,N_4958,N_4964);
nand UO_333 (O_333,N_4955,N_4891);
nand UO_334 (O_334,N_4959,N_4997);
nor UO_335 (O_335,N_4819,N_4975);
and UO_336 (O_336,N_4813,N_4899);
nor UO_337 (O_337,N_4829,N_4981);
or UO_338 (O_338,N_4862,N_4990);
nor UO_339 (O_339,N_4893,N_4912);
nand UO_340 (O_340,N_4832,N_4848);
nand UO_341 (O_341,N_4844,N_4935);
and UO_342 (O_342,N_4920,N_4877);
or UO_343 (O_343,N_4875,N_4984);
or UO_344 (O_344,N_4827,N_4810);
xnor UO_345 (O_345,N_4992,N_4964);
or UO_346 (O_346,N_4886,N_4927);
or UO_347 (O_347,N_4987,N_4851);
xor UO_348 (O_348,N_4819,N_4967);
or UO_349 (O_349,N_4950,N_4814);
nor UO_350 (O_350,N_4924,N_4873);
nor UO_351 (O_351,N_4974,N_4835);
nand UO_352 (O_352,N_4826,N_4921);
nor UO_353 (O_353,N_4908,N_4809);
nand UO_354 (O_354,N_4868,N_4886);
or UO_355 (O_355,N_4890,N_4869);
and UO_356 (O_356,N_4844,N_4939);
and UO_357 (O_357,N_4953,N_4825);
or UO_358 (O_358,N_4916,N_4885);
or UO_359 (O_359,N_4954,N_4910);
or UO_360 (O_360,N_4915,N_4968);
nand UO_361 (O_361,N_4889,N_4913);
nor UO_362 (O_362,N_4880,N_4977);
nor UO_363 (O_363,N_4993,N_4991);
xor UO_364 (O_364,N_4902,N_4882);
or UO_365 (O_365,N_4805,N_4976);
xnor UO_366 (O_366,N_4984,N_4870);
nor UO_367 (O_367,N_4977,N_4896);
and UO_368 (O_368,N_4913,N_4950);
and UO_369 (O_369,N_4988,N_4861);
and UO_370 (O_370,N_4823,N_4838);
or UO_371 (O_371,N_4966,N_4908);
or UO_372 (O_372,N_4856,N_4864);
nor UO_373 (O_373,N_4894,N_4848);
and UO_374 (O_374,N_4877,N_4938);
nand UO_375 (O_375,N_4862,N_4960);
nor UO_376 (O_376,N_4897,N_4830);
or UO_377 (O_377,N_4910,N_4976);
and UO_378 (O_378,N_4859,N_4816);
and UO_379 (O_379,N_4909,N_4829);
nand UO_380 (O_380,N_4955,N_4846);
nand UO_381 (O_381,N_4821,N_4942);
nand UO_382 (O_382,N_4923,N_4870);
nor UO_383 (O_383,N_4803,N_4893);
and UO_384 (O_384,N_4819,N_4930);
nand UO_385 (O_385,N_4931,N_4803);
or UO_386 (O_386,N_4832,N_4989);
nor UO_387 (O_387,N_4801,N_4995);
and UO_388 (O_388,N_4933,N_4936);
nor UO_389 (O_389,N_4953,N_4837);
nor UO_390 (O_390,N_4931,N_4913);
nand UO_391 (O_391,N_4902,N_4849);
and UO_392 (O_392,N_4923,N_4974);
and UO_393 (O_393,N_4947,N_4873);
or UO_394 (O_394,N_4810,N_4873);
xor UO_395 (O_395,N_4912,N_4918);
or UO_396 (O_396,N_4927,N_4989);
nor UO_397 (O_397,N_4857,N_4992);
xor UO_398 (O_398,N_4823,N_4824);
and UO_399 (O_399,N_4833,N_4873);
or UO_400 (O_400,N_4865,N_4907);
nand UO_401 (O_401,N_4875,N_4954);
or UO_402 (O_402,N_4888,N_4920);
nor UO_403 (O_403,N_4959,N_4812);
or UO_404 (O_404,N_4933,N_4819);
and UO_405 (O_405,N_4841,N_4853);
and UO_406 (O_406,N_4974,N_4856);
xor UO_407 (O_407,N_4808,N_4881);
and UO_408 (O_408,N_4816,N_4899);
and UO_409 (O_409,N_4948,N_4882);
nand UO_410 (O_410,N_4815,N_4904);
nor UO_411 (O_411,N_4990,N_4983);
or UO_412 (O_412,N_4859,N_4858);
nor UO_413 (O_413,N_4929,N_4993);
nand UO_414 (O_414,N_4838,N_4937);
or UO_415 (O_415,N_4998,N_4881);
nor UO_416 (O_416,N_4837,N_4850);
nand UO_417 (O_417,N_4946,N_4974);
and UO_418 (O_418,N_4901,N_4920);
nor UO_419 (O_419,N_4873,N_4884);
nand UO_420 (O_420,N_4877,N_4810);
nor UO_421 (O_421,N_4864,N_4854);
nand UO_422 (O_422,N_4986,N_4841);
or UO_423 (O_423,N_4967,N_4901);
and UO_424 (O_424,N_4900,N_4816);
nand UO_425 (O_425,N_4907,N_4833);
or UO_426 (O_426,N_4974,N_4902);
nor UO_427 (O_427,N_4935,N_4879);
xor UO_428 (O_428,N_4809,N_4905);
and UO_429 (O_429,N_4827,N_4845);
nor UO_430 (O_430,N_4953,N_4957);
nand UO_431 (O_431,N_4963,N_4807);
and UO_432 (O_432,N_4893,N_4810);
nand UO_433 (O_433,N_4965,N_4862);
xnor UO_434 (O_434,N_4930,N_4904);
nand UO_435 (O_435,N_4929,N_4957);
nand UO_436 (O_436,N_4981,N_4852);
nor UO_437 (O_437,N_4945,N_4935);
nor UO_438 (O_438,N_4800,N_4807);
and UO_439 (O_439,N_4912,N_4954);
nand UO_440 (O_440,N_4846,N_4853);
xnor UO_441 (O_441,N_4800,N_4991);
and UO_442 (O_442,N_4885,N_4819);
and UO_443 (O_443,N_4911,N_4843);
or UO_444 (O_444,N_4961,N_4893);
nor UO_445 (O_445,N_4956,N_4853);
nor UO_446 (O_446,N_4970,N_4975);
nand UO_447 (O_447,N_4929,N_4819);
or UO_448 (O_448,N_4982,N_4816);
and UO_449 (O_449,N_4840,N_4918);
and UO_450 (O_450,N_4899,N_4855);
nand UO_451 (O_451,N_4829,N_4937);
or UO_452 (O_452,N_4983,N_4855);
and UO_453 (O_453,N_4977,N_4906);
or UO_454 (O_454,N_4981,N_4951);
and UO_455 (O_455,N_4958,N_4836);
or UO_456 (O_456,N_4852,N_4900);
and UO_457 (O_457,N_4902,N_4863);
and UO_458 (O_458,N_4952,N_4844);
or UO_459 (O_459,N_4930,N_4804);
or UO_460 (O_460,N_4998,N_4914);
and UO_461 (O_461,N_4876,N_4989);
or UO_462 (O_462,N_4909,N_4811);
xor UO_463 (O_463,N_4900,N_4899);
nor UO_464 (O_464,N_4813,N_4858);
nor UO_465 (O_465,N_4819,N_4986);
and UO_466 (O_466,N_4923,N_4947);
or UO_467 (O_467,N_4965,N_4885);
and UO_468 (O_468,N_4912,N_4858);
nor UO_469 (O_469,N_4842,N_4851);
nor UO_470 (O_470,N_4981,N_4833);
nand UO_471 (O_471,N_4944,N_4943);
xnor UO_472 (O_472,N_4968,N_4885);
and UO_473 (O_473,N_4947,N_4802);
nand UO_474 (O_474,N_4909,N_4813);
and UO_475 (O_475,N_4979,N_4960);
xor UO_476 (O_476,N_4800,N_4839);
nand UO_477 (O_477,N_4926,N_4979);
nand UO_478 (O_478,N_4833,N_4820);
nor UO_479 (O_479,N_4841,N_4842);
or UO_480 (O_480,N_4862,N_4820);
or UO_481 (O_481,N_4930,N_4801);
nand UO_482 (O_482,N_4943,N_4869);
xor UO_483 (O_483,N_4826,N_4876);
nand UO_484 (O_484,N_4809,N_4823);
or UO_485 (O_485,N_4870,N_4915);
or UO_486 (O_486,N_4865,N_4834);
xor UO_487 (O_487,N_4894,N_4932);
nor UO_488 (O_488,N_4856,N_4917);
or UO_489 (O_489,N_4920,N_4816);
or UO_490 (O_490,N_4992,N_4852);
nor UO_491 (O_491,N_4853,N_4879);
nand UO_492 (O_492,N_4997,N_4949);
or UO_493 (O_493,N_4824,N_4941);
nor UO_494 (O_494,N_4911,N_4998);
xor UO_495 (O_495,N_4825,N_4863);
nor UO_496 (O_496,N_4864,N_4960);
nand UO_497 (O_497,N_4828,N_4829);
and UO_498 (O_498,N_4932,N_4882);
and UO_499 (O_499,N_4876,N_4830);
nand UO_500 (O_500,N_4855,N_4965);
and UO_501 (O_501,N_4995,N_4909);
nand UO_502 (O_502,N_4868,N_4836);
nand UO_503 (O_503,N_4916,N_4877);
and UO_504 (O_504,N_4841,N_4893);
or UO_505 (O_505,N_4879,N_4819);
nor UO_506 (O_506,N_4891,N_4949);
or UO_507 (O_507,N_4931,N_4965);
nand UO_508 (O_508,N_4931,N_4852);
nor UO_509 (O_509,N_4991,N_4986);
nand UO_510 (O_510,N_4898,N_4836);
xnor UO_511 (O_511,N_4972,N_4910);
and UO_512 (O_512,N_4876,N_4945);
or UO_513 (O_513,N_4922,N_4806);
nor UO_514 (O_514,N_4881,N_4948);
nand UO_515 (O_515,N_4842,N_4847);
nand UO_516 (O_516,N_4853,N_4887);
and UO_517 (O_517,N_4845,N_4889);
and UO_518 (O_518,N_4900,N_4806);
or UO_519 (O_519,N_4889,N_4972);
or UO_520 (O_520,N_4972,N_4904);
and UO_521 (O_521,N_4827,N_4821);
and UO_522 (O_522,N_4960,N_4828);
or UO_523 (O_523,N_4911,N_4865);
nor UO_524 (O_524,N_4859,N_4997);
or UO_525 (O_525,N_4968,N_4872);
nor UO_526 (O_526,N_4928,N_4848);
nand UO_527 (O_527,N_4804,N_4834);
xor UO_528 (O_528,N_4947,N_4895);
nand UO_529 (O_529,N_4968,N_4843);
nand UO_530 (O_530,N_4886,N_4814);
nor UO_531 (O_531,N_4980,N_4823);
nor UO_532 (O_532,N_4958,N_4995);
or UO_533 (O_533,N_4887,N_4954);
xnor UO_534 (O_534,N_4939,N_4952);
or UO_535 (O_535,N_4932,N_4869);
nand UO_536 (O_536,N_4871,N_4827);
nand UO_537 (O_537,N_4876,N_4837);
or UO_538 (O_538,N_4863,N_4823);
xnor UO_539 (O_539,N_4993,N_4982);
or UO_540 (O_540,N_4856,N_4819);
xor UO_541 (O_541,N_4985,N_4898);
and UO_542 (O_542,N_4895,N_4991);
or UO_543 (O_543,N_4993,N_4801);
and UO_544 (O_544,N_4985,N_4827);
nand UO_545 (O_545,N_4998,N_4849);
or UO_546 (O_546,N_4870,N_4951);
xnor UO_547 (O_547,N_4885,N_4834);
or UO_548 (O_548,N_4841,N_4917);
nand UO_549 (O_549,N_4978,N_4880);
nor UO_550 (O_550,N_4915,N_4952);
nand UO_551 (O_551,N_4976,N_4992);
nor UO_552 (O_552,N_4863,N_4846);
or UO_553 (O_553,N_4847,N_4975);
and UO_554 (O_554,N_4911,N_4827);
nor UO_555 (O_555,N_4863,N_4964);
xor UO_556 (O_556,N_4847,N_4921);
and UO_557 (O_557,N_4840,N_4978);
or UO_558 (O_558,N_4968,N_4983);
nor UO_559 (O_559,N_4967,N_4875);
or UO_560 (O_560,N_4833,N_4944);
nand UO_561 (O_561,N_4943,N_4840);
nand UO_562 (O_562,N_4943,N_4921);
and UO_563 (O_563,N_4829,N_4863);
or UO_564 (O_564,N_4869,N_4818);
and UO_565 (O_565,N_4926,N_4810);
nand UO_566 (O_566,N_4803,N_4923);
xor UO_567 (O_567,N_4922,N_4890);
xnor UO_568 (O_568,N_4823,N_4843);
nand UO_569 (O_569,N_4872,N_4833);
or UO_570 (O_570,N_4954,N_4886);
and UO_571 (O_571,N_4905,N_4887);
nor UO_572 (O_572,N_4886,N_4893);
nor UO_573 (O_573,N_4879,N_4880);
nand UO_574 (O_574,N_4865,N_4932);
nand UO_575 (O_575,N_4837,N_4975);
nor UO_576 (O_576,N_4841,N_4963);
nor UO_577 (O_577,N_4990,N_4809);
nand UO_578 (O_578,N_4935,N_4813);
nand UO_579 (O_579,N_4871,N_4821);
nor UO_580 (O_580,N_4907,N_4871);
or UO_581 (O_581,N_4878,N_4957);
nor UO_582 (O_582,N_4919,N_4864);
nand UO_583 (O_583,N_4835,N_4884);
nand UO_584 (O_584,N_4999,N_4872);
nand UO_585 (O_585,N_4982,N_4853);
nand UO_586 (O_586,N_4834,N_4805);
nand UO_587 (O_587,N_4866,N_4859);
or UO_588 (O_588,N_4888,N_4912);
xor UO_589 (O_589,N_4946,N_4880);
or UO_590 (O_590,N_4877,N_4850);
and UO_591 (O_591,N_4995,N_4850);
nor UO_592 (O_592,N_4909,N_4902);
nor UO_593 (O_593,N_4912,N_4945);
and UO_594 (O_594,N_4820,N_4987);
nand UO_595 (O_595,N_4849,N_4949);
or UO_596 (O_596,N_4860,N_4891);
nor UO_597 (O_597,N_4802,N_4824);
nor UO_598 (O_598,N_4871,N_4941);
nor UO_599 (O_599,N_4931,N_4801);
and UO_600 (O_600,N_4839,N_4868);
or UO_601 (O_601,N_4976,N_4867);
xnor UO_602 (O_602,N_4944,N_4850);
and UO_603 (O_603,N_4962,N_4919);
nor UO_604 (O_604,N_4960,N_4868);
and UO_605 (O_605,N_4940,N_4923);
xor UO_606 (O_606,N_4863,N_4813);
nand UO_607 (O_607,N_4856,N_4963);
or UO_608 (O_608,N_4862,N_4993);
nand UO_609 (O_609,N_4967,N_4958);
nand UO_610 (O_610,N_4800,N_4939);
and UO_611 (O_611,N_4817,N_4974);
and UO_612 (O_612,N_4966,N_4838);
nor UO_613 (O_613,N_4801,N_4859);
or UO_614 (O_614,N_4918,N_4961);
nor UO_615 (O_615,N_4805,N_4969);
and UO_616 (O_616,N_4872,N_4859);
or UO_617 (O_617,N_4899,N_4981);
nor UO_618 (O_618,N_4939,N_4967);
nand UO_619 (O_619,N_4827,N_4999);
nor UO_620 (O_620,N_4958,N_4904);
or UO_621 (O_621,N_4953,N_4936);
or UO_622 (O_622,N_4944,N_4939);
nand UO_623 (O_623,N_4960,N_4978);
or UO_624 (O_624,N_4969,N_4870);
or UO_625 (O_625,N_4844,N_4890);
nand UO_626 (O_626,N_4873,N_4955);
and UO_627 (O_627,N_4848,N_4930);
nand UO_628 (O_628,N_4889,N_4943);
xnor UO_629 (O_629,N_4973,N_4887);
nor UO_630 (O_630,N_4882,N_4956);
and UO_631 (O_631,N_4866,N_4899);
and UO_632 (O_632,N_4906,N_4943);
and UO_633 (O_633,N_4981,N_4885);
or UO_634 (O_634,N_4848,N_4962);
and UO_635 (O_635,N_4976,N_4971);
and UO_636 (O_636,N_4943,N_4844);
and UO_637 (O_637,N_4977,N_4928);
or UO_638 (O_638,N_4968,N_4868);
and UO_639 (O_639,N_4988,N_4919);
or UO_640 (O_640,N_4808,N_4878);
nand UO_641 (O_641,N_4882,N_4846);
nor UO_642 (O_642,N_4955,N_4867);
and UO_643 (O_643,N_4951,N_4924);
nor UO_644 (O_644,N_4927,N_4895);
xnor UO_645 (O_645,N_4925,N_4914);
nand UO_646 (O_646,N_4816,N_4823);
xor UO_647 (O_647,N_4935,N_4824);
nor UO_648 (O_648,N_4950,N_4805);
and UO_649 (O_649,N_4887,N_4988);
or UO_650 (O_650,N_4904,N_4818);
nand UO_651 (O_651,N_4846,N_4862);
or UO_652 (O_652,N_4847,N_4917);
and UO_653 (O_653,N_4817,N_4903);
or UO_654 (O_654,N_4802,N_4897);
and UO_655 (O_655,N_4823,N_4987);
or UO_656 (O_656,N_4873,N_4811);
and UO_657 (O_657,N_4864,N_4866);
or UO_658 (O_658,N_4843,N_4815);
or UO_659 (O_659,N_4804,N_4833);
or UO_660 (O_660,N_4931,N_4834);
nor UO_661 (O_661,N_4949,N_4821);
or UO_662 (O_662,N_4983,N_4905);
or UO_663 (O_663,N_4823,N_4964);
or UO_664 (O_664,N_4810,N_4864);
and UO_665 (O_665,N_4914,N_4877);
or UO_666 (O_666,N_4886,N_4979);
or UO_667 (O_667,N_4969,N_4904);
or UO_668 (O_668,N_4876,N_4812);
nand UO_669 (O_669,N_4926,N_4998);
or UO_670 (O_670,N_4820,N_4874);
nand UO_671 (O_671,N_4931,N_4848);
nand UO_672 (O_672,N_4833,N_4819);
or UO_673 (O_673,N_4819,N_4928);
nand UO_674 (O_674,N_4918,N_4931);
nor UO_675 (O_675,N_4826,N_4915);
xor UO_676 (O_676,N_4804,N_4900);
nand UO_677 (O_677,N_4809,N_4804);
and UO_678 (O_678,N_4896,N_4860);
and UO_679 (O_679,N_4862,N_4878);
nand UO_680 (O_680,N_4997,N_4944);
and UO_681 (O_681,N_4808,N_4984);
or UO_682 (O_682,N_4958,N_4813);
nor UO_683 (O_683,N_4861,N_4936);
or UO_684 (O_684,N_4946,N_4861);
and UO_685 (O_685,N_4843,N_4963);
nand UO_686 (O_686,N_4933,N_4957);
and UO_687 (O_687,N_4958,N_4823);
nand UO_688 (O_688,N_4901,N_4877);
nor UO_689 (O_689,N_4990,N_4922);
and UO_690 (O_690,N_4975,N_4905);
nor UO_691 (O_691,N_4987,N_4897);
nand UO_692 (O_692,N_4995,N_4925);
xor UO_693 (O_693,N_4945,N_4878);
nand UO_694 (O_694,N_4890,N_4949);
or UO_695 (O_695,N_4863,N_4909);
or UO_696 (O_696,N_4986,N_4997);
nor UO_697 (O_697,N_4836,N_4893);
xnor UO_698 (O_698,N_4973,N_4904);
nand UO_699 (O_699,N_4841,N_4994);
and UO_700 (O_700,N_4949,N_4907);
or UO_701 (O_701,N_4802,N_4892);
xnor UO_702 (O_702,N_4822,N_4808);
nand UO_703 (O_703,N_4925,N_4831);
and UO_704 (O_704,N_4838,N_4929);
nand UO_705 (O_705,N_4830,N_4827);
nor UO_706 (O_706,N_4883,N_4943);
or UO_707 (O_707,N_4887,N_4841);
xor UO_708 (O_708,N_4952,N_4909);
or UO_709 (O_709,N_4960,N_4965);
and UO_710 (O_710,N_4989,N_4942);
nor UO_711 (O_711,N_4857,N_4833);
nand UO_712 (O_712,N_4955,N_4921);
or UO_713 (O_713,N_4802,N_4900);
nand UO_714 (O_714,N_4924,N_4936);
xnor UO_715 (O_715,N_4995,N_4827);
and UO_716 (O_716,N_4984,N_4955);
and UO_717 (O_717,N_4835,N_4882);
nand UO_718 (O_718,N_4891,N_4939);
and UO_719 (O_719,N_4998,N_4841);
or UO_720 (O_720,N_4892,N_4849);
and UO_721 (O_721,N_4802,N_4800);
nand UO_722 (O_722,N_4909,N_4869);
xor UO_723 (O_723,N_4919,N_4804);
or UO_724 (O_724,N_4920,N_4942);
and UO_725 (O_725,N_4857,N_4947);
or UO_726 (O_726,N_4945,N_4982);
nor UO_727 (O_727,N_4888,N_4915);
and UO_728 (O_728,N_4827,N_4948);
and UO_729 (O_729,N_4801,N_4851);
nand UO_730 (O_730,N_4997,N_4906);
or UO_731 (O_731,N_4877,N_4806);
nor UO_732 (O_732,N_4938,N_4921);
nor UO_733 (O_733,N_4804,N_4974);
nand UO_734 (O_734,N_4950,N_4894);
nor UO_735 (O_735,N_4826,N_4814);
and UO_736 (O_736,N_4933,N_4921);
nand UO_737 (O_737,N_4915,N_4828);
or UO_738 (O_738,N_4966,N_4810);
nor UO_739 (O_739,N_4977,N_4875);
xor UO_740 (O_740,N_4976,N_4948);
or UO_741 (O_741,N_4858,N_4803);
and UO_742 (O_742,N_4962,N_4822);
xor UO_743 (O_743,N_4886,N_4919);
or UO_744 (O_744,N_4971,N_4972);
xor UO_745 (O_745,N_4836,N_4999);
or UO_746 (O_746,N_4862,N_4904);
nand UO_747 (O_747,N_4868,N_4812);
and UO_748 (O_748,N_4854,N_4857);
or UO_749 (O_749,N_4915,N_4910);
nand UO_750 (O_750,N_4895,N_4925);
nand UO_751 (O_751,N_4941,N_4878);
nand UO_752 (O_752,N_4991,N_4950);
xnor UO_753 (O_753,N_4822,N_4925);
xnor UO_754 (O_754,N_4833,N_4939);
nand UO_755 (O_755,N_4869,N_4834);
nand UO_756 (O_756,N_4963,N_4846);
nor UO_757 (O_757,N_4888,N_4883);
xnor UO_758 (O_758,N_4936,N_4822);
and UO_759 (O_759,N_4960,N_4971);
nand UO_760 (O_760,N_4870,N_4975);
nand UO_761 (O_761,N_4894,N_4988);
nand UO_762 (O_762,N_4888,N_4928);
and UO_763 (O_763,N_4835,N_4902);
nor UO_764 (O_764,N_4800,N_4979);
xnor UO_765 (O_765,N_4962,N_4980);
nor UO_766 (O_766,N_4850,N_4967);
or UO_767 (O_767,N_4944,N_4851);
or UO_768 (O_768,N_4886,N_4839);
nor UO_769 (O_769,N_4999,N_4821);
or UO_770 (O_770,N_4823,N_4902);
or UO_771 (O_771,N_4806,N_4905);
or UO_772 (O_772,N_4815,N_4812);
or UO_773 (O_773,N_4824,N_4894);
nor UO_774 (O_774,N_4815,N_4960);
or UO_775 (O_775,N_4822,N_4994);
or UO_776 (O_776,N_4957,N_4874);
or UO_777 (O_777,N_4867,N_4856);
nor UO_778 (O_778,N_4873,N_4970);
and UO_779 (O_779,N_4804,N_4891);
xor UO_780 (O_780,N_4893,N_4978);
xor UO_781 (O_781,N_4941,N_4919);
xnor UO_782 (O_782,N_4814,N_4899);
or UO_783 (O_783,N_4825,N_4808);
nand UO_784 (O_784,N_4940,N_4884);
xor UO_785 (O_785,N_4840,N_4832);
nand UO_786 (O_786,N_4819,N_4827);
or UO_787 (O_787,N_4878,N_4908);
xnor UO_788 (O_788,N_4930,N_4866);
nor UO_789 (O_789,N_4973,N_4952);
nand UO_790 (O_790,N_4927,N_4967);
and UO_791 (O_791,N_4846,N_4866);
nand UO_792 (O_792,N_4800,N_4889);
nor UO_793 (O_793,N_4855,N_4882);
nand UO_794 (O_794,N_4842,N_4984);
and UO_795 (O_795,N_4833,N_4918);
nand UO_796 (O_796,N_4899,N_4818);
or UO_797 (O_797,N_4855,N_4809);
nor UO_798 (O_798,N_4860,N_4848);
and UO_799 (O_799,N_4845,N_4967);
xor UO_800 (O_800,N_4976,N_4811);
or UO_801 (O_801,N_4981,N_4937);
nor UO_802 (O_802,N_4969,N_4892);
xnor UO_803 (O_803,N_4907,N_4953);
or UO_804 (O_804,N_4942,N_4849);
nand UO_805 (O_805,N_4976,N_4800);
xor UO_806 (O_806,N_4926,N_4885);
nor UO_807 (O_807,N_4922,N_4893);
or UO_808 (O_808,N_4891,N_4968);
nand UO_809 (O_809,N_4882,N_4943);
xnor UO_810 (O_810,N_4842,N_4923);
xor UO_811 (O_811,N_4801,N_4836);
xor UO_812 (O_812,N_4960,N_4953);
nor UO_813 (O_813,N_4865,N_4954);
nand UO_814 (O_814,N_4936,N_4806);
nand UO_815 (O_815,N_4916,N_4936);
or UO_816 (O_816,N_4808,N_4805);
and UO_817 (O_817,N_4978,N_4853);
nand UO_818 (O_818,N_4962,N_4985);
xnor UO_819 (O_819,N_4914,N_4839);
and UO_820 (O_820,N_4930,N_4952);
and UO_821 (O_821,N_4993,N_4804);
xor UO_822 (O_822,N_4863,N_4908);
nor UO_823 (O_823,N_4935,N_4988);
or UO_824 (O_824,N_4966,N_4977);
xnor UO_825 (O_825,N_4970,N_4904);
nor UO_826 (O_826,N_4971,N_4905);
nand UO_827 (O_827,N_4817,N_4943);
or UO_828 (O_828,N_4835,N_4988);
nand UO_829 (O_829,N_4957,N_4927);
and UO_830 (O_830,N_4902,N_4815);
or UO_831 (O_831,N_4932,N_4988);
and UO_832 (O_832,N_4828,N_4874);
or UO_833 (O_833,N_4881,N_4944);
nor UO_834 (O_834,N_4935,N_4981);
and UO_835 (O_835,N_4836,N_4804);
and UO_836 (O_836,N_4803,N_4809);
nor UO_837 (O_837,N_4943,N_4856);
and UO_838 (O_838,N_4882,N_4944);
or UO_839 (O_839,N_4839,N_4893);
nor UO_840 (O_840,N_4906,N_4982);
or UO_841 (O_841,N_4849,N_4908);
and UO_842 (O_842,N_4880,N_4922);
nand UO_843 (O_843,N_4941,N_4951);
nand UO_844 (O_844,N_4852,N_4875);
nand UO_845 (O_845,N_4946,N_4993);
and UO_846 (O_846,N_4876,N_4900);
nand UO_847 (O_847,N_4930,N_4891);
or UO_848 (O_848,N_4925,N_4946);
or UO_849 (O_849,N_4879,N_4849);
nand UO_850 (O_850,N_4827,N_4813);
and UO_851 (O_851,N_4962,N_4881);
and UO_852 (O_852,N_4973,N_4989);
or UO_853 (O_853,N_4903,N_4844);
nor UO_854 (O_854,N_4928,N_4957);
and UO_855 (O_855,N_4807,N_4905);
nand UO_856 (O_856,N_4925,N_4862);
xnor UO_857 (O_857,N_4944,N_4898);
and UO_858 (O_858,N_4890,N_4859);
or UO_859 (O_859,N_4980,N_4821);
or UO_860 (O_860,N_4940,N_4951);
nor UO_861 (O_861,N_4813,N_4853);
or UO_862 (O_862,N_4964,N_4903);
nor UO_863 (O_863,N_4884,N_4820);
nand UO_864 (O_864,N_4881,N_4846);
and UO_865 (O_865,N_4918,N_4957);
nand UO_866 (O_866,N_4826,N_4896);
or UO_867 (O_867,N_4897,N_4995);
nor UO_868 (O_868,N_4830,N_4924);
xor UO_869 (O_869,N_4874,N_4931);
and UO_870 (O_870,N_4941,N_4879);
nand UO_871 (O_871,N_4895,N_4963);
and UO_872 (O_872,N_4994,N_4931);
xnor UO_873 (O_873,N_4958,N_4890);
nor UO_874 (O_874,N_4888,N_4809);
nand UO_875 (O_875,N_4822,N_4984);
nor UO_876 (O_876,N_4815,N_4821);
or UO_877 (O_877,N_4855,N_4903);
nand UO_878 (O_878,N_4918,N_4969);
and UO_879 (O_879,N_4826,N_4859);
or UO_880 (O_880,N_4881,N_4840);
and UO_881 (O_881,N_4802,N_4939);
xnor UO_882 (O_882,N_4954,N_4919);
or UO_883 (O_883,N_4962,N_4813);
nand UO_884 (O_884,N_4811,N_4860);
or UO_885 (O_885,N_4848,N_4879);
or UO_886 (O_886,N_4905,N_4800);
nand UO_887 (O_887,N_4981,N_4978);
nand UO_888 (O_888,N_4906,N_4846);
nor UO_889 (O_889,N_4946,N_4894);
xor UO_890 (O_890,N_4902,N_4976);
xnor UO_891 (O_891,N_4858,N_4942);
nor UO_892 (O_892,N_4912,N_4995);
nor UO_893 (O_893,N_4830,N_4874);
xor UO_894 (O_894,N_4919,N_4927);
or UO_895 (O_895,N_4805,N_4879);
and UO_896 (O_896,N_4978,N_4920);
and UO_897 (O_897,N_4888,N_4975);
nand UO_898 (O_898,N_4969,N_4875);
nor UO_899 (O_899,N_4958,N_4930);
nand UO_900 (O_900,N_4951,N_4947);
or UO_901 (O_901,N_4808,N_4999);
nor UO_902 (O_902,N_4921,N_4966);
and UO_903 (O_903,N_4988,N_4985);
nand UO_904 (O_904,N_4811,N_4894);
nor UO_905 (O_905,N_4946,N_4863);
and UO_906 (O_906,N_4990,N_4830);
nand UO_907 (O_907,N_4947,N_4833);
nand UO_908 (O_908,N_4878,N_4950);
and UO_909 (O_909,N_4906,N_4963);
or UO_910 (O_910,N_4872,N_4892);
nand UO_911 (O_911,N_4877,N_4933);
nor UO_912 (O_912,N_4894,N_4922);
or UO_913 (O_913,N_4850,N_4802);
or UO_914 (O_914,N_4923,N_4825);
and UO_915 (O_915,N_4869,N_4862);
nand UO_916 (O_916,N_4909,N_4861);
and UO_917 (O_917,N_4868,N_4900);
nor UO_918 (O_918,N_4891,N_4933);
and UO_919 (O_919,N_4807,N_4869);
or UO_920 (O_920,N_4961,N_4912);
or UO_921 (O_921,N_4923,N_4989);
and UO_922 (O_922,N_4926,N_4808);
and UO_923 (O_923,N_4993,N_4858);
or UO_924 (O_924,N_4851,N_4918);
nor UO_925 (O_925,N_4848,N_4831);
nor UO_926 (O_926,N_4953,N_4809);
and UO_927 (O_927,N_4800,N_4985);
nand UO_928 (O_928,N_4880,N_4931);
and UO_929 (O_929,N_4818,N_4946);
nand UO_930 (O_930,N_4898,N_4851);
or UO_931 (O_931,N_4964,N_4949);
and UO_932 (O_932,N_4831,N_4998);
xnor UO_933 (O_933,N_4906,N_4817);
nor UO_934 (O_934,N_4911,N_4924);
nand UO_935 (O_935,N_4873,N_4894);
or UO_936 (O_936,N_4840,N_4989);
nand UO_937 (O_937,N_4897,N_4872);
nand UO_938 (O_938,N_4952,N_4962);
nand UO_939 (O_939,N_4942,N_4972);
and UO_940 (O_940,N_4872,N_4955);
and UO_941 (O_941,N_4906,N_4859);
nor UO_942 (O_942,N_4885,N_4870);
or UO_943 (O_943,N_4843,N_4931);
nor UO_944 (O_944,N_4992,N_4822);
and UO_945 (O_945,N_4910,N_4834);
nor UO_946 (O_946,N_4898,N_4864);
or UO_947 (O_947,N_4818,N_4933);
nand UO_948 (O_948,N_4850,N_4943);
and UO_949 (O_949,N_4951,N_4820);
and UO_950 (O_950,N_4941,N_4848);
or UO_951 (O_951,N_4993,N_4859);
nor UO_952 (O_952,N_4941,N_4954);
nor UO_953 (O_953,N_4801,N_4999);
or UO_954 (O_954,N_4890,N_4806);
and UO_955 (O_955,N_4956,N_4942);
nand UO_956 (O_956,N_4916,N_4876);
nand UO_957 (O_957,N_4939,N_4920);
nor UO_958 (O_958,N_4820,N_4914);
nand UO_959 (O_959,N_4985,N_4983);
or UO_960 (O_960,N_4952,N_4841);
xor UO_961 (O_961,N_4897,N_4857);
nor UO_962 (O_962,N_4899,N_4939);
nor UO_963 (O_963,N_4890,N_4906);
or UO_964 (O_964,N_4900,N_4924);
xnor UO_965 (O_965,N_4858,N_4896);
xor UO_966 (O_966,N_4990,N_4924);
and UO_967 (O_967,N_4919,N_4938);
or UO_968 (O_968,N_4948,N_4932);
nand UO_969 (O_969,N_4905,N_4995);
and UO_970 (O_970,N_4986,N_4927);
xnor UO_971 (O_971,N_4845,N_4820);
nor UO_972 (O_972,N_4854,N_4917);
nor UO_973 (O_973,N_4829,N_4917);
or UO_974 (O_974,N_4915,N_4840);
nor UO_975 (O_975,N_4903,N_4894);
nor UO_976 (O_976,N_4816,N_4952);
nand UO_977 (O_977,N_4847,N_4815);
or UO_978 (O_978,N_4906,N_4919);
and UO_979 (O_979,N_4851,N_4863);
and UO_980 (O_980,N_4970,N_4847);
nand UO_981 (O_981,N_4979,N_4989);
or UO_982 (O_982,N_4924,N_4817);
and UO_983 (O_983,N_4851,N_4914);
nor UO_984 (O_984,N_4808,N_4934);
nor UO_985 (O_985,N_4992,N_4974);
and UO_986 (O_986,N_4897,N_4819);
nor UO_987 (O_987,N_4947,N_4956);
nor UO_988 (O_988,N_4966,N_4824);
nand UO_989 (O_989,N_4861,N_4977);
nor UO_990 (O_990,N_4898,N_4894);
xor UO_991 (O_991,N_4855,N_4996);
nor UO_992 (O_992,N_4933,N_4861);
nand UO_993 (O_993,N_4976,N_4866);
and UO_994 (O_994,N_4995,N_4953);
or UO_995 (O_995,N_4926,N_4802);
and UO_996 (O_996,N_4925,N_4934);
nand UO_997 (O_997,N_4867,N_4987);
nor UO_998 (O_998,N_4865,N_4995);
nand UO_999 (O_999,N_4852,N_4841);
endmodule