module basic_750_5000_1000_25_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_551,In_590);
nand U1 (N_1,In_78,In_416);
nor U2 (N_2,In_707,In_253);
xnor U3 (N_3,In_219,In_576);
nor U4 (N_4,In_43,In_587);
or U5 (N_5,In_380,In_242);
nand U6 (N_6,In_695,In_621);
nor U7 (N_7,In_152,In_421);
or U8 (N_8,In_381,In_641);
or U9 (N_9,In_136,In_492);
or U10 (N_10,In_59,In_368);
nand U11 (N_11,In_203,In_544);
and U12 (N_12,In_573,In_265);
or U13 (N_13,In_190,In_511);
and U14 (N_14,In_16,In_288);
nor U15 (N_15,In_211,In_462);
or U16 (N_16,In_655,In_8);
or U17 (N_17,In_575,In_88);
nor U18 (N_18,In_720,In_128);
or U19 (N_19,In_521,In_374);
nor U20 (N_20,In_310,In_729);
or U21 (N_21,In_578,In_686);
and U22 (N_22,In_391,In_650);
nor U23 (N_23,In_33,In_27);
or U24 (N_24,In_486,In_640);
and U25 (N_25,In_224,In_627);
and U26 (N_26,In_107,In_550);
and U27 (N_27,In_630,In_722);
and U28 (N_28,In_83,In_713);
nor U29 (N_29,In_647,In_563);
or U30 (N_30,In_559,In_495);
and U31 (N_31,In_532,In_217);
or U32 (N_32,In_631,In_681);
nand U33 (N_33,In_129,In_565);
or U34 (N_34,In_212,In_234);
nor U35 (N_35,In_547,In_102);
or U36 (N_36,In_39,In_562);
and U37 (N_37,In_398,In_501);
and U38 (N_38,In_320,In_85);
nand U39 (N_39,In_184,In_618);
nor U40 (N_40,In_719,In_425);
nor U41 (N_41,In_475,In_449);
or U42 (N_42,In_422,In_610);
nand U43 (N_43,In_46,In_245);
or U44 (N_44,In_622,In_546);
and U45 (N_45,In_635,In_543);
nor U46 (N_46,In_468,In_185);
and U47 (N_47,In_336,In_728);
and U48 (N_48,In_510,In_51);
nor U49 (N_49,In_384,In_196);
nor U50 (N_50,In_639,In_315);
or U51 (N_51,In_549,In_414);
nand U52 (N_52,In_92,In_259);
nand U53 (N_53,In_662,In_4);
nand U54 (N_54,In_30,In_322);
nand U55 (N_55,In_619,In_395);
and U56 (N_56,In_418,In_178);
and U57 (N_57,In_527,In_123);
and U58 (N_58,In_7,In_612);
or U59 (N_59,In_36,In_68);
nor U60 (N_60,In_47,In_577);
or U61 (N_61,In_280,In_17);
nand U62 (N_62,In_144,In_323);
or U63 (N_63,In_574,In_455);
nor U64 (N_64,In_67,In_300);
and U65 (N_65,In_285,In_21);
or U66 (N_66,In_114,In_350);
or U67 (N_67,In_167,In_172);
xnor U68 (N_68,In_633,In_493);
and U69 (N_69,In_660,In_693);
and U70 (N_70,In_198,In_415);
or U71 (N_71,In_471,In_403);
and U72 (N_72,In_731,In_487);
or U73 (N_73,In_634,In_221);
nor U74 (N_74,In_72,In_656);
nor U75 (N_75,In_733,In_554);
or U76 (N_76,In_62,In_314);
nor U77 (N_77,In_286,In_588);
nand U78 (N_78,In_456,In_63);
nand U79 (N_79,In_716,In_537);
and U80 (N_80,In_149,In_90);
nor U81 (N_81,In_103,In_111);
and U82 (N_82,In_75,In_266);
or U83 (N_83,In_683,In_239);
nor U84 (N_84,In_268,In_397);
or U85 (N_85,In_741,In_155);
nor U86 (N_86,In_673,In_124);
and U87 (N_87,In_561,In_235);
nor U88 (N_88,In_626,In_735);
nand U89 (N_89,In_324,In_271);
nor U90 (N_90,In_176,In_372);
nor U91 (N_91,In_140,In_187);
and U92 (N_92,In_552,In_31);
nor U93 (N_93,In_296,In_685);
or U94 (N_94,In_709,In_290);
or U95 (N_95,In_512,In_344);
nand U96 (N_96,In_18,In_12);
nand U97 (N_97,In_520,In_137);
and U98 (N_98,In_441,In_363);
nand U99 (N_99,In_367,In_246);
or U100 (N_100,In_452,In_649);
or U101 (N_101,In_451,In_213);
or U102 (N_102,In_230,In_579);
nor U103 (N_103,In_645,In_747);
and U104 (N_104,In_122,In_620);
nand U105 (N_105,In_585,In_566);
or U106 (N_106,In_702,In_2);
and U107 (N_107,In_653,In_156);
xor U108 (N_108,In_465,In_704);
xnor U109 (N_109,In_329,In_121);
nand U110 (N_110,In_688,In_319);
nor U111 (N_111,In_41,In_96);
nand U112 (N_112,In_526,In_179);
or U113 (N_113,In_346,In_229);
and U114 (N_114,In_723,In_478);
nand U115 (N_115,In_423,In_608);
nor U116 (N_116,In_298,In_643);
and U117 (N_117,In_360,In_24);
or U118 (N_118,In_87,In_95);
or U119 (N_119,In_6,In_202);
nand U120 (N_120,In_584,In_556);
nor U121 (N_121,In_613,In_504);
or U122 (N_122,In_283,In_375);
nand U123 (N_123,In_654,In_560);
nor U124 (N_124,In_19,In_316);
and U125 (N_125,In_736,In_602);
nand U126 (N_126,In_49,In_555);
or U127 (N_127,In_480,In_146);
nand U128 (N_128,In_651,In_724);
or U129 (N_129,In_175,In_516);
and U130 (N_130,In_533,In_77);
nor U131 (N_131,In_37,In_58);
nor U132 (N_132,In_714,In_71);
or U133 (N_133,In_409,In_210);
nor U134 (N_134,In_302,In_226);
nand U135 (N_135,In_382,In_601);
nand U136 (N_136,In_410,In_636);
or U137 (N_137,In_181,In_447);
nor U138 (N_138,In_498,In_74);
or U139 (N_139,In_306,In_396);
or U140 (N_140,In_255,In_89);
nor U141 (N_141,In_223,In_592);
nor U142 (N_142,In_529,In_50);
nand U143 (N_143,In_594,In_483);
nor U144 (N_144,In_494,In_154);
nor U145 (N_145,In_503,In_488);
or U146 (N_146,In_118,In_250);
nand U147 (N_147,In_275,In_484);
nand U148 (N_148,In_477,In_466);
and U149 (N_149,In_523,In_605);
or U150 (N_150,In_125,In_744);
nand U151 (N_151,In_370,In_308);
nand U152 (N_152,In_304,In_330);
or U153 (N_153,In_680,In_227);
or U154 (N_154,In_426,In_514);
and U155 (N_155,In_177,In_703);
and U156 (N_156,In_277,In_419);
nor U157 (N_157,In_401,In_109);
and U158 (N_158,In_628,In_117);
nor U159 (N_159,In_343,In_669);
or U160 (N_160,In_359,In_317);
or U161 (N_161,In_473,In_611);
nor U162 (N_162,In_35,In_60);
nand U163 (N_163,In_267,In_127);
and U164 (N_164,In_734,In_205);
or U165 (N_165,In_200,In_215);
nand U166 (N_166,In_366,In_385);
nor U167 (N_167,In_305,In_434);
nor U168 (N_168,In_11,In_119);
nor U169 (N_169,In_97,In_355);
nor U170 (N_170,In_263,In_538);
nand U171 (N_171,In_345,In_690);
and U172 (N_172,In_721,In_297);
nor U173 (N_173,In_105,In_699);
nor U174 (N_174,In_361,In_476);
nor U175 (N_175,In_580,In_134);
nand U176 (N_176,In_353,In_251);
nor U177 (N_177,In_629,In_364);
nor U178 (N_178,In_675,In_5);
or U179 (N_179,In_739,In_28);
or U180 (N_180,In_689,In_38);
or U181 (N_181,In_57,In_571);
nor U182 (N_182,In_108,In_616);
and U183 (N_183,In_338,In_489);
or U184 (N_184,In_670,In_726);
and U185 (N_185,In_417,In_497);
or U186 (N_186,In_727,In_159);
and U187 (N_187,In_48,In_65);
nor U188 (N_188,In_666,In_564);
nor U189 (N_189,In_740,In_593);
or U190 (N_190,In_749,In_443);
or U191 (N_191,In_600,In_94);
nor U192 (N_192,In_53,In_165);
or U193 (N_193,In_248,In_517);
and U194 (N_194,In_148,In_171);
nor U195 (N_195,In_665,In_141);
nor U196 (N_196,In_183,In_524);
or U197 (N_197,In_365,In_379);
and U198 (N_198,In_318,In_499);
and U199 (N_199,In_599,In_191);
and U200 (N_200,In_428,N_161);
nor U201 (N_201,In_143,N_11);
nor U202 (N_202,In_104,In_79);
and U203 (N_203,In_507,In_272);
and U204 (N_204,N_30,N_134);
and U205 (N_205,In_151,In_404);
nand U206 (N_206,N_184,In_525);
or U207 (N_207,N_125,In_204);
nand U208 (N_208,N_90,N_28);
nand U209 (N_209,In_264,N_182);
and U210 (N_210,In_101,In_192);
or U211 (N_211,N_64,In_201);
and U212 (N_212,In_70,In_333);
and U213 (N_213,In_687,In_392);
nor U214 (N_214,In_73,N_103);
or U215 (N_215,In_238,In_188);
and U216 (N_216,In_362,In_531);
nor U217 (N_217,In_553,In_725);
nand U218 (N_218,N_13,In_112);
nor U219 (N_219,N_114,In_182);
nor U220 (N_220,N_129,N_15);
nand U221 (N_221,N_126,In_168);
and U222 (N_222,In_682,N_169);
nand U223 (N_223,In_189,In_389);
nand U224 (N_224,In_158,In_113);
nor U225 (N_225,In_0,N_46);
and U226 (N_226,In_26,In_712);
and U227 (N_227,N_69,In_13);
nor U228 (N_228,N_45,In_442);
nand U229 (N_229,In_160,In_157);
or U230 (N_230,In_717,In_369);
or U231 (N_231,In_312,N_7);
nor U232 (N_232,In_303,N_22);
nor U233 (N_233,In_287,In_698);
and U234 (N_234,In_412,N_74);
or U235 (N_235,In_332,In_371);
and U236 (N_236,N_199,In_742);
and U237 (N_237,In_357,In_582);
nor U238 (N_238,N_20,In_745);
nor U239 (N_239,In_490,In_354);
or U240 (N_240,N_44,In_193);
and U241 (N_241,In_76,In_249);
nand U242 (N_242,In_429,N_140);
nand U243 (N_243,N_9,In_66);
nor U244 (N_244,N_154,In_174);
or U245 (N_245,N_151,N_139);
and U246 (N_246,In_276,In_294);
nor U247 (N_247,In_383,N_73);
nand U248 (N_248,In_513,In_260);
nor U249 (N_249,In_433,In_678);
and U250 (N_250,In_100,N_91);
nor U251 (N_251,In_539,In_659);
nand U252 (N_252,In_166,In_82);
nand U253 (N_253,N_93,In_597);
and U254 (N_254,N_119,N_50);
nor U255 (N_255,In_32,In_625);
or U256 (N_256,N_148,In_390);
nor U257 (N_257,In_252,In_289);
and U258 (N_258,In_56,N_51);
nor U259 (N_259,In_679,N_5);
or U260 (N_260,N_66,In_132);
or U261 (N_261,In_91,In_534);
or U262 (N_262,In_522,N_198);
or U263 (N_263,In_646,In_110);
and U264 (N_264,N_42,In_197);
nor U265 (N_265,N_94,In_233);
nor U266 (N_266,In_106,In_671);
or U267 (N_267,In_377,In_29);
nor U268 (N_268,N_95,N_56);
nand U269 (N_269,In_470,In_23);
nor U270 (N_270,In_748,N_128);
and U271 (N_271,In_301,In_307);
or U272 (N_272,N_52,N_40);
or U273 (N_273,In_325,In_667);
xor U274 (N_274,In_505,In_131);
or U275 (N_275,N_197,In_461);
or U276 (N_276,In_269,In_591);
and U277 (N_277,In_10,In_358);
or U278 (N_278,In_460,In_341);
nand U279 (N_279,N_192,N_43);
nand U280 (N_280,In_491,In_14);
nand U281 (N_281,In_194,N_160);
nor U282 (N_282,In_623,N_152);
nand U283 (N_283,In_430,N_144);
or U284 (N_284,In_254,In_42);
nor U285 (N_285,In_342,In_706);
and U286 (N_286,N_171,In_321);
nor U287 (N_287,N_36,In_145);
and U288 (N_288,In_339,In_262);
nor U289 (N_289,In_274,N_78);
nor U290 (N_290,N_84,In_278);
or U291 (N_291,N_17,In_161);
nand U292 (N_292,In_677,In_220);
and U293 (N_293,In_98,In_347);
or U294 (N_294,In_737,In_232);
and U295 (N_295,In_411,N_65);
or U296 (N_296,N_138,In_438);
nor U297 (N_297,N_135,In_420);
and U298 (N_298,N_32,In_54);
nor U299 (N_299,In_482,N_88);
nand U300 (N_300,N_118,N_54);
nand U301 (N_301,In_93,N_29);
and U302 (N_302,In_258,In_676);
nor U303 (N_303,N_120,In_479);
and U304 (N_304,In_530,In_405);
and U305 (N_305,N_166,N_131);
and U306 (N_306,In_500,In_440);
or U307 (N_307,In_694,N_179);
and U308 (N_308,In_394,In_572);
nor U309 (N_309,N_164,N_193);
nand U310 (N_310,N_153,N_31);
and U311 (N_311,In_351,In_139);
or U312 (N_312,N_57,N_61);
nor U313 (N_313,N_147,N_85);
and U314 (N_314,In_708,In_515);
nand U315 (N_315,In_214,In_373);
and U316 (N_316,N_106,In_454);
and U317 (N_317,N_39,In_496);
or U318 (N_318,N_8,In_206);
nor U319 (N_319,In_664,N_23);
xnor U320 (N_320,In_697,In_349);
or U321 (N_321,In_569,N_136);
nand U322 (N_322,In_474,In_299);
and U323 (N_323,N_75,In_672);
or U324 (N_324,In_446,N_24);
or U325 (N_325,N_187,In_528);
or U326 (N_326,N_108,In_186);
and U327 (N_327,N_77,N_48);
and U328 (N_328,In_209,N_18);
nand U329 (N_329,In_445,In_457);
nor U330 (N_330,In_45,In_352);
and U331 (N_331,In_604,N_109);
nand U332 (N_332,N_175,In_1);
or U333 (N_333,N_14,In_624);
and U334 (N_334,N_63,In_481);
nor U335 (N_335,In_746,N_124);
and U336 (N_336,In_309,In_684);
or U337 (N_337,In_170,N_1);
nand U338 (N_338,In_348,N_71);
or U339 (N_339,N_37,N_68);
nand U340 (N_340,N_137,N_27);
and U341 (N_341,In_164,In_715);
nor U342 (N_342,N_185,N_186);
or U343 (N_343,N_34,In_328);
and U344 (N_344,N_33,In_459);
or U345 (N_345,N_2,In_52);
or U346 (N_346,N_81,In_116);
nor U347 (N_347,In_244,In_437);
and U348 (N_348,In_658,N_188);
or U349 (N_349,In_55,In_293);
nand U350 (N_350,N_16,In_406);
nand U351 (N_351,In_64,N_49);
nand U352 (N_352,In_216,In_463);
nand U353 (N_353,In_282,In_558);
or U354 (N_354,In_701,In_568);
or U355 (N_355,In_25,In_222);
or U356 (N_356,In_400,N_190);
and U357 (N_357,In_652,In_115);
nand U358 (N_358,N_150,N_26);
xor U359 (N_359,N_82,N_10);
and U360 (N_360,In_542,In_663);
and U361 (N_361,N_180,In_540);
nor U362 (N_362,N_107,N_189);
and U363 (N_363,In_256,In_444);
and U364 (N_364,In_617,In_387);
nand U365 (N_365,N_132,In_3);
and U366 (N_366,N_181,In_581);
and U367 (N_367,N_174,In_408);
nor U368 (N_368,In_609,N_62);
or U369 (N_369,N_127,In_133);
or U370 (N_370,In_292,In_44);
nand U371 (N_371,In_509,In_453);
and U372 (N_372,N_110,In_270);
and U373 (N_373,In_502,In_218);
nand U374 (N_374,N_163,In_291);
and U375 (N_375,In_356,N_89);
nor U376 (N_376,In_386,N_162);
nand U377 (N_377,In_138,N_142);
nand U378 (N_378,N_172,In_402);
and U379 (N_379,In_632,In_150);
or U380 (N_380,N_97,In_541);
or U381 (N_381,N_53,N_72);
or U382 (N_382,In_674,In_261);
and U383 (N_383,N_59,In_86);
nor U384 (N_384,N_92,In_80);
or U385 (N_385,In_436,In_464);
and U386 (N_386,N_111,In_126);
nor U387 (N_387,In_467,In_432);
nor U388 (N_388,In_519,N_123);
or U389 (N_389,In_603,N_99);
nand U390 (N_390,N_194,In_180);
and U391 (N_391,In_732,N_167);
nor U392 (N_392,N_98,In_506);
or U393 (N_393,In_334,In_661);
and U394 (N_394,In_710,N_155);
and U395 (N_395,N_47,In_273);
and U396 (N_396,N_146,In_135);
nor U397 (N_397,In_153,In_163);
nor U398 (N_398,In_583,In_606);
nand U399 (N_399,In_730,N_101);
or U400 (N_400,N_311,N_223);
and U401 (N_401,In_130,N_157);
or U402 (N_402,In_705,N_275);
and U403 (N_403,N_254,N_266);
or U404 (N_404,N_242,In_69);
nor U405 (N_405,N_366,N_290);
and U406 (N_406,N_219,N_396);
and U407 (N_407,N_307,In_34);
nor U408 (N_408,N_390,N_116);
or U409 (N_409,N_241,N_331);
nand U410 (N_410,N_381,In_424);
or U411 (N_411,In_692,N_240);
nor U412 (N_412,In_120,N_112);
nor U413 (N_413,In_536,N_354);
or U414 (N_414,In_340,In_243);
nand U415 (N_415,N_38,N_363);
nor U416 (N_416,N_215,In_240);
or U417 (N_417,In_399,In_648);
or U418 (N_418,N_225,N_156);
and U419 (N_419,N_370,In_570);
nor U420 (N_420,N_200,N_121);
or U421 (N_421,N_306,N_228);
nand U422 (N_422,N_352,N_60);
nor U423 (N_423,N_83,N_280);
nand U424 (N_424,In_508,N_268);
nand U425 (N_425,N_105,N_221);
nor U426 (N_426,In_208,In_435);
nor U427 (N_427,N_312,N_207);
nor U428 (N_428,N_329,N_392);
and U429 (N_429,N_227,N_149);
or U430 (N_430,N_388,N_348);
and U431 (N_431,N_378,N_364);
nand U432 (N_432,N_335,In_607);
nor U433 (N_433,N_379,N_230);
nor U434 (N_434,N_293,In_22);
and U435 (N_435,N_372,N_231);
or U436 (N_436,N_353,N_310);
nor U437 (N_437,N_218,N_4);
nand U438 (N_438,N_359,N_346);
and U439 (N_439,N_130,In_40);
nand U440 (N_440,N_308,N_96);
or U441 (N_441,N_236,N_278);
xnor U442 (N_442,N_58,In_598);
and U443 (N_443,In_545,In_431);
or U444 (N_444,N_229,N_341);
or U445 (N_445,N_260,N_70);
and U446 (N_446,N_86,N_334);
and U447 (N_447,N_100,N_177);
or U448 (N_448,N_286,N_232);
and U449 (N_449,In_472,In_195);
and U450 (N_450,N_380,N_234);
and U451 (N_451,N_210,In_326);
and U452 (N_452,N_303,N_371);
or U453 (N_453,In_596,N_355);
nor U454 (N_454,N_249,N_327);
xor U455 (N_455,N_222,N_226);
or U456 (N_456,In_84,In_279);
and U457 (N_457,In_331,N_284);
nor U458 (N_458,N_3,N_339);
nor U459 (N_459,N_253,N_330);
and U460 (N_460,N_321,N_316);
or U461 (N_461,N_237,In_376);
nand U462 (N_462,In_99,N_296);
nor U463 (N_463,In_311,In_20);
and U464 (N_464,N_376,N_272);
or U465 (N_465,In_548,N_235);
nand U466 (N_466,N_333,N_248);
nand U467 (N_467,In_237,In_81);
nand U468 (N_468,N_143,N_269);
or U469 (N_469,In_589,N_305);
nand U470 (N_470,N_12,N_292);
and U471 (N_471,In_313,In_615);
nor U472 (N_472,In_327,N_347);
nor U473 (N_473,N_387,N_337);
or U474 (N_474,N_250,N_158);
nand U475 (N_475,N_19,In_257);
and U476 (N_476,In_162,N_238);
and U477 (N_477,N_313,N_368);
nand U478 (N_478,N_202,N_239);
and U479 (N_479,In_595,N_67);
nor U480 (N_480,In_284,N_297);
nand U481 (N_481,N_314,In_696);
or U482 (N_482,N_277,In_567);
nor U483 (N_483,N_271,N_393);
nor U484 (N_484,N_104,N_183);
and U485 (N_485,N_395,In_557);
nor U486 (N_486,N_35,N_345);
or U487 (N_487,N_324,In_711);
or U488 (N_488,N_115,In_450);
and U489 (N_489,N_398,N_246);
and U490 (N_490,In_407,In_718);
nand U491 (N_491,N_279,N_386);
nand U492 (N_492,N_384,N_176);
or U493 (N_493,In_413,N_141);
and U494 (N_494,N_343,N_385);
nand U495 (N_495,N_288,N_282);
or U496 (N_496,N_389,N_394);
nand U497 (N_497,N_102,N_211);
nor U498 (N_498,N_80,N_342);
or U499 (N_499,N_256,N_262);
nor U500 (N_500,N_257,In_614);
and U501 (N_501,N_217,N_283);
and U502 (N_502,In_295,In_335);
xnor U503 (N_503,N_261,N_133);
or U504 (N_504,In_378,N_325);
or U505 (N_505,In_469,N_328);
nor U506 (N_506,N_322,N_323);
nor U507 (N_507,N_213,N_203);
or U508 (N_508,In_743,N_76);
nor U509 (N_509,N_309,In_637);
and U510 (N_510,In_439,N_270);
and U511 (N_511,N_360,N_205);
or U512 (N_512,N_274,N_245);
nand U513 (N_513,N_168,N_373);
nand U514 (N_514,N_117,In_15);
nor U515 (N_515,N_300,N_291);
xor U516 (N_516,In_231,N_145);
or U517 (N_517,N_170,N_289);
nand U518 (N_518,N_191,In_485);
nor U519 (N_519,N_273,N_209);
and U520 (N_520,N_263,N_336);
nor U521 (N_521,N_369,N_173);
nor U522 (N_522,N_294,N_87);
or U523 (N_523,N_251,N_326);
or U524 (N_524,N_113,In_207);
nor U525 (N_525,N_351,N_201);
or U526 (N_526,N_6,N_382);
nor U527 (N_527,N_255,N_344);
nor U528 (N_528,In_642,In_586);
or U529 (N_529,N_41,N_358);
and U530 (N_530,N_295,N_302);
and U531 (N_531,N_259,N_374);
and U532 (N_532,In_9,N_315);
nand U533 (N_533,In_61,N_247);
nor U534 (N_534,N_122,In_638);
or U535 (N_535,N_233,N_320);
nor U536 (N_536,In_281,In_142);
or U537 (N_537,N_178,N_264);
and U538 (N_538,N_350,N_244);
nor U539 (N_539,N_397,N_281);
nor U540 (N_540,In_199,N_267);
or U541 (N_541,N_55,In_427);
or U542 (N_542,N_224,In_458);
or U543 (N_543,In_228,N_204);
nor U544 (N_544,In_225,N_214);
or U545 (N_545,In_691,N_332);
or U546 (N_546,N_79,N_206);
nor U547 (N_547,In_644,N_276);
nand U548 (N_548,N_159,In_448);
and U549 (N_549,N_216,N_298);
nand U550 (N_550,N_195,N_304);
or U551 (N_551,N_208,N_299);
or U552 (N_552,N_319,N_252);
and U553 (N_553,In_668,N_367);
nor U554 (N_554,N_258,N_375);
and U555 (N_555,N_356,N_165);
and U556 (N_556,N_317,N_301);
nor U557 (N_557,N_361,In_738);
and U558 (N_558,N_287,In_247);
nand U559 (N_559,N_212,In_393);
nor U560 (N_560,In_241,N_0);
nor U561 (N_561,In_657,N_25);
or U562 (N_562,N_318,N_349);
or U563 (N_563,N_340,In_147);
or U564 (N_564,In_337,N_391);
and U565 (N_565,N_220,N_21);
and U566 (N_566,In_700,N_285);
or U567 (N_567,In_173,N_383);
nand U568 (N_568,N_265,N_357);
nand U569 (N_569,In_169,N_362);
and U570 (N_570,N_377,N_196);
nor U571 (N_571,N_399,In_535);
nor U572 (N_572,N_338,N_365);
nand U573 (N_573,In_236,N_243);
nor U574 (N_574,In_518,In_388);
and U575 (N_575,N_385,N_360);
nor U576 (N_576,In_508,In_228);
or U577 (N_577,In_705,In_147);
and U578 (N_578,N_236,N_268);
or U579 (N_579,In_147,N_79);
and U580 (N_580,N_318,N_203);
nor U581 (N_581,N_210,N_122);
and U582 (N_582,N_364,In_327);
nor U583 (N_583,In_326,N_313);
nor U584 (N_584,N_225,N_289);
and U585 (N_585,In_378,N_265);
nor U586 (N_586,N_60,N_121);
nor U587 (N_587,N_113,N_143);
and U588 (N_588,N_12,N_259);
or U589 (N_589,N_149,N_67);
nand U590 (N_590,N_374,N_115);
nand U591 (N_591,In_743,N_387);
nand U592 (N_592,N_385,N_183);
nand U593 (N_593,In_637,N_390);
nor U594 (N_594,N_96,N_345);
nand U595 (N_595,In_169,N_218);
nor U596 (N_596,N_269,N_260);
or U597 (N_597,N_260,In_284);
nor U598 (N_598,N_353,N_105);
and U599 (N_599,N_297,N_326);
or U600 (N_600,N_409,N_427);
nor U601 (N_601,N_522,N_429);
or U602 (N_602,N_509,N_523);
and U603 (N_603,N_494,N_566);
or U604 (N_604,N_421,N_452);
and U605 (N_605,N_428,N_492);
nor U606 (N_606,N_559,N_502);
nor U607 (N_607,N_505,N_479);
xor U608 (N_608,N_581,N_497);
or U609 (N_609,N_466,N_530);
and U610 (N_610,N_503,N_526);
and U611 (N_611,N_487,N_449);
nor U612 (N_612,N_440,N_518);
nor U613 (N_613,N_474,N_496);
and U614 (N_614,N_580,N_463);
nor U615 (N_615,N_471,N_408);
and U616 (N_616,N_462,N_461);
nor U617 (N_617,N_506,N_415);
or U618 (N_618,N_589,N_553);
or U619 (N_619,N_560,N_422);
or U620 (N_620,N_489,N_550);
or U621 (N_621,N_444,N_554);
nor U622 (N_622,N_537,N_406);
or U623 (N_623,N_593,N_570);
nand U624 (N_624,N_431,N_418);
nand U625 (N_625,N_484,N_480);
or U626 (N_626,N_446,N_491);
nor U627 (N_627,N_458,N_533);
nand U628 (N_628,N_598,N_469);
nand U629 (N_629,N_585,N_470);
or U630 (N_630,N_435,N_594);
and U631 (N_631,N_569,N_448);
nand U632 (N_632,N_573,N_528);
or U633 (N_633,N_586,N_407);
nor U634 (N_634,N_430,N_511);
or U635 (N_635,N_411,N_582);
nand U636 (N_636,N_450,N_498);
nor U637 (N_637,N_551,N_515);
nor U638 (N_638,N_562,N_543);
nor U639 (N_639,N_536,N_599);
nand U640 (N_640,N_516,N_504);
nor U641 (N_641,N_565,N_577);
or U642 (N_642,N_552,N_454);
nand U643 (N_643,N_500,N_545);
nand U644 (N_644,N_568,N_524);
nor U645 (N_645,N_433,N_412);
nor U646 (N_646,N_592,N_434);
and U647 (N_647,N_410,N_467);
nand U648 (N_648,N_473,N_538);
and U649 (N_649,N_507,N_529);
nand U650 (N_650,N_597,N_535);
nand U651 (N_651,N_485,N_404);
nor U652 (N_652,N_499,N_447);
nor U653 (N_653,N_417,N_437);
nor U654 (N_654,N_574,N_425);
and U655 (N_655,N_490,N_477);
nor U656 (N_656,N_483,N_482);
or U657 (N_657,N_563,N_520);
nor U658 (N_658,N_420,N_596);
and U659 (N_659,N_546,N_488);
nand U660 (N_660,N_558,N_512);
or U661 (N_661,N_531,N_579);
and U662 (N_662,N_453,N_517);
nand U663 (N_663,N_578,N_424);
or U664 (N_664,N_438,N_541);
nand U665 (N_665,N_584,N_561);
or U666 (N_666,N_501,N_556);
nand U667 (N_667,N_519,N_591);
nand U668 (N_668,N_557,N_590);
nor U669 (N_669,N_583,N_525);
and U670 (N_670,N_400,N_587);
or U671 (N_671,N_575,N_472);
or U672 (N_672,N_401,N_571);
or U673 (N_673,N_459,N_442);
or U674 (N_674,N_495,N_493);
and U675 (N_675,N_481,N_443);
xnor U676 (N_676,N_595,N_478);
or U677 (N_677,N_456,N_521);
nand U678 (N_678,N_436,N_576);
nand U679 (N_679,N_468,N_416);
nand U680 (N_680,N_510,N_527);
and U681 (N_681,N_445,N_441);
and U682 (N_682,N_464,N_532);
or U683 (N_683,N_432,N_402);
or U684 (N_684,N_476,N_564);
and U685 (N_685,N_540,N_414);
and U686 (N_686,N_457,N_567);
nand U687 (N_687,N_413,N_513);
nand U688 (N_688,N_514,N_572);
nand U689 (N_689,N_548,N_403);
and U690 (N_690,N_455,N_547);
nand U691 (N_691,N_460,N_439);
or U692 (N_692,N_549,N_426);
or U693 (N_693,N_451,N_419);
or U694 (N_694,N_542,N_465);
and U695 (N_695,N_539,N_508);
nor U696 (N_696,N_555,N_405);
xor U697 (N_697,N_534,N_486);
nand U698 (N_698,N_588,N_544);
nand U699 (N_699,N_475,N_423);
nand U700 (N_700,N_401,N_485);
and U701 (N_701,N_435,N_479);
nand U702 (N_702,N_527,N_408);
nand U703 (N_703,N_410,N_499);
and U704 (N_704,N_425,N_567);
nand U705 (N_705,N_544,N_454);
or U706 (N_706,N_534,N_433);
and U707 (N_707,N_570,N_429);
or U708 (N_708,N_461,N_592);
or U709 (N_709,N_483,N_400);
nand U710 (N_710,N_529,N_525);
or U711 (N_711,N_402,N_434);
and U712 (N_712,N_406,N_438);
and U713 (N_713,N_542,N_497);
nand U714 (N_714,N_473,N_460);
or U715 (N_715,N_416,N_497);
and U716 (N_716,N_411,N_569);
nor U717 (N_717,N_477,N_579);
and U718 (N_718,N_494,N_451);
nor U719 (N_719,N_528,N_436);
and U720 (N_720,N_587,N_425);
and U721 (N_721,N_430,N_453);
nand U722 (N_722,N_465,N_586);
or U723 (N_723,N_521,N_441);
and U724 (N_724,N_598,N_481);
and U725 (N_725,N_403,N_577);
nand U726 (N_726,N_435,N_409);
or U727 (N_727,N_593,N_401);
and U728 (N_728,N_569,N_506);
nand U729 (N_729,N_454,N_534);
or U730 (N_730,N_436,N_488);
nand U731 (N_731,N_426,N_488);
or U732 (N_732,N_506,N_439);
nor U733 (N_733,N_407,N_587);
and U734 (N_734,N_550,N_441);
and U735 (N_735,N_597,N_491);
nand U736 (N_736,N_441,N_460);
or U737 (N_737,N_499,N_434);
and U738 (N_738,N_465,N_443);
nand U739 (N_739,N_445,N_537);
nor U740 (N_740,N_436,N_560);
or U741 (N_741,N_593,N_454);
or U742 (N_742,N_422,N_548);
nand U743 (N_743,N_433,N_426);
nand U744 (N_744,N_586,N_558);
nand U745 (N_745,N_494,N_483);
nand U746 (N_746,N_539,N_481);
and U747 (N_747,N_496,N_562);
and U748 (N_748,N_403,N_443);
or U749 (N_749,N_500,N_434);
or U750 (N_750,N_504,N_407);
nor U751 (N_751,N_496,N_484);
and U752 (N_752,N_510,N_479);
or U753 (N_753,N_548,N_580);
nor U754 (N_754,N_476,N_596);
nand U755 (N_755,N_582,N_492);
nor U756 (N_756,N_413,N_491);
and U757 (N_757,N_463,N_440);
nand U758 (N_758,N_527,N_598);
nor U759 (N_759,N_562,N_540);
nand U760 (N_760,N_400,N_431);
nand U761 (N_761,N_552,N_471);
nand U762 (N_762,N_430,N_554);
nand U763 (N_763,N_503,N_494);
nor U764 (N_764,N_537,N_561);
nand U765 (N_765,N_523,N_549);
and U766 (N_766,N_524,N_534);
and U767 (N_767,N_415,N_561);
or U768 (N_768,N_504,N_558);
xnor U769 (N_769,N_576,N_566);
nor U770 (N_770,N_533,N_535);
nand U771 (N_771,N_574,N_524);
nor U772 (N_772,N_501,N_454);
nand U773 (N_773,N_560,N_553);
and U774 (N_774,N_563,N_560);
or U775 (N_775,N_460,N_555);
and U776 (N_776,N_598,N_569);
nor U777 (N_777,N_427,N_415);
and U778 (N_778,N_578,N_594);
nor U779 (N_779,N_516,N_550);
and U780 (N_780,N_504,N_442);
nand U781 (N_781,N_544,N_482);
nand U782 (N_782,N_559,N_516);
nand U783 (N_783,N_482,N_573);
or U784 (N_784,N_472,N_507);
or U785 (N_785,N_466,N_534);
or U786 (N_786,N_539,N_505);
and U787 (N_787,N_532,N_591);
or U788 (N_788,N_449,N_457);
and U789 (N_789,N_465,N_557);
and U790 (N_790,N_585,N_534);
and U791 (N_791,N_583,N_514);
or U792 (N_792,N_540,N_542);
nand U793 (N_793,N_452,N_570);
or U794 (N_794,N_554,N_591);
nor U795 (N_795,N_520,N_433);
nand U796 (N_796,N_453,N_428);
and U797 (N_797,N_420,N_477);
and U798 (N_798,N_430,N_490);
and U799 (N_799,N_597,N_532);
nand U800 (N_800,N_661,N_664);
nor U801 (N_801,N_757,N_693);
and U802 (N_802,N_618,N_609);
nor U803 (N_803,N_794,N_717);
or U804 (N_804,N_670,N_614);
and U805 (N_805,N_660,N_784);
or U806 (N_806,N_788,N_774);
or U807 (N_807,N_783,N_778);
nand U808 (N_808,N_793,N_763);
and U809 (N_809,N_699,N_668);
or U810 (N_810,N_600,N_644);
or U811 (N_811,N_650,N_637);
and U812 (N_812,N_713,N_738);
nand U813 (N_813,N_606,N_686);
nand U814 (N_814,N_630,N_617);
and U815 (N_815,N_754,N_762);
nor U816 (N_816,N_781,N_628);
and U817 (N_817,N_641,N_616);
nand U818 (N_818,N_646,N_666);
nor U819 (N_819,N_697,N_712);
or U820 (N_820,N_752,N_761);
or U821 (N_821,N_746,N_651);
or U822 (N_822,N_667,N_772);
or U823 (N_823,N_731,N_698);
or U824 (N_824,N_603,N_716);
or U825 (N_825,N_689,N_755);
or U826 (N_826,N_624,N_747);
or U827 (N_827,N_789,N_608);
nor U828 (N_828,N_739,N_643);
or U829 (N_829,N_741,N_765);
nor U830 (N_830,N_780,N_640);
and U831 (N_831,N_773,N_727);
nand U832 (N_832,N_750,N_657);
nor U833 (N_833,N_740,N_610);
nor U834 (N_834,N_662,N_620);
and U835 (N_835,N_692,N_745);
or U836 (N_836,N_768,N_631);
nand U837 (N_837,N_604,N_714);
nor U838 (N_838,N_766,N_648);
nor U839 (N_839,N_691,N_797);
nor U840 (N_840,N_735,N_695);
nand U841 (N_841,N_736,N_612);
nand U842 (N_842,N_707,N_751);
or U843 (N_843,N_759,N_787);
nor U844 (N_844,N_632,N_626);
or U845 (N_845,N_635,N_785);
and U846 (N_846,N_694,N_709);
nor U847 (N_847,N_673,N_715);
or U848 (N_848,N_654,N_723);
nand U849 (N_849,N_769,N_796);
nor U850 (N_850,N_798,N_671);
or U851 (N_851,N_724,N_615);
nand U852 (N_852,N_685,N_607);
and U853 (N_853,N_672,N_619);
or U854 (N_854,N_658,N_737);
nand U855 (N_855,N_627,N_790);
nand U856 (N_856,N_629,N_786);
and U857 (N_857,N_704,N_748);
nand U858 (N_858,N_705,N_696);
and U859 (N_859,N_756,N_653);
nor U860 (N_860,N_726,N_744);
or U861 (N_861,N_791,N_684);
nor U862 (N_862,N_775,N_681);
and U863 (N_863,N_760,N_636);
or U864 (N_864,N_656,N_734);
nor U865 (N_865,N_719,N_682);
nand U866 (N_866,N_678,N_729);
and U867 (N_867,N_633,N_721);
or U868 (N_868,N_725,N_683);
and U869 (N_869,N_779,N_767);
and U870 (N_870,N_718,N_655);
and U871 (N_871,N_605,N_702);
or U872 (N_872,N_792,N_733);
nor U873 (N_873,N_674,N_758);
nor U874 (N_874,N_776,N_708);
and U875 (N_875,N_669,N_743);
nand U876 (N_876,N_638,N_677);
or U877 (N_877,N_675,N_690);
nand U878 (N_878,N_621,N_659);
and U879 (N_879,N_676,N_728);
and U880 (N_880,N_700,N_665);
nor U881 (N_881,N_799,N_680);
and U882 (N_882,N_611,N_634);
xor U883 (N_883,N_687,N_710);
nor U884 (N_884,N_679,N_642);
nand U885 (N_885,N_602,N_764);
nand U886 (N_886,N_711,N_777);
nand U887 (N_887,N_795,N_645);
or U888 (N_888,N_649,N_742);
nand U889 (N_889,N_770,N_732);
or U890 (N_890,N_703,N_688);
nand U891 (N_891,N_730,N_749);
nand U892 (N_892,N_753,N_706);
nor U893 (N_893,N_622,N_613);
nand U894 (N_894,N_771,N_601);
nor U895 (N_895,N_625,N_652);
or U896 (N_896,N_782,N_720);
nand U897 (N_897,N_647,N_663);
and U898 (N_898,N_623,N_701);
nor U899 (N_899,N_722,N_639);
and U900 (N_900,N_725,N_648);
and U901 (N_901,N_614,N_621);
nor U902 (N_902,N_771,N_650);
nor U903 (N_903,N_758,N_734);
and U904 (N_904,N_661,N_676);
nand U905 (N_905,N_626,N_720);
nand U906 (N_906,N_628,N_746);
nand U907 (N_907,N_798,N_619);
nand U908 (N_908,N_788,N_753);
or U909 (N_909,N_619,N_757);
nand U910 (N_910,N_744,N_653);
or U911 (N_911,N_796,N_784);
nor U912 (N_912,N_616,N_700);
nor U913 (N_913,N_671,N_772);
nor U914 (N_914,N_665,N_625);
or U915 (N_915,N_766,N_799);
nand U916 (N_916,N_761,N_621);
or U917 (N_917,N_743,N_739);
and U918 (N_918,N_632,N_770);
and U919 (N_919,N_687,N_791);
nand U920 (N_920,N_624,N_677);
and U921 (N_921,N_679,N_637);
nor U922 (N_922,N_617,N_756);
nand U923 (N_923,N_637,N_789);
and U924 (N_924,N_714,N_740);
or U925 (N_925,N_727,N_719);
or U926 (N_926,N_742,N_707);
nand U927 (N_927,N_799,N_755);
or U928 (N_928,N_790,N_708);
nor U929 (N_929,N_608,N_618);
nand U930 (N_930,N_756,N_713);
or U931 (N_931,N_633,N_669);
and U932 (N_932,N_754,N_707);
and U933 (N_933,N_796,N_623);
nand U934 (N_934,N_771,N_683);
nor U935 (N_935,N_656,N_719);
or U936 (N_936,N_754,N_603);
or U937 (N_937,N_783,N_620);
and U938 (N_938,N_702,N_773);
or U939 (N_939,N_705,N_740);
or U940 (N_940,N_715,N_710);
and U941 (N_941,N_631,N_746);
nor U942 (N_942,N_774,N_624);
or U943 (N_943,N_602,N_631);
and U944 (N_944,N_673,N_766);
or U945 (N_945,N_626,N_711);
nor U946 (N_946,N_721,N_679);
and U947 (N_947,N_706,N_703);
nor U948 (N_948,N_794,N_731);
nand U949 (N_949,N_700,N_624);
and U950 (N_950,N_631,N_732);
or U951 (N_951,N_713,N_739);
nand U952 (N_952,N_704,N_708);
or U953 (N_953,N_707,N_724);
and U954 (N_954,N_633,N_604);
or U955 (N_955,N_666,N_669);
and U956 (N_956,N_702,N_657);
nand U957 (N_957,N_780,N_775);
or U958 (N_958,N_637,N_666);
and U959 (N_959,N_752,N_686);
nand U960 (N_960,N_759,N_660);
nand U961 (N_961,N_647,N_781);
nor U962 (N_962,N_712,N_669);
and U963 (N_963,N_729,N_764);
nor U964 (N_964,N_644,N_718);
nor U965 (N_965,N_751,N_711);
nor U966 (N_966,N_618,N_728);
and U967 (N_967,N_765,N_670);
nor U968 (N_968,N_763,N_643);
or U969 (N_969,N_667,N_781);
nor U970 (N_970,N_601,N_688);
nor U971 (N_971,N_685,N_711);
nor U972 (N_972,N_767,N_643);
nor U973 (N_973,N_716,N_664);
and U974 (N_974,N_634,N_683);
or U975 (N_975,N_653,N_721);
and U976 (N_976,N_682,N_799);
or U977 (N_977,N_636,N_791);
nor U978 (N_978,N_690,N_699);
and U979 (N_979,N_600,N_785);
nand U980 (N_980,N_723,N_767);
nor U981 (N_981,N_770,N_638);
nand U982 (N_982,N_746,N_672);
nand U983 (N_983,N_615,N_792);
nor U984 (N_984,N_690,N_731);
or U985 (N_985,N_773,N_610);
nand U986 (N_986,N_748,N_665);
nor U987 (N_987,N_717,N_781);
or U988 (N_988,N_642,N_739);
and U989 (N_989,N_650,N_728);
or U990 (N_990,N_788,N_704);
nand U991 (N_991,N_635,N_781);
nand U992 (N_992,N_788,N_705);
nand U993 (N_993,N_738,N_655);
and U994 (N_994,N_729,N_657);
and U995 (N_995,N_762,N_665);
and U996 (N_996,N_730,N_610);
nor U997 (N_997,N_718,N_750);
or U998 (N_998,N_790,N_606);
and U999 (N_999,N_709,N_605);
or U1000 (N_1000,N_962,N_917);
nor U1001 (N_1001,N_963,N_945);
and U1002 (N_1002,N_955,N_912);
nand U1003 (N_1003,N_972,N_967);
nand U1004 (N_1004,N_928,N_965);
or U1005 (N_1005,N_873,N_867);
and U1006 (N_1006,N_875,N_926);
nor U1007 (N_1007,N_956,N_891);
nor U1008 (N_1008,N_971,N_944);
nor U1009 (N_1009,N_843,N_846);
nor U1010 (N_1010,N_813,N_801);
nand U1011 (N_1011,N_897,N_942);
or U1012 (N_1012,N_913,N_816);
or U1013 (N_1013,N_903,N_840);
nand U1014 (N_1014,N_809,N_957);
and U1015 (N_1015,N_894,N_900);
and U1016 (N_1016,N_861,N_905);
nor U1017 (N_1017,N_878,N_828);
and U1018 (N_1018,N_826,N_807);
nand U1019 (N_1019,N_915,N_970);
nand U1020 (N_1020,N_877,N_866);
nand U1021 (N_1021,N_839,N_977);
or U1022 (N_1022,N_858,N_968);
or U1023 (N_1023,N_863,N_918);
and U1024 (N_1024,N_980,N_929);
nor U1025 (N_1025,N_958,N_954);
and U1026 (N_1026,N_989,N_938);
and U1027 (N_1027,N_985,N_857);
nand U1028 (N_1028,N_802,N_998);
and U1029 (N_1029,N_806,N_833);
nor U1030 (N_1030,N_803,N_832);
nor U1031 (N_1031,N_871,N_908);
or U1032 (N_1032,N_898,N_860);
nand U1033 (N_1033,N_911,N_961);
nand U1034 (N_1034,N_808,N_909);
nor U1035 (N_1035,N_814,N_842);
or U1036 (N_1036,N_818,N_889);
and U1037 (N_1037,N_925,N_997);
or U1038 (N_1038,N_995,N_921);
nand U1039 (N_1039,N_827,N_932);
xnor U1040 (N_1040,N_950,N_848);
nor U1041 (N_1041,N_902,N_964);
or U1042 (N_1042,N_831,N_829);
nand U1043 (N_1043,N_988,N_974);
or U1044 (N_1044,N_939,N_890);
nor U1045 (N_1045,N_830,N_941);
nor U1046 (N_1046,N_907,N_914);
and U1047 (N_1047,N_872,N_959);
and U1048 (N_1048,N_948,N_934);
nand U1049 (N_1049,N_966,N_810);
nand U1050 (N_1050,N_947,N_933);
or U1051 (N_1051,N_996,N_820);
or U1052 (N_1052,N_978,N_868);
nand U1053 (N_1053,N_836,N_904);
nor U1054 (N_1054,N_991,N_924);
or U1055 (N_1055,N_823,N_864);
and U1056 (N_1056,N_990,N_804);
nor U1057 (N_1057,N_943,N_800);
and U1058 (N_1058,N_852,N_821);
nand U1059 (N_1059,N_888,N_855);
nand U1060 (N_1060,N_931,N_975);
and U1061 (N_1061,N_880,N_847);
or U1062 (N_1062,N_999,N_984);
nand U1063 (N_1063,N_865,N_979);
or U1064 (N_1064,N_919,N_834);
nor U1065 (N_1065,N_922,N_951);
or U1066 (N_1066,N_853,N_983);
nor U1067 (N_1067,N_850,N_937);
nand U1068 (N_1068,N_936,N_893);
and U1069 (N_1069,N_812,N_920);
or U1070 (N_1070,N_817,N_805);
and U1071 (N_1071,N_841,N_949);
and U1072 (N_1072,N_869,N_859);
or U1073 (N_1073,N_906,N_976);
nor U1074 (N_1074,N_874,N_887);
and U1075 (N_1075,N_883,N_838);
nand U1076 (N_1076,N_835,N_824);
nand U1077 (N_1077,N_899,N_946);
and U1078 (N_1078,N_882,N_892);
or U1079 (N_1079,N_927,N_982);
and U1080 (N_1080,N_876,N_960);
and U1081 (N_1081,N_851,N_885);
or U1082 (N_1082,N_953,N_862);
and U1083 (N_1083,N_849,N_811);
or U1084 (N_1084,N_884,N_923);
nor U1085 (N_1085,N_994,N_910);
nor U1086 (N_1086,N_981,N_895);
nor U1087 (N_1087,N_940,N_952);
and U1088 (N_1088,N_935,N_886);
or U1089 (N_1089,N_870,N_993);
nor U1090 (N_1090,N_896,N_844);
nor U1091 (N_1091,N_825,N_930);
nand U1092 (N_1092,N_822,N_856);
nand U1093 (N_1093,N_881,N_901);
nand U1094 (N_1094,N_837,N_854);
nor U1095 (N_1095,N_916,N_973);
nand U1096 (N_1096,N_986,N_969);
and U1097 (N_1097,N_845,N_819);
and U1098 (N_1098,N_987,N_992);
and U1099 (N_1099,N_815,N_879);
and U1100 (N_1100,N_967,N_977);
nor U1101 (N_1101,N_913,N_902);
nor U1102 (N_1102,N_918,N_801);
and U1103 (N_1103,N_973,N_960);
nand U1104 (N_1104,N_939,N_862);
nor U1105 (N_1105,N_883,N_961);
and U1106 (N_1106,N_804,N_824);
nor U1107 (N_1107,N_874,N_957);
or U1108 (N_1108,N_942,N_997);
nand U1109 (N_1109,N_831,N_917);
or U1110 (N_1110,N_867,N_853);
nor U1111 (N_1111,N_935,N_919);
or U1112 (N_1112,N_887,N_928);
nor U1113 (N_1113,N_893,N_950);
nand U1114 (N_1114,N_884,N_956);
nor U1115 (N_1115,N_907,N_839);
nand U1116 (N_1116,N_874,N_965);
nor U1117 (N_1117,N_894,N_941);
and U1118 (N_1118,N_934,N_920);
nand U1119 (N_1119,N_811,N_854);
and U1120 (N_1120,N_815,N_914);
nor U1121 (N_1121,N_885,N_992);
nand U1122 (N_1122,N_876,N_821);
or U1123 (N_1123,N_847,N_815);
nand U1124 (N_1124,N_915,N_857);
nor U1125 (N_1125,N_854,N_931);
nand U1126 (N_1126,N_992,N_932);
xor U1127 (N_1127,N_915,N_945);
xor U1128 (N_1128,N_819,N_973);
nor U1129 (N_1129,N_889,N_978);
and U1130 (N_1130,N_876,N_957);
nand U1131 (N_1131,N_861,N_808);
or U1132 (N_1132,N_874,N_800);
nor U1133 (N_1133,N_860,N_852);
and U1134 (N_1134,N_856,N_918);
and U1135 (N_1135,N_877,N_955);
or U1136 (N_1136,N_830,N_887);
nor U1137 (N_1137,N_809,N_865);
nor U1138 (N_1138,N_833,N_979);
nand U1139 (N_1139,N_883,N_889);
and U1140 (N_1140,N_821,N_929);
nor U1141 (N_1141,N_828,N_986);
nor U1142 (N_1142,N_850,N_835);
and U1143 (N_1143,N_962,N_933);
nor U1144 (N_1144,N_809,N_903);
nor U1145 (N_1145,N_808,N_809);
and U1146 (N_1146,N_845,N_948);
nor U1147 (N_1147,N_841,N_868);
xnor U1148 (N_1148,N_838,N_968);
and U1149 (N_1149,N_937,N_895);
nand U1150 (N_1150,N_855,N_958);
and U1151 (N_1151,N_921,N_819);
nor U1152 (N_1152,N_949,N_951);
or U1153 (N_1153,N_831,N_929);
or U1154 (N_1154,N_863,N_926);
nor U1155 (N_1155,N_839,N_813);
or U1156 (N_1156,N_966,N_851);
and U1157 (N_1157,N_826,N_912);
nand U1158 (N_1158,N_896,N_857);
nand U1159 (N_1159,N_832,N_913);
or U1160 (N_1160,N_840,N_839);
nand U1161 (N_1161,N_812,N_863);
nand U1162 (N_1162,N_926,N_997);
nand U1163 (N_1163,N_914,N_803);
nor U1164 (N_1164,N_835,N_807);
nand U1165 (N_1165,N_980,N_985);
or U1166 (N_1166,N_861,N_837);
or U1167 (N_1167,N_931,N_892);
and U1168 (N_1168,N_854,N_847);
and U1169 (N_1169,N_847,N_985);
nor U1170 (N_1170,N_987,N_989);
nand U1171 (N_1171,N_827,N_855);
nor U1172 (N_1172,N_963,N_959);
nor U1173 (N_1173,N_882,N_831);
nor U1174 (N_1174,N_982,N_906);
nand U1175 (N_1175,N_867,N_805);
nand U1176 (N_1176,N_880,N_866);
and U1177 (N_1177,N_877,N_938);
or U1178 (N_1178,N_855,N_963);
nand U1179 (N_1179,N_807,N_898);
nor U1180 (N_1180,N_816,N_875);
and U1181 (N_1181,N_993,N_846);
nor U1182 (N_1182,N_970,N_891);
nor U1183 (N_1183,N_883,N_854);
nor U1184 (N_1184,N_960,N_820);
and U1185 (N_1185,N_800,N_941);
or U1186 (N_1186,N_820,N_855);
and U1187 (N_1187,N_920,N_868);
nand U1188 (N_1188,N_850,N_976);
and U1189 (N_1189,N_804,N_979);
nand U1190 (N_1190,N_942,N_954);
nand U1191 (N_1191,N_872,N_885);
nand U1192 (N_1192,N_868,N_905);
xnor U1193 (N_1193,N_833,N_882);
and U1194 (N_1194,N_910,N_907);
or U1195 (N_1195,N_853,N_927);
or U1196 (N_1196,N_966,N_841);
or U1197 (N_1197,N_918,N_882);
and U1198 (N_1198,N_805,N_904);
nor U1199 (N_1199,N_920,N_840);
and U1200 (N_1200,N_1076,N_1187);
and U1201 (N_1201,N_1105,N_1017);
nor U1202 (N_1202,N_1097,N_1140);
nor U1203 (N_1203,N_1142,N_1136);
nor U1204 (N_1204,N_1111,N_1058);
or U1205 (N_1205,N_1163,N_1080);
nor U1206 (N_1206,N_1119,N_1088);
and U1207 (N_1207,N_1192,N_1137);
nand U1208 (N_1208,N_1158,N_1131);
nand U1209 (N_1209,N_1001,N_1059);
or U1210 (N_1210,N_1121,N_1185);
nand U1211 (N_1211,N_1126,N_1063);
or U1212 (N_1212,N_1153,N_1159);
and U1213 (N_1213,N_1188,N_1171);
nor U1214 (N_1214,N_1128,N_1084);
and U1215 (N_1215,N_1167,N_1009);
nor U1216 (N_1216,N_1184,N_1071);
and U1217 (N_1217,N_1056,N_1031);
or U1218 (N_1218,N_1079,N_1177);
and U1219 (N_1219,N_1054,N_1133);
and U1220 (N_1220,N_1070,N_1147);
and U1221 (N_1221,N_1081,N_1166);
nor U1222 (N_1222,N_1003,N_1035);
and U1223 (N_1223,N_1144,N_1149);
nand U1224 (N_1224,N_1049,N_1044);
nand U1225 (N_1225,N_1089,N_1006);
and U1226 (N_1226,N_1183,N_1138);
nand U1227 (N_1227,N_1018,N_1077);
or U1228 (N_1228,N_1132,N_1152);
nand U1229 (N_1229,N_1155,N_1180);
nor U1230 (N_1230,N_1175,N_1050);
nor U1231 (N_1231,N_1117,N_1012);
nor U1232 (N_1232,N_1195,N_1108);
nor U1233 (N_1233,N_1020,N_1019);
and U1234 (N_1234,N_1011,N_1026);
nor U1235 (N_1235,N_1043,N_1186);
and U1236 (N_1236,N_1010,N_1182);
nand U1237 (N_1237,N_1114,N_1040);
or U1238 (N_1238,N_1139,N_1107);
nand U1239 (N_1239,N_1116,N_1156);
or U1240 (N_1240,N_1115,N_1096);
nand U1241 (N_1241,N_1061,N_1085);
or U1242 (N_1242,N_1090,N_1066);
nand U1243 (N_1243,N_1002,N_1099);
xnor U1244 (N_1244,N_1170,N_1073);
nor U1245 (N_1245,N_1038,N_1157);
nand U1246 (N_1246,N_1022,N_1091);
nor U1247 (N_1247,N_1065,N_1094);
or U1248 (N_1248,N_1098,N_1199);
and U1249 (N_1249,N_1027,N_1032);
or U1250 (N_1250,N_1030,N_1179);
nor U1251 (N_1251,N_1150,N_1103);
nor U1252 (N_1252,N_1172,N_1036);
and U1253 (N_1253,N_1135,N_1000);
nor U1254 (N_1254,N_1104,N_1174);
and U1255 (N_1255,N_1191,N_1023);
nor U1256 (N_1256,N_1067,N_1053);
nor U1257 (N_1257,N_1057,N_1196);
nor U1258 (N_1258,N_1148,N_1013);
nand U1259 (N_1259,N_1145,N_1029);
or U1260 (N_1260,N_1072,N_1102);
nor U1261 (N_1261,N_1130,N_1100);
nand U1262 (N_1262,N_1068,N_1169);
or U1263 (N_1263,N_1037,N_1127);
and U1264 (N_1264,N_1123,N_1120);
and U1265 (N_1265,N_1021,N_1124);
nand U1266 (N_1266,N_1194,N_1143);
nand U1267 (N_1267,N_1082,N_1028);
or U1268 (N_1268,N_1198,N_1015);
and U1269 (N_1269,N_1151,N_1062);
or U1270 (N_1270,N_1052,N_1112);
and U1271 (N_1271,N_1095,N_1078);
or U1272 (N_1272,N_1101,N_1046);
xor U1273 (N_1273,N_1181,N_1118);
or U1274 (N_1274,N_1083,N_1055);
and U1275 (N_1275,N_1197,N_1154);
or U1276 (N_1276,N_1164,N_1162);
nor U1277 (N_1277,N_1141,N_1193);
or U1278 (N_1278,N_1113,N_1168);
and U1279 (N_1279,N_1041,N_1069);
or U1280 (N_1280,N_1165,N_1129);
nand U1281 (N_1281,N_1160,N_1014);
and U1282 (N_1282,N_1173,N_1025);
and U1283 (N_1283,N_1039,N_1190);
or U1284 (N_1284,N_1008,N_1051);
xnor U1285 (N_1285,N_1106,N_1134);
or U1286 (N_1286,N_1034,N_1060);
or U1287 (N_1287,N_1176,N_1007);
nor U1288 (N_1288,N_1048,N_1086);
or U1289 (N_1289,N_1004,N_1178);
nor U1290 (N_1290,N_1161,N_1109);
nand U1291 (N_1291,N_1042,N_1024);
nor U1292 (N_1292,N_1087,N_1033);
nand U1293 (N_1293,N_1125,N_1064);
nor U1294 (N_1294,N_1047,N_1092);
and U1295 (N_1295,N_1016,N_1122);
nand U1296 (N_1296,N_1110,N_1189);
or U1297 (N_1297,N_1005,N_1074);
and U1298 (N_1298,N_1045,N_1093);
or U1299 (N_1299,N_1075,N_1146);
nor U1300 (N_1300,N_1009,N_1045);
or U1301 (N_1301,N_1071,N_1113);
or U1302 (N_1302,N_1013,N_1195);
and U1303 (N_1303,N_1061,N_1097);
nand U1304 (N_1304,N_1044,N_1120);
and U1305 (N_1305,N_1168,N_1075);
nand U1306 (N_1306,N_1175,N_1131);
or U1307 (N_1307,N_1040,N_1112);
nand U1308 (N_1308,N_1044,N_1011);
nand U1309 (N_1309,N_1056,N_1087);
nand U1310 (N_1310,N_1029,N_1135);
or U1311 (N_1311,N_1156,N_1070);
nor U1312 (N_1312,N_1031,N_1197);
or U1313 (N_1313,N_1016,N_1163);
or U1314 (N_1314,N_1045,N_1028);
and U1315 (N_1315,N_1026,N_1003);
nor U1316 (N_1316,N_1034,N_1165);
nor U1317 (N_1317,N_1153,N_1155);
and U1318 (N_1318,N_1056,N_1014);
and U1319 (N_1319,N_1046,N_1109);
nor U1320 (N_1320,N_1068,N_1002);
or U1321 (N_1321,N_1028,N_1084);
nand U1322 (N_1322,N_1068,N_1070);
or U1323 (N_1323,N_1003,N_1089);
nor U1324 (N_1324,N_1093,N_1161);
or U1325 (N_1325,N_1152,N_1142);
nand U1326 (N_1326,N_1055,N_1167);
or U1327 (N_1327,N_1145,N_1071);
and U1328 (N_1328,N_1112,N_1035);
xnor U1329 (N_1329,N_1196,N_1116);
and U1330 (N_1330,N_1198,N_1138);
or U1331 (N_1331,N_1032,N_1108);
and U1332 (N_1332,N_1164,N_1141);
and U1333 (N_1333,N_1008,N_1189);
nor U1334 (N_1334,N_1167,N_1188);
and U1335 (N_1335,N_1198,N_1030);
nand U1336 (N_1336,N_1089,N_1071);
nand U1337 (N_1337,N_1057,N_1033);
or U1338 (N_1338,N_1180,N_1168);
or U1339 (N_1339,N_1045,N_1186);
and U1340 (N_1340,N_1011,N_1008);
or U1341 (N_1341,N_1121,N_1112);
nand U1342 (N_1342,N_1095,N_1104);
nand U1343 (N_1343,N_1139,N_1100);
nor U1344 (N_1344,N_1067,N_1041);
nor U1345 (N_1345,N_1190,N_1005);
or U1346 (N_1346,N_1144,N_1044);
and U1347 (N_1347,N_1011,N_1020);
nand U1348 (N_1348,N_1012,N_1171);
or U1349 (N_1349,N_1015,N_1182);
nand U1350 (N_1350,N_1008,N_1134);
or U1351 (N_1351,N_1172,N_1003);
nand U1352 (N_1352,N_1124,N_1085);
nor U1353 (N_1353,N_1046,N_1130);
nor U1354 (N_1354,N_1082,N_1125);
or U1355 (N_1355,N_1157,N_1190);
or U1356 (N_1356,N_1045,N_1025);
or U1357 (N_1357,N_1173,N_1122);
and U1358 (N_1358,N_1021,N_1133);
or U1359 (N_1359,N_1038,N_1190);
and U1360 (N_1360,N_1072,N_1039);
nor U1361 (N_1361,N_1048,N_1010);
nand U1362 (N_1362,N_1185,N_1050);
and U1363 (N_1363,N_1157,N_1199);
and U1364 (N_1364,N_1195,N_1015);
and U1365 (N_1365,N_1040,N_1123);
nor U1366 (N_1366,N_1177,N_1010);
and U1367 (N_1367,N_1128,N_1011);
nand U1368 (N_1368,N_1062,N_1047);
nor U1369 (N_1369,N_1094,N_1035);
and U1370 (N_1370,N_1125,N_1161);
or U1371 (N_1371,N_1169,N_1018);
and U1372 (N_1372,N_1096,N_1151);
nor U1373 (N_1373,N_1034,N_1000);
or U1374 (N_1374,N_1130,N_1180);
and U1375 (N_1375,N_1068,N_1039);
nand U1376 (N_1376,N_1098,N_1194);
nand U1377 (N_1377,N_1089,N_1186);
or U1378 (N_1378,N_1185,N_1088);
or U1379 (N_1379,N_1123,N_1004);
or U1380 (N_1380,N_1161,N_1102);
or U1381 (N_1381,N_1033,N_1020);
or U1382 (N_1382,N_1024,N_1030);
nand U1383 (N_1383,N_1072,N_1085);
or U1384 (N_1384,N_1146,N_1099);
or U1385 (N_1385,N_1118,N_1046);
nand U1386 (N_1386,N_1094,N_1067);
and U1387 (N_1387,N_1045,N_1167);
nand U1388 (N_1388,N_1192,N_1142);
or U1389 (N_1389,N_1114,N_1147);
or U1390 (N_1390,N_1176,N_1066);
nand U1391 (N_1391,N_1151,N_1080);
or U1392 (N_1392,N_1183,N_1156);
and U1393 (N_1393,N_1145,N_1050);
nand U1394 (N_1394,N_1107,N_1162);
nand U1395 (N_1395,N_1169,N_1010);
nor U1396 (N_1396,N_1091,N_1002);
nor U1397 (N_1397,N_1001,N_1160);
nand U1398 (N_1398,N_1061,N_1034);
nor U1399 (N_1399,N_1174,N_1170);
and U1400 (N_1400,N_1225,N_1277);
or U1401 (N_1401,N_1228,N_1287);
or U1402 (N_1402,N_1314,N_1272);
and U1403 (N_1403,N_1239,N_1378);
nand U1404 (N_1404,N_1388,N_1357);
nand U1405 (N_1405,N_1309,N_1211);
and U1406 (N_1406,N_1340,N_1222);
or U1407 (N_1407,N_1216,N_1311);
nor U1408 (N_1408,N_1399,N_1238);
nand U1409 (N_1409,N_1379,N_1358);
or U1410 (N_1410,N_1209,N_1253);
nor U1411 (N_1411,N_1224,N_1231);
nand U1412 (N_1412,N_1296,N_1252);
and U1413 (N_1413,N_1365,N_1278);
nor U1414 (N_1414,N_1327,N_1202);
nor U1415 (N_1415,N_1200,N_1334);
nor U1416 (N_1416,N_1319,N_1391);
nor U1417 (N_1417,N_1249,N_1214);
or U1418 (N_1418,N_1254,N_1341);
nand U1419 (N_1419,N_1303,N_1212);
and U1420 (N_1420,N_1396,N_1285);
nor U1421 (N_1421,N_1307,N_1317);
nor U1422 (N_1422,N_1356,N_1330);
nor U1423 (N_1423,N_1337,N_1367);
or U1424 (N_1424,N_1364,N_1268);
and U1425 (N_1425,N_1218,N_1322);
nand U1426 (N_1426,N_1204,N_1235);
nor U1427 (N_1427,N_1299,N_1382);
and U1428 (N_1428,N_1279,N_1312);
nand U1429 (N_1429,N_1241,N_1350);
nand U1430 (N_1430,N_1210,N_1282);
and U1431 (N_1431,N_1362,N_1257);
nor U1432 (N_1432,N_1261,N_1374);
or U1433 (N_1433,N_1288,N_1292);
or U1434 (N_1434,N_1243,N_1280);
nand U1435 (N_1435,N_1386,N_1208);
nand U1436 (N_1436,N_1283,N_1250);
nand U1437 (N_1437,N_1351,N_1304);
and U1438 (N_1438,N_1255,N_1315);
or U1439 (N_1439,N_1217,N_1259);
nor U1440 (N_1440,N_1264,N_1300);
nor U1441 (N_1441,N_1295,N_1232);
or U1442 (N_1442,N_1286,N_1332);
and U1443 (N_1443,N_1290,N_1236);
nand U1444 (N_1444,N_1389,N_1395);
nor U1445 (N_1445,N_1234,N_1392);
and U1446 (N_1446,N_1333,N_1220);
or U1447 (N_1447,N_1377,N_1335);
nand U1448 (N_1448,N_1294,N_1370);
or U1449 (N_1449,N_1326,N_1383);
nor U1450 (N_1450,N_1273,N_1320);
nand U1451 (N_1451,N_1301,N_1375);
and U1452 (N_1452,N_1274,N_1229);
nor U1453 (N_1453,N_1244,N_1376);
or U1454 (N_1454,N_1305,N_1213);
and U1455 (N_1455,N_1371,N_1384);
nand U1456 (N_1456,N_1360,N_1352);
or U1457 (N_1457,N_1328,N_1348);
or U1458 (N_1458,N_1251,N_1366);
nor U1459 (N_1459,N_1324,N_1267);
nor U1460 (N_1460,N_1205,N_1262);
nand U1461 (N_1461,N_1323,N_1276);
nand U1462 (N_1462,N_1237,N_1381);
or U1463 (N_1463,N_1219,N_1354);
and U1464 (N_1464,N_1223,N_1394);
nor U1465 (N_1465,N_1281,N_1215);
or U1466 (N_1466,N_1336,N_1347);
nand U1467 (N_1467,N_1293,N_1325);
nor U1468 (N_1468,N_1385,N_1372);
nor U1469 (N_1469,N_1310,N_1240);
nor U1470 (N_1470,N_1361,N_1342);
xor U1471 (N_1471,N_1245,N_1398);
and U1472 (N_1472,N_1284,N_1207);
and U1473 (N_1473,N_1206,N_1275);
or U1474 (N_1474,N_1242,N_1380);
and U1475 (N_1475,N_1227,N_1353);
nor U1476 (N_1476,N_1387,N_1390);
nor U1477 (N_1477,N_1368,N_1308);
or U1478 (N_1478,N_1393,N_1346);
or U1479 (N_1479,N_1265,N_1271);
nand U1480 (N_1480,N_1331,N_1291);
nor U1481 (N_1481,N_1343,N_1203);
nor U1482 (N_1482,N_1266,N_1329);
and U1483 (N_1483,N_1339,N_1201);
nor U1484 (N_1484,N_1270,N_1345);
nor U1485 (N_1485,N_1221,N_1297);
or U1486 (N_1486,N_1338,N_1302);
or U1487 (N_1487,N_1230,N_1247);
nand U1488 (N_1488,N_1359,N_1246);
nor U1489 (N_1489,N_1260,N_1373);
nand U1490 (N_1490,N_1233,N_1321);
and U1491 (N_1491,N_1306,N_1248);
or U1492 (N_1492,N_1369,N_1269);
nand U1493 (N_1493,N_1258,N_1298);
nand U1494 (N_1494,N_1363,N_1256);
or U1495 (N_1495,N_1226,N_1289);
and U1496 (N_1496,N_1313,N_1318);
nor U1497 (N_1497,N_1349,N_1344);
or U1498 (N_1498,N_1316,N_1355);
nor U1499 (N_1499,N_1263,N_1397);
or U1500 (N_1500,N_1268,N_1312);
nor U1501 (N_1501,N_1271,N_1217);
nand U1502 (N_1502,N_1311,N_1218);
nor U1503 (N_1503,N_1214,N_1341);
nand U1504 (N_1504,N_1293,N_1250);
and U1505 (N_1505,N_1302,N_1350);
and U1506 (N_1506,N_1297,N_1243);
or U1507 (N_1507,N_1308,N_1256);
nor U1508 (N_1508,N_1370,N_1270);
nand U1509 (N_1509,N_1358,N_1388);
and U1510 (N_1510,N_1360,N_1258);
xnor U1511 (N_1511,N_1274,N_1364);
and U1512 (N_1512,N_1243,N_1299);
nand U1513 (N_1513,N_1207,N_1229);
or U1514 (N_1514,N_1254,N_1249);
nor U1515 (N_1515,N_1214,N_1369);
and U1516 (N_1516,N_1310,N_1307);
nand U1517 (N_1517,N_1357,N_1342);
nor U1518 (N_1518,N_1269,N_1321);
or U1519 (N_1519,N_1206,N_1245);
or U1520 (N_1520,N_1237,N_1348);
or U1521 (N_1521,N_1210,N_1355);
or U1522 (N_1522,N_1230,N_1380);
nand U1523 (N_1523,N_1255,N_1230);
and U1524 (N_1524,N_1366,N_1286);
and U1525 (N_1525,N_1314,N_1345);
or U1526 (N_1526,N_1352,N_1282);
or U1527 (N_1527,N_1267,N_1391);
and U1528 (N_1528,N_1337,N_1300);
or U1529 (N_1529,N_1204,N_1317);
nor U1530 (N_1530,N_1223,N_1252);
xnor U1531 (N_1531,N_1388,N_1344);
nor U1532 (N_1532,N_1269,N_1243);
and U1533 (N_1533,N_1224,N_1341);
and U1534 (N_1534,N_1346,N_1261);
and U1535 (N_1535,N_1384,N_1325);
or U1536 (N_1536,N_1288,N_1226);
nor U1537 (N_1537,N_1372,N_1365);
or U1538 (N_1538,N_1325,N_1392);
or U1539 (N_1539,N_1322,N_1328);
and U1540 (N_1540,N_1391,N_1225);
and U1541 (N_1541,N_1258,N_1237);
and U1542 (N_1542,N_1309,N_1348);
nor U1543 (N_1543,N_1333,N_1287);
and U1544 (N_1544,N_1236,N_1256);
and U1545 (N_1545,N_1220,N_1301);
or U1546 (N_1546,N_1217,N_1326);
or U1547 (N_1547,N_1392,N_1371);
nor U1548 (N_1548,N_1318,N_1206);
nor U1549 (N_1549,N_1295,N_1250);
and U1550 (N_1550,N_1371,N_1227);
and U1551 (N_1551,N_1348,N_1315);
nand U1552 (N_1552,N_1258,N_1367);
nor U1553 (N_1553,N_1286,N_1319);
or U1554 (N_1554,N_1352,N_1357);
or U1555 (N_1555,N_1288,N_1321);
nand U1556 (N_1556,N_1331,N_1369);
nand U1557 (N_1557,N_1368,N_1393);
and U1558 (N_1558,N_1356,N_1319);
or U1559 (N_1559,N_1241,N_1285);
nand U1560 (N_1560,N_1245,N_1375);
or U1561 (N_1561,N_1229,N_1331);
nor U1562 (N_1562,N_1365,N_1202);
or U1563 (N_1563,N_1265,N_1241);
nand U1564 (N_1564,N_1296,N_1204);
nor U1565 (N_1565,N_1381,N_1315);
nand U1566 (N_1566,N_1314,N_1319);
nor U1567 (N_1567,N_1383,N_1335);
nand U1568 (N_1568,N_1303,N_1257);
nor U1569 (N_1569,N_1367,N_1245);
xnor U1570 (N_1570,N_1379,N_1359);
nor U1571 (N_1571,N_1344,N_1374);
nor U1572 (N_1572,N_1244,N_1235);
and U1573 (N_1573,N_1282,N_1372);
nor U1574 (N_1574,N_1334,N_1369);
and U1575 (N_1575,N_1203,N_1296);
nor U1576 (N_1576,N_1332,N_1343);
or U1577 (N_1577,N_1249,N_1284);
or U1578 (N_1578,N_1378,N_1251);
and U1579 (N_1579,N_1349,N_1325);
nand U1580 (N_1580,N_1316,N_1269);
or U1581 (N_1581,N_1254,N_1348);
nand U1582 (N_1582,N_1271,N_1341);
nor U1583 (N_1583,N_1317,N_1333);
nor U1584 (N_1584,N_1256,N_1395);
nand U1585 (N_1585,N_1346,N_1322);
and U1586 (N_1586,N_1259,N_1345);
and U1587 (N_1587,N_1285,N_1296);
nor U1588 (N_1588,N_1240,N_1216);
nor U1589 (N_1589,N_1284,N_1357);
nand U1590 (N_1590,N_1324,N_1350);
and U1591 (N_1591,N_1390,N_1325);
or U1592 (N_1592,N_1354,N_1221);
or U1593 (N_1593,N_1285,N_1320);
and U1594 (N_1594,N_1212,N_1350);
or U1595 (N_1595,N_1383,N_1389);
nand U1596 (N_1596,N_1253,N_1381);
or U1597 (N_1597,N_1305,N_1363);
nand U1598 (N_1598,N_1208,N_1360);
and U1599 (N_1599,N_1397,N_1230);
nor U1600 (N_1600,N_1415,N_1505);
nor U1601 (N_1601,N_1520,N_1417);
or U1602 (N_1602,N_1452,N_1455);
and U1603 (N_1603,N_1515,N_1569);
and U1604 (N_1604,N_1457,N_1446);
and U1605 (N_1605,N_1498,N_1458);
nand U1606 (N_1606,N_1456,N_1459);
nor U1607 (N_1607,N_1516,N_1460);
nor U1608 (N_1608,N_1471,N_1441);
nor U1609 (N_1609,N_1438,N_1556);
nand U1610 (N_1610,N_1574,N_1432);
nand U1611 (N_1611,N_1428,N_1450);
nand U1612 (N_1612,N_1554,N_1511);
nor U1613 (N_1613,N_1496,N_1502);
nand U1614 (N_1614,N_1490,N_1521);
and U1615 (N_1615,N_1422,N_1572);
nand U1616 (N_1616,N_1591,N_1481);
nor U1617 (N_1617,N_1431,N_1531);
or U1618 (N_1618,N_1462,N_1499);
nand U1619 (N_1619,N_1436,N_1468);
nand U1620 (N_1620,N_1587,N_1540);
nor U1621 (N_1621,N_1437,N_1433);
nor U1622 (N_1622,N_1533,N_1461);
nor U1623 (N_1623,N_1578,N_1486);
or U1624 (N_1624,N_1501,N_1477);
nand U1625 (N_1625,N_1472,N_1504);
and U1626 (N_1626,N_1583,N_1558);
nand U1627 (N_1627,N_1416,N_1522);
nor U1628 (N_1628,N_1444,N_1405);
nor U1629 (N_1629,N_1534,N_1495);
and U1630 (N_1630,N_1497,N_1484);
and U1631 (N_1631,N_1403,N_1404);
nand U1632 (N_1632,N_1493,N_1549);
nor U1633 (N_1633,N_1410,N_1421);
and U1634 (N_1634,N_1463,N_1470);
nand U1635 (N_1635,N_1584,N_1527);
and U1636 (N_1636,N_1483,N_1434);
or U1637 (N_1637,N_1445,N_1568);
nand U1638 (N_1638,N_1593,N_1518);
and U1639 (N_1639,N_1443,N_1507);
nor U1640 (N_1640,N_1429,N_1508);
or U1641 (N_1641,N_1546,N_1423);
or U1642 (N_1642,N_1420,N_1412);
nand U1643 (N_1643,N_1494,N_1536);
or U1644 (N_1644,N_1576,N_1553);
and U1645 (N_1645,N_1401,N_1425);
nand U1646 (N_1646,N_1485,N_1476);
and U1647 (N_1647,N_1414,N_1409);
and U1648 (N_1648,N_1487,N_1535);
and U1649 (N_1649,N_1465,N_1560);
nand U1650 (N_1650,N_1528,N_1402);
and U1651 (N_1651,N_1514,N_1552);
nand U1652 (N_1652,N_1563,N_1430);
nand U1653 (N_1653,N_1539,N_1413);
or U1654 (N_1654,N_1474,N_1424);
and U1655 (N_1655,N_1550,N_1588);
nand U1656 (N_1656,N_1543,N_1571);
or U1657 (N_1657,N_1598,N_1542);
nand U1658 (N_1658,N_1454,N_1407);
nand U1659 (N_1659,N_1530,N_1473);
nand U1660 (N_1660,N_1548,N_1564);
xnor U1661 (N_1661,N_1567,N_1582);
nand U1662 (N_1662,N_1488,N_1491);
and U1663 (N_1663,N_1596,N_1559);
and U1664 (N_1664,N_1580,N_1592);
nor U1665 (N_1665,N_1506,N_1435);
and U1666 (N_1666,N_1541,N_1419);
nand U1667 (N_1667,N_1581,N_1492);
or U1668 (N_1668,N_1400,N_1529);
and U1669 (N_1669,N_1503,N_1565);
nor U1670 (N_1670,N_1500,N_1579);
and U1671 (N_1671,N_1509,N_1489);
or U1672 (N_1672,N_1577,N_1532);
or U1673 (N_1673,N_1524,N_1478);
or U1674 (N_1674,N_1545,N_1513);
nor U1675 (N_1675,N_1464,N_1585);
and U1676 (N_1676,N_1519,N_1547);
and U1677 (N_1677,N_1526,N_1480);
or U1678 (N_1678,N_1589,N_1590);
nand U1679 (N_1679,N_1570,N_1538);
and U1680 (N_1680,N_1575,N_1469);
or U1681 (N_1681,N_1411,N_1537);
nor U1682 (N_1682,N_1586,N_1427);
nor U1683 (N_1683,N_1442,N_1561);
nand U1684 (N_1684,N_1466,N_1510);
or U1685 (N_1685,N_1418,N_1551);
nand U1686 (N_1686,N_1451,N_1573);
nor U1687 (N_1687,N_1447,N_1557);
and U1688 (N_1688,N_1594,N_1439);
nand U1689 (N_1689,N_1440,N_1449);
or U1690 (N_1690,N_1595,N_1544);
or U1691 (N_1691,N_1448,N_1479);
and U1692 (N_1692,N_1426,N_1599);
nor U1693 (N_1693,N_1523,N_1467);
and U1694 (N_1694,N_1566,N_1512);
xor U1695 (N_1695,N_1555,N_1475);
nor U1696 (N_1696,N_1408,N_1517);
nor U1697 (N_1697,N_1453,N_1482);
and U1698 (N_1698,N_1597,N_1562);
nor U1699 (N_1699,N_1525,N_1406);
or U1700 (N_1700,N_1421,N_1506);
nor U1701 (N_1701,N_1542,N_1412);
nor U1702 (N_1702,N_1439,N_1591);
nor U1703 (N_1703,N_1568,N_1467);
and U1704 (N_1704,N_1561,N_1539);
and U1705 (N_1705,N_1521,N_1561);
or U1706 (N_1706,N_1497,N_1409);
nor U1707 (N_1707,N_1465,N_1580);
nor U1708 (N_1708,N_1425,N_1517);
nand U1709 (N_1709,N_1568,N_1539);
nand U1710 (N_1710,N_1429,N_1547);
xor U1711 (N_1711,N_1443,N_1551);
and U1712 (N_1712,N_1415,N_1459);
nand U1713 (N_1713,N_1447,N_1575);
nand U1714 (N_1714,N_1465,N_1526);
or U1715 (N_1715,N_1504,N_1425);
and U1716 (N_1716,N_1544,N_1575);
nor U1717 (N_1717,N_1517,N_1406);
or U1718 (N_1718,N_1523,N_1424);
nand U1719 (N_1719,N_1498,N_1556);
nor U1720 (N_1720,N_1541,N_1502);
or U1721 (N_1721,N_1450,N_1448);
or U1722 (N_1722,N_1462,N_1483);
and U1723 (N_1723,N_1579,N_1556);
nand U1724 (N_1724,N_1563,N_1502);
and U1725 (N_1725,N_1549,N_1517);
or U1726 (N_1726,N_1443,N_1541);
or U1727 (N_1727,N_1436,N_1480);
and U1728 (N_1728,N_1428,N_1419);
nand U1729 (N_1729,N_1453,N_1464);
and U1730 (N_1730,N_1404,N_1510);
nand U1731 (N_1731,N_1541,N_1488);
nand U1732 (N_1732,N_1503,N_1588);
and U1733 (N_1733,N_1480,N_1519);
nor U1734 (N_1734,N_1524,N_1499);
or U1735 (N_1735,N_1565,N_1472);
or U1736 (N_1736,N_1537,N_1443);
or U1737 (N_1737,N_1460,N_1526);
nand U1738 (N_1738,N_1506,N_1529);
or U1739 (N_1739,N_1457,N_1466);
nand U1740 (N_1740,N_1571,N_1402);
nor U1741 (N_1741,N_1491,N_1559);
xnor U1742 (N_1742,N_1543,N_1458);
nand U1743 (N_1743,N_1442,N_1535);
or U1744 (N_1744,N_1443,N_1527);
nand U1745 (N_1745,N_1440,N_1553);
nand U1746 (N_1746,N_1435,N_1549);
or U1747 (N_1747,N_1597,N_1548);
and U1748 (N_1748,N_1528,N_1478);
nand U1749 (N_1749,N_1486,N_1569);
nand U1750 (N_1750,N_1552,N_1542);
and U1751 (N_1751,N_1530,N_1577);
and U1752 (N_1752,N_1400,N_1452);
nor U1753 (N_1753,N_1518,N_1580);
or U1754 (N_1754,N_1558,N_1435);
and U1755 (N_1755,N_1429,N_1509);
and U1756 (N_1756,N_1490,N_1590);
nor U1757 (N_1757,N_1545,N_1546);
or U1758 (N_1758,N_1488,N_1421);
and U1759 (N_1759,N_1528,N_1494);
and U1760 (N_1760,N_1596,N_1544);
nand U1761 (N_1761,N_1495,N_1554);
nor U1762 (N_1762,N_1458,N_1594);
or U1763 (N_1763,N_1532,N_1477);
and U1764 (N_1764,N_1471,N_1431);
nand U1765 (N_1765,N_1517,N_1597);
nand U1766 (N_1766,N_1502,N_1434);
nor U1767 (N_1767,N_1495,N_1552);
nand U1768 (N_1768,N_1552,N_1499);
nor U1769 (N_1769,N_1500,N_1533);
and U1770 (N_1770,N_1502,N_1597);
nand U1771 (N_1771,N_1426,N_1530);
and U1772 (N_1772,N_1488,N_1456);
or U1773 (N_1773,N_1545,N_1564);
nor U1774 (N_1774,N_1408,N_1447);
nand U1775 (N_1775,N_1401,N_1426);
and U1776 (N_1776,N_1460,N_1518);
and U1777 (N_1777,N_1530,N_1454);
nand U1778 (N_1778,N_1452,N_1445);
nand U1779 (N_1779,N_1413,N_1455);
or U1780 (N_1780,N_1438,N_1550);
nor U1781 (N_1781,N_1500,N_1524);
or U1782 (N_1782,N_1413,N_1521);
and U1783 (N_1783,N_1402,N_1414);
nand U1784 (N_1784,N_1597,N_1433);
or U1785 (N_1785,N_1579,N_1456);
xnor U1786 (N_1786,N_1471,N_1516);
or U1787 (N_1787,N_1573,N_1428);
or U1788 (N_1788,N_1575,N_1507);
nor U1789 (N_1789,N_1571,N_1495);
and U1790 (N_1790,N_1438,N_1434);
and U1791 (N_1791,N_1400,N_1431);
and U1792 (N_1792,N_1586,N_1452);
and U1793 (N_1793,N_1453,N_1571);
nand U1794 (N_1794,N_1548,N_1518);
or U1795 (N_1795,N_1426,N_1468);
and U1796 (N_1796,N_1458,N_1493);
nand U1797 (N_1797,N_1589,N_1578);
and U1798 (N_1798,N_1494,N_1440);
nand U1799 (N_1799,N_1527,N_1469);
and U1800 (N_1800,N_1647,N_1656);
nand U1801 (N_1801,N_1602,N_1688);
nand U1802 (N_1802,N_1763,N_1653);
nand U1803 (N_1803,N_1787,N_1794);
nor U1804 (N_1804,N_1634,N_1784);
nor U1805 (N_1805,N_1621,N_1755);
and U1806 (N_1806,N_1677,N_1721);
nor U1807 (N_1807,N_1734,N_1754);
nor U1808 (N_1808,N_1773,N_1603);
nand U1809 (N_1809,N_1692,N_1719);
nand U1810 (N_1810,N_1772,N_1633);
nand U1811 (N_1811,N_1795,N_1680);
or U1812 (N_1812,N_1637,N_1673);
nor U1813 (N_1813,N_1701,N_1725);
nand U1814 (N_1814,N_1652,N_1645);
nor U1815 (N_1815,N_1726,N_1799);
or U1816 (N_1816,N_1746,N_1783);
or U1817 (N_1817,N_1761,N_1737);
nand U1818 (N_1818,N_1694,N_1709);
nor U1819 (N_1819,N_1663,N_1622);
nor U1820 (N_1820,N_1796,N_1661);
and U1821 (N_1821,N_1717,N_1628);
and U1822 (N_1822,N_1664,N_1760);
or U1823 (N_1823,N_1779,N_1678);
or U1824 (N_1824,N_1723,N_1789);
nand U1825 (N_1825,N_1611,N_1612);
nand U1826 (N_1826,N_1665,N_1630);
or U1827 (N_1827,N_1790,N_1752);
nor U1828 (N_1828,N_1636,N_1710);
nand U1829 (N_1829,N_1700,N_1606);
nor U1830 (N_1830,N_1659,N_1685);
nand U1831 (N_1831,N_1778,N_1676);
or U1832 (N_1832,N_1728,N_1736);
nand U1833 (N_1833,N_1629,N_1604);
and U1834 (N_1834,N_1600,N_1626);
and U1835 (N_1835,N_1727,N_1627);
nor U1836 (N_1836,N_1732,N_1751);
and U1837 (N_1837,N_1667,N_1650);
nor U1838 (N_1838,N_1646,N_1720);
or U1839 (N_1839,N_1711,N_1780);
nor U1840 (N_1840,N_1797,N_1693);
and U1841 (N_1841,N_1724,N_1733);
nand U1842 (N_1842,N_1689,N_1730);
nor U1843 (N_1843,N_1690,N_1605);
nand U1844 (N_1844,N_1706,N_1696);
nor U1845 (N_1845,N_1642,N_1608);
nor U1846 (N_1846,N_1639,N_1753);
nand U1847 (N_1847,N_1648,N_1671);
and U1848 (N_1848,N_1631,N_1615);
and U1849 (N_1849,N_1699,N_1742);
nand U1850 (N_1850,N_1782,N_1683);
nand U1851 (N_1851,N_1785,N_1749);
nand U1852 (N_1852,N_1731,N_1748);
or U1853 (N_1853,N_1613,N_1617);
and U1854 (N_1854,N_1704,N_1697);
and U1855 (N_1855,N_1607,N_1655);
nor U1856 (N_1856,N_1770,N_1675);
or U1857 (N_1857,N_1764,N_1788);
and U1858 (N_1858,N_1735,N_1691);
nand U1859 (N_1859,N_1669,N_1679);
xor U1860 (N_1860,N_1668,N_1684);
or U1861 (N_1861,N_1712,N_1624);
nand U1862 (N_1862,N_1640,N_1757);
nor U1863 (N_1863,N_1672,N_1705);
and U1864 (N_1864,N_1681,N_1777);
or U1865 (N_1865,N_1738,N_1687);
nand U1866 (N_1866,N_1619,N_1775);
nand U1867 (N_1867,N_1643,N_1695);
nor U1868 (N_1868,N_1616,N_1740);
nand U1869 (N_1869,N_1658,N_1657);
nor U1870 (N_1870,N_1708,N_1632);
nand U1871 (N_1871,N_1707,N_1762);
and U1872 (N_1872,N_1771,N_1798);
nor U1873 (N_1873,N_1774,N_1618);
or U1874 (N_1874,N_1722,N_1641);
nand U1875 (N_1875,N_1729,N_1714);
nor U1876 (N_1876,N_1776,N_1793);
or U1877 (N_1877,N_1644,N_1750);
or U1878 (N_1878,N_1635,N_1662);
and U1879 (N_1879,N_1765,N_1759);
or U1880 (N_1880,N_1768,N_1781);
and U1881 (N_1881,N_1791,N_1767);
and U1882 (N_1882,N_1744,N_1718);
nand U1883 (N_1883,N_1786,N_1620);
and U1884 (N_1884,N_1745,N_1610);
nand U1885 (N_1885,N_1739,N_1625);
and U1886 (N_1886,N_1743,N_1654);
and U1887 (N_1887,N_1747,N_1682);
nor U1888 (N_1888,N_1766,N_1769);
nand U1889 (N_1889,N_1660,N_1703);
and U1890 (N_1890,N_1670,N_1609);
and U1891 (N_1891,N_1741,N_1614);
nand U1892 (N_1892,N_1715,N_1674);
nand U1893 (N_1893,N_1758,N_1649);
nand U1894 (N_1894,N_1651,N_1716);
or U1895 (N_1895,N_1623,N_1792);
or U1896 (N_1896,N_1756,N_1702);
nor U1897 (N_1897,N_1638,N_1666);
nor U1898 (N_1898,N_1698,N_1713);
nand U1899 (N_1899,N_1601,N_1686);
and U1900 (N_1900,N_1711,N_1634);
nand U1901 (N_1901,N_1734,N_1704);
or U1902 (N_1902,N_1726,N_1781);
and U1903 (N_1903,N_1629,N_1775);
and U1904 (N_1904,N_1700,N_1708);
or U1905 (N_1905,N_1779,N_1768);
nor U1906 (N_1906,N_1799,N_1772);
or U1907 (N_1907,N_1700,N_1657);
or U1908 (N_1908,N_1656,N_1616);
nand U1909 (N_1909,N_1765,N_1764);
or U1910 (N_1910,N_1766,N_1649);
nor U1911 (N_1911,N_1643,N_1724);
or U1912 (N_1912,N_1605,N_1753);
or U1913 (N_1913,N_1665,N_1707);
and U1914 (N_1914,N_1678,N_1783);
nor U1915 (N_1915,N_1635,N_1795);
and U1916 (N_1916,N_1761,N_1619);
or U1917 (N_1917,N_1617,N_1766);
or U1918 (N_1918,N_1666,N_1755);
or U1919 (N_1919,N_1666,N_1736);
and U1920 (N_1920,N_1717,N_1621);
and U1921 (N_1921,N_1643,N_1641);
nand U1922 (N_1922,N_1682,N_1788);
and U1923 (N_1923,N_1767,N_1607);
nand U1924 (N_1924,N_1778,N_1631);
nor U1925 (N_1925,N_1793,N_1762);
and U1926 (N_1926,N_1706,N_1766);
and U1927 (N_1927,N_1788,N_1635);
nand U1928 (N_1928,N_1618,N_1642);
and U1929 (N_1929,N_1710,N_1730);
nor U1930 (N_1930,N_1761,N_1739);
nand U1931 (N_1931,N_1745,N_1744);
and U1932 (N_1932,N_1755,N_1732);
nand U1933 (N_1933,N_1619,N_1733);
nor U1934 (N_1934,N_1714,N_1791);
or U1935 (N_1935,N_1768,N_1786);
nor U1936 (N_1936,N_1678,N_1785);
and U1937 (N_1937,N_1690,N_1706);
and U1938 (N_1938,N_1653,N_1635);
and U1939 (N_1939,N_1662,N_1728);
nand U1940 (N_1940,N_1672,N_1709);
nor U1941 (N_1941,N_1665,N_1694);
and U1942 (N_1942,N_1656,N_1771);
or U1943 (N_1943,N_1627,N_1623);
and U1944 (N_1944,N_1717,N_1650);
or U1945 (N_1945,N_1698,N_1727);
nor U1946 (N_1946,N_1692,N_1669);
nor U1947 (N_1947,N_1684,N_1779);
nor U1948 (N_1948,N_1633,N_1639);
nor U1949 (N_1949,N_1786,N_1699);
nor U1950 (N_1950,N_1797,N_1720);
nand U1951 (N_1951,N_1796,N_1632);
nand U1952 (N_1952,N_1656,N_1788);
and U1953 (N_1953,N_1689,N_1691);
or U1954 (N_1954,N_1761,N_1636);
nor U1955 (N_1955,N_1732,N_1745);
xnor U1956 (N_1956,N_1677,N_1760);
or U1957 (N_1957,N_1703,N_1734);
or U1958 (N_1958,N_1696,N_1613);
nor U1959 (N_1959,N_1734,N_1606);
and U1960 (N_1960,N_1770,N_1661);
nand U1961 (N_1961,N_1793,N_1723);
and U1962 (N_1962,N_1732,N_1740);
or U1963 (N_1963,N_1628,N_1621);
and U1964 (N_1964,N_1762,N_1679);
nor U1965 (N_1965,N_1763,N_1711);
xnor U1966 (N_1966,N_1760,N_1708);
and U1967 (N_1967,N_1633,N_1615);
or U1968 (N_1968,N_1780,N_1736);
nand U1969 (N_1969,N_1724,N_1767);
or U1970 (N_1970,N_1736,N_1682);
or U1971 (N_1971,N_1781,N_1660);
xor U1972 (N_1972,N_1674,N_1742);
or U1973 (N_1973,N_1604,N_1711);
and U1974 (N_1974,N_1731,N_1650);
or U1975 (N_1975,N_1789,N_1768);
nand U1976 (N_1976,N_1691,N_1719);
and U1977 (N_1977,N_1744,N_1743);
nand U1978 (N_1978,N_1628,N_1699);
nand U1979 (N_1979,N_1667,N_1688);
nand U1980 (N_1980,N_1741,N_1637);
nor U1981 (N_1981,N_1700,N_1682);
or U1982 (N_1982,N_1769,N_1643);
and U1983 (N_1983,N_1653,N_1740);
nor U1984 (N_1984,N_1688,N_1662);
nor U1985 (N_1985,N_1681,N_1702);
nor U1986 (N_1986,N_1635,N_1793);
or U1987 (N_1987,N_1706,N_1663);
nor U1988 (N_1988,N_1741,N_1657);
nand U1989 (N_1989,N_1695,N_1659);
nand U1990 (N_1990,N_1765,N_1697);
nand U1991 (N_1991,N_1718,N_1763);
and U1992 (N_1992,N_1684,N_1608);
nand U1993 (N_1993,N_1745,N_1793);
and U1994 (N_1994,N_1794,N_1623);
or U1995 (N_1995,N_1784,N_1767);
or U1996 (N_1996,N_1790,N_1604);
or U1997 (N_1997,N_1699,N_1675);
or U1998 (N_1998,N_1642,N_1674);
nand U1999 (N_1999,N_1631,N_1600);
nand U2000 (N_2000,N_1872,N_1888);
and U2001 (N_2001,N_1905,N_1874);
or U2002 (N_2002,N_1812,N_1824);
nor U2003 (N_2003,N_1993,N_1935);
and U2004 (N_2004,N_1934,N_1909);
nor U2005 (N_2005,N_1802,N_1952);
nand U2006 (N_2006,N_1946,N_1844);
nand U2007 (N_2007,N_1890,N_1963);
and U2008 (N_2008,N_1875,N_1931);
nand U2009 (N_2009,N_1868,N_1805);
nor U2010 (N_2010,N_1886,N_1839);
nand U2011 (N_2011,N_1971,N_1806);
or U2012 (N_2012,N_1969,N_1807);
nor U2013 (N_2013,N_1895,N_1927);
or U2014 (N_2014,N_1996,N_1848);
and U2015 (N_2015,N_1871,N_1891);
or U2016 (N_2016,N_1826,N_1995);
and U2017 (N_2017,N_1833,N_1943);
nand U2018 (N_2018,N_1973,N_1831);
nand U2019 (N_2019,N_1843,N_1823);
nand U2020 (N_2020,N_1994,N_1958);
or U2021 (N_2021,N_1900,N_1878);
xor U2022 (N_2022,N_1915,N_1863);
nor U2023 (N_2023,N_1913,N_1827);
or U2024 (N_2024,N_1834,N_1870);
nor U2025 (N_2025,N_1819,N_1979);
xnor U2026 (N_2026,N_1991,N_1883);
nor U2027 (N_2027,N_1907,N_1856);
and U2028 (N_2028,N_1866,N_1939);
xnor U2029 (N_2029,N_1877,N_1904);
nor U2030 (N_2030,N_1947,N_1864);
nand U2031 (N_2031,N_1857,N_1954);
nor U2032 (N_2032,N_1912,N_1898);
nand U2033 (N_2033,N_1862,N_1876);
or U2034 (N_2034,N_1967,N_1949);
or U2035 (N_2035,N_1964,N_1985);
or U2036 (N_2036,N_1879,N_1850);
nand U2037 (N_2037,N_1817,N_1981);
nand U2038 (N_2038,N_1961,N_1861);
nand U2039 (N_2039,N_1873,N_1814);
or U2040 (N_2040,N_1899,N_1855);
and U2041 (N_2041,N_1893,N_1816);
and U2042 (N_2042,N_1923,N_1849);
nor U2043 (N_2043,N_1908,N_1976);
nor U2044 (N_2044,N_1992,N_1968);
nor U2045 (N_2045,N_1903,N_1948);
nand U2046 (N_2046,N_1922,N_1841);
and U2047 (N_2047,N_1830,N_1837);
and U2048 (N_2048,N_1988,N_1936);
and U2049 (N_2049,N_1942,N_1998);
nand U2050 (N_2050,N_1847,N_1854);
nor U2051 (N_2051,N_1938,N_1920);
or U2052 (N_2052,N_1925,N_1986);
nor U2053 (N_2053,N_1828,N_1836);
or U2054 (N_2054,N_1869,N_1808);
or U2055 (N_2055,N_1926,N_1950);
or U2056 (N_2056,N_1822,N_1880);
nor U2057 (N_2057,N_1910,N_1832);
nand U2058 (N_2058,N_1924,N_1919);
nand U2059 (N_2059,N_1937,N_1846);
or U2060 (N_2060,N_1965,N_1842);
nand U2061 (N_2061,N_1956,N_1962);
or U2062 (N_2062,N_1990,N_1881);
nand U2063 (N_2063,N_1820,N_1825);
or U2064 (N_2064,N_1940,N_1860);
and U2065 (N_2065,N_1800,N_1818);
or U2066 (N_2066,N_1972,N_1916);
nand U2067 (N_2067,N_1933,N_1957);
nor U2068 (N_2068,N_1989,N_1953);
nand U2069 (N_2069,N_1983,N_1803);
nor U2070 (N_2070,N_1918,N_1859);
and U2071 (N_2071,N_1987,N_1984);
and U2072 (N_2072,N_1884,N_1980);
and U2073 (N_2073,N_1867,N_1999);
or U2074 (N_2074,N_1889,N_1858);
and U2075 (N_2075,N_1840,N_1838);
and U2076 (N_2076,N_1917,N_1966);
and U2077 (N_2077,N_1813,N_1997);
or U2078 (N_2078,N_1932,N_1928);
or U2079 (N_2079,N_1804,N_1885);
or U2080 (N_2080,N_1851,N_1921);
and U2081 (N_2081,N_1887,N_1975);
or U2082 (N_2082,N_1929,N_1882);
and U2083 (N_2083,N_1978,N_1892);
nand U2084 (N_2084,N_1959,N_1815);
and U2085 (N_2085,N_1977,N_1951);
or U2086 (N_2086,N_1810,N_1865);
and U2087 (N_2087,N_1829,N_1930);
nand U2088 (N_2088,N_1821,N_1974);
or U2089 (N_2089,N_1911,N_1906);
or U2090 (N_2090,N_1901,N_1914);
nor U2091 (N_2091,N_1811,N_1944);
nor U2092 (N_2092,N_1852,N_1853);
nor U2093 (N_2093,N_1809,N_1960);
nor U2094 (N_2094,N_1801,N_1982);
nand U2095 (N_2095,N_1835,N_1945);
nand U2096 (N_2096,N_1970,N_1894);
nand U2097 (N_2097,N_1902,N_1955);
and U2098 (N_2098,N_1845,N_1941);
nand U2099 (N_2099,N_1896,N_1897);
and U2100 (N_2100,N_1964,N_1865);
and U2101 (N_2101,N_1851,N_1901);
and U2102 (N_2102,N_1821,N_1829);
or U2103 (N_2103,N_1990,N_1839);
nand U2104 (N_2104,N_1941,N_1879);
nor U2105 (N_2105,N_1805,N_1865);
nor U2106 (N_2106,N_1984,N_1817);
nand U2107 (N_2107,N_1926,N_1840);
nand U2108 (N_2108,N_1954,N_1859);
nand U2109 (N_2109,N_1877,N_1968);
nand U2110 (N_2110,N_1986,N_1805);
or U2111 (N_2111,N_1841,N_1943);
nor U2112 (N_2112,N_1972,N_1892);
or U2113 (N_2113,N_1935,N_1867);
or U2114 (N_2114,N_1886,N_1947);
nand U2115 (N_2115,N_1965,N_1806);
and U2116 (N_2116,N_1960,N_1980);
nand U2117 (N_2117,N_1841,N_1859);
nor U2118 (N_2118,N_1885,N_1961);
nor U2119 (N_2119,N_1956,N_1873);
and U2120 (N_2120,N_1880,N_1855);
nor U2121 (N_2121,N_1966,N_1801);
nand U2122 (N_2122,N_1863,N_1952);
nand U2123 (N_2123,N_1992,N_1839);
or U2124 (N_2124,N_1990,N_1872);
and U2125 (N_2125,N_1950,N_1851);
nand U2126 (N_2126,N_1932,N_1858);
xor U2127 (N_2127,N_1882,N_1980);
nand U2128 (N_2128,N_1855,N_1944);
nand U2129 (N_2129,N_1854,N_1922);
and U2130 (N_2130,N_1844,N_1870);
or U2131 (N_2131,N_1983,N_1809);
and U2132 (N_2132,N_1995,N_1860);
nand U2133 (N_2133,N_1861,N_1865);
nor U2134 (N_2134,N_1824,N_1989);
nand U2135 (N_2135,N_1801,N_1969);
nand U2136 (N_2136,N_1982,N_1927);
nor U2137 (N_2137,N_1889,N_1929);
nand U2138 (N_2138,N_1937,N_1971);
nor U2139 (N_2139,N_1892,N_1955);
and U2140 (N_2140,N_1979,N_1832);
or U2141 (N_2141,N_1868,N_1970);
or U2142 (N_2142,N_1977,N_1956);
nor U2143 (N_2143,N_1970,N_1952);
or U2144 (N_2144,N_1999,N_1971);
xor U2145 (N_2145,N_1889,N_1992);
nor U2146 (N_2146,N_1837,N_1965);
nor U2147 (N_2147,N_1987,N_1874);
nand U2148 (N_2148,N_1933,N_1968);
or U2149 (N_2149,N_1802,N_1860);
and U2150 (N_2150,N_1828,N_1995);
or U2151 (N_2151,N_1963,N_1982);
nor U2152 (N_2152,N_1814,N_1885);
nor U2153 (N_2153,N_1972,N_1955);
nor U2154 (N_2154,N_1845,N_1801);
xor U2155 (N_2155,N_1873,N_1886);
nand U2156 (N_2156,N_1857,N_1864);
nor U2157 (N_2157,N_1895,N_1849);
and U2158 (N_2158,N_1970,N_1957);
nor U2159 (N_2159,N_1836,N_1842);
nand U2160 (N_2160,N_1978,N_1920);
nand U2161 (N_2161,N_1838,N_1946);
nor U2162 (N_2162,N_1827,N_1894);
and U2163 (N_2163,N_1908,N_1849);
nand U2164 (N_2164,N_1921,N_1886);
or U2165 (N_2165,N_1995,N_1998);
or U2166 (N_2166,N_1876,N_1944);
nor U2167 (N_2167,N_1821,N_1826);
and U2168 (N_2168,N_1804,N_1847);
nor U2169 (N_2169,N_1910,N_1863);
nor U2170 (N_2170,N_1842,N_1824);
nor U2171 (N_2171,N_1941,N_1888);
nor U2172 (N_2172,N_1816,N_1977);
nand U2173 (N_2173,N_1845,N_1874);
or U2174 (N_2174,N_1949,N_1925);
nand U2175 (N_2175,N_1813,N_1949);
nor U2176 (N_2176,N_1989,N_1857);
and U2177 (N_2177,N_1921,N_1812);
nand U2178 (N_2178,N_1919,N_1857);
or U2179 (N_2179,N_1949,N_1906);
and U2180 (N_2180,N_1818,N_1886);
nor U2181 (N_2181,N_1948,N_1846);
nand U2182 (N_2182,N_1988,N_1885);
nand U2183 (N_2183,N_1893,N_1986);
or U2184 (N_2184,N_1928,N_1994);
xnor U2185 (N_2185,N_1966,N_1949);
and U2186 (N_2186,N_1960,N_1885);
or U2187 (N_2187,N_1913,N_1848);
nor U2188 (N_2188,N_1849,N_1822);
or U2189 (N_2189,N_1860,N_1812);
or U2190 (N_2190,N_1856,N_1884);
nor U2191 (N_2191,N_1885,N_1973);
nor U2192 (N_2192,N_1810,N_1925);
nor U2193 (N_2193,N_1923,N_1909);
nand U2194 (N_2194,N_1884,N_1933);
nand U2195 (N_2195,N_1988,N_1802);
nand U2196 (N_2196,N_1856,N_1912);
nor U2197 (N_2197,N_1954,N_1886);
or U2198 (N_2198,N_1806,N_1851);
nor U2199 (N_2199,N_1999,N_1992);
nor U2200 (N_2200,N_2150,N_2191);
or U2201 (N_2201,N_2046,N_2172);
or U2202 (N_2202,N_2096,N_2052);
nand U2203 (N_2203,N_2156,N_2059);
nor U2204 (N_2204,N_2197,N_2027);
or U2205 (N_2205,N_2148,N_2110);
or U2206 (N_2206,N_2058,N_2055);
nand U2207 (N_2207,N_2094,N_2032);
nand U2208 (N_2208,N_2029,N_2076);
nor U2209 (N_2209,N_2111,N_2003);
nor U2210 (N_2210,N_2198,N_2128);
nor U2211 (N_2211,N_2125,N_2109);
and U2212 (N_2212,N_2041,N_2031);
nand U2213 (N_2213,N_2140,N_2165);
nand U2214 (N_2214,N_2025,N_2168);
nor U2215 (N_2215,N_2135,N_2044);
and U2216 (N_2216,N_2078,N_2189);
or U2217 (N_2217,N_2097,N_2192);
nand U2218 (N_2218,N_2034,N_2186);
nor U2219 (N_2219,N_2011,N_2065);
nand U2220 (N_2220,N_2040,N_2139);
nand U2221 (N_2221,N_2091,N_2087);
nor U2222 (N_2222,N_2131,N_2007);
and U2223 (N_2223,N_2107,N_2144);
and U2224 (N_2224,N_2115,N_2101);
and U2225 (N_2225,N_2021,N_2136);
nand U2226 (N_2226,N_2106,N_2030);
and U2227 (N_2227,N_2026,N_2038);
nand U2228 (N_2228,N_2085,N_2169);
nor U2229 (N_2229,N_2105,N_2063);
or U2230 (N_2230,N_2174,N_2133);
nor U2231 (N_2231,N_2014,N_2120);
nor U2232 (N_2232,N_2162,N_2064);
nand U2233 (N_2233,N_2075,N_2121);
and U2234 (N_2234,N_2062,N_2103);
and U2235 (N_2235,N_2153,N_2193);
nor U2236 (N_2236,N_2177,N_2113);
nor U2237 (N_2237,N_2137,N_2171);
nor U2238 (N_2238,N_2123,N_2005);
and U2239 (N_2239,N_2104,N_2082);
nor U2240 (N_2240,N_2188,N_2066);
or U2241 (N_2241,N_2130,N_2024);
nor U2242 (N_2242,N_2159,N_2015);
or U2243 (N_2243,N_2028,N_2074);
nor U2244 (N_2244,N_2114,N_2000);
and U2245 (N_2245,N_2020,N_2077);
nand U2246 (N_2246,N_2184,N_2098);
and U2247 (N_2247,N_2019,N_2017);
nand U2248 (N_2248,N_2069,N_2158);
and U2249 (N_2249,N_2035,N_2146);
nand U2250 (N_2250,N_2023,N_2012);
or U2251 (N_2251,N_2187,N_2164);
nor U2252 (N_2252,N_2093,N_2185);
nand U2253 (N_2253,N_2010,N_2173);
nand U2254 (N_2254,N_2039,N_2132);
or U2255 (N_2255,N_2180,N_2002);
or U2256 (N_2256,N_2151,N_2143);
nand U2257 (N_2257,N_2089,N_2129);
nor U2258 (N_2258,N_2199,N_2149);
or U2259 (N_2259,N_2160,N_2194);
or U2260 (N_2260,N_2006,N_2141);
or U2261 (N_2261,N_2166,N_2154);
and U2262 (N_2262,N_2042,N_2086);
nand U2263 (N_2263,N_2163,N_2004);
or U2264 (N_2264,N_2155,N_2080);
and U2265 (N_2265,N_2161,N_2108);
and U2266 (N_2266,N_2182,N_2157);
xnor U2267 (N_2267,N_2001,N_2119);
and U2268 (N_2268,N_2175,N_2018);
and U2269 (N_2269,N_2099,N_2033);
and U2270 (N_2270,N_2118,N_2047);
nor U2271 (N_2271,N_2178,N_2122);
xnor U2272 (N_2272,N_2022,N_2009);
nor U2273 (N_2273,N_2124,N_2061);
nor U2274 (N_2274,N_2152,N_2037);
nor U2275 (N_2275,N_2053,N_2183);
nor U2276 (N_2276,N_2142,N_2084);
nor U2277 (N_2277,N_2054,N_2117);
or U2278 (N_2278,N_2045,N_2092);
nor U2279 (N_2279,N_2056,N_2013);
nor U2280 (N_2280,N_2179,N_2051);
nor U2281 (N_2281,N_2083,N_2079);
nor U2282 (N_2282,N_2072,N_2145);
nor U2283 (N_2283,N_2126,N_2090);
or U2284 (N_2284,N_2071,N_2100);
or U2285 (N_2285,N_2008,N_2057);
nand U2286 (N_2286,N_2176,N_2049);
or U2287 (N_2287,N_2116,N_2036);
nand U2288 (N_2288,N_2147,N_2196);
nand U2289 (N_2289,N_2190,N_2088);
or U2290 (N_2290,N_2138,N_2043);
and U2291 (N_2291,N_2068,N_2167);
nand U2292 (N_2292,N_2067,N_2112);
and U2293 (N_2293,N_2050,N_2073);
and U2294 (N_2294,N_2070,N_2060);
and U2295 (N_2295,N_2102,N_2016);
nor U2296 (N_2296,N_2170,N_2181);
nor U2297 (N_2297,N_2134,N_2048);
nand U2298 (N_2298,N_2195,N_2081);
nand U2299 (N_2299,N_2095,N_2127);
and U2300 (N_2300,N_2193,N_2073);
and U2301 (N_2301,N_2002,N_2093);
nor U2302 (N_2302,N_2040,N_2191);
and U2303 (N_2303,N_2188,N_2074);
and U2304 (N_2304,N_2030,N_2109);
and U2305 (N_2305,N_2002,N_2066);
or U2306 (N_2306,N_2072,N_2042);
nor U2307 (N_2307,N_2083,N_2119);
nand U2308 (N_2308,N_2174,N_2083);
nor U2309 (N_2309,N_2165,N_2191);
nor U2310 (N_2310,N_2198,N_2137);
nor U2311 (N_2311,N_2174,N_2002);
or U2312 (N_2312,N_2137,N_2168);
or U2313 (N_2313,N_2180,N_2032);
or U2314 (N_2314,N_2121,N_2074);
and U2315 (N_2315,N_2094,N_2155);
or U2316 (N_2316,N_2042,N_2140);
nand U2317 (N_2317,N_2067,N_2180);
nand U2318 (N_2318,N_2010,N_2132);
or U2319 (N_2319,N_2002,N_2139);
nor U2320 (N_2320,N_2090,N_2132);
nand U2321 (N_2321,N_2078,N_2161);
or U2322 (N_2322,N_2111,N_2008);
and U2323 (N_2323,N_2195,N_2022);
or U2324 (N_2324,N_2015,N_2078);
and U2325 (N_2325,N_2142,N_2018);
or U2326 (N_2326,N_2032,N_2188);
nor U2327 (N_2327,N_2166,N_2099);
or U2328 (N_2328,N_2080,N_2024);
and U2329 (N_2329,N_2118,N_2043);
and U2330 (N_2330,N_2162,N_2149);
or U2331 (N_2331,N_2048,N_2031);
or U2332 (N_2332,N_2171,N_2172);
and U2333 (N_2333,N_2073,N_2016);
nor U2334 (N_2334,N_2100,N_2062);
nand U2335 (N_2335,N_2178,N_2078);
nor U2336 (N_2336,N_2172,N_2174);
and U2337 (N_2337,N_2100,N_2163);
nand U2338 (N_2338,N_2014,N_2143);
nand U2339 (N_2339,N_2145,N_2044);
xnor U2340 (N_2340,N_2028,N_2017);
or U2341 (N_2341,N_2109,N_2096);
nand U2342 (N_2342,N_2023,N_2113);
or U2343 (N_2343,N_2193,N_2032);
nor U2344 (N_2344,N_2187,N_2048);
and U2345 (N_2345,N_2156,N_2096);
nand U2346 (N_2346,N_2026,N_2090);
nor U2347 (N_2347,N_2044,N_2071);
or U2348 (N_2348,N_2151,N_2153);
or U2349 (N_2349,N_2028,N_2151);
or U2350 (N_2350,N_2195,N_2182);
and U2351 (N_2351,N_2120,N_2044);
or U2352 (N_2352,N_2173,N_2050);
and U2353 (N_2353,N_2138,N_2080);
or U2354 (N_2354,N_2176,N_2037);
nand U2355 (N_2355,N_2181,N_2135);
nand U2356 (N_2356,N_2039,N_2099);
nor U2357 (N_2357,N_2049,N_2187);
nor U2358 (N_2358,N_2096,N_2100);
or U2359 (N_2359,N_2151,N_2073);
nand U2360 (N_2360,N_2116,N_2132);
and U2361 (N_2361,N_2051,N_2128);
or U2362 (N_2362,N_2155,N_2110);
or U2363 (N_2363,N_2000,N_2118);
nor U2364 (N_2364,N_2039,N_2138);
and U2365 (N_2365,N_2050,N_2051);
and U2366 (N_2366,N_2136,N_2042);
and U2367 (N_2367,N_2167,N_2011);
or U2368 (N_2368,N_2010,N_2195);
or U2369 (N_2369,N_2047,N_2058);
nor U2370 (N_2370,N_2154,N_2014);
nor U2371 (N_2371,N_2133,N_2022);
or U2372 (N_2372,N_2063,N_2100);
nand U2373 (N_2373,N_2149,N_2025);
nand U2374 (N_2374,N_2034,N_2195);
and U2375 (N_2375,N_2191,N_2049);
nand U2376 (N_2376,N_2132,N_2123);
nor U2377 (N_2377,N_2193,N_2141);
and U2378 (N_2378,N_2078,N_2083);
nor U2379 (N_2379,N_2133,N_2103);
nor U2380 (N_2380,N_2091,N_2130);
nand U2381 (N_2381,N_2100,N_2138);
nand U2382 (N_2382,N_2085,N_2033);
or U2383 (N_2383,N_2144,N_2164);
or U2384 (N_2384,N_2026,N_2021);
and U2385 (N_2385,N_2110,N_2096);
and U2386 (N_2386,N_2072,N_2057);
or U2387 (N_2387,N_2124,N_2006);
nor U2388 (N_2388,N_2156,N_2164);
or U2389 (N_2389,N_2097,N_2029);
and U2390 (N_2390,N_2170,N_2037);
nor U2391 (N_2391,N_2172,N_2112);
nor U2392 (N_2392,N_2146,N_2047);
or U2393 (N_2393,N_2006,N_2036);
nor U2394 (N_2394,N_2053,N_2114);
or U2395 (N_2395,N_2195,N_2177);
nor U2396 (N_2396,N_2030,N_2098);
and U2397 (N_2397,N_2149,N_2023);
and U2398 (N_2398,N_2183,N_2015);
nor U2399 (N_2399,N_2086,N_2106);
and U2400 (N_2400,N_2203,N_2365);
nand U2401 (N_2401,N_2294,N_2230);
nand U2402 (N_2402,N_2289,N_2213);
nor U2403 (N_2403,N_2275,N_2246);
nand U2404 (N_2404,N_2308,N_2373);
nor U2405 (N_2405,N_2303,N_2325);
xor U2406 (N_2406,N_2359,N_2361);
or U2407 (N_2407,N_2360,N_2341);
or U2408 (N_2408,N_2277,N_2209);
nand U2409 (N_2409,N_2264,N_2390);
nor U2410 (N_2410,N_2261,N_2336);
or U2411 (N_2411,N_2357,N_2266);
and U2412 (N_2412,N_2338,N_2257);
or U2413 (N_2413,N_2241,N_2304);
nor U2414 (N_2414,N_2355,N_2399);
or U2415 (N_2415,N_2291,N_2343);
nor U2416 (N_2416,N_2340,N_2206);
or U2417 (N_2417,N_2347,N_2364);
or U2418 (N_2418,N_2380,N_2394);
or U2419 (N_2419,N_2398,N_2368);
and U2420 (N_2420,N_2353,N_2306);
nand U2421 (N_2421,N_2218,N_2358);
and U2422 (N_2422,N_2297,N_2345);
or U2423 (N_2423,N_2263,N_2216);
and U2424 (N_2424,N_2256,N_2249);
and U2425 (N_2425,N_2299,N_2222);
and U2426 (N_2426,N_2284,N_2329);
nand U2427 (N_2427,N_2271,N_2248);
and U2428 (N_2428,N_2335,N_2302);
nand U2429 (N_2429,N_2349,N_2370);
nand U2430 (N_2430,N_2376,N_2296);
or U2431 (N_2431,N_2255,N_2348);
and U2432 (N_2432,N_2278,N_2372);
and U2433 (N_2433,N_2207,N_2362);
nand U2434 (N_2434,N_2307,N_2251);
and U2435 (N_2435,N_2392,N_2332);
nor U2436 (N_2436,N_2290,N_2310);
nand U2437 (N_2437,N_2217,N_2272);
and U2438 (N_2438,N_2258,N_2396);
nor U2439 (N_2439,N_2383,N_2238);
nand U2440 (N_2440,N_2267,N_2298);
or U2441 (N_2441,N_2268,N_2344);
xor U2442 (N_2442,N_2242,N_2225);
nand U2443 (N_2443,N_2265,N_2250);
nor U2444 (N_2444,N_2226,N_2346);
and U2445 (N_2445,N_2269,N_2292);
nand U2446 (N_2446,N_2322,N_2293);
and U2447 (N_2447,N_2386,N_2210);
nand U2448 (N_2448,N_2356,N_2212);
nor U2449 (N_2449,N_2211,N_2286);
or U2450 (N_2450,N_2224,N_2323);
nor U2451 (N_2451,N_2252,N_2235);
or U2452 (N_2452,N_2371,N_2244);
and U2453 (N_2453,N_2321,N_2228);
and U2454 (N_2454,N_2202,N_2351);
nor U2455 (N_2455,N_2220,N_2367);
nor U2456 (N_2456,N_2334,N_2350);
nand U2457 (N_2457,N_2391,N_2245);
and U2458 (N_2458,N_2389,N_2254);
nor U2459 (N_2459,N_2208,N_2231);
or U2460 (N_2460,N_2382,N_2219);
or U2461 (N_2461,N_2229,N_2273);
and U2462 (N_2462,N_2259,N_2342);
nor U2463 (N_2463,N_2328,N_2387);
nor U2464 (N_2464,N_2317,N_2375);
or U2465 (N_2465,N_2354,N_2305);
or U2466 (N_2466,N_2232,N_2333);
or U2467 (N_2467,N_2320,N_2221);
or U2468 (N_2468,N_2301,N_2227);
and U2469 (N_2469,N_2295,N_2237);
or U2470 (N_2470,N_2378,N_2287);
or U2471 (N_2471,N_2214,N_2339);
and U2472 (N_2472,N_2201,N_2234);
nand U2473 (N_2473,N_2313,N_2312);
or U2474 (N_2474,N_2282,N_2260);
nor U2475 (N_2475,N_2337,N_2243);
or U2476 (N_2476,N_2377,N_2326);
nand U2477 (N_2477,N_2276,N_2300);
nand U2478 (N_2478,N_2395,N_2324);
or U2479 (N_2479,N_2288,N_2270);
nor U2480 (N_2480,N_2384,N_2200);
nor U2481 (N_2481,N_2215,N_2393);
and U2482 (N_2482,N_2374,N_2285);
and U2483 (N_2483,N_2240,N_2247);
nand U2484 (N_2484,N_2205,N_2204);
and U2485 (N_2485,N_2331,N_2381);
nand U2486 (N_2486,N_2388,N_2318);
and U2487 (N_2487,N_2262,N_2352);
nor U2488 (N_2488,N_2283,N_2280);
or U2489 (N_2489,N_2274,N_2239);
or U2490 (N_2490,N_2279,N_2253);
nor U2491 (N_2491,N_2369,N_2315);
nand U2492 (N_2492,N_2281,N_2233);
and U2493 (N_2493,N_2330,N_2314);
or U2494 (N_2494,N_2319,N_2363);
or U2495 (N_2495,N_2366,N_2316);
nand U2496 (N_2496,N_2223,N_2236);
and U2497 (N_2497,N_2379,N_2311);
nor U2498 (N_2498,N_2327,N_2397);
or U2499 (N_2499,N_2385,N_2309);
or U2500 (N_2500,N_2233,N_2336);
nor U2501 (N_2501,N_2308,N_2248);
and U2502 (N_2502,N_2275,N_2319);
or U2503 (N_2503,N_2333,N_2388);
or U2504 (N_2504,N_2350,N_2244);
nor U2505 (N_2505,N_2223,N_2376);
and U2506 (N_2506,N_2312,N_2287);
nor U2507 (N_2507,N_2261,N_2322);
nand U2508 (N_2508,N_2264,N_2317);
nor U2509 (N_2509,N_2386,N_2340);
or U2510 (N_2510,N_2283,N_2284);
nand U2511 (N_2511,N_2245,N_2335);
nand U2512 (N_2512,N_2299,N_2366);
and U2513 (N_2513,N_2223,N_2345);
nor U2514 (N_2514,N_2364,N_2301);
nor U2515 (N_2515,N_2326,N_2365);
or U2516 (N_2516,N_2310,N_2301);
or U2517 (N_2517,N_2207,N_2242);
nand U2518 (N_2518,N_2274,N_2347);
and U2519 (N_2519,N_2250,N_2280);
nor U2520 (N_2520,N_2391,N_2271);
nand U2521 (N_2521,N_2390,N_2347);
and U2522 (N_2522,N_2217,N_2382);
or U2523 (N_2523,N_2383,N_2216);
nand U2524 (N_2524,N_2322,N_2350);
nor U2525 (N_2525,N_2337,N_2209);
nor U2526 (N_2526,N_2213,N_2347);
nor U2527 (N_2527,N_2282,N_2228);
nand U2528 (N_2528,N_2315,N_2399);
nor U2529 (N_2529,N_2346,N_2241);
nor U2530 (N_2530,N_2255,N_2233);
nand U2531 (N_2531,N_2281,N_2285);
nor U2532 (N_2532,N_2330,N_2296);
or U2533 (N_2533,N_2341,N_2369);
and U2534 (N_2534,N_2260,N_2209);
or U2535 (N_2535,N_2289,N_2225);
and U2536 (N_2536,N_2287,N_2256);
nor U2537 (N_2537,N_2391,N_2352);
nor U2538 (N_2538,N_2278,N_2369);
nand U2539 (N_2539,N_2363,N_2259);
or U2540 (N_2540,N_2261,N_2304);
or U2541 (N_2541,N_2264,N_2298);
and U2542 (N_2542,N_2234,N_2301);
or U2543 (N_2543,N_2260,N_2301);
and U2544 (N_2544,N_2217,N_2391);
nor U2545 (N_2545,N_2333,N_2396);
nand U2546 (N_2546,N_2380,N_2231);
nor U2547 (N_2547,N_2355,N_2381);
or U2548 (N_2548,N_2258,N_2320);
nor U2549 (N_2549,N_2397,N_2303);
and U2550 (N_2550,N_2315,N_2270);
or U2551 (N_2551,N_2297,N_2367);
or U2552 (N_2552,N_2244,N_2361);
nand U2553 (N_2553,N_2309,N_2269);
and U2554 (N_2554,N_2364,N_2202);
nand U2555 (N_2555,N_2367,N_2336);
nor U2556 (N_2556,N_2258,N_2294);
nand U2557 (N_2557,N_2373,N_2228);
or U2558 (N_2558,N_2336,N_2313);
or U2559 (N_2559,N_2293,N_2388);
nand U2560 (N_2560,N_2249,N_2355);
nand U2561 (N_2561,N_2255,N_2217);
nor U2562 (N_2562,N_2301,N_2362);
nand U2563 (N_2563,N_2223,N_2397);
or U2564 (N_2564,N_2253,N_2399);
or U2565 (N_2565,N_2340,N_2234);
nor U2566 (N_2566,N_2296,N_2231);
nand U2567 (N_2567,N_2383,N_2281);
or U2568 (N_2568,N_2252,N_2242);
or U2569 (N_2569,N_2361,N_2372);
nand U2570 (N_2570,N_2232,N_2284);
or U2571 (N_2571,N_2320,N_2317);
and U2572 (N_2572,N_2226,N_2285);
nor U2573 (N_2573,N_2309,N_2241);
and U2574 (N_2574,N_2312,N_2334);
or U2575 (N_2575,N_2330,N_2380);
nand U2576 (N_2576,N_2365,N_2226);
nand U2577 (N_2577,N_2303,N_2284);
nor U2578 (N_2578,N_2274,N_2300);
and U2579 (N_2579,N_2222,N_2304);
and U2580 (N_2580,N_2242,N_2227);
nand U2581 (N_2581,N_2282,N_2345);
or U2582 (N_2582,N_2241,N_2248);
and U2583 (N_2583,N_2331,N_2206);
nand U2584 (N_2584,N_2230,N_2235);
or U2585 (N_2585,N_2372,N_2331);
nor U2586 (N_2586,N_2366,N_2342);
and U2587 (N_2587,N_2313,N_2346);
nand U2588 (N_2588,N_2251,N_2236);
nand U2589 (N_2589,N_2257,N_2242);
nor U2590 (N_2590,N_2399,N_2333);
or U2591 (N_2591,N_2328,N_2302);
nor U2592 (N_2592,N_2306,N_2363);
or U2593 (N_2593,N_2364,N_2206);
nor U2594 (N_2594,N_2320,N_2321);
nor U2595 (N_2595,N_2267,N_2264);
and U2596 (N_2596,N_2211,N_2307);
or U2597 (N_2597,N_2358,N_2250);
and U2598 (N_2598,N_2253,N_2255);
nand U2599 (N_2599,N_2354,N_2322);
or U2600 (N_2600,N_2517,N_2501);
and U2601 (N_2601,N_2494,N_2569);
or U2602 (N_2602,N_2568,N_2413);
and U2603 (N_2603,N_2498,N_2461);
or U2604 (N_2604,N_2554,N_2440);
nand U2605 (N_2605,N_2538,N_2589);
nor U2606 (N_2606,N_2426,N_2452);
nand U2607 (N_2607,N_2504,N_2435);
or U2608 (N_2608,N_2577,N_2508);
nand U2609 (N_2609,N_2427,N_2542);
and U2610 (N_2610,N_2447,N_2464);
or U2611 (N_2611,N_2527,N_2561);
nor U2612 (N_2612,N_2592,N_2553);
and U2613 (N_2613,N_2513,N_2456);
nor U2614 (N_2614,N_2523,N_2436);
nand U2615 (N_2615,N_2432,N_2598);
nand U2616 (N_2616,N_2419,N_2516);
and U2617 (N_2617,N_2591,N_2430);
or U2618 (N_2618,N_2487,N_2422);
nor U2619 (N_2619,N_2578,N_2488);
and U2620 (N_2620,N_2573,N_2449);
nand U2621 (N_2621,N_2550,N_2532);
nand U2622 (N_2622,N_2421,N_2505);
or U2623 (N_2623,N_2511,N_2521);
and U2624 (N_2624,N_2434,N_2579);
and U2625 (N_2625,N_2540,N_2549);
and U2626 (N_2626,N_2567,N_2547);
and U2627 (N_2627,N_2481,N_2507);
or U2628 (N_2628,N_2512,N_2437);
or U2629 (N_2629,N_2420,N_2588);
nor U2630 (N_2630,N_2424,N_2402);
and U2631 (N_2631,N_2478,N_2428);
nand U2632 (N_2632,N_2460,N_2552);
or U2633 (N_2633,N_2454,N_2476);
nor U2634 (N_2634,N_2453,N_2526);
and U2635 (N_2635,N_2416,N_2575);
nor U2636 (N_2636,N_2520,N_2502);
or U2637 (N_2637,N_2403,N_2559);
or U2638 (N_2638,N_2471,N_2407);
and U2639 (N_2639,N_2572,N_2558);
nor U2640 (N_2640,N_2596,N_2586);
nor U2641 (N_2641,N_2433,N_2551);
nor U2642 (N_2642,N_2423,N_2491);
nand U2643 (N_2643,N_2555,N_2493);
nor U2644 (N_2644,N_2593,N_2418);
nor U2645 (N_2645,N_2534,N_2541);
nor U2646 (N_2646,N_2597,N_2484);
or U2647 (N_2647,N_2480,N_2451);
or U2648 (N_2648,N_2510,N_2576);
nand U2649 (N_2649,N_2443,N_2495);
nand U2650 (N_2650,N_2408,N_2528);
nor U2651 (N_2651,N_2529,N_2485);
nand U2652 (N_2652,N_2470,N_2429);
nor U2653 (N_2653,N_2524,N_2531);
nor U2654 (N_2654,N_2455,N_2457);
nand U2655 (N_2655,N_2571,N_2448);
nor U2656 (N_2656,N_2560,N_2506);
or U2657 (N_2657,N_2545,N_2565);
nand U2658 (N_2658,N_2439,N_2497);
or U2659 (N_2659,N_2445,N_2458);
nand U2660 (N_2660,N_2441,N_2486);
and U2661 (N_2661,N_2570,N_2489);
nand U2662 (N_2662,N_2400,N_2466);
or U2663 (N_2663,N_2406,N_2539);
and U2664 (N_2664,N_2474,N_2404);
nand U2665 (N_2665,N_2412,N_2543);
nand U2666 (N_2666,N_2546,N_2515);
or U2667 (N_2667,N_2467,N_2409);
nor U2668 (N_2668,N_2450,N_2425);
or U2669 (N_2669,N_2564,N_2465);
nor U2670 (N_2670,N_2415,N_2496);
nand U2671 (N_2671,N_2584,N_2522);
nand U2672 (N_2672,N_2463,N_2414);
and U2673 (N_2673,N_2599,N_2411);
or U2674 (N_2674,N_2580,N_2509);
and U2675 (N_2675,N_2535,N_2438);
or U2676 (N_2676,N_2525,N_2590);
or U2677 (N_2677,N_2533,N_2556);
nand U2678 (N_2678,N_2574,N_2477);
or U2679 (N_2679,N_2410,N_2500);
and U2680 (N_2680,N_2469,N_2479);
or U2681 (N_2681,N_2583,N_2405);
or U2682 (N_2682,N_2459,N_2446);
nor U2683 (N_2683,N_2518,N_2431);
or U2684 (N_2684,N_2581,N_2537);
nand U2685 (N_2685,N_2401,N_2492);
nand U2686 (N_2686,N_2462,N_2499);
nand U2687 (N_2687,N_2503,N_2548);
or U2688 (N_2688,N_2562,N_2473);
nand U2689 (N_2689,N_2536,N_2594);
or U2690 (N_2690,N_2595,N_2468);
nand U2691 (N_2691,N_2566,N_2530);
or U2692 (N_2692,N_2482,N_2442);
nand U2693 (N_2693,N_2417,N_2563);
or U2694 (N_2694,N_2557,N_2483);
nand U2695 (N_2695,N_2475,N_2472);
nor U2696 (N_2696,N_2585,N_2444);
and U2697 (N_2697,N_2490,N_2519);
nor U2698 (N_2698,N_2514,N_2587);
or U2699 (N_2699,N_2544,N_2582);
nand U2700 (N_2700,N_2480,N_2568);
nor U2701 (N_2701,N_2548,N_2481);
nor U2702 (N_2702,N_2485,N_2555);
nand U2703 (N_2703,N_2579,N_2421);
or U2704 (N_2704,N_2434,N_2598);
or U2705 (N_2705,N_2456,N_2426);
or U2706 (N_2706,N_2490,N_2430);
or U2707 (N_2707,N_2437,N_2414);
and U2708 (N_2708,N_2427,N_2401);
nand U2709 (N_2709,N_2532,N_2534);
or U2710 (N_2710,N_2599,N_2569);
and U2711 (N_2711,N_2479,N_2444);
and U2712 (N_2712,N_2478,N_2461);
nand U2713 (N_2713,N_2596,N_2550);
nand U2714 (N_2714,N_2493,N_2536);
or U2715 (N_2715,N_2527,N_2430);
or U2716 (N_2716,N_2518,N_2589);
nand U2717 (N_2717,N_2592,N_2472);
or U2718 (N_2718,N_2434,N_2486);
nor U2719 (N_2719,N_2464,N_2443);
nand U2720 (N_2720,N_2508,N_2530);
and U2721 (N_2721,N_2447,N_2460);
or U2722 (N_2722,N_2525,N_2486);
and U2723 (N_2723,N_2479,N_2520);
and U2724 (N_2724,N_2402,N_2596);
nand U2725 (N_2725,N_2546,N_2445);
nor U2726 (N_2726,N_2452,N_2507);
nor U2727 (N_2727,N_2431,N_2517);
or U2728 (N_2728,N_2581,N_2406);
nor U2729 (N_2729,N_2409,N_2418);
nand U2730 (N_2730,N_2447,N_2569);
and U2731 (N_2731,N_2441,N_2460);
and U2732 (N_2732,N_2468,N_2558);
nand U2733 (N_2733,N_2459,N_2486);
and U2734 (N_2734,N_2547,N_2413);
nand U2735 (N_2735,N_2482,N_2547);
nand U2736 (N_2736,N_2408,N_2537);
or U2737 (N_2737,N_2551,N_2502);
or U2738 (N_2738,N_2496,N_2515);
or U2739 (N_2739,N_2538,N_2453);
and U2740 (N_2740,N_2498,N_2556);
or U2741 (N_2741,N_2525,N_2579);
or U2742 (N_2742,N_2474,N_2589);
nor U2743 (N_2743,N_2469,N_2591);
or U2744 (N_2744,N_2472,N_2421);
or U2745 (N_2745,N_2557,N_2451);
or U2746 (N_2746,N_2435,N_2594);
and U2747 (N_2747,N_2436,N_2511);
nor U2748 (N_2748,N_2412,N_2558);
or U2749 (N_2749,N_2597,N_2435);
and U2750 (N_2750,N_2527,N_2544);
and U2751 (N_2751,N_2542,N_2445);
nand U2752 (N_2752,N_2435,N_2485);
or U2753 (N_2753,N_2466,N_2475);
or U2754 (N_2754,N_2494,N_2544);
nor U2755 (N_2755,N_2430,N_2474);
nor U2756 (N_2756,N_2558,N_2548);
nor U2757 (N_2757,N_2443,N_2580);
or U2758 (N_2758,N_2431,N_2597);
nor U2759 (N_2759,N_2574,N_2415);
and U2760 (N_2760,N_2556,N_2521);
nor U2761 (N_2761,N_2553,N_2403);
nand U2762 (N_2762,N_2596,N_2462);
or U2763 (N_2763,N_2516,N_2477);
nor U2764 (N_2764,N_2581,N_2422);
and U2765 (N_2765,N_2483,N_2417);
nand U2766 (N_2766,N_2503,N_2580);
nor U2767 (N_2767,N_2487,N_2518);
nand U2768 (N_2768,N_2567,N_2451);
or U2769 (N_2769,N_2505,N_2506);
and U2770 (N_2770,N_2523,N_2442);
xnor U2771 (N_2771,N_2429,N_2519);
and U2772 (N_2772,N_2545,N_2425);
nand U2773 (N_2773,N_2473,N_2587);
nor U2774 (N_2774,N_2422,N_2449);
or U2775 (N_2775,N_2474,N_2414);
and U2776 (N_2776,N_2437,N_2575);
nand U2777 (N_2777,N_2594,N_2480);
and U2778 (N_2778,N_2560,N_2425);
nand U2779 (N_2779,N_2598,N_2562);
or U2780 (N_2780,N_2467,N_2570);
nor U2781 (N_2781,N_2501,N_2533);
or U2782 (N_2782,N_2588,N_2400);
or U2783 (N_2783,N_2472,N_2461);
or U2784 (N_2784,N_2428,N_2555);
nand U2785 (N_2785,N_2553,N_2466);
nand U2786 (N_2786,N_2561,N_2512);
or U2787 (N_2787,N_2583,N_2463);
and U2788 (N_2788,N_2596,N_2421);
nor U2789 (N_2789,N_2432,N_2595);
and U2790 (N_2790,N_2475,N_2539);
and U2791 (N_2791,N_2526,N_2519);
nor U2792 (N_2792,N_2502,N_2548);
nand U2793 (N_2793,N_2596,N_2515);
nand U2794 (N_2794,N_2579,N_2508);
nand U2795 (N_2795,N_2484,N_2489);
or U2796 (N_2796,N_2498,N_2526);
and U2797 (N_2797,N_2507,N_2416);
and U2798 (N_2798,N_2416,N_2407);
and U2799 (N_2799,N_2555,N_2459);
and U2800 (N_2800,N_2722,N_2602);
nand U2801 (N_2801,N_2638,N_2743);
or U2802 (N_2802,N_2697,N_2706);
or U2803 (N_2803,N_2615,N_2704);
or U2804 (N_2804,N_2791,N_2772);
nor U2805 (N_2805,N_2604,N_2628);
and U2806 (N_2806,N_2789,N_2686);
and U2807 (N_2807,N_2627,N_2702);
nor U2808 (N_2808,N_2799,N_2666);
nor U2809 (N_2809,N_2784,N_2732);
nand U2810 (N_2810,N_2660,N_2768);
nand U2811 (N_2811,N_2671,N_2661);
or U2812 (N_2812,N_2770,N_2696);
and U2813 (N_2813,N_2774,N_2657);
or U2814 (N_2814,N_2796,N_2700);
or U2815 (N_2815,N_2771,N_2727);
or U2816 (N_2816,N_2793,N_2668);
or U2817 (N_2817,N_2609,N_2755);
nor U2818 (N_2818,N_2788,N_2699);
nand U2819 (N_2819,N_2749,N_2659);
nand U2820 (N_2820,N_2783,N_2792);
nor U2821 (N_2821,N_2640,N_2782);
or U2822 (N_2822,N_2736,N_2693);
nand U2823 (N_2823,N_2618,N_2787);
nand U2824 (N_2824,N_2712,N_2718);
nor U2825 (N_2825,N_2790,N_2717);
xnor U2826 (N_2826,N_2601,N_2778);
nor U2827 (N_2827,N_2674,N_2715);
nor U2828 (N_2828,N_2742,N_2623);
or U2829 (N_2829,N_2707,N_2720);
nor U2830 (N_2830,N_2769,N_2748);
or U2831 (N_2831,N_2766,N_2621);
and U2832 (N_2832,N_2747,N_2738);
nor U2833 (N_2833,N_2701,N_2635);
nand U2834 (N_2834,N_2681,N_2777);
nand U2835 (N_2835,N_2677,N_2779);
nor U2836 (N_2836,N_2705,N_2644);
nor U2837 (N_2837,N_2654,N_2667);
nor U2838 (N_2838,N_2751,N_2687);
nand U2839 (N_2839,N_2679,N_2762);
nor U2840 (N_2840,N_2685,N_2750);
or U2841 (N_2841,N_2694,N_2690);
and U2842 (N_2842,N_2645,N_2757);
or U2843 (N_2843,N_2622,N_2613);
nand U2844 (N_2844,N_2663,N_2643);
nand U2845 (N_2845,N_2767,N_2775);
xor U2846 (N_2846,N_2744,N_2678);
nand U2847 (N_2847,N_2631,N_2683);
nand U2848 (N_2848,N_2721,N_2676);
nand U2849 (N_2849,N_2633,N_2608);
and U2850 (N_2850,N_2781,N_2626);
nand U2851 (N_2851,N_2662,N_2675);
or U2852 (N_2852,N_2795,N_2763);
nor U2853 (N_2853,N_2632,N_2619);
nor U2854 (N_2854,N_2646,N_2665);
nand U2855 (N_2855,N_2647,N_2691);
and U2856 (N_2856,N_2708,N_2612);
and U2857 (N_2857,N_2656,N_2610);
and U2858 (N_2858,N_2695,N_2684);
and U2859 (N_2859,N_2759,N_2639);
nor U2860 (N_2860,N_2741,N_2620);
nor U2861 (N_2861,N_2740,N_2724);
nand U2862 (N_2862,N_2710,N_2737);
and U2863 (N_2863,N_2669,N_2758);
and U2864 (N_2864,N_2607,N_2786);
nor U2865 (N_2865,N_2765,N_2703);
or U2866 (N_2866,N_2735,N_2723);
or U2867 (N_2867,N_2719,N_2733);
and U2868 (N_2868,N_2606,N_2729);
and U2869 (N_2869,N_2655,N_2726);
nand U2870 (N_2870,N_2746,N_2734);
and U2871 (N_2871,N_2714,N_2670);
or U2872 (N_2872,N_2754,N_2652);
or U2873 (N_2873,N_2653,N_2756);
or U2874 (N_2874,N_2689,N_2611);
nor U2875 (N_2875,N_2629,N_2739);
and U2876 (N_2876,N_2630,N_2673);
nand U2877 (N_2877,N_2680,N_2634);
nor U2878 (N_2878,N_2711,N_2725);
nor U2879 (N_2879,N_2730,N_2637);
or U2880 (N_2880,N_2745,N_2753);
nor U2881 (N_2881,N_2785,N_2650);
nor U2882 (N_2882,N_2617,N_2773);
nand U2883 (N_2883,N_2648,N_2692);
nand U2884 (N_2884,N_2651,N_2641);
nor U2885 (N_2885,N_2752,N_2603);
or U2886 (N_2886,N_2649,N_2600);
or U2887 (N_2887,N_2709,N_2624);
nor U2888 (N_2888,N_2797,N_2794);
nand U2889 (N_2889,N_2713,N_2658);
and U2890 (N_2890,N_2761,N_2672);
or U2891 (N_2891,N_2698,N_2636);
nor U2892 (N_2892,N_2716,N_2760);
or U2893 (N_2893,N_2798,N_2664);
nand U2894 (N_2894,N_2780,N_2642);
and U2895 (N_2895,N_2605,N_2776);
and U2896 (N_2896,N_2614,N_2764);
and U2897 (N_2897,N_2728,N_2688);
and U2898 (N_2898,N_2731,N_2616);
nand U2899 (N_2899,N_2625,N_2682);
nand U2900 (N_2900,N_2750,N_2739);
xor U2901 (N_2901,N_2783,N_2721);
nor U2902 (N_2902,N_2694,N_2649);
nand U2903 (N_2903,N_2672,N_2769);
nand U2904 (N_2904,N_2616,N_2730);
or U2905 (N_2905,N_2766,N_2660);
and U2906 (N_2906,N_2786,N_2664);
and U2907 (N_2907,N_2676,N_2787);
and U2908 (N_2908,N_2608,N_2680);
nand U2909 (N_2909,N_2638,N_2617);
and U2910 (N_2910,N_2716,N_2732);
nor U2911 (N_2911,N_2619,N_2766);
nand U2912 (N_2912,N_2686,N_2727);
nand U2913 (N_2913,N_2664,N_2657);
nand U2914 (N_2914,N_2688,N_2614);
or U2915 (N_2915,N_2645,N_2722);
and U2916 (N_2916,N_2717,N_2657);
and U2917 (N_2917,N_2636,N_2601);
or U2918 (N_2918,N_2659,N_2721);
nand U2919 (N_2919,N_2707,N_2709);
or U2920 (N_2920,N_2651,N_2778);
and U2921 (N_2921,N_2669,N_2763);
and U2922 (N_2922,N_2638,N_2729);
nand U2923 (N_2923,N_2792,N_2600);
nand U2924 (N_2924,N_2724,N_2714);
nor U2925 (N_2925,N_2627,N_2713);
and U2926 (N_2926,N_2722,N_2757);
and U2927 (N_2927,N_2713,N_2606);
and U2928 (N_2928,N_2727,N_2642);
and U2929 (N_2929,N_2665,N_2611);
or U2930 (N_2930,N_2726,N_2650);
nand U2931 (N_2931,N_2772,N_2756);
nor U2932 (N_2932,N_2640,N_2725);
nand U2933 (N_2933,N_2666,N_2655);
nor U2934 (N_2934,N_2642,N_2795);
or U2935 (N_2935,N_2756,N_2642);
and U2936 (N_2936,N_2772,N_2718);
or U2937 (N_2937,N_2772,N_2774);
nand U2938 (N_2938,N_2723,N_2700);
and U2939 (N_2939,N_2728,N_2740);
nand U2940 (N_2940,N_2675,N_2703);
nand U2941 (N_2941,N_2746,N_2614);
nor U2942 (N_2942,N_2764,N_2757);
nand U2943 (N_2943,N_2685,N_2645);
xnor U2944 (N_2944,N_2669,N_2643);
or U2945 (N_2945,N_2671,N_2708);
nor U2946 (N_2946,N_2782,N_2766);
or U2947 (N_2947,N_2632,N_2614);
nor U2948 (N_2948,N_2691,N_2761);
and U2949 (N_2949,N_2716,N_2767);
and U2950 (N_2950,N_2608,N_2761);
nor U2951 (N_2951,N_2638,N_2762);
and U2952 (N_2952,N_2757,N_2680);
nor U2953 (N_2953,N_2765,N_2779);
or U2954 (N_2954,N_2611,N_2644);
nor U2955 (N_2955,N_2785,N_2727);
or U2956 (N_2956,N_2770,N_2718);
nor U2957 (N_2957,N_2628,N_2708);
or U2958 (N_2958,N_2751,N_2644);
xor U2959 (N_2959,N_2710,N_2624);
nor U2960 (N_2960,N_2668,N_2753);
and U2961 (N_2961,N_2630,N_2676);
and U2962 (N_2962,N_2601,N_2699);
or U2963 (N_2963,N_2714,N_2655);
nor U2964 (N_2964,N_2602,N_2795);
or U2965 (N_2965,N_2772,N_2767);
and U2966 (N_2966,N_2668,N_2663);
or U2967 (N_2967,N_2644,N_2788);
and U2968 (N_2968,N_2619,N_2608);
and U2969 (N_2969,N_2751,N_2661);
and U2970 (N_2970,N_2611,N_2636);
or U2971 (N_2971,N_2654,N_2774);
nor U2972 (N_2972,N_2763,N_2641);
and U2973 (N_2973,N_2609,N_2709);
or U2974 (N_2974,N_2758,N_2750);
nand U2975 (N_2975,N_2749,N_2622);
nor U2976 (N_2976,N_2628,N_2685);
nor U2977 (N_2977,N_2608,N_2651);
and U2978 (N_2978,N_2733,N_2644);
and U2979 (N_2979,N_2688,N_2711);
nand U2980 (N_2980,N_2780,N_2709);
nor U2981 (N_2981,N_2795,N_2673);
or U2982 (N_2982,N_2700,N_2621);
nand U2983 (N_2983,N_2789,N_2620);
or U2984 (N_2984,N_2779,N_2661);
or U2985 (N_2985,N_2751,N_2668);
and U2986 (N_2986,N_2696,N_2733);
nor U2987 (N_2987,N_2759,N_2763);
nor U2988 (N_2988,N_2676,N_2651);
and U2989 (N_2989,N_2791,N_2692);
nand U2990 (N_2990,N_2662,N_2641);
nand U2991 (N_2991,N_2712,N_2768);
nand U2992 (N_2992,N_2689,N_2631);
and U2993 (N_2993,N_2670,N_2781);
nand U2994 (N_2994,N_2647,N_2702);
nor U2995 (N_2995,N_2657,N_2790);
and U2996 (N_2996,N_2604,N_2724);
nand U2997 (N_2997,N_2766,N_2787);
nand U2998 (N_2998,N_2757,N_2667);
and U2999 (N_2999,N_2758,N_2769);
and U3000 (N_3000,N_2993,N_2997);
and U3001 (N_3001,N_2821,N_2905);
and U3002 (N_3002,N_2910,N_2970);
and U3003 (N_3003,N_2991,N_2816);
or U3004 (N_3004,N_2873,N_2926);
and U3005 (N_3005,N_2949,N_2874);
and U3006 (N_3006,N_2865,N_2996);
or U3007 (N_3007,N_2870,N_2899);
and U3008 (N_3008,N_2894,N_2888);
and U3009 (N_3009,N_2866,N_2822);
and U3010 (N_3010,N_2927,N_2988);
and U3011 (N_3011,N_2980,N_2815);
nor U3012 (N_3012,N_2922,N_2952);
or U3013 (N_3013,N_2983,N_2962);
or U3014 (N_3014,N_2919,N_2906);
nand U3015 (N_3015,N_2920,N_2936);
nor U3016 (N_3016,N_2841,N_2937);
and U3017 (N_3017,N_2891,N_2860);
nor U3018 (N_3018,N_2989,N_2976);
nor U3019 (N_3019,N_2979,N_2880);
nor U3020 (N_3020,N_2859,N_2858);
nand U3021 (N_3021,N_2802,N_2824);
nand U3022 (N_3022,N_2887,N_2944);
and U3023 (N_3023,N_2975,N_2820);
or U3024 (N_3024,N_2849,N_2957);
and U3025 (N_3025,N_2961,N_2830);
xor U3026 (N_3026,N_2990,N_2800);
nor U3027 (N_3027,N_2892,N_2958);
or U3028 (N_3028,N_2956,N_2907);
nor U3029 (N_3029,N_2939,N_2898);
nand U3030 (N_3030,N_2984,N_2916);
nor U3031 (N_3031,N_2812,N_2813);
and U3032 (N_3032,N_2987,N_2823);
nand U3033 (N_3033,N_2863,N_2878);
nor U3034 (N_3034,N_2917,N_2965);
or U3035 (N_3035,N_2890,N_2933);
nor U3036 (N_3036,N_2950,N_2992);
and U3037 (N_3037,N_2875,N_2843);
nand U3038 (N_3038,N_2804,N_2911);
and U3039 (N_3039,N_2845,N_2834);
and U3040 (N_3040,N_2872,N_2893);
nor U3041 (N_3041,N_2998,N_2901);
nand U3042 (N_3042,N_2930,N_2896);
and U3043 (N_3043,N_2973,N_2908);
or U3044 (N_3044,N_2831,N_2886);
or U3045 (N_3045,N_2971,N_2972);
or U3046 (N_3046,N_2941,N_2842);
and U3047 (N_3047,N_2904,N_2947);
nand U3048 (N_3048,N_2999,N_2951);
or U3049 (N_3049,N_2844,N_2932);
and U3050 (N_3050,N_2817,N_2814);
and U3051 (N_3051,N_2960,N_2964);
and U3052 (N_3052,N_2895,N_2869);
or U3053 (N_3053,N_2837,N_2913);
nor U3054 (N_3054,N_2914,N_2897);
nand U3055 (N_3055,N_2940,N_2977);
and U3056 (N_3056,N_2885,N_2929);
or U3057 (N_3057,N_2839,N_2828);
or U3058 (N_3058,N_2807,N_2969);
or U3059 (N_3059,N_2889,N_2923);
or U3060 (N_3060,N_2928,N_2803);
and U3061 (N_3061,N_2825,N_2959);
xnor U3062 (N_3062,N_2861,N_2931);
nor U3063 (N_3063,N_2945,N_2850);
and U3064 (N_3064,N_2876,N_2966);
nor U3065 (N_3065,N_2943,N_2856);
or U3066 (N_3066,N_2871,N_2801);
or U3067 (N_3067,N_2827,N_2840);
nand U3068 (N_3068,N_2846,N_2835);
and U3069 (N_3069,N_2852,N_2900);
nand U3070 (N_3070,N_2877,N_2806);
or U3071 (N_3071,N_2909,N_2864);
nand U3072 (N_3072,N_2974,N_2925);
nor U3073 (N_3073,N_2954,N_2838);
nand U3074 (N_3074,N_2882,N_2826);
or U3075 (N_3075,N_2855,N_2982);
or U3076 (N_3076,N_2836,N_2968);
and U3077 (N_3077,N_2854,N_2808);
nand U3078 (N_3078,N_2903,N_2857);
nand U3079 (N_3079,N_2868,N_2986);
nand U3080 (N_3080,N_2833,N_2829);
and U3081 (N_3081,N_2884,N_2811);
nand U3082 (N_3082,N_2819,N_2832);
nand U3083 (N_3083,N_2942,N_2948);
nand U3084 (N_3084,N_2883,N_2809);
or U3085 (N_3085,N_2963,N_2924);
and U3086 (N_3086,N_2953,N_2934);
and U3087 (N_3087,N_2818,N_2967);
nand U3088 (N_3088,N_2915,N_2810);
nor U3089 (N_3089,N_2879,N_2981);
nand U3090 (N_3090,N_2902,N_2918);
nand U3091 (N_3091,N_2935,N_2867);
xor U3092 (N_3092,N_2862,N_2853);
nor U3093 (N_3093,N_2851,N_2847);
and U3094 (N_3094,N_2938,N_2995);
nor U3095 (N_3095,N_2848,N_2912);
and U3096 (N_3096,N_2985,N_2955);
and U3097 (N_3097,N_2921,N_2881);
nor U3098 (N_3098,N_2805,N_2946);
or U3099 (N_3099,N_2994,N_2978);
nor U3100 (N_3100,N_2974,N_2856);
and U3101 (N_3101,N_2875,N_2861);
or U3102 (N_3102,N_2923,N_2932);
and U3103 (N_3103,N_2933,N_2963);
and U3104 (N_3104,N_2996,N_2922);
nor U3105 (N_3105,N_2987,N_2887);
nor U3106 (N_3106,N_2846,N_2945);
nand U3107 (N_3107,N_2841,N_2891);
or U3108 (N_3108,N_2928,N_2930);
and U3109 (N_3109,N_2971,N_2836);
nand U3110 (N_3110,N_2872,N_2839);
and U3111 (N_3111,N_2947,N_2871);
or U3112 (N_3112,N_2858,N_2899);
or U3113 (N_3113,N_2844,N_2858);
and U3114 (N_3114,N_2991,N_2860);
and U3115 (N_3115,N_2844,N_2883);
and U3116 (N_3116,N_2881,N_2832);
or U3117 (N_3117,N_2948,N_2941);
or U3118 (N_3118,N_2919,N_2934);
or U3119 (N_3119,N_2880,N_2976);
or U3120 (N_3120,N_2959,N_2960);
nand U3121 (N_3121,N_2882,N_2901);
or U3122 (N_3122,N_2819,N_2826);
nor U3123 (N_3123,N_2919,N_2911);
and U3124 (N_3124,N_2836,N_2811);
nand U3125 (N_3125,N_2869,N_2817);
and U3126 (N_3126,N_2989,N_2857);
and U3127 (N_3127,N_2820,N_2936);
xor U3128 (N_3128,N_2869,N_2987);
nand U3129 (N_3129,N_2923,N_2822);
and U3130 (N_3130,N_2877,N_2930);
xnor U3131 (N_3131,N_2956,N_2934);
or U3132 (N_3132,N_2840,N_2951);
and U3133 (N_3133,N_2830,N_2827);
and U3134 (N_3134,N_2988,N_2931);
nor U3135 (N_3135,N_2929,N_2965);
nor U3136 (N_3136,N_2819,N_2951);
and U3137 (N_3137,N_2816,N_2994);
nor U3138 (N_3138,N_2882,N_2977);
and U3139 (N_3139,N_2982,N_2956);
nor U3140 (N_3140,N_2816,N_2926);
and U3141 (N_3141,N_2903,N_2802);
xor U3142 (N_3142,N_2954,N_2922);
and U3143 (N_3143,N_2893,N_2930);
or U3144 (N_3144,N_2981,N_2832);
and U3145 (N_3145,N_2885,N_2892);
or U3146 (N_3146,N_2904,N_2892);
nand U3147 (N_3147,N_2984,N_2978);
or U3148 (N_3148,N_2924,N_2903);
nand U3149 (N_3149,N_2893,N_2841);
nand U3150 (N_3150,N_2835,N_2957);
nand U3151 (N_3151,N_2945,N_2936);
nor U3152 (N_3152,N_2872,N_2868);
nor U3153 (N_3153,N_2879,N_2982);
and U3154 (N_3154,N_2885,N_2951);
and U3155 (N_3155,N_2990,N_2918);
nor U3156 (N_3156,N_2920,N_2877);
or U3157 (N_3157,N_2814,N_2970);
and U3158 (N_3158,N_2944,N_2826);
or U3159 (N_3159,N_2864,N_2874);
nand U3160 (N_3160,N_2848,N_2947);
nand U3161 (N_3161,N_2889,N_2898);
or U3162 (N_3162,N_2976,N_2981);
nor U3163 (N_3163,N_2834,N_2868);
and U3164 (N_3164,N_2929,N_2863);
nor U3165 (N_3165,N_2813,N_2860);
nand U3166 (N_3166,N_2882,N_2919);
nor U3167 (N_3167,N_2885,N_2836);
nand U3168 (N_3168,N_2887,N_2945);
or U3169 (N_3169,N_2969,N_2839);
and U3170 (N_3170,N_2944,N_2896);
and U3171 (N_3171,N_2991,N_2864);
nand U3172 (N_3172,N_2906,N_2824);
and U3173 (N_3173,N_2896,N_2823);
or U3174 (N_3174,N_2848,N_2931);
or U3175 (N_3175,N_2843,N_2892);
or U3176 (N_3176,N_2893,N_2912);
nand U3177 (N_3177,N_2857,N_2939);
nor U3178 (N_3178,N_2943,N_2979);
or U3179 (N_3179,N_2805,N_2844);
or U3180 (N_3180,N_2896,N_2838);
or U3181 (N_3181,N_2849,N_2993);
and U3182 (N_3182,N_2886,N_2983);
or U3183 (N_3183,N_2810,N_2934);
and U3184 (N_3184,N_2916,N_2808);
or U3185 (N_3185,N_2801,N_2940);
or U3186 (N_3186,N_2970,N_2876);
nor U3187 (N_3187,N_2913,N_2873);
and U3188 (N_3188,N_2834,N_2953);
nor U3189 (N_3189,N_2850,N_2964);
and U3190 (N_3190,N_2970,N_2864);
and U3191 (N_3191,N_2958,N_2953);
and U3192 (N_3192,N_2962,N_2810);
nor U3193 (N_3193,N_2925,N_2887);
and U3194 (N_3194,N_2984,N_2868);
nor U3195 (N_3195,N_2892,N_2957);
nand U3196 (N_3196,N_2966,N_2945);
and U3197 (N_3197,N_2957,N_2871);
nand U3198 (N_3198,N_2895,N_2850);
and U3199 (N_3199,N_2837,N_2840);
nor U3200 (N_3200,N_3118,N_3195);
nor U3201 (N_3201,N_3169,N_3025);
nor U3202 (N_3202,N_3087,N_3011);
or U3203 (N_3203,N_3142,N_3050);
nor U3204 (N_3204,N_3157,N_3190);
nor U3205 (N_3205,N_3199,N_3045);
nor U3206 (N_3206,N_3089,N_3012);
nand U3207 (N_3207,N_3162,N_3160);
and U3208 (N_3208,N_3174,N_3140);
and U3209 (N_3209,N_3004,N_3153);
and U3210 (N_3210,N_3164,N_3146);
nand U3211 (N_3211,N_3161,N_3110);
nor U3212 (N_3212,N_3056,N_3166);
nor U3213 (N_3213,N_3009,N_3120);
or U3214 (N_3214,N_3141,N_3163);
and U3215 (N_3215,N_3171,N_3096);
nand U3216 (N_3216,N_3090,N_3115);
and U3217 (N_3217,N_3083,N_3073);
and U3218 (N_3218,N_3186,N_3010);
or U3219 (N_3219,N_3181,N_3002);
nor U3220 (N_3220,N_3173,N_3137);
or U3221 (N_3221,N_3032,N_3076);
and U3222 (N_3222,N_3084,N_3194);
nor U3223 (N_3223,N_3058,N_3155);
nand U3224 (N_3224,N_3057,N_3114);
nor U3225 (N_3225,N_3097,N_3072);
nand U3226 (N_3226,N_3189,N_3054);
and U3227 (N_3227,N_3132,N_3091);
nor U3228 (N_3228,N_3128,N_3028);
and U3229 (N_3229,N_3018,N_3124);
nor U3230 (N_3230,N_3106,N_3036);
nor U3231 (N_3231,N_3105,N_3191);
nand U3232 (N_3232,N_3168,N_3078);
nand U3233 (N_3233,N_3134,N_3069);
or U3234 (N_3234,N_3129,N_3098);
and U3235 (N_3235,N_3122,N_3188);
nand U3236 (N_3236,N_3031,N_3013);
nand U3237 (N_3237,N_3187,N_3075);
or U3238 (N_3238,N_3099,N_3037);
nor U3239 (N_3239,N_3059,N_3123);
and U3240 (N_3240,N_3086,N_3030);
or U3241 (N_3241,N_3116,N_3065);
or U3242 (N_3242,N_3111,N_3176);
or U3243 (N_3243,N_3074,N_3143);
and U3244 (N_3244,N_3167,N_3094);
nor U3245 (N_3245,N_3127,N_3048);
and U3246 (N_3246,N_3022,N_3046);
and U3247 (N_3247,N_3023,N_3047);
or U3248 (N_3248,N_3034,N_3055);
and U3249 (N_3249,N_3139,N_3049);
nand U3250 (N_3250,N_3066,N_3039);
and U3251 (N_3251,N_3196,N_3130);
and U3252 (N_3252,N_3197,N_3101);
or U3253 (N_3253,N_3136,N_3107);
nand U3254 (N_3254,N_3158,N_3152);
nand U3255 (N_3255,N_3035,N_3180);
nand U3256 (N_3256,N_3016,N_3100);
nand U3257 (N_3257,N_3193,N_3149);
or U3258 (N_3258,N_3185,N_3170);
and U3259 (N_3259,N_3051,N_3053);
nor U3260 (N_3260,N_3156,N_3020);
nor U3261 (N_3261,N_3005,N_3027);
and U3262 (N_3262,N_3081,N_3000);
nand U3263 (N_3263,N_3088,N_3165);
or U3264 (N_3264,N_3024,N_3178);
and U3265 (N_3265,N_3080,N_3085);
nor U3266 (N_3266,N_3126,N_3183);
and U3267 (N_3267,N_3159,N_3095);
and U3268 (N_3268,N_3042,N_3179);
nand U3269 (N_3269,N_3067,N_3079);
nor U3270 (N_3270,N_3198,N_3135);
xnor U3271 (N_3271,N_3092,N_3104);
and U3272 (N_3272,N_3121,N_3001);
and U3273 (N_3273,N_3082,N_3125);
and U3274 (N_3274,N_3133,N_3147);
nand U3275 (N_3275,N_3117,N_3026);
nand U3276 (N_3276,N_3144,N_3063);
nand U3277 (N_3277,N_3102,N_3151);
nand U3278 (N_3278,N_3040,N_3119);
or U3279 (N_3279,N_3015,N_3052);
and U3280 (N_3280,N_3112,N_3154);
nor U3281 (N_3281,N_3093,N_3060);
and U3282 (N_3282,N_3061,N_3021);
nand U3283 (N_3283,N_3175,N_3014);
or U3284 (N_3284,N_3172,N_3003);
nand U3285 (N_3285,N_3033,N_3044);
or U3286 (N_3286,N_3029,N_3006);
and U3287 (N_3287,N_3109,N_3177);
or U3288 (N_3288,N_3041,N_3077);
nand U3289 (N_3289,N_3103,N_3007);
and U3290 (N_3290,N_3192,N_3070);
nor U3291 (N_3291,N_3148,N_3145);
nor U3292 (N_3292,N_3184,N_3182);
nor U3293 (N_3293,N_3019,N_3071);
nand U3294 (N_3294,N_3038,N_3150);
and U3295 (N_3295,N_3068,N_3131);
and U3296 (N_3296,N_3108,N_3138);
or U3297 (N_3297,N_3064,N_3017);
nand U3298 (N_3298,N_3113,N_3062);
nor U3299 (N_3299,N_3043,N_3008);
and U3300 (N_3300,N_3086,N_3089);
nor U3301 (N_3301,N_3047,N_3115);
xnor U3302 (N_3302,N_3006,N_3163);
nand U3303 (N_3303,N_3167,N_3030);
nand U3304 (N_3304,N_3181,N_3187);
and U3305 (N_3305,N_3198,N_3008);
and U3306 (N_3306,N_3083,N_3123);
or U3307 (N_3307,N_3196,N_3020);
or U3308 (N_3308,N_3163,N_3136);
nand U3309 (N_3309,N_3113,N_3038);
and U3310 (N_3310,N_3083,N_3074);
xor U3311 (N_3311,N_3050,N_3177);
and U3312 (N_3312,N_3035,N_3146);
or U3313 (N_3313,N_3102,N_3135);
and U3314 (N_3314,N_3033,N_3104);
nor U3315 (N_3315,N_3124,N_3082);
nand U3316 (N_3316,N_3188,N_3125);
nor U3317 (N_3317,N_3049,N_3009);
nor U3318 (N_3318,N_3157,N_3031);
nand U3319 (N_3319,N_3032,N_3135);
and U3320 (N_3320,N_3020,N_3039);
nor U3321 (N_3321,N_3166,N_3183);
or U3322 (N_3322,N_3122,N_3116);
nand U3323 (N_3323,N_3142,N_3019);
nand U3324 (N_3324,N_3095,N_3057);
nand U3325 (N_3325,N_3007,N_3068);
or U3326 (N_3326,N_3085,N_3057);
nand U3327 (N_3327,N_3178,N_3095);
nor U3328 (N_3328,N_3106,N_3064);
and U3329 (N_3329,N_3185,N_3190);
and U3330 (N_3330,N_3006,N_3017);
nand U3331 (N_3331,N_3194,N_3105);
or U3332 (N_3332,N_3064,N_3187);
or U3333 (N_3333,N_3008,N_3048);
or U3334 (N_3334,N_3181,N_3158);
or U3335 (N_3335,N_3085,N_3194);
nor U3336 (N_3336,N_3018,N_3134);
and U3337 (N_3337,N_3183,N_3136);
or U3338 (N_3338,N_3119,N_3193);
nand U3339 (N_3339,N_3186,N_3129);
nor U3340 (N_3340,N_3026,N_3145);
or U3341 (N_3341,N_3197,N_3016);
nand U3342 (N_3342,N_3179,N_3005);
or U3343 (N_3343,N_3182,N_3064);
and U3344 (N_3344,N_3003,N_3150);
or U3345 (N_3345,N_3040,N_3130);
nor U3346 (N_3346,N_3120,N_3177);
nor U3347 (N_3347,N_3054,N_3162);
and U3348 (N_3348,N_3002,N_3139);
and U3349 (N_3349,N_3121,N_3088);
or U3350 (N_3350,N_3147,N_3086);
nor U3351 (N_3351,N_3151,N_3032);
nor U3352 (N_3352,N_3170,N_3177);
or U3353 (N_3353,N_3025,N_3037);
nor U3354 (N_3354,N_3045,N_3087);
nand U3355 (N_3355,N_3066,N_3192);
nor U3356 (N_3356,N_3160,N_3001);
nand U3357 (N_3357,N_3135,N_3094);
or U3358 (N_3358,N_3023,N_3121);
and U3359 (N_3359,N_3113,N_3102);
nor U3360 (N_3360,N_3095,N_3119);
or U3361 (N_3361,N_3179,N_3157);
or U3362 (N_3362,N_3103,N_3141);
nor U3363 (N_3363,N_3053,N_3041);
and U3364 (N_3364,N_3051,N_3120);
or U3365 (N_3365,N_3115,N_3123);
or U3366 (N_3366,N_3188,N_3058);
and U3367 (N_3367,N_3133,N_3032);
nand U3368 (N_3368,N_3133,N_3051);
or U3369 (N_3369,N_3189,N_3118);
or U3370 (N_3370,N_3047,N_3108);
nand U3371 (N_3371,N_3149,N_3032);
nor U3372 (N_3372,N_3054,N_3122);
nor U3373 (N_3373,N_3124,N_3156);
nor U3374 (N_3374,N_3046,N_3059);
or U3375 (N_3375,N_3058,N_3052);
nand U3376 (N_3376,N_3064,N_3114);
or U3377 (N_3377,N_3094,N_3159);
and U3378 (N_3378,N_3106,N_3070);
or U3379 (N_3379,N_3103,N_3124);
and U3380 (N_3380,N_3067,N_3104);
nand U3381 (N_3381,N_3124,N_3098);
or U3382 (N_3382,N_3065,N_3037);
nor U3383 (N_3383,N_3179,N_3037);
or U3384 (N_3384,N_3043,N_3071);
and U3385 (N_3385,N_3123,N_3018);
or U3386 (N_3386,N_3124,N_3099);
and U3387 (N_3387,N_3100,N_3063);
nand U3388 (N_3388,N_3141,N_3091);
and U3389 (N_3389,N_3127,N_3178);
or U3390 (N_3390,N_3119,N_3128);
and U3391 (N_3391,N_3101,N_3141);
and U3392 (N_3392,N_3083,N_3128);
or U3393 (N_3393,N_3069,N_3125);
and U3394 (N_3394,N_3148,N_3128);
nor U3395 (N_3395,N_3061,N_3153);
and U3396 (N_3396,N_3057,N_3137);
and U3397 (N_3397,N_3126,N_3042);
and U3398 (N_3398,N_3137,N_3007);
nand U3399 (N_3399,N_3024,N_3119);
nor U3400 (N_3400,N_3278,N_3347);
or U3401 (N_3401,N_3385,N_3271);
nor U3402 (N_3402,N_3374,N_3389);
nor U3403 (N_3403,N_3366,N_3203);
nor U3404 (N_3404,N_3226,N_3341);
nand U3405 (N_3405,N_3279,N_3284);
nand U3406 (N_3406,N_3293,N_3204);
nor U3407 (N_3407,N_3301,N_3322);
and U3408 (N_3408,N_3380,N_3230);
or U3409 (N_3409,N_3299,N_3263);
xnor U3410 (N_3410,N_3249,N_3220);
or U3411 (N_3411,N_3340,N_3291);
nand U3412 (N_3412,N_3210,N_3397);
or U3413 (N_3413,N_3202,N_3298);
nor U3414 (N_3414,N_3376,N_3304);
or U3415 (N_3415,N_3213,N_3394);
or U3416 (N_3416,N_3307,N_3209);
nor U3417 (N_3417,N_3267,N_3367);
nor U3418 (N_3418,N_3318,N_3212);
nand U3419 (N_3419,N_3262,N_3388);
and U3420 (N_3420,N_3349,N_3223);
nand U3421 (N_3421,N_3297,N_3275);
nand U3422 (N_3422,N_3254,N_3343);
and U3423 (N_3423,N_3221,N_3260);
nand U3424 (N_3424,N_3342,N_3378);
nor U3425 (N_3425,N_3237,N_3206);
nor U3426 (N_3426,N_3396,N_3384);
nor U3427 (N_3427,N_3353,N_3264);
or U3428 (N_3428,N_3294,N_3258);
nor U3429 (N_3429,N_3346,N_3375);
and U3430 (N_3430,N_3348,N_3320);
or U3431 (N_3431,N_3269,N_3361);
or U3432 (N_3432,N_3280,N_3246);
nand U3433 (N_3433,N_3368,N_3216);
nand U3434 (N_3434,N_3395,N_3285);
and U3435 (N_3435,N_3235,N_3336);
and U3436 (N_3436,N_3356,N_3329);
nor U3437 (N_3437,N_3363,N_3339);
and U3438 (N_3438,N_3370,N_3288);
nor U3439 (N_3439,N_3219,N_3265);
nor U3440 (N_3440,N_3313,N_3252);
nor U3441 (N_3441,N_3350,N_3282);
and U3442 (N_3442,N_3359,N_3222);
and U3443 (N_3443,N_3326,N_3247);
and U3444 (N_3444,N_3305,N_3218);
nand U3445 (N_3445,N_3323,N_3399);
nor U3446 (N_3446,N_3351,N_3215);
and U3447 (N_3447,N_3241,N_3227);
nor U3448 (N_3448,N_3332,N_3200);
nor U3449 (N_3449,N_3311,N_3393);
and U3450 (N_3450,N_3392,N_3387);
nor U3451 (N_3451,N_3268,N_3352);
nor U3452 (N_3452,N_3334,N_3214);
or U3453 (N_3453,N_3328,N_3270);
xor U3454 (N_3454,N_3261,N_3205);
nand U3455 (N_3455,N_3309,N_3242);
nand U3456 (N_3456,N_3228,N_3371);
and U3457 (N_3457,N_3354,N_3233);
or U3458 (N_3458,N_3379,N_3358);
nor U3459 (N_3459,N_3208,N_3245);
nand U3460 (N_3460,N_3300,N_3273);
nand U3461 (N_3461,N_3259,N_3272);
nand U3462 (N_3462,N_3372,N_3256);
nand U3463 (N_3463,N_3250,N_3327);
nor U3464 (N_3464,N_3362,N_3224);
nand U3465 (N_3465,N_3308,N_3355);
nor U3466 (N_3466,N_3234,N_3357);
and U3467 (N_3467,N_3287,N_3330);
or U3468 (N_3468,N_3211,N_3286);
or U3469 (N_3469,N_3325,N_3248);
xor U3470 (N_3470,N_3333,N_3290);
or U3471 (N_3471,N_3314,N_3255);
and U3472 (N_3472,N_3251,N_3281);
nor U3473 (N_3473,N_3289,N_3383);
and U3474 (N_3474,N_3386,N_3344);
nor U3475 (N_3475,N_3390,N_3319);
and U3476 (N_3476,N_3303,N_3257);
or U3477 (N_3477,N_3243,N_3381);
nand U3478 (N_3478,N_3398,N_3312);
or U3479 (N_3479,N_3377,N_3232);
nor U3480 (N_3480,N_3266,N_3217);
nand U3481 (N_3481,N_3292,N_3317);
nand U3482 (N_3482,N_3316,N_3239);
nand U3483 (N_3483,N_3201,N_3240);
or U3484 (N_3484,N_3306,N_3229);
and U3485 (N_3485,N_3382,N_3338);
nand U3486 (N_3486,N_3345,N_3296);
and U3487 (N_3487,N_3364,N_3225);
nor U3488 (N_3488,N_3276,N_3324);
or U3489 (N_3489,N_3277,N_3373);
and U3490 (N_3490,N_3369,N_3321);
and U3491 (N_3491,N_3231,N_3315);
and U3492 (N_3492,N_3302,N_3253);
and U3493 (N_3493,N_3391,N_3274);
nor U3494 (N_3494,N_3337,N_3360);
nand U3495 (N_3495,N_3207,N_3244);
nor U3496 (N_3496,N_3238,N_3310);
nor U3497 (N_3497,N_3331,N_3283);
and U3498 (N_3498,N_3236,N_3365);
or U3499 (N_3499,N_3335,N_3295);
nand U3500 (N_3500,N_3225,N_3360);
and U3501 (N_3501,N_3342,N_3392);
and U3502 (N_3502,N_3352,N_3279);
nor U3503 (N_3503,N_3307,N_3214);
or U3504 (N_3504,N_3249,N_3313);
nand U3505 (N_3505,N_3232,N_3389);
or U3506 (N_3506,N_3395,N_3224);
nor U3507 (N_3507,N_3245,N_3343);
nor U3508 (N_3508,N_3284,N_3344);
nand U3509 (N_3509,N_3355,N_3353);
or U3510 (N_3510,N_3233,N_3243);
and U3511 (N_3511,N_3379,N_3205);
or U3512 (N_3512,N_3297,N_3268);
nand U3513 (N_3513,N_3357,N_3264);
or U3514 (N_3514,N_3218,N_3352);
nor U3515 (N_3515,N_3277,N_3379);
or U3516 (N_3516,N_3264,N_3220);
nand U3517 (N_3517,N_3350,N_3370);
or U3518 (N_3518,N_3247,N_3238);
nor U3519 (N_3519,N_3347,N_3396);
and U3520 (N_3520,N_3367,N_3208);
nand U3521 (N_3521,N_3206,N_3212);
nor U3522 (N_3522,N_3319,N_3316);
and U3523 (N_3523,N_3227,N_3259);
or U3524 (N_3524,N_3246,N_3277);
or U3525 (N_3525,N_3399,N_3317);
nor U3526 (N_3526,N_3228,N_3351);
and U3527 (N_3527,N_3379,N_3382);
nand U3528 (N_3528,N_3264,N_3356);
xnor U3529 (N_3529,N_3345,N_3321);
nand U3530 (N_3530,N_3230,N_3335);
and U3531 (N_3531,N_3389,N_3342);
and U3532 (N_3532,N_3243,N_3366);
and U3533 (N_3533,N_3320,N_3303);
and U3534 (N_3534,N_3257,N_3307);
or U3535 (N_3535,N_3229,N_3232);
nand U3536 (N_3536,N_3361,N_3355);
nand U3537 (N_3537,N_3300,N_3375);
nor U3538 (N_3538,N_3252,N_3342);
and U3539 (N_3539,N_3211,N_3365);
nor U3540 (N_3540,N_3368,N_3330);
and U3541 (N_3541,N_3234,N_3381);
nand U3542 (N_3542,N_3206,N_3326);
nor U3543 (N_3543,N_3364,N_3307);
nor U3544 (N_3544,N_3371,N_3230);
nand U3545 (N_3545,N_3261,N_3378);
and U3546 (N_3546,N_3244,N_3209);
or U3547 (N_3547,N_3255,N_3246);
nand U3548 (N_3548,N_3372,N_3222);
and U3549 (N_3549,N_3236,N_3262);
nor U3550 (N_3550,N_3282,N_3214);
or U3551 (N_3551,N_3210,N_3231);
or U3552 (N_3552,N_3230,N_3363);
or U3553 (N_3553,N_3377,N_3268);
nor U3554 (N_3554,N_3338,N_3240);
or U3555 (N_3555,N_3272,N_3356);
and U3556 (N_3556,N_3233,N_3388);
and U3557 (N_3557,N_3279,N_3239);
or U3558 (N_3558,N_3269,N_3386);
nor U3559 (N_3559,N_3298,N_3256);
and U3560 (N_3560,N_3363,N_3300);
nand U3561 (N_3561,N_3287,N_3315);
or U3562 (N_3562,N_3207,N_3350);
or U3563 (N_3563,N_3351,N_3226);
nor U3564 (N_3564,N_3286,N_3304);
or U3565 (N_3565,N_3359,N_3389);
or U3566 (N_3566,N_3208,N_3271);
or U3567 (N_3567,N_3231,N_3246);
and U3568 (N_3568,N_3381,N_3343);
and U3569 (N_3569,N_3242,N_3270);
and U3570 (N_3570,N_3348,N_3350);
nand U3571 (N_3571,N_3254,N_3212);
or U3572 (N_3572,N_3375,N_3285);
or U3573 (N_3573,N_3323,N_3358);
or U3574 (N_3574,N_3386,N_3222);
nand U3575 (N_3575,N_3322,N_3290);
and U3576 (N_3576,N_3312,N_3233);
or U3577 (N_3577,N_3285,N_3259);
nor U3578 (N_3578,N_3270,N_3367);
or U3579 (N_3579,N_3225,N_3216);
or U3580 (N_3580,N_3362,N_3285);
or U3581 (N_3581,N_3302,N_3274);
or U3582 (N_3582,N_3303,N_3326);
and U3583 (N_3583,N_3393,N_3228);
nand U3584 (N_3584,N_3394,N_3285);
nand U3585 (N_3585,N_3380,N_3309);
nor U3586 (N_3586,N_3368,N_3370);
nand U3587 (N_3587,N_3249,N_3239);
or U3588 (N_3588,N_3273,N_3242);
nor U3589 (N_3589,N_3286,N_3244);
nor U3590 (N_3590,N_3269,N_3374);
or U3591 (N_3591,N_3285,N_3258);
nand U3592 (N_3592,N_3345,N_3357);
nor U3593 (N_3593,N_3367,N_3339);
or U3594 (N_3594,N_3302,N_3310);
or U3595 (N_3595,N_3216,N_3239);
and U3596 (N_3596,N_3254,N_3204);
and U3597 (N_3597,N_3290,N_3382);
nor U3598 (N_3598,N_3289,N_3218);
nand U3599 (N_3599,N_3369,N_3382);
and U3600 (N_3600,N_3537,N_3532);
or U3601 (N_3601,N_3566,N_3491);
and U3602 (N_3602,N_3590,N_3443);
nor U3603 (N_3603,N_3548,N_3448);
nand U3604 (N_3604,N_3488,N_3553);
and U3605 (N_3605,N_3433,N_3504);
nand U3606 (N_3606,N_3586,N_3564);
or U3607 (N_3607,N_3415,N_3527);
nor U3608 (N_3608,N_3544,N_3525);
nor U3609 (N_3609,N_3464,N_3571);
and U3610 (N_3610,N_3402,N_3475);
nand U3611 (N_3611,N_3518,N_3509);
nand U3612 (N_3612,N_3462,N_3523);
and U3613 (N_3613,N_3472,N_3536);
or U3614 (N_3614,N_3439,N_3461);
nor U3615 (N_3615,N_3493,N_3558);
nor U3616 (N_3616,N_3511,N_3519);
or U3617 (N_3617,N_3458,N_3570);
nand U3618 (N_3618,N_3434,N_3427);
and U3619 (N_3619,N_3568,N_3520);
and U3620 (N_3620,N_3560,N_3411);
or U3621 (N_3621,N_3428,N_3572);
nand U3622 (N_3622,N_3487,N_3403);
xnor U3623 (N_3623,N_3492,N_3440);
and U3624 (N_3624,N_3417,N_3438);
nor U3625 (N_3625,N_3524,N_3517);
nand U3626 (N_3626,N_3486,N_3593);
nor U3627 (N_3627,N_3540,N_3578);
nand U3628 (N_3628,N_3460,N_3468);
and U3629 (N_3629,N_3576,N_3422);
or U3630 (N_3630,N_3421,N_3592);
nor U3631 (N_3631,N_3408,N_3552);
or U3632 (N_3632,N_3406,N_3583);
nand U3633 (N_3633,N_3501,N_3424);
or U3634 (N_3634,N_3581,N_3471);
nor U3635 (N_3635,N_3477,N_3530);
nor U3636 (N_3636,N_3426,N_3413);
nand U3637 (N_3637,N_3549,N_3529);
or U3638 (N_3638,N_3589,N_3480);
and U3639 (N_3639,N_3494,N_3412);
nor U3640 (N_3640,N_3534,N_3561);
nor U3641 (N_3641,N_3555,N_3508);
nor U3642 (N_3642,N_3441,N_3409);
nor U3643 (N_3643,N_3510,N_3484);
nor U3644 (N_3644,N_3542,N_3446);
and U3645 (N_3645,N_3505,N_3502);
nand U3646 (N_3646,N_3584,N_3551);
and U3647 (N_3647,N_3420,N_3506);
nor U3648 (N_3648,N_3541,N_3514);
nand U3649 (N_3649,N_3459,N_3585);
nand U3650 (N_3650,N_3538,N_3528);
nor U3651 (N_3651,N_3598,N_3591);
nand U3652 (N_3652,N_3436,N_3457);
nand U3653 (N_3653,N_3483,N_3513);
nor U3654 (N_3654,N_3485,N_3476);
nand U3655 (N_3655,N_3445,N_3473);
nor U3656 (N_3656,N_3414,N_3425);
nor U3657 (N_3657,N_3495,N_3451);
and U3658 (N_3658,N_3569,N_3437);
and U3659 (N_3659,N_3533,N_3587);
and U3660 (N_3660,N_3582,N_3594);
or U3661 (N_3661,N_3467,N_3503);
or U3662 (N_3662,N_3547,N_3469);
xor U3663 (N_3663,N_3565,N_3481);
nand U3664 (N_3664,N_3507,N_3429);
nand U3665 (N_3665,N_3497,N_3496);
and U3666 (N_3666,N_3521,N_3482);
and U3667 (N_3667,N_3450,N_3512);
and U3668 (N_3668,N_3423,N_3595);
or U3669 (N_3669,N_3410,N_3562);
or U3670 (N_3670,N_3474,N_3404);
nor U3671 (N_3671,N_3452,N_3522);
nand U3672 (N_3672,N_3557,N_3577);
nand U3673 (N_3673,N_3454,N_3545);
and U3674 (N_3674,N_3400,N_3419);
and U3675 (N_3675,N_3574,N_3432);
and U3676 (N_3676,N_3435,N_3588);
and U3677 (N_3677,N_3418,N_3563);
nand U3678 (N_3678,N_3431,N_3596);
nand U3679 (N_3679,N_3456,N_3556);
nor U3680 (N_3680,N_3554,N_3559);
nor U3681 (N_3681,N_3453,N_3416);
xor U3682 (N_3682,N_3573,N_3535);
nand U3683 (N_3683,N_3500,N_3567);
nor U3684 (N_3684,N_3599,N_3550);
nor U3685 (N_3685,N_3546,N_3489);
nand U3686 (N_3686,N_3490,N_3444);
and U3687 (N_3687,N_3442,N_3515);
or U3688 (N_3688,N_3580,N_3516);
nor U3689 (N_3689,N_3526,N_3405);
nor U3690 (N_3690,N_3531,N_3401);
and U3691 (N_3691,N_3449,N_3597);
nand U3692 (N_3692,N_3407,N_3478);
xnor U3693 (N_3693,N_3463,N_3539);
or U3694 (N_3694,N_3498,N_3466);
xnor U3695 (N_3695,N_3479,N_3579);
or U3696 (N_3696,N_3430,N_3575);
nor U3697 (N_3697,N_3455,N_3447);
or U3698 (N_3698,N_3465,N_3499);
and U3699 (N_3699,N_3470,N_3543);
nand U3700 (N_3700,N_3574,N_3516);
or U3701 (N_3701,N_3588,N_3404);
and U3702 (N_3702,N_3468,N_3408);
or U3703 (N_3703,N_3505,N_3581);
or U3704 (N_3704,N_3561,N_3466);
nor U3705 (N_3705,N_3589,N_3581);
and U3706 (N_3706,N_3479,N_3444);
and U3707 (N_3707,N_3590,N_3579);
nor U3708 (N_3708,N_3411,N_3507);
or U3709 (N_3709,N_3415,N_3463);
nand U3710 (N_3710,N_3519,N_3476);
nand U3711 (N_3711,N_3491,N_3508);
nand U3712 (N_3712,N_3593,N_3445);
nand U3713 (N_3713,N_3480,N_3538);
nand U3714 (N_3714,N_3416,N_3430);
nand U3715 (N_3715,N_3439,N_3585);
and U3716 (N_3716,N_3437,N_3425);
nor U3717 (N_3717,N_3539,N_3536);
nand U3718 (N_3718,N_3420,N_3594);
nor U3719 (N_3719,N_3543,N_3480);
or U3720 (N_3720,N_3468,N_3509);
nand U3721 (N_3721,N_3519,N_3403);
and U3722 (N_3722,N_3589,N_3563);
or U3723 (N_3723,N_3560,N_3518);
and U3724 (N_3724,N_3505,N_3454);
nand U3725 (N_3725,N_3511,N_3427);
nor U3726 (N_3726,N_3549,N_3438);
nor U3727 (N_3727,N_3425,N_3511);
nor U3728 (N_3728,N_3508,N_3556);
and U3729 (N_3729,N_3566,N_3436);
and U3730 (N_3730,N_3497,N_3546);
and U3731 (N_3731,N_3502,N_3522);
nor U3732 (N_3732,N_3415,N_3405);
nand U3733 (N_3733,N_3485,N_3572);
or U3734 (N_3734,N_3472,N_3476);
or U3735 (N_3735,N_3480,N_3479);
xnor U3736 (N_3736,N_3493,N_3518);
or U3737 (N_3737,N_3472,N_3466);
or U3738 (N_3738,N_3569,N_3401);
nor U3739 (N_3739,N_3439,N_3491);
nand U3740 (N_3740,N_3426,N_3425);
nor U3741 (N_3741,N_3437,N_3440);
nor U3742 (N_3742,N_3492,N_3457);
or U3743 (N_3743,N_3499,N_3537);
nand U3744 (N_3744,N_3585,N_3443);
or U3745 (N_3745,N_3575,N_3496);
nand U3746 (N_3746,N_3567,N_3566);
or U3747 (N_3747,N_3444,N_3437);
and U3748 (N_3748,N_3479,N_3445);
xnor U3749 (N_3749,N_3540,N_3552);
or U3750 (N_3750,N_3565,N_3524);
or U3751 (N_3751,N_3512,N_3582);
nor U3752 (N_3752,N_3493,N_3409);
nor U3753 (N_3753,N_3583,N_3501);
and U3754 (N_3754,N_3453,N_3408);
and U3755 (N_3755,N_3453,N_3518);
or U3756 (N_3756,N_3446,N_3423);
nand U3757 (N_3757,N_3430,N_3497);
nor U3758 (N_3758,N_3427,N_3571);
or U3759 (N_3759,N_3412,N_3587);
and U3760 (N_3760,N_3557,N_3473);
nor U3761 (N_3761,N_3486,N_3524);
nor U3762 (N_3762,N_3428,N_3546);
nor U3763 (N_3763,N_3561,N_3468);
or U3764 (N_3764,N_3510,N_3576);
nor U3765 (N_3765,N_3437,N_3561);
and U3766 (N_3766,N_3578,N_3546);
or U3767 (N_3767,N_3553,N_3554);
nand U3768 (N_3768,N_3595,N_3454);
nor U3769 (N_3769,N_3536,N_3503);
or U3770 (N_3770,N_3564,N_3502);
nor U3771 (N_3771,N_3498,N_3533);
and U3772 (N_3772,N_3476,N_3572);
nor U3773 (N_3773,N_3580,N_3586);
nor U3774 (N_3774,N_3515,N_3474);
and U3775 (N_3775,N_3440,N_3444);
nand U3776 (N_3776,N_3528,N_3516);
nor U3777 (N_3777,N_3440,N_3472);
and U3778 (N_3778,N_3406,N_3585);
nor U3779 (N_3779,N_3488,N_3484);
and U3780 (N_3780,N_3534,N_3577);
nor U3781 (N_3781,N_3470,N_3404);
nor U3782 (N_3782,N_3530,N_3478);
or U3783 (N_3783,N_3501,N_3564);
and U3784 (N_3784,N_3558,N_3528);
nor U3785 (N_3785,N_3532,N_3418);
nor U3786 (N_3786,N_3505,N_3442);
and U3787 (N_3787,N_3572,N_3488);
nor U3788 (N_3788,N_3400,N_3505);
nor U3789 (N_3789,N_3544,N_3412);
or U3790 (N_3790,N_3476,N_3479);
and U3791 (N_3791,N_3452,N_3447);
nand U3792 (N_3792,N_3496,N_3523);
nor U3793 (N_3793,N_3437,N_3465);
or U3794 (N_3794,N_3520,N_3592);
nor U3795 (N_3795,N_3597,N_3539);
and U3796 (N_3796,N_3445,N_3512);
nor U3797 (N_3797,N_3496,N_3475);
nand U3798 (N_3798,N_3582,N_3518);
and U3799 (N_3799,N_3413,N_3558);
nor U3800 (N_3800,N_3632,N_3746);
and U3801 (N_3801,N_3784,N_3645);
nor U3802 (N_3802,N_3748,N_3676);
nand U3803 (N_3803,N_3761,N_3720);
or U3804 (N_3804,N_3765,N_3622);
nand U3805 (N_3805,N_3663,N_3618);
and U3806 (N_3806,N_3722,N_3753);
nor U3807 (N_3807,N_3728,N_3772);
or U3808 (N_3808,N_3656,N_3675);
nand U3809 (N_3809,N_3613,N_3710);
nand U3810 (N_3810,N_3709,N_3660);
nor U3811 (N_3811,N_3705,N_3665);
and U3812 (N_3812,N_3624,N_3747);
nand U3813 (N_3813,N_3732,N_3643);
or U3814 (N_3814,N_3766,N_3630);
nand U3815 (N_3815,N_3777,N_3771);
nor U3816 (N_3816,N_3605,N_3652);
nor U3817 (N_3817,N_3634,N_3730);
or U3818 (N_3818,N_3641,N_3607);
nand U3819 (N_3819,N_3686,N_3773);
nor U3820 (N_3820,N_3754,N_3714);
and U3821 (N_3821,N_3608,N_3621);
or U3822 (N_3822,N_3694,N_3731);
and U3823 (N_3823,N_3651,N_3729);
or U3824 (N_3824,N_3733,N_3637);
or U3825 (N_3825,N_3623,N_3774);
or U3826 (N_3826,N_3795,N_3738);
or U3827 (N_3827,N_3685,N_3752);
or U3828 (N_3828,N_3734,N_3798);
nor U3829 (N_3829,N_3750,N_3677);
nor U3830 (N_3830,N_3679,N_3668);
xnor U3831 (N_3831,N_3716,N_3727);
and U3832 (N_3832,N_3781,N_3755);
nand U3833 (N_3833,N_3620,N_3741);
or U3834 (N_3834,N_3690,N_3662);
or U3835 (N_3835,N_3604,N_3718);
nor U3836 (N_3836,N_3642,N_3737);
nand U3837 (N_3837,N_3786,N_3695);
nand U3838 (N_3838,N_3708,N_3661);
or U3839 (N_3839,N_3745,N_3776);
and U3840 (N_3840,N_3769,N_3768);
and U3841 (N_3841,N_3625,N_3666);
nor U3842 (N_3842,N_3759,N_3749);
or U3843 (N_3843,N_3650,N_3764);
nor U3844 (N_3844,N_3706,N_3793);
and U3845 (N_3845,N_3606,N_3635);
and U3846 (N_3846,N_3636,N_3610);
nor U3847 (N_3847,N_3797,N_3667);
nor U3848 (N_3848,N_3671,N_3654);
and U3849 (N_3849,N_3788,N_3659);
and U3850 (N_3850,N_3664,N_3683);
or U3851 (N_3851,N_3633,N_3682);
and U3852 (N_3852,N_3611,N_3684);
and U3853 (N_3853,N_3619,N_3770);
nand U3854 (N_3854,N_3719,N_3669);
nor U3855 (N_3855,N_3726,N_3778);
or U3856 (N_3856,N_3790,N_3672);
nor U3857 (N_3857,N_3744,N_3615);
or U3858 (N_3858,N_3712,N_3715);
nand U3859 (N_3859,N_3796,N_3678);
nor U3860 (N_3860,N_3758,N_3688);
or U3861 (N_3861,N_3600,N_3603);
nor U3862 (N_3862,N_3681,N_3696);
and U3863 (N_3863,N_3711,N_3789);
nor U3864 (N_3864,N_3780,N_3783);
or U3865 (N_3865,N_3742,N_3787);
and U3866 (N_3866,N_3717,N_3743);
and U3867 (N_3867,N_3617,N_3767);
and U3868 (N_3868,N_3779,N_3639);
and U3869 (N_3869,N_3601,N_3724);
nand U3870 (N_3870,N_3616,N_3785);
nor U3871 (N_3871,N_3707,N_3699);
nor U3872 (N_3872,N_3721,N_3691);
nand U3873 (N_3873,N_3629,N_3698);
and U3874 (N_3874,N_3704,N_3674);
nand U3875 (N_3875,N_3692,N_3614);
or U3876 (N_3876,N_3653,N_3792);
nor U3877 (N_3877,N_3702,N_3757);
nor U3878 (N_3878,N_3638,N_3736);
nand U3879 (N_3879,N_3739,N_3644);
or U3880 (N_3880,N_3701,N_3646);
and U3881 (N_3881,N_3751,N_3612);
and U3882 (N_3882,N_3703,N_3723);
nand U3883 (N_3883,N_3657,N_3647);
or U3884 (N_3884,N_3680,N_3756);
or U3885 (N_3885,N_3640,N_3689);
xor U3886 (N_3886,N_3740,N_3628);
nor U3887 (N_3887,N_3693,N_3775);
and U3888 (N_3888,N_3700,N_3794);
or U3889 (N_3889,N_3627,N_3609);
nand U3890 (N_3890,N_3687,N_3782);
or U3891 (N_3891,N_3649,N_3648);
and U3892 (N_3892,N_3602,N_3658);
and U3893 (N_3893,N_3631,N_3670);
or U3894 (N_3894,N_3735,N_3725);
nor U3895 (N_3895,N_3799,N_3673);
and U3896 (N_3896,N_3655,N_3626);
or U3897 (N_3897,N_3762,N_3791);
nor U3898 (N_3898,N_3713,N_3760);
nand U3899 (N_3899,N_3763,N_3697);
and U3900 (N_3900,N_3755,N_3673);
nor U3901 (N_3901,N_3676,N_3774);
nand U3902 (N_3902,N_3666,N_3752);
nand U3903 (N_3903,N_3652,N_3701);
nand U3904 (N_3904,N_3727,N_3624);
or U3905 (N_3905,N_3783,N_3784);
nor U3906 (N_3906,N_3759,N_3618);
and U3907 (N_3907,N_3605,N_3790);
nor U3908 (N_3908,N_3662,N_3724);
nand U3909 (N_3909,N_3710,N_3693);
nand U3910 (N_3910,N_3621,N_3677);
xnor U3911 (N_3911,N_3718,N_3662);
nand U3912 (N_3912,N_3701,N_3712);
nor U3913 (N_3913,N_3788,N_3729);
or U3914 (N_3914,N_3738,N_3763);
nor U3915 (N_3915,N_3712,N_3772);
and U3916 (N_3916,N_3755,N_3658);
nor U3917 (N_3917,N_3601,N_3705);
and U3918 (N_3918,N_3603,N_3777);
nand U3919 (N_3919,N_3686,N_3622);
nand U3920 (N_3920,N_3693,N_3621);
nand U3921 (N_3921,N_3796,N_3790);
nor U3922 (N_3922,N_3722,N_3631);
and U3923 (N_3923,N_3693,N_3726);
nor U3924 (N_3924,N_3723,N_3739);
nand U3925 (N_3925,N_3618,N_3603);
or U3926 (N_3926,N_3605,N_3686);
nor U3927 (N_3927,N_3648,N_3698);
nor U3928 (N_3928,N_3618,N_3686);
nor U3929 (N_3929,N_3610,N_3624);
or U3930 (N_3930,N_3748,N_3604);
nor U3931 (N_3931,N_3755,N_3715);
nand U3932 (N_3932,N_3615,N_3605);
and U3933 (N_3933,N_3759,N_3789);
nor U3934 (N_3934,N_3652,N_3753);
nand U3935 (N_3935,N_3662,N_3657);
nor U3936 (N_3936,N_3786,N_3626);
nand U3937 (N_3937,N_3637,N_3670);
nor U3938 (N_3938,N_3728,N_3600);
nor U3939 (N_3939,N_3722,N_3776);
and U3940 (N_3940,N_3649,N_3797);
nand U3941 (N_3941,N_3734,N_3706);
and U3942 (N_3942,N_3671,N_3753);
and U3943 (N_3943,N_3723,N_3701);
nor U3944 (N_3944,N_3744,N_3698);
nor U3945 (N_3945,N_3727,N_3600);
and U3946 (N_3946,N_3729,N_3649);
nor U3947 (N_3947,N_3693,N_3774);
nand U3948 (N_3948,N_3644,N_3758);
nand U3949 (N_3949,N_3760,N_3662);
and U3950 (N_3950,N_3759,N_3651);
or U3951 (N_3951,N_3780,N_3747);
xor U3952 (N_3952,N_3628,N_3633);
nand U3953 (N_3953,N_3685,N_3759);
nand U3954 (N_3954,N_3675,N_3652);
nor U3955 (N_3955,N_3785,N_3609);
or U3956 (N_3956,N_3774,N_3609);
and U3957 (N_3957,N_3794,N_3725);
nand U3958 (N_3958,N_3605,N_3704);
and U3959 (N_3959,N_3766,N_3683);
xnor U3960 (N_3960,N_3601,N_3667);
or U3961 (N_3961,N_3777,N_3745);
nand U3962 (N_3962,N_3609,N_3710);
nor U3963 (N_3963,N_3731,N_3758);
or U3964 (N_3964,N_3714,N_3639);
and U3965 (N_3965,N_3625,N_3741);
nor U3966 (N_3966,N_3776,N_3779);
nor U3967 (N_3967,N_3700,N_3699);
or U3968 (N_3968,N_3604,N_3712);
and U3969 (N_3969,N_3638,N_3786);
and U3970 (N_3970,N_3606,N_3600);
or U3971 (N_3971,N_3795,N_3660);
or U3972 (N_3972,N_3792,N_3685);
and U3973 (N_3973,N_3799,N_3633);
nor U3974 (N_3974,N_3770,N_3604);
nor U3975 (N_3975,N_3796,N_3747);
or U3976 (N_3976,N_3640,N_3665);
nor U3977 (N_3977,N_3777,N_3710);
and U3978 (N_3978,N_3621,N_3612);
nand U3979 (N_3979,N_3731,N_3653);
or U3980 (N_3980,N_3675,N_3799);
nand U3981 (N_3981,N_3661,N_3600);
and U3982 (N_3982,N_3742,N_3775);
nand U3983 (N_3983,N_3702,N_3644);
or U3984 (N_3984,N_3731,N_3771);
and U3985 (N_3985,N_3615,N_3643);
nor U3986 (N_3986,N_3621,N_3620);
or U3987 (N_3987,N_3799,N_3674);
nor U3988 (N_3988,N_3706,N_3662);
nor U3989 (N_3989,N_3678,N_3615);
and U3990 (N_3990,N_3678,N_3741);
nand U3991 (N_3991,N_3728,N_3670);
or U3992 (N_3992,N_3655,N_3633);
and U3993 (N_3993,N_3661,N_3745);
nand U3994 (N_3994,N_3689,N_3747);
and U3995 (N_3995,N_3605,N_3725);
nand U3996 (N_3996,N_3600,N_3651);
nand U3997 (N_3997,N_3647,N_3655);
and U3998 (N_3998,N_3644,N_3657);
and U3999 (N_3999,N_3666,N_3687);
nor U4000 (N_4000,N_3822,N_3945);
or U4001 (N_4001,N_3830,N_3898);
nand U4002 (N_4002,N_3856,N_3821);
and U4003 (N_4003,N_3979,N_3932);
nor U4004 (N_4004,N_3926,N_3812);
nor U4005 (N_4005,N_3904,N_3927);
or U4006 (N_4006,N_3862,N_3987);
and U4007 (N_4007,N_3910,N_3915);
nor U4008 (N_4008,N_3917,N_3866);
nor U4009 (N_4009,N_3903,N_3848);
nand U4010 (N_4010,N_3850,N_3899);
or U4011 (N_4011,N_3936,N_3867);
xor U4012 (N_4012,N_3890,N_3801);
and U4013 (N_4013,N_3986,N_3819);
nand U4014 (N_4014,N_3929,N_3994);
or U4015 (N_4015,N_3884,N_3880);
nand U4016 (N_4016,N_3914,N_3882);
and U4017 (N_4017,N_3988,N_3836);
and U4018 (N_4018,N_3922,N_3804);
nor U4019 (N_4019,N_3909,N_3990);
nand U4020 (N_4020,N_3959,N_3870);
or U4021 (N_4021,N_3983,N_3920);
xnor U4022 (N_4022,N_3855,N_3806);
or U4023 (N_4023,N_3967,N_3846);
and U4024 (N_4024,N_3813,N_3940);
and U4025 (N_4025,N_3934,N_3900);
or U4026 (N_4026,N_3951,N_3859);
and U4027 (N_4027,N_3879,N_3984);
nand U4028 (N_4028,N_3919,N_3863);
nor U4029 (N_4029,N_3905,N_3825);
and U4030 (N_4030,N_3996,N_3956);
xor U4031 (N_4031,N_3944,N_3807);
or U4032 (N_4032,N_3977,N_3968);
and U4033 (N_4033,N_3949,N_3823);
nand U4034 (N_4034,N_3876,N_3955);
or U4035 (N_4035,N_3965,N_3924);
or U4036 (N_4036,N_3815,N_3889);
nand U4037 (N_4037,N_3962,N_3958);
and U4038 (N_4038,N_3947,N_3916);
and U4039 (N_4039,N_3891,N_3963);
and U4040 (N_4040,N_3989,N_3953);
nor U4041 (N_4041,N_3998,N_3871);
nor U4042 (N_4042,N_3906,N_3901);
and U4043 (N_4043,N_3839,N_3893);
nand U4044 (N_4044,N_3969,N_3831);
nand U4045 (N_4045,N_3948,N_3816);
or U4046 (N_4046,N_3974,N_3992);
nand U4047 (N_4047,N_3985,N_3809);
nand U4048 (N_4048,N_3802,N_3824);
or U4049 (N_4049,N_3837,N_3960);
or U4050 (N_4050,N_3918,N_3851);
or U4051 (N_4051,N_3852,N_3838);
nor U4052 (N_4052,N_3896,N_3857);
nand U4053 (N_4053,N_3853,N_3895);
or U4054 (N_4054,N_3980,N_3843);
nor U4055 (N_4055,N_3858,N_3943);
xnor U4056 (N_4056,N_3975,N_3805);
and U4057 (N_4057,N_3817,N_3973);
and U4058 (N_4058,N_3810,N_3892);
nand U4059 (N_4059,N_3912,N_3972);
nand U4060 (N_4060,N_3885,N_3941);
nand U4061 (N_4061,N_3829,N_3952);
and U4062 (N_4062,N_3849,N_3868);
or U4063 (N_4063,N_3921,N_3913);
and U4064 (N_4064,N_3835,N_3847);
nand U4065 (N_4065,N_3946,N_3957);
or U4066 (N_4066,N_3902,N_3911);
or U4067 (N_4067,N_3935,N_3997);
and U4068 (N_4068,N_3878,N_3842);
nand U4069 (N_4069,N_3877,N_3828);
and U4070 (N_4070,N_3820,N_3814);
nand U4071 (N_4071,N_3865,N_3961);
and U4072 (N_4072,N_3888,N_3907);
nor U4073 (N_4073,N_3950,N_3887);
or U4074 (N_4074,N_3808,N_3897);
and U4075 (N_4075,N_3861,N_3908);
xnor U4076 (N_4076,N_3864,N_3966);
and U4077 (N_4077,N_3883,N_3845);
nor U4078 (N_4078,N_3970,N_3978);
or U4079 (N_4079,N_3995,N_3931);
and U4080 (N_4080,N_3954,N_3928);
or U4081 (N_4081,N_3872,N_3937);
and U4082 (N_4082,N_3976,N_3818);
and U4083 (N_4083,N_3942,N_3844);
or U4084 (N_4084,N_3939,N_3925);
nor U4085 (N_4085,N_3869,N_3826);
or U4086 (N_4086,N_3860,N_3834);
nor U4087 (N_4087,N_3873,N_3854);
nor U4088 (N_4088,N_3933,N_3827);
and U4089 (N_4089,N_3993,N_3840);
or U4090 (N_4090,N_3938,N_3982);
or U4091 (N_4091,N_3800,N_3991);
or U4092 (N_4092,N_3894,N_3874);
nor U4093 (N_4093,N_3981,N_3964);
nor U4094 (N_4094,N_3841,N_3833);
and U4095 (N_4095,N_3803,N_3811);
nand U4096 (N_4096,N_3930,N_3881);
and U4097 (N_4097,N_3886,N_3923);
and U4098 (N_4098,N_3971,N_3832);
nand U4099 (N_4099,N_3999,N_3875);
and U4100 (N_4100,N_3854,N_3835);
or U4101 (N_4101,N_3914,N_3817);
nand U4102 (N_4102,N_3872,N_3962);
and U4103 (N_4103,N_3896,N_3902);
nor U4104 (N_4104,N_3971,N_3914);
and U4105 (N_4105,N_3823,N_3963);
or U4106 (N_4106,N_3892,N_3977);
and U4107 (N_4107,N_3905,N_3963);
or U4108 (N_4108,N_3888,N_3803);
and U4109 (N_4109,N_3927,N_3858);
and U4110 (N_4110,N_3864,N_3970);
or U4111 (N_4111,N_3893,N_3849);
and U4112 (N_4112,N_3804,N_3840);
or U4113 (N_4113,N_3889,N_3990);
xor U4114 (N_4114,N_3843,N_3818);
nand U4115 (N_4115,N_3856,N_3918);
xor U4116 (N_4116,N_3916,N_3958);
nand U4117 (N_4117,N_3834,N_3958);
nor U4118 (N_4118,N_3829,N_3905);
nor U4119 (N_4119,N_3947,N_3812);
or U4120 (N_4120,N_3846,N_3849);
and U4121 (N_4121,N_3973,N_3861);
or U4122 (N_4122,N_3851,N_3819);
and U4123 (N_4123,N_3805,N_3888);
and U4124 (N_4124,N_3939,N_3984);
nand U4125 (N_4125,N_3959,N_3835);
and U4126 (N_4126,N_3843,N_3905);
and U4127 (N_4127,N_3947,N_3840);
nand U4128 (N_4128,N_3996,N_3937);
nor U4129 (N_4129,N_3905,N_3844);
nor U4130 (N_4130,N_3906,N_3898);
and U4131 (N_4131,N_3919,N_3801);
and U4132 (N_4132,N_3871,N_3970);
and U4133 (N_4133,N_3909,N_3806);
nor U4134 (N_4134,N_3822,N_3848);
nor U4135 (N_4135,N_3870,N_3977);
or U4136 (N_4136,N_3994,N_3894);
or U4137 (N_4137,N_3978,N_3984);
and U4138 (N_4138,N_3847,N_3842);
and U4139 (N_4139,N_3880,N_3877);
nor U4140 (N_4140,N_3925,N_3892);
nand U4141 (N_4141,N_3847,N_3944);
or U4142 (N_4142,N_3990,N_3914);
and U4143 (N_4143,N_3964,N_3944);
nor U4144 (N_4144,N_3876,N_3921);
nor U4145 (N_4145,N_3983,N_3885);
and U4146 (N_4146,N_3818,N_3961);
and U4147 (N_4147,N_3983,N_3907);
and U4148 (N_4148,N_3860,N_3945);
nor U4149 (N_4149,N_3932,N_3893);
and U4150 (N_4150,N_3995,N_3848);
nor U4151 (N_4151,N_3856,N_3920);
and U4152 (N_4152,N_3992,N_3827);
or U4153 (N_4153,N_3907,N_3952);
and U4154 (N_4154,N_3983,N_3971);
or U4155 (N_4155,N_3856,N_3882);
nand U4156 (N_4156,N_3904,N_3892);
or U4157 (N_4157,N_3867,N_3885);
and U4158 (N_4158,N_3849,N_3986);
nand U4159 (N_4159,N_3915,N_3800);
nor U4160 (N_4160,N_3883,N_3930);
nor U4161 (N_4161,N_3863,N_3813);
and U4162 (N_4162,N_3800,N_3826);
nand U4163 (N_4163,N_3801,N_3838);
or U4164 (N_4164,N_3860,N_3814);
and U4165 (N_4165,N_3878,N_3982);
nand U4166 (N_4166,N_3952,N_3886);
nand U4167 (N_4167,N_3917,N_3814);
nand U4168 (N_4168,N_3829,N_3981);
nand U4169 (N_4169,N_3909,N_3893);
nor U4170 (N_4170,N_3906,N_3802);
and U4171 (N_4171,N_3868,N_3952);
and U4172 (N_4172,N_3902,N_3992);
nand U4173 (N_4173,N_3868,N_3878);
nor U4174 (N_4174,N_3812,N_3964);
or U4175 (N_4175,N_3966,N_3815);
nor U4176 (N_4176,N_3980,N_3991);
and U4177 (N_4177,N_3847,N_3889);
and U4178 (N_4178,N_3912,N_3956);
and U4179 (N_4179,N_3963,N_3995);
or U4180 (N_4180,N_3917,N_3910);
and U4181 (N_4181,N_3851,N_3961);
nor U4182 (N_4182,N_3901,N_3923);
or U4183 (N_4183,N_3847,N_3941);
and U4184 (N_4184,N_3811,N_3840);
or U4185 (N_4185,N_3838,N_3905);
and U4186 (N_4186,N_3899,N_3939);
or U4187 (N_4187,N_3821,N_3903);
nand U4188 (N_4188,N_3913,N_3823);
and U4189 (N_4189,N_3911,N_3800);
nand U4190 (N_4190,N_3996,N_3926);
and U4191 (N_4191,N_3968,N_3985);
or U4192 (N_4192,N_3979,N_3847);
and U4193 (N_4193,N_3931,N_3904);
nand U4194 (N_4194,N_3829,N_3957);
nand U4195 (N_4195,N_3980,N_3830);
or U4196 (N_4196,N_3930,N_3936);
nor U4197 (N_4197,N_3867,N_3832);
or U4198 (N_4198,N_3920,N_3842);
and U4199 (N_4199,N_3842,N_3927);
or U4200 (N_4200,N_4163,N_4070);
nand U4201 (N_4201,N_4158,N_4069);
nor U4202 (N_4202,N_4190,N_4109);
or U4203 (N_4203,N_4127,N_4099);
nor U4204 (N_4204,N_4112,N_4128);
nor U4205 (N_4205,N_4122,N_4004);
and U4206 (N_4206,N_4091,N_4040);
xnor U4207 (N_4207,N_4177,N_4056);
nand U4208 (N_4208,N_4125,N_4022);
nand U4209 (N_4209,N_4196,N_4150);
nand U4210 (N_4210,N_4073,N_4159);
nand U4211 (N_4211,N_4083,N_4072);
nor U4212 (N_4212,N_4198,N_4113);
or U4213 (N_4213,N_4088,N_4167);
nand U4214 (N_4214,N_4007,N_4059);
nand U4215 (N_4215,N_4042,N_4143);
xor U4216 (N_4216,N_4185,N_4155);
and U4217 (N_4217,N_4066,N_4027);
and U4218 (N_4218,N_4054,N_4001);
and U4219 (N_4219,N_4005,N_4195);
nor U4220 (N_4220,N_4010,N_4071);
nand U4221 (N_4221,N_4015,N_4009);
nor U4222 (N_4222,N_4117,N_4130);
and U4223 (N_4223,N_4183,N_4063);
and U4224 (N_4224,N_4081,N_4187);
or U4225 (N_4225,N_4030,N_4082);
and U4226 (N_4226,N_4132,N_4120);
or U4227 (N_4227,N_4131,N_4124);
and U4228 (N_4228,N_4067,N_4038);
or U4229 (N_4229,N_4079,N_4115);
or U4230 (N_4230,N_4126,N_4039);
or U4231 (N_4231,N_4094,N_4135);
nor U4232 (N_4232,N_4157,N_4044);
nand U4233 (N_4233,N_4080,N_4019);
or U4234 (N_4234,N_4175,N_4121);
and U4235 (N_4235,N_4003,N_4076);
nand U4236 (N_4236,N_4093,N_4043);
or U4237 (N_4237,N_4160,N_4164);
xnor U4238 (N_4238,N_4100,N_4193);
nand U4239 (N_4239,N_4165,N_4064);
or U4240 (N_4240,N_4045,N_4058);
xor U4241 (N_4241,N_4026,N_4057);
and U4242 (N_4242,N_4114,N_4116);
and U4243 (N_4243,N_4172,N_4171);
or U4244 (N_4244,N_4178,N_4169);
nor U4245 (N_4245,N_4184,N_4013);
or U4246 (N_4246,N_4104,N_4075);
nand U4247 (N_4247,N_4053,N_4181);
or U4248 (N_4248,N_4149,N_4014);
and U4249 (N_4249,N_4021,N_4061);
or U4250 (N_4250,N_4049,N_4096);
nand U4251 (N_4251,N_4050,N_4008);
and U4252 (N_4252,N_4029,N_4188);
or U4253 (N_4253,N_4174,N_4103);
and U4254 (N_4254,N_4134,N_4189);
nand U4255 (N_4255,N_4106,N_4191);
nand U4256 (N_4256,N_4148,N_4145);
and U4257 (N_4257,N_4031,N_4078);
nor U4258 (N_4258,N_4180,N_4118);
nor U4259 (N_4259,N_4192,N_4133);
nor U4260 (N_4260,N_4123,N_4156);
or U4261 (N_4261,N_4085,N_4146);
nand U4262 (N_4262,N_4089,N_4034);
xnor U4263 (N_4263,N_4102,N_4137);
and U4264 (N_4264,N_4147,N_4152);
nand U4265 (N_4265,N_4170,N_4168);
or U4266 (N_4266,N_4154,N_4197);
nor U4267 (N_4267,N_4000,N_4111);
or U4268 (N_4268,N_4176,N_4097);
and U4269 (N_4269,N_4173,N_4016);
or U4270 (N_4270,N_4140,N_4024);
nor U4271 (N_4271,N_4186,N_4153);
and U4272 (N_4272,N_4166,N_4002);
nand U4273 (N_4273,N_4141,N_4144);
or U4274 (N_4274,N_4161,N_4194);
nand U4275 (N_4275,N_4108,N_4138);
and U4276 (N_4276,N_4037,N_4062);
nor U4277 (N_4277,N_4129,N_4139);
and U4278 (N_4278,N_4048,N_4110);
nand U4279 (N_4279,N_4025,N_4199);
nand U4280 (N_4280,N_4006,N_4065);
nor U4281 (N_4281,N_4012,N_4101);
nor U4282 (N_4282,N_4035,N_4020);
and U4283 (N_4283,N_4060,N_4136);
nor U4284 (N_4284,N_4023,N_4107);
nor U4285 (N_4285,N_4046,N_4036);
and U4286 (N_4286,N_4162,N_4182);
or U4287 (N_4287,N_4028,N_4086);
or U4288 (N_4288,N_4032,N_4087);
or U4289 (N_4289,N_4041,N_4051);
nand U4290 (N_4290,N_4068,N_4033);
or U4291 (N_4291,N_4098,N_4017);
nor U4292 (N_4292,N_4092,N_4095);
and U4293 (N_4293,N_4179,N_4142);
nand U4294 (N_4294,N_4011,N_4084);
nor U4295 (N_4295,N_4119,N_4105);
nand U4296 (N_4296,N_4074,N_4090);
or U4297 (N_4297,N_4077,N_4151);
nor U4298 (N_4298,N_4052,N_4047);
nor U4299 (N_4299,N_4018,N_4055);
nand U4300 (N_4300,N_4101,N_4119);
or U4301 (N_4301,N_4047,N_4036);
or U4302 (N_4302,N_4048,N_4111);
nand U4303 (N_4303,N_4084,N_4102);
nand U4304 (N_4304,N_4040,N_4125);
nand U4305 (N_4305,N_4172,N_4164);
nor U4306 (N_4306,N_4009,N_4029);
nor U4307 (N_4307,N_4070,N_4041);
or U4308 (N_4308,N_4192,N_4022);
or U4309 (N_4309,N_4123,N_4108);
and U4310 (N_4310,N_4171,N_4190);
or U4311 (N_4311,N_4009,N_4183);
and U4312 (N_4312,N_4031,N_4083);
nor U4313 (N_4313,N_4008,N_4181);
nor U4314 (N_4314,N_4195,N_4124);
and U4315 (N_4315,N_4041,N_4161);
nand U4316 (N_4316,N_4100,N_4061);
nand U4317 (N_4317,N_4139,N_4007);
or U4318 (N_4318,N_4113,N_4019);
and U4319 (N_4319,N_4056,N_4084);
and U4320 (N_4320,N_4175,N_4028);
or U4321 (N_4321,N_4044,N_4137);
nand U4322 (N_4322,N_4058,N_4010);
nor U4323 (N_4323,N_4037,N_4057);
nor U4324 (N_4324,N_4190,N_4052);
nor U4325 (N_4325,N_4065,N_4016);
nand U4326 (N_4326,N_4059,N_4142);
nand U4327 (N_4327,N_4157,N_4098);
or U4328 (N_4328,N_4193,N_4160);
or U4329 (N_4329,N_4054,N_4102);
nor U4330 (N_4330,N_4059,N_4057);
nor U4331 (N_4331,N_4016,N_4095);
or U4332 (N_4332,N_4071,N_4011);
nor U4333 (N_4333,N_4110,N_4141);
nand U4334 (N_4334,N_4102,N_4174);
nand U4335 (N_4335,N_4032,N_4056);
or U4336 (N_4336,N_4087,N_4129);
and U4337 (N_4337,N_4089,N_4126);
or U4338 (N_4338,N_4016,N_4113);
xor U4339 (N_4339,N_4042,N_4167);
and U4340 (N_4340,N_4198,N_4032);
or U4341 (N_4341,N_4194,N_4140);
and U4342 (N_4342,N_4056,N_4052);
or U4343 (N_4343,N_4185,N_4084);
nand U4344 (N_4344,N_4102,N_4080);
or U4345 (N_4345,N_4040,N_4074);
or U4346 (N_4346,N_4146,N_4088);
and U4347 (N_4347,N_4198,N_4174);
or U4348 (N_4348,N_4095,N_4176);
and U4349 (N_4349,N_4134,N_4037);
nand U4350 (N_4350,N_4121,N_4188);
or U4351 (N_4351,N_4168,N_4156);
and U4352 (N_4352,N_4001,N_4031);
or U4353 (N_4353,N_4177,N_4001);
and U4354 (N_4354,N_4169,N_4064);
nor U4355 (N_4355,N_4097,N_4177);
and U4356 (N_4356,N_4139,N_4080);
nor U4357 (N_4357,N_4016,N_4059);
nand U4358 (N_4358,N_4097,N_4058);
and U4359 (N_4359,N_4132,N_4072);
nand U4360 (N_4360,N_4009,N_4073);
or U4361 (N_4361,N_4070,N_4066);
or U4362 (N_4362,N_4024,N_4058);
nor U4363 (N_4363,N_4141,N_4030);
nand U4364 (N_4364,N_4148,N_4138);
nand U4365 (N_4365,N_4161,N_4033);
nor U4366 (N_4366,N_4130,N_4097);
or U4367 (N_4367,N_4025,N_4133);
nand U4368 (N_4368,N_4003,N_4181);
nand U4369 (N_4369,N_4172,N_4055);
or U4370 (N_4370,N_4037,N_4080);
and U4371 (N_4371,N_4170,N_4080);
nand U4372 (N_4372,N_4104,N_4120);
and U4373 (N_4373,N_4091,N_4109);
or U4374 (N_4374,N_4002,N_4039);
nand U4375 (N_4375,N_4141,N_4149);
and U4376 (N_4376,N_4086,N_4060);
or U4377 (N_4377,N_4080,N_4095);
and U4378 (N_4378,N_4023,N_4096);
nor U4379 (N_4379,N_4144,N_4138);
or U4380 (N_4380,N_4017,N_4015);
nor U4381 (N_4381,N_4197,N_4088);
or U4382 (N_4382,N_4090,N_4068);
and U4383 (N_4383,N_4031,N_4176);
nand U4384 (N_4384,N_4156,N_4196);
or U4385 (N_4385,N_4027,N_4015);
nand U4386 (N_4386,N_4170,N_4192);
nand U4387 (N_4387,N_4072,N_4118);
and U4388 (N_4388,N_4030,N_4191);
or U4389 (N_4389,N_4133,N_4111);
nor U4390 (N_4390,N_4105,N_4087);
and U4391 (N_4391,N_4093,N_4063);
or U4392 (N_4392,N_4045,N_4056);
nand U4393 (N_4393,N_4079,N_4019);
nor U4394 (N_4394,N_4036,N_4027);
nor U4395 (N_4395,N_4108,N_4194);
nor U4396 (N_4396,N_4017,N_4025);
nand U4397 (N_4397,N_4168,N_4065);
nor U4398 (N_4398,N_4190,N_4045);
or U4399 (N_4399,N_4115,N_4000);
or U4400 (N_4400,N_4395,N_4371);
and U4401 (N_4401,N_4361,N_4324);
or U4402 (N_4402,N_4243,N_4200);
and U4403 (N_4403,N_4244,N_4260);
and U4404 (N_4404,N_4331,N_4364);
and U4405 (N_4405,N_4366,N_4261);
and U4406 (N_4406,N_4250,N_4391);
nor U4407 (N_4407,N_4272,N_4202);
nor U4408 (N_4408,N_4320,N_4216);
and U4409 (N_4409,N_4278,N_4349);
nand U4410 (N_4410,N_4303,N_4256);
or U4411 (N_4411,N_4280,N_4231);
and U4412 (N_4412,N_4360,N_4203);
and U4413 (N_4413,N_4228,N_4376);
or U4414 (N_4414,N_4368,N_4362);
and U4415 (N_4415,N_4253,N_4251);
nor U4416 (N_4416,N_4270,N_4227);
nand U4417 (N_4417,N_4305,N_4277);
and U4418 (N_4418,N_4327,N_4212);
or U4419 (N_4419,N_4295,N_4374);
or U4420 (N_4420,N_4334,N_4344);
nand U4421 (N_4421,N_4221,N_4220);
or U4422 (N_4422,N_4313,N_4271);
or U4423 (N_4423,N_4332,N_4259);
nand U4424 (N_4424,N_4241,N_4291);
or U4425 (N_4425,N_4399,N_4343);
or U4426 (N_4426,N_4325,N_4397);
and U4427 (N_4427,N_4205,N_4311);
or U4428 (N_4428,N_4326,N_4201);
nor U4429 (N_4429,N_4316,N_4385);
nand U4430 (N_4430,N_4266,N_4346);
or U4431 (N_4431,N_4392,N_4358);
and U4432 (N_4432,N_4314,N_4281);
and U4433 (N_4433,N_4211,N_4273);
nor U4434 (N_4434,N_4323,N_4245);
nor U4435 (N_4435,N_4351,N_4284);
nand U4436 (N_4436,N_4265,N_4379);
nor U4437 (N_4437,N_4263,N_4370);
nand U4438 (N_4438,N_4276,N_4315);
nand U4439 (N_4439,N_4381,N_4267);
nand U4440 (N_4440,N_4307,N_4290);
nor U4441 (N_4441,N_4369,N_4354);
or U4442 (N_4442,N_4380,N_4269);
nand U4443 (N_4443,N_4347,N_4384);
nand U4444 (N_4444,N_4240,N_4285);
nor U4445 (N_4445,N_4312,N_4268);
and U4446 (N_4446,N_4248,N_4298);
and U4447 (N_4447,N_4318,N_4333);
and U4448 (N_4448,N_4286,N_4338);
or U4449 (N_4449,N_4242,N_4210);
nand U4450 (N_4450,N_4279,N_4218);
nand U4451 (N_4451,N_4302,N_4225);
nand U4452 (N_4452,N_4206,N_4299);
and U4453 (N_4453,N_4319,N_4213);
nor U4454 (N_4454,N_4275,N_4317);
and U4455 (N_4455,N_4350,N_4223);
nand U4456 (N_4456,N_4306,N_4387);
nand U4457 (N_4457,N_4345,N_4356);
or U4458 (N_4458,N_4388,N_4342);
nand U4459 (N_4459,N_4247,N_4304);
or U4460 (N_4460,N_4322,N_4232);
and U4461 (N_4461,N_4217,N_4204);
and U4462 (N_4462,N_4238,N_4235);
and U4463 (N_4463,N_4294,N_4214);
and U4464 (N_4464,N_4289,N_4357);
nand U4465 (N_4465,N_4215,N_4230);
nor U4466 (N_4466,N_4321,N_4383);
and U4467 (N_4467,N_4389,N_4257);
nand U4468 (N_4468,N_4341,N_4352);
and U4469 (N_4469,N_4330,N_4239);
nor U4470 (N_4470,N_4229,N_4394);
nor U4471 (N_4471,N_4309,N_4301);
xnor U4472 (N_4472,N_4249,N_4207);
and U4473 (N_4473,N_4336,N_4372);
nand U4474 (N_4474,N_4282,N_4329);
or U4475 (N_4475,N_4288,N_4258);
nor U4476 (N_4476,N_4373,N_4222);
nand U4477 (N_4477,N_4292,N_4274);
nor U4478 (N_4478,N_4293,N_4308);
and U4479 (N_4479,N_4393,N_4252);
and U4480 (N_4480,N_4339,N_4254);
nand U4481 (N_4481,N_4287,N_4264);
nand U4482 (N_4482,N_4300,N_4390);
or U4483 (N_4483,N_4246,N_4348);
or U4484 (N_4484,N_4296,N_4396);
or U4485 (N_4485,N_4255,N_4233);
and U4486 (N_4486,N_4209,N_4224);
or U4487 (N_4487,N_4353,N_4226);
xnor U4488 (N_4488,N_4355,N_4378);
or U4489 (N_4489,N_4386,N_4262);
nand U4490 (N_4490,N_4377,N_4219);
and U4491 (N_4491,N_4297,N_4310);
or U4492 (N_4492,N_4367,N_4398);
and U4493 (N_4493,N_4340,N_4337);
nor U4494 (N_4494,N_4375,N_4365);
and U4495 (N_4495,N_4363,N_4359);
nand U4496 (N_4496,N_4328,N_4234);
xnor U4497 (N_4497,N_4335,N_4237);
and U4498 (N_4498,N_4208,N_4382);
or U4499 (N_4499,N_4283,N_4236);
or U4500 (N_4500,N_4385,N_4220);
nor U4501 (N_4501,N_4206,N_4272);
or U4502 (N_4502,N_4321,N_4280);
nor U4503 (N_4503,N_4253,N_4328);
and U4504 (N_4504,N_4327,N_4396);
nor U4505 (N_4505,N_4379,N_4206);
nor U4506 (N_4506,N_4360,N_4204);
and U4507 (N_4507,N_4319,N_4309);
nor U4508 (N_4508,N_4222,N_4240);
nor U4509 (N_4509,N_4219,N_4338);
or U4510 (N_4510,N_4280,N_4271);
nor U4511 (N_4511,N_4287,N_4371);
and U4512 (N_4512,N_4203,N_4221);
and U4513 (N_4513,N_4286,N_4276);
nor U4514 (N_4514,N_4206,N_4290);
and U4515 (N_4515,N_4228,N_4299);
or U4516 (N_4516,N_4244,N_4321);
and U4517 (N_4517,N_4244,N_4333);
and U4518 (N_4518,N_4345,N_4312);
nor U4519 (N_4519,N_4354,N_4269);
and U4520 (N_4520,N_4212,N_4266);
and U4521 (N_4521,N_4365,N_4370);
nand U4522 (N_4522,N_4351,N_4264);
nand U4523 (N_4523,N_4216,N_4228);
and U4524 (N_4524,N_4222,N_4273);
nor U4525 (N_4525,N_4374,N_4205);
or U4526 (N_4526,N_4203,N_4369);
nand U4527 (N_4527,N_4342,N_4361);
and U4528 (N_4528,N_4302,N_4315);
nor U4529 (N_4529,N_4227,N_4386);
or U4530 (N_4530,N_4318,N_4359);
or U4531 (N_4531,N_4314,N_4282);
and U4532 (N_4532,N_4253,N_4286);
and U4533 (N_4533,N_4374,N_4334);
or U4534 (N_4534,N_4273,N_4322);
and U4535 (N_4535,N_4201,N_4223);
nor U4536 (N_4536,N_4231,N_4247);
and U4537 (N_4537,N_4348,N_4257);
or U4538 (N_4538,N_4347,N_4389);
or U4539 (N_4539,N_4330,N_4304);
nand U4540 (N_4540,N_4298,N_4333);
and U4541 (N_4541,N_4351,N_4334);
or U4542 (N_4542,N_4378,N_4289);
nand U4543 (N_4543,N_4239,N_4284);
and U4544 (N_4544,N_4368,N_4252);
nor U4545 (N_4545,N_4246,N_4221);
nor U4546 (N_4546,N_4232,N_4253);
nand U4547 (N_4547,N_4287,N_4340);
nor U4548 (N_4548,N_4254,N_4283);
nor U4549 (N_4549,N_4249,N_4359);
and U4550 (N_4550,N_4252,N_4293);
and U4551 (N_4551,N_4288,N_4372);
and U4552 (N_4552,N_4258,N_4369);
and U4553 (N_4553,N_4325,N_4326);
nor U4554 (N_4554,N_4346,N_4234);
nor U4555 (N_4555,N_4306,N_4236);
or U4556 (N_4556,N_4388,N_4315);
nand U4557 (N_4557,N_4256,N_4263);
and U4558 (N_4558,N_4338,N_4227);
or U4559 (N_4559,N_4259,N_4370);
nor U4560 (N_4560,N_4360,N_4395);
nand U4561 (N_4561,N_4384,N_4224);
or U4562 (N_4562,N_4296,N_4362);
nand U4563 (N_4563,N_4213,N_4292);
or U4564 (N_4564,N_4390,N_4326);
nand U4565 (N_4565,N_4268,N_4280);
and U4566 (N_4566,N_4242,N_4318);
nand U4567 (N_4567,N_4325,N_4317);
nand U4568 (N_4568,N_4377,N_4265);
or U4569 (N_4569,N_4366,N_4382);
nand U4570 (N_4570,N_4229,N_4209);
or U4571 (N_4571,N_4362,N_4263);
or U4572 (N_4572,N_4324,N_4372);
or U4573 (N_4573,N_4231,N_4291);
and U4574 (N_4574,N_4291,N_4301);
and U4575 (N_4575,N_4205,N_4316);
and U4576 (N_4576,N_4252,N_4353);
nand U4577 (N_4577,N_4387,N_4377);
or U4578 (N_4578,N_4269,N_4260);
or U4579 (N_4579,N_4382,N_4361);
or U4580 (N_4580,N_4205,N_4289);
nand U4581 (N_4581,N_4367,N_4341);
nor U4582 (N_4582,N_4271,N_4254);
or U4583 (N_4583,N_4257,N_4242);
nor U4584 (N_4584,N_4304,N_4372);
nand U4585 (N_4585,N_4207,N_4317);
nand U4586 (N_4586,N_4216,N_4266);
nand U4587 (N_4587,N_4352,N_4368);
nor U4588 (N_4588,N_4285,N_4270);
or U4589 (N_4589,N_4214,N_4313);
nor U4590 (N_4590,N_4279,N_4324);
nor U4591 (N_4591,N_4389,N_4326);
or U4592 (N_4592,N_4325,N_4387);
nand U4593 (N_4593,N_4373,N_4295);
nand U4594 (N_4594,N_4376,N_4232);
nor U4595 (N_4595,N_4244,N_4388);
nand U4596 (N_4596,N_4282,N_4278);
nand U4597 (N_4597,N_4334,N_4321);
and U4598 (N_4598,N_4303,N_4299);
nor U4599 (N_4599,N_4207,N_4237);
or U4600 (N_4600,N_4521,N_4588);
nor U4601 (N_4601,N_4485,N_4538);
nor U4602 (N_4602,N_4537,N_4554);
nand U4603 (N_4603,N_4489,N_4497);
and U4604 (N_4604,N_4555,N_4490);
nor U4605 (N_4605,N_4518,N_4486);
nor U4606 (N_4606,N_4473,N_4585);
and U4607 (N_4607,N_4587,N_4406);
and U4608 (N_4608,N_4441,N_4590);
or U4609 (N_4609,N_4506,N_4461);
nand U4610 (N_4610,N_4469,N_4524);
nand U4611 (N_4611,N_4424,N_4557);
nor U4612 (N_4612,N_4454,N_4422);
and U4613 (N_4613,N_4581,N_4592);
nor U4614 (N_4614,N_4549,N_4546);
nor U4615 (N_4615,N_4455,N_4478);
and U4616 (N_4616,N_4523,N_4452);
or U4617 (N_4617,N_4453,N_4552);
and U4618 (N_4618,N_4421,N_4551);
or U4619 (N_4619,N_4545,N_4460);
and U4620 (N_4620,N_4423,N_4417);
nor U4621 (N_4621,N_4496,N_4571);
nor U4622 (N_4622,N_4542,N_4475);
nor U4623 (N_4623,N_4566,N_4410);
or U4624 (N_4624,N_4547,N_4465);
or U4625 (N_4625,N_4432,N_4535);
and U4626 (N_4626,N_4540,N_4401);
or U4627 (N_4627,N_4520,N_4408);
and U4628 (N_4628,N_4459,N_4517);
nor U4629 (N_4629,N_4526,N_4400);
nand U4630 (N_4630,N_4505,N_4456);
nor U4631 (N_4631,N_4499,N_4510);
nand U4632 (N_4632,N_4561,N_4580);
or U4633 (N_4633,N_4558,N_4501);
and U4634 (N_4634,N_4425,N_4527);
and U4635 (N_4635,N_4599,N_4576);
and U4636 (N_4636,N_4436,N_4467);
nor U4637 (N_4637,N_4569,N_4414);
or U4638 (N_4638,N_4463,N_4563);
and U4639 (N_4639,N_4420,N_4519);
or U4640 (N_4640,N_4534,N_4528);
or U4641 (N_4641,N_4468,N_4439);
nand U4642 (N_4642,N_4419,N_4462);
or U4643 (N_4643,N_4430,N_4582);
nand U4644 (N_4644,N_4573,N_4470);
nor U4645 (N_4645,N_4553,N_4597);
or U4646 (N_4646,N_4509,N_4416);
or U4647 (N_4647,N_4434,N_4536);
or U4648 (N_4648,N_4435,N_4595);
nor U4649 (N_4649,N_4516,N_4575);
and U4650 (N_4650,N_4570,N_4589);
or U4651 (N_4651,N_4476,N_4507);
and U4652 (N_4652,N_4495,N_4402);
or U4653 (N_4653,N_4531,N_4483);
nor U4654 (N_4654,N_4498,N_4480);
nor U4655 (N_4655,N_4568,N_4513);
and U4656 (N_4656,N_4464,N_4415);
and U4657 (N_4657,N_4488,N_4481);
or U4658 (N_4658,N_4466,N_4446);
or U4659 (N_4659,N_4412,N_4529);
nand U4660 (N_4660,N_4411,N_4550);
nor U4661 (N_4661,N_4404,N_4482);
nor U4662 (N_4662,N_4492,N_4515);
and U4663 (N_4663,N_4562,N_4450);
nor U4664 (N_4664,N_4447,N_4491);
and U4665 (N_4665,N_4451,N_4457);
nand U4666 (N_4666,N_4514,N_4533);
or U4667 (N_4667,N_4591,N_4403);
nand U4668 (N_4668,N_4578,N_4522);
nand U4669 (N_4669,N_4472,N_4502);
and U4670 (N_4670,N_4583,N_4598);
nand U4671 (N_4671,N_4444,N_4572);
and U4672 (N_4672,N_4449,N_4564);
and U4673 (N_4673,N_4503,N_4433);
and U4674 (N_4674,N_4577,N_4500);
and U4675 (N_4675,N_4479,N_4437);
nand U4676 (N_4676,N_4574,N_4541);
or U4677 (N_4677,N_4548,N_4484);
xor U4678 (N_4678,N_4477,N_4442);
nand U4679 (N_4679,N_4458,N_4407);
nand U4680 (N_4680,N_4594,N_4504);
and U4681 (N_4681,N_4487,N_4565);
nand U4682 (N_4682,N_4567,N_4596);
or U4683 (N_4683,N_4443,N_4429);
nor U4684 (N_4684,N_4448,N_4474);
and U4685 (N_4685,N_4438,N_4471);
nand U4686 (N_4686,N_4593,N_4560);
nand U4687 (N_4687,N_4544,N_4579);
or U4688 (N_4688,N_4445,N_4494);
nor U4689 (N_4689,N_4530,N_4508);
nor U4690 (N_4690,N_4512,N_4418);
and U4691 (N_4691,N_4493,N_4413);
nor U4692 (N_4692,N_4511,N_4426);
nor U4693 (N_4693,N_4428,N_4525);
and U4694 (N_4694,N_4409,N_4405);
and U4695 (N_4695,N_4440,N_4431);
and U4696 (N_4696,N_4586,N_4539);
or U4697 (N_4697,N_4559,N_4556);
nor U4698 (N_4698,N_4543,N_4427);
nand U4699 (N_4699,N_4532,N_4584);
or U4700 (N_4700,N_4425,N_4474);
nand U4701 (N_4701,N_4475,N_4555);
or U4702 (N_4702,N_4586,N_4535);
nor U4703 (N_4703,N_4412,N_4464);
nand U4704 (N_4704,N_4502,N_4554);
and U4705 (N_4705,N_4576,N_4447);
and U4706 (N_4706,N_4501,N_4487);
nand U4707 (N_4707,N_4405,N_4520);
nor U4708 (N_4708,N_4588,N_4579);
nand U4709 (N_4709,N_4445,N_4465);
nand U4710 (N_4710,N_4587,N_4516);
or U4711 (N_4711,N_4468,N_4533);
nand U4712 (N_4712,N_4477,N_4545);
nand U4713 (N_4713,N_4445,N_4440);
nand U4714 (N_4714,N_4403,N_4464);
and U4715 (N_4715,N_4591,N_4447);
or U4716 (N_4716,N_4497,N_4435);
nand U4717 (N_4717,N_4466,N_4433);
and U4718 (N_4718,N_4549,N_4562);
nand U4719 (N_4719,N_4553,N_4421);
or U4720 (N_4720,N_4511,N_4430);
nor U4721 (N_4721,N_4477,N_4402);
and U4722 (N_4722,N_4540,N_4449);
nor U4723 (N_4723,N_4478,N_4419);
and U4724 (N_4724,N_4527,N_4536);
or U4725 (N_4725,N_4471,N_4545);
nor U4726 (N_4726,N_4551,N_4460);
or U4727 (N_4727,N_4509,N_4452);
nor U4728 (N_4728,N_4579,N_4570);
nor U4729 (N_4729,N_4493,N_4535);
and U4730 (N_4730,N_4585,N_4556);
and U4731 (N_4731,N_4560,N_4409);
and U4732 (N_4732,N_4519,N_4499);
and U4733 (N_4733,N_4471,N_4533);
nand U4734 (N_4734,N_4506,N_4577);
nand U4735 (N_4735,N_4405,N_4441);
or U4736 (N_4736,N_4571,N_4465);
nand U4737 (N_4737,N_4562,N_4514);
nor U4738 (N_4738,N_4431,N_4444);
nand U4739 (N_4739,N_4453,N_4535);
nand U4740 (N_4740,N_4586,N_4528);
nand U4741 (N_4741,N_4463,N_4434);
and U4742 (N_4742,N_4495,N_4431);
or U4743 (N_4743,N_4550,N_4556);
nand U4744 (N_4744,N_4437,N_4498);
and U4745 (N_4745,N_4589,N_4427);
or U4746 (N_4746,N_4488,N_4410);
nand U4747 (N_4747,N_4482,N_4584);
nor U4748 (N_4748,N_4410,N_4518);
nor U4749 (N_4749,N_4474,N_4504);
nor U4750 (N_4750,N_4437,N_4449);
or U4751 (N_4751,N_4496,N_4537);
or U4752 (N_4752,N_4549,N_4446);
or U4753 (N_4753,N_4514,N_4502);
nor U4754 (N_4754,N_4586,N_4483);
and U4755 (N_4755,N_4514,N_4496);
and U4756 (N_4756,N_4424,N_4430);
nor U4757 (N_4757,N_4483,N_4596);
or U4758 (N_4758,N_4510,N_4593);
nand U4759 (N_4759,N_4546,N_4482);
or U4760 (N_4760,N_4535,N_4468);
xor U4761 (N_4761,N_4599,N_4566);
and U4762 (N_4762,N_4528,N_4478);
xnor U4763 (N_4763,N_4486,N_4571);
or U4764 (N_4764,N_4556,N_4538);
nand U4765 (N_4765,N_4487,N_4512);
and U4766 (N_4766,N_4555,N_4500);
and U4767 (N_4767,N_4541,N_4513);
or U4768 (N_4768,N_4512,N_4497);
nor U4769 (N_4769,N_4584,N_4499);
or U4770 (N_4770,N_4548,N_4530);
nor U4771 (N_4771,N_4542,N_4408);
nor U4772 (N_4772,N_4484,N_4540);
or U4773 (N_4773,N_4466,N_4479);
nor U4774 (N_4774,N_4463,N_4416);
nand U4775 (N_4775,N_4565,N_4566);
and U4776 (N_4776,N_4438,N_4469);
or U4777 (N_4777,N_4507,N_4512);
nand U4778 (N_4778,N_4516,N_4492);
nand U4779 (N_4779,N_4407,N_4584);
nand U4780 (N_4780,N_4514,N_4536);
and U4781 (N_4781,N_4568,N_4490);
nand U4782 (N_4782,N_4573,N_4594);
nand U4783 (N_4783,N_4543,N_4510);
nor U4784 (N_4784,N_4433,N_4489);
nand U4785 (N_4785,N_4477,N_4512);
and U4786 (N_4786,N_4563,N_4509);
and U4787 (N_4787,N_4446,N_4432);
or U4788 (N_4788,N_4440,N_4527);
and U4789 (N_4789,N_4487,N_4579);
nor U4790 (N_4790,N_4407,N_4443);
and U4791 (N_4791,N_4431,N_4491);
and U4792 (N_4792,N_4470,N_4452);
or U4793 (N_4793,N_4414,N_4593);
nand U4794 (N_4794,N_4540,N_4407);
nor U4795 (N_4795,N_4486,N_4477);
nand U4796 (N_4796,N_4560,N_4578);
or U4797 (N_4797,N_4561,N_4513);
nand U4798 (N_4798,N_4494,N_4554);
nand U4799 (N_4799,N_4585,N_4456);
or U4800 (N_4800,N_4603,N_4733);
and U4801 (N_4801,N_4762,N_4671);
or U4802 (N_4802,N_4796,N_4634);
and U4803 (N_4803,N_4629,N_4610);
nand U4804 (N_4804,N_4778,N_4740);
nand U4805 (N_4805,N_4627,N_4709);
and U4806 (N_4806,N_4789,N_4720);
or U4807 (N_4807,N_4798,N_4781);
nand U4808 (N_4808,N_4751,N_4677);
or U4809 (N_4809,N_4769,N_4742);
or U4810 (N_4810,N_4642,N_4719);
nand U4811 (N_4811,N_4646,N_4625);
and U4812 (N_4812,N_4743,N_4647);
nor U4813 (N_4813,N_4685,N_4702);
and U4814 (N_4814,N_4734,N_4665);
nor U4815 (N_4815,N_4669,N_4764);
nor U4816 (N_4816,N_4779,N_4620);
and U4817 (N_4817,N_4790,N_4687);
nor U4818 (N_4818,N_4694,N_4630);
or U4819 (N_4819,N_4739,N_4645);
nand U4820 (N_4820,N_4635,N_4722);
or U4821 (N_4821,N_4639,N_4636);
nand U4822 (N_4822,N_4650,N_4775);
or U4823 (N_4823,N_4651,N_4621);
nand U4824 (N_4824,N_4799,N_4721);
nand U4825 (N_4825,N_4717,N_4699);
nand U4826 (N_4826,N_4772,N_4628);
nor U4827 (N_4827,N_4787,N_4607);
and U4828 (N_4828,N_4725,N_4732);
nand U4829 (N_4829,N_4795,N_4623);
and U4830 (N_4830,N_4667,N_4797);
nand U4831 (N_4831,N_4766,N_4661);
nor U4832 (N_4832,N_4756,N_4640);
or U4833 (N_4833,N_4675,N_4604);
and U4834 (N_4834,N_4767,N_4741);
nor U4835 (N_4835,N_4729,N_4692);
or U4836 (N_4836,N_4689,N_4605);
nor U4837 (N_4837,N_4746,N_4684);
nor U4838 (N_4838,N_4668,N_4674);
nand U4839 (N_4839,N_4761,N_4785);
or U4840 (N_4840,N_4726,N_4637);
and U4841 (N_4841,N_4649,N_4664);
xnor U4842 (N_4842,N_4672,N_4614);
nor U4843 (N_4843,N_4784,N_4666);
nor U4844 (N_4844,N_4690,N_4745);
nor U4845 (N_4845,N_4632,N_4794);
or U4846 (N_4846,N_4612,N_4758);
nor U4847 (N_4847,N_4744,N_4703);
or U4848 (N_4848,N_4648,N_4670);
and U4849 (N_4849,N_4660,N_4633);
nor U4850 (N_4850,N_4792,N_4713);
nand U4851 (N_4851,N_4613,N_4680);
xnor U4852 (N_4852,N_4653,N_4738);
or U4853 (N_4853,N_4723,N_4747);
nand U4854 (N_4854,N_4724,N_4788);
nand U4855 (N_4855,N_4754,N_4735);
nor U4856 (N_4856,N_4730,N_4695);
nor U4857 (N_4857,N_4654,N_4652);
nand U4858 (N_4858,N_4656,N_4683);
or U4859 (N_4859,N_4609,N_4773);
nor U4860 (N_4860,N_4774,N_4716);
nor U4861 (N_4861,N_4658,N_4622);
or U4862 (N_4862,N_4606,N_4707);
nor U4863 (N_4863,N_4749,N_4748);
nor U4864 (N_4864,N_4678,N_4700);
and U4865 (N_4865,N_4681,N_4731);
or U4866 (N_4866,N_4686,N_4736);
and U4867 (N_4867,N_4641,N_4710);
and U4868 (N_4868,N_4701,N_4611);
nor U4869 (N_4869,N_4698,N_4659);
and U4870 (N_4870,N_4617,N_4624);
or U4871 (N_4871,N_4616,N_4708);
nor U4872 (N_4872,N_4786,N_4688);
or U4873 (N_4873,N_4768,N_4791);
and U4874 (N_4874,N_4602,N_4760);
and U4875 (N_4875,N_4759,N_4679);
nand U4876 (N_4876,N_4752,N_4601);
nand U4877 (N_4877,N_4780,N_4697);
or U4878 (N_4878,N_4608,N_4793);
xor U4879 (N_4879,N_4631,N_4643);
nor U4880 (N_4880,N_4655,N_4638);
nor U4881 (N_4881,N_4783,N_4691);
nand U4882 (N_4882,N_4676,N_4753);
nor U4883 (N_4883,N_4657,N_4704);
nand U4884 (N_4884,N_4619,N_4737);
nand U4885 (N_4885,N_4693,N_4770);
nand U4886 (N_4886,N_4711,N_4662);
nand U4887 (N_4887,N_4618,N_4600);
or U4888 (N_4888,N_4755,N_4705);
nand U4889 (N_4889,N_4615,N_4718);
nor U4890 (N_4890,N_4771,N_4763);
and U4891 (N_4891,N_4706,N_4782);
nand U4892 (N_4892,N_4626,N_4727);
and U4893 (N_4893,N_4696,N_4682);
and U4894 (N_4894,N_4728,N_4712);
or U4895 (N_4895,N_4714,N_4644);
nand U4896 (N_4896,N_4765,N_4663);
or U4897 (N_4897,N_4757,N_4777);
and U4898 (N_4898,N_4750,N_4776);
and U4899 (N_4899,N_4715,N_4673);
nand U4900 (N_4900,N_4746,N_4679);
or U4901 (N_4901,N_4725,N_4619);
nor U4902 (N_4902,N_4743,N_4714);
and U4903 (N_4903,N_4679,N_4637);
nand U4904 (N_4904,N_4688,N_4611);
nor U4905 (N_4905,N_4694,N_4732);
and U4906 (N_4906,N_4697,N_4687);
and U4907 (N_4907,N_4685,N_4679);
and U4908 (N_4908,N_4773,N_4635);
nand U4909 (N_4909,N_4738,N_4730);
and U4910 (N_4910,N_4604,N_4607);
and U4911 (N_4911,N_4647,N_4744);
nand U4912 (N_4912,N_4711,N_4628);
or U4913 (N_4913,N_4724,N_4719);
nor U4914 (N_4914,N_4618,N_4656);
nor U4915 (N_4915,N_4649,N_4633);
or U4916 (N_4916,N_4630,N_4708);
xnor U4917 (N_4917,N_4763,N_4633);
nor U4918 (N_4918,N_4722,N_4771);
and U4919 (N_4919,N_4743,N_4637);
nand U4920 (N_4920,N_4630,N_4706);
nor U4921 (N_4921,N_4771,N_4768);
nand U4922 (N_4922,N_4740,N_4761);
and U4923 (N_4923,N_4665,N_4723);
nand U4924 (N_4924,N_4791,N_4687);
or U4925 (N_4925,N_4775,N_4694);
and U4926 (N_4926,N_4664,N_4797);
nor U4927 (N_4927,N_4694,N_4607);
nand U4928 (N_4928,N_4693,N_4732);
nor U4929 (N_4929,N_4744,N_4684);
or U4930 (N_4930,N_4728,N_4694);
and U4931 (N_4931,N_4774,N_4664);
or U4932 (N_4932,N_4617,N_4792);
and U4933 (N_4933,N_4656,N_4660);
nor U4934 (N_4934,N_4621,N_4605);
nor U4935 (N_4935,N_4672,N_4675);
nor U4936 (N_4936,N_4672,N_4756);
and U4937 (N_4937,N_4667,N_4637);
nand U4938 (N_4938,N_4684,N_4789);
nor U4939 (N_4939,N_4793,N_4656);
and U4940 (N_4940,N_4606,N_4794);
nand U4941 (N_4941,N_4648,N_4707);
or U4942 (N_4942,N_4712,N_4658);
and U4943 (N_4943,N_4735,N_4621);
nor U4944 (N_4944,N_4701,N_4646);
nor U4945 (N_4945,N_4778,N_4780);
or U4946 (N_4946,N_4619,N_4611);
and U4947 (N_4947,N_4760,N_4731);
or U4948 (N_4948,N_4602,N_4651);
or U4949 (N_4949,N_4611,N_4618);
and U4950 (N_4950,N_4620,N_4716);
or U4951 (N_4951,N_4609,N_4634);
nand U4952 (N_4952,N_4666,N_4695);
nor U4953 (N_4953,N_4699,N_4680);
and U4954 (N_4954,N_4734,N_4691);
or U4955 (N_4955,N_4746,N_4750);
and U4956 (N_4956,N_4600,N_4702);
nor U4957 (N_4957,N_4723,N_4660);
nor U4958 (N_4958,N_4647,N_4799);
nor U4959 (N_4959,N_4617,N_4641);
nor U4960 (N_4960,N_4731,N_4645);
and U4961 (N_4961,N_4749,N_4655);
nor U4962 (N_4962,N_4602,N_4728);
nand U4963 (N_4963,N_4757,N_4635);
and U4964 (N_4964,N_4678,N_4611);
nor U4965 (N_4965,N_4750,N_4600);
and U4966 (N_4966,N_4750,N_4642);
nor U4967 (N_4967,N_4689,N_4625);
nor U4968 (N_4968,N_4612,N_4688);
or U4969 (N_4969,N_4610,N_4684);
nor U4970 (N_4970,N_4775,N_4783);
and U4971 (N_4971,N_4734,N_4736);
or U4972 (N_4972,N_4711,N_4776);
nand U4973 (N_4973,N_4732,N_4642);
or U4974 (N_4974,N_4635,N_4680);
nor U4975 (N_4975,N_4689,N_4600);
nor U4976 (N_4976,N_4771,N_4637);
nor U4977 (N_4977,N_4789,N_4708);
and U4978 (N_4978,N_4734,N_4613);
nand U4979 (N_4979,N_4714,N_4682);
and U4980 (N_4980,N_4714,N_4648);
or U4981 (N_4981,N_4704,N_4628);
nand U4982 (N_4982,N_4646,N_4731);
and U4983 (N_4983,N_4612,N_4728);
nor U4984 (N_4984,N_4776,N_4708);
nor U4985 (N_4985,N_4722,N_4751);
and U4986 (N_4986,N_4763,N_4681);
and U4987 (N_4987,N_4629,N_4631);
nor U4988 (N_4988,N_4627,N_4626);
or U4989 (N_4989,N_4746,N_4673);
or U4990 (N_4990,N_4685,N_4771);
and U4991 (N_4991,N_4672,N_4741);
and U4992 (N_4992,N_4715,N_4656);
nand U4993 (N_4993,N_4610,N_4701);
and U4994 (N_4994,N_4608,N_4700);
nand U4995 (N_4995,N_4712,N_4605);
nand U4996 (N_4996,N_4734,N_4792);
nor U4997 (N_4997,N_4726,N_4620);
or U4998 (N_4998,N_4684,N_4669);
nor U4999 (N_4999,N_4642,N_4783);
nor UO_0 (O_0,N_4819,N_4890);
nor UO_1 (O_1,N_4872,N_4905);
nand UO_2 (O_2,N_4839,N_4931);
nand UO_3 (O_3,N_4945,N_4984);
or UO_4 (O_4,N_4871,N_4996);
nor UO_5 (O_5,N_4937,N_4950);
and UO_6 (O_6,N_4850,N_4900);
or UO_7 (O_7,N_4969,N_4926);
and UO_8 (O_8,N_4800,N_4877);
nand UO_9 (O_9,N_4814,N_4927);
or UO_10 (O_10,N_4939,N_4868);
or UO_11 (O_11,N_4976,N_4902);
and UO_12 (O_12,N_4979,N_4854);
or UO_13 (O_13,N_4878,N_4919);
and UO_14 (O_14,N_4894,N_4887);
or UO_15 (O_15,N_4915,N_4823);
nand UO_16 (O_16,N_4825,N_4867);
nand UO_17 (O_17,N_4965,N_4882);
nor UO_18 (O_18,N_4893,N_4956);
or UO_19 (O_19,N_4891,N_4827);
nand UO_20 (O_20,N_4832,N_4949);
or UO_21 (O_21,N_4941,N_4855);
and UO_22 (O_22,N_4994,N_4828);
and UO_23 (O_23,N_4876,N_4859);
or UO_24 (O_24,N_4858,N_4865);
or UO_25 (O_25,N_4880,N_4920);
and UO_26 (O_26,N_4993,N_4845);
nor UO_27 (O_27,N_4881,N_4972);
nand UO_28 (O_28,N_4988,N_4982);
nand UO_29 (O_29,N_4930,N_4966);
nor UO_30 (O_30,N_4943,N_4816);
nor UO_31 (O_31,N_4909,N_4959);
and UO_32 (O_32,N_4961,N_4999);
nor UO_33 (O_33,N_4973,N_4852);
nand UO_34 (O_34,N_4960,N_4842);
and UO_35 (O_35,N_4903,N_4983);
or UO_36 (O_36,N_4913,N_4953);
nand UO_37 (O_37,N_4952,N_4862);
nand UO_38 (O_38,N_4992,N_4813);
nand UO_39 (O_39,N_4817,N_4940);
and UO_40 (O_40,N_4829,N_4808);
and UO_41 (O_41,N_4904,N_4921);
and UO_42 (O_42,N_4860,N_4818);
and UO_43 (O_43,N_4947,N_4998);
or UO_44 (O_44,N_4951,N_4923);
nor UO_45 (O_45,N_4869,N_4815);
nor UO_46 (O_46,N_4853,N_4824);
and UO_47 (O_47,N_4826,N_4901);
and UO_48 (O_48,N_4971,N_4884);
and UO_49 (O_49,N_4908,N_4886);
or UO_50 (O_50,N_4821,N_4914);
nand UO_51 (O_51,N_4948,N_4811);
or UO_52 (O_52,N_4985,N_4957);
or UO_53 (O_53,N_4989,N_4833);
or UO_54 (O_54,N_4840,N_4944);
nand UO_55 (O_55,N_4990,N_4954);
nand UO_56 (O_56,N_4977,N_4963);
nand UO_57 (O_57,N_4899,N_4975);
nor UO_58 (O_58,N_4929,N_4964);
or UO_59 (O_59,N_4834,N_4805);
and UO_60 (O_60,N_4968,N_4911);
or UO_61 (O_61,N_4883,N_4942);
and UO_62 (O_62,N_4897,N_4981);
xnor UO_63 (O_63,N_4925,N_4803);
and UO_64 (O_64,N_4922,N_4935);
nor UO_65 (O_65,N_4846,N_4932);
nor UO_66 (O_66,N_4830,N_4822);
nor UO_67 (O_67,N_4843,N_4831);
xnor UO_68 (O_68,N_4804,N_4916);
and UO_69 (O_69,N_4870,N_4906);
nor UO_70 (O_70,N_4807,N_4910);
nor UO_71 (O_71,N_4934,N_4851);
and UO_72 (O_72,N_4885,N_4962);
or UO_73 (O_73,N_4946,N_4907);
or UO_74 (O_74,N_4933,N_4918);
nor UO_75 (O_75,N_4812,N_4806);
and UO_76 (O_76,N_4837,N_4892);
nor UO_77 (O_77,N_4980,N_4866);
nor UO_78 (O_78,N_4874,N_4928);
nor UO_79 (O_79,N_4863,N_4848);
xor UO_80 (O_80,N_4967,N_4849);
or UO_81 (O_81,N_4889,N_4924);
nand UO_82 (O_82,N_4987,N_4912);
or UO_83 (O_83,N_4879,N_4856);
nor UO_84 (O_84,N_4802,N_4955);
or UO_85 (O_85,N_4978,N_4861);
nand UO_86 (O_86,N_4835,N_4917);
or UO_87 (O_87,N_4838,N_4898);
or UO_88 (O_88,N_4809,N_4896);
and UO_89 (O_89,N_4974,N_4936);
or UO_90 (O_90,N_4847,N_4970);
and UO_91 (O_91,N_4995,N_4888);
or UO_92 (O_92,N_4864,N_4841);
nor UO_93 (O_93,N_4991,N_4875);
and UO_94 (O_94,N_4836,N_4938);
nor UO_95 (O_95,N_4997,N_4873);
nor UO_96 (O_96,N_4810,N_4801);
nand UO_97 (O_97,N_4844,N_4895);
nor UO_98 (O_98,N_4857,N_4986);
and UO_99 (O_99,N_4958,N_4820);
nor UO_100 (O_100,N_4817,N_4945);
nor UO_101 (O_101,N_4837,N_4801);
and UO_102 (O_102,N_4996,N_4867);
and UO_103 (O_103,N_4861,N_4941);
nor UO_104 (O_104,N_4996,N_4997);
nand UO_105 (O_105,N_4916,N_4844);
nor UO_106 (O_106,N_4952,N_4842);
or UO_107 (O_107,N_4998,N_4889);
nor UO_108 (O_108,N_4938,N_4960);
and UO_109 (O_109,N_4866,N_4806);
and UO_110 (O_110,N_4965,N_4817);
and UO_111 (O_111,N_4882,N_4871);
nand UO_112 (O_112,N_4985,N_4855);
nor UO_113 (O_113,N_4826,N_4928);
and UO_114 (O_114,N_4932,N_4875);
nor UO_115 (O_115,N_4871,N_4838);
and UO_116 (O_116,N_4827,N_4999);
nand UO_117 (O_117,N_4842,N_4965);
or UO_118 (O_118,N_4882,N_4830);
and UO_119 (O_119,N_4960,N_4806);
or UO_120 (O_120,N_4875,N_4882);
or UO_121 (O_121,N_4850,N_4895);
or UO_122 (O_122,N_4811,N_4830);
or UO_123 (O_123,N_4810,N_4817);
nand UO_124 (O_124,N_4881,N_4853);
and UO_125 (O_125,N_4819,N_4866);
or UO_126 (O_126,N_4811,N_4941);
and UO_127 (O_127,N_4824,N_4862);
nand UO_128 (O_128,N_4803,N_4858);
and UO_129 (O_129,N_4892,N_4968);
or UO_130 (O_130,N_4992,N_4998);
nor UO_131 (O_131,N_4909,N_4806);
nand UO_132 (O_132,N_4835,N_4919);
or UO_133 (O_133,N_4897,N_4952);
and UO_134 (O_134,N_4869,N_4918);
or UO_135 (O_135,N_4972,N_4868);
and UO_136 (O_136,N_4983,N_4931);
or UO_137 (O_137,N_4950,N_4906);
and UO_138 (O_138,N_4927,N_4892);
nor UO_139 (O_139,N_4958,N_4844);
and UO_140 (O_140,N_4855,N_4809);
nor UO_141 (O_141,N_4877,N_4859);
and UO_142 (O_142,N_4865,N_4862);
or UO_143 (O_143,N_4847,N_4978);
nand UO_144 (O_144,N_4838,N_4851);
and UO_145 (O_145,N_4843,N_4997);
or UO_146 (O_146,N_4999,N_4839);
nor UO_147 (O_147,N_4898,N_4964);
or UO_148 (O_148,N_4871,N_4862);
nor UO_149 (O_149,N_4987,N_4835);
and UO_150 (O_150,N_4819,N_4899);
and UO_151 (O_151,N_4911,N_4988);
nand UO_152 (O_152,N_4938,N_4849);
nor UO_153 (O_153,N_4905,N_4876);
and UO_154 (O_154,N_4976,N_4819);
or UO_155 (O_155,N_4868,N_4922);
and UO_156 (O_156,N_4825,N_4947);
or UO_157 (O_157,N_4846,N_4989);
and UO_158 (O_158,N_4849,N_4925);
nand UO_159 (O_159,N_4946,N_4977);
nand UO_160 (O_160,N_4842,N_4982);
and UO_161 (O_161,N_4953,N_4926);
nor UO_162 (O_162,N_4965,N_4891);
or UO_163 (O_163,N_4909,N_4902);
nand UO_164 (O_164,N_4903,N_4821);
or UO_165 (O_165,N_4815,N_4935);
nor UO_166 (O_166,N_4967,N_4985);
nand UO_167 (O_167,N_4944,N_4979);
nor UO_168 (O_168,N_4866,N_4933);
and UO_169 (O_169,N_4967,N_4945);
and UO_170 (O_170,N_4814,N_4910);
nor UO_171 (O_171,N_4993,N_4800);
or UO_172 (O_172,N_4831,N_4892);
nand UO_173 (O_173,N_4891,N_4979);
nand UO_174 (O_174,N_4824,N_4977);
nand UO_175 (O_175,N_4999,N_4867);
or UO_176 (O_176,N_4852,N_4920);
and UO_177 (O_177,N_4884,N_4925);
nand UO_178 (O_178,N_4801,N_4853);
and UO_179 (O_179,N_4972,N_4804);
nand UO_180 (O_180,N_4864,N_4806);
and UO_181 (O_181,N_4919,N_4928);
nor UO_182 (O_182,N_4868,N_4892);
or UO_183 (O_183,N_4929,N_4895);
nor UO_184 (O_184,N_4899,N_4843);
and UO_185 (O_185,N_4889,N_4939);
nand UO_186 (O_186,N_4979,N_4916);
and UO_187 (O_187,N_4862,N_4954);
or UO_188 (O_188,N_4839,N_4994);
nand UO_189 (O_189,N_4844,N_4968);
or UO_190 (O_190,N_4947,N_4931);
nand UO_191 (O_191,N_4805,N_4923);
or UO_192 (O_192,N_4988,N_4996);
or UO_193 (O_193,N_4877,N_4885);
nor UO_194 (O_194,N_4820,N_4907);
or UO_195 (O_195,N_4850,N_4831);
nand UO_196 (O_196,N_4929,N_4876);
and UO_197 (O_197,N_4903,N_4824);
nor UO_198 (O_198,N_4915,N_4818);
nand UO_199 (O_199,N_4917,N_4905);
and UO_200 (O_200,N_4983,N_4933);
or UO_201 (O_201,N_4956,N_4959);
nand UO_202 (O_202,N_4915,N_4993);
and UO_203 (O_203,N_4839,N_4809);
or UO_204 (O_204,N_4937,N_4887);
and UO_205 (O_205,N_4908,N_4990);
or UO_206 (O_206,N_4842,N_4891);
and UO_207 (O_207,N_4834,N_4966);
xnor UO_208 (O_208,N_4894,N_4909);
nor UO_209 (O_209,N_4947,N_4859);
or UO_210 (O_210,N_4817,N_4939);
or UO_211 (O_211,N_4983,N_4955);
nand UO_212 (O_212,N_4906,N_4810);
nor UO_213 (O_213,N_4882,N_4909);
or UO_214 (O_214,N_4898,N_4951);
or UO_215 (O_215,N_4860,N_4876);
and UO_216 (O_216,N_4983,N_4888);
or UO_217 (O_217,N_4803,N_4903);
or UO_218 (O_218,N_4954,N_4981);
nand UO_219 (O_219,N_4956,N_4807);
or UO_220 (O_220,N_4898,N_4926);
nand UO_221 (O_221,N_4974,N_4887);
nand UO_222 (O_222,N_4858,N_4825);
and UO_223 (O_223,N_4807,N_4928);
or UO_224 (O_224,N_4800,N_4824);
and UO_225 (O_225,N_4935,N_4954);
or UO_226 (O_226,N_4944,N_4808);
nor UO_227 (O_227,N_4973,N_4987);
or UO_228 (O_228,N_4946,N_4962);
nand UO_229 (O_229,N_4896,N_4929);
and UO_230 (O_230,N_4918,N_4993);
nor UO_231 (O_231,N_4860,N_4995);
or UO_232 (O_232,N_4932,N_4818);
or UO_233 (O_233,N_4898,N_4808);
nand UO_234 (O_234,N_4814,N_4930);
nand UO_235 (O_235,N_4883,N_4801);
or UO_236 (O_236,N_4864,N_4973);
nor UO_237 (O_237,N_4848,N_4884);
nand UO_238 (O_238,N_4877,N_4840);
or UO_239 (O_239,N_4989,N_4982);
nand UO_240 (O_240,N_4847,N_4854);
nor UO_241 (O_241,N_4951,N_4837);
nor UO_242 (O_242,N_4802,N_4819);
and UO_243 (O_243,N_4852,N_4991);
nor UO_244 (O_244,N_4892,N_4877);
nand UO_245 (O_245,N_4823,N_4892);
or UO_246 (O_246,N_4810,N_4960);
and UO_247 (O_247,N_4871,N_4902);
nand UO_248 (O_248,N_4915,N_4902);
or UO_249 (O_249,N_4913,N_4979);
nor UO_250 (O_250,N_4832,N_4945);
or UO_251 (O_251,N_4906,N_4926);
nor UO_252 (O_252,N_4872,N_4871);
nor UO_253 (O_253,N_4931,N_4909);
nand UO_254 (O_254,N_4949,N_4923);
nand UO_255 (O_255,N_4804,N_4991);
or UO_256 (O_256,N_4833,N_4970);
xor UO_257 (O_257,N_4843,N_4812);
and UO_258 (O_258,N_4850,N_4902);
nand UO_259 (O_259,N_4994,N_4933);
nor UO_260 (O_260,N_4863,N_4914);
nand UO_261 (O_261,N_4933,N_4985);
and UO_262 (O_262,N_4865,N_4998);
nor UO_263 (O_263,N_4843,N_4977);
nor UO_264 (O_264,N_4942,N_4872);
nor UO_265 (O_265,N_4954,N_4833);
nand UO_266 (O_266,N_4865,N_4833);
or UO_267 (O_267,N_4886,N_4966);
and UO_268 (O_268,N_4874,N_4939);
and UO_269 (O_269,N_4954,N_4942);
and UO_270 (O_270,N_4818,N_4877);
nor UO_271 (O_271,N_4823,N_4984);
or UO_272 (O_272,N_4952,N_4861);
nand UO_273 (O_273,N_4831,N_4914);
nor UO_274 (O_274,N_4933,N_4915);
and UO_275 (O_275,N_4823,N_4943);
or UO_276 (O_276,N_4872,N_4953);
xor UO_277 (O_277,N_4946,N_4980);
and UO_278 (O_278,N_4979,N_4820);
nor UO_279 (O_279,N_4900,N_4950);
nand UO_280 (O_280,N_4834,N_4816);
nor UO_281 (O_281,N_4860,N_4884);
and UO_282 (O_282,N_4929,N_4980);
nand UO_283 (O_283,N_4844,N_4849);
nor UO_284 (O_284,N_4992,N_4911);
and UO_285 (O_285,N_4837,N_4901);
or UO_286 (O_286,N_4964,N_4850);
or UO_287 (O_287,N_4875,N_4934);
or UO_288 (O_288,N_4817,N_4926);
and UO_289 (O_289,N_4950,N_4851);
or UO_290 (O_290,N_4830,N_4999);
or UO_291 (O_291,N_4821,N_4961);
and UO_292 (O_292,N_4826,N_4833);
and UO_293 (O_293,N_4973,N_4935);
nand UO_294 (O_294,N_4992,N_4943);
or UO_295 (O_295,N_4821,N_4846);
and UO_296 (O_296,N_4995,N_4865);
nand UO_297 (O_297,N_4944,N_4829);
and UO_298 (O_298,N_4814,N_4911);
or UO_299 (O_299,N_4820,N_4960);
or UO_300 (O_300,N_4894,N_4840);
and UO_301 (O_301,N_4959,N_4876);
or UO_302 (O_302,N_4990,N_4880);
and UO_303 (O_303,N_4887,N_4966);
nor UO_304 (O_304,N_4976,N_4804);
and UO_305 (O_305,N_4903,N_4907);
or UO_306 (O_306,N_4902,N_4953);
nor UO_307 (O_307,N_4934,N_4896);
or UO_308 (O_308,N_4890,N_4820);
or UO_309 (O_309,N_4898,N_4891);
nor UO_310 (O_310,N_4921,N_4805);
and UO_311 (O_311,N_4975,N_4951);
and UO_312 (O_312,N_4853,N_4809);
nor UO_313 (O_313,N_4837,N_4900);
or UO_314 (O_314,N_4968,N_4852);
nand UO_315 (O_315,N_4880,N_4884);
nor UO_316 (O_316,N_4843,N_4873);
nand UO_317 (O_317,N_4988,N_4998);
nor UO_318 (O_318,N_4901,N_4944);
and UO_319 (O_319,N_4985,N_4825);
xor UO_320 (O_320,N_4852,N_4954);
nand UO_321 (O_321,N_4858,N_4938);
nand UO_322 (O_322,N_4889,N_4874);
nand UO_323 (O_323,N_4878,N_4855);
and UO_324 (O_324,N_4910,N_4903);
and UO_325 (O_325,N_4848,N_4895);
xnor UO_326 (O_326,N_4948,N_4825);
xnor UO_327 (O_327,N_4972,N_4986);
nor UO_328 (O_328,N_4991,N_4839);
nand UO_329 (O_329,N_4944,N_4981);
and UO_330 (O_330,N_4940,N_4961);
nor UO_331 (O_331,N_4961,N_4998);
or UO_332 (O_332,N_4856,N_4830);
nand UO_333 (O_333,N_4978,N_4858);
nand UO_334 (O_334,N_4805,N_4943);
nor UO_335 (O_335,N_4832,N_4985);
nor UO_336 (O_336,N_4993,N_4990);
and UO_337 (O_337,N_4876,N_4925);
or UO_338 (O_338,N_4947,N_4959);
nand UO_339 (O_339,N_4884,N_4986);
nor UO_340 (O_340,N_4948,N_4991);
or UO_341 (O_341,N_4898,N_4821);
nand UO_342 (O_342,N_4886,N_4943);
nand UO_343 (O_343,N_4879,N_4961);
nor UO_344 (O_344,N_4802,N_4839);
nor UO_345 (O_345,N_4924,N_4919);
or UO_346 (O_346,N_4902,N_4961);
nor UO_347 (O_347,N_4965,N_4930);
nor UO_348 (O_348,N_4970,N_4997);
and UO_349 (O_349,N_4834,N_4901);
and UO_350 (O_350,N_4961,N_4820);
or UO_351 (O_351,N_4922,N_4906);
nor UO_352 (O_352,N_4983,N_4920);
nand UO_353 (O_353,N_4805,N_4987);
nor UO_354 (O_354,N_4826,N_4987);
nor UO_355 (O_355,N_4963,N_4876);
and UO_356 (O_356,N_4983,N_4880);
nor UO_357 (O_357,N_4966,N_4816);
nand UO_358 (O_358,N_4959,N_4967);
nand UO_359 (O_359,N_4971,N_4863);
nand UO_360 (O_360,N_4829,N_4870);
or UO_361 (O_361,N_4851,N_4873);
nor UO_362 (O_362,N_4919,N_4870);
or UO_363 (O_363,N_4813,N_4859);
or UO_364 (O_364,N_4976,N_4941);
nand UO_365 (O_365,N_4989,N_4949);
or UO_366 (O_366,N_4983,N_4934);
nor UO_367 (O_367,N_4908,N_4826);
nor UO_368 (O_368,N_4849,N_4896);
or UO_369 (O_369,N_4990,N_4915);
nand UO_370 (O_370,N_4952,N_4889);
nor UO_371 (O_371,N_4994,N_4932);
and UO_372 (O_372,N_4910,N_4849);
or UO_373 (O_373,N_4992,N_4901);
nor UO_374 (O_374,N_4894,N_4821);
or UO_375 (O_375,N_4854,N_4859);
and UO_376 (O_376,N_4810,N_4990);
and UO_377 (O_377,N_4974,N_4814);
nand UO_378 (O_378,N_4910,N_4941);
nand UO_379 (O_379,N_4987,N_4964);
nand UO_380 (O_380,N_4835,N_4926);
and UO_381 (O_381,N_4853,N_4938);
nor UO_382 (O_382,N_4990,N_4921);
nor UO_383 (O_383,N_4955,N_4828);
nand UO_384 (O_384,N_4803,N_4820);
nand UO_385 (O_385,N_4809,N_4967);
or UO_386 (O_386,N_4879,N_4901);
or UO_387 (O_387,N_4826,N_4829);
nand UO_388 (O_388,N_4811,N_4931);
nor UO_389 (O_389,N_4837,N_4987);
or UO_390 (O_390,N_4911,N_4842);
or UO_391 (O_391,N_4853,N_4816);
and UO_392 (O_392,N_4972,N_4979);
nor UO_393 (O_393,N_4930,N_4873);
nand UO_394 (O_394,N_4878,N_4815);
and UO_395 (O_395,N_4931,N_4888);
nor UO_396 (O_396,N_4862,N_4892);
nor UO_397 (O_397,N_4932,N_4935);
nor UO_398 (O_398,N_4948,N_4821);
and UO_399 (O_399,N_4971,N_4846);
nand UO_400 (O_400,N_4947,N_4991);
and UO_401 (O_401,N_4811,N_4923);
nand UO_402 (O_402,N_4907,N_4807);
nor UO_403 (O_403,N_4916,N_4870);
or UO_404 (O_404,N_4995,N_4881);
or UO_405 (O_405,N_4828,N_4891);
nor UO_406 (O_406,N_4882,N_4985);
nand UO_407 (O_407,N_4871,N_4869);
nand UO_408 (O_408,N_4901,N_4871);
and UO_409 (O_409,N_4995,N_4937);
nand UO_410 (O_410,N_4972,N_4831);
or UO_411 (O_411,N_4906,N_4878);
or UO_412 (O_412,N_4988,N_4939);
nand UO_413 (O_413,N_4821,N_4923);
nand UO_414 (O_414,N_4839,N_4950);
nand UO_415 (O_415,N_4965,N_4872);
or UO_416 (O_416,N_4871,N_4940);
nor UO_417 (O_417,N_4996,N_4986);
nand UO_418 (O_418,N_4938,N_4870);
xnor UO_419 (O_419,N_4949,N_4964);
or UO_420 (O_420,N_4952,N_4893);
and UO_421 (O_421,N_4930,N_4904);
or UO_422 (O_422,N_4905,N_4912);
and UO_423 (O_423,N_4841,N_4970);
nand UO_424 (O_424,N_4937,N_4990);
nor UO_425 (O_425,N_4984,N_4836);
nor UO_426 (O_426,N_4932,N_4967);
and UO_427 (O_427,N_4933,N_4832);
nor UO_428 (O_428,N_4987,N_4857);
or UO_429 (O_429,N_4934,N_4923);
or UO_430 (O_430,N_4951,N_4850);
nor UO_431 (O_431,N_4823,N_4830);
nor UO_432 (O_432,N_4910,N_4960);
and UO_433 (O_433,N_4954,N_4839);
nor UO_434 (O_434,N_4814,N_4894);
and UO_435 (O_435,N_4826,N_4878);
and UO_436 (O_436,N_4917,N_4889);
and UO_437 (O_437,N_4851,N_4963);
and UO_438 (O_438,N_4929,N_4962);
nor UO_439 (O_439,N_4889,N_4996);
and UO_440 (O_440,N_4880,N_4955);
and UO_441 (O_441,N_4917,N_4983);
nor UO_442 (O_442,N_4871,N_4860);
nand UO_443 (O_443,N_4953,N_4860);
nor UO_444 (O_444,N_4976,N_4883);
xor UO_445 (O_445,N_4811,N_4969);
nor UO_446 (O_446,N_4986,N_4965);
or UO_447 (O_447,N_4812,N_4895);
nor UO_448 (O_448,N_4980,N_4856);
nor UO_449 (O_449,N_4848,N_4988);
and UO_450 (O_450,N_4822,N_4800);
or UO_451 (O_451,N_4807,N_4986);
nor UO_452 (O_452,N_4838,N_4864);
or UO_453 (O_453,N_4872,N_4969);
or UO_454 (O_454,N_4889,N_4902);
and UO_455 (O_455,N_4972,N_4871);
and UO_456 (O_456,N_4927,N_4813);
nand UO_457 (O_457,N_4966,N_4804);
or UO_458 (O_458,N_4828,N_4841);
and UO_459 (O_459,N_4872,N_4810);
and UO_460 (O_460,N_4800,N_4948);
nand UO_461 (O_461,N_4853,N_4983);
and UO_462 (O_462,N_4827,N_4852);
or UO_463 (O_463,N_4802,N_4886);
or UO_464 (O_464,N_4846,N_4980);
and UO_465 (O_465,N_4836,N_4998);
nand UO_466 (O_466,N_4878,N_4993);
nand UO_467 (O_467,N_4842,N_4846);
nor UO_468 (O_468,N_4905,N_4907);
nor UO_469 (O_469,N_4866,N_4932);
nand UO_470 (O_470,N_4957,N_4963);
nand UO_471 (O_471,N_4945,N_4846);
nor UO_472 (O_472,N_4849,N_4980);
and UO_473 (O_473,N_4991,N_4945);
nand UO_474 (O_474,N_4831,N_4981);
and UO_475 (O_475,N_4959,N_4969);
nor UO_476 (O_476,N_4924,N_4974);
nand UO_477 (O_477,N_4922,N_4927);
or UO_478 (O_478,N_4863,N_4937);
nor UO_479 (O_479,N_4912,N_4871);
or UO_480 (O_480,N_4842,N_4953);
nand UO_481 (O_481,N_4844,N_4886);
and UO_482 (O_482,N_4994,N_4920);
nor UO_483 (O_483,N_4966,N_4972);
nand UO_484 (O_484,N_4961,N_4964);
or UO_485 (O_485,N_4920,N_4842);
and UO_486 (O_486,N_4925,N_4813);
or UO_487 (O_487,N_4861,N_4841);
or UO_488 (O_488,N_4829,N_4966);
nor UO_489 (O_489,N_4811,N_4925);
nor UO_490 (O_490,N_4983,N_4816);
and UO_491 (O_491,N_4882,N_4993);
nor UO_492 (O_492,N_4871,N_4890);
or UO_493 (O_493,N_4890,N_4802);
or UO_494 (O_494,N_4847,N_4897);
nor UO_495 (O_495,N_4977,N_4990);
or UO_496 (O_496,N_4809,N_4867);
and UO_497 (O_497,N_4837,N_4932);
nand UO_498 (O_498,N_4963,N_4894);
nand UO_499 (O_499,N_4969,N_4846);
nor UO_500 (O_500,N_4983,N_4843);
nand UO_501 (O_501,N_4871,N_4837);
nand UO_502 (O_502,N_4860,N_4887);
nor UO_503 (O_503,N_4835,N_4973);
or UO_504 (O_504,N_4977,N_4936);
nor UO_505 (O_505,N_4891,N_4853);
nor UO_506 (O_506,N_4863,N_4807);
or UO_507 (O_507,N_4964,N_4924);
or UO_508 (O_508,N_4865,N_4892);
nand UO_509 (O_509,N_4949,N_4903);
or UO_510 (O_510,N_4970,N_4864);
nor UO_511 (O_511,N_4969,N_4995);
and UO_512 (O_512,N_4878,N_4890);
nand UO_513 (O_513,N_4914,N_4843);
nand UO_514 (O_514,N_4875,N_4863);
or UO_515 (O_515,N_4996,N_4891);
or UO_516 (O_516,N_4910,N_4994);
or UO_517 (O_517,N_4839,N_4920);
nand UO_518 (O_518,N_4919,N_4984);
nor UO_519 (O_519,N_4848,N_4938);
and UO_520 (O_520,N_4936,N_4806);
or UO_521 (O_521,N_4870,N_4841);
and UO_522 (O_522,N_4908,N_4945);
nand UO_523 (O_523,N_4927,N_4995);
nand UO_524 (O_524,N_4801,N_4902);
and UO_525 (O_525,N_4844,N_4871);
nor UO_526 (O_526,N_4804,N_4872);
nor UO_527 (O_527,N_4864,N_4924);
nor UO_528 (O_528,N_4955,N_4939);
nand UO_529 (O_529,N_4828,N_4812);
nor UO_530 (O_530,N_4813,N_4822);
nor UO_531 (O_531,N_4821,N_4924);
nor UO_532 (O_532,N_4959,N_4994);
nor UO_533 (O_533,N_4916,N_4909);
nor UO_534 (O_534,N_4852,N_4976);
or UO_535 (O_535,N_4887,N_4825);
nor UO_536 (O_536,N_4994,N_4988);
or UO_537 (O_537,N_4951,N_4823);
and UO_538 (O_538,N_4845,N_4898);
nand UO_539 (O_539,N_4972,N_4939);
or UO_540 (O_540,N_4951,N_4962);
nand UO_541 (O_541,N_4927,N_4948);
or UO_542 (O_542,N_4839,N_4858);
or UO_543 (O_543,N_4898,N_4837);
and UO_544 (O_544,N_4849,N_4816);
nor UO_545 (O_545,N_4895,N_4898);
or UO_546 (O_546,N_4813,N_4867);
nor UO_547 (O_547,N_4840,N_4990);
and UO_548 (O_548,N_4860,N_4848);
and UO_549 (O_549,N_4952,N_4969);
and UO_550 (O_550,N_4848,N_4872);
and UO_551 (O_551,N_4905,N_4913);
and UO_552 (O_552,N_4913,N_4986);
and UO_553 (O_553,N_4857,N_4930);
or UO_554 (O_554,N_4907,N_4956);
and UO_555 (O_555,N_4846,N_4931);
and UO_556 (O_556,N_4977,N_4840);
nand UO_557 (O_557,N_4957,N_4966);
nand UO_558 (O_558,N_4815,N_4981);
nand UO_559 (O_559,N_4985,N_4870);
or UO_560 (O_560,N_4997,N_4815);
nand UO_561 (O_561,N_4874,N_4908);
nor UO_562 (O_562,N_4845,N_4818);
nand UO_563 (O_563,N_4951,N_4833);
nor UO_564 (O_564,N_4972,N_4968);
and UO_565 (O_565,N_4814,N_4913);
nor UO_566 (O_566,N_4965,N_4966);
and UO_567 (O_567,N_4859,N_4872);
nand UO_568 (O_568,N_4837,N_4953);
and UO_569 (O_569,N_4838,N_4868);
nand UO_570 (O_570,N_4888,N_4915);
nor UO_571 (O_571,N_4800,N_4977);
and UO_572 (O_572,N_4907,N_4869);
nor UO_573 (O_573,N_4826,N_4891);
nor UO_574 (O_574,N_4901,N_4881);
or UO_575 (O_575,N_4856,N_4976);
or UO_576 (O_576,N_4835,N_4887);
or UO_577 (O_577,N_4826,N_4980);
and UO_578 (O_578,N_4851,N_4900);
nand UO_579 (O_579,N_4944,N_4922);
nor UO_580 (O_580,N_4852,N_4849);
nand UO_581 (O_581,N_4968,N_4817);
or UO_582 (O_582,N_4820,N_4983);
nand UO_583 (O_583,N_4862,N_4975);
nand UO_584 (O_584,N_4821,N_4925);
nand UO_585 (O_585,N_4984,N_4873);
nor UO_586 (O_586,N_4837,N_4922);
or UO_587 (O_587,N_4832,N_4911);
nor UO_588 (O_588,N_4998,N_4872);
nor UO_589 (O_589,N_4807,N_4901);
nor UO_590 (O_590,N_4810,N_4896);
and UO_591 (O_591,N_4823,N_4838);
nor UO_592 (O_592,N_4914,N_4855);
nor UO_593 (O_593,N_4827,N_4830);
nand UO_594 (O_594,N_4978,N_4971);
and UO_595 (O_595,N_4934,N_4878);
and UO_596 (O_596,N_4844,N_4811);
nand UO_597 (O_597,N_4974,N_4962);
nand UO_598 (O_598,N_4894,N_4988);
nor UO_599 (O_599,N_4915,N_4942);
or UO_600 (O_600,N_4997,N_4856);
nor UO_601 (O_601,N_4866,N_4975);
or UO_602 (O_602,N_4960,N_4975);
and UO_603 (O_603,N_4907,N_4865);
and UO_604 (O_604,N_4976,N_4855);
and UO_605 (O_605,N_4935,N_4837);
nor UO_606 (O_606,N_4911,N_4876);
nand UO_607 (O_607,N_4949,N_4822);
and UO_608 (O_608,N_4907,N_4866);
nand UO_609 (O_609,N_4867,N_4846);
nor UO_610 (O_610,N_4956,N_4809);
nor UO_611 (O_611,N_4929,N_4863);
or UO_612 (O_612,N_4830,N_4866);
nor UO_613 (O_613,N_4809,N_4898);
nor UO_614 (O_614,N_4992,N_4969);
or UO_615 (O_615,N_4983,N_4817);
nor UO_616 (O_616,N_4949,N_4915);
nor UO_617 (O_617,N_4849,N_4841);
nor UO_618 (O_618,N_4996,N_4838);
nor UO_619 (O_619,N_4832,N_4817);
or UO_620 (O_620,N_4970,N_4886);
and UO_621 (O_621,N_4819,N_4959);
and UO_622 (O_622,N_4995,N_4914);
or UO_623 (O_623,N_4888,N_4887);
or UO_624 (O_624,N_4850,N_4944);
or UO_625 (O_625,N_4895,N_4836);
nand UO_626 (O_626,N_4859,N_4988);
or UO_627 (O_627,N_4942,N_4936);
nand UO_628 (O_628,N_4922,N_4831);
nor UO_629 (O_629,N_4947,N_4873);
and UO_630 (O_630,N_4920,N_4838);
and UO_631 (O_631,N_4869,N_4823);
nand UO_632 (O_632,N_4813,N_4857);
nand UO_633 (O_633,N_4926,N_4859);
or UO_634 (O_634,N_4836,N_4855);
or UO_635 (O_635,N_4889,N_4887);
nand UO_636 (O_636,N_4905,N_4916);
nor UO_637 (O_637,N_4866,N_4936);
nand UO_638 (O_638,N_4903,N_4970);
nor UO_639 (O_639,N_4900,N_4912);
and UO_640 (O_640,N_4942,N_4902);
nor UO_641 (O_641,N_4899,N_4847);
and UO_642 (O_642,N_4995,N_4862);
nand UO_643 (O_643,N_4915,N_4812);
or UO_644 (O_644,N_4986,N_4937);
or UO_645 (O_645,N_4851,N_4841);
and UO_646 (O_646,N_4999,N_4918);
nor UO_647 (O_647,N_4909,N_4805);
nand UO_648 (O_648,N_4991,N_4812);
nand UO_649 (O_649,N_4883,N_4987);
and UO_650 (O_650,N_4871,N_4977);
nand UO_651 (O_651,N_4877,N_4918);
nand UO_652 (O_652,N_4899,N_4889);
nand UO_653 (O_653,N_4866,N_4909);
nand UO_654 (O_654,N_4961,N_4900);
nand UO_655 (O_655,N_4967,N_4803);
nand UO_656 (O_656,N_4854,N_4965);
and UO_657 (O_657,N_4879,N_4862);
and UO_658 (O_658,N_4933,N_4996);
and UO_659 (O_659,N_4866,N_4950);
or UO_660 (O_660,N_4874,N_4905);
and UO_661 (O_661,N_4897,N_4950);
or UO_662 (O_662,N_4837,N_4804);
or UO_663 (O_663,N_4836,N_4915);
nor UO_664 (O_664,N_4857,N_4834);
nand UO_665 (O_665,N_4968,N_4926);
and UO_666 (O_666,N_4972,N_4865);
or UO_667 (O_667,N_4970,N_4920);
nor UO_668 (O_668,N_4911,N_4852);
nor UO_669 (O_669,N_4921,N_4910);
nand UO_670 (O_670,N_4834,N_4935);
nor UO_671 (O_671,N_4905,N_4816);
or UO_672 (O_672,N_4979,N_4930);
nor UO_673 (O_673,N_4813,N_4825);
and UO_674 (O_674,N_4979,N_4864);
and UO_675 (O_675,N_4841,N_4961);
nor UO_676 (O_676,N_4823,N_4891);
and UO_677 (O_677,N_4895,N_4810);
and UO_678 (O_678,N_4922,N_4822);
or UO_679 (O_679,N_4858,N_4962);
nor UO_680 (O_680,N_4946,N_4821);
or UO_681 (O_681,N_4959,N_4892);
nor UO_682 (O_682,N_4937,N_4892);
nor UO_683 (O_683,N_4933,N_4955);
and UO_684 (O_684,N_4881,N_4894);
nor UO_685 (O_685,N_4905,N_4992);
and UO_686 (O_686,N_4900,N_4889);
and UO_687 (O_687,N_4824,N_4905);
nor UO_688 (O_688,N_4955,N_4919);
nor UO_689 (O_689,N_4836,N_4817);
nor UO_690 (O_690,N_4912,N_4881);
nand UO_691 (O_691,N_4843,N_4963);
or UO_692 (O_692,N_4896,N_4867);
and UO_693 (O_693,N_4839,N_4915);
nor UO_694 (O_694,N_4945,N_4985);
nor UO_695 (O_695,N_4895,N_4843);
or UO_696 (O_696,N_4868,N_4882);
and UO_697 (O_697,N_4986,N_4821);
xnor UO_698 (O_698,N_4957,N_4816);
and UO_699 (O_699,N_4906,N_4821);
or UO_700 (O_700,N_4971,N_4907);
or UO_701 (O_701,N_4977,N_4802);
or UO_702 (O_702,N_4907,N_4873);
or UO_703 (O_703,N_4940,N_4986);
nor UO_704 (O_704,N_4855,N_4987);
nand UO_705 (O_705,N_4843,N_4810);
nand UO_706 (O_706,N_4841,N_4835);
nor UO_707 (O_707,N_4920,N_4840);
or UO_708 (O_708,N_4940,N_4882);
or UO_709 (O_709,N_4991,N_4850);
and UO_710 (O_710,N_4934,N_4981);
or UO_711 (O_711,N_4918,N_4952);
and UO_712 (O_712,N_4872,N_4889);
nor UO_713 (O_713,N_4858,N_4994);
or UO_714 (O_714,N_4951,N_4999);
and UO_715 (O_715,N_4992,N_4828);
nand UO_716 (O_716,N_4871,N_4892);
and UO_717 (O_717,N_4852,N_4875);
or UO_718 (O_718,N_4841,N_4882);
nor UO_719 (O_719,N_4929,N_4933);
nand UO_720 (O_720,N_4863,N_4907);
or UO_721 (O_721,N_4903,N_4918);
nor UO_722 (O_722,N_4989,N_4968);
and UO_723 (O_723,N_4998,N_4966);
nor UO_724 (O_724,N_4983,N_4987);
nand UO_725 (O_725,N_4998,N_4804);
and UO_726 (O_726,N_4833,N_4987);
nor UO_727 (O_727,N_4986,N_4825);
or UO_728 (O_728,N_4883,N_4893);
or UO_729 (O_729,N_4885,N_4880);
and UO_730 (O_730,N_4969,N_4937);
or UO_731 (O_731,N_4851,N_4919);
nand UO_732 (O_732,N_4862,N_4909);
or UO_733 (O_733,N_4942,N_4847);
and UO_734 (O_734,N_4869,N_4954);
nor UO_735 (O_735,N_4802,N_4830);
nor UO_736 (O_736,N_4900,N_4997);
nor UO_737 (O_737,N_4818,N_4896);
and UO_738 (O_738,N_4960,N_4905);
nor UO_739 (O_739,N_4852,N_4987);
nor UO_740 (O_740,N_4970,N_4822);
nor UO_741 (O_741,N_4857,N_4885);
nor UO_742 (O_742,N_4837,N_4855);
or UO_743 (O_743,N_4909,N_4884);
and UO_744 (O_744,N_4957,N_4810);
or UO_745 (O_745,N_4802,N_4984);
and UO_746 (O_746,N_4997,N_4893);
and UO_747 (O_747,N_4913,N_4981);
nor UO_748 (O_748,N_4935,N_4803);
or UO_749 (O_749,N_4980,N_4858);
or UO_750 (O_750,N_4928,N_4950);
nand UO_751 (O_751,N_4979,N_4887);
and UO_752 (O_752,N_4803,N_4808);
and UO_753 (O_753,N_4818,N_4828);
and UO_754 (O_754,N_4905,N_4926);
or UO_755 (O_755,N_4882,N_4977);
and UO_756 (O_756,N_4815,N_4810);
nand UO_757 (O_757,N_4869,N_4880);
or UO_758 (O_758,N_4917,N_4968);
or UO_759 (O_759,N_4965,N_4916);
and UO_760 (O_760,N_4947,N_4960);
nor UO_761 (O_761,N_4898,N_4819);
and UO_762 (O_762,N_4928,N_4966);
nor UO_763 (O_763,N_4825,N_4945);
nor UO_764 (O_764,N_4817,N_4823);
or UO_765 (O_765,N_4840,N_4889);
and UO_766 (O_766,N_4877,N_4923);
xor UO_767 (O_767,N_4865,N_4983);
nand UO_768 (O_768,N_4836,N_4801);
nand UO_769 (O_769,N_4981,N_4972);
nor UO_770 (O_770,N_4853,N_4840);
nand UO_771 (O_771,N_4955,N_4985);
and UO_772 (O_772,N_4924,N_4887);
nor UO_773 (O_773,N_4859,N_4811);
or UO_774 (O_774,N_4904,N_4848);
or UO_775 (O_775,N_4820,N_4878);
and UO_776 (O_776,N_4892,N_4810);
nor UO_777 (O_777,N_4805,N_4842);
nor UO_778 (O_778,N_4953,N_4978);
nor UO_779 (O_779,N_4865,N_4853);
and UO_780 (O_780,N_4916,N_4831);
nand UO_781 (O_781,N_4807,N_4892);
nor UO_782 (O_782,N_4819,N_4888);
and UO_783 (O_783,N_4892,N_4817);
nand UO_784 (O_784,N_4975,N_4938);
nor UO_785 (O_785,N_4801,N_4981);
nor UO_786 (O_786,N_4917,N_4804);
nand UO_787 (O_787,N_4907,N_4947);
nand UO_788 (O_788,N_4876,N_4935);
and UO_789 (O_789,N_4888,N_4863);
nor UO_790 (O_790,N_4844,N_4866);
nand UO_791 (O_791,N_4937,N_4945);
nand UO_792 (O_792,N_4976,N_4980);
nor UO_793 (O_793,N_4980,N_4817);
and UO_794 (O_794,N_4822,N_4831);
and UO_795 (O_795,N_4986,N_4907);
or UO_796 (O_796,N_4962,N_4818);
nand UO_797 (O_797,N_4969,N_4896);
or UO_798 (O_798,N_4905,N_4937);
and UO_799 (O_799,N_4841,N_4920);
nor UO_800 (O_800,N_4854,N_4840);
nand UO_801 (O_801,N_4834,N_4919);
or UO_802 (O_802,N_4922,N_4842);
and UO_803 (O_803,N_4936,N_4913);
and UO_804 (O_804,N_4959,N_4992);
xor UO_805 (O_805,N_4966,N_4913);
nand UO_806 (O_806,N_4955,N_4960);
or UO_807 (O_807,N_4943,N_4973);
or UO_808 (O_808,N_4840,N_4942);
nor UO_809 (O_809,N_4898,N_4815);
nand UO_810 (O_810,N_4859,N_4932);
nand UO_811 (O_811,N_4812,N_4914);
and UO_812 (O_812,N_4868,N_4983);
nand UO_813 (O_813,N_4848,N_4817);
and UO_814 (O_814,N_4886,N_4973);
nor UO_815 (O_815,N_4804,N_4820);
nor UO_816 (O_816,N_4845,N_4819);
and UO_817 (O_817,N_4958,N_4853);
and UO_818 (O_818,N_4972,N_4954);
or UO_819 (O_819,N_4846,N_4941);
nor UO_820 (O_820,N_4889,N_4967);
or UO_821 (O_821,N_4888,N_4932);
and UO_822 (O_822,N_4832,N_4829);
and UO_823 (O_823,N_4931,N_4850);
nor UO_824 (O_824,N_4985,N_4998);
or UO_825 (O_825,N_4934,N_4999);
nand UO_826 (O_826,N_4896,N_4971);
or UO_827 (O_827,N_4856,N_4861);
nand UO_828 (O_828,N_4827,N_4855);
or UO_829 (O_829,N_4967,N_4822);
nand UO_830 (O_830,N_4889,N_4810);
nor UO_831 (O_831,N_4918,N_4942);
or UO_832 (O_832,N_4963,N_4992);
or UO_833 (O_833,N_4825,N_4960);
nand UO_834 (O_834,N_4869,N_4906);
and UO_835 (O_835,N_4929,N_4830);
nor UO_836 (O_836,N_4853,N_4962);
nor UO_837 (O_837,N_4812,N_4907);
nand UO_838 (O_838,N_4865,N_4917);
and UO_839 (O_839,N_4805,N_4827);
nand UO_840 (O_840,N_4845,N_4922);
nand UO_841 (O_841,N_4880,N_4804);
nor UO_842 (O_842,N_4873,N_4864);
or UO_843 (O_843,N_4890,N_4985);
and UO_844 (O_844,N_4831,N_4860);
nor UO_845 (O_845,N_4936,N_4986);
or UO_846 (O_846,N_4959,N_4874);
nand UO_847 (O_847,N_4856,N_4866);
nor UO_848 (O_848,N_4823,N_4801);
nand UO_849 (O_849,N_4888,N_4893);
nand UO_850 (O_850,N_4801,N_4950);
and UO_851 (O_851,N_4870,N_4956);
or UO_852 (O_852,N_4832,N_4840);
or UO_853 (O_853,N_4892,N_4850);
nor UO_854 (O_854,N_4810,N_4935);
nor UO_855 (O_855,N_4855,N_4828);
and UO_856 (O_856,N_4895,N_4874);
nor UO_857 (O_857,N_4816,N_4960);
or UO_858 (O_858,N_4973,N_4846);
or UO_859 (O_859,N_4800,N_4915);
or UO_860 (O_860,N_4840,N_4811);
nand UO_861 (O_861,N_4964,N_4954);
nand UO_862 (O_862,N_4911,N_4877);
nand UO_863 (O_863,N_4871,N_4885);
nand UO_864 (O_864,N_4879,N_4926);
nand UO_865 (O_865,N_4874,N_4988);
nor UO_866 (O_866,N_4919,N_4842);
nand UO_867 (O_867,N_4999,N_4968);
and UO_868 (O_868,N_4963,N_4831);
and UO_869 (O_869,N_4859,N_4810);
nor UO_870 (O_870,N_4813,N_4923);
or UO_871 (O_871,N_4916,N_4927);
and UO_872 (O_872,N_4943,N_4920);
and UO_873 (O_873,N_4892,N_4993);
nand UO_874 (O_874,N_4800,N_4944);
or UO_875 (O_875,N_4886,N_4867);
nand UO_876 (O_876,N_4821,N_4853);
or UO_877 (O_877,N_4964,N_4860);
and UO_878 (O_878,N_4889,N_4821);
nand UO_879 (O_879,N_4861,N_4881);
or UO_880 (O_880,N_4837,N_4860);
and UO_881 (O_881,N_4982,N_4828);
or UO_882 (O_882,N_4818,N_4832);
xnor UO_883 (O_883,N_4968,N_4995);
xor UO_884 (O_884,N_4843,N_4828);
or UO_885 (O_885,N_4817,N_4978);
and UO_886 (O_886,N_4891,N_4800);
nor UO_887 (O_887,N_4959,N_4900);
and UO_888 (O_888,N_4997,N_4886);
nor UO_889 (O_889,N_4807,N_4988);
or UO_890 (O_890,N_4889,N_4905);
nand UO_891 (O_891,N_4891,N_4870);
and UO_892 (O_892,N_4866,N_4961);
xnor UO_893 (O_893,N_4973,N_4832);
nand UO_894 (O_894,N_4808,N_4912);
or UO_895 (O_895,N_4934,N_4928);
nor UO_896 (O_896,N_4916,N_4901);
or UO_897 (O_897,N_4844,N_4888);
nand UO_898 (O_898,N_4932,N_4946);
nor UO_899 (O_899,N_4924,N_4871);
or UO_900 (O_900,N_4866,N_4956);
nor UO_901 (O_901,N_4837,N_4877);
nand UO_902 (O_902,N_4820,N_4941);
nor UO_903 (O_903,N_4805,N_4861);
and UO_904 (O_904,N_4814,N_4900);
and UO_905 (O_905,N_4867,N_4895);
nand UO_906 (O_906,N_4839,N_4832);
nor UO_907 (O_907,N_4982,N_4831);
nand UO_908 (O_908,N_4935,N_4934);
and UO_909 (O_909,N_4884,N_4885);
nor UO_910 (O_910,N_4844,N_4855);
nand UO_911 (O_911,N_4935,N_4843);
or UO_912 (O_912,N_4944,N_4902);
xnor UO_913 (O_913,N_4817,N_4846);
or UO_914 (O_914,N_4948,N_4971);
and UO_915 (O_915,N_4925,N_4916);
and UO_916 (O_916,N_4803,N_4960);
nand UO_917 (O_917,N_4849,N_4847);
nor UO_918 (O_918,N_4938,N_4894);
and UO_919 (O_919,N_4978,N_4804);
and UO_920 (O_920,N_4945,N_4894);
and UO_921 (O_921,N_4937,N_4864);
nor UO_922 (O_922,N_4915,N_4935);
or UO_923 (O_923,N_4831,N_4824);
nand UO_924 (O_924,N_4907,N_4917);
and UO_925 (O_925,N_4960,N_4850);
nand UO_926 (O_926,N_4941,N_4975);
or UO_927 (O_927,N_4865,N_4887);
nand UO_928 (O_928,N_4930,N_4883);
or UO_929 (O_929,N_4977,N_4954);
nand UO_930 (O_930,N_4907,N_4994);
nor UO_931 (O_931,N_4828,N_4852);
or UO_932 (O_932,N_4962,N_4972);
and UO_933 (O_933,N_4930,N_4937);
nand UO_934 (O_934,N_4929,N_4915);
nor UO_935 (O_935,N_4950,N_4970);
or UO_936 (O_936,N_4960,N_4922);
nor UO_937 (O_937,N_4852,N_4810);
nor UO_938 (O_938,N_4951,N_4991);
nor UO_939 (O_939,N_4926,N_4890);
and UO_940 (O_940,N_4846,N_4922);
nor UO_941 (O_941,N_4828,N_4804);
nor UO_942 (O_942,N_4986,N_4843);
or UO_943 (O_943,N_4831,N_4933);
and UO_944 (O_944,N_4885,N_4830);
nor UO_945 (O_945,N_4855,N_4975);
or UO_946 (O_946,N_4996,N_4813);
nor UO_947 (O_947,N_4971,N_4920);
nor UO_948 (O_948,N_4843,N_4878);
or UO_949 (O_949,N_4860,N_4986);
or UO_950 (O_950,N_4951,N_4965);
or UO_951 (O_951,N_4975,N_4800);
or UO_952 (O_952,N_4910,N_4897);
or UO_953 (O_953,N_4839,N_4972);
nand UO_954 (O_954,N_4884,N_4904);
nand UO_955 (O_955,N_4988,N_4949);
and UO_956 (O_956,N_4938,N_4814);
or UO_957 (O_957,N_4974,N_4951);
nand UO_958 (O_958,N_4865,N_4812);
and UO_959 (O_959,N_4916,N_4986);
and UO_960 (O_960,N_4901,N_4921);
and UO_961 (O_961,N_4885,N_4950);
or UO_962 (O_962,N_4940,N_4966);
and UO_963 (O_963,N_4974,N_4857);
or UO_964 (O_964,N_4980,N_4981);
nand UO_965 (O_965,N_4808,N_4816);
nand UO_966 (O_966,N_4874,N_4926);
nor UO_967 (O_967,N_4907,N_4853);
and UO_968 (O_968,N_4948,N_4981);
nand UO_969 (O_969,N_4978,N_4863);
and UO_970 (O_970,N_4847,N_4889);
and UO_971 (O_971,N_4804,N_4913);
and UO_972 (O_972,N_4857,N_4928);
nor UO_973 (O_973,N_4989,N_4948);
or UO_974 (O_974,N_4800,N_4918);
and UO_975 (O_975,N_4980,N_4893);
nor UO_976 (O_976,N_4916,N_4864);
nand UO_977 (O_977,N_4821,N_4874);
or UO_978 (O_978,N_4839,N_4814);
nand UO_979 (O_979,N_4998,N_4928);
or UO_980 (O_980,N_4959,N_4981);
or UO_981 (O_981,N_4915,N_4873);
or UO_982 (O_982,N_4883,N_4900);
nor UO_983 (O_983,N_4941,N_4909);
or UO_984 (O_984,N_4856,N_4867);
nor UO_985 (O_985,N_4817,N_4911);
and UO_986 (O_986,N_4874,N_4972);
or UO_987 (O_987,N_4886,N_4803);
and UO_988 (O_988,N_4880,N_4874);
and UO_989 (O_989,N_4939,N_4887);
or UO_990 (O_990,N_4901,N_4995);
nor UO_991 (O_991,N_4861,N_4849);
nor UO_992 (O_992,N_4832,N_4977);
or UO_993 (O_993,N_4896,N_4845);
and UO_994 (O_994,N_4930,N_4936);
and UO_995 (O_995,N_4964,N_4846);
and UO_996 (O_996,N_4932,N_4827);
and UO_997 (O_997,N_4859,N_4890);
or UO_998 (O_998,N_4997,N_4887);
or UO_999 (O_999,N_4812,N_4845);
endmodule