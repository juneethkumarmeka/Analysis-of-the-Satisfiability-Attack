module basic_2500_25000_3000_40_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_619,In_1970);
nand U1 (N_1,In_1313,In_896);
nor U2 (N_2,In_2252,In_1965);
nand U3 (N_3,In_2471,In_197);
or U4 (N_4,In_2305,In_26);
or U5 (N_5,In_2018,In_106);
or U6 (N_6,In_480,In_53);
or U7 (N_7,In_125,In_1726);
nand U8 (N_8,In_55,In_229);
nor U9 (N_9,In_782,In_18);
or U10 (N_10,In_16,In_117);
nor U11 (N_11,In_189,In_2247);
and U12 (N_12,In_1865,In_736);
or U13 (N_13,In_1287,In_2191);
nor U14 (N_14,In_1729,In_533);
xor U15 (N_15,In_1648,In_2007);
xnor U16 (N_16,In_439,In_1988);
xnor U17 (N_17,In_1170,In_1282);
nor U18 (N_18,In_2364,In_52);
or U19 (N_19,In_2081,In_295);
nand U20 (N_20,In_1624,In_573);
nand U21 (N_21,In_1740,In_1336);
xor U22 (N_22,In_37,In_2053);
and U23 (N_23,In_1422,In_1542);
nand U24 (N_24,In_705,In_1375);
nor U25 (N_25,In_742,In_2172);
nand U26 (N_26,In_1208,In_458);
or U27 (N_27,In_522,In_321);
and U28 (N_28,In_2192,In_1436);
nand U29 (N_29,In_2254,In_1310);
nand U30 (N_30,In_2112,In_1901);
and U31 (N_31,In_730,In_889);
xor U32 (N_32,In_2258,In_922);
or U33 (N_33,In_1519,In_387);
or U34 (N_34,In_1420,In_1312);
or U35 (N_35,In_729,In_1296);
or U36 (N_36,In_245,In_30);
or U37 (N_37,In_1508,In_1917);
nor U38 (N_38,In_2203,In_1891);
nor U39 (N_39,In_1687,In_2242);
xnor U40 (N_40,In_1702,In_1378);
or U41 (N_41,In_1189,In_1290);
nand U42 (N_42,In_1720,In_2066);
nand U43 (N_43,In_1869,In_301);
or U44 (N_44,In_440,In_98);
or U45 (N_45,In_652,In_1589);
nor U46 (N_46,In_2197,In_2331);
or U47 (N_47,In_720,In_559);
xnor U48 (N_48,In_989,In_317);
xnor U49 (N_49,In_792,In_2131);
xnor U50 (N_50,In_1110,In_1320);
nor U51 (N_51,In_94,In_1139);
nor U52 (N_52,In_1164,In_1305);
and U53 (N_53,In_2162,In_1458);
nand U54 (N_54,In_908,In_1428);
xor U55 (N_55,In_2399,In_395);
nand U56 (N_56,In_929,In_2138);
nand U57 (N_57,In_745,In_1265);
xor U58 (N_58,In_1475,In_2015);
and U59 (N_59,In_1331,In_1317);
nor U60 (N_60,In_860,In_1625);
and U61 (N_61,In_102,In_1196);
xnor U62 (N_62,In_632,In_2363);
xnor U63 (N_63,In_2375,In_886);
or U64 (N_64,In_1578,In_1506);
or U65 (N_65,In_1468,In_497);
and U66 (N_66,In_988,In_917);
or U67 (N_67,In_1714,In_1486);
nand U68 (N_68,In_99,In_1772);
xnor U69 (N_69,In_269,In_1738);
nor U70 (N_70,In_529,In_778);
or U71 (N_71,In_369,In_916);
xnor U72 (N_72,In_2054,In_796);
nor U73 (N_73,In_1845,In_793);
xor U74 (N_74,In_262,In_1062);
or U75 (N_75,In_224,In_912);
nand U76 (N_76,In_2347,In_1018);
nand U77 (N_77,In_2251,In_1138);
or U78 (N_78,In_856,In_1014);
xor U79 (N_79,In_2064,In_773);
nand U80 (N_80,In_888,In_177);
xor U81 (N_81,In_2256,In_338);
nand U82 (N_82,In_952,In_334);
xor U83 (N_83,In_2308,In_1258);
or U84 (N_84,In_1431,In_453);
and U85 (N_85,In_2359,In_893);
xor U86 (N_86,In_1850,In_2445);
xor U87 (N_87,In_1048,In_288);
nor U88 (N_88,In_830,In_325);
nand U89 (N_89,In_1511,In_79);
nand U90 (N_90,In_928,In_2259);
and U91 (N_91,In_204,In_1715);
xnor U92 (N_92,In_1273,In_1924);
and U93 (N_93,In_1448,In_1543);
xor U94 (N_94,In_1728,In_2133);
nor U95 (N_95,In_1945,In_633);
nand U96 (N_96,In_1716,In_1179);
xor U97 (N_97,In_1408,In_375);
and U98 (N_98,In_123,In_394);
xor U99 (N_99,In_2052,In_384);
xnor U100 (N_100,In_2354,In_2026);
nor U101 (N_101,In_2279,In_1377);
or U102 (N_102,In_920,In_1992);
nand U103 (N_103,In_378,In_2187);
xnor U104 (N_104,In_948,In_2361);
nand U105 (N_105,In_1597,In_1045);
nor U106 (N_106,In_1700,In_216);
xor U107 (N_107,In_2050,In_2451);
and U108 (N_108,In_2250,In_690);
nand U109 (N_109,In_227,In_1609);
xnor U110 (N_110,In_521,In_236);
or U111 (N_111,In_157,In_1193);
xnor U112 (N_112,In_305,In_196);
and U113 (N_113,In_2379,In_1564);
nor U114 (N_114,In_1149,In_193);
or U115 (N_115,In_2412,In_1175);
xnor U116 (N_116,In_1509,In_469);
nand U117 (N_117,In_1710,In_502);
nor U118 (N_118,In_1278,In_1293);
and U119 (N_119,In_605,In_273);
and U120 (N_120,In_1822,In_1166);
or U121 (N_121,In_1051,In_1387);
and U122 (N_122,In_868,In_1315);
nor U123 (N_123,In_76,In_564);
or U124 (N_124,In_1060,In_1148);
and U125 (N_125,In_2395,In_1569);
and U126 (N_126,In_1212,In_242);
xnor U127 (N_127,In_462,In_2088);
nand U128 (N_128,In_501,In_776);
xnor U129 (N_129,In_65,In_804);
nor U130 (N_130,In_1993,In_281);
nor U131 (N_131,In_1309,In_1701);
xnor U132 (N_132,In_1111,In_133);
xor U133 (N_133,In_1692,In_1492);
nor U134 (N_134,In_560,In_1931);
nor U135 (N_135,In_302,In_1064);
xor U136 (N_136,In_1560,In_306);
xor U137 (N_137,In_2057,In_1639);
nor U138 (N_138,In_142,In_419);
nand U139 (N_139,In_1288,In_1386);
or U140 (N_140,In_698,In_1214);
or U141 (N_141,In_983,In_2420);
xor U142 (N_142,In_202,In_822);
nor U143 (N_143,In_1198,In_2327);
xor U144 (N_144,In_1673,In_155);
nor U145 (N_145,In_1178,In_1882);
nor U146 (N_146,In_261,In_1391);
or U147 (N_147,In_2045,In_2294);
and U148 (N_148,In_554,In_1144);
nor U149 (N_149,In_1626,In_1926);
xnor U150 (N_150,In_19,In_1426);
xnor U151 (N_151,In_1024,In_1071);
xnor U152 (N_152,In_1430,In_162);
nor U153 (N_153,In_757,In_1435);
nor U154 (N_154,In_2167,In_1142);
and U155 (N_155,In_320,In_2457);
nor U156 (N_156,In_691,In_1215);
nand U157 (N_157,In_862,In_2313);
nor U158 (N_158,In_432,In_256);
nor U159 (N_159,In_641,In_1722);
and U160 (N_160,In_2013,In_672);
nand U161 (N_161,In_70,In_1327);
xor U162 (N_162,In_28,In_938);
nor U163 (N_163,In_2468,In_1656);
nand U164 (N_164,In_1608,In_2208);
xnor U165 (N_165,In_1104,In_2207);
xnor U166 (N_166,In_1368,In_2366);
and U167 (N_167,In_175,In_96);
or U168 (N_168,In_1335,In_354);
nand U169 (N_169,In_2410,In_1030);
and U170 (N_170,In_2315,In_885);
nand U171 (N_171,In_2290,In_1217);
and U172 (N_172,In_2209,In_971);
nor U173 (N_173,In_1711,In_1634);
nor U174 (N_174,In_991,In_1128);
nor U175 (N_175,In_1994,In_1016);
and U176 (N_176,In_324,In_170);
or U177 (N_177,In_1848,In_1115);
nand U178 (N_178,In_215,In_1944);
xnor U179 (N_179,In_591,In_158);
nand U180 (N_180,In_1963,In_358);
or U181 (N_181,In_1957,In_1971);
or U182 (N_182,In_1763,In_476);
or U183 (N_183,In_944,In_60);
nor U184 (N_184,In_2150,In_1319);
or U185 (N_185,In_639,In_2286);
nand U186 (N_186,In_391,In_1878);
or U187 (N_187,In_1499,In_528);
nand U188 (N_188,In_1363,In_1080);
and U189 (N_189,In_2337,In_1995);
nor U190 (N_190,In_1053,In_2266);
xor U191 (N_191,In_762,In_1253);
nor U192 (N_192,In_1539,In_2389);
nand U193 (N_193,In_819,In_2429);
xnor U194 (N_194,In_2486,In_577);
nand U195 (N_195,In_699,In_1675);
xor U196 (N_196,In_1640,In_114);
nand U197 (N_197,In_2097,In_1579);
and U198 (N_198,In_1690,In_2326);
and U199 (N_199,In_704,In_1165);
nand U200 (N_200,In_1923,In_1513);
or U201 (N_201,In_630,In_2368);
xor U202 (N_202,In_1998,In_2070);
nor U203 (N_203,In_17,In_2411);
and U204 (N_204,In_2293,In_602);
and U205 (N_205,In_919,In_1834);
or U206 (N_206,In_2019,In_167);
or U207 (N_207,In_1122,In_894);
or U208 (N_208,In_2204,In_146);
nand U209 (N_209,In_601,In_209);
xor U210 (N_210,In_1304,In_2426);
and U211 (N_211,In_111,In_1987);
nand U212 (N_212,In_83,In_2303);
xor U213 (N_213,In_1061,In_1935);
xnor U214 (N_214,In_775,In_1999);
and U215 (N_215,In_2194,In_688);
nand U216 (N_216,In_1552,In_1762);
xor U217 (N_217,In_1875,In_2212);
nand U218 (N_218,In_459,In_596);
nor U219 (N_219,In_1480,In_1405);
nand U220 (N_220,In_427,In_1314);
nand U221 (N_221,In_1825,In_186);
or U222 (N_222,In_1081,In_1440);
nand U223 (N_223,In_1678,In_1223);
xor U224 (N_224,In_1330,In_41);
or U225 (N_225,In_292,In_315);
xnor U226 (N_226,In_1200,In_1655);
nand U227 (N_227,In_1580,In_654);
nand U228 (N_228,In_192,In_1880);
or U229 (N_229,In_2033,In_612);
nand U230 (N_230,In_1514,In_435);
nand U231 (N_231,In_808,In_707);
xor U232 (N_232,In_486,In_1830);
xnor U233 (N_233,In_1551,In_2367);
xor U234 (N_234,In_90,In_1867);
nand U235 (N_235,In_802,In_814);
xnor U236 (N_236,In_748,In_2008);
nor U237 (N_237,In_156,In_335);
nor U238 (N_238,In_2236,In_1154);
and U239 (N_239,In_198,In_2283);
or U240 (N_240,In_608,In_403);
and U241 (N_241,In_1835,In_932);
nand U242 (N_242,In_1783,In_1745);
or U243 (N_243,In_1750,In_2029);
or U244 (N_244,In_1191,In_323);
nand U245 (N_245,In_179,In_1614);
or U246 (N_246,In_1739,In_765);
nor U247 (N_247,In_225,In_285);
nand U248 (N_248,In_210,In_420);
and U249 (N_249,In_1503,In_1941);
xnor U250 (N_250,In_2160,In_598);
or U251 (N_251,In_1786,In_801);
nand U252 (N_252,In_2484,In_1916);
nor U253 (N_253,In_407,In_2092);
nand U254 (N_254,In_1811,In_86);
or U255 (N_255,In_1870,In_904);
nand U256 (N_256,In_869,In_247);
xnor U257 (N_257,In_405,In_1973);
or U258 (N_258,In_2069,In_950);
nor U259 (N_259,In_2168,In_959);
xor U260 (N_260,In_2496,In_1112);
xor U261 (N_261,In_723,In_1156);
or U262 (N_262,In_2022,In_680);
nor U263 (N_263,In_1488,In_2023);
and U264 (N_264,In_2104,In_1123);
or U265 (N_265,In_2086,In_2270);
or U266 (N_266,In_265,In_1004);
nor U267 (N_267,In_337,In_2431);
or U268 (N_268,In_1407,In_2017);
xor U269 (N_269,In_2102,In_2415);
or U270 (N_270,In_322,In_2287);
nand U271 (N_271,In_648,In_1765);
xnor U272 (N_272,In_289,In_1982);
nor U273 (N_273,In_714,In_1298);
nor U274 (N_274,In_582,In_393);
and U275 (N_275,In_2413,In_367);
nor U276 (N_276,In_2320,In_2295);
nand U277 (N_277,In_362,In_2149);
xnor U278 (N_278,In_546,In_1383);
or U279 (N_279,In_905,In_1694);
or U280 (N_280,In_91,In_1339);
nand U281 (N_281,In_2460,In_424);
nand U282 (N_282,In_219,In_506);
or U283 (N_283,In_172,In_1977);
or U284 (N_284,In_1810,In_31);
or U285 (N_285,In_2436,In_2271);
nor U286 (N_286,In_61,In_1211);
or U287 (N_287,In_2483,In_1704);
nor U288 (N_288,In_927,In_275);
or U289 (N_289,In_768,In_532);
and U290 (N_290,In_1360,In_1927);
or U291 (N_291,In_1418,In_1252);
or U292 (N_292,In_212,In_1529);
and U293 (N_293,In_264,In_949);
or U294 (N_294,In_34,In_1180);
and U295 (N_295,In_626,In_2463);
xnor U296 (N_296,In_622,In_597);
nor U297 (N_297,In_344,In_1902);
and U298 (N_298,In_1686,In_863);
or U299 (N_299,In_2227,In_653);
and U300 (N_300,In_1844,In_260);
or U301 (N_301,In_1549,In_2198);
and U302 (N_302,In_1346,In_383);
nor U303 (N_303,In_492,In_1113);
or U304 (N_304,In_2307,In_1662);
nand U305 (N_305,In_1533,In_1683);
nand U306 (N_306,In_1647,In_2079);
nand U307 (N_307,In_280,In_1344);
nor U308 (N_308,In_973,In_1752);
and U309 (N_309,In_2152,In_112);
nor U310 (N_310,In_518,In_738);
and U311 (N_311,In_1607,In_2459);
or U312 (N_312,In_2322,In_414);
and U313 (N_313,In_2180,In_2105);
or U314 (N_314,In_716,In_1501);
xor U315 (N_315,In_2346,In_482);
nor U316 (N_316,In_1836,In_625);
or U317 (N_317,In_2311,In_956);
and U318 (N_318,In_1755,In_2228);
nand U319 (N_319,In_2369,In_2492);
xnor U320 (N_320,In_444,In_1434);
xor U321 (N_321,In_1137,In_556);
xor U322 (N_322,In_513,In_1190);
or U323 (N_323,In_254,In_1197);
xnor U324 (N_324,In_24,In_1909);
and U325 (N_325,In_872,In_1698);
nand U326 (N_326,In_2155,In_116);
xor U327 (N_327,In_696,In_221);
xnor U328 (N_328,In_1133,In_1131);
xnor U329 (N_329,In_1900,In_2456);
xnor U330 (N_330,In_381,In_1797);
or U331 (N_331,In_1620,In_1753);
nand U332 (N_332,In_1600,In_734);
or U333 (N_333,In_1406,In_1233);
nand U334 (N_334,In_1912,In_1976);
or U335 (N_335,In_2365,In_2119);
xor U336 (N_336,In_1685,In_517);
and U337 (N_337,In_1660,In_426);
and U338 (N_338,In_2243,In_2376);
xnor U339 (N_339,In_2268,In_962);
and U340 (N_340,In_1877,In_2239);
xnor U341 (N_341,In_2284,In_2325);
or U342 (N_342,In_416,In_794);
and U343 (N_343,In_1325,In_709);
nor U344 (N_344,In_2473,In_972);
nand U345 (N_345,In_1140,In_408);
and U346 (N_346,In_1059,In_771);
and U347 (N_347,In_744,In_485);
nand U348 (N_348,In_311,In_566);
xor U349 (N_349,In_279,In_543);
and U350 (N_350,In_1228,In_182);
and U351 (N_351,In_11,In_1754);
nand U352 (N_352,In_1372,In_2164);
nor U353 (N_353,In_1838,In_758);
nand U354 (N_354,In_2126,In_342);
xor U355 (N_355,In_964,In_2186);
or U356 (N_356,In_1617,In_2355);
nand U357 (N_357,In_1452,In_569);
nor U358 (N_358,In_866,In_900);
nor U359 (N_359,In_2257,In_494);
nand U360 (N_360,In_879,In_694);
nor U361 (N_361,In_1021,In_537);
nand U362 (N_362,In_92,In_1118);
nor U363 (N_363,In_578,In_1297);
nand U364 (N_364,In_1362,In_788);
or U365 (N_365,In_356,In_1771);
xor U366 (N_366,In_755,In_1540);
and U367 (N_367,In_1856,In_2391);
or U368 (N_368,In_2272,In_2358);
and U369 (N_369,In_882,In_516);
nand U370 (N_370,In_1000,In_1896);
xor U371 (N_371,In_2446,In_1795);
nor U372 (N_372,In_884,In_1151);
or U373 (N_373,In_1359,In_1760);
and U374 (N_374,In_609,In_1404);
nor U375 (N_375,In_2061,In_1099);
xor U376 (N_376,In_2114,In_1855);
nor U377 (N_377,In_113,In_800);
nand U378 (N_378,In_735,In_1558);
and U379 (N_379,In_1351,In_438);
or U380 (N_380,In_610,In_726);
nor U381 (N_381,In_1496,In_1324);
and U382 (N_382,In_456,In_719);
xnor U383 (N_383,In_1251,In_2195);
or U384 (N_384,In_891,In_535);
nand U385 (N_385,In_1459,In_1152);
xor U386 (N_386,In_2374,In_1277);
nand U387 (N_387,In_918,In_2224);
xor U388 (N_388,In_2036,In_368);
and U389 (N_389,In_218,In_163);
and U390 (N_390,In_1644,In_1813);
and U391 (N_391,In_78,In_550);
and U392 (N_392,In_1669,In_906);
nand U393 (N_393,In_923,In_2384);
xor U394 (N_394,In_861,In_763);
nand U395 (N_395,In_1604,In_2184);
nand U396 (N_396,In_2465,In_1316);
xnor U397 (N_397,In_1990,In_1065);
and U398 (N_398,In_95,In_780);
or U399 (N_399,In_1329,In_1466);
nor U400 (N_400,In_2439,In_833);
nor U401 (N_401,In_2230,In_2106);
nand U402 (N_402,In_865,In_2078);
nor U403 (N_403,In_1559,In_2166);
and U404 (N_404,In_1311,In_851);
and U405 (N_405,In_1078,In_1457);
or U406 (N_406,In_1244,In_722);
and U407 (N_407,In_1553,In_541);
xnor U408 (N_408,In_1802,In_353);
nand U409 (N_409,In_2060,In_134);
nand U410 (N_410,In_1735,In_713);
or U411 (N_411,In_1649,In_1507);
and U412 (N_412,In_536,In_1664);
nor U413 (N_413,In_2144,In_881);
or U414 (N_414,In_66,In_2350);
xor U415 (N_415,In_1479,In_933);
nand U416 (N_416,In_1780,In_40);
xor U417 (N_417,In_996,In_1725);
or U418 (N_418,In_1474,In_2083);
nand U419 (N_419,In_1518,In_1670);
xor U420 (N_420,In_466,In_2056);
xor U421 (N_421,In_1415,In_1618);
or U422 (N_422,In_422,In_168);
and U423 (N_423,In_2109,In_1095);
nand U424 (N_424,In_319,In_231);
xor U425 (N_425,In_296,In_1732);
nor U426 (N_426,In_309,In_2099);
nand U427 (N_427,In_2025,In_1733);
and U428 (N_428,In_446,In_498);
or U429 (N_429,In_1032,In_1932);
or U430 (N_430,In_33,In_1576);
or U431 (N_431,In_2244,In_2235);
nor U432 (N_432,In_1385,In_697);
nor U433 (N_433,In_1605,In_1642);
and U434 (N_434,In_1570,In_1220);
xor U435 (N_435,In_2034,In_1271);
or U436 (N_436,In_141,In_2348);
nand U437 (N_437,In_825,In_984);
and U438 (N_438,In_2454,In_1953);
xor U439 (N_439,In_561,In_2043);
or U440 (N_440,In_662,In_2222);
nor U441 (N_441,In_1283,In_1495);
nor U442 (N_442,In_656,In_415);
nor U443 (N_443,In_943,In_600);
nand U444 (N_444,In_207,In_1601);
and U445 (N_445,In_777,In_2014);
xor U446 (N_446,In_208,In_2177);
xor U447 (N_447,In_149,In_1933);
xnor U448 (N_448,In_428,In_593);
xnor U449 (N_449,In_781,In_1731);
xor U450 (N_450,In_1427,In_140);
and U451 (N_451,In_1695,In_1424);
and U452 (N_452,In_2206,In_1043);
and U453 (N_453,In_1490,In_1381);
nor U454 (N_454,In_1879,In_1120);
nor U455 (N_455,In_1467,In_1086);
nand U456 (N_456,In_2111,In_658);
xor U457 (N_457,In_431,In_239);
nand U458 (N_458,In_411,In_1785);
nand U459 (N_459,In_774,In_437);
xor U460 (N_460,In_2418,In_1585);
and U461 (N_461,In_1260,In_1746);
and U462 (N_462,In_805,In_646);
xnor U463 (N_463,In_503,In_417);
or U464 (N_464,In_2010,In_1814);
nand U465 (N_465,In_1056,In_1221);
nor U466 (N_466,In_687,In_2202);
xnor U467 (N_467,In_510,In_1592);
or U468 (N_468,In_1744,In_2096);
nand U469 (N_469,In_9,In_1846);
or U470 (N_470,In_749,In_1801);
nand U471 (N_471,In_404,In_1102);
nor U472 (N_472,In_2127,In_1161);
nand U473 (N_473,In_940,In_1937);
nand U474 (N_474,In_1243,In_1055);
or U475 (N_475,In_636,In_756);
xnor U476 (N_476,In_1764,In_1799);
and U477 (N_477,In_519,In_1380);
or U478 (N_478,In_2245,In_668);
and U479 (N_479,In_1135,In_443);
nand U480 (N_480,In_139,In_448);
or U481 (N_481,In_1526,In_43);
nand U482 (N_482,In_2498,In_2107);
nor U483 (N_483,In_57,In_1679);
nor U484 (N_484,In_511,In_1920);
nor U485 (N_485,In_447,In_545);
nor U486 (N_486,In_1124,In_1779);
nor U487 (N_487,In_1275,In_2046);
and U488 (N_488,In_2332,In_1535);
and U489 (N_489,In_766,In_1441);
nor U490 (N_490,In_1862,In_361);
xor U491 (N_491,In_2122,In_1790);
or U492 (N_492,In_1972,In_1007);
or U493 (N_493,In_1632,In_2118);
nor U494 (N_494,In_790,In_1237);
nand U495 (N_495,In_1623,In_2282);
and U496 (N_496,In_421,In_824);
or U497 (N_497,In_1079,In_1603);
xor U498 (N_498,In_1584,In_1172);
nand U499 (N_499,In_883,In_1129);
and U500 (N_500,In_1348,In_921);
and U501 (N_501,In_1054,In_1839);
nand U502 (N_502,In_784,In_1465);
or U503 (N_503,In_620,In_1910);
and U504 (N_504,In_230,In_213);
xnor U505 (N_505,In_910,In_2216);
xor U506 (N_506,In_1538,In_514);
xor U507 (N_507,In_1411,In_2442);
nand U508 (N_508,In_2255,In_753);
nand U509 (N_509,In_1593,In_2467);
nor U510 (N_510,In_1853,In_2146);
nor U511 (N_511,In_308,In_667);
nand U512 (N_512,In_77,In_71);
nor U513 (N_513,In_2425,In_1682);
nand U514 (N_514,In_1003,In_1697);
nor U515 (N_515,In_2285,In_1946);
nand U516 (N_516,In_942,In_235);
nand U517 (N_517,In_349,In_496);
nor U518 (N_518,In_1826,In_702);
nand U519 (N_519,In_246,In_1807);
nor U520 (N_520,In_2440,In_700);
and U521 (N_521,In_852,In_1069);
nand U522 (N_522,In_38,In_2499);
nor U523 (N_523,In_1712,In_1017);
and U524 (N_524,In_746,In_1);
xnor U525 (N_525,In_160,In_1192);
nor U526 (N_526,In_604,In_840);
or U527 (N_527,In_2020,In_2485);
nor U528 (N_528,In_1703,In_1087);
xor U529 (N_529,In_634,In_552);
xor U530 (N_530,In_2240,In_191);
xor U531 (N_531,In_467,In_1693);
xnor U532 (N_532,In_1093,In_1473);
nor U533 (N_533,In_346,In_731);
and U534 (N_534,In_188,In_1471);
xor U535 (N_535,In_1195,In_252);
or U536 (N_536,In_2382,In_1804);
xor U537 (N_537,In_594,In_835);
xor U538 (N_538,In_563,In_201);
and U539 (N_539,In_2419,In_1872);
or U540 (N_540,In_733,In_1899);
and U541 (N_541,In_1345,In_1938);
nand U542 (N_542,In_531,In_1724);
nand U543 (N_543,In_2136,In_64);
nor U544 (N_544,In_1888,In_1425);
nor U545 (N_545,In_621,In_176);
nor U546 (N_546,In_442,In_478);
nand U547 (N_547,In_2174,In_464);
xor U548 (N_548,In_1103,In_2404);
nor U549 (N_549,In_806,In_1903);
nand U550 (N_550,In_571,In_436);
and U551 (N_551,In_957,In_298);
or U552 (N_552,In_1402,In_1438);
and U553 (N_553,In_684,In_1416);
nand U554 (N_554,In_237,In_82);
xor U555 (N_555,In_572,In_1159);
xnor U556 (N_556,In_372,In_1340);
nor U557 (N_557,In_931,In_392);
nand U558 (N_558,In_1677,In_1485);
xor U559 (N_559,In_637,In_2085);
xnor U560 (N_560,In_1232,In_1985);
and U561 (N_561,In_1883,In_924);
or U562 (N_562,In_2360,In_1602);
xnor U563 (N_563,In_1766,In_452);
xnor U564 (N_564,In_222,In_1188);
nor U565 (N_565,In_907,In_1107);
xor U566 (N_566,In_895,In_351);
xor U567 (N_567,In_147,In_1510);
nand U568 (N_568,In_670,In_1796);
nor U569 (N_569,In_1761,In_2214);
nand U570 (N_570,In_187,In_715);
nand U571 (N_571,In_1672,In_2193);
or U572 (N_572,In_836,In_2217);
xnor U573 (N_573,In_1816,In_2477);
nand U574 (N_574,In_504,In_1394);
nand U575 (N_575,In_586,In_2458);
nor U576 (N_576,In_2414,In_607);
or U577 (N_577,In_2229,In_1979);
nor U578 (N_578,In_747,In_240);
and U579 (N_579,In_1652,In_2387);
nand U580 (N_580,In_708,In_1153);
nor U581 (N_581,In_2082,In_899);
or U582 (N_582,In_624,In_1858);
xnor U583 (N_583,In_1350,In_1136);
or U584 (N_584,In_2408,In_1996);
xor U585 (N_585,In_1171,In_1606);
nor U586 (N_586,In_1279,In_2095);
or U587 (N_587,In_651,In_2141);
nor U588 (N_588,In_1788,In_1011);
or U589 (N_589,In_1812,In_1125);
or U590 (N_590,In_551,In_1447);
and U591 (N_591,In_2336,In_303);
and U592 (N_592,In_903,In_2474);
and U593 (N_593,In_472,In_360);
xnor U594 (N_594,In_2487,In_2093);
xnor U595 (N_595,In_939,In_2495);
and U596 (N_596,In_803,In_993);
or U597 (N_597,In_1389,In_461);
or U598 (N_598,In_2356,In_846);
xnor U599 (N_599,In_2269,In_220);
nor U600 (N_600,In_1691,In_579);
nor U601 (N_601,In_2169,In_1074);
nor U602 (N_602,In_382,In_1815);
nor U603 (N_603,In_2005,In_2011);
and U604 (N_604,In_982,In_1583);
xnor U605 (N_605,In_2397,In_477);
nor U606 (N_606,In_2334,In_2394);
nor U607 (N_607,In_581,In_1379);
or U608 (N_608,In_479,In_1777);
nand U609 (N_609,In_359,In_1020);
nand U610 (N_610,In_1983,In_638);
nand U611 (N_611,In_2289,In_1259);
or U612 (N_612,In_1337,In_1637);
and U613 (N_613,In_93,In_2100);
nand U614 (N_614,In_875,In_1284);
and U615 (N_615,In_2120,In_1235);
or U616 (N_616,In_795,In_474);
nand U617 (N_617,In_331,In_1266);
nor U618 (N_618,In_363,In_1374);
and U619 (N_619,In_871,In_307);
xnor U620 (N_620,In_547,In_1638);
nand U621 (N_621,In_115,In_1307);
nor U622 (N_622,In_673,In_567);
nand U623 (N_623,In_925,In_583);
and U624 (N_624,In_399,In_2383);
and U625 (N_625,In_1759,N_457);
and U626 (N_626,In_1219,In_2300);
nand U627 (N_627,In_1949,N_494);
or U628 (N_628,In_374,In_418);
and U629 (N_629,In_1091,In_1049);
or U630 (N_630,N_93,In_2051);
nor U631 (N_631,In_2301,N_581);
nand U632 (N_632,N_169,N_595);
nand U633 (N_633,In_1322,In_542);
nand U634 (N_634,In_659,In_2433);
or U635 (N_635,N_372,In_1758);
nand U636 (N_636,N_73,N_299);
and U637 (N_637,N_621,N_541);
nor U638 (N_638,In_1906,N_405);
or U639 (N_639,In_1073,In_300);
or U640 (N_640,N_281,In_2464);
and U641 (N_641,In_1827,In_857);
nand U642 (N_642,In_44,In_500);
nand U643 (N_643,N_580,N_455);
and U644 (N_644,In_979,In_1823);
xor U645 (N_645,In_650,In_1803);
or U646 (N_646,In_2403,In_2044);
nand U647 (N_647,In_1914,In_647);
nor U648 (N_648,In_935,N_257);
xnor U649 (N_649,In_1462,In_1478);
xnor U650 (N_650,In_2161,In_629);
or U651 (N_651,In_834,In_505);
nand U652 (N_652,N_232,In_1419);
or U653 (N_653,N_212,N_310);
nor U654 (N_654,In_491,In_844);
and U655 (N_655,N_397,In_2328);
nor U656 (N_656,N_450,In_1022);
and U657 (N_657,In_1075,In_2241);
xnor U658 (N_658,In_108,In_874);
nor U659 (N_659,In_434,N_529);
xnor U660 (N_660,N_7,In_2153);
nand U661 (N_661,In_1203,In_35);
nor U662 (N_662,In_59,In_1876);
nand U663 (N_663,In_2281,N_521);
and U664 (N_664,In_1226,In_1554);
nor U665 (N_665,In_406,In_732);
and U666 (N_666,In_837,In_2273);
xor U667 (N_667,N_308,In_2199);
xnor U668 (N_668,In_58,N_249);
or U669 (N_669,N_138,In_2434);
nand U670 (N_670,In_1229,In_570);
and U671 (N_671,N_586,In_1532);
xnor U672 (N_672,N_479,In_409);
nand U673 (N_673,In_74,In_1082);
or U674 (N_674,N_606,In_997);
nand U675 (N_675,N_305,N_599);
nor U676 (N_676,N_272,In_1205);
or U677 (N_677,In_1676,In_1594);
xor U678 (N_678,In_1096,In_1665);
xnor U679 (N_679,N_129,N_221);
nand U680 (N_680,In_986,In_159);
or U681 (N_681,In_1098,N_164);
or U682 (N_682,In_1524,In_12);
nor U683 (N_683,In_2351,N_561);
or U684 (N_684,N_512,N_542);
and U685 (N_685,In_2028,In_283);
or U686 (N_686,In_2037,In_1413);
nand U687 (N_687,N_559,In_2306);
xnor U688 (N_688,In_1666,N_360);
nor U689 (N_689,In_199,N_188);
nor U690 (N_690,In_2154,N_395);
nand U691 (N_691,In_1143,In_1824);
or U692 (N_692,In_2089,N_190);
and U693 (N_693,In_1361,In_2263);
xor U694 (N_694,N_551,In_2323);
and U695 (N_695,In_1778,N_195);
nor U696 (N_696,N_403,N_300);
and U697 (N_697,In_873,In_1399);
xnor U698 (N_698,N_312,N_436);
nand U699 (N_699,N_474,In_345);
nor U700 (N_700,In_995,In_87);
xnor U701 (N_701,In_1500,In_1332);
or U702 (N_702,In_1031,N_445);
nor U703 (N_703,N_336,N_84);
and U704 (N_704,N_260,N_112);
or U705 (N_705,In_1433,In_1121);
and U706 (N_706,N_252,In_2213);
nor U707 (N_707,In_2221,In_655);
nor U708 (N_708,N_286,N_532);
nand U709 (N_709,In_1757,In_1001);
and U710 (N_710,N_226,N_456);
and U711 (N_711,In_618,In_2139);
nand U712 (N_712,In_1070,In_1042);
nand U713 (N_713,In_2316,In_433);
nor U714 (N_714,In_150,N_544);
nand U715 (N_715,N_63,N_483);
nor U716 (N_716,In_1263,N_213);
nor U717 (N_717,N_52,In_2024);
nor U718 (N_718,In_1306,In_1536);
nand U719 (N_719,In_1747,In_1216);
and U720 (N_720,N_589,In_787);
and U721 (N_721,In_1134,In_2261);
and U722 (N_722,N_88,In_2423);
nor U723 (N_723,In_1874,In_611);
or U724 (N_724,In_739,In_1942);
or U725 (N_725,In_1444,In_994);
and U726 (N_726,In_2058,N_295);
nor U727 (N_727,In_1157,N_374);
and U728 (N_728,N_613,N_177);
nor U729 (N_729,N_4,N_16);
and U730 (N_730,N_283,N_133);
and U731 (N_731,In_2466,N_167);
nor U732 (N_732,In_259,In_2232);
or U733 (N_733,In_791,In_926);
xnor U734 (N_734,In_1541,In_1036);
nor U735 (N_735,In_934,N_390);
or U736 (N_736,N_371,In_901);
nand U737 (N_737,In_136,In_481);
nor U738 (N_738,In_1635,N_46);
nand U739 (N_739,In_2377,In_299);
or U740 (N_740,N_368,N_464);
and U741 (N_741,N_21,In_1150);
and U742 (N_742,In_388,In_674);
and U743 (N_743,In_1489,N_543);
xor U744 (N_744,N_500,N_615);
or U745 (N_745,N_503,In_1155);
nand U746 (N_746,In_1147,In_1256);
nand U747 (N_747,In_1050,In_2179);
and U748 (N_748,N_473,In_412);
nand U749 (N_749,N_350,In_2182);
and U750 (N_750,In_223,In_664);
and U751 (N_751,In_2218,N_104);
nor U752 (N_752,In_1077,In_1450);
nor U753 (N_753,In_1227,N_202);
xnor U754 (N_754,In_1806,In_2201);
and U755 (N_755,In_1213,N_179);
or U756 (N_756,In_1491,In_1961);
or U757 (N_757,In_1116,In_1206);
or U758 (N_758,N_11,In_1950);
or U759 (N_759,In_1952,N_435);
nand U760 (N_760,In_751,In_2312);
or U761 (N_761,N_223,In_2163);
or U762 (N_762,In_2002,N_406);
nand U763 (N_763,N_279,N_3);
nor U764 (N_764,N_602,In_724);
nand U765 (N_765,In_2219,In_1469);
nor U766 (N_766,In_2121,In_676);
nor U767 (N_767,N_524,In_692);
and U768 (N_768,In_1868,In_1482);
or U769 (N_769,In_1333,N_23);
nand U770 (N_770,In_789,In_1709);
and U771 (N_771,In_1484,In_1066);
and U772 (N_772,In_2156,N_562);
or U773 (N_773,In_42,In_1596);
nand U774 (N_774,In_1328,In_2183);
nand U775 (N_775,In_1588,In_2345);
nand U776 (N_776,In_50,N_477);
or U777 (N_777,In_2006,In_2210);
nand U778 (N_778,In_587,In_21);
nand U779 (N_779,In_1546,In_1775);
nor U780 (N_780,N_578,In_969);
nor U781 (N_781,In_297,In_1705);
xnor U782 (N_782,In_2134,In_1365);
or U783 (N_783,N_346,In_364);
nor U784 (N_784,In_2490,N_377);
or U785 (N_785,In_214,In_2205);
xnor U786 (N_786,In_1442,N_345);
and U787 (N_787,In_1498,N_351);
nand U788 (N_788,N_198,N_236);
and U789 (N_789,In_2470,N_619);
nand U790 (N_790,In_282,In_812);
nor U791 (N_791,In_244,In_1674);
nand U792 (N_792,In_1567,In_947);
xor U793 (N_793,In_2343,In_1119);
or U794 (N_794,In_1231,N_258);
and U795 (N_795,N_45,In_2430);
and U796 (N_796,N_175,In_2339);
or U797 (N_797,In_257,In_512);
or U798 (N_798,N_100,N_97);
xnor U799 (N_799,In_69,In_1719);
nand U800 (N_800,In_1202,N_488);
nor U801 (N_801,In_955,In_1555);
nor U802 (N_802,In_785,In_1616);
or U803 (N_803,N_442,In_2385);
nand U804 (N_804,In_549,N_446);
or U805 (N_805,In_1851,In_1864);
and U806 (N_806,In_1837,In_1034);
or U807 (N_807,In_1100,In_471);
and U808 (N_808,In_1800,In_1410);
xnor U809 (N_809,N_553,In_2478);
xor U810 (N_810,In_976,In_816);
nand U811 (N_811,In_1299,In_1088);
nand U812 (N_812,In_2277,In_1308);
xnor U813 (N_813,In_1843,In_48);
and U814 (N_814,In_249,In_1707);
or U815 (N_815,In_968,N_623);
or U816 (N_816,N_614,In_10);
xor U817 (N_817,In_1421,N_72);
nor U818 (N_818,In_185,In_1067);
nor U819 (N_819,N_507,In_2314);
nor U820 (N_820,N_402,N_91);
and U821 (N_821,N_552,In_1680);
nand U822 (N_822,In_1352,In_701);
nand U823 (N_823,In_1456,In_1006);
nor U824 (N_824,In_2469,N_163);
nand U825 (N_825,In_1857,In_73);
and U826 (N_826,In_6,N_15);
or U827 (N_827,N_591,In_855);
nor U828 (N_828,In_2159,In_592);
nand U829 (N_829,In_530,In_144);
nor U830 (N_830,In_1991,N_160);
nand U831 (N_831,N_496,N_191);
nor U832 (N_832,In_1630,In_562);
xor U833 (N_833,In_2042,In_1727);
nor U834 (N_834,In_1530,In_276);
or U835 (N_835,N_17,In_1967);
nor U836 (N_836,N_329,N_38);
nand U837 (N_837,In_1557,N_287);
nand U838 (N_838,In_1828,In_798);
nand U839 (N_839,In_2123,In_2288);
xor U840 (N_840,In_911,In_890);
and U841 (N_841,In_1922,In_1254);
xor U842 (N_842,In_870,In_770);
or U843 (N_843,In_2299,In_23);
nand U844 (N_844,In_831,In_1793);
and U845 (N_845,In_1587,In_2402);
and U846 (N_846,In_740,In_234);
or U847 (N_847,N_51,N_416);
nor U848 (N_848,N_585,In_228);
nor U849 (N_849,In_1276,N_366);
and U850 (N_850,In_1357,In_2409);
and U851 (N_851,In_821,N_135);
nor U852 (N_852,N_34,N_69);
nand U853 (N_853,N_352,In_2329);
nor U854 (N_854,N_419,In_2267);
nand U855 (N_855,In_1898,In_663);
nor U856 (N_856,In_413,In_1581);
xnor U857 (N_857,In_721,In_2333);
nand U858 (N_858,In_1437,N_441);
nand U859 (N_859,In_685,In_340);
xor U860 (N_860,N_127,In_2398);
and U861 (N_861,In_1493,N_570);
nor U862 (N_862,In_2388,In_1038);
nor U863 (N_863,N_335,N_487);
nor U864 (N_864,N_605,N_504);
xor U865 (N_865,N_134,In_1453);
or U866 (N_866,In_725,N_564);
nor U867 (N_867,In_2265,In_47);
and U868 (N_868,N_367,In_1833);
and U869 (N_869,In_1717,In_902);
nand U870 (N_870,In_2441,In_1781);
and U871 (N_871,N_68,In_2424);
and U872 (N_872,In_2378,N_444);
xor U873 (N_873,N_101,In_1210);
and U874 (N_874,In_2130,In_813);
and U875 (N_875,In_154,In_1773);
nand U876 (N_876,N_196,In_2489);
or U877 (N_877,In_1063,In_985);
nand U878 (N_878,N_56,N_86);
xor U879 (N_879,In_1561,N_276);
nand U880 (N_880,N_180,N_582);
xor U881 (N_881,In_2176,In_767);
and U882 (N_882,In_195,N_370);
nand U883 (N_883,In_1300,N_81);
xor U884 (N_884,In_1400,N_307);
xor U885 (N_885,In_558,In_379);
or U886 (N_886,In_2406,N_251);
nor U887 (N_887,In_487,N_262);
and U888 (N_888,N_24,In_1565);
or U889 (N_889,In_2117,In_2225);
nor U890 (N_890,In_617,N_9);
nor U891 (N_891,In_2237,In_1449);
or U892 (N_892,In_2493,In_145);
and U893 (N_893,In_2178,In_643);
nand U894 (N_894,N_224,In_2040);
nor U895 (N_895,N_398,In_2041);
or U896 (N_896,N_332,In_1681);
and U897 (N_897,In_2165,In_1873);
or U898 (N_898,In_1439,In_1502);
xnor U899 (N_899,In_2373,N_568);
or U900 (N_900,N_57,In_2448);
and U901 (N_901,N_596,N_274);
xor U902 (N_902,In_2137,In_1841);
or U903 (N_903,In_1808,N_492);
xnor U904 (N_904,In_2000,In_1366);
nor U905 (N_905,In_527,In_278);
nand U906 (N_906,In_1005,In_2087);
and U907 (N_907,In_1904,In_313);
or U908 (N_908,In_169,N_522);
xor U909 (N_909,In_975,In_1269);
nand U910 (N_910,N_18,N_383);
and U911 (N_911,In_270,In_1209);
and U912 (N_912,In_67,N_269);
and U913 (N_913,N_119,N_128);
and U914 (N_914,In_1918,N_569);
or U915 (N_915,N_467,In_754);
xor U916 (N_916,In_761,In_0);
nand U917 (N_917,In_105,In_1866);
xnor U918 (N_918,N_29,In_557);
or U919 (N_919,N_420,In_2450);
or U920 (N_920,N_617,In_811);
xnor U921 (N_921,In_1571,In_330);
and U922 (N_922,In_4,In_1989);
or U923 (N_923,In_1068,In_1566);
and U924 (N_924,In_2067,N_327);
nor U925 (N_925,In_1859,In_1980);
or U926 (N_926,In_2342,In_1622);
or U927 (N_927,N_253,In_1023);
or U928 (N_928,N_89,N_110);
nor U929 (N_929,In_253,N_254);
nand U930 (N_930,In_2113,In_355);
nand U931 (N_931,In_2249,N_192);
xor U932 (N_932,In_1572,In_1169);
and U933 (N_933,In_1052,In_2233);
and U934 (N_934,N_121,In_1887);
and U935 (N_935,In_2437,In_1981);
xor U936 (N_936,N_139,In_1894);
xnor U937 (N_937,N_290,In_827);
nand U938 (N_938,N_314,N_426);
and U939 (N_939,In_25,In_1497);
and U940 (N_940,In_1512,N_338);
xor U941 (N_941,In_135,N_489);
xor U942 (N_942,In_1009,N_65);
nor U943 (N_943,In_2488,In_1186);
xnor U944 (N_944,In_312,In_1183);
nand U945 (N_945,In_1829,N_391);
and U946 (N_946,N_355,N_587);
or U947 (N_947,In_1928,N_28);
and U948 (N_948,In_2321,In_1562);
nor U949 (N_949,In_2292,In_2253);
or U950 (N_950,N_75,In_1058);
or U951 (N_951,N_206,In_809);
xnor U952 (N_952,In_15,N_131);
xnor U953 (N_953,In_1534,N_10);
or U954 (N_954,In_371,In_980);
or U955 (N_955,In_1072,N_622);
or U956 (N_956,In_616,In_1940);
xor U957 (N_957,In_1699,In_615);
nand U958 (N_958,In_590,In_122);
xnor U959 (N_959,N_44,In_2074);
nand U960 (N_960,In_2234,In_1358);
and U961 (N_961,N_58,In_84);
nand U962 (N_962,In_2291,In_2386);
nand U963 (N_963,In_1046,N_19);
or U964 (N_964,N_594,In_2084);
xnor U965 (N_965,In_2405,In_1083);
nor U966 (N_966,N_389,In_2278);
or U967 (N_967,N_470,In_490);
and U968 (N_968,In_657,In_341);
and U969 (N_969,In_2101,In_20);
nor U970 (N_970,N_523,In_1784);
nand U971 (N_971,In_1141,In_2098);
and U972 (N_972,N_322,In_45);
nor U973 (N_973,In_2352,In_1249);
nor U974 (N_974,N_227,In_132);
nor U975 (N_975,N_539,N_126);
nor U976 (N_976,N_311,N_574);
nor U977 (N_977,In_1382,N_407);
or U978 (N_978,N_536,N_540);
xnor U979 (N_979,In_1629,N_533);
xnor U980 (N_980,In_1769,N_590);
xor U981 (N_981,In_1262,In_967);
or U982 (N_982,In_854,In_1338);
or U983 (N_983,In_1341,In_1861);
and U984 (N_984,In_343,N_40);
nand U985 (N_985,In_2038,In_1028);
nor U986 (N_986,In_248,In_580);
nand U987 (N_987,In_786,In_1092);
and U988 (N_988,In_1343,In_2338);
xnor U989 (N_989,In_2400,N_264);
or U990 (N_990,In_2223,N_458);
xor U991 (N_991,N_430,In_1886);
and U992 (N_992,In_1145,In_2476);
nor U993 (N_993,In_2157,N_178);
xor U994 (N_994,N_476,In_1792);
or U995 (N_995,In_489,In_2189);
or U996 (N_996,In_1667,N_531);
or U997 (N_997,In_2059,N_598);
xnor U998 (N_998,In_138,N_132);
or U999 (N_999,In_2171,In_499);
xnor U1000 (N_1000,In_2185,N_501);
and U1001 (N_1001,In_293,N_55);
or U1002 (N_1002,In_250,In_2215);
nor U1003 (N_1003,N_187,In_3);
or U1004 (N_1004,N_365,In_1443);
xor U1005 (N_1005,In_2370,In_1168);
or U1006 (N_1006,N_59,In_1117);
nand U1007 (N_1007,N_462,In_1636);
and U1008 (N_1008,In_22,In_1915);
nor U1009 (N_1009,N_603,In_946);
xnor U1010 (N_1010,N_185,In_206);
nand U1011 (N_1011,In_1651,In_2196);
nand U1012 (N_1012,In_2422,N_94);
xor U1013 (N_1013,In_1461,In_2497);
or U1014 (N_1014,N_8,In_2181);
and U1015 (N_1015,In_1347,In_645);
nor U1016 (N_1016,In_1356,N_502);
nor U1017 (N_1017,N_173,In_759);
nor U1018 (N_1018,In_1403,In_666);
nor U1019 (N_1019,N_362,In_1460);
and U1020 (N_1020,N_47,In_1090);
nor U1021 (N_1021,In_843,In_470);
or U1022 (N_1022,N_171,In_1225);
nor U1023 (N_1023,In_1204,In_1737);
or U1024 (N_1024,In_1721,In_575);
xor U1025 (N_1025,In_32,In_1013);
nor U1026 (N_1026,In_1654,In_1964);
and U1027 (N_1027,In_2447,N_242);
and U1028 (N_1028,N_418,In_396);
nand U1029 (N_1029,In_1483,In_2090);
nand U1030 (N_1030,N_439,N_197);
nor U1031 (N_1031,In_1663,In_565);
xnor U1032 (N_1032,In_2401,In_727);
nand U1033 (N_1033,In_54,N_328);
nor U1034 (N_1034,In_1286,In_951);
and U1035 (N_1035,In_1951,N_215);
nand U1036 (N_1036,In_287,In_1890);
nor U1037 (N_1037,N_348,In_1026);
or U1038 (N_1038,In_954,N_151);
and U1039 (N_1039,In_1751,In_385);
or U1040 (N_1040,In_373,N_159);
or U1041 (N_1041,N_415,N_155);
nor U1042 (N_1042,In_2,In_1521);
and U1043 (N_1043,N_82,N_388);
nor U1044 (N_1044,In_1794,In_1743);
nor U1045 (N_1045,N_379,N_288);
xnor U1046 (N_1046,In_760,N_392);
or U1047 (N_1047,N_199,N_575);
nand U1048 (N_1048,N_537,In_810);
and U1049 (N_1049,In_1832,In_2135);
or U1050 (N_1050,In_1285,N_145);
and U1051 (N_1051,In_1106,In_1446);
xor U1052 (N_1052,N_194,In_178);
and U1053 (N_1053,N_296,In_1657);
xnor U1054 (N_1054,In_2393,In_7);
xnor U1055 (N_1055,In_2475,In_858);
or U1056 (N_1056,In_1057,In_818);
or U1057 (N_1057,In_1598,In_2262);
and U1058 (N_1058,N_71,In_820);
nand U1059 (N_1059,In_574,In_1321);
or U1060 (N_1060,In_2047,In_1631);
xor U1061 (N_1061,In_152,N_200);
xor U1062 (N_1062,In_402,In_1696);
and U1063 (N_1063,In_1921,In_1911);
nand U1064 (N_1064,In_1010,In_2129);
and U1065 (N_1065,In_1295,N_363);
and U1066 (N_1066,N_41,In_1653);
and U1067 (N_1067,In_1842,In_89);
xnor U1068 (N_1068,N_528,N_548);
nor U1069 (N_1069,In_752,N_149);
nand U1070 (N_1070,In_2073,In_180);
nor U1071 (N_1071,N_204,In_46);
or U1072 (N_1072,In_243,N_193);
or U1073 (N_1073,N_560,N_485);
and U1074 (N_1074,N_181,In_1671);
nand U1075 (N_1075,In_1907,In_1628);
nor U1076 (N_1076,In_1934,N_233);
nand U1077 (N_1077,In_1247,N_231);
nand U1078 (N_1078,N_333,N_111);
nor U1079 (N_1079,In_450,In_842);
nor U1080 (N_1080,In_1274,In_1956);
or U1081 (N_1081,In_1897,N_255);
or U1082 (N_1082,In_217,N_292);
nand U1083 (N_1083,In_1367,In_540);
or U1084 (N_1084,N_184,In_2417);
nor U1085 (N_1085,N_109,N_36);
xnor U1086 (N_1086,In_85,N_318);
nor U1087 (N_1087,In_1101,In_1713);
and U1088 (N_1088,N_27,In_1162);
and U1089 (N_1089,N_214,In_1948);
nor U1090 (N_1090,N_510,N_584);
and U1091 (N_1091,In_1831,In_665);
or U1092 (N_1092,N_125,In_660);
or U1093 (N_1093,In_2304,In_127);
or U1094 (N_1094,In_2274,In_109);
or U1095 (N_1095,In_1289,In_2444);
or U1096 (N_1096,In_1684,In_1393);
and U1097 (N_1097,In_741,N_422);
xnor U1098 (N_1098,In_173,In_347);
nand U1099 (N_1099,In_718,In_1621);
nand U1100 (N_1100,In_2452,In_1218);
nor U1101 (N_1101,In_1105,In_981);
nand U1102 (N_1102,In_1860,N_513);
or U1103 (N_1103,In_544,In_1033);
or U1104 (N_1104,In_2220,In_51);
xnor U1105 (N_1105,In_2080,In_555);
nand U1106 (N_1106,In_1261,N_240);
xnor U1107 (N_1107,In_675,N_428);
xor U1108 (N_1108,N_535,N_344);
nor U1109 (N_1109,In_377,In_460);
and U1110 (N_1110,In_1742,In_2068);
or U1111 (N_1111,In_2275,In_327);
and U1112 (N_1112,In_445,N_484);
xnor U1113 (N_1113,In_2147,In_1659);
xnor U1114 (N_1114,In_1199,In_1291);
nor U1115 (N_1115,N_271,In_2151);
or U1116 (N_1116,In_2324,In_268);
nand U1117 (N_1117,In_797,In_1236);
xnor U1118 (N_1118,In_750,N_518);
nand U1119 (N_1119,In_859,In_2009);
nand U1120 (N_1120,In_1525,In_1968);
nand U1121 (N_1121,In_2432,In_1429);
or U1122 (N_1122,N_273,In_390);
xnor U1123 (N_1123,In_2416,N_530);
or U1124 (N_1124,In_1240,N_219);
xor U1125 (N_1125,In_850,In_515);
xnor U1126 (N_1126,N_172,In_233);
nand U1127 (N_1127,In_2062,In_1893);
xor U1128 (N_1128,In_1574,N_583);
nand U1129 (N_1129,N_394,N_113);
xor U1130 (N_1130,In_1871,In_507);
or U1131 (N_1131,N_294,In_164);
nor U1132 (N_1132,In_1047,N_618);
xor U1133 (N_1133,In_304,In_1040);
and U1134 (N_1134,N_417,N_443);
and U1135 (N_1135,In_2110,N_607);
and U1136 (N_1136,N_432,In_1207);
xor U1137 (N_1137,N_404,In_1817);
or U1138 (N_1138,N_373,N_592);
or U1139 (N_1139,In_266,In_1364);
nor U1140 (N_1140,In_203,In_1187);
nand U1141 (N_1141,In_669,In_1035);
nor U1142 (N_1142,In_271,In_683);
nor U1143 (N_1143,In_2115,N_620);
nand U1144 (N_1144,In_1749,N_571);
or U1145 (N_1145,In_1863,In_644);
nor U1146 (N_1146,In_2143,N_13);
xnor U1147 (N_1147,In_603,In_161);
and U1148 (N_1148,In_1997,N_573);
nand U1149 (N_1149,N_284,In_1591);
nor U1150 (N_1150,In_961,In_987);
or U1151 (N_1151,In_2340,In_1182);
or U1152 (N_1152,In_877,N_463);
nor U1153 (N_1153,N_554,N_316);
nand U1154 (N_1154,In_1342,N_339);
or U1155 (N_1155,N_22,In_483);
and U1156 (N_1156,In_454,In_2453);
and U1157 (N_1157,N_604,In_992);
nand U1158 (N_1158,N_497,In_1318);
nor U1159 (N_1159,In_75,N_517);
xnor U1160 (N_1160,In_1925,In_121);
xor U1161 (N_1161,In_2004,In_2140);
or U1162 (N_1162,N_225,In_548);
or U1163 (N_1163,In_2016,N_556);
xnor U1164 (N_1164,N_140,In_640);
or U1165 (N_1165,In_845,N_421);
or U1166 (N_1166,In_1246,In_1905);
xnor U1167 (N_1167,N_566,In_817);
or U1168 (N_1168,N_230,N_414);
and U1169 (N_1169,N_120,In_1736);
nand U1170 (N_1170,N_340,N_106);
or U1171 (N_1171,In_1847,In_1939);
or U1172 (N_1172,N_491,In_1390);
and U1173 (N_1173,N_64,N_380);
or U1174 (N_1174,In_853,In_2065);
nand U1175 (N_1175,N_186,In_1019);
nor U1176 (N_1176,N_506,In_1173);
nor U1177 (N_1177,N_449,In_1323);
xor U1178 (N_1178,N_136,N_347);
and U1179 (N_1179,In_1414,In_2075);
and U1180 (N_1180,In_1936,In_526);
nor U1181 (N_1181,N_235,N_505);
and U1182 (N_1182,In_2027,In_848);
nor U1183 (N_1183,In_1146,In_2148);
nor U1184 (N_1184,N_337,In_36);
nand U1185 (N_1185,N_245,In_2246);
nor U1186 (N_1186,In_2407,N_152);
or U1187 (N_1187,N_270,N_247);
or U1188 (N_1188,In_2132,In_2438);
nor U1189 (N_1189,In_1782,In_63);
nor U1190 (N_1190,N_342,In_2309);
xnor U1191 (N_1191,N_205,N_107);
or U1192 (N_1192,N_399,In_1470);
and U1193 (N_1193,In_451,In_241);
xor U1194 (N_1194,In_1476,N_538);
xnor U1195 (N_1195,In_682,In_151);
xor U1196 (N_1196,In_181,N_396);
nand U1197 (N_1197,In_712,N_92);
xnor U1198 (N_1198,In_2142,In_2443);
or U1199 (N_1199,In_826,In_2260);
or U1200 (N_1200,In_430,In_1455);
nor U1201 (N_1201,N_354,In_1369);
nor U1202 (N_1202,N_166,In_1528);
nand U1203 (N_1203,N_30,N_429);
xnor U1204 (N_1204,N_453,In_1257);
nand U1205 (N_1205,In_128,In_357);
and U1206 (N_1206,In_1349,In_1613);
nand U1207 (N_1207,N_146,In_1586);
or U1208 (N_1208,In_8,N_624);
or U1209 (N_1209,In_1370,In_488);
xnor U1210 (N_1210,In_1376,N_610);
nand U1211 (N_1211,In_1158,In_2390);
nor U1212 (N_1212,N_309,N_546);
nor U1213 (N_1213,N_85,In_2302);
or U1214 (N_1214,In_1550,N_208);
nand U1215 (N_1215,In_2349,In_137);
nand U1216 (N_1216,N_408,In_1234);
or U1217 (N_1217,In_1776,In_2428);
nand U1218 (N_1218,In_284,In_352);
nand U1219 (N_1219,N_150,N_519);
xnor U1220 (N_1220,In_1292,In_1774);
or U1221 (N_1221,In_1798,In_258);
xnor U1222 (N_1222,N_425,In_1612);
nand U1223 (N_1223,In_635,In_828);
xnor U1224 (N_1224,In_876,In_1930);
and U1225 (N_1225,In_823,In_1929);
xor U1226 (N_1226,In_171,In_1268);
or U1227 (N_1227,In_1966,In_1039);
or U1228 (N_1228,N_67,In_1610);
and U1229 (N_1229,N_170,In_350);
nand U1230 (N_1230,In_386,N_498);
nand U1231 (N_1231,In_508,In_915);
or U1232 (N_1232,N_37,In_129);
nor U1233 (N_1233,N_77,In_457);
xor U1234 (N_1234,In_2032,In_1954);
nor U1235 (N_1235,N_579,In_847);
and U1236 (N_1236,In_1723,In_166);
xnor U1237 (N_1237,N_115,In_568);
nand U1238 (N_1238,N_130,In_661);
and U1239 (N_1239,N_256,N_156);
xnor U1240 (N_1240,N_356,N_465);
nand U1241 (N_1241,In_534,In_1481);
or U1242 (N_1242,N_478,In_1025);
nor U1243 (N_1243,N_278,In_1919);
or U1244 (N_1244,In_2380,N_609);
nor U1245 (N_1245,N_369,In_1423);
nand U1246 (N_1246,In_2072,In_62);
xnor U1247 (N_1247,N_102,In_779);
nand U1248 (N_1248,In_348,In_263);
nor U1249 (N_1249,In_2481,In_119);
nand U1250 (N_1250,In_49,N_508);
and U1251 (N_1251,In_1029,N_749);
nor U1252 (N_1252,N_495,N_1056);
nand U1253 (N_1253,N_1236,In_2012);
xor U1254 (N_1254,In_2077,In_2211);
or U1255 (N_1255,N_87,N_1149);
nor U1256 (N_1256,N_1057,In_81);
or U1257 (N_1257,In_277,N_401);
or U1258 (N_1258,N_1148,N_637);
xor U1259 (N_1259,N_886,In_1960);
and U1260 (N_1260,N_726,N_990);
nor U1261 (N_1261,N_1136,N_343);
nor U1262 (N_1262,N_90,In_1353);
nor U1263 (N_1263,N_878,In_1163);
and U1264 (N_1264,N_557,N_1027);
or U1265 (N_1265,N_772,In_1599);
and U1266 (N_1266,In_2421,N_838);
xor U1267 (N_1267,N_781,In_1176);
and U1268 (N_1268,N_1020,N_386);
xnor U1269 (N_1269,N_829,In_72);
and U1270 (N_1270,N_1205,N_731);
nor U1271 (N_1271,N_835,N_625);
nor U1272 (N_1272,In_1527,N_1069);
and U1273 (N_1273,N_1007,N_845);
nor U1274 (N_1274,In_764,N_822);
xnor U1275 (N_1275,N_672,In_1556);
xor U1276 (N_1276,N_1146,N_854);
and U1277 (N_1277,N_1066,In_143);
nand U1278 (N_1278,In_468,N_649);
nor U1279 (N_1279,N_945,In_1184);
nor U1280 (N_1280,In_1326,N_677);
nand U1281 (N_1281,N_447,In_131);
and U1282 (N_1282,N_1188,N_968);
nor U1283 (N_1283,N_411,In_1127);
nand U1284 (N_1284,N_974,N_1117);
nand U1285 (N_1285,N_960,N_963);
or U1286 (N_1286,In_1085,N_1154);
or U1287 (N_1287,In_2031,N_689);
and U1288 (N_1288,N_83,N_770);
and U1289 (N_1289,N_1097,N_910);
nor U1290 (N_1290,N_1121,N_810);
nor U1291 (N_1291,N_1110,In_1239);
nor U1292 (N_1292,In_1464,N_750);
nor U1293 (N_1293,In_2021,In_584);
nor U1294 (N_1294,In_68,N_987);
and U1295 (N_1295,N_1050,N_1132);
or U1296 (N_1296,In_1884,In_523);
or U1297 (N_1297,N_1091,In_553);
xor U1298 (N_1298,N_753,N_704);
or U1299 (N_1299,In_1986,N_480);
and U1300 (N_1300,N_853,In_892);
xnor U1301 (N_1301,N_766,N_955);
and U1302 (N_1302,In_1245,N_1224);
or U1303 (N_1303,N_948,N_889);
xor U1304 (N_1304,N_1003,N_685);
or U1305 (N_1305,In_441,N_26);
nand U1306 (N_1306,N_263,In_326);
or U1307 (N_1307,N_268,N_410);
nand U1308 (N_1308,In_310,In_1301);
nand U1309 (N_1309,N_1158,In_1545);
and U1310 (N_1310,N_636,N_239);
and U1311 (N_1311,N_448,N_1130);
nor U1312 (N_1312,N_741,N_1118);
or U1313 (N_1313,In_124,N_839);
and U1314 (N_1314,N_147,N_710);
or U1315 (N_1315,N_785,N_451);
xnor U1316 (N_1316,N_248,In_272);
nand U1317 (N_1317,N_760,N_1037);
nor U1318 (N_1318,N_979,In_2298);
and U1319 (N_1319,N_877,In_1294);
xor U1320 (N_1320,N_122,N_777);
nand U1321 (N_1321,N_819,N_567);
xnor U1322 (N_1322,N_857,N_1026);
and U1323 (N_1323,N_944,N_216);
nand U1324 (N_1324,N_836,In_878);
nor U1325 (N_1325,In_110,N_201);
nand U1326 (N_1326,N_203,N_905);
nand U1327 (N_1327,In_2035,N_1193);
or U1328 (N_1328,N_79,N_863);
nand U1329 (N_1329,N_1035,N_209);
or U1330 (N_1330,In_88,N_802);
nand U1331 (N_1331,In_126,In_2076);
nor U1332 (N_1332,N_746,N_875);
and U1333 (N_1333,In_1819,N_323);
nand U1334 (N_1334,In_153,In_524);
nand U1335 (N_1335,In_101,In_2048);
and U1336 (N_1336,In_423,N_951);
nand U1337 (N_1337,In_1355,N_971);
or U1338 (N_1338,N_1145,N_783);
nand U1339 (N_1339,In_2094,N_246);
nor U1340 (N_1340,N_137,N_959);
and U1341 (N_1341,N_918,N_250);
nand U1342 (N_1342,N_1072,N_572);
nand U1343 (N_1343,N_999,In_290);
nand U1344 (N_1344,In_2371,N_493);
or U1345 (N_1345,N_933,N_881);
and U1346 (N_1346,In_838,N_545);
nand U1347 (N_1347,N_1153,N_709);
nand U1348 (N_1348,In_473,N_1024);
and U1349 (N_1349,N_734,N_1089);
xor U1350 (N_1350,N_699,N_1046);
nor U1351 (N_1351,N_289,In_401);
nor U1352 (N_1352,N_1184,In_1392);
or U1353 (N_1353,N_972,In_1563);
and U1354 (N_1354,N_956,In_1646);
or U1355 (N_1355,N_847,N_1225);
nand U1356 (N_1356,N_313,N_744);
or U1357 (N_1357,In_966,N_259);
nand U1358 (N_1358,In_29,In_815);
and U1359 (N_1359,N_1206,In_1627);
or U1360 (N_1360,In_449,In_14);
and U1361 (N_1361,N_326,N_1126);
nor U1362 (N_1362,N_158,In_39);
nand U1363 (N_1363,N_942,In_1027);
xnor U1364 (N_1364,N_742,In_783);
and U1365 (N_1365,N_54,N_841);
nor U1366 (N_1366,N_1036,N_775);
or U1367 (N_1367,N_930,N_816);
nor U1368 (N_1368,N_923,N_748);
nor U1369 (N_1369,N_647,In_1619);
or U1370 (N_1370,N_330,N_995);
nand U1371 (N_1371,In_1547,N_1100);
xnor U1372 (N_1372,In_484,N_1226);
xor U1373 (N_1373,N_1210,N_1157);
nand U1374 (N_1374,N_499,N_349);
or U1375 (N_1375,N_558,N_325);
nand U1376 (N_1376,N_95,N_1084);
xor U1377 (N_1377,N_826,In_1820);
and U1378 (N_1378,N_920,In_1978);
nand U1379 (N_1379,N_936,N_550);
nor U1380 (N_1380,In_232,In_1689);
and U1381 (N_1381,In_1505,In_693);
xnor U1382 (N_1382,N_901,N_49);
nand U1383 (N_1383,In_2280,In_1885);
or U1384 (N_1384,In_677,N_645);
or U1385 (N_1385,In_614,In_13);
xnor U1386 (N_1386,In_1222,In_1412);
xor U1387 (N_1387,In_194,In_2296);
or U1388 (N_1388,N_1237,N_1015);
nand U1389 (N_1389,N_682,N_424);
and U1390 (N_1390,N_803,In_1840);
nor U1391 (N_1391,N_285,N_1219);
nand U1392 (N_1392,N_220,N_745);
or U1393 (N_1393,N_393,N_1107);
and U1394 (N_1394,N_1022,N_302);
and U1395 (N_1395,N_1180,In_465);
xor U1396 (N_1396,In_1537,In_999);
nand U1397 (N_1397,In_1454,N_1160);
and U1398 (N_1398,In_318,N_916);
or U1399 (N_1399,N_1212,In_291);
or U1400 (N_1400,In_2170,In_2344);
or U1401 (N_1401,N_1101,N_732);
xor U1402 (N_1402,N_702,N_969);
nand U1403 (N_1403,N_795,N_638);
xor U1404 (N_1404,N_358,In_717);
or U1405 (N_1405,N_593,N_1085);
or U1406 (N_1406,N_830,N_143);
and U1407 (N_1407,In_2372,N_118);
nand U1408 (N_1408,N_1079,N_756);
or U1409 (N_1409,In_960,In_799);
or U1410 (N_1410,In_2001,N_828);
and U1411 (N_1411,In_1041,N_757);
or U1412 (N_1412,N_1033,N_1208);
and U1413 (N_1413,In_2297,In_839);
and U1414 (N_1414,N_752,N_914);
and U1415 (N_1415,N_353,N_985);
nor U1416 (N_1416,N_1109,In_2318);
and U1417 (N_1417,N_1175,N_1242);
nand U1418 (N_1418,N_992,N_658);
or U1419 (N_1419,In_1270,N_953);
or U1420 (N_1420,N_669,In_589);
or U1421 (N_1421,N_207,N_891);
and U1422 (N_1422,N_879,N_873);
nand U1423 (N_1423,N_1065,N_33);
or U1424 (N_1424,N_1195,N_526);
or U1425 (N_1425,N_698,N_703);
or U1426 (N_1426,N_600,N_947);
nand U1427 (N_1427,N_931,N_475);
and U1428 (N_1428,N_176,N_315);
and U1429 (N_1429,In_1494,In_2039);
or U1430 (N_1430,In_463,In_1913);
xnor U1431 (N_1431,N_921,In_2264);
and U1432 (N_1432,N_1231,N_641);
and U1433 (N_1433,N_275,N_1131);
nand U1434 (N_1434,N_737,N_688);
nand U1435 (N_1435,In_710,In_103);
xor U1436 (N_1436,In_2427,In_2125);
or U1437 (N_1437,N_1115,N_1070);
and U1438 (N_1438,N_161,N_812);
xor U1439 (N_1439,In_2055,N_1172);
nand U1440 (N_1440,In_120,N_78);
and U1441 (N_1441,N_1238,N_642);
and U1442 (N_1442,In_1650,In_1012);
or U1443 (N_1443,N_320,N_1176);
nand U1444 (N_1444,N_1241,N_481);
or U1445 (N_1445,N_722,In_1373);
nor U1446 (N_1446,N_1207,N_154);
xnor U1447 (N_1447,In_978,N_1189);
nand U1448 (N_1448,N_509,In_1515);
nor U1449 (N_1449,N_1080,N_1152);
nor U1450 (N_1450,N_1049,N_954);
nand U1451 (N_1451,In_2392,In_104);
or U1452 (N_1452,N_1128,N_427);
or U1453 (N_1453,In_294,N_1106);
xnor U1454 (N_1454,N_764,In_1267);
nor U1455 (N_1455,N_1090,N_776);
nand U1456 (N_1456,N_694,N_1209);
xnor U1457 (N_1457,N_676,N_1082);
nand U1458 (N_1458,N_162,N_984);
nor U1459 (N_1459,N_639,In_339);
nor U1460 (N_1460,In_689,N_844);
nor U1461 (N_1461,In_267,N_626);
nand U1462 (N_1462,N_317,In_772);
nand U1463 (N_1463,In_370,In_963);
or U1464 (N_1464,In_1962,N_687);
nand U1465 (N_1465,N_970,N_423);
xnor U1466 (N_1466,In_2030,In_165);
xnor U1467 (N_1467,In_495,N_952);
xnor U1468 (N_1468,N_880,N_157);
or U1469 (N_1469,N_1161,N_471);
nor U1470 (N_1470,N_740,N_1245);
xnor U1471 (N_1471,N_1034,N_1139);
and U1472 (N_1472,In_2449,N_640);
xor U1473 (N_1473,N_997,N_988);
nand U1474 (N_1474,In_1487,N_516);
xnor U1475 (N_1475,In_1264,N_723);
nand U1476 (N_1476,In_397,In_649);
nor U1477 (N_1477,N_1196,N_60);
nor U1478 (N_1478,N_228,N_1083);
and U1479 (N_1479,In_686,In_1384);
or U1480 (N_1480,N_1230,N_693);
nand U1481 (N_1481,N_800,N_413);
and U1482 (N_1482,N_62,N_243);
xnor U1483 (N_1483,In_200,N_1054);
nand U1484 (N_1484,N_720,In_226);
nand U1485 (N_1485,In_1248,N_902);
nand U1486 (N_1486,In_631,N_1102);
or U1487 (N_1487,N_1,In_1577);
or U1488 (N_1488,N_707,In_1037);
nand U1489 (N_1489,N_1029,N_1051);
or U1490 (N_1490,N_792,N_1190);
nor U1491 (N_1491,N_1221,N_341);
and U1492 (N_1492,N_381,In_174);
and U1493 (N_1493,N_789,N_461);
nor U1494 (N_1494,N_981,N_460);
nor U1495 (N_1495,N_635,N_103);
nand U1496 (N_1496,N_899,N_779);
nand U1497 (N_1497,N_865,In_493);
or U1498 (N_1498,N_12,N_747);
and U1499 (N_1499,N_66,N_1047);
or U1500 (N_1500,In_1645,In_2341);
xnor U1501 (N_1501,N_941,N_105);
and U1502 (N_1502,N_1048,In_2494);
and U1503 (N_1503,N_1204,In_255);
xor U1504 (N_1504,N_1181,In_2491);
and U1505 (N_1505,In_1523,N_928);
xor U1506 (N_1506,In_897,In_898);
xor U1507 (N_1507,N_695,N_466);
nor U1508 (N_1508,In_190,In_1544);
nand U1509 (N_1509,N_858,N_434);
xor U1510 (N_1510,In_1397,N_713);
nand U1511 (N_1511,N_1201,In_274);
xnor U1512 (N_1512,In_1181,N_763);
xnor U1513 (N_1513,In_1084,N_525);
or U1514 (N_1514,N_986,In_913);
and U1515 (N_1515,N_431,N_25);
and U1516 (N_1516,N_627,N_994);
and U1517 (N_1517,In_2175,In_1708);
nand U1518 (N_1518,N_1138,N_1004);
or U1519 (N_1519,N_1099,N_364);
or U1520 (N_1520,N_1010,In_1167);
xnor U1521 (N_1521,N_794,In_585);
nor U1522 (N_1522,In_97,N_1017);
and U1523 (N_1523,N_739,N_189);
or U1524 (N_1524,N_1232,N_733);
nor U1525 (N_1525,N_1140,N_238);
and U1526 (N_1526,N_1187,N_1009);
nand U1527 (N_1527,N_382,N_821);
or U1528 (N_1528,N_728,In_1959);
xnor U1529 (N_1529,N_0,N_868);
nor U1530 (N_1530,In_880,In_613);
and U1531 (N_1531,In_1002,N_904);
nor U1532 (N_1532,In_945,In_1395);
and U1533 (N_1533,In_1658,N_906);
and U1534 (N_1534,N_165,In_2145);
nand U1535 (N_1535,N_996,N_629);
and U1536 (N_1536,N_743,N_1246);
nor U1537 (N_1537,N_666,N_1018);
nor U1538 (N_1538,N_861,In_1595);
or U1539 (N_1539,N_400,N_874);
xnor U1540 (N_1540,In_2108,N_946);
xnor U1541 (N_1541,In_737,In_1718);
nand U1542 (N_1542,N_966,N_1218);
nand U1543 (N_1543,In_1590,N_261);
nor U1544 (N_1544,N_872,N_690);
xor U1545 (N_1545,N_39,In_1334);
or U1546 (N_1546,N_643,N_304);
nand U1547 (N_1547,N_769,In_1984);
nor U1548 (N_1548,N_1213,N_277);
and U1549 (N_1549,N_1093,N_885);
and U1550 (N_1550,In_2128,In_2173);
xnor U1551 (N_1551,N_706,In_623);
nor U1552 (N_1552,N_1071,N_818);
xnor U1553 (N_1553,In_251,N_1227);
or U1554 (N_1554,N_1075,N_267);
or U1555 (N_1555,N_1067,N_866);
nor U1556 (N_1556,N_1192,In_455);
or U1557 (N_1557,N_1223,N_896);
and U1558 (N_1558,In_425,N_1215);
or U1559 (N_1559,N_611,N_5);
nor U1560 (N_1560,N_934,N_962);
nor U1561 (N_1561,N_375,In_841);
and U1562 (N_1562,N_1214,N_412);
xnor U1563 (N_1563,N_937,N_1055);
nor U1564 (N_1564,N_727,N_1133);
nand U1565 (N_1565,N_1191,In_184);
xnor U1566 (N_1566,N_576,N_949);
or U1567 (N_1567,N_20,N_870);
and U1568 (N_1568,In_1854,N_124);
xnor U1569 (N_1569,In_642,N_565);
or U1570 (N_1570,N_925,In_1445);
xor U1571 (N_1571,N_793,In_332);
or U1572 (N_1572,N_1038,In_1611);
nor U1573 (N_1573,N_982,N_1030);
and U1574 (N_1574,N_1179,N_1222);
xor U1575 (N_1575,N_1229,N_1244);
or U1576 (N_1576,In_909,N_940);
and U1577 (N_1577,N_1194,N_869);
xnor U1578 (N_1578,N_490,N_924);
xor U1579 (N_1579,N_814,N_796);
and U1580 (N_1580,N_909,N_673);
xor U1581 (N_1581,N_108,In_1194);
or U1582 (N_1582,In_1741,N_759);
or U1583 (N_1583,In_2319,N_993);
nand U1584 (N_1584,N_1170,N_1073);
nand U1585 (N_1585,N_114,In_118);
nor U1586 (N_1586,N_1078,N_1144);
nor U1587 (N_1587,N_831,N_1105);
nor U1588 (N_1588,In_333,N_588);
or U1589 (N_1589,N_1013,N_837);
xor U1590 (N_1590,N_659,N_751);
or U1591 (N_1591,N_468,In_1520);
nor U1592 (N_1592,N_534,N_630);
or U1593 (N_1593,N_334,In_389);
nand U1594 (N_1594,N_244,N_1199);
and U1595 (N_1595,N_833,In_1908);
nor U1596 (N_1596,N_683,In_728);
xor U1597 (N_1597,In_1582,In_953);
xor U1598 (N_1598,N_1098,N_633);
nand U1599 (N_1599,In_887,In_1516);
or U1600 (N_1600,N_980,N_153);
xnor U1601 (N_1601,N_1177,N_1127);
nor U1602 (N_1602,N_851,In_627);
nor U1603 (N_1603,In_366,In_148);
nor U1604 (N_1604,In_2353,In_1517);
or U1605 (N_1605,N_1165,N_1124);
or U1606 (N_1606,In_2200,In_1280);
nand U1607 (N_1607,N_1239,N_1040);
nor U1608 (N_1608,N_711,N_74);
and U1609 (N_1609,In_681,N_547);
and U1610 (N_1610,In_807,N_771);
xor U1611 (N_1611,N_1041,In_525);
or U1612 (N_1612,N_652,In_628);
or U1613 (N_1613,N_1182,N_701);
nor U1614 (N_1614,N_549,N_670);
or U1615 (N_1615,In_1643,N_385);
xnor U1616 (N_1616,N_1156,N_459);
or U1617 (N_1617,N_820,N_628);
or U1618 (N_1618,N_116,In_958);
nand U1619 (N_1619,In_2330,In_2063);
and U1620 (N_1620,N_671,N_842);
nor U1621 (N_1621,N_1217,N_663);
nand U1622 (N_1622,In_539,In_1432);
and U1623 (N_1623,N_846,N_35);
or U1624 (N_1624,In_2435,In_1201);
xor U1625 (N_1625,In_2335,In_2472);
or U1626 (N_1626,N_96,In_2461);
nor U1627 (N_1627,N_736,N_1059);
nand U1628 (N_1628,N_1248,N_1045);
or U1629 (N_1629,In_1388,N_700);
xnor U1630 (N_1630,N_50,N_897);
xnor U1631 (N_1631,N_714,In_1241);
or U1632 (N_1632,N_882,In_1809);
or U1633 (N_1633,In_671,N_319);
nor U1634 (N_1634,N_1120,N_849);
or U1635 (N_1635,N_938,N_1125);
nand U1636 (N_1636,In_974,N_804);
or U1637 (N_1637,N_1032,N_843);
nand U1638 (N_1638,N_1167,N_718);
nand U1639 (N_1639,In_678,N_1006);
nand U1640 (N_1640,N_1129,N_656);
or U1641 (N_1641,In_1789,N_321);
xnor U1642 (N_1642,N_667,N_1053);
and U1643 (N_1643,In_1975,N_514);
or U1644 (N_1644,N_123,N_331);
xnor U1645 (N_1645,N_1141,N_825);
nor U1646 (N_1646,N_1081,N_211);
or U1647 (N_1647,In_286,N_801);
and U1648 (N_1648,N_61,N_1174);
nand U1649 (N_1649,N_597,N_651);
xor U1650 (N_1650,N_1092,N_957);
and U1651 (N_1651,N_222,N_650);
nor U1652 (N_1652,N_1135,N_939);
or U1653 (N_1653,N_817,In_606);
nand U1654 (N_1654,In_376,N_1216);
or U1655 (N_1655,N_1086,In_1477);
nor U1656 (N_1656,N_1062,N_680);
or U1657 (N_1657,N_32,N_915);
nand U1658 (N_1658,N_520,In_1185);
nor U1659 (N_1659,N_14,In_1943);
nor U1660 (N_1660,In_1401,N_1123);
or U1661 (N_1661,N_827,In_1132);
and U1662 (N_1662,N_117,N_438);
nand U1663 (N_1663,N_908,In_1730);
xor U1664 (N_1664,In_1818,In_1969);
nor U1665 (N_1665,N_991,N_1134);
or U1666 (N_1666,In_1076,N_376);
and U1667 (N_1667,N_1119,N_1052);
nor U1668 (N_1668,N_983,N_665);
nor U1669 (N_1669,N_686,N_1198);
nand U1670 (N_1670,N_1200,In_2455);
or U1671 (N_1671,N_965,In_1126);
or U1672 (N_1672,N_42,In_1947);
or U1673 (N_1673,N_648,N_1094);
nand U1674 (N_1674,N_234,N_266);
nor U1675 (N_1675,In_2158,In_1661);
xnor U1676 (N_1676,In_1748,In_595);
xor U1677 (N_1677,In_1108,In_2462);
nand U1678 (N_1678,In_130,N_387);
nand U1679 (N_1679,In_1230,In_706);
or U1680 (N_1680,In_2116,N_721);
or U1681 (N_1681,N_469,In_1568);
and U1682 (N_1682,N_511,In_2480);
and U1683 (N_1683,N_437,N_813);
and U1684 (N_1684,N_834,In_1889);
nor U1685 (N_1685,N_1162,In_998);
or U1686 (N_1686,N_608,In_1130);
and U1687 (N_1687,N_716,In_1522);
nand U1688 (N_1688,N_1058,N_1183);
and U1689 (N_1689,N_472,N_890);
xor U1690 (N_1690,In_2317,N_1112);
nand U1691 (N_1691,N_1005,N_1186);
or U1692 (N_1692,N_917,N_799);
xnor U1693 (N_1693,N_735,N_324);
nand U1694 (N_1694,In_1575,In_1160);
and U1695 (N_1695,In_1398,In_2396);
or U1696 (N_1696,N_832,N_778);
nor U1697 (N_1697,N_780,N_977);
nand U1698 (N_1698,In_1044,N_1023);
xor U1699 (N_1699,N_210,N_912);
xor U1700 (N_1700,In_1177,N_378);
or U1701 (N_1701,N_976,N_2);
and U1702 (N_1702,N_359,N_612);
xnor U1703 (N_1703,N_712,In_1224);
nand U1704 (N_1704,N_855,N_99);
or U1705 (N_1705,N_409,In_1409);
or U1706 (N_1706,N_929,N_848);
nor U1707 (N_1707,In_1238,In_100);
nand U1708 (N_1708,N_926,N_1008);
xor U1709 (N_1709,In_329,In_2190);
nand U1710 (N_1710,In_429,N_927);
or U1711 (N_1711,N_563,N_48);
or U1712 (N_1712,N_903,N_898);
nor U1713 (N_1713,In_2381,N_31);
and U1714 (N_1714,N_678,In_599);
nor U1715 (N_1715,N_237,N_301);
nand U1716 (N_1716,In_914,In_965);
or U1717 (N_1717,N_767,In_1633);
and U1718 (N_1718,N_717,N_357);
xor U1719 (N_1719,N_998,N_291);
nor U1720 (N_1720,N_755,N_768);
and U1721 (N_1721,N_1243,In_1094);
nor U1722 (N_1722,In_2357,N_76);
xor U1723 (N_1723,In_2362,In_1852);
nor U1724 (N_1724,N_893,N_911);
or U1725 (N_1725,In_56,N_265);
nand U1726 (N_1726,N_144,In_1354);
nand U1727 (N_1727,N_871,In_2310);
nand U1728 (N_1728,N_482,N_303);
xnor U1729 (N_1729,N_70,In_1089);
nand U1730 (N_1730,In_1734,N_907);
nor U1731 (N_1731,N_452,N_1197);
nand U1732 (N_1732,N_1228,N_486);
and U1733 (N_1733,N_788,In_1805);
or U1734 (N_1734,N_1108,In_1451);
nor U1735 (N_1735,In_977,N_280);
nor U1736 (N_1736,In_1895,In_1531);
or U1737 (N_1737,N_815,N_1095);
or U1738 (N_1738,N_217,In_211);
and U1739 (N_1739,In_1768,N_1202);
xor U1740 (N_1740,In_769,N_634);
or U1741 (N_1741,In_1791,In_400);
and U1742 (N_1742,N_1074,N_856);
nor U1743 (N_1743,N_1011,In_588);
xnor U1744 (N_1744,N_668,N_1044);
nor U1745 (N_1745,N_892,In_2479);
and U1746 (N_1746,In_107,N_1021);
and U1747 (N_1747,N_895,N_616);
nand U1748 (N_1748,N_798,N_900);
nor U1749 (N_1749,N_174,In_1302);
and U1750 (N_1750,In_380,N_894);
nor U1751 (N_1751,In_1955,N_1211);
or U1752 (N_1752,In_1881,In_520);
nand U1753 (N_1753,N_229,In_2049);
and U1754 (N_1754,N_852,N_1155);
or U1755 (N_1755,In_183,In_398);
nand U1756 (N_1756,N_824,N_791);
and U1757 (N_1757,N_555,N_1166);
and U1758 (N_1758,In_829,N_724);
or U1759 (N_1759,N_1063,N_1143);
or U1760 (N_1760,N_527,N_681);
nor U1761 (N_1761,N_715,N_98);
or U1762 (N_1762,N_1151,N_631);
or U1763 (N_1763,In_1463,N_888);
xnor U1764 (N_1764,N_148,N_1185);
nor U1765 (N_1765,N_675,N_765);
and U1766 (N_1766,N_691,In_2231);
and U1767 (N_1767,In_1892,N_1114);
or U1768 (N_1768,N_913,In_1242);
nor U1769 (N_1769,N_1235,N_218);
or U1770 (N_1770,In_867,N_697);
and U1771 (N_1771,N_664,N_297);
or U1772 (N_1772,N_730,N_705);
nor U1773 (N_1773,In_1114,N_1068);
or U1774 (N_1774,In_2238,N_975);
or U1775 (N_1775,In_849,In_1548);
nand U1776 (N_1776,N_692,In_1008);
or U1777 (N_1777,N_864,N_657);
nand U1778 (N_1778,N_811,N_883);
nand U1779 (N_1779,N_797,In_2188);
and U1780 (N_1780,In_314,In_1668);
nor U1781 (N_1781,In_538,N_684);
or U1782 (N_1782,N_1159,N_973);
nor U1783 (N_1783,N_1249,In_1706);
or U1784 (N_1784,N_919,N_679);
xnor U1785 (N_1785,N_282,N_1147);
or U1786 (N_1786,N_1064,In_1974);
nand U1787 (N_1787,N_1088,N_808);
xor U1788 (N_1788,N_719,In_27);
nor U1789 (N_1789,In_1396,N_1028);
nand U1790 (N_1790,N_967,In_238);
or U1791 (N_1791,N_1234,N_1116);
and U1792 (N_1792,N_1096,In_1015);
nand U1793 (N_1793,In_1281,N_293);
nand U1794 (N_1794,N_1150,N_762);
nor U1795 (N_1795,N_1014,N_876);
nand U1796 (N_1796,N_989,In_336);
xnor U1797 (N_1797,N_298,In_475);
or U1798 (N_1798,N_1104,In_80);
nand U1799 (N_1799,N_80,N_1173);
or U1800 (N_1800,N_1016,In_937);
nand U1801 (N_1801,In_509,N_168);
and U1802 (N_1802,N_1025,N_43);
xnor U1803 (N_1803,In_316,In_1250);
nand U1804 (N_1804,N_1060,N_1233);
xnor U1805 (N_1805,N_859,In_2003);
nor U1806 (N_1806,N_662,N_805);
and U1807 (N_1807,In_703,N_964);
nand U1808 (N_1808,N_577,N_1077);
and U1809 (N_1809,N_807,In_941);
xor U1810 (N_1810,N_1164,In_936);
xnor U1811 (N_1811,N_932,N_823);
or U1812 (N_1812,N_1043,N_840);
and U1813 (N_1813,N_1247,In_743);
nand U1814 (N_1814,In_2124,N_809);
nor U1815 (N_1815,N_754,In_576);
or U1816 (N_1816,N_6,In_1615);
nand U1817 (N_1817,In_5,N_784);
nand U1818 (N_1818,In_990,In_930);
or U1819 (N_1819,In_1787,N_1002);
and U1820 (N_1820,In_1756,N_922);
nor U1821 (N_1821,In_2091,N_654);
xnor U1822 (N_1822,N_1076,N_515);
nand U1823 (N_1823,In_1097,In_1504);
xnor U1824 (N_1824,N_306,N_1142);
or U1825 (N_1825,In_328,In_1417);
nand U1826 (N_1826,N_1122,N_761);
or U1827 (N_1827,N_884,In_1472);
xor U1828 (N_1828,In_1767,N_1168);
and U1829 (N_1829,In_1272,N_1169);
and U1830 (N_1830,In_1821,N_696);
nand U1831 (N_1831,N_782,N_142);
nand U1832 (N_1832,N_660,N_141);
or U1833 (N_1833,N_433,N_655);
nand U1834 (N_1834,N_790,N_1061);
nand U1835 (N_1835,N_850,N_1087);
or U1836 (N_1836,N_1137,In_1958);
and U1837 (N_1837,N_887,N_786);
nand U1838 (N_1838,N_183,In_2071);
and U1839 (N_1839,In_711,N_601);
xnor U1840 (N_1840,N_787,In_410);
nand U1841 (N_1841,N_935,N_1203);
nand U1842 (N_1842,In_1255,N_729);
and U1843 (N_1843,N_773,N_1113);
and U1844 (N_1844,N_806,N_454);
xor U1845 (N_1845,N_867,N_440);
or U1846 (N_1846,N_774,In_1688);
or U1847 (N_1847,In_1109,In_1573);
nor U1848 (N_1848,N_241,In_2276);
xnor U1849 (N_1849,N_862,N_646);
or U1850 (N_1850,N_943,In_2248);
xnor U1851 (N_1851,N_53,N_1178);
and U1852 (N_1852,N_1039,N_653);
nand U1853 (N_1853,N_1001,N_632);
and U1854 (N_1854,N_961,N_860);
and U1855 (N_1855,N_1031,In_2103);
nor U1856 (N_1856,In_1371,N_1163);
or U1857 (N_1857,N_758,N_1012);
and U1858 (N_1858,In_679,N_738);
nand U1859 (N_1859,N_708,N_661);
nor U1860 (N_1860,N_1019,N_182);
and U1861 (N_1861,N_361,N_725);
and U1862 (N_1862,In_1770,In_1641);
xnor U1863 (N_1863,N_674,In_1174);
nand U1864 (N_1864,N_950,N_958);
nor U1865 (N_1865,N_1240,N_1171);
and U1866 (N_1866,N_1042,N_1000);
nand U1867 (N_1867,In_864,In_970);
nand U1868 (N_1868,N_1111,In_832);
nand U1869 (N_1869,In_2226,N_384);
xnor U1870 (N_1870,N_978,In_695);
or U1871 (N_1871,N_1103,In_365);
and U1872 (N_1872,N_1220,In_1849);
nor U1873 (N_1873,In_205,N_644);
or U1874 (N_1874,In_2482,In_1303);
and U1875 (N_1875,N_1252,N_1497);
xnor U1876 (N_1876,N_1477,N_1427);
nand U1877 (N_1877,N_1370,N_1860);
nor U1878 (N_1878,N_1544,N_1369);
xnor U1879 (N_1879,N_1396,N_1290);
nor U1880 (N_1880,N_1743,N_1635);
nor U1881 (N_1881,N_1400,N_1853);
and U1882 (N_1882,N_1298,N_1613);
xor U1883 (N_1883,N_1271,N_1593);
xor U1884 (N_1884,N_1414,N_1406);
nor U1885 (N_1885,N_1817,N_1456);
and U1886 (N_1886,N_1655,N_1380);
nand U1887 (N_1887,N_1728,N_1539);
or U1888 (N_1888,N_1818,N_1630);
and U1889 (N_1889,N_1831,N_1717);
nor U1890 (N_1890,N_1779,N_1789);
xor U1891 (N_1891,N_1736,N_1698);
xor U1892 (N_1892,N_1425,N_1337);
nor U1893 (N_1893,N_1725,N_1361);
nand U1894 (N_1894,N_1807,N_1714);
nor U1895 (N_1895,N_1352,N_1318);
or U1896 (N_1896,N_1602,N_1854);
xor U1897 (N_1897,N_1546,N_1598);
nand U1898 (N_1898,N_1504,N_1667);
and U1899 (N_1899,N_1757,N_1604);
or U1900 (N_1900,N_1267,N_1439);
nor U1901 (N_1901,N_1769,N_1798);
or U1902 (N_1902,N_1569,N_1381);
xnor U1903 (N_1903,N_1773,N_1761);
nand U1904 (N_1904,N_1415,N_1550);
or U1905 (N_1905,N_1741,N_1416);
xnor U1906 (N_1906,N_1649,N_1404);
xnor U1907 (N_1907,N_1850,N_1264);
and U1908 (N_1908,N_1484,N_1537);
or U1909 (N_1909,N_1745,N_1557);
xnor U1910 (N_1910,N_1475,N_1579);
or U1911 (N_1911,N_1302,N_1658);
or U1912 (N_1912,N_1827,N_1446);
or U1913 (N_1913,N_1314,N_1357);
nor U1914 (N_1914,N_1813,N_1841);
nor U1915 (N_1915,N_1481,N_1444);
or U1916 (N_1916,N_1382,N_1363);
nand U1917 (N_1917,N_1344,N_1268);
xor U1918 (N_1918,N_1830,N_1601);
xor U1919 (N_1919,N_1677,N_1781);
xor U1920 (N_1920,N_1760,N_1388);
nor U1921 (N_1921,N_1723,N_1608);
or U1922 (N_1922,N_1636,N_1589);
nand U1923 (N_1923,N_1258,N_1826);
and U1924 (N_1924,N_1345,N_1808);
nor U1925 (N_1925,N_1595,N_1863);
xor U1926 (N_1926,N_1772,N_1413);
nor U1927 (N_1927,N_1606,N_1324);
or U1928 (N_1928,N_1403,N_1842);
nor U1929 (N_1929,N_1701,N_1681);
or U1930 (N_1930,N_1751,N_1801);
xor U1931 (N_1931,N_1639,N_1583);
and U1932 (N_1932,N_1443,N_1257);
xnor U1933 (N_1933,N_1800,N_1263);
and U1934 (N_1934,N_1836,N_1855);
nand U1935 (N_1935,N_1699,N_1847);
nor U1936 (N_1936,N_1351,N_1837);
nand U1937 (N_1937,N_1542,N_1768);
nand U1938 (N_1938,N_1488,N_1685);
xnor U1939 (N_1939,N_1684,N_1501);
and U1940 (N_1940,N_1748,N_1561);
xnor U1941 (N_1941,N_1350,N_1543);
and U1942 (N_1942,N_1430,N_1311);
or U1943 (N_1943,N_1647,N_1587);
and U1944 (N_1944,N_1300,N_1678);
xor U1945 (N_1945,N_1642,N_1829);
nor U1946 (N_1946,N_1700,N_1548);
or U1947 (N_1947,N_1646,N_1291);
xnor U1948 (N_1948,N_1765,N_1766);
nor U1949 (N_1949,N_1422,N_1609);
and U1950 (N_1950,N_1463,N_1449);
or U1951 (N_1951,N_1605,N_1839);
nand U1952 (N_1952,N_1571,N_1355);
and U1953 (N_1953,N_1848,N_1358);
nand U1954 (N_1954,N_1686,N_1653);
and U1955 (N_1955,N_1657,N_1336);
xnor U1956 (N_1956,N_1553,N_1412);
and U1957 (N_1957,N_1669,N_1820);
nand U1958 (N_1958,N_1372,N_1424);
xor U1959 (N_1959,N_1476,N_1517);
or U1960 (N_1960,N_1465,N_1624);
or U1961 (N_1961,N_1260,N_1718);
xor U1962 (N_1962,N_1832,N_1662);
or U1963 (N_1963,N_1523,N_1573);
nor U1964 (N_1964,N_1467,N_1767);
and U1965 (N_1965,N_1762,N_1423);
xor U1966 (N_1966,N_1399,N_1865);
or U1967 (N_1967,N_1323,N_1474);
or U1968 (N_1968,N_1558,N_1472);
or U1969 (N_1969,N_1277,N_1692);
nor U1970 (N_1970,N_1656,N_1627);
nand U1971 (N_1971,N_1821,N_1572);
and U1972 (N_1972,N_1868,N_1334);
nand U1973 (N_1973,N_1375,N_1721);
or U1974 (N_1974,N_1815,N_1834);
and U1975 (N_1975,N_1659,N_1331);
nor U1976 (N_1976,N_1788,N_1280);
or U1977 (N_1977,N_1308,N_1417);
xnor U1978 (N_1978,N_1274,N_1575);
and U1979 (N_1979,N_1644,N_1509);
or U1980 (N_1980,N_1521,N_1451);
nor U1981 (N_1981,N_1459,N_1464);
or U1982 (N_1982,N_1862,N_1531);
nand U1983 (N_1983,N_1840,N_1724);
nand U1984 (N_1984,N_1784,N_1590);
and U1985 (N_1985,N_1554,N_1420);
xnor U1986 (N_1986,N_1356,N_1460);
nor U1987 (N_1987,N_1709,N_1733);
and U1988 (N_1988,N_1565,N_1809);
xnor U1989 (N_1989,N_1547,N_1645);
and U1990 (N_1990,N_1683,N_1637);
or U1991 (N_1991,N_1578,N_1833);
nand U1992 (N_1992,N_1785,N_1435);
nor U1993 (N_1993,N_1397,N_1253);
or U1994 (N_1994,N_1391,N_1442);
and U1995 (N_1995,N_1858,N_1694);
xnor U1996 (N_1996,N_1259,N_1514);
or U1997 (N_1997,N_1401,N_1874);
or U1998 (N_1998,N_1690,N_1266);
nor U1999 (N_1999,N_1688,N_1480);
nor U2000 (N_2000,N_1254,N_1433);
or U2001 (N_2001,N_1262,N_1675);
nand U2002 (N_2002,N_1511,N_1279);
nor U2003 (N_2003,N_1434,N_1385);
and U2004 (N_2004,N_1735,N_1510);
xor U2005 (N_2005,N_1545,N_1742);
nor U2006 (N_2006,N_1533,N_1654);
or U2007 (N_2007,N_1462,N_1270);
and U2008 (N_2008,N_1555,N_1367);
nand U2009 (N_2009,N_1261,N_1486);
nor U2010 (N_2010,N_1586,N_1679);
nor U2011 (N_2011,N_1696,N_1431);
or U2012 (N_2012,N_1440,N_1774);
nor U2013 (N_2013,N_1339,N_1532);
and U2014 (N_2014,N_1770,N_1756);
and U2015 (N_2015,N_1373,N_1626);
and U2016 (N_2016,N_1607,N_1814);
or U2017 (N_2017,N_1771,N_1625);
nand U2018 (N_2018,N_1332,N_1568);
xnor U2019 (N_2019,N_1780,N_1612);
and U2020 (N_2020,N_1461,N_1597);
and U2021 (N_2021,N_1719,N_1529);
or U2022 (N_2022,N_1371,N_1740);
or U2023 (N_2023,N_1284,N_1468);
nor U2024 (N_2024,N_1652,N_1661);
and U2025 (N_2025,N_1835,N_1294);
nand U2026 (N_2026,N_1870,N_1507);
nor U2027 (N_2027,N_1343,N_1628);
or U2028 (N_2028,N_1845,N_1864);
xnor U2029 (N_2029,N_1487,N_1594);
nand U2030 (N_2030,N_1347,N_1303);
xor U2031 (N_2031,N_1411,N_1445);
and U2032 (N_2032,N_1287,N_1438);
nand U2033 (N_2033,N_1713,N_1640);
xnor U2034 (N_2034,N_1436,N_1641);
or U2035 (N_2035,N_1856,N_1377);
nor U2036 (N_2036,N_1429,N_1787);
nor U2037 (N_2037,N_1410,N_1275);
nand U2038 (N_2038,N_1540,N_1360);
or U2039 (N_2039,N_1710,N_1421);
and U2040 (N_2040,N_1705,N_1794);
and U2041 (N_2041,N_1552,N_1492);
and U2042 (N_2042,N_1499,N_1493);
and U2043 (N_2043,N_1738,N_1668);
xor U2044 (N_2044,N_1392,N_1320);
nor U2045 (N_2045,N_1322,N_1764);
xor U2046 (N_2046,N_1538,N_1691);
nand U2047 (N_2047,N_1793,N_1731);
or U2048 (N_2048,N_1365,N_1824);
nor U2049 (N_2049,N_1567,N_1873);
or U2050 (N_2050,N_1516,N_1680);
nor U2051 (N_2051,N_1620,N_1674);
nor U2052 (N_2052,N_1282,N_1610);
xor U2053 (N_2053,N_1621,N_1432);
xor U2054 (N_2054,N_1374,N_1469);
and U2055 (N_2055,N_1273,N_1796);
xnor U2056 (N_2056,N_1285,N_1697);
and U2057 (N_2057,N_1328,N_1634);
nand U2058 (N_2058,N_1600,N_1763);
nand U2059 (N_2059,N_1269,N_1671);
and U2060 (N_2060,N_1295,N_1797);
or U2061 (N_2061,N_1478,N_1502);
xor U2062 (N_2062,N_1506,N_1470);
or U2063 (N_2063,N_1576,N_1292);
nand U2064 (N_2064,N_1265,N_1250);
and U2065 (N_2065,N_1305,N_1408);
or U2066 (N_2066,N_1489,N_1580);
xor U2067 (N_2067,N_1663,N_1739);
nand U2068 (N_2068,N_1524,N_1255);
and U2069 (N_2069,N_1485,N_1682);
and U2070 (N_2070,N_1660,N_1618);
and U2071 (N_2071,N_1353,N_1389);
xor U2072 (N_2072,N_1526,N_1729);
or U2073 (N_2073,N_1378,N_1689);
and U2074 (N_2074,N_1490,N_1437);
nand U2075 (N_2075,N_1251,N_1278);
and U2076 (N_2076,N_1466,N_1619);
nor U2077 (N_2077,N_1455,N_1299);
nor U2078 (N_2078,N_1491,N_1326);
nor U2079 (N_2079,N_1732,N_1843);
or U2080 (N_2080,N_1319,N_1665);
and U2081 (N_2081,N_1289,N_1549);
and U2082 (N_2082,N_1327,N_1670);
nor U2083 (N_2083,N_1819,N_1338);
and U2084 (N_2084,N_1712,N_1457);
and U2085 (N_2085,N_1726,N_1498);
and U2086 (N_2086,N_1707,N_1711);
or U2087 (N_2087,N_1321,N_1276);
nand U2088 (N_2088,N_1823,N_1428);
nor U2089 (N_2089,N_1615,N_1746);
and U2090 (N_2090,N_1359,N_1500);
and U2091 (N_2091,N_1846,N_1816);
nand U2092 (N_2092,N_1599,N_1368);
or U2093 (N_2093,N_1851,N_1702);
nor U2094 (N_2094,N_1281,N_1584);
and U2095 (N_2095,N_1483,N_1309);
or U2096 (N_2096,N_1560,N_1301);
xor U2097 (N_2097,N_1825,N_1782);
nand U2098 (N_2098,N_1857,N_1582);
nand U2099 (N_2099,N_1349,N_1452);
or U2100 (N_2100,N_1342,N_1871);
nor U2101 (N_2101,N_1304,N_1570);
xor U2102 (N_2102,N_1448,N_1852);
or U2103 (N_2103,N_1563,N_1631);
nand U2104 (N_2104,N_1454,N_1795);
xor U2105 (N_2105,N_1664,N_1828);
and U2106 (N_2106,N_1325,N_1307);
nand U2107 (N_2107,N_1426,N_1716);
or U2108 (N_2108,N_1783,N_1346);
and U2109 (N_2109,N_1758,N_1394);
nand U2110 (N_2110,N_1384,N_1643);
nor U2111 (N_2111,N_1390,N_1799);
or U2112 (N_2112,N_1747,N_1737);
xor U2113 (N_2113,N_1706,N_1859);
nor U2114 (N_2114,N_1804,N_1838);
or U2115 (N_2115,N_1530,N_1727);
and U2116 (N_2116,N_1722,N_1534);
xor U2117 (N_2117,N_1447,N_1541);
or U2118 (N_2118,N_1503,N_1775);
xnor U2119 (N_2119,N_1348,N_1849);
nor U2120 (N_2120,N_1810,N_1383);
or U2121 (N_2121,N_1450,N_1759);
nand U2122 (N_2122,N_1617,N_1512);
and U2123 (N_2123,N_1364,N_1708);
and U2124 (N_2124,N_1869,N_1622);
xnor U2125 (N_2125,N_1296,N_1293);
and U2126 (N_2126,N_1693,N_1528);
xor U2127 (N_2127,N_1398,N_1333);
xor U2128 (N_2128,N_1754,N_1536);
or U2129 (N_2129,N_1844,N_1519);
or U2130 (N_2130,N_1687,N_1297);
xor U2131 (N_2131,N_1395,N_1603);
nand U2132 (N_2132,N_1419,N_1715);
or U2133 (N_2133,N_1402,N_1376);
nor U2134 (N_2134,N_1564,N_1473);
and U2135 (N_2135,N_1458,N_1340);
and U2136 (N_2136,N_1496,N_1790);
nand U2137 (N_2137,N_1632,N_1409);
nand U2138 (N_2138,N_1574,N_1518);
nor U2139 (N_2139,N_1577,N_1777);
and U2140 (N_2140,N_1744,N_1866);
xnor U2141 (N_2141,N_1592,N_1453);
nor U2142 (N_2142,N_1676,N_1792);
and U2143 (N_2143,N_1272,N_1312);
nor U2144 (N_2144,N_1527,N_1651);
and U2145 (N_2145,N_1581,N_1556);
and U2146 (N_2146,N_1805,N_1330);
nor U2147 (N_2147,N_1749,N_1335);
nand U2148 (N_2148,N_1525,N_1317);
and U2149 (N_2149,N_1776,N_1672);
and U2150 (N_2150,N_1791,N_1703);
and U2151 (N_2151,N_1316,N_1585);
or U2152 (N_2152,N_1362,N_1614);
and U2153 (N_2153,N_1306,N_1666);
xnor U2154 (N_2154,N_1386,N_1822);
nor U2155 (N_2155,N_1379,N_1811);
nand U2156 (N_2156,N_1734,N_1495);
xnor U2157 (N_2157,N_1623,N_1616);
nand U2158 (N_2158,N_1867,N_1535);
and U2159 (N_2159,N_1752,N_1720);
and U2160 (N_2160,N_1633,N_1418);
and U2161 (N_2161,N_1482,N_1559);
or U2162 (N_2162,N_1611,N_1315);
and U2163 (N_2163,N_1508,N_1313);
or U2164 (N_2164,N_1522,N_1704);
nand U2165 (N_2165,N_1566,N_1650);
nand U2166 (N_2166,N_1520,N_1812);
and U2167 (N_2167,N_1393,N_1872);
xor U2168 (N_2168,N_1286,N_1673);
and U2169 (N_2169,N_1778,N_1588);
xnor U2170 (N_2170,N_1479,N_1802);
or U2171 (N_2171,N_1730,N_1354);
nand U2172 (N_2172,N_1755,N_1648);
and U2173 (N_2173,N_1310,N_1629);
nand U2174 (N_2174,N_1471,N_1329);
and U2175 (N_2175,N_1515,N_1505);
xor U2176 (N_2176,N_1405,N_1256);
nand U2177 (N_2177,N_1806,N_1551);
nor U2178 (N_2178,N_1786,N_1753);
and U2179 (N_2179,N_1366,N_1441);
and U2180 (N_2180,N_1638,N_1695);
or U2181 (N_2181,N_1288,N_1513);
and U2182 (N_2182,N_1387,N_1407);
or U2183 (N_2183,N_1861,N_1283);
or U2184 (N_2184,N_1750,N_1803);
xor U2185 (N_2185,N_1596,N_1494);
or U2186 (N_2186,N_1341,N_1591);
nand U2187 (N_2187,N_1562,N_1539);
nor U2188 (N_2188,N_1485,N_1442);
or U2189 (N_2189,N_1498,N_1353);
nand U2190 (N_2190,N_1510,N_1297);
xor U2191 (N_2191,N_1610,N_1296);
xor U2192 (N_2192,N_1814,N_1304);
nor U2193 (N_2193,N_1416,N_1473);
and U2194 (N_2194,N_1393,N_1513);
xnor U2195 (N_2195,N_1700,N_1715);
nor U2196 (N_2196,N_1834,N_1701);
nor U2197 (N_2197,N_1813,N_1719);
nor U2198 (N_2198,N_1276,N_1636);
nand U2199 (N_2199,N_1866,N_1386);
xor U2200 (N_2200,N_1648,N_1382);
xor U2201 (N_2201,N_1351,N_1605);
or U2202 (N_2202,N_1318,N_1625);
nor U2203 (N_2203,N_1679,N_1834);
xor U2204 (N_2204,N_1314,N_1373);
xor U2205 (N_2205,N_1579,N_1348);
or U2206 (N_2206,N_1300,N_1551);
nand U2207 (N_2207,N_1803,N_1776);
or U2208 (N_2208,N_1502,N_1265);
nand U2209 (N_2209,N_1438,N_1503);
and U2210 (N_2210,N_1851,N_1365);
and U2211 (N_2211,N_1292,N_1862);
or U2212 (N_2212,N_1674,N_1360);
nand U2213 (N_2213,N_1361,N_1291);
or U2214 (N_2214,N_1321,N_1481);
xor U2215 (N_2215,N_1786,N_1511);
nand U2216 (N_2216,N_1376,N_1783);
and U2217 (N_2217,N_1510,N_1326);
and U2218 (N_2218,N_1859,N_1707);
nor U2219 (N_2219,N_1830,N_1565);
nor U2220 (N_2220,N_1314,N_1847);
or U2221 (N_2221,N_1579,N_1797);
xor U2222 (N_2222,N_1436,N_1279);
and U2223 (N_2223,N_1682,N_1841);
nor U2224 (N_2224,N_1734,N_1745);
or U2225 (N_2225,N_1750,N_1432);
nor U2226 (N_2226,N_1456,N_1427);
and U2227 (N_2227,N_1323,N_1711);
and U2228 (N_2228,N_1275,N_1363);
nand U2229 (N_2229,N_1341,N_1560);
or U2230 (N_2230,N_1446,N_1864);
nor U2231 (N_2231,N_1444,N_1301);
xor U2232 (N_2232,N_1466,N_1829);
nand U2233 (N_2233,N_1686,N_1605);
or U2234 (N_2234,N_1796,N_1746);
and U2235 (N_2235,N_1788,N_1590);
nor U2236 (N_2236,N_1722,N_1322);
xor U2237 (N_2237,N_1504,N_1729);
nor U2238 (N_2238,N_1829,N_1698);
or U2239 (N_2239,N_1261,N_1516);
nor U2240 (N_2240,N_1795,N_1317);
nor U2241 (N_2241,N_1359,N_1796);
and U2242 (N_2242,N_1397,N_1325);
nand U2243 (N_2243,N_1786,N_1287);
nand U2244 (N_2244,N_1736,N_1411);
and U2245 (N_2245,N_1641,N_1833);
nor U2246 (N_2246,N_1442,N_1659);
xnor U2247 (N_2247,N_1394,N_1815);
and U2248 (N_2248,N_1542,N_1660);
nand U2249 (N_2249,N_1665,N_1710);
nor U2250 (N_2250,N_1820,N_1672);
xor U2251 (N_2251,N_1674,N_1393);
or U2252 (N_2252,N_1401,N_1839);
xnor U2253 (N_2253,N_1758,N_1769);
xnor U2254 (N_2254,N_1409,N_1359);
nand U2255 (N_2255,N_1355,N_1837);
or U2256 (N_2256,N_1560,N_1736);
nor U2257 (N_2257,N_1817,N_1576);
or U2258 (N_2258,N_1725,N_1327);
and U2259 (N_2259,N_1426,N_1836);
nor U2260 (N_2260,N_1474,N_1652);
nand U2261 (N_2261,N_1355,N_1699);
xor U2262 (N_2262,N_1753,N_1737);
xor U2263 (N_2263,N_1788,N_1265);
xnor U2264 (N_2264,N_1268,N_1707);
nand U2265 (N_2265,N_1600,N_1873);
nand U2266 (N_2266,N_1489,N_1298);
xor U2267 (N_2267,N_1552,N_1645);
nand U2268 (N_2268,N_1470,N_1365);
nor U2269 (N_2269,N_1375,N_1820);
xor U2270 (N_2270,N_1456,N_1288);
nand U2271 (N_2271,N_1468,N_1641);
and U2272 (N_2272,N_1733,N_1840);
nor U2273 (N_2273,N_1307,N_1697);
nor U2274 (N_2274,N_1253,N_1507);
nor U2275 (N_2275,N_1410,N_1293);
nand U2276 (N_2276,N_1485,N_1622);
nor U2277 (N_2277,N_1810,N_1704);
nor U2278 (N_2278,N_1528,N_1802);
nor U2279 (N_2279,N_1868,N_1670);
nand U2280 (N_2280,N_1506,N_1458);
xor U2281 (N_2281,N_1739,N_1559);
and U2282 (N_2282,N_1665,N_1566);
nor U2283 (N_2283,N_1403,N_1567);
xor U2284 (N_2284,N_1528,N_1697);
nor U2285 (N_2285,N_1634,N_1348);
nor U2286 (N_2286,N_1852,N_1488);
and U2287 (N_2287,N_1781,N_1377);
nand U2288 (N_2288,N_1415,N_1427);
or U2289 (N_2289,N_1822,N_1437);
or U2290 (N_2290,N_1554,N_1857);
nor U2291 (N_2291,N_1566,N_1570);
nand U2292 (N_2292,N_1425,N_1420);
nor U2293 (N_2293,N_1613,N_1692);
xor U2294 (N_2294,N_1473,N_1841);
and U2295 (N_2295,N_1751,N_1452);
nor U2296 (N_2296,N_1478,N_1677);
and U2297 (N_2297,N_1530,N_1762);
xnor U2298 (N_2298,N_1547,N_1355);
nor U2299 (N_2299,N_1549,N_1445);
nor U2300 (N_2300,N_1544,N_1868);
xnor U2301 (N_2301,N_1665,N_1535);
and U2302 (N_2302,N_1407,N_1566);
nand U2303 (N_2303,N_1291,N_1627);
xnor U2304 (N_2304,N_1806,N_1474);
nand U2305 (N_2305,N_1254,N_1394);
xnor U2306 (N_2306,N_1485,N_1455);
nor U2307 (N_2307,N_1852,N_1764);
and U2308 (N_2308,N_1391,N_1808);
nand U2309 (N_2309,N_1540,N_1438);
nand U2310 (N_2310,N_1395,N_1262);
xnor U2311 (N_2311,N_1256,N_1513);
and U2312 (N_2312,N_1302,N_1651);
nand U2313 (N_2313,N_1453,N_1372);
nor U2314 (N_2314,N_1421,N_1486);
nor U2315 (N_2315,N_1690,N_1705);
or U2316 (N_2316,N_1272,N_1732);
nor U2317 (N_2317,N_1743,N_1820);
nand U2318 (N_2318,N_1259,N_1598);
nor U2319 (N_2319,N_1741,N_1392);
xnor U2320 (N_2320,N_1507,N_1333);
or U2321 (N_2321,N_1656,N_1801);
and U2322 (N_2322,N_1300,N_1799);
nand U2323 (N_2323,N_1438,N_1596);
and U2324 (N_2324,N_1484,N_1836);
or U2325 (N_2325,N_1440,N_1715);
and U2326 (N_2326,N_1253,N_1821);
and U2327 (N_2327,N_1853,N_1466);
xnor U2328 (N_2328,N_1582,N_1555);
or U2329 (N_2329,N_1650,N_1668);
nand U2330 (N_2330,N_1780,N_1586);
or U2331 (N_2331,N_1432,N_1602);
nand U2332 (N_2332,N_1414,N_1255);
nand U2333 (N_2333,N_1666,N_1673);
and U2334 (N_2334,N_1462,N_1411);
xnor U2335 (N_2335,N_1834,N_1588);
xor U2336 (N_2336,N_1364,N_1637);
nor U2337 (N_2337,N_1428,N_1733);
nor U2338 (N_2338,N_1434,N_1620);
nand U2339 (N_2339,N_1288,N_1735);
xor U2340 (N_2340,N_1539,N_1748);
nand U2341 (N_2341,N_1577,N_1778);
nor U2342 (N_2342,N_1568,N_1870);
and U2343 (N_2343,N_1251,N_1411);
and U2344 (N_2344,N_1343,N_1810);
nor U2345 (N_2345,N_1430,N_1463);
and U2346 (N_2346,N_1652,N_1696);
xnor U2347 (N_2347,N_1482,N_1830);
and U2348 (N_2348,N_1293,N_1746);
or U2349 (N_2349,N_1694,N_1667);
and U2350 (N_2350,N_1288,N_1530);
nand U2351 (N_2351,N_1368,N_1557);
nor U2352 (N_2352,N_1581,N_1418);
nand U2353 (N_2353,N_1642,N_1359);
or U2354 (N_2354,N_1512,N_1412);
xor U2355 (N_2355,N_1673,N_1707);
nand U2356 (N_2356,N_1737,N_1733);
nor U2357 (N_2357,N_1517,N_1865);
xor U2358 (N_2358,N_1672,N_1437);
or U2359 (N_2359,N_1540,N_1350);
and U2360 (N_2360,N_1365,N_1253);
and U2361 (N_2361,N_1749,N_1538);
nor U2362 (N_2362,N_1816,N_1791);
nand U2363 (N_2363,N_1314,N_1764);
or U2364 (N_2364,N_1712,N_1301);
nand U2365 (N_2365,N_1508,N_1703);
and U2366 (N_2366,N_1658,N_1833);
nor U2367 (N_2367,N_1317,N_1758);
nor U2368 (N_2368,N_1629,N_1838);
or U2369 (N_2369,N_1616,N_1505);
nand U2370 (N_2370,N_1522,N_1319);
xor U2371 (N_2371,N_1453,N_1832);
nor U2372 (N_2372,N_1609,N_1610);
and U2373 (N_2373,N_1682,N_1550);
xor U2374 (N_2374,N_1617,N_1851);
xor U2375 (N_2375,N_1692,N_1870);
nor U2376 (N_2376,N_1465,N_1333);
nand U2377 (N_2377,N_1691,N_1476);
xnor U2378 (N_2378,N_1820,N_1685);
xor U2379 (N_2379,N_1661,N_1354);
nand U2380 (N_2380,N_1864,N_1325);
and U2381 (N_2381,N_1257,N_1381);
or U2382 (N_2382,N_1870,N_1585);
xnor U2383 (N_2383,N_1258,N_1553);
or U2384 (N_2384,N_1392,N_1848);
nor U2385 (N_2385,N_1382,N_1512);
nand U2386 (N_2386,N_1680,N_1779);
or U2387 (N_2387,N_1657,N_1498);
or U2388 (N_2388,N_1303,N_1336);
nor U2389 (N_2389,N_1594,N_1853);
xor U2390 (N_2390,N_1723,N_1390);
and U2391 (N_2391,N_1530,N_1477);
xor U2392 (N_2392,N_1670,N_1825);
nand U2393 (N_2393,N_1360,N_1536);
nor U2394 (N_2394,N_1823,N_1377);
nand U2395 (N_2395,N_1835,N_1435);
nand U2396 (N_2396,N_1517,N_1873);
nand U2397 (N_2397,N_1338,N_1639);
or U2398 (N_2398,N_1817,N_1721);
xnor U2399 (N_2399,N_1802,N_1728);
or U2400 (N_2400,N_1303,N_1828);
and U2401 (N_2401,N_1713,N_1806);
and U2402 (N_2402,N_1326,N_1530);
and U2403 (N_2403,N_1576,N_1540);
xor U2404 (N_2404,N_1831,N_1429);
nand U2405 (N_2405,N_1355,N_1469);
xor U2406 (N_2406,N_1265,N_1867);
xor U2407 (N_2407,N_1407,N_1586);
nor U2408 (N_2408,N_1874,N_1722);
and U2409 (N_2409,N_1262,N_1722);
or U2410 (N_2410,N_1874,N_1645);
nand U2411 (N_2411,N_1523,N_1606);
and U2412 (N_2412,N_1795,N_1343);
or U2413 (N_2413,N_1488,N_1421);
nand U2414 (N_2414,N_1507,N_1764);
nor U2415 (N_2415,N_1684,N_1622);
nor U2416 (N_2416,N_1536,N_1683);
nand U2417 (N_2417,N_1800,N_1648);
or U2418 (N_2418,N_1538,N_1641);
xor U2419 (N_2419,N_1706,N_1517);
xor U2420 (N_2420,N_1440,N_1485);
nor U2421 (N_2421,N_1821,N_1322);
or U2422 (N_2422,N_1449,N_1680);
nor U2423 (N_2423,N_1370,N_1854);
nand U2424 (N_2424,N_1698,N_1508);
or U2425 (N_2425,N_1783,N_1630);
nand U2426 (N_2426,N_1374,N_1849);
and U2427 (N_2427,N_1503,N_1462);
nand U2428 (N_2428,N_1669,N_1456);
nand U2429 (N_2429,N_1808,N_1650);
xor U2430 (N_2430,N_1798,N_1459);
nor U2431 (N_2431,N_1617,N_1331);
and U2432 (N_2432,N_1555,N_1627);
nand U2433 (N_2433,N_1597,N_1754);
and U2434 (N_2434,N_1735,N_1468);
xor U2435 (N_2435,N_1533,N_1261);
xnor U2436 (N_2436,N_1436,N_1713);
nand U2437 (N_2437,N_1284,N_1624);
or U2438 (N_2438,N_1510,N_1540);
and U2439 (N_2439,N_1273,N_1468);
nor U2440 (N_2440,N_1662,N_1400);
and U2441 (N_2441,N_1828,N_1460);
xnor U2442 (N_2442,N_1785,N_1797);
nand U2443 (N_2443,N_1524,N_1865);
or U2444 (N_2444,N_1606,N_1443);
nor U2445 (N_2445,N_1649,N_1322);
nor U2446 (N_2446,N_1353,N_1278);
xor U2447 (N_2447,N_1282,N_1263);
xor U2448 (N_2448,N_1639,N_1570);
and U2449 (N_2449,N_1767,N_1631);
and U2450 (N_2450,N_1869,N_1619);
xnor U2451 (N_2451,N_1459,N_1377);
nor U2452 (N_2452,N_1634,N_1460);
nor U2453 (N_2453,N_1722,N_1709);
or U2454 (N_2454,N_1286,N_1523);
nor U2455 (N_2455,N_1367,N_1527);
and U2456 (N_2456,N_1338,N_1623);
nand U2457 (N_2457,N_1831,N_1354);
or U2458 (N_2458,N_1435,N_1531);
xnor U2459 (N_2459,N_1425,N_1550);
xnor U2460 (N_2460,N_1351,N_1808);
nor U2461 (N_2461,N_1659,N_1846);
xor U2462 (N_2462,N_1801,N_1401);
xor U2463 (N_2463,N_1334,N_1756);
nor U2464 (N_2464,N_1811,N_1620);
or U2465 (N_2465,N_1472,N_1481);
or U2466 (N_2466,N_1623,N_1722);
and U2467 (N_2467,N_1779,N_1425);
or U2468 (N_2468,N_1699,N_1344);
or U2469 (N_2469,N_1305,N_1413);
nand U2470 (N_2470,N_1457,N_1793);
or U2471 (N_2471,N_1287,N_1683);
nand U2472 (N_2472,N_1543,N_1850);
nand U2473 (N_2473,N_1813,N_1754);
and U2474 (N_2474,N_1723,N_1456);
nand U2475 (N_2475,N_1733,N_1533);
or U2476 (N_2476,N_1458,N_1574);
nor U2477 (N_2477,N_1855,N_1370);
nor U2478 (N_2478,N_1749,N_1448);
nand U2479 (N_2479,N_1464,N_1585);
and U2480 (N_2480,N_1717,N_1405);
xor U2481 (N_2481,N_1453,N_1613);
xnor U2482 (N_2482,N_1679,N_1421);
nor U2483 (N_2483,N_1374,N_1653);
and U2484 (N_2484,N_1664,N_1861);
nand U2485 (N_2485,N_1853,N_1708);
or U2486 (N_2486,N_1553,N_1784);
nor U2487 (N_2487,N_1724,N_1720);
and U2488 (N_2488,N_1488,N_1455);
nand U2489 (N_2489,N_1485,N_1265);
nand U2490 (N_2490,N_1572,N_1534);
and U2491 (N_2491,N_1654,N_1759);
nor U2492 (N_2492,N_1805,N_1405);
or U2493 (N_2493,N_1860,N_1517);
or U2494 (N_2494,N_1506,N_1322);
xnor U2495 (N_2495,N_1819,N_1629);
or U2496 (N_2496,N_1604,N_1349);
or U2497 (N_2497,N_1820,N_1816);
xor U2498 (N_2498,N_1430,N_1468);
and U2499 (N_2499,N_1571,N_1712);
and U2500 (N_2500,N_2308,N_2107);
nand U2501 (N_2501,N_2353,N_2434);
nor U2502 (N_2502,N_2208,N_2478);
or U2503 (N_2503,N_2030,N_2426);
nor U2504 (N_2504,N_2130,N_2008);
nand U2505 (N_2505,N_1965,N_2165);
nor U2506 (N_2506,N_2329,N_2444);
nor U2507 (N_2507,N_2438,N_2479);
or U2508 (N_2508,N_2446,N_2418);
xnor U2509 (N_2509,N_1968,N_1910);
or U2510 (N_2510,N_1947,N_2455);
xnor U2511 (N_2511,N_1991,N_2183);
and U2512 (N_2512,N_2062,N_2201);
and U2513 (N_2513,N_2496,N_2382);
or U2514 (N_2514,N_2138,N_2487);
and U2515 (N_2515,N_2284,N_2139);
or U2516 (N_2516,N_2423,N_2300);
and U2517 (N_2517,N_2059,N_2070);
or U2518 (N_2518,N_2347,N_2217);
or U2519 (N_2519,N_2026,N_1894);
xnor U2520 (N_2520,N_2311,N_2095);
and U2521 (N_2521,N_2089,N_2274);
xnor U2522 (N_2522,N_1911,N_2228);
or U2523 (N_2523,N_2358,N_2072);
nor U2524 (N_2524,N_2482,N_1973);
nor U2525 (N_2525,N_1970,N_2331);
xnor U2526 (N_2526,N_2472,N_2024);
xor U2527 (N_2527,N_2133,N_2015);
xor U2528 (N_2528,N_2324,N_1901);
nor U2529 (N_2529,N_1898,N_2047);
and U2530 (N_2530,N_2330,N_2497);
nor U2531 (N_2531,N_2083,N_1932);
xor U2532 (N_2532,N_2129,N_2189);
nor U2533 (N_2533,N_2425,N_2099);
and U2534 (N_2534,N_2368,N_2086);
and U2535 (N_2535,N_2104,N_1888);
and U2536 (N_2536,N_2152,N_2112);
xnor U2537 (N_2537,N_2336,N_1889);
or U2538 (N_2538,N_2389,N_2388);
nand U2539 (N_2539,N_1939,N_2312);
xor U2540 (N_2540,N_2052,N_2454);
or U2541 (N_2541,N_2394,N_2279);
nor U2542 (N_2542,N_2204,N_2432);
and U2543 (N_2543,N_1950,N_1875);
or U2544 (N_2544,N_2441,N_2280);
xor U2545 (N_2545,N_2198,N_1885);
nand U2546 (N_2546,N_2137,N_2258);
nand U2547 (N_2547,N_2398,N_1995);
xnor U2548 (N_2548,N_2214,N_2465);
nand U2549 (N_2549,N_2163,N_2292);
and U2550 (N_2550,N_2436,N_2351);
nor U2551 (N_2551,N_2449,N_2209);
nor U2552 (N_2552,N_2117,N_1963);
or U2553 (N_2553,N_2064,N_2428);
or U2554 (N_2554,N_2241,N_2013);
xnor U2555 (N_2555,N_2158,N_2459);
xor U2556 (N_2556,N_1944,N_2169);
or U2557 (N_2557,N_2196,N_1907);
and U2558 (N_2558,N_2363,N_2076);
or U2559 (N_2559,N_2435,N_2273);
and U2560 (N_2560,N_1990,N_1892);
or U2561 (N_2561,N_2186,N_2345);
or U2562 (N_2562,N_2247,N_2451);
nand U2563 (N_2563,N_2249,N_2493);
or U2564 (N_2564,N_2342,N_2022);
or U2565 (N_2565,N_2243,N_2355);
nor U2566 (N_2566,N_2341,N_2275);
nor U2567 (N_2567,N_2227,N_2050);
nand U2568 (N_2568,N_2145,N_2039);
nor U2569 (N_2569,N_2021,N_2172);
xnor U2570 (N_2570,N_1940,N_2271);
nand U2571 (N_2571,N_2097,N_1976);
nand U2572 (N_2572,N_2126,N_2340);
xor U2573 (N_2573,N_2109,N_2309);
xor U2574 (N_2574,N_2159,N_2025);
xor U2575 (N_2575,N_2245,N_2409);
nand U2576 (N_2576,N_2365,N_2492);
nand U2577 (N_2577,N_2257,N_2301);
xnor U2578 (N_2578,N_2202,N_2289);
nor U2579 (N_2579,N_2181,N_1928);
and U2580 (N_2580,N_2298,N_2352);
xnor U2581 (N_2581,N_2113,N_1984);
xnor U2582 (N_2582,N_2185,N_2404);
nor U2583 (N_2583,N_1884,N_2297);
nor U2584 (N_2584,N_2458,N_2085);
and U2585 (N_2585,N_2223,N_1993);
nand U2586 (N_2586,N_2264,N_2461);
nor U2587 (N_2587,N_2171,N_2067);
and U2588 (N_2588,N_2002,N_2216);
nor U2589 (N_2589,N_2387,N_2147);
or U2590 (N_2590,N_2207,N_2043);
and U2591 (N_2591,N_2381,N_1877);
and U2592 (N_2592,N_2313,N_2157);
or U2593 (N_2593,N_2370,N_2038);
nand U2594 (N_2594,N_2422,N_2054);
or U2595 (N_2595,N_1997,N_2253);
nor U2596 (N_2596,N_1926,N_2287);
and U2597 (N_2597,N_2488,N_2176);
and U2598 (N_2598,N_1902,N_2489);
xor U2599 (N_2599,N_1903,N_2255);
nand U2600 (N_2600,N_2326,N_2069);
nor U2601 (N_2601,N_1977,N_2048);
and U2602 (N_2602,N_2001,N_2009);
xor U2603 (N_2603,N_2467,N_2178);
or U2604 (N_2604,N_1879,N_2403);
nor U2605 (N_2605,N_2037,N_1938);
and U2606 (N_2606,N_2131,N_2276);
nand U2607 (N_2607,N_2357,N_2266);
nor U2608 (N_2608,N_2491,N_1921);
and U2609 (N_2609,N_1943,N_1996);
or U2610 (N_2610,N_2079,N_2150);
or U2611 (N_2611,N_2018,N_2075);
or U2612 (N_2612,N_2246,N_2111);
xnor U2613 (N_2613,N_2173,N_2367);
nor U2614 (N_2614,N_2269,N_1908);
and U2615 (N_2615,N_2121,N_2058);
and U2616 (N_2616,N_2384,N_2195);
nand U2617 (N_2617,N_2203,N_2392);
xnor U2618 (N_2618,N_1953,N_2055);
xor U2619 (N_2619,N_2480,N_1880);
nor U2620 (N_2620,N_2304,N_1933);
nor U2621 (N_2621,N_1983,N_2260);
nor U2622 (N_2622,N_1952,N_2310);
or U2623 (N_2623,N_2302,N_2452);
and U2624 (N_2624,N_2374,N_2360);
or U2625 (N_2625,N_1899,N_2191);
xor U2626 (N_2626,N_2250,N_2221);
and U2627 (N_2627,N_2366,N_2102);
nor U2628 (N_2628,N_2386,N_1958);
nor U2629 (N_2629,N_2061,N_2453);
and U2630 (N_2630,N_2262,N_2421);
or U2631 (N_2631,N_2164,N_2268);
or U2632 (N_2632,N_2475,N_2407);
nand U2633 (N_2633,N_2463,N_2256);
nor U2634 (N_2634,N_2417,N_2125);
or U2635 (N_2635,N_2031,N_2495);
xnor U2636 (N_2636,N_2232,N_1915);
xor U2637 (N_2637,N_2115,N_2020);
nand U2638 (N_2638,N_2393,N_2252);
or U2639 (N_2639,N_2141,N_1917);
and U2640 (N_2640,N_1900,N_2242);
and U2641 (N_2641,N_2041,N_2476);
and U2642 (N_2642,N_2044,N_2071);
and U2643 (N_2643,N_2328,N_2019);
xor U2644 (N_2644,N_1951,N_2212);
nor U2645 (N_2645,N_2205,N_1955);
and U2646 (N_2646,N_1986,N_2361);
xnor U2647 (N_2647,N_2144,N_2261);
nand U2648 (N_2648,N_2410,N_2066);
nand U2649 (N_2649,N_1989,N_2042);
or U2650 (N_2650,N_2464,N_1896);
nor U2651 (N_2651,N_2143,N_1937);
and U2652 (N_2652,N_1936,N_1927);
nand U2653 (N_2653,N_1945,N_2036);
and U2654 (N_2654,N_2429,N_2317);
or U2655 (N_2655,N_2265,N_2315);
nor U2656 (N_2656,N_1883,N_2396);
and U2657 (N_2657,N_2343,N_1886);
or U2658 (N_2658,N_2296,N_2140);
nor U2659 (N_2659,N_2395,N_2231);
or U2660 (N_2660,N_2094,N_2119);
or U2661 (N_2661,N_1916,N_1920);
or U2662 (N_2662,N_1975,N_2151);
xnor U2663 (N_2663,N_2327,N_2337);
or U2664 (N_2664,N_2096,N_1878);
and U2665 (N_2665,N_2288,N_1956);
nor U2666 (N_2666,N_1905,N_2226);
nand U2667 (N_2667,N_1890,N_2391);
nand U2668 (N_2668,N_2029,N_2084);
or U2669 (N_2669,N_2179,N_2194);
or U2670 (N_2670,N_2053,N_2499);
nand U2671 (N_2671,N_2068,N_2263);
xnor U2672 (N_2672,N_2373,N_2457);
nand U2673 (N_2673,N_2128,N_2177);
nand U2674 (N_2674,N_1967,N_2108);
or U2675 (N_2675,N_2033,N_2371);
and U2676 (N_2676,N_2259,N_2320);
nand U2677 (N_2677,N_2132,N_2375);
and U2678 (N_2678,N_2267,N_2012);
or U2679 (N_2679,N_2136,N_2142);
or U2680 (N_2680,N_2023,N_2080);
or U2681 (N_2681,N_1982,N_2106);
and U2682 (N_2682,N_2161,N_2057);
or U2683 (N_2683,N_2364,N_2045);
and U2684 (N_2684,N_2469,N_2498);
or U2685 (N_2685,N_2462,N_2248);
nor U2686 (N_2686,N_1946,N_1931);
xor U2687 (N_2687,N_1985,N_1957);
xnor U2688 (N_2688,N_2087,N_2174);
nand U2689 (N_2689,N_2486,N_2065);
nand U2690 (N_2690,N_2149,N_2040);
xnor U2691 (N_2691,N_1897,N_1994);
or U2692 (N_2692,N_2322,N_1919);
nand U2693 (N_2693,N_1923,N_2291);
and U2694 (N_2694,N_2445,N_2011);
nand U2695 (N_2695,N_2474,N_2127);
or U2696 (N_2696,N_2416,N_2154);
nor U2697 (N_2697,N_1929,N_2063);
nor U2698 (N_2698,N_2146,N_2431);
or U2699 (N_2699,N_2110,N_2318);
nor U2700 (N_2700,N_1922,N_2397);
nand U2701 (N_2701,N_2448,N_2222);
xor U2702 (N_2702,N_2003,N_2028);
or U2703 (N_2703,N_2319,N_2210);
and U2704 (N_2704,N_2286,N_2293);
xor U2705 (N_2705,N_2335,N_1942);
or U2706 (N_2706,N_2447,N_2372);
and U2707 (N_2707,N_2272,N_2197);
nor U2708 (N_2708,N_2348,N_2412);
xnor U2709 (N_2709,N_2218,N_2419);
and U2710 (N_2710,N_2359,N_2439);
nor U2711 (N_2711,N_1934,N_2237);
and U2712 (N_2712,N_2035,N_1969);
xnor U2713 (N_2713,N_2323,N_2299);
nand U2714 (N_2714,N_2215,N_2004);
nand U2715 (N_2715,N_2424,N_2090);
nand U2716 (N_2716,N_2000,N_1974);
and U2717 (N_2717,N_2346,N_2098);
or U2718 (N_2718,N_1941,N_2334);
and U2719 (N_2719,N_1999,N_2032);
nor U2720 (N_2720,N_1949,N_2116);
and U2721 (N_2721,N_2402,N_2182);
or U2722 (N_2722,N_2277,N_2483);
nand U2723 (N_2723,N_2200,N_2490);
nand U2724 (N_2724,N_2321,N_2017);
and U2725 (N_2725,N_2333,N_2155);
and U2726 (N_2726,N_2187,N_1992);
and U2727 (N_2727,N_2376,N_2184);
or U2728 (N_2728,N_2484,N_2006);
nor U2729 (N_2729,N_1906,N_2362);
or U2730 (N_2730,N_1914,N_2219);
and U2731 (N_2731,N_1964,N_2225);
and U2732 (N_2732,N_2339,N_2056);
nor U2733 (N_2733,N_2400,N_2105);
or U2734 (N_2734,N_2356,N_2332);
and U2735 (N_2735,N_2156,N_2206);
nand U2736 (N_2736,N_2338,N_2168);
xnor U2737 (N_2737,N_2118,N_2238);
nor U2738 (N_2738,N_1979,N_2406);
or U2739 (N_2739,N_2316,N_2103);
nor U2740 (N_2740,N_1876,N_2390);
nor U2741 (N_2741,N_1978,N_1913);
nor U2742 (N_2742,N_2046,N_2073);
nor U2743 (N_2743,N_2007,N_2034);
and U2744 (N_2744,N_2060,N_1882);
and U2745 (N_2745,N_1981,N_1948);
or U2746 (N_2746,N_2167,N_2443);
nand U2747 (N_2747,N_2229,N_2470);
or U2748 (N_2748,N_2213,N_2354);
nand U2749 (N_2749,N_1935,N_2411);
xnor U2750 (N_2750,N_2082,N_2283);
nand U2751 (N_2751,N_2192,N_2405);
and U2752 (N_2752,N_1998,N_2401);
nand U2753 (N_2753,N_1980,N_2385);
nand U2754 (N_2754,N_1904,N_2437);
or U2755 (N_2755,N_2166,N_2220);
nor U2756 (N_2756,N_2124,N_2100);
nor U2757 (N_2757,N_1966,N_2314);
or U2758 (N_2758,N_2440,N_1962);
or U2759 (N_2759,N_2077,N_2383);
and U2760 (N_2760,N_2074,N_2380);
xor U2761 (N_2761,N_1930,N_1891);
nor U2762 (N_2762,N_2399,N_2433);
and U2763 (N_2763,N_2450,N_1893);
nand U2764 (N_2764,N_2175,N_2254);
xor U2765 (N_2765,N_1988,N_2281);
xnor U2766 (N_2766,N_2369,N_1971);
and U2767 (N_2767,N_2211,N_2442);
xnor U2768 (N_2768,N_2122,N_2239);
xnor U2769 (N_2769,N_2224,N_2290);
nand U2770 (N_2770,N_2456,N_2134);
and U2771 (N_2771,N_2153,N_2088);
xnor U2772 (N_2772,N_2190,N_1912);
and U2773 (N_2773,N_2430,N_2344);
nor U2774 (N_2774,N_2466,N_2236);
nor U2775 (N_2775,N_2471,N_2473);
or U2776 (N_2776,N_2170,N_2305);
or U2777 (N_2777,N_2240,N_1881);
or U2778 (N_2778,N_1895,N_2349);
and U2779 (N_2779,N_2091,N_1924);
or U2780 (N_2780,N_2306,N_2278);
xor U2781 (N_2781,N_2408,N_2234);
nor U2782 (N_2782,N_2420,N_2123);
nor U2783 (N_2783,N_2485,N_2350);
nor U2784 (N_2784,N_2180,N_1972);
nor U2785 (N_2785,N_2494,N_1954);
nand U2786 (N_2786,N_1960,N_2377);
xor U2787 (N_2787,N_2005,N_2078);
or U2788 (N_2788,N_2016,N_2244);
nor U2789 (N_2789,N_2160,N_2101);
nand U2790 (N_2790,N_2188,N_2148);
xnor U2791 (N_2791,N_2295,N_2081);
nor U2792 (N_2792,N_2378,N_2135);
nand U2793 (N_2793,N_2379,N_2120);
nand U2794 (N_2794,N_2415,N_2460);
nor U2795 (N_2795,N_2251,N_2162);
or U2796 (N_2796,N_1918,N_2233);
nor U2797 (N_2797,N_2014,N_2307);
xnor U2798 (N_2798,N_2199,N_2027);
nand U2799 (N_2799,N_2049,N_2285);
and U2800 (N_2800,N_1959,N_1909);
and U2801 (N_2801,N_2413,N_2093);
and U2802 (N_2802,N_2193,N_2481);
nor U2803 (N_2803,N_1987,N_2282);
and U2804 (N_2804,N_2468,N_2270);
xor U2805 (N_2805,N_2477,N_1925);
nor U2806 (N_2806,N_2092,N_1961);
and U2807 (N_2807,N_2414,N_2235);
and U2808 (N_2808,N_2010,N_2051);
and U2809 (N_2809,N_2325,N_2114);
nand U2810 (N_2810,N_2230,N_2303);
nand U2811 (N_2811,N_1887,N_2427);
nand U2812 (N_2812,N_2294,N_2234);
and U2813 (N_2813,N_1988,N_2255);
xnor U2814 (N_2814,N_2427,N_2404);
or U2815 (N_2815,N_2044,N_2426);
nand U2816 (N_2816,N_2232,N_2142);
or U2817 (N_2817,N_2394,N_2354);
xor U2818 (N_2818,N_2421,N_2251);
and U2819 (N_2819,N_2189,N_2012);
nor U2820 (N_2820,N_2024,N_2264);
xnor U2821 (N_2821,N_1910,N_2294);
nor U2822 (N_2822,N_2365,N_2175);
nand U2823 (N_2823,N_1892,N_1967);
xnor U2824 (N_2824,N_2060,N_2033);
and U2825 (N_2825,N_1897,N_1901);
nor U2826 (N_2826,N_2029,N_2282);
nor U2827 (N_2827,N_1964,N_1901);
and U2828 (N_2828,N_2394,N_2355);
xnor U2829 (N_2829,N_2298,N_2065);
and U2830 (N_2830,N_2001,N_1877);
and U2831 (N_2831,N_1895,N_1976);
nand U2832 (N_2832,N_1992,N_2118);
nand U2833 (N_2833,N_2319,N_2396);
nor U2834 (N_2834,N_2426,N_2374);
or U2835 (N_2835,N_2409,N_2303);
nor U2836 (N_2836,N_2469,N_2203);
nor U2837 (N_2837,N_2081,N_2363);
or U2838 (N_2838,N_2434,N_2230);
xnor U2839 (N_2839,N_2405,N_2386);
or U2840 (N_2840,N_2110,N_2126);
or U2841 (N_2841,N_2319,N_1876);
nand U2842 (N_2842,N_2077,N_2168);
nand U2843 (N_2843,N_1994,N_2035);
xor U2844 (N_2844,N_2049,N_2234);
xor U2845 (N_2845,N_2373,N_2088);
nand U2846 (N_2846,N_2139,N_2030);
and U2847 (N_2847,N_2108,N_2089);
nand U2848 (N_2848,N_2025,N_2104);
nand U2849 (N_2849,N_2487,N_2397);
and U2850 (N_2850,N_2148,N_2292);
nand U2851 (N_2851,N_2030,N_2357);
xor U2852 (N_2852,N_2068,N_2075);
xnor U2853 (N_2853,N_1910,N_2383);
xor U2854 (N_2854,N_2104,N_1968);
xnor U2855 (N_2855,N_1954,N_2005);
nor U2856 (N_2856,N_2266,N_1928);
nor U2857 (N_2857,N_2169,N_2105);
nand U2858 (N_2858,N_2386,N_2219);
nand U2859 (N_2859,N_2204,N_2408);
nand U2860 (N_2860,N_2476,N_2407);
nand U2861 (N_2861,N_2090,N_2402);
and U2862 (N_2862,N_2443,N_2278);
nor U2863 (N_2863,N_1910,N_2492);
nor U2864 (N_2864,N_2408,N_1995);
nand U2865 (N_2865,N_2455,N_2406);
or U2866 (N_2866,N_1910,N_2262);
and U2867 (N_2867,N_1884,N_2240);
nor U2868 (N_2868,N_2482,N_1990);
and U2869 (N_2869,N_2070,N_2290);
nand U2870 (N_2870,N_2072,N_1966);
and U2871 (N_2871,N_2187,N_2412);
and U2872 (N_2872,N_1921,N_2271);
and U2873 (N_2873,N_2287,N_2296);
and U2874 (N_2874,N_2316,N_2147);
or U2875 (N_2875,N_2368,N_2122);
nand U2876 (N_2876,N_2045,N_2151);
or U2877 (N_2877,N_2084,N_1980);
or U2878 (N_2878,N_2256,N_2369);
nand U2879 (N_2879,N_2417,N_2027);
nor U2880 (N_2880,N_1937,N_1992);
or U2881 (N_2881,N_2230,N_2076);
nand U2882 (N_2882,N_2351,N_2212);
and U2883 (N_2883,N_2391,N_2145);
xor U2884 (N_2884,N_1992,N_2054);
or U2885 (N_2885,N_2391,N_2497);
xor U2886 (N_2886,N_2461,N_1909);
xnor U2887 (N_2887,N_2049,N_2444);
nand U2888 (N_2888,N_2327,N_2490);
or U2889 (N_2889,N_2118,N_2453);
nand U2890 (N_2890,N_2160,N_2213);
xnor U2891 (N_2891,N_2350,N_2035);
nand U2892 (N_2892,N_2214,N_2463);
nand U2893 (N_2893,N_2069,N_2243);
and U2894 (N_2894,N_2034,N_2310);
nand U2895 (N_2895,N_2334,N_2232);
or U2896 (N_2896,N_2222,N_2321);
or U2897 (N_2897,N_2072,N_2055);
nor U2898 (N_2898,N_1972,N_2312);
nand U2899 (N_2899,N_2304,N_2050);
nand U2900 (N_2900,N_2454,N_2103);
xor U2901 (N_2901,N_2026,N_2397);
nand U2902 (N_2902,N_2470,N_2158);
or U2903 (N_2903,N_1990,N_1978);
nor U2904 (N_2904,N_2217,N_2490);
and U2905 (N_2905,N_2134,N_2114);
xor U2906 (N_2906,N_2055,N_2422);
nand U2907 (N_2907,N_2225,N_2403);
and U2908 (N_2908,N_2074,N_2179);
nand U2909 (N_2909,N_2330,N_2382);
or U2910 (N_2910,N_1923,N_2087);
nor U2911 (N_2911,N_1894,N_2368);
or U2912 (N_2912,N_1924,N_1945);
or U2913 (N_2913,N_2012,N_1895);
and U2914 (N_2914,N_2301,N_2049);
xnor U2915 (N_2915,N_2357,N_1879);
and U2916 (N_2916,N_1881,N_2313);
nor U2917 (N_2917,N_2115,N_2166);
xnor U2918 (N_2918,N_1901,N_2374);
nor U2919 (N_2919,N_2098,N_2092);
nor U2920 (N_2920,N_2053,N_2143);
nand U2921 (N_2921,N_2132,N_2018);
or U2922 (N_2922,N_2219,N_2063);
or U2923 (N_2923,N_2278,N_2393);
nor U2924 (N_2924,N_1987,N_2061);
or U2925 (N_2925,N_2120,N_2101);
and U2926 (N_2926,N_2249,N_2324);
nor U2927 (N_2927,N_2427,N_2400);
and U2928 (N_2928,N_2403,N_2002);
or U2929 (N_2929,N_2013,N_1978);
or U2930 (N_2930,N_2309,N_2420);
nor U2931 (N_2931,N_1960,N_1959);
nor U2932 (N_2932,N_2108,N_2110);
nand U2933 (N_2933,N_2297,N_2350);
xnor U2934 (N_2934,N_2046,N_2417);
nor U2935 (N_2935,N_2124,N_1887);
nand U2936 (N_2936,N_2351,N_2338);
or U2937 (N_2937,N_2224,N_2078);
or U2938 (N_2938,N_2448,N_2387);
xor U2939 (N_2939,N_1946,N_2454);
and U2940 (N_2940,N_2446,N_2392);
and U2941 (N_2941,N_2098,N_2216);
or U2942 (N_2942,N_2404,N_2289);
nand U2943 (N_2943,N_2193,N_1916);
or U2944 (N_2944,N_2497,N_1979);
nand U2945 (N_2945,N_2214,N_2183);
nor U2946 (N_2946,N_2214,N_2116);
nor U2947 (N_2947,N_2381,N_2433);
xnor U2948 (N_2948,N_2271,N_2097);
or U2949 (N_2949,N_2271,N_2306);
xor U2950 (N_2950,N_2001,N_2470);
nor U2951 (N_2951,N_2248,N_2456);
nor U2952 (N_2952,N_2058,N_2333);
xor U2953 (N_2953,N_2364,N_2496);
nor U2954 (N_2954,N_1969,N_2064);
xnor U2955 (N_2955,N_1902,N_2313);
nand U2956 (N_2956,N_2013,N_1887);
xor U2957 (N_2957,N_2378,N_2286);
and U2958 (N_2958,N_2011,N_2194);
nand U2959 (N_2959,N_2484,N_2410);
nor U2960 (N_2960,N_2427,N_1959);
and U2961 (N_2961,N_2463,N_2379);
xor U2962 (N_2962,N_2438,N_1990);
or U2963 (N_2963,N_1997,N_1960);
and U2964 (N_2964,N_1932,N_2103);
nor U2965 (N_2965,N_2132,N_1881);
nor U2966 (N_2966,N_1992,N_1907);
xor U2967 (N_2967,N_2320,N_2234);
and U2968 (N_2968,N_2397,N_2226);
and U2969 (N_2969,N_2050,N_2482);
nand U2970 (N_2970,N_1912,N_2496);
nor U2971 (N_2971,N_1900,N_2158);
and U2972 (N_2972,N_2147,N_1946);
nand U2973 (N_2973,N_2170,N_2155);
or U2974 (N_2974,N_2189,N_2188);
nor U2975 (N_2975,N_2109,N_2482);
xnor U2976 (N_2976,N_2058,N_1878);
or U2977 (N_2977,N_2356,N_2158);
xnor U2978 (N_2978,N_2159,N_2334);
nand U2979 (N_2979,N_1958,N_2474);
nor U2980 (N_2980,N_2288,N_2284);
xor U2981 (N_2981,N_2114,N_2355);
xor U2982 (N_2982,N_2499,N_2294);
xnor U2983 (N_2983,N_1886,N_2179);
or U2984 (N_2984,N_2056,N_2178);
and U2985 (N_2985,N_1915,N_2462);
nand U2986 (N_2986,N_2037,N_1964);
nor U2987 (N_2987,N_2148,N_2315);
and U2988 (N_2988,N_2376,N_2386);
nand U2989 (N_2989,N_2186,N_1998);
xnor U2990 (N_2990,N_1948,N_2454);
nand U2991 (N_2991,N_2443,N_2348);
nand U2992 (N_2992,N_2314,N_2020);
and U2993 (N_2993,N_2443,N_1950);
or U2994 (N_2994,N_2055,N_2310);
nand U2995 (N_2995,N_2134,N_1978);
xnor U2996 (N_2996,N_1973,N_2151);
nand U2997 (N_2997,N_2307,N_2103);
nor U2998 (N_2998,N_1971,N_2240);
nor U2999 (N_2999,N_1929,N_1884);
nor U3000 (N_3000,N_2490,N_1919);
or U3001 (N_3001,N_2449,N_2292);
xnor U3002 (N_3002,N_2298,N_1882);
nor U3003 (N_3003,N_2221,N_2006);
nor U3004 (N_3004,N_2026,N_2375);
nor U3005 (N_3005,N_2306,N_2107);
and U3006 (N_3006,N_2275,N_2119);
nor U3007 (N_3007,N_2046,N_2062);
nor U3008 (N_3008,N_2440,N_2067);
and U3009 (N_3009,N_2004,N_2050);
xnor U3010 (N_3010,N_2060,N_1886);
nor U3011 (N_3011,N_2120,N_2013);
xnor U3012 (N_3012,N_2100,N_2333);
nor U3013 (N_3013,N_2299,N_2343);
xnor U3014 (N_3014,N_2217,N_2338);
nor U3015 (N_3015,N_2353,N_2195);
and U3016 (N_3016,N_2272,N_1879);
nand U3017 (N_3017,N_1900,N_2032);
xor U3018 (N_3018,N_1991,N_2091);
and U3019 (N_3019,N_2051,N_2368);
nand U3020 (N_3020,N_1875,N_2108);
nor U3021 (N_3021,N_2145,N_2256);
nor U3022 (N_3022,N_2331,N_2492);
and U3023 (N_3023,N_2477,N_2376);
xnor U3024 (N_3024,N_1970,N_2071);
nor U3025 (N_3025,N_2253,N_2215);
nor U3026 (N_3026,N_2068,N_2371);
and U3027 (N_3027,N_2321,N_2036);
and U3028 (N_3028,N_2318,N_2019);
nor U3029 (N_3029,N_2386,N_2004);
nor U3030 (N_3030,N_2061,N_2125);
and U3031 (N_3031,N_1994,N_2122);
nor U3032 (N_3032,N_2126,N_2251);
and U3033 (N_3033,N_2020,N_2019);
or U3034 (N_3034,N_2419,N_2152);
xor U3035 (N_3035,N_2153,N_2405);
and U3036 (N_3036,N_1878,N_1991);
or U3037 (N_3037,N_1901,N_2411);
or U3038 (N_3038,N_2178,N_2097);
nand U3039 (N_3039,N_2231,N_1934);
nand U3040 (N_3040,N_1900,N_2200);
or U3041 (N_3041,N_2001,N_2277);
or U3042 (N_3042,N_2411,N_2148);
nor U3043 (N_3043,N_1910,N_2108);
nor U3044 (N_3044,N_2485,N_2023);
nand U3045 (N_3045,N_2385,N_2439);
and U3046 (N_3046,N_2162,N_2284);
xnor U3047 (N_3047,N_1995,N_2013);
nand U3048 (N_3048,N_2369,N_2276);
and U3049 (N_3049,N_2062,N_2335);
nand U3050 (N_3050,N_1979,N_2183);
nand U3051 (N_3051,N_2212,N_2357);
xor U3052 (N_3052,N_1994,N_2445);
nand U3053 (N_3053,N_2359,N_2405);
and U3054 (N_3054,N_2189,N_1980);
nand U3055 (N_3055,N_2356,N_2322);
xnor U3056 (N_3056,N_1946,N_2400);
nor U3057 (N_3057,N_1926,N_2156);
xor U3058 (N_3058,N_2339,N_2069);
nor U3059 (N_3059,N_2048,N_2278);
xnor U3060 (N_3060,N_2234,N_1922);
nor U3061 (N_3061,N_2468,N_2144);
nor U3062 (N_3062,N_2423,N_1994);
and U3063 (N_3063,N_2242,N_2239);
xor U3064 (N_3064,N_2039,N_1994);
or U3065 (N_3065,N_2455,N_1981);
nand U3066 (N_3066,N_2348,N_2312);
and U3067 (N_3067,N_2202,N_2134);
xor U3068 (N_3068,N_2204,N_2008);
nand U3069 (N_3069,N_1972,N_1978);
xnor U3070 (N_3070,N_2173,N_2382);
and U3071 (N_3071,N_2218,N_2350);
or U3072 (N_3072,N_2453,N_1984);
nand U3073 (N_3073,N_2048,N_1905);
nor U3074 (N_3074,N_2207,N_2305);
nand U3075 (N_3075,N_1918,N_2013);
and U3076 (N_3076,N_2375,N_2152);
xor U3077 (N_3077,N_2073,N_2290);
or U3078 (N_3078,N_2083,N_2356);
nand U3079 (N_3079,N_2122,N_1970);
xnor U3080 (N_3080,N_2253,N_2401);
nor U3081 (N_3081,N_2311,N_2122);
or U3082 (N_3082,N_2327,N_2471);
and U3083 (N_3083,N_1940,N_2072);
xnor U3084 (N_3084,N_1953,N_2160);
or U3085 (N_3085,N_1998,N_1923);
nand U3086 (N_3086,N_2248,N_2366);
or U3087 (N_3087,N_1963,N_2105);
nand U3088 (N_3088,N_2107,N_2118);
nand U3089 (N_3089,N_2343,N_1915);
or U3090 (N_3090,N_2386,N_1875);
nor U3091 (N_3091,N_2476,N_1971);
and U3092 (N_3092,N_2126,N_2033);
nand U3093 (N_3093,N_2468,N_2066);
or U3094 (N_3094,N_1962,N_2434);
xnor U3095 (N_3095,N_1880,N_1895);
and U3096 (N_3096,N_2040,N_2164);
xnor U3097 (N_3097,N_2221,N_2496);
nand U3098 (N_3098,N_2081,N_2033);
xnor U3099 (N_3099,N_2155,N_2417);
nand U3100 (N_3100,N_2203,N_2277);
nor U3101 (N_3101,N_1895,N_2113);
nand U3102 (N_3102,N_2496,N_2497);
or U3103 (N_3103,N_2124,N_2287);
nand U3104 (N_3104,N_1987,N_2432);
nor U3105 (N_3105,N_1890,N_2218);
nand U3106 (N_3106,N_1981,N_2218);
nor U3107 (N_3107,N_1978,N_2233);
nand U3108 (N_3108,N_2492,N_2032);
and U3109 (N_3109,N_2094,N_2067);
or U3110 (N_3110,N_2417,N_2115);
nor U3111 (N_3111,N_2189,N_1982);
nand U3112 (N_3112,N_2360,N_1945);
nor U3113 (N_3113,N_1974,N_2014);
nor U3114 (N_3114,N_2041,N_2404);
and U3115 (N_3115,N_2175,N_2417);
and U3116 (N_3116,N_1890,N_2462);
and U3117 (N_3117,N_2328,N_2077);
or U3118 (N_3118,N_1876,N_2245);
xor U3119 (N_3119,N_2135,N_2036);
nor U3120 (N_3120,N_2029,N_1931);
nand U3121 (N_3121,N_2115,N_2121);
xnor U3122 (N_3122,N_1961,N_2329);
xor U3123 (N_3123,N_2007,N_1989);
xnor U3124 (N_3124,N_2019,N_2029);
and U3125 (N_3125,N_3110,N_2678);
nor U3126 (N_3126,N_2600,N_2525);
nand U3127 (N_3127,N_2539,N_3076);
and U3128 (N_3128,N_2542,N_2711);
nor U3129 (N_3129,N_2992,N_2758);
nor U3130 (N_3130,N_2624,N_2683);
nor U3131 (N_3131,N_2805,N_3109);
xor U3132 (N_3132,N_2519,N_2569);
nand U3133 (N_3133,N_2800,N_3031);
nand U3134 (N_3134,N_2911,N_2703);
nor U3135 (N_3135,N_3048,N_3094);
nor U3136 (N_3136,N_3055,N_3034);
and U3137 (N_3137,N_3000,N_2796);
xnor U3138 (N_3138,N_2851,N_3095);
nor U3139 (N_3139,N_3015,N_2852);
xnor U3140 (N_3140,N_2652,N_2513);
xnor U3141 (N_3141,N_3027,N_2535);
nand U3142 (N_3142,N_3052,N_2508);
or U3143 (N_3143,N_2865,N_2933);
nor U3144 (N_3144,N_2716,N_2505);
nor U3145 (N_3145,N_2787,N_2616);
and U3146 (N_3146,N_2854,N_2580);
nor U3147 (N_3147,N_2672,N_2896);
xor U3148 (N_3148,N_2515,N_2629);
xnor U3149 (N_3149,N_2993,N_3041);
and U3150 (N_3150,N_2808,N_2862);
and U3151 (N_3151,N_2700,N_2951);
or U3152 (N_3152,N_2605,N_2615);
and U3153 (N_3153,N_2832,N_2744);
nor U3154 (N_3154,N_3099,N_2870);
nand U3155 (N_3155,N_2528,N_2633);
xor U3156 (N_3156,N_2734,N_2770);
nor U3157 (N_3157,N_2756,N_2562);
xnor U3158 (N_3158,N_2594,N_2721);
and U3159 (N_3159,N_3006,N_2708);
xnor U3160 (N_3160,N_2799,N_2861);
or U3161 (N_3161,N_2867,N_3085);
or U3162 (N_3162,N_2655,N_2897);
xnor U3163 (N_3163,N_2658,N_2641);
and U3164 (N_3164,N_2934,N_2783);
nand U3165 (N_3165,N_3014,N_2893);
xor U3166 (N_3166,N_3045,N_2737);
and U3167 (N_3167,N_2841,N_2617);
and U3168 (N_3168,N_2809,N_2524);
and U3169 (N_3169,N_2776,N_2907);
xnor U3170 (N_3170,N_2803,N_2604);
xor U3171 (N_3171,N_2802,N_2696);
nand U3172 (N_3172,N_2559,N_2793);
or U3173 (N_3173,N_2686,N_2974);
and U3174 (N_3174,N_2750,N_2961);
xnor U3175 (N_3175,N_2845,N_2684);
nor U3176 (N_3176,N_2685,N_2731);
nor U3177 (N_3177,N_2578,N_2664);
xnor U3178 (N_3178,N_2925,N_2522);
xor U3179 (N_3179,N_3082,N_2648);
nand U3180 (N_3180,N_3001,N_3043);
nor U3181 (N_3181,N_3040,N_2975);
or U3182 (N_3182,N_2697,N_3111);
xnor U3183 (N_3183,N_2614,N_2811);
xnor U3184 (N_3184,N_2673,N_2835);
or U3185 (N_3185,N_3103,N_2838);
and U3186 (N_3186,N_3080,N_2608);
nor U3187 (N_3187,N_2691,N_2848);
nor U3188 (N_3188,N_2837,N_2806);
nor U3189 (N_3189,N_2695,N_2602);
or U3190 (N_3190,N_2530,N_2613);
xor U3191 (N_3191,N_3112,N_2928);
nand U3192 (N_3192,N_2692,N_2903);
xnor U3193 (N_3193,N_2989,N_2637);
nand U3194 (N_3194,N_2693,N_2757);
nor U3195 (N_3195,N_3039,N_2581);
nor U3196 (N_3196,N_2959,N_2509);
nand U3197 (N_3197,N_2639,N_2831);
or U3198 (N_3198,N_2814,N_2858);
and U3199 (N_3199,N_2970,N_2883);
or U3200 (N_3200,N_2926,N_2937);
xor U3201 (N_3201,N_3011,N_2636);
or U3202 (N_3202,N_2909,N_2628);
or U3203 (N_3203,N_2801,N_3056);
and U3204 (N_3204,N_2726,N_2709);
xnor U3205 (N_3205,N_3046,N_2634);
nor U3206 (N_3206,N_2548,N_2815);
nor U3207 (N_3207,N_3054,N_3021);
nand U3208 (N_3208,N_2900,N_2775);
and U3209 (N_3209,N_3102,N_2753);
nor U3210 (N_3210,N_2784,N_2729);
nand U3211 (N_3211,N_2556,N_2752);
nor U3212 (N_3212,N_3049,N_3051);
xnor U3213 (N_3213,N_2665,N_2844);
nor U3214 (N_3214,N_2751,N_2719);
and U3215 (N_3215,N_2789,N_3067);
nor U3216 (N_3216,N_2606,N_2518);
nand U3217 (N_3217,N_2923,N_2612);
and U3218 (N_3218,N_2620,N_2586);
or U3219 (N_3219,N_3088,N_2743);
nand U3220 (N_3220,N_2874,N_2813);
nor U3221 (N_3221,N_3115,N_2792);
nor U3222 (N_3222,N_2982,N_3122);
nand U3223 (N_3223,N_2998,N_2681);
nor U3224 (N_3224,N_2866,N_2521);
or U3225 (N_3225,N_2710,N_2856);
xor U3226 (N_3226,N_2849,N_2557);
nand U3227 (N_3227,N_2918,N_2772);
or U3228 (N_3228,N_2999,N_2882);
nand U3229 (N_3229,N_2912,N_2980);
nor U3230 (N_3230,N_2847,N_2887);
nand U3231 (N_3231,N_2917,N_2952);
or U3232 (N_3232,N_2836,N_2820);
and U3233 (N_3233,N_2859,N_2654);
xnor U3234 (N_3234,N_2596,N_2643);
xnor U3235 (N_3235,N_2707,N_2574);
or U3236 (N_3236,N_2924,N_2759);
or U3237 (N_3237,N_2694,N_2979);
nand U3238 (N_3238,N_2771,N_2584);
and U3239 (N_3239,N_3053,N_2798);
xnor U3240 (N_3240,N_2794,N_2857);
and U3241 (N_3241,N_2864,N_3119);
xor U3242 (N_3242,N_3118,N_2516);
nand U3243 (N_3243,N_2607,N_2780);
nand U3244 (N_3244,N_2589,N_2736);
and U3245 (N_3245,N_2902,N_2778);
or U3246 (N_3246,N_2948,N_2941);
or U3247 (N_3247,N_2843,N_2646);
or U3248 (N_3248,N_2564,N_2728);
and U3249 (N_3249,N_2537,N_2938);
and U3250 (N_3250,N_3108,N_2632);
xnor U3251 (N_3251,N_2609,N_2939);
nand U3252 (N_3252,N_3037,N_3042);
xor U3253 (N_3253,N_2830,N_3057);
or U3254 (N_3254,N_2571,N_2833);
nor U3255 (N_3255,N_2791,N_2669);
and U3256 (N_3256,N_2875,N_2825);
nand U3257 (N_3257,N_2877,N_2619);
or U3258 (N_3258,N_2610,N_3065);
and U3259 (N_3259,N_2774,N_3093);
and U3260 (N_3260,N_2949,N_3038);
or U3261 (N_3261,N_2720,N_3050);
or U3262 (N_3262,N_2567,N_3008);
xnor U3263 (N_3263,N_2807,N_2839);
nand U3264 (N_3264,N_2790,N_2898);
xor U3265 (N_3265,N_3107,N_2527);
nor U3266 (N_3266,N_3114,N_2576);
and U3267 (N_3267,N_2512,N_2585);
and U3268 (N_3268,N_2546,N_2593);
and U3269 (N_3269,N_2915,N_2745);
nand U3270 (N_3270,N_2985,N_2676);
and U3271 (N_3271,N_2657,N_2741);
xnor U3272 (N_3272,N_3070,N_2573);
xnor U3273 (N_3273,N_3026,N_2510);
or U3274 (N_3274,N_2929,N_2520);
and U3275 (N_3275,N_2829,N_2552);
or U3276 (N_3276,N_2551,N_2554);
nand U3277 (N_3277,N_2812,N_2868);
and U3278 (N_3278,N_2943,N_2880);
nor U3279 (N_3279,N_2595,N_2818);
nand U3280 (N_3280,N_2717,N_2969);
xor U3281 (N_3281,N_2653,N_2671);
nand U3282 (N_3282,N_2855,N_3081);
nor U3283 (N_3283,N_3068,N_2922);
or U3284 (N_3284,N_3092,N_2765);
nand U3285 (N_3285,N_2725,N_3061);
nand U3286 (N_3286,N_3100,N_2647);
xor U3287 (N_3287,N_3084,N_3060);
or U3288 (N_3288,N_2531,N_2821);
xnor U3289 (N_3289,N_2819,N_2704);
nand U3290 (N_3290,N_3018,N_2740);
nor U3291 (N_3291,N_2591,N_2876);
nand U3292 (N_3292,N_3071,N_2699);
xnor U3293 (N_3293,N_3032,N_2529);
and U3294 (N_3294,N_3097,N_2895);
and U3295 (N_3295,N_2713,N_2885);
and U3296 (N_3296,N_2860,N_2538);
nor U3297 (N_3297,N_2566,N_3012);
or U3298 (N_3298,N_2964,N_2781);
xor U3299 (N_3299,N_2588,N_2611);
or U3300 (N_3300,N_2890,N_3098);
or U3301 (N_3301,N_2582,N_3105);
xor U3302 (N_3302,N_2755,N_2668);
nand U3303 (N_3303,N_3120,N_3007);
xnor U3304 (N_3304,N_2931,N_3101);
nand U3305 (N_3305,N_2545,N_3091);
xnor U3306 (N_3306,N_2735,N_2732);
nand U3307 (N_3307,N_2804,N_2638);
nand U3308 (N_3308,N_2879,N_3069);
or U3309 (N_3309,N_2718,N_2727);
and U3310 (N_3310,N_2599,N_3009);
xor U3311 (N_3311,N_2984,N_3005);
nor U3312 (N_3312,N_2677,N_2987);
xor U3313 (N_3313,N_2598,N_2666);
or U3314 (N_3314,N_3023,N_2826);
nor U3315 (N_3315,N_2797,N_2966);
and U3316 (N_3316,N_2635,N_2627);
nor U3317 (N_3317,N_2660,N_3121);
nand U3318 (N_3318,N_3017,N_2722);
nor U3319 (N_3319,N_2506,N_2850);
nand U3320 (N_3320,N_2945,N_2878);
xor U3321 (N_3321,N_2523,N_3064);
and U3322 (N_3322,N_2560,N_2702);
or U3323 (N_3323,N_2511,N_2988);
xor U3324 (N_3324,N_2502,N_2978);
and U3325 (N_3325,N_2714,N_2983);
xor U3326 (N_3326,N_2640,N_2682);
nand U3327 (N_3327,N_2561,N_2942);
xnor U3328 (N_3328,N_2822,N_2568);
nand U3329 (N_3329,N_3030,N_3073);
nand U3330 (N_3330,N_2763,N_2997);
nor U3331 (N_3331,N_2863,N_2563);
nand U3332 (N_3332,N_2908,N_2846);
or U3333 (N_3333,N_2921,N_2881);
or U3334 (N_3334,N_2533,N_2946);
xor U3335 (N_3335,N_2760,N_2786);
nand U3336 (N_3336,N_2958,N_2904);
nor U3337 (N_3337,N_3117,N_2587);
and U3338 (N_3338,N_2603,N_3090);
nand U3339 (N_3339,N_3078,N_3003);
or U3340 (N_3340,N_2575,N_2723);
xor U3341 (N_3341,N_2824,N_2621);
and U3342 (N_3342,N_3033,N_2944);
or U3343 (N_3343,N_2549,N_2504);
xor U3344 (N_3344,N_2910,N_2656);
xor U3345 (N_3345,N_2746,N_2782);
nand U3346 (N_3346,N_2749,N_2828);
nand U3347 (N_3347,N_2543,N_3116);
nor U3348 (N_3348,N_3020,N_2739);
and U3349 (N_3349,N_2661,N_3044);
nor U3350 (N_3350,N_3002,N_2674);
or U3351 (N_3351,N_2583,N_2873);
and U3352 (N_3352,N_2884,N_2947);
nor U3353 (N_3353,N_2555,N_2690);
or U3354 (N_3354,N_3087,N_3013);
or U3355 (N_3355,N_2761,N_2935);
nand U3356 (N_3356,N_2834,N_2767);
or U3357 (N_3357,N_2747,N_2748);
nor U3358 (N_3358,N_2577,N_2892);
nor U3359 (N_3359,N_2572,N_2842);
nand U3360 (N_3360,N_2894,N_2706);
and U3361 (N_3361,N_2905,N_2590);
nand U3362 (N_3362,N_2940,N_3025);
nor U3363 (N_3363,N_2623,N_2971);
xnor U3364 (N_3364,N_2899,N_2766);
nand U3365 (N_3365,N_2667,N_2977);
nor U3366 (N_3366,N_3059,N_2630);
nand U3367 (N_3367,N_2779,N_2965);
and U3368 (N_3368,N_2994,N_2827);
xor U3369 (N_3369,N_2517,N_2990);
xnor U3370 (N_3370,N_3123,N_3047);
and U3371 (N_3371,N_2954,N_3106);
nand U3372 (N_3372,N_2514,N_2995);
nand U3373 (N_3373,N_2795,N_3074);
nor U3374 (N_3374,N_2730,N_3024);
and U3375 (N_3375,N_2651,N_2626);
nor U3376 (N_3376,N_2622,N_2631);
nor U3377 (N_3377,N_3066,N_2769);
and U3378 (N_3378,N_2930,N_2962);
nand U3379 (N_3379,N_2953,N_2932);
and U3380 (N_3380,N_2565,N_3075);
and U3381 (N_3381,N_2742,N_3036);
nand U3382 (N_3382,N_2976,N_2705);
nor U3383 (N_3383,N_2956,N_2888);
nor U3384 (N_3384,N_2810,N_2500);
nor U3385 (N_3385,N_2936,N_3010);
nor U3386 (N_3386,N_2871,N_2916);
nand U3387 (N_3387,N_2724,N_2972);
xor U3388 (N_3388,N_3104,N_2986);
and U3389 (N_3389,N_3019,N_2579);
xor U3390 (N_3390,N_3029,N_2601);
nand U3391 (N_3391,N_2853,N_2960);
or U3392 (N_3392,N_2663,N_3058);
nand U3393 (N_3393,N_2872,N_2715);
xnor U3394 (N_3394,N_2503,N_3077);
nand U3395 (N_3395,N_2913,N_2973);
nor U3396 (N_3396,N_2688,N_2625);
xor U3397 (N_3397,N_2967,N_3016);
or U3398 (N_3398,N_3062,N_2501);
xor U3399 (N_3399,N_3063,N_2869);
nor U3400 (N_3400,N_2906,N_2679);
and U3401 (N_3401,N_2963,N_2649);
xor U3402 (N_3402,N_2957,N_2689);
nand U3403 (N_3403,N_2701,N_2886);
and U3404 (N_3404,N_2642,N_2823);
nor U3405 (N_3405,N_3035,N_2991);
xnor U3406 (N_3406,N_2680,N_2532);
xnor U3407 (N_3407,N_2950,N_2785);
or U3408 (N_3408,N_2536,N_2526);
nor U3409 (N_3409,N_2891,N_2534);
or U3410 (N_3410,N_2920,N_2670);
xor U3411 (N_3411,N_2981,N_2550);
or U3412 (N_3412,N_2816,N_2840);
and U3413 (N_3413,N_3004,N_3089);
nor U3414 (N_3414,N_3028,N_2659);
and U3415 (N_3415,N_3072,N_3079);
xnor U3416 (N_3416,N_2927,N_2955);
xnor U3417 (N_3417,N_2996,N_2889);
and U3418 (N_3418,N_2773,N_3022);
xnor U3419 (N_3419,N_2675,N_2817);
and U3420 (N_3420,N_2540,N_2738);
nor U3421 (N_3421,N_2764,N_2788);
xnor U3422 (N_3422,N_2547,N_2618);
and U3423 (N_3423,N_2762,N_2644);
and U3424 (N_3424,N_3086,N_2768);
and U3425 (N_3425,N_2733,N_2698);
nand U3426 (N_3426,N_2553,N_2687);
xnor U3427 (N_3427,N_2507,N_2754);
nand U3428 (N_3428,N_2541,N_2650);
nor U3429 (N_3429,N_2592,N_2558);
nand U3430 (N_3430,N_2712,N_2777);
nor U3431 (N_3431,N_2914,N_2544);
nand U3432 (N_3432,N_3083,N_2645);
and U3433 (N_3433,N_2968,N_3124);
xnor U3434 (N_3434,N_2901,N_2570);
and U3435 (N_3435,N_2597,N_2919);
nor U3436 (N_3436,N_3096,N_2662);
nor U3437 (N_3437,N_3113,N_3085);
nor U3438 (N_3438,N_2766,N_2840);
and U3439 (N_3439,N_2667,N_2695);
nor U3440 (N_3440,N_2780,N_2580);
or U3441 (N_3441,N_2577,N_2810);
and U3442 (N_3442,N_2711,N_2831);
and U3443 (N_3443,N_2658,N_3044);
and U3444 (N_3444,N_2879,N_2983);
nand U3445 (N_3445,N_2812,N_2937);
or U3446 (N_3446,N_2797,N_2965);
nand U3447 (N_3447,N_3116,N_2612);
xor U3448 (N_3448,N_2573,N_3092);
or U3449 (N_3449,N_2609,N_2877);
or U3450 (N_3450,N_2752,N_3074);
nor U3451 (N_3451,N_2747,N_2710);
xnor U3452 (N_3452,N_2642,N_2974);
xnor U3453 (N_3453,N_2877,N_2978);
xor U3454 (N_3454,N_2553,N_2882);
nor U3455 (N_3455,N_2943,N_3036);
and U3456 (N_3456,N_2743,N_3052);
xnor U3457 (N_3457,N_2675,N_2623);
or U3458 (N_3458,N_3000,N_2758);
nor U3459 (N_3459,N_2811,N_2534);
xnor U3460 (N_3460,N_2820,N_2989);
xor U3461 (N_3461,N_2506,N_2955);
or U3462 (N_3462,N_2680,N_2959);
or U3463 (N_3463,N_2722,N_2792);
or U3464 (N_3464,N_2838,N_2857);
nor U3465 (N_3465,N_3049,N_3024);
and U3466 (N_3466,N_2964,N_2808);
nor U3467 (N_3467,N_2919,N_2613);
and U3468 (N_3468,N_2814,N_2513);
xor U3469 (N_3469,N_2510,N_3018);
nor U3470 (N_3470,N_3034,N_2937);
nor U3471 (N_3471,N_2750,N_2807);
nor U3472 (N_3472,N_2766,N_2716);
nor U3473 (N_3473,N_2642,N_2645);
nor U3474 (N_3474,N_3022,N_2648);
and U3475 (N_3475,N_2779,N_2605);
or U3476 (N_3476,N_2761,N_2658);
and U3477 (N_3477,N_2633,N_2863);
nor U3478 (N_3478,N_2735,N_2970);
and U3479 (N_3479,N_2793,N_2680);
xor U3480 (N_3480,N_2671,N_2555);
xnor U3481 (N_3481,N_2637,N_2856);
and U3482 (N_3482,N_2590,N_3055);
and U3483 (N_3483,N_2579,N_2511);
xnor U3484 (N_3484,N_2755,N_2702);
nand U3485 (N_3485,N_3069,N_2858);
and U3486 (N_3486,N_2606,N_2967);
xnor U3487 (N_3487,N_2964,N_3013);
nor U3488 (N_3488,N_2819,N_2866);
xnor U3489 (N_3489,N_2649,N_2788);
or U3490 (N_3490,N_2799,N_2928);
nand U3491 (N_3491,N_2782,N_2656);
and U3492 (N_3492,N_2844,N_3096);
nor U3493 (N_3493,N_2679,N_2963);
and U3494 (N_3494,N_2960,N_2772);
xnor U3495 (N_3495,N_2807,N_2932);
xnor U3496 (N_3496,N_2862,N_2944);
or U3497 (N_3497,N_2616,N_3035);
xnor U3498 (N_3498,N_2965,N_2518);
or U3499 (N_3499,N_2796,N_2988);
or U3500 (N_3500,N_2777,N_2526);
nor U3501 (N_3501,N_2586,N_2685);
nand U3502 (N_3502,N_2675,N_2925);
nor U3503 (N_3503,N_2579,N_2696);
or U3504 (N_3504,N_3053,N_3091);
nor U3505 (N_3505,N_2866,N_2576);
nor U3506 (N_3506,N_2796,N_2673);
nand U3507 (N_3507,N_3119,N_2992);
nor U3508 (N_3508,N_2935,N_2734);
or U3509 (N_3509,N_2688,N_2526);
or U3510 (N_3510,N_3094,N_2578);
nor U3511 (N_3511,N_2846,N_2931);
nand U3512 (N_3512,N_3025,N_3105);
nor U3513 (N_3513,N_2954,N_2825);
or U3514 (N_3514,N_2515,N_2972);
or U3515 (N_3515,N_2566,N_2702);
or U3516 (N_3516,N_2656,N_2860);
or U3517 (N_3517,N_2552,N_3114);
nor U3518 (N_3518,N_2579,N_2668);
and U3519 (N_3519,N_2786,N_2633);
or U3520 (N_3520,N_2669,N_2898);
and U3521 (N_3521,N_2809,N_3116);
xnor U3522 (N_3522,N_2756,N_2834);
nand U3523 (N_3523,N_2806,N_2932);
or U3524 (N_3524,N_2527,N_2863);
nor U3525 (N_3525,N_2678,N_2877);
nand U3526 (N_3526,N_3043,N_3048);
or U3527 (N_3527,N_2548,N_2651);
or U3528 (N_3528,N_2851,N_3027);
xnor U3529 (N_3529,N_3105,N_2723);
nand U3530 (N_3530,N_2876,N_2889);
and U3531 (N_3531,N_3086,N_2517);
nor U3532 (N_3532,N_2704,N_2653);
nand U3533 (N_3533,N_2717,N_3102);
nand U3534 (N_3534,N_2516,N_2683);
nor U3535 (N_3535,N_2910,N_2633);
nor U3536 (N_3536,N_2738,N_2704);
xor U3537 (N_3537,N_2638,N_2692);
or U3538 (N_3538,N_2606,N_3011);
or U3539 (N_3539,N_2895,N_3010);
nor U3540 (N_3540,N_2682,N_2646);
xor U3541 (N_3541,N_2857,N_2534);
and U3542 (N_3542,N_2927,N_3053);
xnor U3543 (N_3543,N_2586,N_2584);
nor U3544 (N_3544,N_2968,N_2859);
xor U3545 (N_3545,N_2559,N_3069);
or U3546 (N_3546,N_2882,N_2976);
or U3547 (N_3547,N_3082,N_3086);
nor U3548 (N_3548,N_2626,N_3010);
nor U3549 (N_3549,N_3082,N_2756);
or U3550 (N_3550,N_2847,N_2979);
and U3551 (N_3551,N_3030,N_2538);
xnor U3552 (N_3552,N_3092,N_2998);
or U3553 (N_3553,N_2969,N_3050);
xor U3554 (N_3554,N_2876,N_2648);
and U3555 (N_3555,N_2513,N_2970);
and U3556 (N_3556,N_2527,N_2603);
nor U3557 (N_3557,N_2617,N_2994);
and U3558 (N_3558,N_2698,N_2762);
and U3559 (N_3559,N_2738,N_2688);
and U3560 (N_3560,N_2908,N_2501);
xor U3561 (N_3561,N_3024,N_2500);
nor U3562 (N_3562,N_3096,N_2658);
nand U3563 (N_3563,N_2525,N_3100);
nor U3564 (N_3564,N_2794,N_2559);
xor U3565 (N_3565,N_3097,N_2754);
nand U3566 (N_3566,N_2855,N_2934);
and U3567 (N_3567,N_2940,N_2975);
or U3568 (N_3568,N_3015,N_2927);
nor U3569 (N_3569,N_3080,N_2969);
xnor U3570 (N_3570,N_2707,N_2651);
nand U3571 (N_3571,N_3052,N_2964);
or U3572 (N_3572,N_2911,N_2721);
xnor U3573 (N_3573,N_2605,N_2693);
nor U3574 (N_3574,N_2770,N_2974);
xor U3575 (N_3575,N_2853,N_2873);
nor U3576 (N_3576,N_2634,N_2864);
nor U3577 (N_3577,N_2607,N_2913);
and U3578 (N_3578,N_2880,N_3030);
nand U3579 (N_3579,N_2636,N_3015);
xnor U3580 (N_3580,N_2903,N_2680);
or U3581 (N_3581,N_3096,N_2846);
xnor U3582 (N_3582,N_2967,N_2900);
or U3583 (N_3583,N_2538,N_3020);
xor U3584 (N_3584,N_2882,N_2517);
and U3585 (N_3585,N_2736,N_3049);
nand U3586 (N_3586,N_2861,N_2875);
and U3587 (N_3587,N_2984,N_2662);
and U3588 (N_3588,N_2696,N_2520);
nand U3589 (N_3589,N_3044,N_2851);
and U3590 (N_3590,N_3048,N_2636);
and U3591 (N_3591,N_2534,N_2522);
xor U3592 (N_3592,N_2886,N_2910);
and U3593 (N_3593,N_2721,N_2704);
xor U3594 (N_3594,N_2963,N_2610);
xnor U3595 (N_3595,N_2508,N_2976);
nand U3596 (N_3596,N_2799,N_2788);
xor U3597 (N_3597,N_3107,N_2712);
and U3598 (N_3598,N_2867,N_2552);
nand U3599 (N_3599,N_2598,N_2928);
or U3600 (N_3600,N_2632,N_2544);
and U3601 (N_3601,N_2601,N_3104);
nand U3602 (N_3602,N_3072,N_2742);
nor U3603 (N_3603,N_2649,N_2905);
nand U3604 (N_3604,N_2970,N_2808);
and U3605 (N_3605,N_2931,N_2534);
nand U3606 (N_3606,N_2615,N_2810);
nor U3607 (N_3607,N_2705,N_2882);
xor U3608 (N_3608,N_2642,N_3000);
nor U3609 (N_3609,N_2574,N_2818);
xnor U3610 (N_3610,N_3082,N_2763);
or U3611 (N_3611,N_2799,N_2564);
nor U3612 (N_3612,N_2813,N_2703);
xnor U3613 (N_3613,N_2879,N_3025);
nand U3614 (N_3614,N_2640,N_2779);
xnor U3615 (N_3615,N_3024,N_2570);
xor U3616 (N_3616,N_2683,N_3074);
or U3617 (N_3617,N_2546,N_2660);
xnor U3618 (N_3618,N_2920,N_2911);
xnor U3619 (N_3619,N_2588,N_2710);
xor U3620 (N_3620,N_2624,N_2618);
nor U3621 (N_3621,N_2627,N_2735);
xnor U3622 (N_3622,N_2552,N_3088);
or U3623 (N_3623,N_2620,N_2988);
xnor U3624 (N_3624,N_2892,N_3086);
nand U3625 (N_3625,N_3002,N_2991);
xor U3626 (N_3626,N_3084,N_3002);
nor U3627 (N_3627,N_2840,N_2603);
nor U3628 (N_3628,N_2839,N_2587);
nand U3629 (N_3629,N_2745,N_2759);
nor U3630 (N_3630,N_3009,N_2911);
and U3631 (N_3631,N_2675,N_2504);
nand U3632 (N_3632,N_2784,N_2633);
or U3633 (N_3633,N_2574,N_2558);
or U3634 (N_3634,N_2758,N_2914);
xor U3635 (N_3635,N_2611,N_2772);
nand U3636 (N_3636,N_3032,N_2720);
and U3637 (N_3637,N_2731,N_2542);
nand U3638 (N_3638,N_2618,N_3104);
nor U3639 (N_3639,N_2944,N_2789);
nor U3640 (N_3640,N_2754,N_2897);
nand U3641 (N_3641,N_2574,N_2530);
nand U3642 (N_3642,N_2965,N_2685);
or U3643 (N_3643,N_2549,N_2793);
and U3644 (N_3644,N_2659,N_3008);
nor U3645 (N_3645,N_2676,N_2751);
or U3646 (N_3646,N_3087,N_2808);
or U3647 (N_3647,N_2924,N_2818);
xnor U3648 (N_3648,N_2890,N_3118);
nor U3649 (N_3649,N_2890,N_2625);
nand U3650 (N_3650,N_2649,N_2816);
or U3651 (N_3651,N_2678,N_2539);
or U3652 (N_3652,N_2610,N_3019);
and U3653 (N_3653,N_2504,N_2958);
nand U3654 (N_3654,N_2919,N_2864);
nor U3655 (N_3655,N_3104,N_2685);
xnor U3656 (N_3656,N_2975,N_2650);
nor U3657 (N_3657,N_3120,N_2841);
xor U3658 (N_3658,N_2998,N_2501);
xnor U3659 (N_3659,N_2763,N_2941);
nand U3660 (N_3660,N_2599,N_2825);
nor U3661 (N_3661,N_2731,N_2793);
and U3662 (N_3662,N_2536,N_2980);
and U3663 (N_3663,N_2571,N_2583);
nor U3664 (N_3664,N_2670,N_2850);
nand U3665 (N_3665,N_2883,N_2617);
or U3666 (N_3666,N_2992,N_3072);
xnor U3667 (N_3667,N_2877,N_2981);
nand U3668 (N_3668,N_2968,N_2571);
and U3669 (N_3669,N_2807,N_2885);
and U3670 (N_3670,N_2512,N_2829);
and U3671 (N_3671,N_2532,N_2645);
xnor U3672 (N_3672,N_2527,N_3028);
or U3673 (N_3673,N_2931,N_2720);
and U3674 (N_3674,N_2649,N_2696);
and U3675 (N_3675,N_2561,N_3047);
or U3676 (N_3676,N_2606,N_2850);
nand U3677 (N_3677,N_2568,N_3052);
nor U3678 (N_3678,N_2873,N_2766);
and U3679 (N_3679,N_3070,N_3108);
or U3680 (N_3680,N_2945,N_2573);
nand U3681 (N_3681,N_2878,N_2969);
nor U3682 (N_3682,N_2800,N_2517);
xor U3683 (N_3683,N_3073,N_3122);
nor U3684 (N_3684,N_2639,N_2847);
or U3685 (N_3685,N_2778,N_2770);
or U3686 (N_3686,N_2965,N_2922);
nand U3687 (N_3687,N_2683,N_2562);
xor U3688 (N_3688,N_2829,N_2817);
and U3689 (N_3689,N_2574,N_2886);
xor U3690 (N_3690,N_2869,N_3066);
or U3691 (N_3691,N_2836,N_2828);
or U3692 (N_3692,N_2505,N_2537);
nor U3693 (N_3693,N_3071,N_2996);
or U3694 (N_3694,N_2529,N_2843);
and U3695 (N_3695,N_2741,N_2523);
nand U3696 (N_3696,N_2661,N_2623);
nand U3697 (N_3697,N_2750,N_3012);
xnor U3698 (N_3698,N_2955,N_2940);
nand U3699 (N_3699,N_2919,N_2979);
or U3700 (N_3700,N_3091,N_2775);
and U3701 (N_3701,N_2603,N_2886);
nand U3702 (N_3702,N_2739,N_2695);
or U3703 (N_3703,N_2608,N_2574);
and U3704 (N_3704,N_2560,N_2969);
xor U3705 (N_3705,N_2543,N_2795);
xnor U3706 (N_3706,N_3026,N_3025);
nand U3707 (N_3707,N_2744,N_2994);
or U3708 (N_3708,N_3108,N_2506);
nand U3709 (N_3709,N_2566,N_2668);
nor U3710 (N_3710,N_2921,N_2592);
nor U3711 (N_3711,N_2505,N_2575);
xnor U3712 (N_3712,N_2933,N_3002);
nand U3713 (N_3713,N_2788,N_2839);
or U3714 (N_3714,N_2615,N_3018);
or U3715 (N_3715,N_3091,N_2909);
nand U3716 (N_3716,N_2773,N_2735);
xor U3717 (N_3717,N_2843,N_3094);
or U3718 (N_3718,N_2761,N_2741);
xnor U3719 (N_3719,N_3078,N_3019);
nand U3720 (N_3720,N_2930,N_2891);
or U3721 (N_3721,N_2860,N_2861);
or U3722 (N_3722,N_2581,N_3091);
or U3723 (N_3723,N_2529,N_2969);
nor U3724 (N_3724,N_2633,N_2659);
and U3725 (N_3725,N_2675,N_2894);
xnor U3726 (N_3726,N_3066,N_2587);
xnor U3727 (N_3727,N_2585,N_2502);
nor U3728 (N_3728,N_2582,N_2557);
nand U3729 (N_3729,N_2637,N_2893);
xnor U3730 (N_3730,N_3111,N_2975);
and U3731 (N_3731,N_2614,N_3073);
or U3732 (N_3732,N_3109,N_2980);
or U3733 (N_3733,N_2936,N_2574);
or U3734 (N_3734,N_2747,N_3072);
nor U3735 (N_3735,N_3006,N_2919);
or U3736 (N_3736,N_2509,N_2663);
nand U3737 (N_3737,N_2513,N_2997);
or U3738 (N_3738,N_2571,N_2577);
or U3739 (N_3739,N_2508,N_2983);
xnor U3740 (N_3740,N_3079,N_2586);
xnor U3741 (N_3741,N_2722,N_2829);
nand U3742 (N_3742,N_2650,N_2582);
xor U3743 (N_3743,N_2943,N_2583);
and U3744 (N_3744,N_2508,N_2757);
nand U3745 (N_3745,N_2780,N_3095);
and U3746 (N_3746,N_3059,N_2875);
and U3747 (N_3747,N_2894,N_2658);
and U3748 (N_3748,N_3005,N_2748);
or U3749 (N_3749,N_3113,N_3103);
and U3750 (N_3750,N_3388,N_3300);
xnor U3751 (N_3751,N_3439,N_3688);
and U3752 (N_3752,N_3650,N_3176);
xnor U3753 (N_3753,N_3391,N_3721);
or U3754 (N_3754,N_3153,N_3734);
nand U3755 (N_3755,N_3622,N_3178);
nor U3756 (N_3756,N_3307,N_3319);
or U3757 (N_3757,N_3390,N_3656);
nand U3758 (N_3758,N_3355,N_3548);
xnor U3759 (N_3759,N_3418,N_3161);
or U3760 (N_3760,N_3647,N_3185);
nand U3761 (N_3761,N_3683,N_3360);
or U3762 (N_3762,N_3210,N_3347);
or U3763 (N_3763,N_3340,N_3395);
and U3764 (N_3764,N_3484,N_3362);
xnor U3765 (N_3765,N_3242,N_3557);
or U3766 (N_3766,N_3387,N_3254);
or U3767 (N_3767,N_3130,N_3728);
xor U3768 (N_3768,N_3280,N_3173);
and U3769 (N_3769,N_3371,N_3268);
nor U3770 (N_3770,N_3188,N_3495);
and U3771 (N_3771,N_3632,N_3199);
nand U3772 (N_3772,N_3708,N_3434);
or U3773 (N_3773,N_3715,N_3139);
nor U3774 (N_3774,N_3284,N_3513);
nand U3775 (N_3775,N_3403,N_3462);
and U3776 (N_3776,N_3672,N_3614);
nand U3777 (N_3777,N_3579,N_3616);
or U3778 (N_3778,N_3287,N_3446);
nand U3779 (N_3779,N_3681,N_3179);
or U3780 (N_3780,N_3271,N_3617);
and U3781 (N_3781,N_3601,N_3432);
nor U3782 (N_3782,N_3259,N_3248);
and U3783 (N_3783,N_3564,N_3592);
and U3784 (N_3784,N_3430,N_3456);
nand U3785 (N_3785,N_3381,N_3441);
xnor U3786 (N_3786,N_3234,N_3237);
or U3787 (N_3787,N_3276,N_3565);
nor U3788 (N_3788,N_3674,N_3584);
nand U3789 (N_3789,N_3166,N_3704);
xor U3790 (N_3790,N_3748,N_3405);
or U3791 (N_3791,N_3301,N_3465);
nand U3792 (N_3792,N_3180,N_3596);
and U3793 (N_3793,N_3215,N_3163);
nand U3794 (N_3794,N_3710,N_3687);
nand U3795 (N_3795,N_3290,N_3620);
or U3796 (N_3796,N_3431,N_3494);
xor U3797 (N_3797,N_3639,N_3745);
nor U3798 (N_3798,N_3701,N_3192);
xnor U3799 (N_3799,N_3299,N_3643);
or U3800 (N_3800,N_3197,N_3401);
and U3801 (N_3801,N_3326,N_3516);
xnor U3802 (N_3802,N_3341,N_3330);
nand U3803 (N_3803,N_3133,N_3746);
or U3804 (N_3804,N_3365,N_3413);
nand U3805 (N_3805,N_3537,N_3527);
nor U3806 (N_3806,N_3295,N_3566);
nor U3807 (N_3807,N_3500,N_3306);
or U3808 (N_3808,N_3478,N_3244);
and U3809 (N_3809,N_3682,N_3706);
and U3810 (N_3810,N_3212,N_3555);
xnor U3811 (N_3811,N_3277,N_3291);
xor U3812 (N_3812,N_3172,N_3397);
and U3813 (N_3813,N_3183,N_3634);
or U3814 (N_3814,N_3556,N_3148);
or U3815 (N_3815,N_3132,N_3747);
and U3816 (N_3816,N_3597,N_3587);
nand U3817 (N_3817,N_3694,N_3547);
or U3818 (N_3818,N_3677,N_3417);
nand U3819 (N_3819,N_3470,N_3402);
or U3820 (N_3820,N_3396,N_3366);
nand U3821 (N_3821,N_3157,N_3458);
nand U3822 (N_3822,N_3506,N_3350);
xor U3823 (N_3823,N_3705,N_3385);
nand U3824 (N_3824,N_3283,N_3320);
nand U3825 (N_3825,N_3569,N_3651);
or U3826 (N_3826,N_3345,N_3539);
nor U3827 (N_3827,N_3375,N_3194);
or U3828 (N_3828,N_3658,N_3526);
or U3829 (N_3829,N_3296,N_3258);
nand U3830 (N_3830,N_3489,N_3145);
nor U3831 (N_3831,N_3571,N_3731);
or U3832 (N_3832,N_3618,N_3522);
and U3833 (N_3833,N_3243,N_3697);
nand U3834 (N_3834,N_3187,N_3600);
nand U3835 (N_3835,N_3655,N_3154);
xnor U3836 (N_3836,N_3570,N_3454);
xnor U3837 (N_3837,N_3236,N_3136);
nand U3838 (N_3838,N_3314,N_3393);
nor U3839 (N_3839,N_3333,N_3127);
and U3840 (N_3840,N_3604,N_3225);
xnor U3841 (N_3841,N_3585,N_3263);
nor U3842 (N_3842,N_3275,N_3498);
and U3843 (N_3843,N_3216,N_3593);
or U3844 (N_3844,N_3129,N_3691);
xor U3845 (N_3845,N_3572,N_3503);
or U3846 (N_3846,N_3423,N_3738);
nand U3847 (N_3847,N_3680,N_3631);
or U3848 (N_3848,N_3181,N_3313);
or U3849 (N_3849,N_3128,N_3329);
nand U3850 (N_3850,N_3214,N_3382);
or U3851 (N_3851,N_3449,N_3661);
xnor U3852 (N_3852,N_3558,N_3599);
nor U3853 (N_3853,N_3357,N_3536);
nand U3854 (N_3854,N_3359,N_3486);
nor U3855 (N_3855,N_3170,N_3147);
or U3856 (N_3856,N_3499,N_3190);
or U3857 (N_3857,N_3664,N_3560);
nor U3858 (N_3858,N_3591,N_3512);
and U3859 (N_3859,N_3137,N_3636);
xnor U3860 (N_3860,N_3709,N_3264);
and U3861 (N_3861,N_3448,N_3702);
xnor U3862 (N_3862,N_3722,N_3713);
or U3863 (N_3863,N_3553,N_3255);
xor U3864 (N_3864,N_3392,N_3220);
and U3865 (N_3865,N_3175,N_3514);
or U3866 (N_3866,N_3207,N_3652);
or U3867 (N_3867,N_3281,N_3383);
xnor U3868 (N_3868,N_3228,N_3420);
nor U3869 (N_3869,N_3668,N_3628);
xnor U3870 (N_3870,N_3676,N_3335);
xor U3871 (N_3871,N_3703,N_3156);
xor U3872 (N_3872,N_3318,N_3338);
nand U3873 (N_3873,N_3331,N_3224);
or U3874 (N_3874,N_3640,N_3419);
and U3875 (N_3875,N_3266,N_3437);
nand U3876 (N_3876,N_3546,N_3240);
and U3877 (N_3877,N_3693,N_3429);
or U3878 (N_3878,N_3576,N_3409);
and U3879 (N_3879,N_3246,N_3654);
or U3880 (N_3880,N_3377,N_3411);
xor U3881 (N_3881,N_3292,N_3563);
nand U3882 (N_3882,N_3191,N_3229);
xor U3883 (N_3883,N_3635,N_3155);
and U3884 (N_3884,N_3531,N_3743);
xnor U3885 (N_3885,N_3312,N_3151);
nand U3886 (N_3886,N_3740,N_3718);
and U3887 (N_3887,N_3325,N_3638);
nor U3888 (N_3888,N_3644,N_3646);
xor U3889 (N_3889,N_3208,N_3349);
or U3890 (N_3890,N_3669,N_3444);
xnor U3891 (N_3891,N_3552,N_3358);
nand U3892 (N_3892,N_3311,N_3406);
or U3893 (N_3893,N_3186,N_3719);
and U3894 (N_3894,N_3519,N_3233);
xnor U3895 (N_3895,N_3450,N_3256);
or U3896 (N_3896,N_3630,N_3467);
nor U3897 (N_3897,N_3222,N_3245);
and U3898 (N_3898,N_3162,N_3424);
or U3899 (N_3899,N_3700,N_3545);
or U3900 (N_3900,N_3729,N_3445);
or U3901 (N_3901,N_3665,N_3535);
nand U3902 (N_3902,N_3165,N_3414);
xnor U3903 (N_3903,N_3568,N_3485);
and U3904 (N_3904,N_3201,N_3442);
or U3905 (N_3905,N_3493,N_3158);
nor U3906 (N_3906,N_3466,N_3641);
nor U3907 (N_3907,N_3373,N_3581);
or U3908 (N_3908,N_3135,N_3407);
nand U3909 (N_3909,N_3321,N_3374);
nor U3910 (N_3910,N_3737,N_3260);
and U3911 (N_3911,N_3720,N_3297);
xor U3912 (N_3912,N_3394,N_3356);
nor U3913 (N_3913,N_3226,N_3611);
and U3914 (N_3914,N_3663,N_3613);
and U3915 (N_3915,N_3690,N_3742);
nor U3916 (N_3916,N_3131,N_3623);
or U3917 (N_3917,N_3138,N_3505);
and U3918 (N_3918,N_3447,N_3525);
xnor U3919 (N_3919,N_3274,N_3744);
and U3920 (N_3920,N_3404,N_3464);
xnor U3921 (N_3921,N_3657,N_3699);
nand U3922 (N_3922,N_3689,N_3339);
xor U3923 (N_3923,N_3438,N_3629);
nor U3924 (N_3924,N_3267,N_3412);
nor U3925 (N_3925,N_3534,N_3459);
nand U3926 (N_3926,N_3189,N_3304);
nor U3927 (N_3927,N_3473,N_3554);
nor U3928 (N_3928,N_3262,N_3421);
xnor U3929 (N_3929,N_3583,N_3574);
nand U3930 (N_3930,N_3471,N_3230);
or U3931 (N_3931,N_3559,N_3144);
xnor U3932 (N_3932,N_3344,N_3353);
nor U3933 (N_3933,N_3294,N_3384);
or U3934 (N_3934,N_3483,N_3184);
nor U3935 (N_3935,N_3491,N_3685);
nor U3936 (N_3936,N_3303,N_3348);
xor U3937 (N_3937,N_3741,N_3195);
nand U3938 (N_3938,N_3502,N_3482);
nor U3939 (N_3939,N_3218,N_3714);
nand U3940 (N_3940,N_3182,N_3528);
nand U3941 (N_3941,N_3272,N_3726);
nor U3942 (N_3942,N_3247,N_3352);
and U3943 (N_3943,N_3501,N_3322);
or U3944 (N_3944,N_3477,N_3125);
or U3945 (N_3945,N_3278,N_3435);
or U3946 (N_3946,N_3542,N_3562);
nor U3947 (N_3947,N_3608,N_3490);
nor U3948 (N_3948,N_3678,N_3143);
or U3949 (N_3949,N_3370,N_3368);
or U3950 (N_3950,N_3717,N_3152);
nor U3951 (N_3951,N_3141,N_3317);
nor U3952 (N_3952,N_3428,N_3440);
nand U3953 (N_3953,N_3507,N_3509);
nor U3954 (N_3954,N_3198,N_3455);
or U3955 (N_3955,N_3621,N_3213);
or U3956 (N_3956,N_3270,N_3219);
nand U3957 (N_3957,N_3269,N_3436);
nand U3958 (N_3958,N_3649,N_3733);
and U3959 (N_3959,N_3251,N_3305);
nand U3960 (N_3960,N_3487,N_3625);
nor U3961 (N_3961,N_3204,N_3686);
and U3962 (N_3962,N_3540,N_3206);
nor U3963 (N_3963,N_3279,N_3160);
nor U3964 (N_3964,N_3232,N_3324);
and U3965 (N_3965,N_3530,N_3711);
or U3966 (N_3966,N_3543,N_3126);
and U3967 (N_3967,N_3361,N_3725);
xnor U3968 (N_3968,N_3150,N_3732);
and U3969 (N_3969,N_3241,N_3457);
nand U3970 (N_3970,N_3205,N_3595);
xnor U3971 (N_3971,N_3451,N_3386);
nor U3972 (N_3972,N_3476,N_3351);
xnor U3973 (N_3973,N_3475,N_3425);
nand U3974 (N_3974,N_3520,N_3567);
nand U3975 (N_3975,N_3615,N_3415);
xor U3976 (N_3976,N_3480,N_3698);
or U3977 (N_3977,N_3354,N_3364);
nor U3978 (N_3978,N_3550,N_3169);
and U3979 (N_3979,N_3538,N_3452);
xor U3980 (N_3980,N_3342,N_3399);
xor U3981 (N_3981,N_3316,N_3586);
nor U3982 (N_3982,N_3217,N_3410);
or U3983 (N_3983,N_3315,N_3252);
nor U3984 (N_3984,N_3497,N_3261);
or U3985 (N_3985,N_3508,N_3168);
or U3986 (N_3986,N_3203,N_3416);
and U3987 (N_3987,N_3177,N_3749);
or U3988 (N_3988,N_3510,N_3521);
nor U3989 (N_3989,N_3285,N_3588);
xor U3990 (N_3990,N_3633,N_3167);
or U3991 (N_3991,N_3492,N_3609);
nand U3992 (N_3992,N_3221,N_3472);
xnor U3993 (N_3993,N_3610,N_3605);
nor U3994 (N_3994,N_3273,N_3727);
or U3995 (N_3995,N_3288,N_3679);
or U3996 (N_3996,N_3134,N_3529);
xnor U3997 (N_3997,N_3544,N_3735);
nor U3998 (N_3998,N_3675,N_3479);
or U3999 (N_3999,N_3164,N_3627);
xnor U4000 (N_4000,N_3524,N_3561);
and U4001 (N_4001,N_3235,N_3739);
and U4002 (N_4002,N_3606,N_3376);
or U4003 (N_4003,N_3696,N_3298);
xor U4004 (N_4004,N_3662,N_3642);
nor U4005 (N_4005,N_3323,N_3551);
and U4006 (N_4006,N_3202,N_3603);
or U4007 (N_4007,N_3174,N_3712);
nor U4008 (N_4008,N_3140,N_3575);
nand U4009 (N_4009,N_3238,N_3346);
nand U4010 (N_4010,N_3293,N_3308);
nor U4011 (N_4011,N_3626,N_3193);
or U4012 (N_4012,N_3211,N_3372);
xor U4013 (N_4013,N_3289,N_3253);
xor U4014 (N_4014,N_3343,N_3453);
nand U4015 (N_4015,N_3209,N_3648);
or U4016 (N_4016,N_3523,N_3337);
nor U4017 (N_4017,N_3334,N_3671);
nand U4018 (N_4018,N_3310,N_3624);
and U4019 (N_4019,N_3619,N_3443);
nand U4020 (N_4020,N_3496,N_3504);
and U4021 (N_4021,N_3426,N_3653);
and U4022 (N_4022,N_3573,N_3332);
nand U4023 (N_4023,N_3474,N_3670);
and U4024 (N_4024,N_3286,N_3637);
xnor U4025 (N_4025,N_3723,N_3692);
nor U4026 (N_4026,N_3363,N_3239);
nor U4027 (N_4027,N_3302,N_3380);
xor U4028 (N_4028,N_3645,N_3666);
xor U4029 (N_4029,N_3673,N_3590);
nor U4030 (N_4030,N_3367,N_3607);
or U4031 (N_4031,N_3142,N_3146);
nand U4032 (N_4032,N_3265,N_3309);
nand U4033 (N_4033,N_3196,N_3149);
and U4034 (N_4034,N_3518,N_3379);
nand U4035 (N_4035,N_3400,N_3378);
nand U4036 (N_4036,N_3577,N_3223);
nor U4037 (N_4037,N_3257,N_3336);
nor U4038 (N_4038,N_3327,N_3578);
or U4039 (N_4039,N_3589,N_3469);
and U4040 (N_4040,N_3730,N_3171);
or U4041 (N_4041,N_3408,N_3549);
nand U4042 (N_4042,N_3481,N_3541);
xor U4043 (N_4043,N_3580,N_3460);
nand U4044 (N_4044,N_3461,N_3398);
nor U4045 (N_4045,N_3612,N_3463);
xnor U4046 (N_4046,N_3427,N_3598);
xor U4047 (N_4047,N_3250,N_3369);
nand U4048 (N_4048,N_3200,N_3659);
nor U4049 (N_4049,N_3716,N_3660);
nor U4050 (N_4050,N_3515,N_3389);
xor U4051 (N_4051,N_3231,N_3227);
xnor U4052 (N_4052,N_3511,N_3422);
or U4053 (N_4053,N_3488,N_3594);
or U4054 (N_4054,N_3517,N_3724);
nor U4055 (N_4055,N_3433,N_3468);
nand U4056 (N_4056,N_3684,N_3736);
or U4057 (N_4057,N_3602,N_3707);
xnor U4058 (N_4058,N_3695,N_3667);
nor U4059 (N_4059,N_3249,N_3328);
nand U4060 (N_4060,N_3533,N_3532);
and U4061 (N_4061,N_3159,N_3282);
nor U4062 (N_4062,N_3582,N_3624);
and U4063 (N_4063,N_3364,N_3338);
and U4064 (N_4064,N_3156,N_3198);
xnor U4065 (N_4065,N_3612,N_3511);
and U4066 (N_4066,N_3432,N_3673);
or U4067 (N_4067,N_3686,N_3388);
nor U4068 (N_4068,N_3141,N_3282);
nand U4069 (N_4069,N_3715,N_3376);
xnor U4070 (N_4070,N_3500,N_3746);
xor U4071 (N_4071,N_3292,N_3307);
xnor U4072 (N_4072,N_3657,N_3175);
or U4073 (N_4073,N_3640,N_3587);
nand U4074 (N_4074,N_3158,N_3350);
and U4075 (N_4075,N_3148,N_3423);
xnor U4076 (N_4076,N_3594,N_3210);
xnor U4077 (N_4077,N_3656,N_3433);
nand U4078 (N_4078,N_3718,N_3370);
nand U4079 (N_4079,N_3201,N_3643);
or U4080 (N_4080,N_3480,N_3421);
nor U4081 (N_4081,N_3315,N_3241);
or U4082 (N_4082,N_3412,N_3328);
and U4083 (N_4083,N_3681,N_3489);
and U4084 (N_4084,N_3738,N_3484);
or U4085 (N_4085,N_3722,N_3366);
nor U4086 (N_4086,N_3347,N_3706);
xnor U4087 (N_4087,N_3734,N_3727);
and U4088 (N_4088,N_3430,N_3382);
nand U4089 (N_4089,N_3343,N_3177);
xnor U4090 (N_4090,N_3355,N_3260);
and U4091 (N_4091,N_3604,N_3542);
xnor U4092 (N_4092,N_3539,N_3226);
nand U4093 (N_4093,N_3182,N_3184);
xor U4094 (N_4094,N_3643,N_3573);
and U4095 (N_4095,N_3325,N_3183);
nand U4096 (N_4096,N_3643,N_3469);
nand U4097 (N_4097,N_3566,N_3564);
and U4098 (N_4098,N_3167,N_3557);
and U4099 (N_4099,N_3543,N_3195);
xnor U4100 (N_4100,N_3428,N_3398);
nand U4101 (N_4101,N_3613,N_3501);
nand U4102 (N_4102,N_3412,N_3612);
nor U4103 (N_4103,N_3231,N_3143);
nor U4104 (N_4104,N_3482,N_3496);
xnor U4105 (N_4105,N_3269,N_3389);
nand U4106 (N_4106,N_3309,N_3567);
and U4107 (N_4107,N_3383,N_3361);
xor U4108 (N_4108,N_3323,N_3225);
nor U4109 (N_4109,N_3142,N_3727);
nand U4110 (N_4110,N_3664,N_3359);
or U4111 (N_4111,N_3481,N_3478);
xnor U4112 (N_4112,N_3586,N_3146);
xnor U4113 (N_4113,N_3267,N_3608);
nor U4114 (N_4114,N_3704,N_3261);
nand U4115 (N_4115,N_3587,N_3345);
nor U4116 (N_4116,N_3644,N_3316);
and U4117 (N_4117,N_3217,N_3356);
xor U4118 (N_4118,N_3160,N_3525);
or U4119 (N_4119,N_3406,N_3586);
nor U4120 (N_4120,N_3521,N_3412);
nor U4121 (N_4121,N_3647,N_3687);
xor U4122 (N_4122,N_3590,N_3225);
xnor U4123 (N_4123,N_3562,N_3696);
and U4124 (N_4124,N_3656,N_3356);
xor U4125 (N_4125,N_3273,N_3445);
and U4126 (N_4126,N_3567,N_3485);
xnor U4127 (N_4127,N_3421,N_3571);
nor U4128 (N_4128,N_3575,N_3357);
xor U4129 (N_4129,N_3733,N_3325);
xnor U4130 (N_4130,N_3673,N_3287);
xnor U4131 (N_4131,N_3318,N_3733);
or U4132 (N_4132,N_3654,N_3437);
nor U4133 (N_4133,N_3162,N_3231);
nand U4134 (N_4134,N_3527,N_3457);
and U4135 (N_4135,N_3425,N_3163);
or U4136 (N_4136,N_3571,N_3226);
nand U4137 (N_4137,N_3489,N_3418);
and U4138 (N_4138,N_3749,N_3522);
or U4139 (N_4139,N_3187,N_3186);
nand U4140 (N_4140,N_3273,N_3235);
xor U4141 (N_4141,N_3720,N_3278);
nor U4142 (N_4142,N_3717,N_3460);
xor U4143 (N_4143,N_3582,N_3735);
nand U4144 (N_4144,N_3529,N_3649);
nor U4145 (N_4145,N_3306,N_3273);
xor U4146 (N_4146,N_3724,N_3672);
and U4147 (N_4147,N_3475,N_3561);
nand U4148 (N_4148,N_3173,N_3412);
and U4149 (N_4149,N_3266,N_3718);
xnor U4150 (N_4150,N_3444,N_3242);
nand U4151 (N_4151,N_3611,N_3618);
nor U4152 (N_4152,N_3193,N_3327);
and U4153 (N_4153,N_3510,N_3675);
or U4154 (N_4154,N_3323,N_3287);
nand U4155 (N_4155,N_3381,N_3499);
xor U4156 (N_4156,N_3281,N_3325);
and U4157 (N_4157,N_3368,N_3676);
xor U4158 (N_4158,N_3419,N_3169);
xor U4159 (N_4159,N_3718,N_3359);
xor U4160 (N_4160,N_3598,N_3230);
xor U4161 (N_4161,N_3325,N_3639);
nand U4162 (N_4162,N_3591,N_3624);
xnor U4163 (N_4163,N_3193,N_3444);
xor U4164 (N_4164,N_3413,N_3589);
xnor U4165 (N_4165,N_3633,N_3127);
and U4166 (N_4166,N_3566,N_3200);
and U4167 (N_4167,N_3738,N_3482);
or U4168 (N_4168,N_3190,N_3337);
and U4169 (N_4169,N_3314,N_3359);
nand U4170 (N_4170,N_3550,N_3720);
nand U4171 (N_4171,N_3688,N_3661);
xor U4172 (N_4172,N_3473,N_3496);
xor U4173 (N_4173,N_3570,N_3418);
and U4174 (N_4174,N_3352,N_3239);
nand U4175 (N_4175,N_3315,N_3209);
or U4176 (N_4176,N_3496,N_3348);
and U4177 (N_4177,N_3452,N_3334);
nor U4178 (N_4178,N_3731,N_3222);
nor U4179 (N_4179,N_3685,N_3353);
nand U4180 (N_4180,N_3272,N_3640);
nand U4181 (N_4181,N_3343,N_3675);
and U4182 (N_4182,N_3154,N_3467);
or U4183 (N_4183,N_3414,N_3569);
or U4184 (N_4184,N_3286,N_3132);
nand U4185 (N_4185,N_3696,N_3553);
and U4186 (N_4186,N_3451,N_3307);
nor U4187 (N_4187,N_3147,N_3143);
xor U4188 (N_4188,N_3232,N_3734);
xnor U4189 (N_4189,N_3632,N_3200);
and U4190 (N_4190,N_3598,N_3191);
nor U4191 (N_4191,N_3196,N_3258);
xor U4192 (N_4192,N_3747,N_3464);
xor U4193 (N_4193,N_3689,N_3255);
xor U4194 (N_4194,N_3666,N_3377);
or U4195 (N_4195,N_3240,N_3620);
nand U4196 (N_4196,N_3708,N_3711);
or U4197 (N_4197,N_3262,N_3432);
nor U4198 (N_4198,N_3300,N_3584);
or U4199 (N_4199,N_3515,N_3558);
and U4200 (N_4200,N_3441,N_3523);
and U4201 (N_4201,N_3203,N_3426);
nand U4202 (N_4202,N_3198,N_3341);
or U4203 (N_4203,N_3549,N_3490);
xor U4204 (N_4204,N_3559,N_3392);
and U4205 (N_4205,N_3552,N_3402);
and U4206 (N_4206,N_3543,N_3516);
nor U4207 (N_4207,N_3201,N_3189);
nand U4208 (N_4208,N_3517,N_3487);
or U4209 (N_4209,N_3367,N_3333);
or U4210 (N_4210,N_3243,N_3493);
nor U4211 (N_4211,N_3474,N_3403);
xnor U4212 (N_4212,N_3555,N_3639);
xor U4213 (N_4213,N_3284,N_3415);
xor U4214 (N_4214,N_3168,N_3384);
nand U4215 (N_4215,N_3716,N_3306);
nand U4216 (N_4216,N_3229,N_3499);
or U4217 (N_4217,N_3161,N_3431);
or U4218 (N_4218,N_3301,N_3369);
nor U4219 (N_4219,N_3377,N_3732);
xor U4220 (N_4220,N_3219,N_3159);
xnor U4221 (N_4221,N_3480,N_3420);
nand U4222 (N_4222,N_3302,N_3374);
or U4223 (N_4223,N_3566,N_3211);
xor U4224 (N_4224,N_3504,N_3264);
xor U4225 (N_4225,N_3404,N_3268);
or U4226 (N_4226,N_3623,N_3225);
nand U4227 (N_4227,N_3188,N_3493);
or U4228 (N_4228,N_3243,N_3317);
or U4229 (N_4229,N_3577,N_3253);
nand U4230 (N_4230,N_3422,N_3334);
or U4231 (N_4231,N_3414,N_3332);
and U4232 (N_4232,N_3460,N_3520);
nor U4233 (N_4233,N_3711,N_3332);
nand U4234 (N_4234,N_3326,N_3368);
xnor U4235 (N_4235,N_3435,N_3602);
or U4236 (N_4236,N_3468,N_3175);
nor U4237 (N_4237,N_3400,N_3527);
nor U4238 (N_4238,N_3709,N_3649);
nor U4239 (N_4239,N_3693,N_3341);
xor U4240 (N_4240,N_3137,N_3531);
nor U4241 (N_4241,N_3377,N_3560);
nor U4242 (N_4242,N_3227,N_3420);
nor U4243 (N_4243,N_3531,N_3706);
xor U4244 (N_4244,N_3709,N_3667);
xor U4245 (N_4245,N_3211,N_3180);
and U4246 (N_4246,N_3315,N_3692);
nor U4247 (N_4247,N_3525,N_3616);
nand U4248 (N_4248,N_3377,N_3713);
nand U4249 (N_4249,N_3295,N_3555);
nand U4250 (N_4250,N_3270,N_3388);
or U4251 (N_4251,N_3544,N_3175);
xnor U4252 (N_4252,N_3374,N_3485);
xnor U4253 (N_4253,N_3531,N_3184);
and U4254 (N_4254,N_3735,N_3725);
nand U4255 (N_4255,N_3521,N_3577);
or U4256 (N_4256,N_3481,N_3565);
or U4257 (N_4257,N_3395,N_3501);
and U4258 (N_4258,N_3301,N_3593);
nor U4259 (N_4259,N_3445,N_3707);
or U4260 (N_4260,N_3505,N_3283);
or U4261 (N_4261,N_3373,N_3697);
xnor U4262 (N_4262,N_3492,N_3228);
xor U4263 (N_4263,N_3501,N_3130);
or U4264 (N_4264,N_3523,N_3344);
and U4265 (N_4265,N_3219,N_3643);
nand U4266 (N_4266,N_3163,N_3487);
xnor U4267 (N_4267,N_3311,N_3688);
xnor U4268 (N_4268,N_3621,N_3599);
and U4269 (N_4269,N_3583,N_3264);
nor U4270 (N_4270,N_3292,N_3627);
nor U4271 (N_4271,N_3636,N_3313);
and U4272 (N_4272,N_3555,N_3501);
nand U4273 (N_4273,N_3230,N_3499);
or U4274 (N_4274,N_3676,N_3206);
or U4275 (N_4275,N_3606,N_3347);
or U4276 (N_4276,N_3152,N_3468);
nand U4277 (N_4277,N_3749,N_3165);
xor U4278 (N_4278,N_3688,N_3644);
xor U4279 (N_4279,N_3497,N_3689);
nor U4280 (N_4280,N_3209,N_3710);
and U4281 (N_4281,N_3653,N_3643);
nor U4282 (N_4282,N_3303,N_3301);
nand U4283 (N_4283,N_3724,N_3413);
or U4284 (N_4284,N_3486,N_3496);
and U4285 (N_4285,N_3231,N_3206);
or U4286 (N_4286,N_3220,N_3398);
or U4287 (N_4287,N_3211,N_3215);
xor U4288 (N_4288,N_3548,N_3216);
nand U4289 (N_4289,N_3694,N_3313);
and U4290 (N_4290,N_3504,N_3728);
xor U4291 (N_4291,N_3245,N_3276);
or U4292 (N_4292,N_3681,N_3400);
or U4293 (N_4293,N_3732,N_3453);
nor U4294 (N_4294,N_3562,N_3587);
nand U4295 (N_4295,N_3461,N_3747);
and U4296 (N_4296,N_3377,N_3524);
xor U4297 (N_4297,N_3366,N_3696);
and U4298 (N_4298,N_3151,N_3222);
and U4299 (N_4299,N_3355,N_3591);
nor U4300 (N_4300,N_3321,N_3259);
and U4301 (N_4301,N_3630,N_3392);
xor U4302 (N_4302,N_3194,N_3516);
nor U4303 (N_4303,N_3182,N_3198);
or U4304 (N_4304,N_3724,N_3319);
and U4305 (N_4305,N_3602,N_3271);
nand U4306 (N_4306,N_3573,N_3357);
nor U4307 (N_4307,N_3210,N_3129);
nand U4308 (N_4308,N_3441,N_3346);
and U4309 (N_4309,N_3149,N_3242);
or U4310 (N_4310,N_3516,N_3709);
and U4311 (N_4311,N_3174,N_3199);
nor U4312 (N_4312,N_3489,N_3211);
or U4313 (N_4313,N_3652,N_3589);
nor U4314 (N_4314,N_3364,N_3424);
nor U4315 (N_4315,N_3419,N_3549);
nand U4316 (N_4316,N_3265,N_3749);
nand U4317 (N_4317,N_3336,N_3406);
nor U4318 (N_4318,N_3452,N_3313);
nor U4319 (N_4319,N_3423,N_3556);
xnor U4320 (N_4320,N_3279,N_3413);
xor U4321 (N_4321,N_3398,N_3748);
or U4322 (N_4322,N_3420,N_3581);
nand U4323 (N_4323,N_3407,N_3320);
or U4324 (N_4324,N_3163,N_3341);
nand U4325 (N_4325,N_3587,N_3475);
xor U4326 (N_4326,N_3476,N_3336);
nor U4327 (N_4327,N_3712,N_3350);
xor U4328 (N_4328,N_3334,N_3627);
and U4329 (N_4329,N_3222,N_3467);
or U4330 (N_4330,N_3288,N_3494);
or U4331 (N_4331,N_3229,N_3176);
or U4332 (N_4332,N_3156,N_3359);
nor U4333 (N_4333,N_3609,N_3251);
and U4334 (N_4334,N_3486,N_3710);
or U4335 (N_4335,N_3315,N_3475);
nor U4336 (N_4336,N_3210,N_3657);
nor U4337 (N_4337,N_3342,N_3659);
xor U4338 (N_4338,N_3635,N_3551);
xor U4339 (N_4339,N_3552,N_3662);
nand U4340 (N_4340,N_3504,N_3249);
nor U4341 (N_4341,N_3749,N_3464);
nor U4342 (N_4342,N_3349,N_3198);
or U4343 (N_4343,N_3746,N_3358);
xor U4344 (N_4344,N_3365,N_3440);
xnor U4345 (N_4345,N_3258,N_3688);
nand U4346 (N_4346,N_3639,N_3206);
nor U4347 (N_4347,N_3735,N_3474);
or U4348 (N_4348,N_3270,N_3510);
and U4349 (N_4349,N_3379,N_3713);
and U4350 (N_4350,N_3462,N_3417);
nand U4351 (N_4351,N_3608,N_3571);
nand U4352 (N_4352,N_3526,N_3619);
nor U4353 (N_4353,N_3253,N_3656);
or U4354 (N_4354,N_3645,N_3714);
xor U4355 (N_4355,N_3716,N_3696);
xnor U4356 (N_4356,N_3607,N_3175);
and U4357 (N_4357,N_3349,N_3592);
nand U4358 (N_4358,N_3322,N_3177);
or U4359 (N_4359,N_3730,N_3594);
nor U4360 (N_4360,N_3400,N_3391);
nand U4361 (N_4361,N_3744,N_3147);
and U4362 (N_4362,N_3584,N_3695);
xor U4363 (N_4363,N_3480,N_3273);
or U4364 (N_4364,N_3192,N_3295);
nand U4365 (N_4365,N_3266,N_3197);
xnor U4366 (N_4366,N_3535,N_3165);
or U4367 (N_4367,N_3596,N_3388);
nor U4368 (N_4368,N_3660,N_3234);
or U4369 (N_4369,N_3566,N_3382);
xnor U4370 (N_4370,N_3341,N_3645);
or U4371 (N_4371,N_3423,N_3228);
and U4372 (N_4372,N_3365,N_3152);
or U4373 (N_4373,N_3127,N_3245);
xnor U4374 (N_4374,N_3448,N_3494);
or U4375 (N_4375,N_4360,N_3823);
or U4376 (N_4376,N_4278,N_3781);
nor U4377 (N_4377,N_3861,N_3853);
nand U4378 (N_4378,N_3836,N_4192);
or U4379 (N_4379,N_4059,N_3865);
nand U4380 (N_4380,N_3899,N_4023);
xnor U4381 (N_4381,N_3972,N_4353);
and U4382 (N_4382,N_3875,N_4131);
and U4383 (N_4383,N_4259,N_4168);
or U4384 (N_4384,N_3835,N_4204);
nand U4385 (N_4385,N_4033,N_4336);
xor U4386 (N_4386,N_4157,N_4241);
or U4387 (N_4387,N_4311,N_4319);
or U4388 (N_4388,N_4374,N_4301);
or U4389 (N_4389,N_4046,N_4169);
and U4390 (N_4390,N_4048,N_4290);
and U4391 (N_4391,N_4367,N_4300);
nand U4392 (N_4392,N_4293,N_3780);
nor U4393 (N_4393,N_4020,N_4053);
and U4394 (N_4394,N_3815,N_3832);
xor U4395 (N_4395,N_3802,N_3943);
xor U4396 (N_4396,N_3866,N_4189);
nor U4397 (N_4397,N_3950,N_3918);
and U4398 (N_4398,N_4337,N_3812);
xor U4399 (N_4399,N_4183,N_3882);
xnor U4400 (N_4400,N_4151,N_4282);
or U4401 (N_4401,N_3818,N_4264);
or U4402 (N_4402,N_3798,N_3952);
or U4403 (N_4403,N_4056,N_4086);
nor U4404 (N_4404,N_3940,N_4087);
or U4405 (N_4405,N_3775,N_3880);
and U4406 (N_4406,N_4182,N_4312);
xnor U4407 (N_4407,N_3816,N_4012);
xor U4408 (N_4408,N_4158,N_4320);
nor U4409 (N_4409,N_3784,N_4295);
nand U4410 (N_4410,N_3762,N_4141);
nor U4411 (N_4411,N_3975,N_4016);
nand U4412 (N_4412,N_3929,N_4093);
nor U4413 (N_4413,N_4283,N_4231);
or U4414 (N_4414,N_3826,N_4036);
nor U4415 (N_4415,N_3951,N_4260);
xor U4416 (N_4416,N_3825,N_3855);
nand U4417 (N_4417,N_3752,N_3821);
or U4418 (N_4418,N_4124,N_4212);
xnor U4419 (N_4419,N_3787,N_4326);
and U4420 (N_4420,N_4196,N_4116);
and U4421 (N_4421,N_4040,N_4126);
or U4422 (N_4422,N_3834,N_4115);
nor U4423 (N_4423,N_3953,N_3849);
or U4424 (N_4424,N_4111,N_3892);
or U4425 (N_4425,N_3936,N_4345);
nor U4426 (N_4426,N_4245,N_4099);
nor U4427 (N_4427,N_4167,N_3898);
or U4428 (N_4428,N_4247,N_4058);
and U4429 (N_4429,N_4230,N_4346);
and U4430 (N_4430,N_4054,N_4011);
xnor U4431 (N_4431,N_4330,N_3799);
nor U4432 (N_4432,N_4163,N_3765);
xnor U4433 (N_4433,N_3938,N_3924);
nand U4434 (N_4434,N_3981,N_4074);
xor U4435 (N_4435,N_4223,N_4318);
or U4436 (N_4436,N_4370,N_4195);
nor U4437 (N_4437,N_4096,N_4242);
xnor U4438 (N_4438,N_4339,N_3988);
nor U4439 (N_4439,N_4085,N_3805);
nor U4440 (N_4440,N_3770,N_4051);
nand U4441 (N_4441,N_3997,N_4049);
nor U4442 (N_4442,N_4275,N_4200);
or U4443 (N_4443,N_3911,N_3901);
nor U4444 (N_4444,N_4171,N_4215);
and U4445 (N_4445,N_4310,N_4080);
nand U4446 (N_4446,N_4135,N_4348);
xor U4447 (N_4447,N_4137,N_4075);
and U4448 (N_4448,N_4237,N_4334);
nand U4449 (N_4449,N_4229,N_3904);
xor U4450 (N_4450,N_3846,N_4338);
xor U4451 (N_4451,N_3862,N_3960);
nand U4452 (N_4452,N_4184,N_4072);
xor U4453 (N_4453,N_4327,N_4366);
xnor U4454 (N_4454,N_3779,N_3927);
nor U4455 (N_4455,N_4209,N_3800);
nor U4456 (N_4456,N_4324,N_3791);
or U4457 (N_4457,N_4057,N_3813);
or U4458 (N_4458,N_4153,N_3778);
xnor U4459 (N_4459,N_4240,N_4173);
xor U4460 (N_4460,N_4206,N_3999);
nor U4461 (N_4461,N_4025,N_4018);
nor U4462 (N_4462,N_3771,N_3996);
and U4463 (N_4463,N_4226,N_4006);
or U4464 (N_4464,N_3839,N_4187);
nand U4465 (N_4465,N_4090,N_3900);
nor U4466 (N_4466,N_4152,N_4081);
nor U4467 (N_4467,N_4066,N_4165);
or U4468 (N_4468,N_3974,N_3989);
or U4469 (N_4469,N_4084,N_4021);
nand U4470 (N_4470,N_3970,N_3944);
nor U4471 (N_4471,N_4001,N_4091);
nand U4472 (N_4472,N_3908,N_4325);
nand U4473 (N_4473,N_3930,N_3810);
xor U4474 (N_4474,N_3777,N_3844);
nand U4475 (N_4475,N_3962,N_4107);
and U4476 (N_4476,N_4292,N_4101);
nor U4477 (N_4477,N_4331,N_4009);
and U4478 (N_4478,N_4274,N_4332);
xor U4479 (N_4479,N_4267,N_3905);
nor U4480 (N_4480,N_4164,N_4019);
nor U4481 (N_4481,N_4067,N_4306);
and U4482 (N_4482,N_4233,N_4239);
nor U4483 (N_4483,N_4217,N_4007);
nand U4484 (N_4484,N_3751,N_3947);
and U4485 (N_4485,N_3754,N_4342);
and U4486 (N_4486,N_3889,N_4052);
nand U4487 (N_4487,N_3969,N_4284);
nor U4488 (N_4488,N_4110,N_4253);
or U4489 (N_4489,N_4362,N_4299);
or U4490 (N_4490,N_4022,N_4106);
nand U4491 (N_4491,N_4202,N_4155);
xor U4492 (N_4492,N_3942,N_4039);
and U4493 (N_4493,N_3856,N_4280);
or U4494 (N_4494,N_4102,N_4122);
xor U4495 (N_4495,N_3897,N_3760);
nor U4496 (N_4496,N_4246,N_3967);
and U4497 (N_4497,N_3830,N_4361);
and U4498 (N_4498,N_4079,N_4243);
nor U4499 (N_4499,N_4294,N_3803);
or U4500 (N_4500,N_3890,N_4277);
or U4501 (N_4501,N_4117,N_3776);
nor U4502 (N_4502,N_4272,N_3923);
or U4503 (N_4503,N_3842,N_4088);
or U4504 (N_4504,N_3946,N_3966);
xor U4505 (N_4505,N_3759,N_4030);
and U4506 (N_4506,N_4143,N_4061);
or U4507 (N_4507,N_4045,N_3873);
nand U4508 (N_4508,N_3829,N_3837);
or U4509 (N_4509,N_3790,N_3789);
and U4510 (N_4510,N_4269,N_4043);
nand U4511 (N_4511,N_4266,N_4364);
xor U4512 (N_4512,N_3932,N_4149);
nand U4513 (N_4513,N_4322,N_3785);
nor U4514 (N_4514,N_4094,N_4077);
and U4515 (N_4515,N_3991,N_4238);
nor U4516 (N_4516,N_4150,N_4186);
nand U4517 (N_4517,N_3902,N_4014);
nand U4518 (N_4518,N_4136,N_4130);
and U4519 (N_4519,N_3976,N_3934);
xnor U4520 (N_4520,N_4317,N_4236);
xor U4521 (N_4521,N_4095,N_4034);
xnor U4522 (N_4522,N_3896,N_3757);
xor U4523 (N_4523,N_4100,N_4287);
and U4524 (N_4524,N_3949,N_3995);
or U4525 (N_4525,N_3961,N_4028);
xnor U4526 (N_4526,N_4357,N_3912);
xor U4527 (N_4527,N_3801,N_4365);
or U4528 (N_4528,N_4128,N_4015);
or U4529 (N_4529,N_4340,N_4358);
nor U4530 (N_4530,N_4328,N_4174);
nand U4531 (N_4531,N_3761,N_4175);
and U4532 (N_4532,N_3982,N_3870);
nand U4533 (N_4533,N_4097,N_3913);
xor U4534 (N_4534,N_4305,N_4222);
or U4535 (N_4535,N_4344,N_3895);
nand U4536 (N_4536,N_4197,N_4113);
nor U4537 (N_4537,N_4350,N_4145);
and U4538 (N_4538,N_4321,N_4055);
nor U4539 (N_4539,N_4304,N_4207);
or U4540 (N_4540,N_4323,N_4178);
and U4541 (N_4541,N_4368,N_3786);
and U4542 (N_4542,N_3851,N_3917);
and U4543 (N_4543,N_3774,N_3994);
nor U4544 (N_4544,N_3845,N_4308);
nor U4545 (N_4545,N_3828,N_4142);
nand U4546 (N_4546,N_3841,N_4258);
nand U4547 (N_4547,N_4144,N_4347);
nor U4548 (N_4548,N_4121,N_4286);
or U4549 (N_4549,N_4162,N_4276);
and U4550 (N_4550,N_3782,N_4176);
or U4551 (N_4551,N_3804,N_4216);
and U4552 (N_4552,N_3964,N_3753);
and U4553 (N_4553,N_4218,N_4146);
nand U4554 (N_4554,N_4147,N_4132);
or U4555 (N_4555,N_3919,N_4127);
nor U4556 (N_4556,N_3788,N_4351);
xor U4557 (N_4557,N_4017,N_3986);
nand U4558 (N_4558,N_3885,N_4227);
nor U4559 (N_4559,N_4041,N_3817);
nand U4560 (N_4560,N_3928,N_3992);
nor U4561 (N_4561,N_4109,N_3858);
xor U4562 (N_4562,N_4148,N_4129);
nor U4563 (N_4563,N_4172,N_3850);
nand U4564 (N_4564,N_4031,N_3959);
or U4565 (N_4565,N_3956,N_3783);
or U4566 (N_4566,N_3809,N_4208);
and U4567 (N_4567,N_3948,N_4114);
xnor U4568 (N_4568,N_3848,N_3750);
nand U4569 (N_4569,N_4032,N_3883);
or U4570 (N_4570,N_3811,N_4044);
nand U4571 (N_4571,N_3859,N_3756);
and U4572 (N_4572,N_4268,N_4062);
or U4573 (N_4573,N_3794,N_3876);
xor U4574 (N_4574,N_3833,N_3773);
or U4575 (N_4575,N_4355,N_3874);
nand U4576 (N_4576,N_4297,N_4125);
xor U4577 (N_4577,N_3863,N_4273);
xnor U4578 (N_4578,N_3763,N_4159);
xor U4579 (N_4579,N_3922,N_4303);
nand U4580 (N_4580,N_4234,N_3808);
nand U4581 (N_4581,N_4251,N_4082);
xor U4582 (N_4582,N_3840,N_3925);
xnor U4583 (N_4583,N_4279,N_3824);
or U4584 (N_4584,N_4291,N_4289);
nor U4585 (N_4585,N_4252,N_4271);
and U4586 (N_4586,N_3937,N_4068);
nand U4587 (N_4587,N_4219,N_3820);
nor U4588 (N_4588,N_4185,N_3764);
and U4589 (N_4589,N_3767,N_4352);
or U4590 (N_4590,N_4356,N_4248);
or U4591 (N_4591,N_3990,N_3926);
nand U4592 (N_4592,N_4213,N_3935);
nand U4593 (N_4593,N_4134,N_3864);
xor U4594 (N_4594,N_3814,N_4298);
or U4595 (N_4595,N_3879,N_4069);
xnor U4596 (N_4596,N_3945,N_3916);
xor U4597 (N_4597,N_4083,N_4177);
xnor U4598 (N_4598,N_3906,N_4140);
nand U4599 (N_4599,N_4024,N_3758);
nand U4600 (N_4600,N_4029,N_4042);
xor U4601 (N_4601,N_4005,N_4078);
nor U4602 (N_4602,N_3827,N_3910);
xnor U4603 (N_4603,N_4089,N_3984);
nand U4604 (N_4604,N_3755,N_4359);
or U4605 (N_4605,N_4118,N_4073);
nand U4606 (N_4606,N_3857,N_4008);
and U4607 (N_4607,N_3854,N_3843);
nand U4608 (N_4608,N_4092,N_4249);
and U4609 (N_4609,N_3979,N_4281);
xnor U4610 (N_4610,N_3766,N_3957);
xor U4611 (N_4611,N_4335,N_3980);
xor U4612 (N_4612,N_3954,N_3983);
xnor U4613 (N_4613,N_3931,N_3886);
xnor U4614 (N_4614,N_4156,N_3993);
nor U4615 (N_4615,N_4035,N_3772);
xnor U4616 (N_4616,N_4027,N_3939);
nor U4617 (N_4617,N_3958,N_3941);
nor U4618 (N_4618,N_4261,N_3881);
nand U4619 (N_4619,N_3998,N_4250);
and U4620 (N_4620,N_3893,N_3867);
xnor U4621 (N_4621,N_4228,N_4120);
and U4622 (N_4622,N_4210,N_4315);
nand U4623 (N_4623,N_4104,N_3978);
nor U4624 (N_4624,N_4288,N_4313);
xor U4625 (N_4625,N_4050,N_4065);
xnor U4626 (N_4626,N_4254,N_3914);
xor U4627 (N_4627,N_4138,N_4373);
nand U4628 (N_4628,N_4191,N_4179);
xor U4629 (N_4629,N_4307,N_4166);
and U4630 (N_4630,N_3888,N_4194);
or U4631 (N_4631,N_4198,N_4193);
xnor U4632 (N_4632,N_4369,N_4003);
and U4633 (N_4633,N_3838,N_4302);
nand U4634 (N_4634,N_3903,N_4064);
nand U4635 (N_4635,N_4119,N_4105);
nor U4636 (N_4636,N_4244,N_4098);
or U4637 (N_4637,N_3872,N_3965);
nor U4638 (N_4638,N_3915,N_4203);
xnor U4639 (N_4639,N_4180,N_4205);
and U4640 (N_4640,N_3768,N_4263);
or U4641 (N_4641,N_4343,N_4220);
xor U4642 (N_4642,N_4038,N_4224);
nor U4643 (N_4643,N_4354,N_3920);
or U4644 (N_4644,N_3792,N_4232);
nand U4645 (N_4645,N_4363,N_3955);
xor U4646 (N_4646,N_3884,N_4071);
xnor U4647 (N_4647,N_3819,N_4214);
nand U4648 (N_4648,N_4341,N_4181);
or U4649 (N_4649,N_3796,N_3868);
or U4650 (N_4650,N_3894,N_4010);
nand U4651 (N_4651,N_4262,N_4002);
nor U4652 (N_4652,N_4257,N_4037);
xnor U4653 (N_4653,N_4123,N_4372);
nor U4654 (N_4654,N_3871,N_4316);
nor U4655 (N_4655,N_4000,N_4170);
or U4656 (N_4656,N_4026,N_3877);
nor U4657 (N_4657,N_4255,N_3847);
nand U4658 (N_4658,N_4047,N_4103);
and U4659 (N_4659,N_4139,N_4349);
or U4660 (N_4660,N_3852,N_4004);
and U4661 (N_4661,N_4190,N_4256);
nor U4662 (N_4662,N_3878,N_3891);
or U4663 (N_4663,N_4161,N_4221);
nor U4664 (N_4664,N_4160,N_4265);
or U4665 (N_4665,N_4235,N_3909);
nor U4666 (N_4666,N_4270,N_3797);
nor U4667 (N_4667,N_3869,N_4060);
and U4668 (N_4668,N_4199,N_4296);
nor U4669 (N_4669,N_4112,N_4225);
nand U4670 (N_4670,N_3807,N_4314);
nor U4671 (N_4671,N_3963,N_3806);
xnor U4672 (N_4672,N_4063,N_4013);
nor U4673 (N_4673,N_3971,N_3769);
nand U4674 (N_4674,N_4329,N_3793);
and U4675 (N_4675,N_3795,N_4133);
nand U4676 (N_4676,N_3822,N_4309);
and U4677 (N_4677,N_3968,N_3860);
nand U4678 (N_4678,N_4108,N_4285);
xnor U4679 (N_4679,N_3887,N_4371);
nor U4680 (N_4680,N_4154,N_3921);
or U4681 (N_4681,N_3985,N_3977);
and U4682 (N_4682,N_3933,N_4076);
xor U4683 (N_4683,N_3973,N_3907);
and U4684 (N_4684,N_4201,N_3987);
nor U4685 (N_4685,N_4188,N_4211);
nand U4686 (N_4686,N_3831,N_4070);
nand U4687 (N_4687,N_4333,N_3937);
xnor U4688 (N_4688,N_3750,N_4147);
nand U4689 (N_4689,N_4221,N_3944);
nor U4690 (N_4690,N_4175,N_4354);
or U4691 (N_4691,N_3828,N_3869);
nand U4692 (N_4692,N_3776,N_3797);
or U4693 (N_4693,N_3896,N_4331);
or U4694 (N_4694,N_4116,N_4221);
or U4695 (N_4695,N_4177,N_4206);
nor U4696 (N_4696,N_3833,N_4115);
nand U4697 (N_4697,N_4269,N_4330);
xnor U4698 (N_4698,N_3958,N_4295);
xnor U4699 (N_4699,N_3977,N_3946);
nand U4700 (N_4700,N_4017,N_3771);
xor U4701 (N_4701,N_3884,N_3753);
xor U4702 (N_4702,N_3812,N_4305);
and U4703 (N_4703,N_4135,N_4008);
nand U4704 (N_4704,N_4265,N_4287);
nand U4705 (N_4705,N_4039,N_3924);
and U4706 (N_4706,N_4126,N_3799);
nand U4707 (N_4707,N_4010,N_3795);
nor U4708 (N_4708,N_4252,N_4191);
nor U4709 (N_4709,N_3860,N_3958);
xor U4710 (N_4710,N_3818,N_3876);
nor U4711 (N_4711,N_3961,N_3832);
nand U4712 (N_4712,N_3870,N_4251);
xnor U4713 (N_4713,N_3807,N_3928);
and U4714 (N_4714,N_4365,N_3933);
or U4715 (N_4715,N_4237,N_3912);
xor U4716 (N_4716,N_4298,N_3846);
nor U4717 (N_4717,N_4090,N_3888);
or U4718 (N_4718,N_4144,N_4299);
nand U4719 (N_4719,N_4037,N_4366);
nor U4720 (N_4720,N_3846,N_4127);
xor U4721 (N_4721,N_3875,N_4322);
xnor U4722 (N_4722,N_3802,N_4004);
and U4723 (N_4723,N_3764,N_4297);
nor U4724 (N_4724,N_4187,N_4142);
xnor U4725 (N_4725,N_3819,N_3865);
or U4726 (N_4726,N_4226,N_3928);
nand U4727 (N_4727,N_3751,N_4008);
or U4728 (N_4728,N_3815,N_4135);
or U4729 (N_4729,N_3933,N_4334);
or U4730 (N_4730,N_4373,N_4144);
and U4731 (N_4731,N_3856,N_3918);
xnor U4732 (N_4732,N_4158,N_3921);
or U4733 (N_4733,N_3879,N_3902);
nor U4734 (N_4734,N_4185,N_3767);
nand U4735 (N_4735,N_4352,N_4055);
nor U4736 (N_4736,N_4109,N_4343);
and U4737 (N_4737,N_3796,N_4122);
xor U4738 (N_4738,N_3837,N_4373);
and U4739 (N_4739,N_4266,N_3984);
or U4740 (N_4740,N_4075,N_3853);
or U4741 (N_4741,N_3912,N_4142);
and U4742 (N_4742,N_3915,N_3919);
nand U4743 (N_4743,N_4353,N_3937);
and U4744 (N_4744,N_4115,N_3987);
or U4745 (N_4745,N_3931,N_3932);
nand U4746 (N_4746,N_4346,N_4214);
xnor U4747 (N_4747,N_3887,N_3842);
nand U4748 (N_4748,N_4064,N_3772);
and U4749 (N_4749,N_4095,N_4016);
nor U4750 (N_4750,N_3912,N_4220);
nor U4751 (N_4751,N_3911,N_3902);
nor U4752 (N_4752,N_4029,N_3848);
xor U4753 (N_4753,N_4261,N_4144);
and U4754 (N_4754,N_4259,N_4122);
or U4755 (N_4755,N_4227,N_4058);
or U4756 (N_4756,N_4155,N_3811);
or U4757 (N_4757,N_4161,N_4176);
and U4758 (N_4758,N_3758,N_4164);
and U4759 (N_4759,N_4204,N_4095);
and U4760 (N_4760,N_3773,N_3923);
nor U4761 (N_4761,N_4364,N_4208);
or U4762 (N_4762,N_4149,N_3784);
and U4763 (N_4763,N_3954,N_3843);
nand U4764 (N_4764,N_3810,N_4221);
or U4765 (N_4765,N_3765,N_3932);
xnor U4766 (N_4766,N_4323,N_4205);
or U4767 (N_4767,N_4213,N_4180);
nor U4768 (N_4768,N_3752,N_4306);
xor U4769 (N_4769,N_4010,N_4121);
nor U4770 (N_4770,N_4281,N_4171);
or U4771 (N_4771,N_4101,N_4164);
and U4772 (N_4772,N_3917,N_4087);
and U4773 (N_4773,N_4155,N_3994);
nor U4774 (N_4774,N_4013,N_4167);
nand U4775 (N_4775,N_4076,N_4232);
or U4776 (N_4776,N_3799,N_3844);
or U4777 (N_4777,N_4145,N_3835);
nor U4778 (N_4778,N_3836,N_4265);
nor U4779 (N_4779,N_4006,N_4091);
xnor U4780 (N_4780,N_4277,N_3980);
xnor U4781 (N_4781,N_3849,N_4047);
xnor U4782 (N_4782,N_3775,N_3755);
nand U4783 (N_4783,N_3778,N_4245);
nand U4784 (N_4784,N_4292,N_4160);
or U4785 (N_4785,N_3889,N_4135);
nand U4786 (N_4786,N_3887,N_4292);
xnor U4787 (N_4787,N_3893,N_4269);
xnor U4788 (N_4788,N_3957,N_3883);
and U4789 (N_4789,N_4130,N_3896);
and U4790 (N_4790,N_3771,N_4370);
nor U4791 (N_4791,N_4036,N_3961);
xor U4792 (N_4792,N_4102,N_4168);
and U4793 (N_4793,N_4369,N_4361);
nand U4794 (N_4794,N_4055,N_4199);
nand U4795 (N_4795,N_3975,N_4112);
nand U4796 (N_4796,N_4047,N_4105);
and U4797 (N_4797,N_4213,N_4102);
xor U4798 (N_4798,N_3896,N_4205);
and U4799 (N_4799,N_4288,N_4032);
or U4800 (N_4800,N_4085,N_4160);
and U4801 (N_4801,N_3762,N_4257);
xnor U4802 (N_4802,N_4212,N_4170);
xnor U4803 (N_4803,N_4268,N_3885);
nor U4804 (N_4804,N_4018,N_3868);
nand U4805 (N_4805,N_3898,N_3973);
nor U4806 (N_4806,N_4171,N_3827);
xor U4807 (N_4807,N_4287,N_4247);
nor U4808 (N_4808,N_4143,N_3862);
or U4809 (N_4809,N_4244,N_4055);
and U4810 (N_4810,N_3942,N_4040);
xnor U4811 (N_4811,N_4026,N_4086);
xnor U4812 (N_4812,N_3939,N_3791);
nor U4813 (N_4813,N_4342,N_3919);
nor U4814 (N_4814,N_4085,N_4213);
xor U4815 (N_4815,N_4315,N_4352);
nand U4816 (N_4816,N_3756,N_3842);
or U4817 (N_4817,N_4050,N_3835);
and U4818 (N_4818,N_4186,N_4220);
xor U4819 (N_4819,N_4012,N_4021);
or U4820 (N_4820,N_4000,N_4363);
xnor U4821 (N_4821,N_4136,N_3839);
nor U4822 (N_4822,N_3842,N_3846);
nand U4823 (N_4823,N_4224,N_4322);
and U4824 (N_4824,N_3945,N_4002);
xor U4825 (N_4825,N_4155,N_4217);
nand U4826 (N_4826,N_3907,N_4264);
nand U4827 (N_4827,N_3930,N_3989);
or U4828 (N_4828,N_4205,N_4057);
nor U4829 (N_4829,N_4275,N_3833);
nand U4830 (N_4830,N_3866,N_4223);
xor U4831 (N_4831,N_3768,N_4334);
nand U4832 (N_4832,N_4121,N_4289);
and U4833 (N_4833,N_4046,N_3983);
or U4834 (N_4834,N_4037,N_3976);
or U4835 (N_4835,N_4068,N_4100);
and U4836 (N_4836,N_4325,N_4048);
nand U4837 (N_4837,N_3787,N_4187);
or U4838 (N_4838,N_3896,N_4183);
or U4839 (N_4839,N_3905,N_4339);
and U4840 (N_4840,N_4326,N_3816);
or U4841 (N_4841,N_4008,N_4101);
or U4842 (N_4842,N_3909,N_4357);
xor U4843 (N_4843,N_4030,N_4128);
nand U4844 (N_4844,N_3790,N_4041);
nor U4845 (N_4845,N_4067,N_4103);
nor U4846 (N_4846,N_4099,N_3924);
nor U4847 (N_4847,N_4010,N_3898);
or U4848 (N_4848,N_3884,N_3938);
xor U4849 (N_4849,N_4279,N_3814);
nor U4850 (N_4850,N_3814,N_4248);
and U4851 (N_4851,N_4373,N_4287);
nor U4852 (N_4852,N_3882,N_4201);
nor U4853 (N_4853,N_3842,N_4296);
nor U4854 (N_4854,N_4080,N_4302);
nand U4855 (N_4855,N_3924,N_4231);
or U4856 (N_4856,N_3998,N_4063);
xor U4857 (N_4857,N_3762,N_4103);
nor U4858 (N_4858,N_3930,N_4215);
nand U4859 (N_4859,N_4316,N_3999);
xnor U4860 (N_4860,N_3956,N_3852);
xnor U4861 (N_4861,N_3989,N_4034);
or U4862 (N_4862,N_3885,N_4336);
xnor U4863 (N_4863,N_4064,N_4363);
or U4864 (N_4864,N_4265,N_4137);
xor U4865 (N_4865,N_3835,N_4022);
and U4866 (N_4866,N_3905,N_4328);
xnor U4867 (N_4867,N_4284,N_4148);
and U4868 (N_4868,N_4235,N_3752);
nor U4869 (N_4869,N_3914,N_4250);
and U4870 (N_4870,N_4196,N_4218);
or U4871 (N_4871,N_4063,N_3951);
nor U4872 (N_4872,N_4062,N_3840);
nor U4873 (N_4873,N_4242,N_4325);
and U4874 (N_4874,N_4126,N_3821);
nor U4875 (N_4875,N_3959,N_3805);
nand U4876 (N_4876,N_3970,N_3987);
nor U4877 (N_4877,N_4233,N_4351);
xor U4878 (N_4878,N_3982,N_4277);
or U4879 (N_4879,N_4227,N_3939);
nand U4880 (N_4880,N_3949,N_4215);
nor U4881 (N_4881,N_4235,N_3893);
and U4882 (N_4882,N_3894,N_4019);
nand U4883 (N_4883,N_4319,N_4188);
or U4884 (N_4884,N_4251,N_4090);
and U4885 (N_4885,N_4004,N_4201);
nor U4886 (N_4886,N_3954,N_3865);
and U4887 (N_4887,N_3988,N_4312);
nand U4888 (N_4888,N_4113,N_3829);
and U4889 (N_4889,N_3768,N_3896);
nand U4890 (N_4890,N_3901,N_4181);
nand U4891 (N_4891,N_4344,N_4311);
and U4892 (N_4892,N_4078,N_4025);
nand U4893 (N_4893,N_4055,N_3752);
nand U4894 (N_4894,N_4184,N_4007);
and U4895 (N_4895,N_4031,N_3955);
or U4896 (N_4896,N_3957,N_3781);
nand U4897 (N_4897,N_3869,N_4035);
or U4898 (N_4898,N_4202,N_4199);
or U4899 (N_4899,N_3925,N_4074);
xnor U4900 (N_4900,N_4338,N_4358);
nor U4901 (N_4901,N_4293,N_4127);
xnor U4902 (N_4902,N_4137,N_4058);
nor U4903 (N_4903,N_3892,N_4332);
or U4904 (N_4904,N_3897,N_4370);
nand U4905 (N_4905,N_4321,N_4269);
nor U4906 (N_4906,N_4071,N_4313);
or U4907 (N_4907,N_3986,N_4110);
xnor U4908 (N_4908,N_4166,N_3793);
or U4909 (N_4909,N_3919,N_4089);
xor U4910 (N_4910,N_3819,N_4139);
nor U4911 (N_4911,N_4368,N_3864);
or U4912 (N_4912,N_4147,N_4023);
or U4913 (N_4913,N_4253,N_3958);
xor U4914 (N_4914,N_4271,N_4185);
or U4915 (N_4915,N_4111,N_4086);
nand U4916 (N_4916,N_3957,N_4158);
nor U4917 (N_4917,N_3982,N_4265);
nand U4918 (N_4918,N_4132,N_3959);
and U4919 (N_4919,N_4146,N_4264);
xnor U4920 (N_4920,N_4185,N_3758);
or U4921 (N_4921,N_4343,N_3782);
nor U4922 (N_4922,N_4305,N_4114);
xnor U4923 (N_4923,N_4289,N_4349);
xnor U4924 (N_4924,N_4029,N_4352);
nor U4925 (N_4925,N_4057,N_4207);
nand U4926 (N_4926,N_4076,N_3822);
and U4927 (N_4927,N_4263,N_4196);
and U4928 (N_4928,N_4107,N_4317);
nand U4929 (N_4929,N_3758,N_4050);
and U4930 (N_4930,N_4326,N_4234);
nand U4931 (N_4931,N_4335,N_4092);
nor U4932 (N_4932,N_4331,N_4329);
nand U4933 (N_4933,N_4305,N_3884);
xnor U4934 (N_4934,N_3831,N_4348);
or U4935 (N_4935,N_4068,N_3759);
nor U4936 (N_4936,N_4313,N_4133);
and U4937 (N_4937,N_4242,N_3818);
xor U4938 (N_4938,N_4148,N_3843);
and U4939 (N_4939,N_3979,N_3875);
nor U4940 (N_4940,N_4083,N_4171);
and U4941 (N_4941,N_3933,N_4200);
or U4942 (N_4942,N_3820,N_4127);
xor U4943 (N_4943,N_3928,N_4293);
xnor U4944 (N_4944,N_3786,N_3894);
nand U4945 (N_4945,N_3996,N_4138);
nand U4946 (N_4946,N_4071,N_3876);
and U4947 (N_4947,N_4367,N_4285);
nand U4948 (N_4948,N_4176,N_3814);
or U4949 (N_4949,N_4193,N_3788);
xor U4950 (N_4950,N_3854,N_3786);
xor U4951 (N_4951,N_3995,N_3765);
xnor U4952 (N_4952,N_4024,N_4351);
or U4953 (N_4953,N_3914,N_4129);
nand U4954 (N_4954,N_4057,N_4075);
and U4955 (N_4955,N_3818,N_3907);
nor U4956 (N_4956,N_4284,N_4083);
xor U4957 (N_4957,N_4272,N_3999);
nand U4958 (N_4958,N_4125,N_3856);
nand U4959 (N_4959,N_3817,N_3948);
or U4960 (N_4960,N_3769,N_4192);
or U4961 (N_4961,N_4356,N_4144);
and U4962 (N_4962,N_3760,N_3951);
nor U4963 (N_4963,N_4297,N_4111);
nor U4964 (N_4964,N_3761,N_4090);
xnor U4965 (N_4965,N_3934,N_3829);
nor U4966 (N_4966,N_4265,N_4331);
or U4967 (N_4967,N_3757,N_4276);
nor U4968 (N_4968,N_4225,N_4272);
and U4969 (N_4969,N_4279,N_4102);
nor U4970 (N_4970,N_3833,N_4256);
xor U4971 (N_4971,N_4061,N_4212);
and U4972 (N_4972,N_3996,N_4038);
or U4973 (N_4973,N_4355,N_4080);
nor U4974 (N_4974,N_4124,N_4200);
or U4975 (N_4975,N_4139,N_3906);
nand U4976 (N_4976,N_4232,N_4024);
nor U4977 (N_4977,N_4358,N_3889);
and U4978 (N_4978,N_3983,N_4340);
xor U4979 (N_4979,N_4023,N_3951);
xor U4980 (N_4980,N_3951,N_3876);
nand U4981 (N_4981,N_3753,N_4248);
and U4982 (N_4982,N_4265,N_4294);
nor U4983 (N_4983,N_4236,N_4193);
xnor U4984 (N_4984,N_3967,N_4003);
or U4985 (N_4985,N_4257,N_3855);
xor U4986 (N_4986,N_3804,N_4339);
nor U4987 (N_4987,N_3935,N_4350);
and U4988 (N_4988,N_4155,N_4218);
xor U4989 (N_4989,N_4299,N_4166);
nor U4990 (N_4990,N_4180,N_4080);
and U4991 (N_4991,N_3892,N_4182);
nand U4992 (N_4992,N_3923,N_4035);
and U4993 (N_4993,N_3795,N_4243);
nand U4994 (N_4994,N_3988,N_3841);
xor U4995 (N_4995,N_3883,N_3909);
and U4996 (N_4996,N_4001,N_3873);
nand U4997 (N_4997,N_4171,N_3882);
or U4998 (N_4998,N_4210,N_4013);
and U4999 (N_4999,N_4103,N_4071);
and U5000 (N_5000,N_4620,N_4770);
xor U5001 (N_5001,N_4919,N_4767);
or U5002 (N_5002,N_4570,N_4898);
xnor U5003 (N_5003,N_4588,N_4580);
and U5004 (N_5004,N_4894,N_4934);
and U5005 (N_5005,N_4468,N_4702);
xor U5006 (N_5006,N_4715,N_4523);
or U5007 (N_5007,N_4509,N_4382);
or U5008 (N_5008,N_4585,N_4577);
or U5009 (N_5009,N_4976,N_4911);
and U5010 (N_5010,N_4895,N_4747);
and U5011 (N_5011,N_4482,N_4410);
nand U5012 (N_5012,N_4994,N_4875);
and U5013 (N_5013,N_4579,N_4662);
nand U5014 (N_5014,N_4917,N_4874);
nand U5015 (N_5015,N_4800,N_4700);
xnor U5016 (N_5016,N_4415,N_4461);
and U5017 (N_5017,N_4560,N_4479);
nor U5018 (N_5018,N_4661,N_4707);
nor U5019 (N_5019,N_4780,N_4634);
or U5020 (N_5020,N_4591,N_4690);
nor U5021 (N_5021,N_4996,N_4948);
and U5022 (N_5022,N_4838,N_4613);
nor U5023 (N_5023,N_4398,N_4547);
nor U5024 (N_5024,N_4553,N_4563);
or U5025 (N_5025,N_4820,N_4552);
nand U5026 (N_5026,N_4982,N_4471);
nor U5027 (N_5027,N_4896,N_4678);
nor U5028 (N_5028,N_4663,N_4670);
or U5029 (N_5029,N_4947,N_4392);
and U5030 (N_5030,N_4564,N_4680);
nor U5031 (N_5031,N_4604,N_4644);
or U5032 (N_5032,N_4951,N_4512);
xnor U5033 (N_5033,N_4386,N_4477);
and U5034 (N_5034,N_4501,N_4754);
xnor U5035 (N_5035,N_4544,N_4836);
nand U5036 (N_5036,N_4810,N_4759);
and U5037 (N_5037,N_4799,N_4632);
and U5038 (N_5038,N_4495,N_4883);
or U5039 (N_5039,N_4457,N_4961);
and U5040 (N_5040,N_4945,N_4614);
and U5041 (N_5041,N_4744,N_4757);
xnor U5042 (N_5042,N_4381,N_4658);
nor U5043 (N_5043,N_4722,N_4655);
nor U5044 (N_5044,N_4387,N_4912);
and U5045 (N_5045,N_4651,N_4992);
nand U5046 (N_5046,N_4854,N_4921);
nand U5047 (N_5047,N_4904,N_4397);
nor U5048 (N_5048,N_4531,N_4646);
nand U5049 (N_5049,N_4454,N_4877);
xnor U5050 (N_5050,N_4955,N_4782);
xnor U5051 (N_5051,N_4498,N_4652);
or U5052 (N_5052,N_4411,N_4803);
and U5053 (N_5053,N_4428,N_4882);
xnor U5054 (N_5054,N_4638,N_4606);
or U5055 (N_5055,N_4811,N_4872);
and U5056 (N_5056,N_4953,N_4740);
and U5057 (N_5057,N_4970,N_4944);
nand U5058 (N_5058,N_4657,N_4987);
nor U5059 (N_5059,N_4698,N_4407);
xnor U5060 (N_5060,N_4907,N_4485);
nor U5061 (N_5061,N_4504,N_4633);
or U5062 (N_5062,N_4596,N_4781);
nand U5063 (N_5063,N_4988,N_4396);
xnor U5064 (N_5064,N_4460,N_4764);
nand U5065 (N_5065,N_4593,N_4624);
and U5066 (N_5066,N_4816,N_4536);
xnor U5067 (N_5067,N_4419,N_4888);
xor U5068 (N_5068,N_4809,N_4611);
xor U5069 (N_5069,N_4727,N_4629);
xor U5070 (N_5070,N_4760,N_4761);
xor U5071 (N_5071,N_4738,N_4766);
or U5072 (N_5072,N_4659,N_4557);
and U5073 (N_5073,N_4926,N_4422);
xnor U5074 (N_5074,N_4431,N_4795);
nor U5075 (N_5075,N_4984,N_4493);
xor U5076 (N_5076,N_4699,N_4693);
xor U5077 (N_5077,N_4941,N_4494);
nand U5078 (N_5078,N_4516,N_4607);
nor U5079 (N_5079,N_4960,N_4434);
or U5080 (N_5080,N_4551,N_4681);
nand U5081 (N_5081,N_4418,N_4685);
nor U5082 (N_5082,N_4807,N_4584);
and U5083 (N_5083,N_4432,N_4814);
or U5084 (N_5084,N_4804,N_4384);
and U5085 (N_5085,N_4393,N_4910);
or U5086 (N_5086,N_4676,N_4447);
nand U5087 (N_5087,N_4927,N_4840);
or U5088 (N_5088,N_4899,N_4426);
nor U5089 (N_5089,N_4435,N_4576);
nor U5090 (N_5090,N_4842,N_4409);
nor U5091 (N_5091,N_4540,N_4445);
or U5092 (N_5092,N_4880,N_4954);
and U5093 (N_5093,N_4828,N_4390);
nand U5094 (N_5094,N_4776,N_4403);
nor U5095 (N_5095,N_4790,N_4515);
or U5096 (N_5096,N_4873,N_4949);
and U5097 (N_5097,N_4891,N_4753);
and U5098 (N_5098,N_4714,N_4789);
nand U5099 (N_5099,N_4510,N_4908);
xor U5100 (N_5100,N_4731,N_4855);
and U5101 (N_5101,N_4935,N_4721);
nor U5102 (N_5102,N_4723,N_4379);
and U5103 (N_5103,N_4710,N_4687);
xor U5104 (N_5104,N_4733,N_4443);
nor U5105 (N_5105,N_4528,N_4535);
nor U5106 (N_5106,N_4548,N_4959);
xor U5107 (N_5107,N_4656,N_4466);
and U5108 (N_5108,N_4946,N_4826);
xnor U5109 (N_5109,N_4973,N_4413);
nor U5110 (N_5110,N_4550,N_4859);
or U5111 (N_5111,N_4701,N_4725);
and U5112 (N_5112,N_4694,N_4441);
or U5113 (N_5113,N_4666,N_4871);
or U5114 (N_5114,N_4446,N_4546);
nor U5115 (N_5115,N_4845,N_4476);
xnor U5116 (N_5116,N_4487,N_4755);
xor U5117 (N_5117,N_4879,N_4712);
nand U5118 (N_5118,N_4451,N_4602);
xnor U5119 (N_5119,N_4705,N_4488);
xor U5120 (N_5120,N_4601,N_4915);
or U5121 (N_5121,N_4470,N_4672);
xor U5122 (N_5122,N_4503,N_4756);
or U5123 (N_5123,N_4818,N_4650);
and U5124 (N_5124,N_4566,N_4985);
nand U5125 (N_5125,N_4572,N_4983);
nor U5126 (N_5126,N_4968,N_4892);
nand U5127 (N_5127,N_4438,N_4928);
or U5128 (N_5128,N_4555,N_4682);
nand U5129 (N_5129,N_4711,N_4545);
and U5130 (N_5130,N_4376,N_4936);
or U5131 (N_5131,N_4797,N_4957);
and U5132 (N_5132,N_4905,N_4683);
nand U5133 (N_5133,N_4724,N_4796);
xor U5134 (N_5134,N_4554,N_4497);
nor U5135 (N_5135,N_4843,N_4444);
nand U5136 (N_5136,N_4929,N_4886);
and U5137 (N_5137,N_4956,N_4631);
nand U5138 (N_5138,N_4743,N_4783);
and U5139 (N_5139,N_4716,N_4395);
nor U5140 (N_5140,N_4508,N_4605);
nand U5141 (N_5141,N_4537,N_4452);
xor U5142 (N_5142,N_4639,N_4442);
and U5143 (N_5143,N_4459,N_4831);
xnor U5144 (N_5144,N_4742,N_4610);
and U5145 (N_5145,N_4645,N_4677);
nand U5146 (N_5146,N_4745,N_4616);
and U5147 (N_5147,N_4401,N_4514);
xnor U5148 (N_5148,N_4771,N_4837);
nand U5149 (N_5149,N_4792,N_4964);
nor U5150 (N_5150,N_4990,N_4785);
nor U5151 (N_5151,N_4590,N_4600);
nor U5152 (N_5152,N_4794,N_4586);
nor U5153 (N_5153,N_4775,N_4385);
nand U5154 (N_5154,N_4408,N_4991);
nand U5155 (N_5155,N_4708,N_4943);
or U5156 (N_5156,N_4865,N_4823);
nor U5157 (N_5157,N_4526,N_4473);
nor U5158 (N_5158,N_4746,N_4621);
nand U5159 (N_5159,N_4925,N_4541);
xor U5160 (N_5160,N_4784,N_4587);
and U5161 (N_5161,N_4965,N_4399);
xnor U5162 (N_5162,N_4768,N_4664);
and U5163 (N_5163,N_4749,N_4862);
nand U5164 (N_5164,N_4900,N_4686);
xnor U5165 (N_5165,N_4997,N_4730);
nand U5166 (N_5166,N_4518,N_4825);
and U5167 (N_5167,N_4732,N_4618);
xor U5168 (N_5168,N_4913,N_4542);
and U5169 (N_5169,N_4706,N_4671);
and U5170 (N_5170,N_4932,N_4801);
or U5171 (N_5171,N_4822,N_4846);
nand U5172 (N_5172,N_4832,N_4748);
nand U5173 (N_5173,N_4806,N_4737);
nor U5174 (N_5174,N_4808,N_4425);
nor U5175 (N_5175,N_4532,N_4647);
nor U5176 (N_5176,N_4567,N_4713);
and U5177 (N_5177,N_4923,N_4841);
or U5178 (N_5178,N_4405,N_4417);
nor U5179 (N_5179,N_4649,N_4857);
and U5180 (N_5180,N_4424,N_4617);
xnor U5181 (N_5181,N_4868,N_4971);
nor U5182 (N_5182,N_4974,N_4480);
nand U5183 (N_5183,N_4615,N_4967);
xnor U5184 (N_5184,N_4918,N_4769);
nor U5185 (N_5185,N_4628,N_4937);
or U5186 (N_5186,N_4852,N_4958);
xor U5187 (N_5187,N_4375,N_4522);
and U5188 (N_5188,N_4718,N_4430);
or U5189 (N_5189,N_4709,N_4599);
xnor U5190 (N_5190,N_4952,N_4582);
nand U5191 (N_5191,N_4734,N_4692);
or U5192 (N_5192,N_4429,N_4870);
nand U5193 (N_5193,N_4561,N_4674);
xor U5194 (N_5194,N_4993,N_4995);
nand U5195 (N_5195,N_4890,N_4729);
or U5196 (N_5196,N_4455,N_4612);
nor U5197 (N_5197,N_4777,N_4450);
or U5198 (N_5198,N_4848,N_4653);
xor U5199 (N_5199,N_4660,N_4830);
nor U5200 (N_5200,N_4787,N_4630);
xor U5201 (N_5201,N_4589,N_4404);
nand U5202 (N_5202,N_4719,N_4758);
or U5203 (N_5203,N_4774,N_4641);
nand U5204 (N_5204,N_4433,N_4697);
and U5205 (N_5205,N_4920,N_4463);
nand U5206 (N_5206,N_4458,N_4668);
xnor U5207 (N_5207,N_4999,N_4977);
xor U5208 (N_5208,N_4665,N_4981);
nand U5209 (N_5209,N_4608,N_4829);
xor U5210 (N_5210,N_4583,N_4568);
nor U5211 (N_5211,N_4813,N_4380);
nor U5212 (N_5212,N_4798,N_4578);
xor U5213 (N_5213,N_4884,N_4978);
and U5214 (N_5214,N_4394,N_4619);
nor U5215 (N_5215,N_4812,N_4691);
and U5216 (N_5216,N_4924,N_4623);
nor U5217 (N_5217,N_4565,N_4728);
xnor U5218 (N_5218,N_4939,N_4648);
and U5219 (N_5219,N_4496,N_4817);
xnor U5220 (N_5220,N_4505,N_4673);
xnor U5221 (N_5221,N_4938,N_4517);
or U5222 (N_5222,N_4860,N_4856);
and U5223 (N_5223,N_4834,N_4499);
nor U5224 (N_5224,N_4741,N_4490);
xnor U5225 (N_5225,N_4511,N_4791);
nor U5226 (N_5226,N_4878,N_4881);
and U5227 (N_5227,N_4864,N_4669);
xnor U5228 (N_5228,N_4421,N_4575);
or U5229 (N_5229,N_4867,N_4717);
or U5230 (N_5230,N_4489,N_4689);
nand U5231 (N_5231,N_4998,N_4627);
nor U5232 (N_5232,N_4773,N_4636);
nor U5233 (N_5233,N_4835,N_4556);
nand U5234 (N_5234,N_4484,N_4400);
nand U5235 (N_5235,N_4462,N_4849);
nor U5236 (N_5236,N_4642,N_4427);
and U5237 (N_5237,N_4688,N_4940);
and U5238 (N_5238,N_4412,N_4562);
and U5239 (N_5239,N_4901,N_4750);
or U5240 (N_5240,N_4598,N_4802);
nand U5241 (N_5241,N_4597,N_4377);
or U5242 (N_5242,N_4839,N_4475);
xnor U5243 (N_5243,N_4464,N_4383);
xor U5244 (N_5244,N_4439,N_4833);
nor U5245 (N_5245,N_4861,N_4513);
or U5246 (N_5246,N_4440,N_4569);
xor U5247 (N_5247,N_4696,N_4851);
nor U5248 (N_5248,N_4520,N_4863);
and U5249 (N_5249,N_4388,N_4893);
and U5250 (N_5250,N_4736,N_4695);
nand U5251 (N_5251,N_4772,N_4963);
or U5252 (N_5252,N_4850,N_4595);
xnor U5253 (N_5253,N_4916,N_4474);
nand U5254 (N_5254,N_4975,N_4456);
xnor U5255 (N_5255,N_4472,N_4887);
or U5256 (N_5256,N_4592,N_4530);
nor U5257 (N_5257,N_4966,N_4989);
xnor U5258 (N_5258,N_4469,N_4726);
nand U5259 (N_5259,N_4414,N_4897);
xor U5260 (N_5260,N_4423,N_4558);
nor U5261 (N_5261,N_4391,N_4574);
nor U5262 (N_5262,N_4525,N_4378);
and U5263 (N_5263,N_4765,N_4853);
or U5264 (N_5264,N_4720,N_4524);
nor U5265 (N_5265,N_4762,N_4805);
or U5266 (N_5266,N_4640,N_4885);
and U5267 (N_5267,N_4704,N_4389);
and U5268 (N_5268,N_4559,N_4869);
nor U5269 (N_5269,N_4549,N_4876);
xnor U5270 (N_5270,N_4972,N_4643);
nand U5271 (N_5271,N_4679,N_4406);
or U5272 (N_5272,N_4436,N_4821);
and U5273 (N_5273,N_4483,N_4521);
nor U5274 (N_5274,N_4763,N_4793);
and U5275 (N_5275,N_4622,N_4507);
and U5276 (N_5276,N_4903,N_4635);
nor U5277 (N_5277,N_4573,N_4667);
and U5278 (N_5278,N_4486,N_4684);
nor U5279 (N_5279,N_4779,N_4933);
or U5280 (N_5280,N_4402,N_4625);
xor U5281 (N_5281,N_4527,N_4752);
xnor U5282 (N_5282,N_4739,N_4979);
or U5283 (N_5283,N_4420,N_4778);
nand U5284 (N_5284,N_4931,N_4889);
nand U5285 (N_5285,N_4819,N_4751);
nand U5286 (N_5286,N_4534,N_4827);
or U5287 (N_5287,N_4844,N_4539);
xor U5288 (N_5288,N_4416,N_4788);
and U5289 (N_5289,N_4478,N_4922);
xnor U5290 (N_5290,N_4909,N_4609);
nand U5291 (N_5291,N_4465,N_4594);
xor U5292 (N_5292,N_4654,N_4914);
or U5293 (N_5293,N_4502,N_4467);
nor U5294 (N_5294,N_4491,N_4538);
nand U5295 (N_5295,N_4448,N_4675);
and U5296 (N_5296,N_4533,N_4824);
nand U5297 (N_5297,N_4437,N_4786);
or U5298 (N_5298,N_4506,N_4815);
nand U5299 (N_5299,N_4481,N_4519);
and U5300 (N_5300,N_4902,N_4930);
or U5301 (N_5301,N_4942,N_4986);
and U5302 (N_5302,N_4703,N_4847);
xnor U5303 (N_5303,N_4980,N_4529);
nand U5304 (N_5304,N_4962,N_4626);
and U5305 (N_5305,N_4571,N_4969);
or U5306 (N_5306,N_4543,N_4500);
and U5307 (N_5307,N_4637,N_4906);
nand U5308 (N_5308,N_4603,N_4858);
and U5309 (N_5309,N_4449,N_4950);
nand U5310 (N_5310,N_4492,N_4735);
and U5311 (N_5311,N_4453,N_4581);
xnor U5312 (N_5312,N_4866,N_4744);
nor U5313 (N_5313,N_4745,N_4739);
nor U5314 (N_5314,N_4437,N_4502);
nor U5315 (N_5315,N_4450,N_4519);
and U5316 (N_5316,N_4487,N_4589);
nor U5317 (N_5317,N_4412,N_4815);
xor U5318 (N_5318,N_4419,N_4429);
nor U5319 (N_5319,N_4950,N_4471);
nand U5320 (N_5320,N_4545,N_4714);
nand U5321 (N_5321,N_4667,N_4598);
xor U5322 (N_5322,N_4829,N_4818);
nand U5323 (N_5323,N_4672,N_4600);
nand U5324 (N_5324,N_4768,N_4564);
and U5325 (N_5325,N_4823,N_4976);
and U5326 (N_5326,N_4428,N_4635);
or U5327 (N_5327,N_4994,N_4624);
xor U5328 (N_5328,N_4579,N_4551);
and U5329 (N_5329,N_4461,N_4610);
and U5330 (N_5330,N_4673,N_4853);
or U5331 (N_5331,N_4642,N_4411);
nor U5332 (N_5332,N_4442,N_4928);
nand U5333 (N_5333,N_4451,N_4906);
and U5334 (N_5334,N_4985,N_4493);
nor U5335 (N_5335,N_4808,N_4417);
nor U5336 (N_5336,N_4568,N_4382);
nand U5337 (N_5337,N_4414,N_4906);
nor U5338 (N_5338,N_4543,N_4779);
xor U5339 (N_5339,N_4404,N_4516);
xor U5340 (N_5340,N_4784,N_4939);
and U5341 (N_5341,N_4704,N_4562);
or U5342 (N_5342,N_4401,N_4967);
xor U5343 (N_5343,N_4656,N_4668);
or U5344 (N_5344,N_4802,N_4765);
nand U5345 (N_5345,N_4977,N_4624);
xor U5346 (N_5346,N_4672,N_4708);
nand U5347 (N_5347,N_4611,N_4949);
nand U5348 (N_5348,N_4395,N_4431);
nand U5349 (N_5349,N_4893,N_4650);
and U5350 (N_5350,N_4512,N_4717);
nor U5351 (N_5351,N_4583,N_4508);
xor U5352 (N_5352,N_4591,N_4708);
xor U5353 (N_5353,N_4418,N_4615);
nor U5354 (N_5354,N_4666,N_4916);
or U5355 (N_5355,N_4994,N_4574);
nor U5356 (N_5356,N_4870,N_4688);
nand U5357 (N_5357,N_4618,N_4671);
xnor U5358 (N_5358,N_4743,N_4874);
nor U5359 (N_5359,N_4715,N_4604);
nor U5360 (N_5360,N_4541,N_4927);
xor U5361 (N_5361,N_4423,N_4492);
nor U5362 (N_5362,N_4619,N_4553);
nor U5363 (N_5363,N_4667,N_4988);
xnor U5364 (N_5364,N_4863,N_4947);
or U5365 (N_5365,N_4961,N_4911);
xnor U5366 (N_5366,N_4628,N_4699);
or U5367 (N_5367,N_4917,N_4502);
or U5368 (N_5368,N_4976,N_4537);
nor U5369 (N_5369,N_4752,N_4897);
nand U5370 (N_5370,N_4593,N_4607);
nand U5371 (N_5371,N_4817,N_4881);
nand U5372 (N_5372,N_4938,N_4456);
and U5373 (N_5373,N_4974,N_4809);
and U5374 (N_5374,N_4439,N_4534);
xnor U5375 (N_5375,N_4504,N_4677);
nor U5376 (N_5376,N_4679,N_4584);
and U5377 (N_5377,N_4722,N_4561);
or U5378 (N_5378,N_4746,N_4652);
and U5379 (N_5379,N_4958,N_4900);
and U5380 (N_5380,N_4643,N_4741);
nor U5381 (N_5381,N_4577,N_4573);
nor U5382 (N_5382,N_4429,N_4683);
xor U5383 (N_5383,N_4523,N_4782);
and U5384 (N_5384,N_4917,N_4858);
or U5385 (N_5385,N_4665,N_4765);
xor U5386 (N_5386,N_4613,N_4924);
nand U5387 (N_5387,N_4563,N_4801);
nor U5388 (N_5388,N_4544,N_4650);
or U5389 (N_5389,N_4376,N_4769);
and U5390 (N_5390,N_4764,N_4573);
xor U5391 (N_5391,N_4784,N_4524);
xor U5392 (N_5392,N_4787,N_4385);
xor U5393 (N_5393,N_4737,N_4728);
nand U5394 (N_5394,N_4839,N_4712);
xnor U5395 (N_5395,N_4769,N_4531);
xnor U5396 (N_5396,N_4448,N_4437);
and U5397 (N_5397,N_4443,N_4384);
nand U5398 (N_5398,N_4390,N_4722);
or U5399 (N_5399,N_4938,N_4586);
xnor U5400 (N_5400,N_4971,N_4659);
or U5401 (N_5401,N_4637,N_4854);
nand U5402 (N_5402,N_4457,N_4420);
and U5403 (N_5403,N_4980,N_4595);
and U5404 (N_5404,N_4611,N_4614);
nor U5405 (N_5405,N_4796,N_4755);
xor U5406 (N_5406,N_4696,N_4437);
nand U5407 (N_5407,N_4965,N_4417);
nand U5408 (N_5408,N_4654,N_4376);
xor U5409 (N_5409,N_4826,N_4660);
and U5410 (N_5410,N_4474,N_4706);
and U5411 (N_5411,N_4549,N_4648);
and U5412 (N_5412,N_4823,N_4951);
and U5413 (N_5413,N_4381,N_4419);
and U5414 (N_5414,N_4815,N_4436);
or U5415 (N_5415,N_4744,N_4492);
nor U5416 (N_5416,N_4644,N_4393);
xnor U5417 (N_5417,N_4430,N_4844);
nor U5418 (N_5418,N_4893,N_4927);
nor U5419 (N_5419,N_4757,N_4743);
and U5420 (N_5420,N_4755,N_4853);
xor U5421 (N_5421,N_4697,N_4948);
nor U5422 (N_5422,N_4882,N_4996);
nand U5423 (N_5423,N_4773,N_4580);
nand U5424 (N_5424,N_4810,N_4639);
or U5425 (N_5425,N_4699,N_4651);
nand U5426 (N_5426,N_4893,N_4883);
nand U5427 (N_5427,N_4902,N_4416);
xnor U5428 (N_5428,N_4979,N_4883);
nor U5429 (N_5429,N_4835,N_4846);
nand U5430 (N_5430,N_4418,N_4697);
nand U5431 (N_5431,N_4998,N_4416);
nor U5432 (N_5432,N_4662,N_4638);
nor U5433 (N_5433,N_4616,N_4837);
or U5434 (N_5434,N_4990,N_4984);
xnor U5435 (N_5435,N_4830,N_4549);
or U5436 (N_5436,N_4555,N_4752);
nand U5437 (N_5437,N_4843,N_4434);
or U5438 (N_5438,N_4425,N_4931);
nand U5439 (N_5439,N_4513,N_4925);
or U5440 (N_5440,N_4821,N_4649);
nand U5441 (N_5441,N_4569,N_4736);
nand U5442 (N_5442,N_4392,N_4538);
nor U5443 (N_5443,N_4842,N_4476);
nand U5444 (N_5444,N_4619,N_4631);
or U5445 (N_5445,N_4879,N_4889);
xor U5446 (N_5446,N_4784,N_4674);
xnor U5447 (N_5447,N_4759,N_4614);
or U5448 (N_5448,N_4498,N_4456);
xnor U5449 (N_5449,N_4875,N_4644);
nand U5450 (N_5450,N_4653,N_4487);
nor U5451 (N_5451,N_4910,N_4588);
xnor U5452 (N_5452,N_4831,N_4734);
or U5453 (N_5453,N_4996,N_4766);
or U5454 (N_5454,N_4548,N_4889);
nor U5455 (N_5455,N_4823,N_4399);
or U5456 (N_5456,N_4762,N_4458);
nor U5457 (N_5457,N_4954,N_4446);
xor U5458 (N_5458,N_4563,N_4873);
xnor U5459 (N_5459,N_4436,N_4614);
and U5460 (N_5460,N_4493,N_4837);
nor U5461 (N_5461,N_4863,N_4790);
and U5462 (N_5462,N_4854,N_4817);
or U5463 (N_5463,N_4807,N_4836);
or U5464 (N_5464,N_4854,N_4729);
or U5465 (N_5465,N_4822,N_4777);
nand U5466 (N_5466,N_4862,N_4659);
nand U5467 (N_5467,N_4411,N_4686);
xor U5468 (N_5468,N_4661,N_4451);
and U5469 (N_5469,N_4791,N_4942);
and U5470 (N_5470,N_4841,N_4898);
xnor U5471 (N_5471,N_4677,N_4791);
or U5472 (N_5472,N_4866,N_4597);
nand U5473 (N_5473,N_4806,N_4872);
nand U5474 (N_5474,N_4828,N_4725);
and U5475 (N_5475,N_4689,N_4763);
nand U5476 (N_5476,N_4580,N_4699);
or U5477 (N_5477,N_4872,N_4563);
nand U5478 (N_5478,N_4950,N_4451);
nand U5479 (N_5479,N_4996,N_4861);
nand U5480 (N_5480,N_4517,N_4931);
nand U5481 (N_5481,N_4607,N_4836);
xor U5482 (N_5482,N_4842,N_4964);
xnor U5483 (N_5483,N_4849,N_4953);
nand U5484 (N_5484,N_4778,N_4437);
nand U5485 (N_5485,N_4700,N_4516);
nor U5486 (N_5486,N_4983,N_4537);
xor U5487 (N_5487,N_4810,N_4407);
or U5488 (N_5488,N_4385,N_4752);
or U5489 (N_5489,N_4503,N_4397);
xnor U5490 (N_5490,N_4514,N_4594);
nand U5491 (N_5491,N_4665,N_4817);
and U5492 (N_5492,N_4382,N_4935);
and U5493 (N_5493,N_4560,N_4687);
xnor U5494 (N_5494,N_4738,N_4897);
or U5495 (N_5495,N_4440,N_4555);
or U5496 (N_5496,N_4762,N_4583);
nor U5497 (N_5497,N_4390,N_4381);
nand U5498 (N_5498,N_4629,N_4838);
and U5499 (N_5499,N_4797,N_4908);
or U5500 (N_5500,N_4791,N_4693);
xor U5501 (N_5501,N_4723,N_4816);
xor U5502 (N_5502,N_4421,N_4470);
or U5503 (N_5503,N_4541,N_4692);
xor U5504 (N_5504,N_4640,N_4528);
or U5505 (N_5505,N_4748,N_4669);
nor U5506 (N_5506,N_4386,N_4738);
nor U5507 (N_5507,N_4581,N_4837);
and U5508 (N_5508,N_4705,N_4741);
nor U5509 (N_5509,N_4583,N_4698);
or U5510 (N_5510,N_4729,N_4850);
nand U5511 (N_5511,N_4464,N_4980);
nand U5512 (N_5512,N_4684,N_4834);
nand U5513 (N_5513,N_4405,N_4536);
nand U5514 (N_5514,N_4557,N_4542);
xnor U5515 (N_5515,N_4950,N_4624);
xnor U5516 (N_5516,N_4573,N_4980);
nor U5517 (N_5517,N_4517,N_4656);
nand U5518 (N_5518,N_4462,N_4882);
nor U5519 (N_5519,N_4445,N_4561);
or U5520 (N_5520,N_4874,N_4673);
or U5521 (N_5521,N_4676,N_4485);
nand U5522 (N_5522,N_4689,N_4948);
nand U5523 (N_5523,N_4686,N_4757);
and U5524 (N_5524,N_4948,N_4576);
and U5525 (N_5525,N_4543,N_4830);
xnor U5526 (N_5526,N_4944,N_4806);
or U5527 (N_5527,N_4949,N_4461);
nor U5528 (N_5528,N_4781,N_4959);
nand U5529 (N_5529,N_4884,N_4870);
nand U5530 (N_5530,N_4376,N_4906);
nand U5531 (N_5531,N_4944,N_4567);
xnor U5532 (N_5532,N_4755,N_4393);
nor U5533 (N_5533,N_4783,N_4396);
and U5534 (N_5534,N_4585,N_4505);
and U5535 (N_5535,N_4408,N_4496);
nor U5536 (N_5536,N_4444,N_4613);
nor U5537 (N_5537,N_4379,N_4592);
nor U5538 (N_5538,N_4949,N_4662);
or U5539 (N_5539,N_4768,N_4419);
xor U5540 (N_5540,N_4671,N_4382);
nor U5541 (N_5541,N_4432,N_4417);
nor U5542 (N_5542,N_4820,N_4729);
or U5543 (N_5543,N_4628,N_4889);
xnor U5544 (N_5544,N_4765,N_4396);
and U5545 (N_5545,N_4730,N_4771);
and U5546 (N_5546,N_4409,N_4990);
xor U5547 (N_5547,N_4940,N_4580);
nand U5548 (N_5548,N_4687,N_4793);
or U5549 (N_5549,N_4929,N_4733);
xor U5550 (N_5550,N_4835,N_4501);
or U5551 (N_5551,N_4442,N_4558);
nand U5552 (N_5552,N_4515,N_4508);
or U5553 (N_5553,N_4687,N_4768);
nand U5554 (N_5554,N_4477,N_4747);
xor U5555 (N_5555,N_4667,N_4726);
or U5556 (N_5556,N_4675,N_4426);
xnor U5557 (N_5557,N_4729,N_4520);
nor U5558 (N_5558,N_4526,N_4794);
and U5559 (N_5559,N_4389,N_4889);
or U5560 (N_5560,N_4442,N_4596);
nand U5561 (N_5561,N_4645,N_4912);
or U5562 (N_5562,N_4734,N_4659);
nand U5563 (N_5563,N_4514,N_4875);
nand U5564 (N_5564,N_4676,N_4564);
and U5565 (N_5565,N_4861,N_4479);
xor U5566 (N_5566,N_4474,N_4589);
nand U5567 (N_5567,N_4455,N_4981);
nor U5568 (N_5568,N_4506,N_4390);
xor U5569 (N_5569,N_4836,N_4751);
xor U5570 (N_5570,N_4729,N_4606);
nand U5571 (N_5571,N_4867,N_4406);
and U5572 (N_5572,N_4768,N_4375);
nor U5573 (N_5573,N_4710,N_4844);
xor U5574 (N_5574,N_4885,N_4406);
xor U5575 (N_5575,N_4862,N_4668);
nand U5576 (N_5576,N_4606,N_4784);
and U5577 (N_5577,N_4413,N_4969);
nor U5578 (N_5578,N_4787,N_4578);
xnor U5579 (N_5579,N_4929,N_4534);
nand U5580 (N_5580,N_4504,N_4973);
nand U5581 (N_5581,N_4966,N_4782);
nor U5582 (N_5582,N_4661,N_4998);
and U5583 (N_5583,N_4573,N_4581);
or U5584 (N_5584,N_4520,N_4582);
nor U5585 (N_5585,N_4845,N_4824);
and U5586 (N_5586,N_4460,N_4686);
nor U5587 (N_5587,N_4466,N_4866);
and U5588 (N_5588,N_4988,N_4420);
and U5589 (N_5589,N_4892,N_4715);
xor U5590 (N_5590,N_4918,N_4890);
and U5591 (N_5591,N_4635,N_4422);
nor U5592 (N_5592,N_4985,N_4788);
nand U5593 (N_5593,N_4860,N_4545);
nand U5594 (N_5594,N_4377,N_4801);
or U5595 (N_5595,N_4960,N_4959);
or U5596 (N_5596,N_4614,N_4990);
or U5597 (N_5597,N_4699,N_4907);
nor U5598 (N_5598,N_4574,N_4400);
and U5599 (N_5599,N_4767,N_4959);
xor U5600 (N_5600,N_4454,N_4479);
or U5601 (N_5601,N_4460,N_4690);
xor U5602 (N_5602,N_4590,N_4621);
xnor U5603 (N_5603,N_4753,N_4602);
nor U5604 (N_5604,N_4688,N_4640);
and U5605 (N_5605,N_4846,N_4753);
and U5606 (N_5606,N_4779,N_4995);
nand U5607 (N_5607,N_4978,N_4587);
nor U5608 (N_5608,N_4776,N_4468);
nand U5609 (N_5609,N_4658,N_4913);
nand U5610 (N_5610,N_4436,N_4459);
and U5611 (N_5611,N_4424,N_4987);
nand U5612 (N_5612,N_4544,N_4413);
or U5613 (N_5613,N_4555,N_4707);
nor U5614 (N_5614,N_4505,N_4999);
nand U5615 (N_5615,N_4899,N_4423);
or U5616 (N_5616,N_4790,N_4654);
and U5617 (N_5617,N_4431,N_4837);
nand U5618 (N_5618,N_4707,N_4406);
xor U5619 (N_5619,N_4720,N_4827);
and U5620 (N_5620,N_4777,N_4569);
and U5621 (N_5621,N_4410,N_4578);
and U5622 (N_5622,N_4655,N_4839);
nand U5623 (N_5623,N_4877,N_4730);
nor U5624 (N_5624,N_4375,N_4720);
or U5625 (N_5625,N_5338,N_5608);
nor U5626 (N_5626,N_5045,N_5326);
or U5627 (N_5627,N_5605,N_5490);
nor U5628 (N_5628,N_5414,N_5455);
xor U5629 (N_5629,N_5537,N_5301);
or U5630 (N_5630,N_5111,N_5117);
xnor U5631 (N_5631,N_5385,N_5059);
nor U5632 (N_5632,N_5554,N_5528);
nor U5633 (N_5633,N_5363,N_5170);
nor U5634 (N_5634,N_5074,N_5478);
or U5635 (N_5635,N_5467,N_5371);
xnor U5636 (N_5636,N_5067,N_5546);
xor U5637 (N_5637,N_5116,N_5163);
xor U5638 (N_5638,N_5173,N_5123);
and U5639 (N_5639,N_5542,N_5539);
and U5640 (N_5640,N_5482,N_5292);
nand U5641 (N_5641,N_5114,N_5598);
or U5642 (N_5642,N_5094,N_5257);
nand U5643 (N_5643,N_5136,N_5193);
nand U5644 (N_5644,N_5535,N_5509);
and U5645 (N_5645,N_5603,N_5079);
xnor U5646 (N_5646,N_5082,N_5147);
and U5647 (N_5647,N_5392,N_5597);
and U5648 (N_5648,N_5453,N_5515);
or U5649 (N_5649,N_5565,N_5017);
and U5650 (N_5650,N_5579,N_5126);
nand U5651 (N_5651,N_5112,N_5167);
nand U5652 (N_5652,N_5459,N_5584);
or U5653 (N_5653,N_5177,N_5236);
xor U5654 (N_5654,N_5374,N_5581);
nand U5655 (N_5655,N_5550,N_5233);
nand U5656 (N_5656,N_5072,N_5344);
and U5657 (N_5657,N_5100,N_5190);
nor U5658 (N_5658,N_5346,N_5533);
or U5659 (N_5659,N_5577,N_5093);
xor U5660 (N_5660,N_5090,N_5355);
xnor U5661 (N_5661,N_5446,N_5360);
and U5662 (N_5662,N_5370,N_5500);
nand U5663 (N_5663,N_5138,N_5336);
xor U5664 (N_5664,N_5569,N_5368);
nand U5665 (N_5665,N_5150,N_5381);
xor U5666 (N_5666,N_5434,N_5510);
nand U5667 (N_5667,N_5599,N_5521);
xor U5668 (N_5668,N_5057,N_5526);
and U5669 (N_5669,N_5578,N_5146);
or U5670 (N_5670,N_5419,N_5293);
xnor U5671 (N_5671,N_5279,N_5408);
nand U5672 (N_5672,N_5042,N_5475);
xor U5673 (N_5673,N_5454,N_5296);
nor U5674 (N_5674,N_5283,N_5372);
and U5675 (N_5675,N_5342,N_5216);
xnor U5676 (N_5676,N_5213,N_5506);
nor U5677 (N_5677,N_5602,N_5243);
xnor U5678 (N_5678,N_5202,N_5396);
or U5679 (N_5679,N_5566,N_5516);
xnor U5680 (N_5680,N_5601,N_5388);
or U5681 (N_5681,N_5558,N_5435);
nor U5682 (N_5682,N_5592,N_5261);
nand U5683 (N_5683,N_5286,N_5472);
nand U5684 (N_5684,N_5483,N_5544);
nand U5685 (N_5685,N_5137,N_5092);
nand U5686 (N_5686,N_5189,N_5530);
nand U5687 (N_5687,N_5125,N_5572);
or U5688 (N_5688,N_5448,N_5259);
or U5689 (N_5689,N_5449,N_5295);
and U5690 (N_5690,N_5540,N_5505);
and U5691 (N_5691,N_5507,N_5549);
or U5692 (N_5692,N_5450,N_5423);
and U5693 (N_5693,N_5149,N_5021);
nor U5694 (N_5694,N_5444,N_5143);
or U5695 (N_5695,N_5054,N_5252);
or U5696 (N_5696,N_5024,N_5386);
nor U5697 (N_5697,N_5442,N_5426);
nand U5698 (N_5698,N_5564,N_5573);
and U5699 (N_5699,N_5560,N_5473);
or U5700 (N_5700,N_5495,N_5347);
xor U5701 (N_5701,N_5181,N_5369);
nand U5702 (N_5702,N_5254,N_5425);
nor U5703 (N_5703,N_5586,N_5618);
nor U5704 (N_5704,N_5310,N_5152);
xnor U5705 (N_5705,N_5334,N_5345);
or U5706 (N_5706,N_5003,N_5348);
or U5707 (N_5707,N_5328,N_5036);
xnor U5708 (N_5708,N_5018,N_5262);
nand U5709 (N_5709,N_5195,N_5489);
or U5710 (N_5710,N_5307,N_5591);
or U5711 (N_5711,N_5184,N_5553);
and U5712 (N_5712,N_5557,N_5140);
xor U5713 (N_5713,N_5161,N_5232);
or U5714 (N_5714,N_5031,N_5337);
nor U5715 (N_5715,N_5231,N_5273);
xnor U5716 (N_5716,N_5617,N_5321);
nand U5717 (N_5717,N_5397,N_5380);
and U5718 (N_5718,N_5356,N_5316);
or U5719 (N_5719,N_5587,N_5044);
xnor U5720 (N_5720,N_5576,N_5314);
nor U5721 (N_5721,N_5413,N_5221);
or U5722 (N_5722,N_5135,N_5128);
xor U5723 (N_5723,N_5352,N_5364);
and U5724 (N_5724,N_5215,N_5005);
or U5725 (N_5725,N_5134,N_5407);
and U5726 (N_5726,N_5623,N_5606);
xor U5727 (N_5727,N_5165,N_5080);
or U5728 (N_5728,N_5375,N_5524);
and U5729 (N_5729,N_5101,N_5154);
nor U5730 (N_5730,N_5520,N_5399);
xor U5731 (N_5731,N_5319,N_5604);
nor U5732 (N_5732,N_5480,N_5272);
nor U5733 (N_5733,N_5494,N_5329);
xnor U5734 (N_5734,N_5308,N_5323);
xor U5735 (N_5735,N_5313,N_5585);
or U5736 (N_5736,N_5561,N_5387);
or U5737 (N_5737,N_5568,N_5162);
nor U5738 (N_5738,N_5452,N_5282);
xor U5739 (N_5739,N_5476,N_5046);
or U5740 (N_5740,N_5619,N_5570);
and U5741 (N_5741,N_5290,N_5098);
xnor U5742 (N_5742,N_5532,N_5029);
nand U5743 (N_5743,N_5513,N_5271);
nand U5744 (N_5744,N_5622,N_5225);
and U5745 (N_5745,N_5353,N_5085);
nor U5746 (N_5746,N_5235,N_5491);
or U5747 (N_5747,N_5103,N_5266);
or U5748 (N_5748,N_5034,N_5188);
nand U5749 (N_5749,N_5304,N_5590);
nor U5750 (N_5750,N_5253,N_5543);
or U5751 (N_5751,N_5120,N_5400);
or U5752 (N_5752,N_5139,N_5595);
xnor U5753 (N_5753,N_5280,N_5268);
nand U5754 (N_5754,N_5501,N_5411);
and U5755 (N_5755,N_5217,N_5027);
xor U5756 (N_5756,N_5518,N_5209);
and U5757 (N_5757,N_5084,N_5479);
nor U5758 (N_5758,N_5600,N_5264);
xnor U5759 (N_5759,N_5324,N_5312);
or U5760 (N_5760,N_5325,N_5499);
nand U5761 (N_5761,N_5060,N_5199);
nand U5762 (N_5762,N_5294,N_5541);
nand U5763 (N_5763,N_5341,N_5456);
and U5764 (N_5764,N_5488,N_5169);
or U5765 (N_5765,N_5095,N_5485);
or U5766 (N_5766,N_5359,N_5358);
nand U5767 (N_5767,N_5153,N_5056);
nor U5768 (N_5768,N_5088,N_5129);
xnor U5769 (N_5769,N_5551,N_5401);
nand U5770 (N_5770,N_5439,N_5200);
nor U5771 (N_5771,N_5234,N_5222);
and U5772 (N_5772,N_5115,N_5192);
nor U5773 (N_5773,N_5545,N_5285);
xnor U5774 (N_5774,N_5350,N_5615);
xnor U5775 (N_5775,N_5620,N_5463);
xnor U5776 (N_5776,N_5119,N_5144);
or U5777 (N_5777,N_5409,N_5208);
nor U5778 (N_5778,N_5429,N_5068);
nand U5779 (N_5779,N_5109,N_5267);
nand U5780 (N_5780,N_5228,N_5251);
and U5781 (N_5781,N_5322,N_5083);
xnor U5782 (N_5782,N_5441,N_5069);
or U5783 (N_5783,N_5269,N_5151);
or U5784 (N_5784,N_5502,N_5405);
nor U5785 (N_5785,N_5365,N_5614);
nand U5786 (N_5786,N_5611,N_5302);
nand U5787 (N_5787,N_5394,N_5504);
nor U5788 (N_5788,N_5062,N_5340);
xor U5789 (N_5789,N_5171,N_5182);
and U5790 (N_5790,N_5023,N_5191);
nor U5791 (N_5791,N_5010,N_5514);
or U5792 (N_5792,N_5206,N_5108);
nand U5793 (N_5793,N_5610,N_5274);
xor U5794 (N_5794,N_5469,N_5053);
xnor U5795 (N_5795,N_5041,N_5168);
and U5796 (N_5796,N_5536,N_5327);
or U5797 (N_5797,N_5404,N_5297);
and U5798 (N_5798,N_5461,N_5354);
or U5799 (N_5799,N_5025,N_5107);
nor U5800 (N_5800,N_5220,N_5175);
and U5801 (N_5801,N_5012,N_5582);
nand U5802 (N_5802,N_5527,N_5007);
nor U5803 (N_5803,N_5052,N_5097);
or U5804 (N_5804,N_5159,N_5481);
or U5805 (N_5805,N_5204,N_5548);
xor U5806 (N_5806,N_5214,N_5180);
xnor U5807 (N_5807,N_5291,N_5196);
and U5808 (N_5808,N_5486,N_5594);
xor U5809 (N_5809,N_5349,N_5157);
and U5810 (N_5810,N_5309,N_5066);
nor U5811 (N_5811,N_5002,N_5563);
xnor U5812 (N_5812,N_5240,N_5468);
nand U5813 (N_5813,N_5246,N_5086);
or U5814 (N_5814,N_5624,N_5522);
nand U5815 (N_5815,N_5470,N_5218);
nor U5816 (N_5816,N_5104,N_5258);
or U5817 (N_5817,N_5030,N_5160);
nand U5818 (N_5818,N_5547,N_5078);
nor U5819 (N_5819,N_5008,N_5471);
and U5820 (N_5820,N_5462,N_5198);
nor U5821 (N_5821,N_5164,N_5447);
nand U5822 (N_5822,N_5418,N_5122);
nor U5823 (N_5823,N_5299,N_5607);
and U5824 (N_5824,N_5589,N_5277);
xnor U5825 (N_5825,N_5131,N_5288);
and U5826 (N_5826,N_5332,N_5099);
xor U5827 (N_5827,N_5102,N_5048);
and U5828 (N_5828,N_5289,N_5087);
and U5829 (N_5829,N_5050,N_5178);
and U5830 (N_5830,N_5305,N_5616);
and U5831 (N_5831,N_5121,N_5567);
and U5832 (N_5832,N_5432,N_5512);
or U5833 (N_5833,N_5421,N_5593);
or U5834 (N_5834,N_5106,N_5427);
nor U5835 (N_5835,N_5298,N_5303);
or U5836 (N_5836,N_5384,N_5194);
nor U5837 (N_5837,N_5105,N_5166);
xor U5838 (N_5838,N_5367,N_5433);
and U5839 (N_5839,N_5156,N_5612);
xor U5840 (N_5840,N_5362,N_5148);
xnor U5841 (N_5841,N_5431,N_5185);
nand U5842 (N_5842,N_5398,N_5333);
nor U5843 (N_5843,N_5076,N_5032);
nor U5844 (N_5844,N_5065,N_5311);
and U5845 (N_5845,N_5124,N_5040);
xnor U5846 (N_5846,N_5265,N_5422);
and U5847 (N_5847,N_5037,N_5226);
xor U5848 (N_5848,N_5534,N_5075);
or U5849 (N_5849,N_5508,N_5239);
nand U5850 (N_5850,N_5278,N_5588);
and U5851 (N_5851,N_5255,N_5357);
and U5852 (N_5852,N_5529,N_5403);
and U5853 (N_5853,N_5130,N_5416);
nor U5854 (N_5854,N_5016,N_5306);
and U5855 (N_5855,N_5517,N_5028);
nand U5856 (N_5856,N_5058,N_5402);
or U5857 (N_5857,N_5317,N_5460);
and U5858 (N_5858,N_5559,N_5377);
or U5859 (N_5859,N_5064,N_5227);
nand U5860 (N_5860,N_5263,N_5430);
nor U5861 (N_5861,N_5465,N_5496);
nand U5862 (N_5862,N_5051,N_5113);
xor U5863 (N_5863,N_5256,N_5621);
xor U5864 (N_5864,N_5223,N_5061);
nand U5865 (N_5865,N_5212,N_5006);
nor U5866 (N_5866,N_5466,N_5420);
nand U5867 (N_5867,N_5343,N_5428);
xnor U5868 (N_5868,N_5335,N_5519);
and U5869 (N_5869,N_5457,N_5415);
nand U5870 (N_5870,N_5033,N_5141);
nor U5871 (N_5871,N_5183,N_5276);
xor U5872 (N_5872,N_5211,N_5300);
nand U5873 (N_5873,N_5244,N_5315);
nor U5874 (N_5874,N_5406,N_5014);
nor U5875 (N_5875,N_5571,N_5237);
nor U5876 (N_5876,N_5555,N_5248);
or U5877 (N_5877,N_5039,N_5474);
xnor U5878 (N_5878,N_5390,N_5609);
and U5879 (N_5879,N_5424,N_5020);
or U5880 (N_5880,N_5376,N_5081);
nand U5881 (N_5881,N_5155,N_5210);
and U5882 (N_5882,N_5320,N_5270);
nor U5883 (N_5883,N_5205,N_5260);
or U5884 (N_5884,N_5331,N_5132);
nand U5885 (N_5885,N_5484,N_5613);
xnor U5886 (N_5886,N_5238,N_5110);
and U5887 (N_5887,N_5458,N_5525);
nand U5888 (N_5888,N_5219,N_5245);
xor U5889 (N_5889,N_5022,N_5580);
xnor U5890 (N_5890,N_5229,N_5049);
xor U5891 (N_5891,N_5201,N_5395);
xor U5892 (N_5892,N_5436,N_5583);
xnor U5893 (N_5893,N_5247,N_5179);
xor U5894 (N_5894,N_5497,N_5176);
nand U5895 (N_5895,N_5410,N_5538);
nand U5896 (N_5896,N_5063,N_5035);
xnor U5897 (N_5897,N_5445,N_5096);
nand U5898 (N_5898,N_5503,N_5531);
or U5899 (N_5899,N_5242,N_5142);
or U5900 (N_5900,N_5241,N_5281);
or U5901 (N_5901,N_5145,N_5464);
nand U5902 (N_5902,N_5207,N_5230);
xnor U5903 (N_5903,N_5378,N_5562);
nor U5904 (N_5904,N_5477,N_5574);
nor U5905 (N_5905,N_5366,N_5158);
and U5906 (N_5906,N_5001,N_5373);
nand U5907 (N_5907,N_5118,N_5172);
nand U5908 (N_5908,N_5026,N_5187);
or U5909 (N_5909,N_5284,N_5047);
or U5910 (N_5910,N_5019,N_5127);
or U5911 (N_5911,N_5015,N_5197);
or U5912 (N_5912,N_5556,N_5437);
nand U5913 (N_5913,N_5275,N_5339);
nand U5914 (N_5914,N_5318,N_5575);
nor U5915 (N_5915,N_5077,N_5379);
or U5916 (N_5916,N_5000,N_5091);
nor U5917 (N_5917,N_5055,N_5443);
xor U5918 (N_5918,N_5330,N_5412);
nor U5919 (N_5919,N_5361,N_5596);
and U5920 (N_5920,N_5011,N_5287);
or U5921 (N_5921,N_5487,N_5383);
nand U5922 (N_5922,N_5174,N_5043);
nand U5923 (N_5923,N_5493,N_5073);
or U5924 (N_5924,N_5004,N_5552);
xnor U5925 (N_5925,N_5009,N_5440);
and U5926 (N_5926,N_5071,N_5089);
and U5927 (N_5927,N_5133,N_5203);
xnor U5928 (N_5928,N_5511,N_5038);
nor U5929 (N_5929,N_5013,N_5249);
xnor U5930 (N_5930,N_5186,N_5070);
xnor U5931 (N_5931,N_5498,N_5224);
and U5932 (N_5932,N_5523,N_5351);
or U5933 (N_5933,N_5492,N_5250);
nor U5934 (N_5934,N_5389,N_5382);
nand U5935 (N_5935,N_5393,N_5438);
xnor U5936 (N_5936,N_5451,N_5391);
and U5937 (N_5937,N_5417,N_5274);
xor U5938 (N_5938,N_5354,N_5432);
nor U5939 (N_5939,N_5517,N_5081);
and U5940 (N_5940,N_5137,N_5517);
nand U5941 (N_5941,N_5104,N_5337);
xnor U5942 (N_5942,N_5200,N_5619);
nand U5943 (N_5943,N_5437,N_5236);
nand U5944 (N_5944,N_5358,N_5251);
and U5945 (N_5945,N_5037,N_5449);
nor U5946 (N_5946,N_5523,N_5299);
nor U5947 (N_5947,N_5018,N_5553);
xnor U5948 (N_5948,N_5116,N_5278);
and U5949 (N_5949,N_5138,N_5133);
or U5950 (N_5950,N_5346,N_5607);
or U5951 (N_5951,N_5542,N_5029);
xnor U5952 (N_5952,N_5168,N_5502);
and U5953 (N_5953,N_5186,N_5398);
nor U5954 (N_5954,N_5446,N_5344);
nand U5955 (N_5955,N_5390,N_5350);
xnor U5956 (N_5956,N_5554,N_5433);
xor U5957 (N_5957,N_5214,N_5113);
nor U5958 (N_5958,N_5475,N_5558);
nor U5959 (N_5959,N_5322,N_5534);
xor U5960 (N_5960,N_5597,N_5549);
or U5961 (N_5961,N_5456,N_5063);
and U5962 (N_5962,N_5532,N_5340);
and U5963 (N_5963,N_5238,N_5105);
nand U5964 (N_5964,N_5575,N_5302);
and U5965 (N_5965,N_5384,N_5569);
or U5966 (N_5966,N_5254,N_5365);
or U5967 (N_5967,N_5503,N_5190);
and U5968 (N_5968,N_5527,N_5548);
nand U5969 (N_5969,N_5092,N_5330);
and U5970 (N_5970,N_5344,N_5620);
or U5971 (N_5971,N_5228,N_5071);
nor U5972 (N_5972,N_5307,N_5581);
or U5973 (N_5973,N_5186,N_5620);
or U5974 (N_5974,N_5328,N_5537);
xnor U5975 (N_5975,N_5266,N_5490);
or U5976 (N_5976,N_5586,N_5480);
and U5977 (N_5977,N_5241,N_5454);
and U5978 (N_5978,N_5517,N_5543);
and U5979 (N_5979,N_5291,N_5376);
nand U5980 (N_5980,N_5245,N_5077);
nand U5981 (N_5981,N_5170,N_5367);
xor U5982 (N_5982,N_5496,N_5029);
xnor U5983 (N_5983,N_5537,N_5035);
nor U5984 (N_5984,N_5268,N_5231);
or U5985 (N_5985,N_5267,N_5247);
and U5986 (N_5986,N_5463,N_5033);
nand U5987 (N_5987,N_5223,N_5203);
nor U5988 (N_5988,N_5317,N_5381);
nor U5989 (N_5989,N_5471,N_5284);
and U5990 (N_5990,N_5106,N_5277);
or U5991 (N_5991,N_5230,N_5458);
or U5992 (N_5992,N_5020,N_5006);
nand U5993 (N_5993,N_5521,N_5166);
xnor U5994 (N_5994,N_5353,N_5543);
nor U5995 (N_5995,N_5239,N_5163);
nand U5996 (N_5996,N_5035,N_5365);
and U5997 (N_5997,N_5561,N_5180);
or U5998 (N_5998,N_5290,N_5140);
nor U5999 (N_5999,N_5175,N_5106);
xnor U6000 (N_6000,N_5469,N_5130);
and U6001 (N_6001,N_5462,N_5334);
and U6002 (N_6002,N_5607,N_5485);
and U6003 (N_6003,N_5080,N_5049);
and U6004 (N_6004,N_5622,N_5020);
xnor U6005 (N_6005,N_5328,N_5312);
and U6006 (N_6006,N_5130,N_5397);
nor U6007 (N_6007,N_5524,N_5376);
or U6008 (N_6008,N_5193,N_5488);
nand U6009 (N_6009,N_5327,N_5312);
xor U6010 (N_6010,N_5528,N_5262);
nand U6011 (N_6011,N_5450,N_5176);
nor U6012 (N_6012,N_5302,N_5438);
xor U6013 (N_6013,N_5125,N_5035);
nor U6014 (N_6014,N_5113,N_5610);
and U6015 (N_6015,N_5600,N_5341);
nor U6016 (N_6016,N_5391,N_5437);
or U6017 (N_6017,N_5056,N_5299);
and U6018 (N_6018,N_5161,N_5307);
or U6019 (N_6019,N_5457,N_5483);
or U6020 (N_6020,N_5583,N_5090);
xnor U6021 (N_6021,N_5192,N_5478);
and U6022 (N_6022,N_5331,N_5481);
xor U6023 (N_6023,N_5510,N_5198);
nand U6024 (N_6024,N_5614,N_5288);
or U6025 (N_6025,N_5228,N_5622);
or U6026 (N_6026,N_5566,N_5401);
and U6027 (N_6027,N_5294,N_5144);
nor U6028 (N_6028,N_5142,N_5154);
nand U6029 (N_6029,N_5011,N_5089);
or U6030 (N_6030,N_5545,N_5109);
or U6031 (N_6031,N_5617,N_5241);
nor U6032 (N_6032,N_5139,N_5245);
and U6033 (N_6033,N_5392,N_5486);
or U6034 (N_6034,N_5454,N_5387);
nand U6035 (N_6035,N_5353,N_5532);
nor U6036 (N_6036,N_5383,N_5386);
or U6037 (N_6037,N_5042,N_5157);
or U6038 (N_6038,N_5194,N_5162);
or U6039 (N_6039,N_5061,N_5482);
or U6040 (N_6040,N_5559,N_5438);
and U6041 (N_6041,N_5258,N_5419);
nand U6042 (N_6042,N_5024,N_5132);
and U6043 (N_6043,N_5344,N_5445);
xor U6044 (N_6044,N_5245,N_5426);
and U6045 (N_6045,N_5442,N_5054);
xor U6046 (N_6046,N_5017,N_5298);
nor U6047 (N_6047,N_5501,N_5545);
and U6048 (N_6048,N_5373,N_5507);
nand U6049 (N_6049,N_5577,N_5550);
nor U6050 (N_6050,N_5368,N_5366);
nand U6051 (N_6051,N_5292,N_5612);
or U6052 (N_6052,N_5125,N_5586);
nor U6053 (N_6053,N_5552,N_5357);
or U6054 (N_6054,N_5257,N_5588);
nand U6055 (N_6055,N_5609,N_5505);
xor U6056 (N_6056,N_5396,N_5315);
nand U6057 (N_6057,N_5543,N_5176);
and U6058 (N_6058,N_5073,N_5110);
nor U6059 (N_6059,N_5380,N_5157);
nor U6060 (N_6060,N_5066,N_5486);
or U6061 (N_6061,N_5138,N_5115);
or U6062 (N_6062,N_5576,N_5563);
nand U6063 (N_6063,N_5543,N_5384);
and U6064 (N_6064,N_5178,N_5129);
nand U6065 (N_6065,N_5404,N_5061);
nand U6066 (N_6066,N_5474,N_5011);
or U6067 (N_6067,N_5133,N_5108);
xnor U6068 (N_6068,N_5377,N_5267);
and U6069 (N_6069,N_5328,N_5258);
xor U6070 (N_6070,N_5117,N_5522);
xnor U6071 (N_6071,N_5407,N_5428);
or U6072 (N_6072,N_5305,N_5286);
and U6073 (N_6073,N_5390,N_5460);
xnor U6074 (N_6074,N_5064,N_5152);
nor U6075 (N_6075,N_5472,N_5292);
nor U6076 (N_6076,N_5066,N_5412);
nand U6077 (N_6077,N_5232,N_5565);
xor U6078 (N_6078,N_5461,N_5040);
nor U6079 (N_6079,N_5587,N_5130);
xnor U6080 (N_6080,N_5260,N_5614);
nor U6081 (N_6081,N_5302,N_5131);
and U6082 (N_6082,N_5357,N_5123);
nand U6083 (N_6083,N_5444,N_5279);
or U6084 (N_6084,N_5532,N_5309);
or U6085 (N_6085,N_5493,N_5023);
xnor U6086 (N_6086,N_5304,N_5033);
nor U6087 (N_6087,N_5276,N_5040);
nor U6088 (N_6088,N_5375,N_5544);
and U6089 (N_6089,N_5603,N_5397);
or U6090 (N_6090,N_5540,N_5099);
nand U6091 (N_6091,N_5233,N_5432);
xnor U6092 (N_6092,N_5362,N_5116);
xnor U6093 (N_6093,N_5144,N_5040);
nand U6094 (N_6094,N_5438,N_5498);
nor U6095 (N_6095,N_5467,N_5136);
or U6096 (N_6096,N_5255,N_5429);
xor U6097 (N_6097,N_5508,N_5546);
nor U6098 (N_6098,N_5056,N_5554);
xor U6099 (N_6099,N_5132,N_5389);
nor U6100 (N_6100,N_5312,N_5322);
or U6101 (N_6101,N_5566,N_5107);
xor U6102 (N_6102,N_5501,N_5097);
nand U6103 (N_6103,N_5041,N_5315);
xor U6104 (N_6104,N_5599,N_5349);
or U6105 (N_6105,N_5313,N_5174);
and U6106 (N_6106,N_5191,N_5489);
xor U6107 (N_6107,N_5412,N_5099);
xnor U6108 (N_6108,N_5372,N_5487);
or U6109 (N_6109,N_5148,N_5616);
and U6110 (N_6110,N_5246,N_5010);
nor U6111 (N_6111,N_5115,N_5582);
nand U6112 (N_6112,N_5452,N_5247);
or U6113 (N_6113,N_5023,N_5546);
or U6114 (N_6114,N_5194,N_5555);
nor U6115 (N_6115,N_5263,N_5379);
xor U6116 (N_6116,N_5417,N_5431);
or U6117 (N_6117,N_5482,N_5412);
and U6118 (N_6118,N_5290,N_5506);
and U6119 (N_6119,N_5544,N_5097);
xor U6120 (N_6120,N_5445,N_5622);
nor U6121 (N_6121,N_5227,N_5164);
or U6122 (N_6122,N_5051,N_5451);
nand U6123 (N_6123,N_5425,N_5087);
or U6124 (N_6124,N_5379,N_5254);
nand U6125 (N_6125,N_5374,N_5600);
and U6126 (N_6126,N_5410,N_5522);
xor U6127 (N_6127,N_5457,N_5207);
and U6128 (N_6128,N_5310,N_5079);
nand U6129 (N_6129,N_5515,N_5455);
nor U6130 (N_6130,N_5434,N_5381);
xnor U6131 (N_6131,N_5491,N_5550);
or U6132 (N_6132,N_5108,N_5442);
nand U6133 (N_6133,N_5463,N_5515);
nor U6134 (N_6134,N_5250,N_5384);
and U6135 (N_6135,N_5458,N_5357);
and U6136 (N_6136,N_5308,N_5466);
xnor U6137 (N_6137,N_5147,N_5514);
or U6138 (N_6138,N_5470,N_5105);
nand U6139 (N_6139,N_5029,N_5463);
or U6140 (N_6140,N_5157,N_5622);
and U6141 (N_6141,N_5164,N_5593);
and U6142 (N_6142,N_5463,N_5606);
xor U6143 (N_6143,N_5269,N_5050);
nand U6144 (N_6144,N_5262,N_5258);
or U6145 (N_6145,N_5521,N_5165);
nand U6146 (N_6146,N_5340,N_5269);
nand U6147 (N_6147,N_5400,N_5447);
xnor U6148 (N_6148,N_5291,N_5307);
nand U6149 (N_6149,N_5298,N_5175);
nor U6150 (N_6150,N_5263,N_5047);
or U6151 (N_6151,N_5048,N_5394);
xor U6152 (N_6152,N_5367,N_5012);
and U6153 (N_6153,N_5161,N_5600);
nor U6154 (N_6154,N_5421,N_5125);
nand U6155 (N_6155,N_5147,N_5398);
xnor U6156 (N_6156,N_5479,N_5353);
nor U6157 (N_6157,N_5180,N_5087);
xor U6158 (N_6158,N_5413,N_5130);
or U6159 (N_6159,N_5519,N_5255);
xor U6160 (N_6160,N_5576,N_5200);
xnor U6161 (N_6161,N_5201,N_5062);
nand U6162 (N_6162,N_5451,N_5574);
and U6163 (N_6163,N_5392,N_5197);
xnor U6164 (N_6164,N_5039,N_5169);
nand U6165 (N_6165,N_5014,N_5352);
nor U6166 (N_6166,N_5458,N_5352);
xor U6167 (N_6167,N_5037,N_5281);
xnor U6168 (N_6168,N_5418,N_5591);
and U6169 (N_6169,N_5037,N_5218);
xor U6170 (N_6170,N_5191,N_5118);
xor U6171 (N_6171,N_5117,N_5357);
nand U6172 (N_6172,N_5620,N_5095);
or U6173 (N_6173,N_5308,N_5024);
xnor U6174 (N_6174,N_5218,N_5553);
and U6175 (N_6175,N_5566,N_5215);
or U6176 (N_6176,N_5205,N_5489);
or U6177 (N_6177,N_5234,N_5027);
nand U6178 (N_6178,N_5178,N_5213);
or U6179 (N_6179,N_5201,N_5210);
nand U6180 (N_6180,N_5345,N_5421);
and U6181 (N_6181,N_5200,N_5415);
and U6182 (N_6182,N_5413,N_5430);
or U6183 (N_6183,N_5325,N_5367);
or U6184 (N_6184,N_5539,N_5616);
nand U6185 (N_6185,N_5054,N_5597);
and U6186 (N_6186,N_5386,N_5384);
and U6187 (N_6187,N_5401,N_5205);
nor U6188 (N_6188,N_5560,N_5220);
xnor U6189 (N_6189,N_5122,N_5367);
or U6190 (N_6190,N_5162,N_5547);
nor U6191 (N_6191,N_5545,N_5237);
and U6192 (N_6192,N_5456,N_5605);
and U6193 (N_6193,N_5240,N_5038);
nand U6194 (N_6194,N_5348,N_5621);
and U6195 (N_6195,N_5081,N_5329);
and U6196 (N_6196,N_5375,N_5131);
nand U6197 (N_6197,N_5247,N_5113);
and U6198 (N_6198,N_5539,N_5208);
and U6199 (N_6199,N_5154,N_5562);
nand U6200 (N_6200,N_5011,N_5278);
nor U6201 (N_6201,N_5528,N_5228);
nor U6202 (N_6202,N_5580,N_5540);
and U6203 (N_6203,N_5223,N_5602);
and U6204 (N_6204,N_5269,N_5152);
or U6205 (N_6205,N_5622,N_5347);
or U6206 (N_6206,N_5559,N_5030);
and U6207 (N_6207,N_5610,N_5501);
nand U6208 (N_6208,N_5147,N_5309);
and U6209 (N_6209,N_5134,N_5138);
and U6210 (N_6210,N_5239,N_5411);
and U6211 (N_6211,N_5021,N_5403);
nand U6212 (N_6212,N_5341,N_5044);
nand U6213 (N_6213,N_5458,N_5346);
xor U6214 (N_6214,N_5317,N_5140);
xnor U6215 (N_6215,N_5473,N_5128);
nor U6216 (N_6216,N_5578,N_5381);
xnor U6217 (N_6217,N_5305,N_5031);
or U6218 (N_6218,N_5343,N_5454);
xor U6219 (N_6219,N_5503,N_5426);
nand U6220 (N_6220,N_5487,N_5417);
nor U6221 (N_6221,N_5476,N_5463);
xor U6222 (N_6222,N_5469,N_5254);
and U6223 (N_6223,N_5297,N_5014);
nand U6224 (N_6224,N_5224,N_5089);
or U6225 (N_6225,N_5044,N_5124);
nand U6226 (N_6226,N_5593,N_5452);
or U6227 (N_6227,N_5376,N_5252);
and U6228 (N_6228,N_5151,N_5139);
nor U6229 (N_6229,N_5184,N_5393);
nor U6230 (N_6230,N_5597,N_5554);
nor U6231 (N_6231,N_5355,N_5084);
nor U6232 (N_6232,N_5551,N_5468);
or U6233 (N_6233,N_5224,N_5321);
nor U6234 (N_6234,N_5565,N_5433);
or U6235 (N_6235,N_5034,N_5231);
nor U6236 (N_6236,N_5460,N_5222);
or U6237 (N_6237,N_5136,N_5261);
and U6238 (N_6238,N_5233,N_5098);
xor U6239 (N_6239,N_5243,N_5031);
xor U6240 (N_6240,N_5450,N_5148);
xnor U6241 (N_6241,N_5195,N_5113);
nor U6242 (N_6242,N_5303,N_5602);
nor U6243 (N_6243,N_5362,N_5347);
and U6244 (N_6244,N_5535,N_5615);
nor U6245 (N_6245,N_5032,N_5091);
nor U6246 (N_6246,N_5451,N_5020);
xor U6247 (N_6247,N_5508,N_5512);
nor U6248 (N_6248,N_5229,N_5382);
nand U6249 (N_6249,N_5153,N_5498);
xor U6250 (N_6250,N_6054,N_6061);
nor U6251 (N_6251,N_5698,N_6083);
nor U6252 (N_6252,N_5962,N_6130);
and U6253 (N_6253,N_6105,N_6027);
or U6254 (N_6254,N_5897,N_6089);
nand U6255 (N_6255,N_6087,N_5978);
xor U6256 (N_6256,N_6114,N_5695);
nor U6257 (N_6257,N_5968,N_5664);
or U6258 (N_6258,N_5999,N_6245);
nand U6259 (N_6259,N_5697,N_5668);
nor U6260 (N_6260,N_5754,N_6071);
nor U6261 (N_6261,N_6204,N_6188);
or U6262 (N_6262,N_5822,N_5790);
or U6263 (N_6263,N_5824,N_5844);
or U6264 (N_6264,N_5920,N_5975);
or U6265 (N_6265,N_5735,N_5864);
and U6266 (N_6266,N_6079,N_5817);
or U6267 (N_6267,N_6058,N_5915);
and U6268 (N_6268,N_5748,N_6214);
nand U6269 (N_6269,N_5659,N_5758);
nand U6270 (N_6270,N_6246,N_5686);
nand U6271 (N_6271,N_5926,N_6136);
nor U6272 (N_6272,N_6032,N_5843);
or U6273 (N_6273,N_5811,N_5728);
and U6274 (N_6274,N_5712,N_5996);
xnor U6275 (N_6275,N_5929,N_5831);
xnor U6276 (N_6276,N_5903,N_5910);
xor U6277 (N_6277,N_6034,N_6148);
and U6278 (N_6278,N_5655,N_5784);
nor U6279 (N_6279,N_5694,N_6218);
or U6280 (N_6280,N_5855,N_5781);
and U6281 (N_6281,N_5626,N_6103);
or U6282 (N_6282,N_5902,N_5932);
and U6283 (N_6283,N_5840,N_6059);
nand U6284 (N_6284,N_6025,N_6197);
nor U6285 (N_6285,N_5923,N_6176);
or U6286 (N_6286,N_6137,N_5858);
and U6287 (N_6287,N_5990,N_5636);
or U6288 (N_6288,N_5885,N_6039);
nand U6289 (N_6289,N_5802,N_6097);
and U6290 (N_6290,N_5800,N_6207);
and U6291 (N_6291,N_6019,N_6146);
or U6292 (N_6292,N_6240,N_5684);
and U6293 (N_6293,N_6026,N_6140);
and U6294 (N_6294,N_5647,N_6196);
xnor U6295 (N_6295,N_6002,N_6011);
and U6296 (N_6296,N_5988,N_5709);
nand U6297 (N_6297,N_6141,N_5770);
nand U6298 (N_6298,N_5820,N_5997);
xor U6299 (N_6299,N_5813,N_6219);
and U6300 (N_6300,N_5936,N_5736);
nand U6301 (N_6301,N_6050,N_5846);
and U6302 (N_6302,N_5702,N_6180);
xnor U6303 (N_6303,N_6093,N_5752);
or U6304 (N_6304,N_5699,N_6117);
or U6305 (N_6305,N_6175,N_6161);
or U6306 (N_6306,N_5856,N_5906);
xor U6307 (N_6307,N_5727,N_6088);
xnor U6308 (N_6308,N_5768,N_6139);
xnor U6309 (N_6309,N_5964,N_5927);
xor U6310 (N_6310,N_5871,N_6086);
nand U6311 (N_6311,N_6178,N_6100);
xnor U6312 (N_6312,N_5714,N_5872);
nand U6313 (N_6313,N_6211,N_5795);
and U6314 (N_6314,N_5774,N_6224);
and U6315 (N_6315,N_5653,N_6084);
or U6316 (N_6316,N_5630,N_6000);
xor U6317 (N_6317,N_6158,N_6151);
or U6318 (N_6318,N_5751,N_6183);
nand U6319 (N_6319,N_5646,N_6080);
or U6320 (N_6320,N_6051,N_6015);
and U6321 (N_6321,N_5961,N_6123);
nand U6322 (N_6322,N_5991,N_5656);
xor U6323 (N_6323,N_6138,N_5755);
nor U6324 (N_6324,N_6206,N_6202);
and U6325 (N_6325,N_6067,N_5738);
and U6326 (N_6326,N_6205,N_6220);
and U6327 (N_6327,N_5682,N_5966);
or U6328 (N_6328,N_5776,N_5842);
xnor U6329 (N_6329,N_5974,N_5950);
xor U6330 (N_6330,N_5853,N_5984);
or U6331 (N_6331,N_5805,N_6031);
nor U6332 (N_6332,N_5658,N_6213);
or U6333 (N_6333,N_5971,N_5868);
or U6334 (N_6334,N_5878,N_5866);
or U6335 (N_6335,N_6085,N_5625);
nor U6336 (N_6336,N_5716,N_5870);
or U6337 (N_6337,N_6028,N_5704);
xnor U6338 (N_6338,N_6073,N_6249);
and U6339 (N_6339,N_5983,N_6153);
nand U6340 (N_6340,N_5806,N_5976);
nand U6341 (N_6341,N_5772,N_5977);
or U6342 (N_6342,N_5663,N_5803);
or U6343 (N_6343,N_5881,N_5737);
and U6344 (N_6344,N_5725,N_5877);
or U6345 (N_6345,N_6185,N_5690);
xnor U6346 (N_6346,N_6234,N_5845);
nand U6347 (N_6347,N_5912,N_6150);
and U6348 (N_6348,N_6223,N_6056);
nor U6349 (N_6349,N_5786,N_6237);
nand U6350 (N_6350,N_5639,N_5821);
or U6351 (N_6351,N_5746,N_5979);
and U6352 (N_6352,N_5830,N_5633);
xnor U6353 (N_6353,N_6003,N_6216);
or U6354 (N_6354,N_5807,N_6167);
nand U6355 (N_6355,N_5718,N_5762);
and U6356 (N_6356,N_5838,N_5723);
nand U6357 (N_6357,N_6238,N_6242);
or U6358 (N_6358,N_5930,N_6109);
nor U6359 (N_6359,N_6008,N_5994);
and U6360 (N_6360,N_5722,N_5969);
nor U6361 (N_6361,N_5992,N_5917);
nand U6362 (N_6362,N_5940,N_5710);
nor U6363 (N_6363,N_6060,N_5960);
and U6364 (N_6364,N_5884,N_6235);
and U6365 (N_6365,N_5879,N_6181);
xnor U6366 (N_6366,N_6247,N_5671);
nand U6367 (N_6367,N_5804,N_6164);
or U6368 (N_6368,N_6037,N_6190);
nand U6369 (N_6369,N_5944,N_6023);
nor U6370 (N_6370,N_5891,N_6094);
or U6371 (N_6371,N_6052,N_5829);
nor U6372 (N_6372,N_6228,N_6095);
xnor U6373 (N_6373,N_5701,N_6182);
and U6374 (N_6374,N_5798,N_5933);
nor U6375 (N_6375,N_5757,N_5850);
nand U6376 (N_6376,N_5687,N_6106);
xor U6377 (N_6377,N_5836,N_5677);
and U6378 (N_6378,N_6009,N_6040);
nor U6379 (N_6379,N_6169,N_6159);
nor U6380 (N_6380,N_5995,N_6135);
or U6381 (N_6381,N_5854,N_6033);
and U6382 (N_6382,N_5678,N_5908);
nand U6383 (N_6383,N_6113,N_5819);
nor U6384 (N_6384,N_5681,N_6121);
or U6385 (N_6385,N_6074,N_5833);
and U6386 (N_6386,N_6045,N_5700);
xor U6387 (N_6387,N_5892,N_5660);
nand U6388 (N_6388,N_5711,N_5753);
or U6389 (N_6389,N_5794,N_5631);
nand U6390 (N_6390,N_5680,N_6192);
and U6391 (N_6391,N_5739,N_6070);
or U6392 (N_6392,N_6195,N_5652);
and U6393 (N_6393,N_5672,N_5889);
xor U6394 (N_6394,N_5981,N_6006);
or U6395 (N_6395,N_5869,N_5775);
and U6396 (N_6396,N_5779,N_5987);
xnor U6397 (N_6397,N_6022,N_5764);
and U6398 (N_6398,N_6166,N_6124);
xnor U6399 (N_6399,N_6145,N_5632);
xor U6400 (N_6400,N_5967,N_6203);
or U6401 (N_6401,N_6001,N_5789);
xnor U6402 (N_6402,N_6239,N_5665);
xnor U6403 (N_6403,N_5922,N_5715);
nand U6404 (N_6404,N_5860,N_5675);
nand U6405 (N_6405,N_5769,N_5899);
nor U6406 (N_6406,N_6099,N_6063);
and U6407 (N_6407,N_6013,N_5792);
or U6408 (N_6408,N_6171,N_6017);
xor U6409 (N_6409,N_5828,N_6077);
and U6410 (N_6410,N_5857,N_5980);
nand U6411 (N_6411,N_6082,N_5852);
or U6412 (N_6412,N_6173,N_5662);
or U6413 (N_6413,N_5919,N_6018);
xor U6414 (N_6414,N_5706,N_5849);
xor U6415 (N_6415,N_5673,N_5777);
and U6416 (N_6416,N_5628,N_6016);
and U6417 (N_6417,N_5904,N_6090);
nor U6418 (N_6418,N_5670,N_5782);
xor U6419 (N_6419,N_5900,N_6029);
or U6420 (N_6420,N_5669,N_6098);
xnor U6421 (N_6421,N_5947,N_5679);
nand U6422 (N_6422,N_5880,N_5685);
or U6423 (N_6423,N_6221,N_6069);
nand U6424 (N_6424,N_5676,N_6142);
or U6425 (N_6425,N_6122,N_5839);
or U6426 (N_6426,N_5771,N_5861);
nor U6427 (N_6427,N_5890,N_5651);
nand U6428 (N_6428,N_5657,N_5693);
nor U6429 (N_6429,N_5692,N_5705);
xor U6430 (N_6430,N_5924,N_6119);
and U6431 (N_6431,N_6076,N_5907);
nor U6432 (N_6432,N_5888,N_6186);
nor U6433 (N_6433,N_6134,N_5661);
nand U6434 (N_6434,N_6064,N_5973);
nand U6435 (N_6435,N_6007,N_5951);
xnor U6436 (N_6436,N_5859,N_5745);
nand U6437 (N_6437,N_5882,N_6155);
nor U6438 (N_6438,N_6162,N_6004);
and U6439 (N_6439,N_5948,N_6232);
nand U6440 (N_6440,N_5749,N_5939);
or U6441 (N_6441,N_6057,N_6200);
nor U6442 (N_6442,N_5946,N_5949);
xor U6443 (N_6443,N_5742,N_5744);
or U6444 (N_6444,N_6030,N_5816);
xor U6445 (N_6445,N_6231,N_5740);
xor U6446 (N_6446,N_5637,N_5865);
or U6447 (N_6447,N_5873,N_6147);
or U6448 (N_6448,N_6233,N_5766);
nand U6449 (N_6449,N_6035,N_6209);
nor U6450 (N_6450,N_6133,N_6110);
xor U6451 (N_6451,N_6160,N_5894);
or U6452 (N_6452,N_5887,N_6091);
nand U6453 (N_6453,N_5837,N_5759);
xor U6454 (N_6454,N_6226,N_6217);
nor U6455 (N_6455,N_5761,N_5952);
and U6456 (N_6456,N_5788,N_5953);
or U6457 (N_6457,N_6210,N_5954);
nand U6458 (N_6458,N_5627,N_5874);
xnor U6459 (N_6459,N_5724,N_6152);
nand U6460 (N_6460,N_6174,N_5862);
xnor U6461 (N_6461,N_5925,N_5750);
and U6462 (N_6462,N_6081,N_5696);
nand U6463 (N_6463,N_5832,N_5921);
nand U6464 (N_6464,N_6230,N_5703);
nor U6465 (N_6465,N_5941,N_5935);
and U6466 (N_6466,N_5972,N_6005);
nand U6467 (N_6467,N_5898,N_6041);
xnor U6468 (N_6468,N_6143,N_5913);
nor U6469 (N_6469,N_6179,N_5689);
and U6470 (N_6470,N_5928,N_5767);
and U6471 (N_6471,N_5886,N_6154);
and U6472 (N_6472,N_6012,N_5825);
nor U6473 (N_6473,N_6131,N_6248);
nand U6474 (N_6474,N_6184,N_6048);
nor U6475 (N_6475,N_6062,N_5911);
and U6476 (N_6476,N_6236,N_6065);
xor U6477 (N_6477,N_6047,N_6132);
nand U6478 (N_6478,N_5895,N_5733);
or U6479 (N_6479,N_6043,N_5629);
xnor U6480 (N_6480,N_5916,N_6053);
xor U6481 (N_6481,N_6038,N_5787);
xnor U6482 (N_6482,N_6193,N_5645);
nor U6483 (N_6483,N_5810,N_6189);
and U6484 (N_6484,N_5943,N_6010);
and U6485 (N_6485,N_6156,N_6092);
xnor U6486 (N_6486,N_5959,N_6116);
or U6487 (N_6487,N_6170,N_5638);
and U6488 (N_6488,N_6227,N_5955);
nor U6489 (N_6489,N_6096,N_5641);
or U6490 (N_6490,N_6144,N_6111);
nand U6491 (N_6491,N_5848,N_5778);
xnor U6492 (N_6492,N_5893,N_5783);
nand U6493 (N_6493,N_5741,N_5998);
nor U6494 (N_6494,N_5814,N_5938);
or U6495 (N_6495,N_6177,N_5815);
xnor U6496 (N_6496,N_6014,N_5876);
xor U6497 (N_6497,N_5986,N_6036);
nor U6498 (N_6498,N_5847,N_5914);
nand U6499 (N_6499,N_6066,N_6120);
xnor U6500 (N_6500,N_6229,N_5937);
nand U6501 (N_6501,N_5834,N_5763);
nor U6502 (N_6502,N_5640,N_5765);
and U6503 (N_6503,N_6172,N_5957);
nand U6504 (N_6504,N_6075,N_6102);
nand U6505 (N_6505,N_5809,N_6187);
and U6506 (N_6506,N_6055,N_5791);
or U6507 (N_6507,N_5643,N_5958);
xnor U6508 (N_6508,N_6222,N_5732);
and U6509 (N_6509,N_6024,N_6042);
or U6510 (N_6510,N_5883,N_5797);
or U6511 (N_6511,N_5896,N_5993);
nand U6512 (N_6512,N_5965,N_5729);
and U6513 (N_6513,N_5867,N_6128);
nor U6514 (N_6514,N_6021,N_5708);
xnor U6515 (N_6515,N_5707,N_5863);
nor U6516 (N_6516,N_6129,N_5747);
xor U6517 (N_6517,N_5818,N_6157);
nor U6518 (N_6518,N_6241,N_6127);
and U6519 (N_6519,N_5982,N_5667);
or U6520 (N_6520,N_6072,N_5942);
nor U6521 (N_6521,N_5808,N_5760);
nor U6522 (N_6522,N_6149,N_5796);
xnor U6523 (N_6523,N_6168,N_6244);
xor U6524 (N_6524,N_5719,N_5666);
nor U6525 (N_6525,N_6201,N_5726);
or U6526 (N_6526,N_5931,N_5720);
and U6527 (N_6527,N_5835,N_5827);
nor U6528 (N_6528,N_6078,N_6049);
nand U6529 (N_6529,N_5730,N_5721);
and U6530 (N_6530,N_5743,N_5909);
nand U6531 (N_6531,N_5851,N_6046);
and U6532 (N_6532,N_6212,N_6101);
nor U6533 (N_6533,N_6194,N_5654);
xnor U6534 (N_6534,N_5945,N_5793);
nor U6535 (N_6535,N_6020,N_6199);
and U6536 (N_6536,N_6115,N_5970);
or U6537 (N_6537,N_5780,N_6104);
or U6538 (N_6538,N_5634,N_5649);
or U6539 (N_6539,N_6165,N_5688);
xor U6540 (N_6540,N_5713,N_6243);
nor U6541 (N_6541,N_5918,N_5734);
or U6542 (N_6542,N_6208,N_5650);
nor U6543 (N_6543,N_5731,N_5989);
nand U6544 (N_6544,N_5901,N_5773);
nand U6545 (N_6545,N_6126,N_5756);
or U6546 (N_6546,N_6068,N_6044);
xor U6547 (N_6547,N_5635,N_5956);
and U6548 (N_6548,N_5905,N_5717);
and U6549 (N_6549,N_5785,N_5799);
xor U6550 (N_6550,N_5934,N_5812);
and U6551 (N_6551,N_6163,N_5648);
nor U6552 (N_6552,N_5674,N_6118);
nand U6553 (N_6553,N_6198,N_6225);
nand U6554 (N_6554,N_5683,N_6125);
and U6555 (N_6555,N_5985,N_5963);
nor U6556 (N_6556,N_6215,N_5691);
xor U6557 (N_6557,N_5642,N_6112);
and U6558 (N_6558,N_5644,N_5826);
nor U6559 (N_6559,N_5841,N_5823);
or U6560 (N_6560,N_6108,N_6191);
and U6561 (N_6561,N_6107,N_5801);
or U6562 (N_6562,N_5875,N_5719);
and U6563 (N_6563,N_5998,N_5985);
xor U6564 (N_6564,N_5932,N_6133);
nand U6565 (N_6565,N_5683,N_5839);
nand U6566 (N_6566,N_5966,N_5865);
nand U6567 (N_6567,N_5705,N_5979);
or U6568 (N_6568,N_5639,N_6082);
nor U6569 (N_6569,N_5907,N_6020);
nand U6570 (N_6570,N_6132,N_6040);
or U6571 (N_6571,N_5831,N_5697);
or U6572 (N_6572,N_5826,N_6236);
nor U6573 (N_6573,N_5962,N_6053);
and U6574 (N_6574,N_6170,N_5717);
or U6575 (N_6575,N_5966,N_6148);
or U6576 (N_6576,N_5935,N_5677);
nand U6577 (N_6577,N_5912,N_5745);
xor U6578 (N_6578,N_5922,N_5863);
and U6579 (N_6579,N_6233,N_6218);
or U6580 (N_6580,N_6085,N_6094);
and U6581 (N_6581,N_5878,N_5988);
and U6582 (N_6582,N_5996,N_5784);
nand U6583 (N_6583,N_6076,N_6008);
or U6584 (N_6584,N_5960,N_5928);
nor U6585 (N_6585,N_6060,N_5983);
xor U6586 (N_6586,N_5876,N_6129);
and U6587 (N_6587,N_5672,N_5761);
nor U6588 (N_6588,N_6167,N_6062);
and U6589 (N_6589,N_5768,N_5749);
or U6590 (N_6590,N_5877,N_5985);
nor U6591 (N_6591,N_6122,N_5929);
nor U6592 (N_6592,N_5758,N_6156);
xor U6593 (N_6593,N_5953,N_5764);
or U6594 (N_6594,N_6180,N_5718);
xnor U6595 (N_6595,N_5859,N_6100);
nor U6596 (N_6596,N_6229,N_5850);
and U6597 (N_6597,N_6153,N_6038);
xor U6598 (N_6598,N_5761,N_6145);
nand U6599 (N_6599,N_5874,N_6061);
and U6600 (N_6600,N_5978,N_5825);
nor U6601 (N_6601,N_6035,N_5672);
xnor U6602 (N_6602,N_5923,N_5851);
nand U6603 (N_6603,N_6002,N_5751);
nor U6604 (N_6604,N_5900,N_5943);
xnor U6605 (N_6605,N_5920,N_5985);
nand U6606 (N_6606,N_5890,N_5805);
and U6607 (N_6607,N_6123,N_5994);
nor U6608 (N_6608,N_5770,N_5950);
nor U6609 (N_6609,N_6086,N_5918);
and U6610 (N_6610,N_5768,N_5991);
nand U6611 (N_6611,N_5694,N_5668);
nand U6612 (N_6612,N_5915,N_6217);
nand U6613 (N_6613,N_6185,N_6023);
xor U6614 (N_6614,N_5654,N_5655);
and U6615 (N_6615,N_5642,N_5726);
and U6616 (N_6616,N_6228,N_6015);
nand U6617 (N_6617,N_5725,N_6224);
nand U6618 (N_6618,N_6139,N_5649);
or U6619 (N_6619,N_5922,N_5793);
and U6620 (N_6620,N_5959,N_5823);
nor U6621 (N_6621,N_6141,N_6143);
or U6622 (N_6622,N_6159,N_6187);
nand U6623 (N_6623,N_6186,N_5720);
or U6624 (N_6624,N_6043,N_5789);
nand U6625 (N_6625,N_6129,N_5826);
or U6626 (N_6626,N_6084,N_5974);
xnor U6627 (N_6627,N_5874,N_5743);
xor U6628 (N_6628,N_5761,N_6159);
or U6629 (N_6629,N_5896,N_5639);
nor U6630 (N_6630,N_5630,N_5680);
and U6631 (N_6631,N_5866,N_6029);
nor U6632 (N_6632,N_5916,N_6016);
or U6633 (N_6633,N_5829,N_6151);
or U6634 (N_6634,N_5817,N_6058);
nor U6635 (N_6635,N_5647,N_5735);
nand U6636 (N_6636,N_5882,N_6097);
nand U6637 (N_6637,N_5669,N_6153);
and U6638 (N_6638,N_6046,N_5912);
or U6639 (N_6639,N_6186,N_6175);
nor U6640 (N_6640,N_5949,N_6047);
nand U6641 (N_6641,N_6175,N_6177);
nand U6642 (N_6642,N_5854,N_5988);
or U6643 (N_6643,N_6019,N_6026);
xnor U6644 (N_6644,N_6092,N_5776);
and U6645 (N_6645,N_6053,N_5907);
or U6646 (N_6646,N_6114,N_5731);
and U6647 (N_6647,N_5822,N_5630);
nand U6648 (N_6648,N_5823,N_5790);
or U6649 (N_6649,N_5651,N_6185);
or U6650 (N_6650,N_6109,N_5836);
nor U6651 (N_6651,N_6028,N_6073);
nor U6652 (N_6652,N_5911,N_5652);
and U6653 (N_6653,N_6181,N_5626);
and U6654 (N_6654,N_6197,N_6194);
nor U6655 (N_6655,N_6168,N_6235);
nand U6656 (N_6656,N_5797,N_6023);
xor U6657 (N_6657,N_5901,N_6130);
and U6658 (N_6658,N_5930,N_5687);
nor U6659 (N_6659,N_5770,N_5867);
nand U6660 (N_6660,N_5949,N_6092);
or U6661 (N_6661,N_5900,N_5690);
xor U6662 (N_6662,N_6074,N_5952);
and U6663 (N_6663,N_6073,N_6185);
or U6664 (N_6664,N_6135,N_6237);
nand U6665 (N_6665,N_6017,N_5631);
and U6666 (N_6666,N_5882,N_5798);
nor U6667 (N_6667,N_6111,N_5957);
xor U6668 (N_6668,N_5626,N_5844);
nor U6669 (N_6669,N_6137,N_5983);
and U6670 (N_6670,N_5883,N_5682);
xor U6671 (N_6671,N_5881,N_5997);
xor U6672 (N_6672,N_5968,N_6165);
or U6673 (N_6673,N_5704,N_6175);
or U6674 (N_6674,N_5875,N_5746);
nand U6675 (N_6675,N_5947,N_6144);
or U6676 (N_6676,N_6067,N_5741);
and U6677 (N_6677,N_6017,N_5735);
xor U6678 (N_6678,N_5680,N_6015);
or U6679 (N_6679,N_6160,N_6034);
nor U6680 (N_6680,N_5668,N_5797);
nand U6681 (N_6681,N_5709,N_6013);
nand U6682 (N_6682,N_6128,N_5859);
xnor U6683 (N_6683,N_6232,N_5868);
and U6684 (N_6684,N_5900,N_6173);
nand U6685 (N_6685,N_6248,N_5748);
and U6686 (N_6686,N_5957,N_5811);
nand U6687 (N_6687,N_5870,N_5888);
nor U6688 (N_6688,N_5861,N_6047);
or U6689 (N_6689,N_6161,N_5783);
and U6690 (N_6690,N_5864,N_6144);
or U6691 (N_6691,N_5661,N_6086);
and U6692 (N_6692,N_5941,N_6047);
or U6693 (N_6693,N_5728,N_5826);
or U6694 (N_6694,N_6214,N_5989);
nor U6695 (N_6695,N_5972,N_5968);
nand U6696 (N_6696,N_6148,N_6139);
xor U6697 (N_6697,N_5642,N_5638);
and U6698 (N_6698,N_6082,N_5741);
or U6699 (N_6699,N_5925,N_5683);
nor U6700 (N_6700,N_6240,N_5676);
nand U6701 (N_6701,N_5790,N_5872);
nand U6702 (N_6702,N_5843,N_6120);
xor U6703 (N_6703,N_6062,N_5869);
or U6704 (N_6704,N_5802,N_6046);
and U6705 (N_6705,N_6102,N_5767);
nand U6706 (N_6706,N_5948,N_5676);
nand U6707 (N_6707,N_6050,N_5704);
xnor U6708 (N_6708,N_5839,N_5898);
or U6709 (N_6709,N_6185,N_5843);
or U6710 (N_6710,N_5688,N_5980);
and U6711 (N_6711,N_6012,N_6053);
nand U6712 (N_6712,N_6236,N_5686);
nand U6713 (N_6713,N_5907,N_5644);
nand U6714 (N_6714,N_5772,N_5629);
nand U6715 (N_6715,N_5847,N_6107);
nor U6716 (N_6716,N_5773,N_6135);
nand U6717 (N_6717,N_5971,N_5715);
nand U6718 (N_6718,N_6027,N_5895);
nand U6719 (N_6719,N_5851,N_5833);
nand U6720 (N_6720,N_6227,N_6139);
nand U6721 (N_6721,N_6236,N_5631);
nand U6722 (N_6722,N_5841,N_5921);
nor U6723 (N_6723,N_6123,N_5908);
and U6724 (N_6724,N_5861,N_6118);
nand U6725 (N_6725,N_6104,N_6060);
or U6726 (N_6726,N_5917,N_5851);
or U6727 (N_6727,N_5798,N_6145);
nand U6728 (N_6728,N_5843,N_5713);
nand U6729 (N_6729,N_6098,N_6156);
and U6730 (N_6730,N_6179,N_5761);
or U6731 (N_6731,N_5871,N_5650);
nor U6732 (N_6732,N_5832,N_6212);
and U6733 (N_6733,N_5948,N_5849);
xnor U6734 (N_6734,N_5721,N_5772);
and U6735 (N_6735,N_5956,N_5985);
and U6736 (N_6736,N_6220,N_6025);
and U6737 (N_6737,N_5916,N_5812);
and U6738 (N_6738,N_6178,N_5815);
or U6739 (N_6739,N_6079,N_6096);
nand U6740 (N_6740,N_6197,N_5804);
or U6741 (N_6741,N_6202,N_6217);
nor U6742 (N_6742,N_5858,N_6241);
nor U6743 (N_6743,N_6053,N_5771);
and U6744 (N_6744,N_5851,N_5752);
xnor U6745 (N_6745,N_5845,N_5781);
nor U6746 (N_6746,N_6188,N_6093);
nor U6747 (N_6747,N_6189,N_5875);
and U6748 (N_6748,N_5700,N_6228);
nand U6749 (N_6749,N_5763,N_6105);
and U6750 (N_6750,N_5943,N_5737);
and U6751 (N_6751,N_5681,N_5863);
or U6752 (N_6752,N_5662,N_6029);
nand U6753 (N_6753,N_6051,N_5997);
nand U6754 (N_6754,N_5804,N_6027);
nand U6755 (N_6755,N_6116,N_5653);
and U6756 (N_6756,N_5818,N_5690);
and U6757 (N_6757,N_6244,N_5691);
nor U6758 (N_6758,N_6044,N_6118);
xor U6759 (N_6759,N_6238,N_6228);
and U6760 (N_6760,N_5737,N_5850);
nor U6761 (N_6761,N_5747,N_5798);
or U6762 (N_6762,N_5817,N_6155);
nand U6763 (N_6763,N_5790,N_5776);
nand U6764 (N_6764,N_6224,N_5994);
nor U6765 (N_6765,N_6197,N_5859);
and U6766 (N_6766,N_6017,N_6226);
nor U6767 (N_6767,N_6033,N_6195);
nor U6768 (N_6768,N_6076,N_5838);
nand U6769 (N_6769,N_5901,N_5842);
xnor U6770 (N_6770,N_6187,N_5891);
nor U6771 (N_6771,N_5719,N_5911);
xnor U6772 (N_6772,N_5793,N_6007);
or U6773 (N_6773,N_6138,N_6157);
xnor U6774 (N_6774,N_6157,N_6120);
xnor U6775 (N_6775,N_5833,N_5938);
nand U6776 (N_6776,N_5866,N_5673);
nand U6777 (N_6777,N_5893,N_6016);
and U6778 (N_6778,N_5926,N_5956);
nand U6779 (N_6779,N_6171,N_6002);
nand U6780 (N_6780,N_5909,N_5843);
xnor U6781 (N_6781,N_5786,N_5756);
nor U6782 (N_6782,N_5952,N_6097);
nor U6783 (N_6783,N_5995,N_6105);
nand U6784 (N_6784,N_6097,N_5850);
nand U6785 (N_6785,N_5762,N_6189);
xor U6786 (N_6786,N_6090,N_5847);
or U6787 (N_6787,N_6031,N_6084);
xor U6788 (N_6788,N_6080,N_6239);
and U6789 (N_6789,N_6167,N_5632);
and U6790 (N_6790,N_6229,N_5810);
and U6791 (N_6791,N_5977,N_5837);
nor U6792 (N_6792,N_5850,N_6207);
or U6793 (N_6793,N_6245,N_6136);
and U6794 (N_6794,N_5979,N_5736);
nand U6795 (N_6795,N_6166,N_5666);
nor U6796 (N_6796,N_5743,N_5706);
and U6797 (N_6797,N_5926,N_5679);
nor U6798 (N_6798,N_5830,N_5900);
nand U6799 (N_6799,N_5761,N_6066);
nand U6800 (N_6800,N_5654,N_5987);
nand U6801 (N_6801,N_6041,N_5631);
nor U6802 (N_6802,N_5757,N_5862);
nand U6803 (N_6803,N_5847,N_5965);
xor U6804 (N_6804,N_6132,N_6212);
nand U6805 (N_6805,N_6099,N_5842);
nor U6806 (N_6806,N_5786,N_5681);
nor U6807 (N_6807,N_5779,N_5937);
nand U6808 (N_6808,N_5851,N_5672);
and U6809 (N_6809,N_6199,N_6130);
nand U6810 (N_6810,N_6154,N_6087);
nand U6811 (N_6811,N_5988,N_5892);
and U6812 (N_6812,N_5762,N_5737);
or U6813 (N_6813,N_5789,N_6241);
nor U6814 (N_6814,N_5629,N_6182);
nor U6815 (N_6815,N_6052,N_6072);
and U6816 (N_6816,N_6175,N_5783);
nand U6817 (N_6817,N_6019,N_5651);
xor U6818 (N_6818,N_6072,N_6086);
nor U6819 (N_6819,N_5660,N_5807);
xor U6820 (N_6820,N_6013,N_5997);
or U6821 (N_6821,N_5782,N_6098);
nor U6822 (N_6822,N_5881,N_6118);
xor U6823 (N_6823,N_5678,N_5869);
xnor U6824 (N_6824,N_6119,N_5907);
nor U6825 (N_6825,N_5721,N_6178);
or U6826 (N_6826,N_6111,N_5986);
nor U6827 (N_6827,N_6053,N_5805);
nor U6828 (N_6828,N_5730,N_6072);
nand U6829 (N_6829,N_5665,N_6143);
xnor U6830 (N_6830,N_5701,N_6131);
or U6831 (N_6831,N_6065,N_6061);
nand U6832 (N_6832,N_5887,N_6224);
and U6833 (N_6833,N_6121,N_5664);
and U6834 (N_6834,N_5649,N_5936);
xor U6835 (N_6835,N_6089,N_5849);
and U6836 (N_6836,N_5964,N_5893);
nor U6837 (N_6837,N_5861,N_5735);
nor U6838 (N_6838,N_6223,N_5683);
nor U6839 (N_6839,N_6219,N_5990);
nand U6840 (N_6840,N_6108,N_5773);
nor U6841 (N_6841,N_6115,N_5910);
or U6842 (N_6842,N_6075,N_6019);
nand U6843 (N_6843,N_5780,N_5753);
nor U6844 (N_6844,N_6244,N_5855);
or U6845 (N_6845,N_6238,N_5842);
xnor U6846 (N_6846,N_6141,N_6196);
nor U6847 (N_6847,N_5812,N_6138);
xor U6848 (N_6848,N_5823,N_6173);
xor U6849 (N_6849,N_5962,N_5842);
nor U6850 (N_6850,N_6008,N_6023);
and U6851 (N_6851,N_5931,N_5805);
xor U6852 (N_6852,N_5909,N_6100);
nand U6853 (N_6853,N_5670,N_5880);
xor U6854 (N_6854,N_5896,N_5750);
and U6855 (N_6855,N_6232,N_6028);
or U6856 (N_6856,N_6173,N_5637);
or U6857 (N_6857,N_5681,N_5924);
nand U6858 (N_6858,N_6226,N_5727);
nand U6859 (N_6859,N_6051,N_5985);
or U6860 (N_6860,N_6023,N_5886);
xor U6861 (N_6861,N_5669,N_5699);
xor U6862 (N_6862,N_5924,N_6061);
nand U6863 (N_6863,N_5950,N_6102);
or U6864 (N_6864,N_5833,N_6035);
nand U6865 (N_6865,N_6243,N_5769);
and U6866 (N_6866,N_5761,N_5919);
or U6867 (N_6867,N_5669,N_6022);
xor U6868 (N_6868,N_6098,N_5865);
xor U6869 (N_6869,N_5719,N_6028);
or U6870 (N_6870,N_5951,N_5692);
and U6871 (N_6871,N_5642,N_5976);
nand U6872 (N_6872,N_5924,N_6199);
or U6873 (N_6873,N_6232,N_5924);
and U6874 (N_6874,N_5990,N_5773);
nor U6875 (N_6875,N_6604,N_6685);
and U6876 (N_6876,N_6674,N_6869);
and U6877 (N_6877,N_6323,N_6689);
nand U6878 (N_6878,N_6422,N_6738);
nor U6879 (N_6879,N_6602,N_6428);
nand U6880 (N_6880,N_6487,N_6719);
xnor U6881 (N_6881,N_6650,N_6541);
or U6882 (N_6882,N_6306,N_6308);
nand U6883 (N_6883,N_6739,N_6839);
nand U6884 (N_6884,N_6459,N_6601);
nor U6885 (N_6885,N_6744,N_6835);
nor U6886 (N_6886,N_6451,N_6591);
or U6887 (N_6887,N_6542,N_6646);
and U6888 (N_6888,N_6395,N_6412);
or U6889 (N_6889,N_6423,N_6379);
nand U6890 (N_6890,N_6778,N_6256);
and U6891 (N_6891,N_6587,N_6663);
xnor U6892 (N_6892,N_6455,N_6818);
xor U6893 (N_6893,N_6293,N_6571);
xnor U6894 (N_6894,N_6438,N_6552);
xnor U6895 (N_6895,N_6311,N_6425);
or U6896 (N_6896,N_6672,N_6509);
nand U6897 (N_6897,N_6496,N_6697);
nor U6898 (N_6898,N_6703,N_6456);
nand U6899 (N_6899,N_6613,N_6720);
and U6900 (N_6900,N_6777,N_6670);
xnor U6901 (N_6901,N_6305,N_6765);
and U6902 (N_6902,N_6819,N_6847);
xor U6903 (N_6903,N_6253,N_6516);
nor U6904 (N_6904,N_6784,N_6301);
or U6905 (N_6905,N_6734,N_6594);
xor U6906 (N_6906,N_6483,N_6763);
and U6907 (N_6907,N_6327,N_6649);
or U6908 (N_6908,N_6475,N_6748);
nand U6909 (N_6909,N_6299,N_6679);
and U6910 (N_6910,N_6733,N_6832);
xor U6911 (N_6911,N_6866,N_6749);
nand U6912 (N_6912,N_6429,N_6651);
nor U6913 (N_6913,N_6848,N_6314);
nand U6914 (N_6914,N_6279,N_6692);
xor U6915 (N_6915,N_6261,N_6268);
and U6916 (N_6916,N_6675,N_6368);
xnor U6917 (N_6917,N_6351,N_6399);
xor U6918 (N_6918,N_6406,N_6362);
nor U6919 (N_6919,N_6295,N_6736);
nor U6920 (N_6920,N_6329,N_6389);
xor U6921 (N_6921,N_6330,N_6392);
nand U6922 (N_6922,N_6870,N_6417);
and U6923 (N_6923,N_6440,N_6641);
nand U6924 (N_6924,N_6677,N_6501);
or U6925 (N_6925,N_6338,N_6654);
nand U6926 (N_6926,N_6278,N_6700);
or U6927 (N_6927,N_6787,N_6630);
or U6928 (N_6928,N_6762,N_6753);
and U6929 (N_6929,N_6502,N_6657);
xor U6930 (N_6930,N_6536,N_6662);
nand U6931 (N_6931,N_6504,N_6312);
xor U6932 (N_6932,N_6551,N_6806);
xor U6933 (N_6933,N_6569,N_6708);
xnor U6934 (N_6934,N_6384,N_6310);
xnor U6935 (N_6935,N_6729,N_6332);
nor U6936 (N_6936,N_6628,N_6537);
or U6937 (N_6937,N_6514,N_6726);
nand U6938 (N_6938,N_6798,N_6757);
xor U6939 (N_6939,N_6653,N_6617);
nor U6940 (N_6940,N_6859,N_6524);
xor U6941 (N_6941,N_6370,N_6860);
or U6942 (N_6942,N_6386,N_6359);
nor U6943 (N_6943,N_6627,N_6290);
or U6944 (N_6944,N_6764,N_6498);
and U6945 (N_6945,N_6326,N_6793);
nand U6946 (N_6946,N_6714,N_6358);
and U6947 (N_6947,N_6799,N_6631);
nor U6948 (N_6948,N_6446,N_6385);
xor U6949 (N_6949,N_6792,N_6579);
nor U6950 (N_6950,N_6336,N_6534);
nand U6951 (N_6951,N_6302,N_6797);
xor U6952 (N_6952,N_6411,N_6444);
and U6953 (N_6953,N_6255,N_6767);
nor U6954 (N_6954,N_6741,N_6852);
or U6955 (N_6955,N_6759,N_6668);
and U6956 (N_6956,N_6289,N_6269);
xor U6957 (N_6957,N_6790,N_6723);
xnor U6958 (N_6958,N_6560,N_6251);
xor U6959 (N_6959,N_6372,N_6466);
nor U6960 (N_6960,N_6825,N_6292);
and U6961 (N_6961,N_6666,N_6671);
xnor U6962 (N_6962,N_6600,N_6297);
or U6963 (N_6963,N_6315,N_6391);
and U6964 (N_6964,N_6805,N_6851);
or U6965 (N_6965,N_6575,N_6356);
xor U6966 (N_6966,N_6680,N_6783);
nand U6967 (N_6967,N_6846,N_6706);
xnor U6968 (N_6968,N_6343,N_6394);
xor U6969 (N_6969,N_6402,N_6661);
nand U6970 (N_6970,N_6383,N_6773);
nor U6971 (N_6971,N_6335,N_6333);
xor U6972 (N_6972,N_6469,N_6262);
xor U6973 (N_6973,N_6341,N_6340);
xnor U6974 (N_6974,N_6543,N_6450);
and U6975 (N_6975,N_6530,N_6861);
xnor U6976 (N_6976,N_6864,N_6441);
nor U6977 (N_6977,N_6453,N_6334);
or U6978 (N_6978,N_6296,N_6486);
or U6979 (N_6979,N_6622,N_6484);
nand U6980 (N_6980,N_6642,N_6510);
and U6981 (N_6981,N_6270,N_6461);
or U6982 (N_6982,N_6562,N_6271);
nand U6983 (N_6983,N_6698,N_6865);
or U6984 (N_6984,N_6563,N_6813);
or U6985 (N_6985,N_6694,N_6621);
nor U6986 (N_6986,N_6452,N_6521);
and U6987 (N_6987,N_6527,N_6645);
nor U6988 (N_6988,N_6837,N_6775);
nor U6989 (N_6989,N_6515,N_6303);
and U6990 (N_6990,N_6812,N_6388);
and U6991 (N_6991,N_6477,N_6490);
nor U6992 (N_6992,N_6842,N_6324);
nor U6993 (N_6993,N_6566,N_6488);
and U6994 (N_6994,N_6795,N_6285);
nor U6995 (N_6995,N_6442,N_6637);
nand U6996 (N_6996,N_6616,N_6274);
and U6997 (N_6997,N_6476,N_6618);
nor U6998 (N_6998,N_6347,N_6580);
or U6999 (N_6999,N_6766,N_6458);
nand U7000 (N_7000,N_6508,N_6478);
nor U7001 (N_7001,N_6593,N_6578);
nor U7002 (N_7002,N_6400,N_6381);
nand U7003 (N_7003,N_6321,N_6715);
or U7004 (N_7004,N_6531,N_6322);
or U7005 (N_7005,N_6361,N_6364);
and U7006 (N_7006,N_6871,N_6686);
and U7007 (N_7007,N_6320,N_6590);
nor U7008 (N_7008,N_6768,N_6644);
and U7009 (N_7009,N_6266,N_6307);
and U7010 (N_7010,N_6319,N_6448);
nor U7011 (N_7011,N_6711,N_6817);
nor U7012 (N_7012,N_6664,N_6667);
or U7013 (N_7013,N_6647,N_6827);
xnor U7014 (N_7014,N_6619,N_6868);
nand U7015 (N_7015,N_6522,N_6610);
xor U7016 (N_7016,N_6769,N_6529);
nor U7017 (N_7017,N_6577,N_6781);
and U7018 (N_7018,N_6855,N_6660);
nand U7019 (N_7019,N_6743,N_6615);
and U7020 (N_7020,N_6607,N_6526);
or U7021 (N_7021,N_6405,N_6665);
nand U7022 (N_7022,N_6695,N_6873);
xnor U7023 (N_7023,N_6779,N_6833);
or U7024 (N_7024,N_6756,N_6474);
nor U7025 (N_7025,N_6275,N_6598);
nor U7026 (N_7026,N_6432,N_6648);
or U7027 (N_7027,N_6583,N_6513);
and U7028 (N_7028,N_6313,N_6471);
nand U7029 (N_7029,N_6856,N_6449);
nand U7030 (N_7030,N_6809,N_6863);
nand U7031 (N_7031,N_6512,N_6457);
nor U7032 (N_7032,N_6853,N_6273);
nand U7033 (N_7033,N_6624,N_6393);
or U7034 (N_7034,N_6603,N_6655);
and U7035 (N_7035,N_6494,N_6345);
nand U7036 (N_7036,N_6377,N_6761);
nor U7037 (N_7037,N_6460,N_6731);
and U7038 (N_7038,N_6331,N_6802);
and U7039 (N_7039,N_6557,N_6640);
nand U7040 (N_7040,N_6408,N_6712);
and U7041 (N_7041,N_6633,N_6612);
and U7042 (N_7042,N_6831,N_6472);
or U7043 (N_7043,N_6673,N_6443);
or U7044 (N_7044,N_6467,N_6874);
and U7045 (N_7045,N_6844,N_6634);
xnor U7046 (N_7046,N_6782,N_6470);
nand U7047 (N_7047,N_6858,N_6599);
and U7048 (N_7048,N_6420,N_6317);
nor U7049 (N_7049,N_6823,N_6540);
xnor U7050 (N_7050,N_6367,N_6822);
and U7051 (N_7051,N_6403,N_6463);
or U7052 (N_7052,N_6482,N_6639);
and U7053 (N_7053,N_6742,N_6713);
nand U7054 (N_7054,N_6716,N_6427);
nand U7055 (N_7055,N_6804,N_6493);
and U7056 (N_7056,N_6691,N_6752);
nor U7057 (N_7057,N_6586,N_6505);
and U7058 (N_7058,N_6298,N_6725);
and U7059 (N_7059,N_6597,N_6786);
nand U7060 (N_7060,N_6533,N_6464);
or U7061 (N_7061,N_6506,N_6528);
xor U7062 (N_7062,N_6337,N_6605);
nand U7063 (N_7063,N_6280,N_6554);
xor U7064 (N_7064,N_6772,N_6789);
or U7065 (N_7065,N_6410,N_6572);
or U7066 (N_7066,N_6318,N_6730);
nand U7067 (N_7067,N_6485,N_6576);
nor U7068 (N_7068,N_6500,N_6264);
xnor U7069 (N_7069,N_6820,N_6770);
xor U7070 (N_7070,N_6588,N_6746);
xnor U7071 (N_7071,N_6265,N_6520);
or U7072 (N_7072,N_6658,N_6676);
xnor U7073 (N_7073,N_6561,N_6415);
nor U7074 (N_7074,N_6595,N_6371);
nor U7075 (N_7075,N_6433,N_6854);
nand U7076 (N_7076,N_6636,N_6532);
or U7077 (N_7077,N_6840,N_6499);
and U7078 (N_7078,N_6824,N_6788);
and U7079 (N_7079,N_6465,N_6652);
and U7080 (N_7080,N_6365,N_6325);
nand U7081 (N_7081,N_6544,N_6735);
and U7082 (N_7082,N_6404,N_6702);
nand U7083 (N_7083,N_6491,N_6407);
xnor U7084 (N_7084,N_6418,N_6750);
xnor U7085 (N_7085,N_6355,N_6416);
nand U7086 (N_7086,N_6304,N_6821);
nor U7087 (N_7087,N_6565,N_6751);
nor U7088 (N_7088,N_6814,N_6549);
or U7089 (N_7089,N_6387,N_6747);
xor U7090 (N_7090,N_6539,N_6838);
nor U7091 (N_7091,N_6369,N_6608);
or U7092 (N_7092,N_6807,N_6545);
nand U7093 (N_7093,N_6260,N_6431);
or U7094 (N_7094,N_6836,N_6643);
or U7095 (N_7095,N_6287,N_6737);
and U7096 (N_7096,N_6573,N_6845);
and U7097 (N_7097,N_6776,N_6468);
xor U7098 (N_7098,N_6473,N_6632);
and U7099 (N_7099,N_6678,N_6780);
or U7100 (N_7100,N_6254,N_6732);
nand U7101 (N_7101,N_6707,N_6867);
xnor U7102 (N_7102,N_6426,N_6360);
xnor U7103 (N_7103,N_6517,N_6830);
nand U7104 (N_7104,N_6559,N_6348);
and U7105 (N_7105,N_6462,N_6376);
and U7106 (N_7106,N_6291,N_6437);
nand U7107 (N_7107,N_6727,N_6259);
and U7108 (N_7108,N_6611,N_6589);
nand U7109 (N_7109,N_6519,N_6872);
or U7110 (N_7110,N_6635,N_6445);
nor U7111 (N_7111,N_6489,N_6669);
nor U7112 (N_7112,N_6585,N_6592);
xor U7113 (N_7113,N_6841,N_6277);
nor U7114 (N_7114,N_6396,N_6771);
or U7115 (N_7115,N_6681,N_6350);
or U7116 (N_7116,N_6758,N_6862);
nand U7117 (N_7117,N_6564,N_6284);
nor U7118 (N_7118,N_6553,N_6492);
nand U7119 (N_7119,N_6479,N_6346);
nand U7120 (N_7120,N_6606,N_6309);
and U7121 (N_7121,N_6850,N_6421);
nor U7122 (N_7122,N_6547,N_6693);
and U7123 (N_7123,N_6574,N_6558);
or U7124 (N_7124,N_6857,N_6826);
or U7125 (N_7125,N_6447,N_6811);
nand U7126 (N_7126,N_6829,N_6375);
xor U7127 (N_7127,N_6511,N_6688);
and U7128 (N_7128,N_6570,N_6555);
or U7129 (N_7129,N_6609,N_6282);
and U7130 (N_7130,N_6808,N_6436);
or U7131 (N_7131,N_6803,N_6556);
xor U7132 (N_7132,N_6283,N_6409);
or U7133 (N_7133,N_6728,N_6378);
or U7134 (N_7134,N_6354,N_6701);
or U7135 (N_7135,N_6363,N_6272);
nor U7136 (N_7136,N_6709,N_6755);
and U7137 (N_7137,N_6801,N_6791);
nand U7138 (N_7138,N_6849,N_6373);
and U7139 (N_7139,N_6276,N_6687);
nor U7140 (N_7140,N_6357,N_6286);
nor U7141 (N_7141,N_6816,N_6518);
or U7142 (N_7142,N_6722,N_6828);
nand U7143 (N_7143,N_6339,N_6414);
nand U7144 (N_7144,N_6745,N_6774);
and U7145 (N_7145,N_6374,N_6690);
xor U7146 (N_7146,N_6810,N_6550);
or U7147 (N_7147,N_6413,N_6740);
nand U7148 (N_7148,N_6538,N_6638);
nor U7149 (N_7149,N_6721,N_6581);
xor U7150 (N_7150,N_6481,N_6454);
nor U7151 (N_7151,N_6382,N_6380);
and U7152 (N_7152,N_6718,N_6258);
or U7153 (N_7153,N_6704,N_6439);
nor U7154 (N_7154,N_6684,N_6342);
nand U7155 (N_7155,N_6316,N_6656);
or U7156 (N_7156,N_6401,N_6435);
or U7157 (N_7157,N_6567,N_6397);
or U7158 (N_7158,N_6366,N_6705);
xor U7159 (N_7159,N_6710,N_6390);
nand U7160 (N_7160,N_6699,N_6250);
nand U7161 (N_7161,N_6503,N_6815);
nor U7162 (N_7162,N_6625,N_6683);
or U7163 (N_7163,N_6263,N_6344);
nor U7164 (N_7164,N_6614,N_6257);
and U7165 (N_7165,N_6252,N_6430);
and U7166 (N_7166,N_6328,N_6834);
and U7167 (N_7167,N_6620,N_6267);
nand U7168 (N_7168,N_6596,N_6582);
xor U7169 (N_7169,N_6760,N_6629);
nand U7170 (N_7170,N_6696,N_6523);
xor U7171 (N_7171,N_6419,N_6349);
xnor U7172 (N_7172,N_6495,N_6352);
xnor U7173 (N_7173,N_6300,N_6525);
and U7174 (N_7174,N_6353,N_6754);
and U7175 (N_7175,N_6546,N_6398);
nand U7176 (N_7176,N_6568,N_6507);
nor U7177 (N_7177,N_6480,N_6535);
nor U7178 (N_7178,N_6434,N_6659);
nand U7179 (N_7179,N_6424,N_6294);
nor U7180 (N_7180,N_6623,N_6843);
or U7181 (N_7181,N_6497,N_6796);
or U7182 (N_7182,N_6682,N_6281);
nand U7183 (N_7183,N_6288,N_6724);
nand U7184 (N_7184,N_6584,N_6794);
xnor U7185 (N_7185,N_6626,N_6548);
or U7186 (N_7186,N_6785,N_6717);
nor U7187 (N_7187,N_6800,N_6344);
nand U7188 (N_7188,N_6296,N_6573);
or U7189 (N_7189,N_6340,N_6674);
nor U7190 (N_7190,N_6376,N_6555);
xor U7191 (N_7191,N_6771,N_6307);
nor U7192 (N_7192,N_6572,N_6831);
or U7193 (N_7193,N_6296,N_6414);
xnor U7194 (N_7194,N_6547,N_6606);
xnor U7195 (N_7195,N_6757,N_6546);
and U7196 (N_7196,N_6565,N_6252);
nand U7197 (N_7197,N_6521,N_6475);
or U7198 (N_7198,N_6741,N_6670);
nand U7199 (N_7199,N_6265,N_6456);
or U7200 (N_7200,N_6709,N_6272);
nand U7201 (N_7201,N_6306,N_6771);
or U7202 (N_7202,N_6701,N_6398);
and U7203 (N_7203,N_6593,N_6307);
nor U7204 (N_7204,N_6792,N_6381);
or U7205 (N_7205,N_6731,N_6676);
and U7206 (N_7206,N_6853,N_6373);
and U7207 (N_7207,N_6584,N_6565);
nor U7208 (N_7208,N_6860,N_6794);
and U7209 (N_7209,N_6584,N_6649);
nand U7210 (N_7210,N_6725,N_6370);
and U7211 (N_7211,N_6782,N_6662);
and U7212 (N_7212,N_6829,N_6304);
nor U7213 (N_7213,N_6835,N_6753);
nand U7214 (N_7214,N_6252,N_6858);
and U7215 (N_7215,N_6631,N_6426);
and U7216 (N_7216,N_6849,N_6440);
or U7217 (N_7217,N_6375,N_6425);
xnor U7218 (N_7218,N_6777,N_6327);
nand U7219 (N_7219,N_6262,N_6659);
xor U7220 (N_7220,N_6580,N_6326);
nand U7221 (N_7221,N_6786,N_6747);
or U7222 (N_7222,N_6328,N_6865);
and U7223 (N_7223,N_6813,N_6312);
or U7224 (N_7224,N_6609,N_6588);
nor U7225 (N_7225,N_6260,N_6473);
nor U7226 (N_7226,N_6294,N_6604);
nand U7227 (N_7227,N_6849,N_6626);
nand U7228 (N_7228,N_6583,N_6475);
and U7229 (N_7229,N_6362,N_6730);
or U7230 (N_7230,N_6746,N_6690);
or U7231 (N_7231,N_6825,N_6603);
or U7232 (N_7232,N_6338,N_6312);
xnor U7233 (N_7233,N_6303,N_6583);
xor U7234 (N_7234,N_6794,N_6318);
or U7235 (N_7235,N_6741,N_6463);
and U7236 (N_7236,N_6862,N_6372);
or U7237 (N_7237,N_6712,N_6512);
nor U7238 (N_7238,N_6832,N_6508);
nor U7239 (N_7239,N_6824,N_6522);
or U7240 (N_7240,N_6460,N_6613);
nor U7241 (N_7241,N_6731,N_6843);
or U7242 (N_7242,N_6851,N_6773);
or U7243 (N_7243,N_6753,N_6442);
nand U7244 (N_7244,N_6687,N_6863);
and U7245 (N_7245,N_6303,N_6302);
and U7246 (N_7246,N_6812,N_6754);
nor U7247 (N_7247,N_6772,N_6584);
or U7248 (N_7248,N_6315,N_6850);
and U7249 (N_7249,N_6842,N_6854);
xnor U7250 (N_7250,N_6754,N_6707);
or U7251 (N_7251,N_6360,N_6825);
xor U7252 (N_7252,N_6739,N_6359);
and U7253 (N_7253,N_6793,N_6865);
nor U7254 (N_7254,N_6529,N_6728);
or U7255 (N_7255,N_6468,N_6689);
nor U7256 (N_7256,N_6556,N_6312);
nor U7257 (N_7257,N_6429,N_6502);
and U7258 (N_7258,N_6442,N_6298);
xor U7259 (N_7259,N_6565,N_6367);
nand U7260 (N_7260,N_6384,N_6677);
nor U7261 (N_7261,N_6779,N_6572);
nand U7262 (N_7262,N_6796,N_6272);
nor U7263 (N_7263,N_6427,N_6251);
nor U7264 (N_7264,N_6582,N_6708);
xor U7265 (N_7265,N_6366,N_6346);
xor U7266 (N_7266,N_6485,N_6815);
nand U7267 (N_7267,N_6410,N_6738);
or U7268 (N_7268,N_6762,N_6800);
xor U7269 (N_7269,N_6513,N_6463);
and U7270 (N_7270,N_6822,N_6398);
nor U7271 (N_7271,N_6754,N_6670);
and U7272 (N_7272,N_6640,N_6286);
nand U7273 (N_7273,N_6661,N_6657);
nor U7274 (N_7274,N_6283,N_6419);
xnor U7275 (N_7275,N_6695,N_6848);
and U7276 (N_7276,N_6652,N_6689);
and U7277 (N_7277,N_6437,N_6550);
nor U7278 (N_7278,N_6576,N_6782);
nor U7279 (N_7279,N_6620,N_6579);
nor U7280 (N_7280,N_6844,N_6261);
nor U7281 (N_7281,N_6669,N_6254);
or U7282 (N_7282,N_6272,N_6423);
nand U7283 (N_7283,N_6288,N_6664);
and U7284 (N_7284,N_6759,N_6715);
nor U7285 (N_7285,N_6750,N_6802);
or U7286 (N_7286,N_6450,N_6479);
or U7287 (N_7287,N_6358,N_6265);
and U7288 (N_7288,N_6721,N_6334);
xor U7289 (N_7289,N_6653,N_6804);
and U7290 (N_7290,N_6480,N_6449);
or U7291 (N_7291,N_6835,N_6599);
and U7292 (N_7292,N_6791,N_6699);
or U7293 (N_7293,N_6379,N_6598);
or U7294 (N_7294,N_6648,N_6354);
or U7295 (N_7295,N_6715,N_6741);
xnor U7296 (N_7296,N_6649,N_6401);
nor U7297 (N_7297,N_6666,N_6802);
or U7298 (N_7298,N_6856,N_6820);
nand U7299 (N_7299,N_6864,N_6313);
or U7300 (N_7300,N_6448,N_6691);
or U7301 (N_7301,N_6828,N_6530);
nor U7302 (N_7302,N_6341,N_6639);
nand U7303 (N_7303,N_6734,N_6874);
xnor U7304 (N_7304,N_6519,N_6306);
and U7305 (N_7305,N_6479,N_6639);
xnor U7306 (N_7306,N_6633,N_6464);
or U7307 (N_7307,N_6677,N_6330);
xor U7308 (N_7308,N_6712,N_6532);
nor U7309 (N_7309,N_6341,N_6806);
nor U7310 (N_7310,N_6799,N_6312);
and U7311 (N_7311,N_6765,N_6738);
nand U7312 (N_7312,N_6297,N_6455);
nor U7313 (N_7313,N_6828,N_6619);
and U7314 (N_7314,N_6767,N_6850);
nor U7315 (N_7315,N_6612,N_6826);
nand U7316 (N_7316,N_6304,N_6605);
nor U7317 (N_7317,N_6341,N_6609);
xor U7318 (N_7318,N_6753,N_6551);
or U7319 (N_7319,N_6745,N_6365);
nor U7320 (N_7320,N_6511,N_6502);
and U7321 (N_7321,N_6263,N_6814);
nand U7322 (N_7322,N_6561,N_6572);
xnor U7323 (N_7323,N_6486,N_6758);
nand U7324 (N_7324,N_6861,N_6649);
xnor U7325 (N_7325,N_6428,N_6269);
nor U7326 (N_7326,N_6690,N_6529);
nand U7327 (N_7327,N_6732,N_6376);
and U7328 (N_7328,N_6858,N_6767);
nor U7329 (N_7329,N_6310,N_6771);
nand U7330 (N_7330,N_6465,N_6532);
nor U7331 (N_7331,N_6500,N_6295);
and U7332 (N_7332,N_6691,N_6711);
nand U7333 (N_7333,N_6341,N_6389);
or U7334 (N_7334,N_6693,N_6528);
nor U7335 (N_7335,N_6537,N_6749);
xnor U7336 (N_7336,N_6664,N_6351);
or U7337 (N_7337,N_6588,N_6327);
nand U7338 (N_7338,N_6679,N_6765);
xnor U7339 (N_7339,N_6676,N_6865);
nand U7340 (N_7340,N_6286,N_6254);
xnor U7341 (N_7341,N_6471,N_6537);
xnor U7342 (N_7342,N_6566,N_6744);
and U7343 (N_7343,N_6416,N_6452);
and U7344 (N_7344,N_6667,N_6370);
nor U7345 (N_7345,N_6329,N_6821);
or U7346 (N_7346,N_6795,N_6461);
or U7347 (N_7347,N_6598,N_6609);
or U7348 (N_7348,N_6479,N_6478);
and U7349 (N_7349,N_6744,N_6840);
and U7350 (N_7350,N_6363,N_6747);
xor U7351 (N_7351,N_6253,N_6637);
nor U7352 (N_7352,N_6732,N_6796);
nor U7353 (N_7353,N_6581,N_6374);
nor U7354 (N_7354,N_6778,N_6847);
xor U7355 (N_7355,N_6747,N_6731);
nand U7356 (N_7356,N_6603,N_6796);
nand U7357 (N_7357,N_6826,N_6289);
or U7358 (N_7358,N_6871,N_6600);
or U7359 (N_7359,N_6723,N_6678);
or U7360 (N_7360,N_6329,N_6544);
and U7361 (N_7361,N_6417,N_6595);
xor U7362 (N_7362,N_6309,N_6266);
or U7363 (N_7363,N_6305,N_6320);
nor U7364 (N_7364,N_6297,N_6498);
and U7365 (N_7365,N_6291,N_6612);
xor U7366 (N_7366,N_6764,N_6633);
or U7367 (N_7367,N_6655,N_6722);
nand U7368 (N_7368,N_6355,N_6798);
nor U7369 (N_7369,N_6591,N_6280);
or U7370 (N_7370,N_6750,N_6495);
or U7371 (N_7371,N_6643,N_6795);
and U7372 (N_7372,N_6361,N_6629);
xor U7373 (N_7373,N_6572,N_6553);
and U7374 (N_7374,N_6355,N_6780);
xor U7375 (N_7375,N_6694,N_6803);
nand U7376 (N_7376,N_6531,N_6418);
nor U7377 (N_7377,N_6467,N_6464);
xnor U7378 (N_7378,N_6805,N_6842);
or U7379 (N_7379,N_6812,N_6330);
nor U7380 (N_7380,N_6367,N_6662);
nand U7381 (N_7381,N_6774,N_6574);
xor U7382 (N_7382,N_6461,N_6609);
nor U7383 (N_7383,N_6866,N_6325);
xor U7384 (N_7384,N_6403,N_6749);
nand U7385 (N_7385,N_6271,N_6860);
or U7386 (N_7386,N_6546,N_6802);
or U7387 (N_7387,N_6440,N_6721);
and U7388 (N_7388,N_6361,N_6429);
nor U7389 (N_7389,N_6412,N_6681);
xor U7390 (N_7390,N_6407,N_6822);
or U7391 (N_7391,N_6722,N_6378);
nand U7392 (N_7392,N_6489,N_6729);
xor U7393 (N_7393,N_6669,N_6495);
and U7394 (N_7394,N_6383,N_6724);
or U7395 (N_7395,N_6662,N_6351);
xor U7396 (N_7396,N_6873,N_6730);
nor U7397 (N_7397,N_6325,N_6702);
or U7398 (N_7398,N_6865,N_6419);
or U7399 (N_7399,N_6789,N_6547);
nand U7400 (N_7400,N_6366,N_6645);
or U7401 (N_7401,N_6438,N_6439);
xnor U7402 (N_7402,N_6821,N_6396);
or U7403 (N_7403,N_6739,N_6770);
nand U7404 (N_7404,N_6678,N_6659);
nor U7405 (N_7405,N_6434,N_6874);
nor U7406 (N_7406,N_6775,N_6650);
xnor U7407 (N_7407,N_6286,N_6477);
nand U7408 (N_7408,N_6342,N_6357);
or U7409 (N_7409,N_6282,N_6617);
and U7410 (N_7410,N_6656,N_6768);
xor U7411 (N_7411,N_6422,N_6595);
nand U7412 (N_7412,N_6328,N_6689);
xnor U7413 (N_7413,N_6608,N_6853);
nor U7414 (N_7414,N_6410,N_6440);
and U7415 (N_7415,N_6534,N_6430);
xnor U7416 (N_7416,N_6550,N_6293);
or U7417 (N_7417,N_6403,N_6801);
nand U7418 (N_7418,N_6370,N_6523);
xor U7419 (N_7419,N_6684,N_6490);
nand U7420 (N_7420,N_6360,N_6570);
nand U7421 (N_7421,N_6436,N_6833);
nand U7422 (N_7422,N_6515,N_6725);
xnor U7423 (N_7423,N_6435,N_6597);
and U7424 (N_7424,N_6451,N_6335);
and U7425 (N_7425,N_6437,N_6341);
and U7426 (N_7426,N_6452,N_6664);
nor U7427 (N_7427,N_6850,N_6748);
and U7428 (N_7428,N_6334,N_6788);
nor U7429 (N_7429,N_6782,N_6699);
and U7430 (N_7430,N_6263,N_6856);
or U7431 (N_7431,N_6350,N_6299);
nand U7432 (N_7432,N_6834,N_6271);
and U7433 (N_7433,N_6479,N_6574);
and U7434 (N_7434,N_6315,N_6742);
xnor U7435 (N_7435,N_6761,N_6448);
and U7436 (N_7436,N_6625,N_6796);
nor U7437 (N_7437,N_6545,N_6721);
xnor U7438 (N_7438,N_6614,N_6719);
or U7439 (N_7439,N_6476,N_6367);
and U7440 (N_7440,N_6451,N_6480);
nand U7441 (N_7441,N_6696,N_6615);
and U7442 (N_7442,N_6408,N_6648);
xor U7443 (N_7443,N_6370,N_6382);
and U7444 (N_7444,N_6868,N_6252);
and U7445 (N_7445,N_6843,N_6692);
and U7446 (N_7446,N_6273,N_6365);
and U7447 (N_7447,N_6841,N_6325);
xnor U7448 (N_7448,N_6851,N_6668);
and U7449 (N_7449,N_6499,N_6443);
and U7450 (N_7450,N_6825,N_6774);
or U7451 (N_7451,N_6825,N_6406);
nand U7452 (N_7452,N_6638,N_6569);
nand U7453 (N_7453,N_6685,N_6536);
nand U7454 (N_7454,N_6542,N_6664);
nand U7455 (N_7455,N_6530,N_6642);
or U7456 (N_7456,N_6331,N_6656);
or U7457 (N_7457,N_6286,N_6708);
nor U7458 (N_7458,N_6678,N_6342);
nor U7459 (N_7459,N_6551,N_6853);
and U7460 (N_7460,N_6416,N_6284);
or U7461 (N_7461,N_6750,N_6573);
and U7462 (N_7462,N_6466,N_6264);
nor U7463 (N_7463,N_6347,N_6495);
nand U7464 (N_7464,N_6758,N_6613);
xor U7465 (N_7465,N_6831,N_6287);
nand U7466 (N_7466,N_6257,N_6766);
and U7467 (N_7467,N_6748,N_6791);
or U7468 (N_7468,N_6739,N_6829);
xor U7469 (N_7469,N_6440,N_6445);
or U7470 (N_7470,N_6304,N_6723);
nor U7471 (N_7471,N_6273,N_6432);
nor U7472 (N_7472,N_6476,N_6699);
nor U7473 (N_7473,N_6698,N_6365);
xnor U7474 (N_7474,N_6560,N_6253);
or U7475 (N_7475,N_6644,N_6259);
nand U7476 (N_7476,N_6853,N_6317);
and U7477 (N_7477,N_6825,N_6442);
xor U7478 (N_7478,N_6604,N_6562);
and U7479 (N_7479,N_6557,N_6298);
nand U7480 (N_7480,N_6305,N_6270);
nor U7481 (N_7481,N_6820,N_6302);
or U7482 (N_7482,N_6791,N_6592);
nor U7483 (N_7483,N_6430,N_6431);
or U7484 (N_7484,N_6335,N_6310);
or U7485 (N_7485,N_6755,N_6846);
or U7486 (N_7486,N_6447,N_6355);
nor U7487 (N_7487,N_6336,N_6762);
nor U7488 (N_7488,N_6762,N_6369);
and U7489 (N_7489,N_6439,N_6804);
nor U7490 (N_7490,N_6709,N_6558);
xor U7491 (N_7491,N_6396,N_6660);
xnor U7492 (N_7492,N_6650,N_6451);
nor U7493 (N_7493,N_6854,N_6558);
or U7494 (N_7494,N_6723,N_6552);
xor U7495 (N_7495,N_6801,N_6376);
and U7496 (N_7496,N_6268,N_6646);
xnor U7497 (N_7497,N_6613,N_6297);
or U7498 (N_7498,N_6575,N_6306);
or U7499 (N_7499,N_6616,N_6303);
xor U7500 (N_7500,N_7476,N_7436);
nor U7501 (N_7501,N_7194,N_7428);
nand U7502 (N_7502,N_7251,N_6906);
and U7503 (N_7503,N_6997,N_7368);
nand U7504 (N_7504,N_7367,N_6977);
or U7505 (N_7505,N_7112,N_7475);
and U7506 (N_7506,N_7373,N_7406);
and U7507 (N_7507,N_7175,N_7489);
xor U7508 (N_7508,N_7087,N_6975);
nor U7509 (N_7509,N_7197,N_6953);
nand U7510 (N_7510,N_6955,N_7347);
nand U7511 (N_7511,N_6973,N_7437);
and U7512 (N_7512,N_7139,N_6959);
and U7513 (N_7513,N_7479,N_6923);
nand U7514 (N_7514,N_7072,N_7138);
nor U7515 (N_7515,N_7375,N_7046);
nor U7516 (N_7516,N_7008,N_6907);
and U7517 (N_7517,N_6887,N_7136);
and U7518 (N_7518,N_7103,N_7441);
and U7519 (N_7519,N_6946,N_7385);
xnor U7520 (N_7520,N_7022,N_7192);
nand U7521 (N_7521,N_7255,N_6929);
nor U7522 (N_7522,N_7092,N_7277);
and U7523 (N_7523,N_7419,N_7259);
and U7524 (N_7524,N_7080,N_6879);
and U7525 (N_7525,N_7315,N_6875);
nand U7526 (N_7526,N_7451,N_7405);
nand U7527 (N_7527,N_7497,N_6981);
or U7528 (N_7528,N_7356,N_7300);
or U7529 (N_7529,N_7210,N_7317);
nand U7530 (N_7530,N_6942,N_7253);
and U7531 (N_7531,N_6976,N_6993);
nor U7532 (N_7532,N_7389,N_7477);
nand U7533 (N_7533,N_7301,N_7323);
xnor U7534 (N_7534,N_7453,N_7361);
and U7535 (N_7535,N_7307,N_7382);
and U7536 (N_7536,N_7393,N_7180);
nor U7537 (N_7537,N_7126,N_7042);
or U7538 (N_7538,N_7474,N_6990);
nand U7539 (N_7539,N_7450,N_7073);
or U7540 (N_7540,N_7338,N_7294);
nand U7541 (N_7541,N_7156,N_7454);
xor U7542 (N_7542,N_6908,N_7293);
nor U7543 (N_7543,N_7067,N_7026);
nand U7544 (N_7544,N_7006,N_6893);
or U7545 (N_7545,N_7131,N_7214);
and U7546 (N_7546,N_7309,N_7151);
nand U7547 (N_7547,N_7040,N_7161);
or U7548 (N_7548,N_7423,N_7190);
and U7549 (N_7549,N_7005,N_7117);
and U7550 (N_7550,N_7314,N_7155);
nand U7551 (N_7551,N_6918,N_7220);
nor U7552 (N_7552,N_7238,N_6986);
nor U7553 (N_7553,N_7229,N_7047);
or U7554 (N_7554,N_7207,N_7485);
or U7555 (N_7555,N_6922,N_7234);
nor U7556 (N_7556,N_7014,N_7213);
or U7557 (N_7557,N_7366,N_6913);
xnor U7558 (N_7558,N_7057,N_7304);
nand U7559 (N_7559,N_7009,N_6916);
xnor U7560 (N_7560,N_7459,N_7212);
nor U7561 (N_7561,N_7209,N_6969);
nand U7562 (N_7562,N_7033,N_7106);
nand U7563 (N_7563,N_7358,N_7204);
or U7564 (N_7564,N_7110,N_7283);
xor U7565 (N_7565,N_7312,N_7100);
or U7566 (N_7566,N_7374,N_7426);
nor U7567 (N_7567,N_7364,N_6994);
nor U7568 (N_7568,N_6896,N_7061);
nor U7569 (N_7569,N_7240,N_7381);
nor U7570 (N_7570,N_6950,N_6898);
nand U7571 (N_7571,N_7333,N_7051);
or U7572 (N_7572,N_7226,N_7482);
or U7573 (N_7573,N_7000,N_6979);
nand U7574 (N_7574,N_6967,N_7020);
nor U7575 (N_7575,N_6971,N_7111);
or U7576 (N_7576,N_7411,N_7181);
nor U7577 (N_7577,N_7402,N_7044);
xnor U7578 (N_7578,N_7230,N_7410);
xnor U7579 (N_7579,N_6938,N_6933);
and U7580 (N_7580,N_7062,N_7035);
nor U7581 (N_7581,N_6897,N_7342);
nand U7582 (N_7582,N_7254,N_7025);
or U7583 (N_7583,N_7457,N_7266);
xor U7584 (N_7584,N_7037,N_7143);
nand U7585 (N_7585,N_7086,N_7289);
nand U7586 (N_7586,N_7055,N_7007);
nand U7587 (N_7587,N_7414,N_7354);
xnor U7588 (N_7588,N_6949,N_7372);
or U7589 (N_7589,N_7228,N_6941);
or U7590 (N_7590,N_7049,N_7052);
xnor U7591 (N_7591,N_7455,N_6883);
nand U7592 (N_7592,N_7119,N_7202);
and U7593 (N_7593,N_7132,N_7446);
or U7594 (N_7594,N_7195,N_7286);
nor U7595 (N_7595,N_7463,N_7442);
nand U7596 (N_7596,N_6876,N_6945);
nor U7597 (N_7597,N_7282,N_7396);
xor U7598 (N_7598,N_7427,N_7438);
or U7599 (N_7599,N_7129,N_7499);
xor U7600 (N_7600,N_7248,N_7233);
nand U7601 (N_7601,N_7348,N_7247);
and U7602 (N_7602,N_7326,N_6937);
nor U7603 (N_7603,N_7335,N_7150);
nand U7604 (N_7604,N_7352,N_7193);
or U7605 (N_7605,N_6978,N_7429);
nor U7606 (N_7606,N_7425,N_7386);
nor U7607 (N_7607,N_7440,N_7256);
nor U7608 (N_7608,N_7388,N_7153);
xnor U7609 (N_7609,N_6983,N_6935);
xnor U7610 (N_7610,N_7239,N_7071);
nand U7611 (N_7611,N_6928,N_7257);
nor U7612 (N_7612,N_7174,N_7187);
nand U7613 (N_7613,N_7223,N_7343);
nand U7614 (N_7614,N_7029,N_7468);
or U7615 (N_7615,N_7308,N_7324);
nor U7616 (N_7616,N_7310,N_7465);
nor U7617 (N_7617,N_7268,N_7083);
nor U7618 (N_7618,N_7134,N_7345);
xor U7619 (N_7619,N_7169,N_7043);
or U7620 (N_7620,N_7376,N_7113);
xor U7621 (N_7621,N_7391,N_7404);
or U7622 (N_7622,N_7299,N_7095);
nor U7623 (N_7623,N_7152,N_7462);
nand U7624 (N_7624,N_7217,N_7305);
xnor U7625 (N_7625,N_6882,N_7068);
nand U7626 (N_7626,N_7246,N_7449);
or U7627 (N_7627,N_6980,N_7091);
xor U7628 (N_7628,N_7004,N_6904);
nor U7629 (N_7629,N_6903,N_7178);
nor U7630 (N_7630,N_6999,N_7144);
nand U7631 (N_7631,N_7048,N_7179);
nand U7632 (N_7632,N_7215,N_7149);
nand U7633 (N_7633,N_7355,N_7176);
or U7634 (N_7634,N_7291,N_7464);
nand U7635 (N_7635,N_6934,N_7168);
or U7636 (N_7636,N_7206,N_7019);
or U7637 (N_7637,N_7002,N_6886);
or U7638 (N_7638,N_7408,N_7433);
nand U7639 (N_7639,N_7265,N_7350);
xor U7640 (N_7640,N_7261,N_7056);
and U7641 (N_7641,N_6960,N_7218);
nor U7642 (N_7642,N_7023,N_7216);
or U7643 (N_7643,N_7357,N_6914);
nand U7644 (N_7644,N_7330,N_7456);
xor U7645 (N_7645,N_7390,N_7447);
and U7646 (N_7646,N_7377,N_7297);
nor U7647 (N_7647,N_7295,N_7413);
xnor U7648 (N_7648,N_7221,N_7045);
nand U7649 (N_7649,N_7311,N_7146);
nor U7650 (N_7650,N_7141,N_7339);
or U7651 (N_7651,N_7400,N_7109);
or U7652 (N_7652,N_7344,N_7362);
nand U7653 (N_7653,N_7183,N_7398);
nor U7654 (N_7654,N_7182,N_7365);
and U7655 (N_7655,N_7205,N_7084);
and U7656 (N_7656,N_7010,N_7270);
xnor U7657 (N_7657,N_7066,N_7353);
nand U7658 (N_7658,N_7001,N_7125);
and U7659 (N_7659,N_6889,N_7290);
xor U7660 (N_7660,N_6926,N_7371);
and U7661 (N_7661,N_7079,N_7082);
nor U7662 (N_7662,N_6905,N_7363);
nand U7663 (N_7663,N_7196,N_6998);
nand U7664 (N_7664,N_6884,N_7321);
or U7665 (N_7665,N_7191,N_7279);
or U7666 (N_7666,N_7050,N_7164);
nor U7667 (N_7667,N_6968,N_7318);
nand U7668 (N_7668,N_7065,N_7016);
or U7669 (N_7669,N_7021,N_6951);
or U7670 (N_7670,N_7041,N_7015);
or U7671 (N_7671,N_7250,N_6974);
or U7672 (N_7672,N_7172,N_7473);
nand U7673 (N_7673,N_7424,N_7287);
nor U7674 (N_7674,N_7093,N_7232);
xnor U7675 (N_7675,N_7154,N_7167);
xnor U7676 (N_7676,N_7135,N_7378);
xnor U7677 (N_7677,N_7085,N_7395);
xnor U7678 (N_7678,N_7208,N_7285);
or U7679 (N_7679,N_7104,N_6912);
nand U7680 (N_7680,N_7252,N_6996);
nand U7681 (N_7681,N_7235,N_6915);
nor U7682 (N_7682,N_6965,N_7069);
nor U7683 (N_7683,N_7325,N_6880);
or U7684 (N_7684,N_7470,N_6961);
nand U7685 (N_7685,N_7128,N_7278);
and U7686 (N_7686,N_7349,N_7058);
nor U7687 (N_7687,N_7157,N_6956);
or U7688 (N_7688,N_6958,N_7262);
xor U7689 (N_7689,N_7272,N_7031);
and U7690 (N_7690,N_7346,N_6901);
and U7691 (N_7691,N_6924,N_7432);
xnor U7692 (N_7692,N_7292,N_7296);
nor U7693 (N_7693,N_7162,N_7403);
xor U7694 (N_7694,N_6962,N_7076);
nand U7695 (N_7695,N_7137,N_7075);
xor U7696 (N_7696,N_6947,N_6911);
xor U7697 (N_7697,N_7416,N_7120);
nand U7698 (N_7698,N_7483,N_7469);
nand U7699 (N_7699,N_6964,N_7490);
nor U7700 (N_7700,N_6995,N_7458);
or U7701 (N_7701,N_7185,N_6930);
and U7702 (N_7702,N_6931,N_7370);
nand U7703 (N_7703,N_7090,N_7332);
or U7704 (N_7704,N_7306,N_7188);
or U7705 (N_7705,N_7124,N_7224);
nor U7706 (N_7706,N_7337,N_6932);
or U7707 (N_7707,N_7322,N_7418);
nor U7708 (N_7708,N_7467,N_7460);
and U7709 (N_7709,N_7472,N_7302);
nor U7710 (N_7710,N_7030,N_7313);
and U7711 (N_7711,N_7273,N_7243);
nor U7712 (N_7712,N_6987,N_7145);
or U7713 (N_7713,N_7122,N_7431);
and U7714 (N_7714,N_7077,N_7108);
and U7715 (N_7715,N_6891,N_7166);
nor U7716 (N_7716,N_7269,N_7303);
or U7717 (N_7717,N_6900,N_7171);
nor U7718 (N_7718,N_6888,N_7039);
and U7719 (N_7719,N_7121,N_7481);
nand U7720 (N_7720,N_6948,N_7280);
nand U7721 (N_7721,N_6878,N_7341);
xnor U7722 (N_7722,N_7018,N_7495);
nand U7723 (N_7723,N_6984,N_7244);
nor U7724 (N_7724,N_7105,N_6881);
nor U7725 (N_7725,N_7412,N_6988);
nand U7726 (N_7726,N_7496,N_7351);
nor U7727 (N_7727,N_7003,N_6917);
nand U7728 (N_7728,N_7130,N_7012);
xor U7729 (N_7729,N_6894,N_6919);
or U7730 (N_7730,N_7227,N_7340);
or U7731 (N_7731,N_7028,N_6954);
and U7732 (N_7732,N_7165,N_7133);
nand U7733 (N_7733,N_7211,N_7123);
and U7734 (N_7734,N_7434,N_7369);
and U7735 (N_7735,N_6952,N_7444);
nand U7736 (N_7736,N_7494,N_7115);
or U7737 (N_7737,N_7127,N_7445);
nand U7738 (N_7738,N_7466,N_7160);
nand U7739 (N_7739,N_7334,N_7471);
nand U7740 (N_7740,N_7487,N_6963);
nor U7741 (N_7741,N_7219,N_7284);
xnor U7742 (N_7742,N_7097,N_7189);
or U7743 (N_7743,N_7493,N_7407);
nand U7744 (N_7744,N_7379,N_6936);
or U7745 (N_7745,N_7435,N_7140);
or U7746 (N_7746,N_7486,N_7298);
or U7747 (N_7747,N_7081,N_7142);
nand U7748 (N_7748,N_7102,N_7118);
xnor U7749 (N_7749,N_7387,N_6899);
and U7750 (N_7750,N_7148,N_7163);
nand U7751 (N_7751,N_6920,N_7036);
or U7752 (N_7752,N_6925,N_7114);
and U7753 (N_7753,N_7380,N_7064);
nor U7754 (N_7754,N_7439,N_7383);
and U7755 (N_7755,N_7203,N_7274);
nand U7756 (N_7756,N_6991,N_6957);
and U7757 (N_7757,N_7237,N_7401);
or U7758 (N_7758,N_7098,N_7397);
nand U7759 (N_7759,N_7319,N_6943);
and U7760 (N_7760,N_6921,N_7498);
xnor U7761 (N_7761,N_7316,N_7034);
or U7762 (N_7762,N_7417,N_7480);
nand U7763 (N_7763,N_7443,N_7392);
or U7764 (N_7764,N_7484,N_7276);
or U7765 (N_7765,N_7116,N_7200);
nor U7766 (N_7766,N_7059,N_7336);
or U7767 (N_7767,N_7245,N_7288);
nand U7768 (N_7768,N_7038,N_7328);
xnor U7769 (N_7769,N_7107,N_7070);
and U7770 (N_7770,N_7184,N_7096);
and U7771 (N_7771,N_7271,N_7099);
nor U7772 (N_7772,N_7074,N_7384);
or U7773 (N_7773,N_6910,N_7260);
or U7774 (N_7774,N_7394,N_6890);
and U7775 (N_7775,N_7409,N_7170);
nand U7776 (N_7776,N_6877,N_7222);
or U7777 (N_7777,N_7478,N_7024);
and U7778 (N_7778,N_7242,N_7275);
or U7779 (N_7779,N_7177,N_7094);
nand U7780 (N_7780,N_6972,N_7186);
xnor U7781 (N_7781,N_7263,N_7461);
nand U7782 (N_7782,N_7078,N_6982);
nand U7783 (N_7783,N_7329,N_6939);
nor U7784 (N_7784,N_7264,N_7249);
nor U7785 (N_7785,N_7089,N_6992);
nor U7786 (N_7786,N_7231,N_6966);
or U7787 (N_7787,N_6944,N_7452);
xnor U7788 (N_7788,N_7063,N_7430);
xnor U7789 (N_7789,N_7331,N_7199);
or U7790 (N_7790,N_7088,N_7491);
or U7791 (N_7791,N_6940,N_7359);
nand U7792 (N_7792,N_7421,N_6909);
xnor U7793 (N_7793,N_7225,N_7415);
nand U7794 (N_7794,N_7198,N_6970);
nor U7795 (N_7795,N_6985,N_7236);
xnor U7796 (N_7796,N_7422,N_7492);
and U7797 (N_7797,N_7399,N_6885);
xnor U7798 (N_7798,N_7053,N_7488);
nand U7799 (N_7799,N_7281,N_7032);
and U7800 (N_7800,N_7320,N_7360);
or U7801 (N_7801,N_7158,N_7420);
or U7802 (N_7802,N_6902,N_7159);
nor U7803 (N_7803,N_7017,N_7201);
xnor U7804 (N_7804,N_7448,N_7327);
nor U7805 (N_7805,N_6895,N_7147);
and U7806 (N_7806,N_6892,N_7101);
and U7807 (N_7807,N_6989,N_7054);
nand U7808 (N_7808,N_7241,N_7258);
nor U7809 (N_7809,N_7060,N_7011);
nor U7810 (N_7810,N_7267,N_7173);
xnor U7811 (N_7811,N_6927,N_7013);
nor U7812 (N_7812,N_7027,N_7085);
or U7813 (N_7813,N_7249,N_7165);
xor U7814 (N_7814,N_7174,N_7352);
and U7815 (N_7815,N_7154,N_7029);
nand U7816 (N_7816,N_7223,N_6915);
or U7817 (N_7817,N_7275,N_7454);
nand U7818 (N_7818,N_7249,N_7047);
nand U7819 (N_7819,N_7430,N_7409);
and U7820 (N_7820,N_7175,N_7081);
or U7821 (N_7821,N_7112,N_7373);
xor U7822 (N_7822,N_7398,N_7019);
xnor U7823 (N_7823,N_6921,N_7328);
nand U7824 (N_7824,N_7488,N_7063);
nor U7825 (N_7825,N_6990,N_7160);
nand U7826 (N_7826,N_6888,N_7366);
nor U7827 (N_7827,N_7369,N_7453);
nand U7828 (N_7828,N_7428,N_7318);
and U7829 (N_7829,N_7386,N_7029);
nand U7830 (N_7830,N_7458,N_6942);
or U7831 (N_7831,N_7249,N_7098);
xnor U7832 (N_7832,N_7182,N_7384);
or U7833 (N_7833,N_6963,N_7139);
or U7834 (N_7834,N_7306,N_7213);
xor U7835 (N_7835,N_7407,N_7203);
xnor U7836 (N_7836,N_7010,N_7340);
and U7837 (N_7837,N_7368,N_6959);
or U7838 (N_7838,N_7053,N_7297);
or U7839 (N_7839,N_7084,N_7257);
and U7840 (N_7840,N_7016,N_7423);
xor U7841 (N_7841,N_7360,N_7445);
or U7842 (N_7842,N_7293,N_6943);
xor U7843 (N_7843,N_7285,N_6902);
xnor U7844 (N_7844,N_6883,N_7015);
xnor U7845 (N_7845,N_7186,N_7134);
or U7846 (N_7846,N_7324,N_7056);
xor U7847 (N_7847,N_7135,N_7012);
nor U7848 (N_7848,N_7158,N_7294);
and U7849 (N_7849,N_7222,N_7303);
and U7850 (N_7850,N_7148,N_7092);
nand U7851 (N_7851,N_7135,N_7250);
nand U7852 (N_7852,N_6900,N_7150);
and U7853 (N_7853,N_7485,N_7177);
nand U7854 (N_7854,N_7462,N_6940);
xnor U7855 (N_7855,N_7364,N_7114);
nand U7856 (N_7856,N_7040,N_7388);
xnor U7857 (N_7857,N_7076,N_7354);
xnor U7858 (N_7858,N_7266,N_7439);
nand U7859 (N_7859,N_6939,N_6931);
xor U7860 (N_7860,N_6875,N_7372);
nor U7861 (N_7861,N_7258,N_7237);
and U7862 (N_7862,N_7098,N_7061);
or U7863 (N_7863,N_7344,N_7402);
and U7864 (N_7864,N_7334,N_6931);
or U7865 (N_7865,N_7027,N_7158);
nor U7866 (N_7866,N_7431,N_7285);
or U7867 (N_7867,N_7018,N_6956);
and U7868 (N_7868,N_7151,N_7225);
nand U7869 (N_7869,N_7349,N_7122);
and U7870 (N_7870,N_7200,N_7359);
nand U7871 (N_7871,N_7431,N_7179);
and U7872 (N_7872,N_7168,N_7448);
nand U7873 (N_7873,N_7048,N_7057);
nor U7874 (N_7874,N_6975,N_7400);
or U7875 (N_7875,N_7106,N_7165);
nand U7876 (N_7876,N_7479,N_7031);
xor U7877 (N_7877,N_7472,N_6887);
nand U7878 (N_7878,N_6957,N_7010);
and U7879 (N_7879,N_7054,N_6950);
or U7880 (N_7880,N_7161,N_7165);
and U7881 (N_7881,N_7107,N_7034);
xor U7882 (N_7882,N_7076,N_7439);
or U7883 (N_7883,N_7113,N_6976);
nand U7884 (N_7884,N_7458,N_7119);
and U7885 (N_7885,N_7329,N_7031);
or U7886 (N_7886,N_7051,N_7295);
and U7887 (N_7887,N_7259,N_7450);
nor U7888 (N_7888,N_7298,N_7351);
nor U7889 (N_7889,N_6982,N_6909);
nand U7890 (N_7890,N_6875,N_7000);
or U7891 (N_7891,N_6979,N_7038);
or U7892 (N_7892,N_7172,N_6967);
xor U7893 (N_7893,N_7124,N_7303);
nor U7894 (N_7894,N_7405,N_7035);
xnor U7895 (N_7895,N_7288,N_7248);
nor U7896 (N_7896,N_7072,N_7487);
and U7897 (N_7897,N_7245,N_7233);
or U7898 (N_7898,N_7416,N_7132);
and U7899 (N_7899,N_7074,N_7003);
and U7900 (N_7900,N_6989,N_7308);
nand U7901 (N_7901,N_7001,N_6881);
xor U7902 (N_7902,N_7049,N_7053);
nor U7903 (N_7903,N_7249,N_7070);
and U7904 (N_7904,N_7034,N_6913);
and U7905 (N_7905,N_7447,N_7490);
or U7906 (N_7906,N_6977,N_7327);
xnor U7907 (N_7907,N_7301,N_7006);
xnor U7908 (N_7908,N_7305,N_7014);
xor U7909 (N_7909,N_6912,N_7066);
nand U7910 (N_7910,N_7381,N_6984);
nand U7911 (N_7911,N_7360,N_6989);
or U7912 (N_7912,N_7141,N_7324);
and U7913 (N_7913,N_7242,N_7110);
nand U7914 (N_7914,N_6901,N_7067);
xor U7915 (N_7915,N_7135,N_7023);
nor U7916 (N_7916,N_7427,N_7134);
nand U7917 (N_7917,N_7227,N_6905);
or U7918 (N_7918,N_7465,N_6957);
nor U7919 (N_7919,N_7265,N_7140);
nand U7920 (N_7920,N_6937,N_7156);
and U7921 (N_7921,N_7358,N_7263);
nand U7922 (N_7922,N_6981,N_7236);
nand U7923 (N_7923,N_7352,N_7097);
and U7924 (N_7924,N_7065,N_7371);
xnor U7925 (N_7925,N_7258,N_7179);
nor U7926 (N_7926,N_7390,N_7184);
xor U7927 (N_7927,N_6937,N_7228);
and U7928 (N_7928,N_7398,N_7440);
xnor U7929 (N_7929,N_6878,N_7273);
or U7930 (N_7930,N_7390,N_7386);
or U7931 (N_7931,N_7325,N_7278);
and U7932 (N_7932,N_7197,N_7205);
or U7933 (N_7933,N_7198,N_7274);
xnor U7934 (N_7934,N_7251,N_6885);
xor U7935 (N_7935,N_7449,N_7188);
and U7936 (N_7936,N_7206,N_7319);
or U7937 (N_7937,N_7450,N_6930);
nor U7938 (N_7938,N_6884,N_7290);
nor U7939 (N_7939,N_7099,N_6907);
nand U7940 (N_7940,N_7470,N_7469);
xnor U7941 (N_7941,N_7372,N_7235);
xor U7942 (N_7942,N_6877,N_7493);
xor U7943 (N_7943,N_7241,N_6909);
and U7944 (N_7944,N_6999,N_7268);
and U7945 (N_7945,N_7352,N_7423);
or U7946 (N_7946,N_7121,N_7164);
nor U7947 (N_7947,N_7461,N_7297);
or U7948 (N_7948,N_6987,N_7083);
nor U7949 (N_7949,N_7484,N_7219);
and U7950 (N_7950,N_7382,N_7209);
or U7951 (N_7951,N_7045,N_7402);
xor U7952 (N_7952,N_7037,N_6989);
nand U7953 (N_7953,N_7353,N_6888);
xor U7954 (N_7954,N_7205,N_6982);
xor U7955 (N_7955,N_7461,N_7037);
nor U7956 (N_7956,N_7321,N_7020);
nor U7957 (N_7957,N_7493,N_7254);
or U7958 (N_7958,N_6913,N_6888);
and U7959 (N_7959,N_7371,N_7340);
and U7960 (N_7960,N_7131,N_7034);
or U7961 (N_7961,N_7466,N_7061);
nand U7962 (N_7962,N_7080,N_7205);
and U7963 (N_7963,N_7176,N_6988);
or U7964 (N_7964,N_7048,N_7058);
xnor U7965 (N_7965,N_6936,N_6965);
xnor U7966 (N_7966,N_7234,N_7338);
or U7967 (N_7967,N_7152,N_7301);
and U7968 (N_7968,N_6923,N_7016);
or U7969 (N_7969,N_7292,N_7423);
or U7970 (N_7970,N_6891,N_7135);
xnor U7971 (N_7971,N_6953,N_7225);
and U7972 (N_7972,N_7243,N_7123);
nand U7973 (N_7973,N_7437,N_7151);
or U7974 (N_7974,N_7088,N_7180);
or U7975 (N_7975,N_7428,N_7451);
and U7976 (N_7976,N_7279,N_6968);
nand U7977 (N_7977,N_7248,N_7218);
or U7978 (N_7978,N_7029,N_7104);
and U7979 (N_7979,N_7034,N_7496);
nor U7980 (N_7980,N_6880,N_7337);
or U7981 (N_7981,N_7155,N_7103);
and U7982 (N_7982,N_6980,N_6921);
and U7983 (N_7983,N_7168,N_7232);
and U7984 (N_7984,N_7327,N_6890);
or U7985 (N_7985,N_7369,N_7109);
and U7986 (N_7986,N_7298,N_7444);
xnor U7987 (N_7987,N_7024,N_7250);
and U7988 (N_7988,N_7455,N_7386);
or U7989 (N_7989,N_7482,N_7221);
nand U7990 (N_7990,N_7293,N_7221);
and U7991 (N_7991,N_6876,N_7003);
xnor U7992 (N_7992,N_7222,N_7497);
nor U7993 (N_7993,N_7452,N_7454);
and U7994 (N_7994,N_7380,N_7248);
or U7995 (N_7995,N_7351,N_7294);
xor U7996 (N_7996,N_7269,N_7332);
or U7997 (N_7997,N_7133,N_7379);
and U7998 (N_7998,N_7110,N_7307);
or U7999 (N_7999,N_7258,N_7465);
and U8000 (N_8000,N_7222,N_7196);
nand U8001 (N_8001,N_7417,N_7110);
nand U8002 (N_8002,N_6903,N_7110);
or U8003 (N_8003,N_7064,N_7033);
and U8004 (N_8004,N_7416,N_7303);
or U8005 (N_8005,N_7294,N_7163);
xor U8006 (N_8006,N_7433,N_7180);
xor U8007 (N_8007,N_6992,N_7077);
and U8008 (N_8008,N_7117,N_7346);
xnor U8009 (N_8009,N_7419,N_7476);
nand U8010 (N_8010,N_7195,N_7155);
nand U8011 (N_8011,N_7066,N_7194);
xor U8012 (N_8012,N_6977,N_7164);
or U8013 (N_8013,N_7490,N_7253);
xnor U8014 (N_8014,N_7081,N_7344);
or U8015 (N_8015,N_7421,N_7069);
nor U8016 (N_8016,N_7137,N_7482);
or U8017 (N_8017,N_7445,N_7400);
and U8018 (N_8018,N_7321,N_7497);
nor U8019 (N_8019,N_7429,N_7002);
nand U8020 (N_8020,N_6988,N_7157);
and U8021 (N_8021,N_6922,N_6876);
nor U8022 (N_8022,N_7201,N_7098);
nand U8023 (N_8023,N_6996,N_7191);
nor U8024 (N_8024,N_7453,N_6979);
or U8025 (N_8025,N_7344,N_7123);
xor U8026 (N_8026,N_7118,N_6931);
nand U8027 (N_8027,N_7191,N_7356);
nor U8028 (N_8028,N_6918,N_7489);
nor U8029 (N_8029,N_7461,N_6956);
xor U8030 (N_8030,N_7179,N_7037);
and U8031 (N_8031,N_7112,N_7049);
xor U8032 (N_8032,N_7295,N_6889);
xnor U8033 (N_8033,N_6966,N_7455);
nand U8034 (N_8034,N_6947,N_7374);
nor U8035 (N_8035,N_6915,N_7038);
or U8036 (N_8036,N_7065,N_7359);
or U8037 (N_8037,N_7259,N_7094);
nor U8038 (N_8038,N_7133,N_6932);
nand U8039 (N_8039,N_7005,N_7010);
nor U8040 (N_8040,N_6921,N_7301);
and U8041 (N_8041,N_6879,N_7362);
nor U8042 (N_8042,N_7308,N_7247);
and U8043 (N_8043,N_7001,N_7203);
and U8044 (N_8044,N_7128,N_7291);
xnor U8045 (N_8045,N_7426,N_7027);
xor U8046 (N_8046,N_7123,N_6960);
nand U8047 (N_8047,N_7365,N_7212);
and U8048 (N_8048,N_7492,N_7380);
or U8049 (N_8049,N_7150,N_7329);
nand U8050 (N_8050,N_7027,N_7050);
nand U8051 (N_8051,N_7087,N_6908);
nor U8052 (N_8052,N_7107,N_7008);
or U8053 (N_8053,N_7333,N_7230);
nor U8054 (N_8054,N_7454,N_7054);
and U8055 (N_8055,N_6890,N_7378);
nand U8056 (N_8056,N_7327,N_6883);
nand U8057 (N_8057,N_7406,N_7019);
nor U8058 (N_8058,N_6911,N_7334);
xnor U8059 (N_8059,N_7383,N_7072);
nor U8060 (N_8060,N_6988,N_7416);
or U8061 (N_8061,N_7239,N_6950);
xnor U8062 (N_8062,N_7057,N_7469);
and U8063 (N_8063,N_7147,N_7478);
nor U8064 (N_8064,N_6888,N_6895);
or U8065 (N_8065,N_7166,N_7157);
nand U8066 (N_8066,N_7220,N_7148);
xnor U8067 (N_8067,N_6878,N_7001);
or U8068 (N_8068,N_7135,N_7397);
nand U8069 (N_8069,N_7010,N_7399);
nand U8070 (N_8070,N_6898,N_7184);
nand U8071 (N_8071,N_7269,N_7163);
and U8072 (N_8072,N_6964,N_7085);
nor U8073 (N_8073,N_6985,N_6976);
nor U8074 (N_8074,N_7337,N_7324);
nor U8075 (N_8075,N_6937,N_6879);
and U8076 (N_8076,N_7202,N_7260);
and U8077 (N_8077,N_6903,N_7216);
nor U8078 (N_8078,N_7216,N_7162);
and U8079 (N_8079,N_7049,N_7116);
or U8080 (N_8080,N_6899,N_7321);
nand U8081 (N_8081,N_7430,N_6978);
and U8082 (N_8082,N_7060,N_7057);
xor U8083 (N_8083,N_7047,N_6944);
nor U8084 (N_8084,N_7411,N_7451);
nor U8085 (N_8085,N_7045,N_7365);
and U8086 (N_8086,N_6882,N_7198);
nor U8087 (N_8087,N_7046,N_6957);
nand U8088 (N_8088,N_7250,N_7131);
and U8089 (N_8089,N_7492,N_6975);
and U8090 (N_8090,N_6877,N_6888);
nand U8091 (N_8091,N_7457,N_7472);
nor U8092 (N_8092,N_7120,N_6952);
xnor U8093 (N_8093,N_7409,N_7021);
or U8094 (N_8094,N_7320,N_7058);
nor U8095 (N_8095,N_6884,N_7055);
nand U8096 (N_8096,N_7056,N_7192);
nor U8097 (N_8097,N_7037,N_6887);
and U8098 (N_8098,N_7420,N_7046);
xor U8099 (N_8099,N_7025,N_7323);
nor U8100 (N_8100,N_7344,N_7306);
nand U8101 (N_8101,N_7306,N_7257);
nand U8102 (N_8102,N_7028,N_6977);
xnor U8103 (N_8103,N_7085,N_7241);
or U8104 (N_8104,N_7020,N_6903);
xor U8105 (N_8105,N_7185,N_7139);
nand U8106 (N_8106,N_7088,N_7131);
or U8107 (N_8107,N_7386,N_7146);
nor U8108 (N_8108,N_7348,N_6944);
nor U8109 (N_8109,N_6936,N_7053);
nand U8110 (N_8110,N_6903,N_7061);
nor U8111 (N_8111,N_7185,N_6971);
or U8112 (N_8112,N_6948,N_6962);
nand U8113 (N_8113,N_7450,N_7331);
nand U8114 (N_8114,N_7134,N_7097);
or U8115 (N_8115,N_6919,N_7408);
or U8116 (N_8116,N_6880,N_7112);
nand U8117 (N_8117,N_6898,N_7132);
xnor U8118 (N_8118,N_7244,N_7303);
xnor U8119 (N_8119,N_7043,N_7483);
xnor U8120 (N_8120,N_7061,N_7344);
nor U8121 (N_8121,N_7225,N_7289);
or U8122 (N_8122,N_7437,N_7099);
nand U8123 (N_8123,N_7263,N_7342);
xor U8124 (N_8124,N_6939,N_7394);
nor U8125 (N_8125,N_7512,N_7780);
xnor U8126 (N_8126,N_7667,N_7980);
or U8127 (N_8127,N_8062,N_7905);
nand U8128 (N_8128,N_7990,N_8102);
and U8129 (N_8129,N_7576,N_7888);
nor U8130 (N_8130,N_7540,N_8040);
or U8131 (N_8131,N_7515,N_8099);
or U8132 (N_8132,N_7580,N_7859);
and U8133 (N_8133,N_7665,N_7509);
and U8134 (N_8134,N_7839,N_7851);
and U8135 (N_8135,N_7841,N_8006);
xor U8136 (N_8136,N_8095,N_7877);
xor U8137 (N_8137,N_8088,N_7510);
nor U8138 (N_8138,N_7744,N_7717);
and U8139 (N_8139,N_7567,N_7982);
nand U8140 (N_8140,N_8120,N_8078);
nand U8141 (N_8141,N_7882,N_7796);
nand U8142 (N_8142,N_7828,N_7874);
nand U8143 (N_8143,N_7958,N_7899);
nor U8144 (N_8144,N_7765,N_7528);
nor U8145 (N_8145,N_8104,N_7811);
nand U8146 (N_8146,N_7908,N_8009);
or U8147 (N_8147,N_7670,N_7645);
xor U8148 (N_8148,N_7994,N_7909);
xnor U8149 (N_8149,N_7834,N_7729);
or U8150 (N_8150,N_7936,N_7588);
or U8151 (N_8151,N_7624,N_7976);
nand U8152 (N_8152,N_7916,N_7803);
nand U8153 (N_8153,N_7770,N_7548);
nand U8154 (N_8154,N_7687,N_7832);
or U8155 (N_8155,N_7883,N_7594);
nor U8156 (N_8156,N_7894,N_7791);
nor U8157 (N_8157,N_7947,N_7955);
nand U8158 (N_8158,N_7995,N_7745);
nor U8159 (N_8159,N_7607,N_7904);
or U8160 (N_8160,N_7983,N_7733);
and U8161 (N_8161,N_7961,N_7919);
or U8162 (N_8162,N_7924,N_7578);
or U8163 (N_8163,N_7783,N_7569);
nand U8164 (N_8164,N_7560,N_7853);
xor U8165 (N_8165,N_7655,N_7820);
and U8166 (N_8166,N_7866,N_7558);
or U8167 (N_8167,N_7819,N_7704);
and U8168 (N_8168,N_7572,N_7684);
xor U8169 (N_8169,N_7554,N_7668);
and U8170 (N_8170,N_7561,N_8085);
xnor U8171 (N_8171,N_7547,N_7511);
xor U8172 (N_8172,N_7603,N_8034);
and U8173 (N_8173,N_7968,N_8056);
nor U8174 (N_8174,N_7914,N_7585);
xnor U8175 (N_8175,N_8019,N_7997);
or U8176 (N_8176,N_7829,N_7731);
and U8177 (N_8177,N_7844,N_7570);
nor U8178 (N_8178,N_7973,N_8101);
and U8179 (N_8179,N_8110,N_7868);
xnor U8180 (N_8180,N_7775,N_8048);
nor U8181 (N_8181,N_7934,N_7969);
and U8182 (N_8182,N_8025,N_7971);
nand U8183 (N_8183,N_7940,N_8045);
xnor U8184 (N_8184,N_7505,N_7598);
nand U8185 (N_8185,N_8115,N_8039);
nor U8186 (N_8186,N_7503,N_7777);
and U8187 (N_8187,N_7930,N_7771);
nor U8188 (N_8188,N_7690,N_7843);
and U8189 (N_8189,N_7565,N_8058);
xnor U8190 (N_8190,N_7628,N_7721);
nand U8191 (N_8191,N_7521,N_7525);
nand U8192 (N_8192,N_7761,N_8026);
nor U8193 (N_8193,N_8066,N_7998);
or U8194 (N_8194,N_7591,N_7692);
or U8195 (N_8195,N_7822,N_7858);
nand U8196 (N_8196,N_7630,N_7825);
nand U8197 (N_8197,N_7933,N_8046);
and U8198 (N_8198,N_7517,N_7694);
nand U8199 (N_8199,N_7575,N_7666);
nor U8200 (N_8200,N_7946,N_8005);
nand U8201 (N_8201,N_8043,N_7880);
nor U8202 (N_8202,N_8053,N_8057);
xnor U8203 (N_8203,N_7629,N_7647);
xnor U8204 (N_8204,N_7559,N_8084);
or U8205 (N_8205,N_7649,N_7696);
nand U8206 (N_8206,N_7891,N_7810);
xnor U8207 (N_8207,N_7680,N_7600);
and U8208 (N_8208,N_7732,N_8074);
nand U8209 (N_8209,N_7508,N_7582);
nor U8210 (N_8210,N_8021,N_7621);
nor U8211 (N_8211,N_7974,N_7720);
or U8212 (N_8212,N_7644,N_7773);
and U8213 (N_8213,N_7938,N_7897);
or U8214 (N_8214,N_7781,N_7756);
xnor U8215 (N_8215,N_7746,N_7650);
nor U8216 (N_8216,N_8018,N_7623);
nand U8217 (N_8217,N_7957,N_7590);
and U8218 (N_8218,N_7748,N_7960);
or U8219 (N_8219,N_8013,N_7929);
xor U8220 (N_8220,N_7823,N_7710);
xor U8221 (N_8221,N_7817,N_7906);
nor U8222 (N_8222,N_7893,N_7790);
and U8223 (N_8223,N_8028,N_7978);
and U8224 (N_8224,N_8059,N_8033);
xor U8225 (N_8225,N_7776,N_7619);
nand U8226 (N_8226,N_8075,N_7672);
nor U8227 (N_8227,N_7656,N_7869);
nor U8228 (N_8228,N_7543,N_7638);
nand U8229 (N_8229,N_7852,N_7555);
xor U8230 (N_8230,N_7573,N_7737);
nand U8231 (N_8231,N_7513,N_7681);
or U8232 (N_8232,N_7949,N_8086);
and U8233 (N_8233,N_7798,N_7945);
nor U8234 (N_8234,N_7967,N_7760);
xnor U8235 (N_8235,N_7890,N_8041);
or U8236 (N_8236,N_7674,N_7571);
nor U8237 (N_8237,N_7531,N_7743);
nor U8238 (N_8238,N_7682,N_7956);
and U8239 (N_8239,N_7886,N_7802);
xnor U8240 (N_8240,N_7614,N_7609);
or U8241 (N_8241,N_7845,N_7700);
nor U8242 (N_8242,N_7794,N_7661);
nand U8243 (N_8243,N_8098,N_7759);
or U8244 (N_8244,N_7730,N_7912);
xor U8245 (N_8245,N_7651,N_8010);
xor U8246 (N_8246,N_8068,N_7975);
and U8247 (N_8247,N_8094,N_7738);
or U8248 (N_8248,N_7856,N_7596);
xnor U8249 (N_8249,N_7915,N_7636);
xnor U8250 (N_8250,N_7863,N_8001);
nor U8251 (N_8251,N_7734,N_7787);
or U8252 (N_8252,N_7762,N_7772);
xor U8253 (N_8253,N_7532,N_7586);
nor U8254 (N_8254,N_8020,N_8035);
or U8255 (N_8255,N_7988,N_8014);
or U8256 (N_8256,N_7950,N_7814);
nor U8257 (N_8257,N_7827,N_7602);
nor U8258 (N_8258,N_7935,N_7993);
nor U8259 (N_8259,N_7617,N_7754);
xor U8260 (N_8260,N_7835,N_7952);
xnor U8261 (N_8261,N_7922,N_7766);
nand U8262 (N_8262,N_7657,N_8060);
nor U8263 (N_8263,N_7648,N_7689);
nand U8264 (N_8264,N_7574,N_7695);
xor U8265 (N_8265,N_7769,N_7778);
or U8266 (N_8266,N_7849,N_7907);
xnor U8267 (N_8267,N_7707,N_7847);
nor U8268 (N_8268,N_8063,N_8073);
nor U8269 (N_8269,N_8114,N_7826);
or U8270 (N_8270,N_7941,N_7895);
nor U8271 (N_8271,N_7615,N_7669);
xnor U8272 (N_8272,N_7688,N_8113);
or U8273 (N_8273,N_7693,N_8089);
xor U8274 (N_8274,N_8090,N_7753);
or U8275 (N_8275,N_8122,N_7719);
xor U8276 (N_8276,N_8007,N_7676);
xor U8277 (N_8277,N_7501,N_7706);
or U8278 (N_8278,N_8012,N_7870);
xnor U8279 (N_8279,N_7943,N_8047);
xnor U8280 (N_8280,N_7901,N_7979);
and U8281 (N_8281,N_7923,N_7833);
xnor U8282 (N_8282,N_7807,N_7885);
or U8283 (N_8283,N_7857,N_7726);
xnor U8284 (N_8284,N_8118,N_7599);
or U8285 (N_8285,N_7631,N_7544);
or U8286 (N_8286,N_7673,N_8091);
nand U8287 (N_8287,N_7812,N_7884);
nand U8288 (N_8288,N_7824,N_7653);
and U8289 (N_8289,N_8016,N_7537);
and U8290 (N_8290,N_7677,N_7821);
xnor U8291 (N_8291,N_7966,N_7768);
nor U8292 (N_8292,N_8002,N_8017);
and U8293 (N_8293,N_7984,N_7724);
or U8294 (N_8294,N_7577,N_7813);
nor U8295 (N_8295,N_7881,N_8054);
or U8296 (N_8296,N_7977,N_8042);
and U8297 (N_8297,N_7605,N_8107);
nand U8298 (N_8298,N_7900,N_7774);
or U8299 (N_8299,N_7937,N_7878);
nor U8300 (N_8300,N_7529,N_7523);
and U8301 (N_8301,N_7757,N_7889);
or U8302 (N_8302,N_7806,N_7535);
xnor U8303 (N_8303,N_7522,N_8079);
and U8304 (N_8304,N_7864,N_7902);
nand U8305 (N_8305,N_8105,N_7542);
or U8306 (N_8306,N_7948,N_7725);
and U8307 (N_8307,N_7683,N_7991);
nor U8308 (N_8308,N_7727,N_7646);
xnor U8309 (N_8309,N_7972,N_7658);
nand U8310 (N_8310,N_7742,N_7703);
nor U8311 (N_8311,N_8011,N_7691);
nand U8312 (N_8312,N_8067,N_7604);
xnor U8313 (N_8313,N_7622,N_7837);
nor U8314 (N_8314,N_7541,N_7705);
nor U8315 (N_8315,N_7792,N_7557);
and U8316 (N_8316,N_8087,N_7662);
nand U8317 (N_8317,N_7855,N_7723);
nor U8318 (N_8318,N_7583,N_7921);
or U8319 (N_8319,N_7981,N_7925);
or U8320 (N_8320,N_7939,N_8071);
nor U8321 (N_8321,N_7504,N_7763);
xnor U8322 (N_8322,N_7740,N_7741);
or U8323 (N_8323,N_7992,N_7799);
and U8324 (N_8324,N_7838,N_7698);
xnor U8325 (N_8325,N_7809,N_8032);
or U8326 (N_8326,N_7918,N_8050);
nor U8327 (N_8327,N_7788,N_7536);
xor U8328 (N_8328,N_7702,N_7663);
xnor U8329 (N_8329,N_7711,N_7533);
nand U8330 (N_8330,N_7808,N_8061);
xnor U8331 (N_8331,N_7751,N_8037);
nor U8332 (N_8332,N_7597,N_8072);
or U8333 (N_8333,N_7618,N_7749);
or U8334 (N_8334,N_7970,N_7678);
and U8335 (N_8335,N_7875,N_7767);
nand U8336 (N_8336,N_7516,N_7660);
and U8337 (N_8337,N_8038,N_7758);
nor U8338 (N_8338,N_8024,N_7860);
nand U8339 (N_8339,N_7962,N_7639);
xor U8340 (N_8340,N_7551,N_7625);
or U8341 (N_8341,N_8109,N_7716);
nand U8342 (N_8342,N_8022,N_7611);
or U8343 (N_8343,N_7926,N_7944);
nor U8344 (N_8344,N_7502,N_7739);
and U8345 (N_8345,N_7785,N_8000);
nand U8346 (N_8346,N_7862,N_7552);
and U8347 (N_8347,N_7584,N_7816);
and U8348 (N_8348,N_7932,N_7784);
nand U8349 (N_8349,N_7804,N_7831);
and U8350 (N_8350,N_7654,N_8029);
or U8351 (N_8351,N_7910,N_7954);
and U8352 (N_8352,N_7718,N_7527);
xnor U8353 (N_8353,N_7846,N_7592);
and U8354 (N_8354,N_7634,N_7854);
nand U8355 (N_8355,N_7500,N_7755);
nor U8356 (N_8356,N_7850,N_7587);
or U8357 (N_8357,N_7986,N_7985);
and U8358 (N_8358,N_8082,N_7606);
xor U8359 (N_8359,N_8030,N_7610);
xor U8360 (N_8360,N_8117,N_7715);
and U8361 (N_8361,N_7612,N_7556);
and U8362 (N_8362,N_8097,N_7818);
nand U8363 (N_8363,N_8027,N_7671);
nor U8364 (N_8364,N_7686,N_8015);
nand U8365 (N_8365,N_8003,N_7633);
nor U8366 (N_8366,N_8069,N_7830);
nand U8367 (N_8367,N_8051,N_7876);
and U8368 (N_8368,N_8064,N_7728);
or U8369 (N_8369,N_7538,N_8055);
xor U8370 (N_8370,N_7566,N_7911);
xor U8371 (N_8371,N_8083,N_7913);
nand U8372 (N_8372,N_7616,N_7549);
xnor U8373 (N_8373,N_7917,N_7514);
or U8374 (N_8374,N_8008,N_7519);
or U8375 (N_8375,N_8036,N_7959);
or U8376 (N_8376,N_8103,N_8044);
xor U8377 (N_8377,N_7652,N_8081);
xnor U8378 (N_8378,N_7736,N_7953);
or U8379 (N_8379,N_7563,N_7685);
and U8380 (N_8380,N_7553,N_7534);
and U8381 (N_8381,N_7550,N_7701);
and U8382 (N_8382,N_7805,N_7848);
and U8383 (N_8383,N_7530,N_8116);
and U8384 (N_8384,N_7581,N_7659);
xnor U8385 (N_8385,N_7896,N_8106);
or U8386 (N_8386,N_7520,N_7632);
and U8387 (N_8387,N_7708,N_7524);
nand U8388 (N_8388,N_8124,N_7526);
or U8389 (N_8389,N_7815,N_7562);
nor U8390 (N_8390,N_8080,N_7867);
and U8391 (N_8391,N_8100,N_7795);
nor U8392 (N_8392,N_7786,N_8093);
and U8393 (N_8393,N_7965,N_8004);
and U8394 (N_8394,N_7920,N_7989);
xnor U8395 (N_8395,N_8031,N_7518);
xor U8396 (N_8396,N_7507,N_7879);
nand U8397 (N_8397,N_7564,N_8092);
nand U8398 (N_8398,N_7568,N_7903);
and U8399 (N_8399,N_7842,N_7620);
and U8400 (N_8400,N_7865,N_8112);
or U8401 (N_8401,N_7931,N_7699);
nor U8402 (N_8402,N_8065,N_7928);
nor U8403 (N_8403,N_7840,N_7709);
or U8404 (N_8404,N_8076,N_7861);
nand U8405 (N_8405,N_7964,N_7873);
nand U8406 (N_8406,N_7735,N_7963);
nor U8407 (N_8407,N_7872,N_8096);
nand U8408 (N_8408,N_7539,N_7892);
nand U8409 (N_8409,N_7898,N_7797);
or U8410 (N_8410,N_7640,N_7627);
nand U8411 (N_8411,N_7579,N_7764);
nor U8412 (N_8412,N_7595,N_7793);
and U8413 (N_8413,N_7800,N_7675);
or U8414 (N_8414,N_7601,N_7545);
or U8415 (N_8415,N_7801,N_7608);
xnor U8416 (N_8416,N_7871,N_8070);
and U8417 (N_8417,N_7643,N_7836);
xnor U8418 (N_8418,N_7782,N_8023);
or U8419 (N_8419,N_7546,N_8119);
and U8420 (N_8420,N_7752,N_7999);
or U8421 (N_8421,N_7712,N_7642);
and U8422 (N_8422,N_7626,N_8077);
xnor U8423 (N_8423,N_7714,N_8111);
nor U8424 (N_8424,N_7613,N_7951);
or U8425 (N_8425,N_7713,N_7789);
xnor U8426 (N_8426,N_8121,N_7747);
nor U8427 (N_8427,N_7722,N_7589);
or U8428 (N_8428,N_7987,N_7697);
and U8429 (N_8429,N_7750,N_8108);
nor U8430 (N_8430,N_7635,N_7679);
nor U8431 (N_8431,N_7593,N_7942);
or U8432 (N_8432,N_7887,N_7927);
or U8433 (N_8433,N_8123,N_7641);
nand U8434 (N_8434,N_8049,N_7664);
nor U8435 (N_8435,N_8052,N_7506);
xor U8436 (N_8436,N_7996,N_7779);
and U8437 (N_8437,N_7637,N_7987);
and U8438 (N_8438,N_7853,N_7716);
nand U8439 (N_8439,N_8008,N_7681);
or U8440 (N_8440,N_8097,N_7544);
or U8441 (N_8441,N_7988,N_7930);
xnor U8442 (N_8442,N_8038,N_8045);
or U8443 (N_8443,N_8088,N_7563);
nand U8444 (N_8444,N_7643,N_8067);
nand U8445 (N_8445,N_7804,N_7891);
nand U8446 (N_8446,N_7647,N_7926);
or U8447 (N_8447,N_7892,N_8112);
nor U8448 (N_8448,N_7614,N_7668);
and U8449 (N_8449,N_7723,N_7555);
nand U8450 (N_8450,N_8066,N_7545);
or U8451 (N_8451,N_7738,N_7876);
and U8452 (N_8452,N_7937,N_7992);
nor U8453 (N_8453,N_7676,N_7597);
and U8454 (N_8454,N_7673,N_7681);
nor U8455 (N_8455,N_7694,N_7528);
and U8456 (N_8456,N_7859,N_7972);
and U8457 (N_8457,N_7523,N_7694);
xnor U8458 (N_8458,N_7638,N_7583);
nand U8459 (N_8459,N_7880,N_7803);
or U8460 (N_8460,N_8063,N_7954);
nor U8461 (N_8461,N_7762,N_7602);
nor U8462 (N_8462,N_7550,N_7813);
nand U8463 (N_8463,N_7889,N_7857);
nand U8464 (N_8464,N_7579,N_8020);
xnor U8465 (N_8465,N_7769,N_7809);
nor U8466 (N_8466,N_7817,N_7827);
nand U8467 (N_8467,N_7963,N_7907);
or U8468 (N_8468,N_8047,N_7554);
nand U8469 (N_8469,N_7759,N_7668);
xor U8470 (N_8470,N_7945,N_7643);
xor U8471 (N_8471,N_8037,N_7916);
xnor U8472 (N_8472,N_7831,N_7617);
nand U8473 (N_8473,N_7852,N_7674);
nand U8474 (N_8474,N_7813,N_8100);
and U8475 (N_8475,N_7813,N_7837);
xor U8476 (N_8476,N_7739,N_7906);
xor U8477 (N_8477,N_7536,N_8027);
or U8478 (N_8478,N_7634,N_7514);
and U8479 (N_8479,N_7782,N_8046);
nand U8480 (N_8480,N_7538,N_7999);
nand U8481 (N_8481,N_7905,N_7668);
xor U8482 (N_8482,N_7695,N_7969);
nor U8483 (N_8483,N_7531,N_7577);
nor U8484 (N_8484,N_7958,N_7804);
nor U8485 (N_8485,N_7516,N_7982);
nor U8486 (N_8486,N_7520,N_7642);
or U8487 (N_8487,N_7730,N_7909);
nor U8488 (N_8488,N_7975,N_7865);
nor U8489 (N_8489,N_7535,N_7504);
or U8490 (N_8490,N_7756,N_7805);
and U8491 (N_8491,N_7601,N_7658);
or U8492 (N_8492,N_8116,N_7630);
nor U8493 (N_8493,N_8065,N_7909);
nand U8494 (N_8494,N_7967,N_7880);
and U8495 (N_8495,N_7896,N_7850);
nor U8496 (N_8496,N_8005,N_7936);
xnor U8497 (N_8497,N_7506,N_7959);
and U8498 (N_8498,N_8044,N_7661);
nand U8499 (N_8499,N_7717,N_7509);
or U8500 (N_8500,N_7974,N_7951);
nand U8501 (N_8501,N_7528,N_7639);
nand U8502 (N_8502,N_8094,N_7904);
xor U8503 (N_8503,N_7577,N_8083);
and U8504 (N_8504,N_7749,N_8015);
and U8505 (N_8505,N_7921,N_7709);
or U8506 (N_8506,N_7707,N_7776);
nor U8507 (N_8507,N_7929,N_8064);
nand U8508 (N_8508,N_7947,N_7690);
nand U8509 (N_8509,N_7870,N_8040);
nand U8510 (N_8510,N_7910,N_8059);
and U8511 (N_8511,N_7724,N_7913);
nand U8512 (N_8512,N_7707,N_7580);
nand U8513 (N_8513,N_7803,N_7924);
or U8514 (N_8514,N_8085,N_7926);
nand U8515 (N_8515,N_7529,N_7838);
nand U8516 (N_8516,N_7996,N_7522);
and U8517 (N_8517,N_7516,N_7634);
nand U8518 (N_8518,N_7599,N_7973);
nand U8519 (N_8519,N_7532,N_7995);
nor U8520 (N_8520,N_8023,N_7875);
nor U8521 (N_8521,N_7589,N_7666);
nand U8522 (N_8522,N_7529,N_8034);
nand U8523 (N_8523,N_7589,N_7967);
or U8524 (N_8524,N_7986,N_7718);
nand U8525 (N_8525,N_7956,N_7963);
xor U8526 (N_8526,N_7942,N_7652);
xnor U8527 (N_8527,N_7946,N_7991);
nand U8528 (N_8528,N_8031,N_7763);
nor U8529 (N_8529,N_7784,N_7720);
or U8530 (N_8530,N_8051,N_7666);
and U8531 (N_8531,N_8035,N_7930);
and U8532 (N_8532,N_8115,N_7705);
nand U8533 (N_8533,N_8087,N_7627);
nand U8534 (N_8534,N_8102,N_7925);
xor U8535 (N_8535,N_7922,N_7924);
or U8536 (N_8536,N_7621,N_8039);
or U8537 (N_8537,N_7634,N_7815);
xnor U8538 (N_8538,N_7509,N_7973);
nand U8539 (N_8539,N_7544,N_7710);
nor U8540 (N_8540,N_7724,N_8078);
or U8541 (N_8541,N_7864,N_7550);
xor U8542 (N_8542,N_7720,N_7757);
or U8543 (N_8543,N_7531,N_7704);
or U8544 (N_8544,N_7580,N_7637);
nand U8545 (N_8545,N_7636,N_7761);
nand U8546 (N_8546,N_7951,N_7770);
xor U8547 (N_8547,N_8007,N_7787);
and U8548 (N_8548,N_7854,N_7585);
xor U8549 (N_8549,N_7926,N_7690);
and U8550 (N_8550,N_8065,N_7862);
or U8551 (N_8551,N_7581,N_7520);
and U8552 (N_8552,N_8050,N_7544);
xnor U8553 (N_8553,N_7631,N_7643);
nand U8554 (N_8554,N_7793,N_8018);
nand U8555 (N_8555,N_7704,N_7716);
and U8556 (N_8556,N_7905,N_7987);
nor U8557 (N_8557,N_7569,N_8073);
nand U8558 (N_8558,N_8077,N_7853);
nand U8559 (N_8559,N_8084,N_8022);
nor U8560 (N_8560,N_8121,N_7926);
nand U8561 (N_8561,N_7611,N_7948);
and U8562 (N_8562,N_7812,N_7848);
or U8563 (N_8563,N_8044,N_7881);
xnor U8564 (N_8564,N_7866,N_7503);
and U8565 (N_8565,N_8049,N_7863);
nor U8566 (N_8566,N_7797,N_7866);
xor U8567 (N_8567,N_7858,N_7618);
nor U8568 (N_8568,N_7868,N_7564);
nand U8569 (N_8569,N_8035,N_7835);
nand U8570 (N_8570,N_7692,N_7894);
nand U8571 (N_8571,N_8021,N_7584);
nand U8572 (N_8572,N_7964,N_8108);
or U8573 (N_8573,N_7762,N_7633);
nand U8574 (N_8574,N_8068,N_7516);
nand U8575 (N_8575,N_8086,N_7969);
and U8576 (N_8576,N_7724,N_7675);
or U8577 (N_8577,N_7658,N_7976);
or U8578 (N_8578,N_7681,N_8116);
and U8579 (N_8579,N_7790,N_7761);
and U8580 (N_8580,N_7976,N_7715);
xnor U8581 (N_8581,N_8085,N_7530);
xor U8582 (N_8582,N_8100,N_7989);
and U8583 (N_8583,N_7653,N_7512);
xor U8584 (N_8584,N_7842,N_8061);
and U8585 (N_8585,N_7511,N_7917);
xor U8586 (N_8586,N_7737,N_7605);
nand U8587 (N_8587,N_8079,N_7697);
nor U8588 (N_8588,N_7598,N_7923);
and U8589 (N_8589,N_7825,N_7692);
xor U8590 (N_8590,N_7939,N_7821);
and U8591 (N_8591,N_7629,N_7718);
nor U8592 (N_8592,N_7690,N_8000);
xnor U8593 (N_8593,N_7638,N_7827);
or U8594 (N_8594,N_7932,N_7752);
or U8595 (N_8595,N_7842,N_7507);
nand U8596 (N_8596,N_8038,N_7981);
nor U8597 (N_8597,N_7855,N_7612);
and U8598 (N_8598,N_8034,N_7699);
xnor U8599 (N_8599,N_7503,N_7621);
or U8600 (N_8600,N_7977,N_7845);
nor U8601 (N_8601,N_7817,N_7900);
or U8602 (N_8602,N_7820,N_8081);
nor U8603 (N_8603,N_7823,N_7837);
xnor U8604 (N_8604,N_7747,N_7722);
or U8605 (N_8605,N_7851,N_7910);
or U8606 (N_8606,N_7724,N_7700);
nor U8607 (N_8607,N_7865,N_7591);
nand U8608 (N_8608,N_8089,N_7554);
xnor U8609 (N_8609,N_8017,N_7824);
nand U8610 (N_8610,N_7716,N_7786);
and U8611 (N_8611,N_8018,N_7681);
xnor U8612 (N_8612,N_7754,N_7788);
xnor U8613 (N_8613,N_7502,N_7892);
and U8614 (N_8614,N_7654,N_7521);
or U8615 (N_8615,N_7885,N_7751);
and U8616 (N_8616,N_8079,N_7983);
nor U8617 (N_8617,N_7896,N_8025);
or U8618 (N_8618,N_7756,N_7501);
or U8619 (N_8619,N_8102,N_8077);
and U8620 (N_8620,N_7705,N_8034);
nand U8621 (N_8621,N_7710,N_8028);
nor U8622 (N_8622,N_7824,N_7805);
or U8623 (N_8623,N_8094,N_8007);
or U8624 (N_8624,N_7878,N_7739);
nor U8625 (N_8625,N_7503,N_7793);
nor U8626 (N_8626,N_8079,N_7934);
xnor U8627 (N_8627,N_7859,N_7533);
and U8628 (N_8628,N_7962,N_7783);
nand U8629 (N_8629,N_8073,N_7711);
nand U8630 (N_8630,N_8119,N_7563);
and U8631 (N_8631,N_7572,N_7774);
or U8632 (N_8632,N_7906,N_7823);
nor U8633 (N_8633,N_7751,N_7511);
or U8634 (N_8634,N_7522,N_7568);
and U8635 (N_8635,N_7518,N_7509);
nand U8636 (N_8636,N_7845,N_7703);
nor U8637 (N_8637,N_7716,N_7838);
nor U8638 (N_8638,N_7634,N_8073);
or U8639 (N_8639,N_7736,N_7890);
and U8640 (N_8640,N_7693,N_7873);
nand U8641 (N_8641,N_8020,N_7830);
xnor U8642 (N_8642,N_7547,N_7889);
nand U8643 (N_8643,N_7824,N_7679);
xor U8644 (N_8644,N_7953,N_7810);
nand U8645 (N_8645,N_7983,N_7885);
nand U8646 (N_8646,N_7647,N_7667);
and U8647 (N_8647,N_7540,N_7557);
nor U8648 (N_8648,N_7894,N_8009);
and U8649 (N_8649,N_7524,N_8053);
nor U8650 (N_8650,N_7672,N_7946);
or U8651 (N_8651,N_7912,N_8056);
or U8652 (N_8652,N_7719,N_8016);
and U8653 (N_8653,N_7747,N_7691);
xnor U8654 (N_8654,N_7660,N_7710);
or U8655 (N_8655,N_8049,N_8041);
nand U8656 (N_8656,N_7740,N_8105);
nor U8657 (N_8657,N_8118,N_7922);
xor U8658 (N_8658,N_7548,N_7692);
xor U8659 (N_8659,N_7676,N_7748);
nand U8660 (N_8660,N_7861,N_7981);
nor U8661 (N_8661,N_8089,N_7639);
xor U8662 (N_8662,N_7665,N_7577);
xor U8663 (N_8663,N_8050,N_8035);
xor U8664 (N_8664,N_7848,N_7840);
nor U8665 (N_8665,N_7907,N_8100);
xor U8666 (N_8666,N_8104,N_8013);
xnor U8667 (N_8667,N_7622,N_7639);
xnor U8668 (N_8668,N_7622,N_7892);
or U8669 (N_8669,N_7877,N_8037);
nand U8670 (N_8670,N_7599,N_7902);
and U8671 (N_8671,N_7869,N_7710);
or U8672 (N_8672,N_7580,N_7760);
nor U8673 (N_8673,N_7895,N_7571);
and U8674 (N_8674,N_7679,N_8073);
and U8675 (N_8675,N_7976,N_7794);
nand U8676 (N_8676,N_7719,N_7879);
and U8677 (N_8677,N_8056,N_7577);
xor U8678 (N_8678,N_8101,N_7526);
nand U8679 (N_8679,N_7906,N_7653);
nand U8680 (N_8680,N_7621,N_7907);
nor U8681 (N_8681,N_7743,N_7879);
nor U8682 (N_8682,N_7814,N_7900);
and U8683 (N_8683,N_7525,N_8103);
nand U8684 (N_8684,N_8036,N_7675);
or U8685 (N_8685,N_7988,N_8097);
nand U8686 (N_8686,N_7646,N_8009);
and U8687 (N_8687,N_7679,N_8065);
xnor U8688 (N_8688,N_7636,N_7611);
xor U8689 (N_8689,N_7645,N_7692);
nor U8690 (N_8690,N_7601,N_7953);
nand U8691 (N_8691,N_8098,N_7944);
nand U8692 (N_8692,N_7731,N_7504);
and U8693 (N_8693,N_8096,N_8052);
and U8694 (N_8694,N_7939,N_7850);
nand U8695 (N_8695,N_7585,N_8099);
nor U8696 (N_8696,N_7853,N_7619);
nor U8697 (N_8697,N_7619,N_7505);
and U8698 (N_8698,N_7711,N_7546);
nor U8699 (N_8699,N_8071,N_7506);
xnor U8700 (N_8700,N_7626,N_7749);
nor U8701 (N_8701,N_7608,N_7897);
or U8702 (N_8702,N_7935,N_7744);
and U8703 (N_8703,N_7630,N_7641);
xnor U8704 (N_8704,N_7923,N_7652);
nand U8705 (N_8705,N_7788,N_7779);
nor U8706 (N_8706,N_7989,N_8039);
or U8707 (N_8707,N_7956,N_8008);
nand U8708 (N_8708,N_7948,N_7636);
nor U8709 (N_8709,N_7906,N_7836);
and U8710 (N_8710,N_7746,N_7769);
or U8711 (N_8711,N_7568,N_7904);
nor U8712 (N_8712,N_7745,N_7881);
or U8713 (N_8713,N_7955,N_7656);
xor U8714 (N_8714,N_7523,N_7579);
and U8715 (N_8715,N_7601,N_7705);
and U8716 (N_8716,N_7690,N_7635);
xor U8717 (N_8717,N_7676,N_7690);
and U8718 (N_8718,N_7741,N_7607);
nor U8719 (N_8719,N_8072,N_7571);
and U8720 (N_8720,N_8010,N_8048);
xor U8721 (N_8721,N_7833,N_7552);
nand U8722 (N_8722,N_8097,N_7600);
and U8723 (N_8723,N_7926,N_7595);
and U8724 (N_8724,N_8110,N_7920);
xnor U8725 (N_8725,N_7681,N_7601);
nor U8726 (N_8726,N_7777,N_8087);
nor U8727 (N_8727,N_7688,N_8003);
or U8728 (N_8728,N_7825,N_7640);
and U8729 (N_8729,N_7819,N_7862);
and U8730 (N_8730,N_8025,N_7572);
nor U8731 (N_8731,N_7933,N_8008);
and U8732 (N_8732,N_7771,N_7986);
nand U8733 (N_8733,N_7562,N_8017);
or U8734 (N_8734,N_8032,N_7641);
nand U8735 (N_8735,N_7679,N_8096);
or U8736 (N_8736,N_8122,N_7980);
or U8737 (N_8737,N_7956,N_8015);
or U8738 (N_8738,N_7876,N_7503);
xor U8739 (N_8739,N_7652,N_8105);
nand U8740 (N_8740,N_7663,N_7635);
nor U8741 (N_8741,N_7933,N_7960);
nand U8742 (N_8742,N_7832,N_7620);
and U8743 (N_8743,N_7620,N_7936);
nand U8744 (N_8744,N_7719,N_8029);
xnor U8745 (N_8745,N_7856,N_7658);
nor U8746 (N_8746,N_7703,N_7764);
or U8747 (N_8747,N_7560,N_7658);
nor U8748 (N_8748,N_7527,N_7924);
xor U8749 (N_8749,N_7771,N_7678);
nor U8750 (N_8750,N_8638,N_8126);
nand U8751 (N_8751,N_8357,N_8710);
nor U8752 (N_8752,N_8146,N_8263);
nor U8753 (N_8753,N_8628,N_8240);
or U8754 (N_8754,N_8483,N_8714);
nand U8755 (N_8755,N_8190,N_8595);
xnor U8756 (N_8756,N_8382,N_8722);
nor U8757 (N_8757,N_8518,N_8301);
and U8758 (N_8758,N_8400,N_8545);
nor U8759 (N_8759,N_8337,N_8432);
xor U8760 (N_8760,N_8627,N_8205);
and U8761 (N_8761,N_8459,N_8224);
nor U8762 (N_8762,N_8286,N_8364);
xor U8763 (N_8763,N_8642,N_8623);
or U8764 (N_8764,N_8150,N_8635);
xor U8765 (N_8765,N_8244,N_8179);
or U8766 (N_8766,N_8560,N_8725);
nand U8767 (N_8767,N_8164,N_8365);
xor U8768 (N_8768,N_8236,N_8239);
and U8769 (N_8769,N_8485,N_8167);
and U8770 (N_8770,N_8324,N_8686);
xor U8771 (N_8771,N_8130,N_8320);
and U8772 (N_8772,N_8267,N_8367);
nand U8773 (N_8773,N_8542,N_8478);
or U8774 (N_8774,N_8437,N_8407);
and U8775 (N_8775,N_8298,N_8730);
xor U8776 (N_8776,N_8335,N_8685);
and U8777 (N_8777,N_8598,N_8664);
and U8778 (N_8778,N_8720,N_8403);
and U8779 (N_8779,N_8350,N_8184);
xnor U8780 (N_8780,N_8345,N_8278);
nor U8781 (N_8781,N_8741,N_8674);
or U8782 (N_8782,N_8393,N_8472);
xor U8783 (N_8783,N_8353,N_8457);
nor U8784 (N_8784,N_8426,N_8151);
and U8785 (N_8785,N_8719,N_8712);
nand U8786 (N_8786,N_8463,N_8321);
and U8787 (N_8787,N_8625,N_8141);
or U8788 (N_8788,N_8469,N_8140);
or U8789 (N_8789,N_8160,N_8229);
nand U8790 (N_8790,N_8441,N_8523);
nor U8791 (N_8791,N_8338,N_8691);
nand U8792 (N_8792,N_8621,N_8656);
and U8793 (N_8793,N_8187,N_8166);
or U8794 (N_8794,N_8139,N_8138);
nor U8795 (N_8795,N_8667,N_8492);
xor U8796 (N_8796,N_8445,N_8423);
nand U8797 (N_8797,N_8454,N_8415);
or U8798 (N_8798,N_8653,N_8550);
xnor U8799 (N_8799,N_8270,N_8650);
and U8800 (N_8800,N_8433,N_8608);
and U8801 (N_8801,N_8732,N_8496);
and U8802 (N_8802,N_8199,N_8487);
xor U8803 (N_8803,N_8737,N_8692);
xor U8804 (N_8804,N_8438,N_8501);
xor U8805 (N_8805,N_8534,N_8145);
and U8806 (N_8806,N_8255,N_8134);
nand U8807 (N_8807,N_8616,N_8196);
or U8808 (N_8808,N_8597,N_8195);
xnor U8809 (N_8809,N_8673,N_8261);
nor U8810 (N_8810,N_8573,N_8273);
or U8811 (N_8811,N_8171,N_8589);
xnor U8812 (N_8812,N_8362,N_8183);
xor U8813 (N_8813,N_8431,N_8388);
or U8814 (N_8814,N_8617,N_8319);
nor U8815 (N_8815,N_8554,N_8652);
xor U8816 (N_8816,N_8634,N_8356);
and U8817 (N_8817,N_8210,N_8733);
and U8818 (N_8818,N_8484,N_8194);
nor U8819 (N_8819,N_8624,N_8579);
xor U8820 (N_8820,N_8551,N_8152);
or U8821 (N_8821,N_8208,N_8749);
or U8822 (N_8822,N_8748,N_8569);
nand U8823 (N_8823,N_8611,N_8746);
or U8824 (N_8824,N_8174,N_8520);
xnor U8825 (N_8825,N_8460,N_8371);
and U8826 (N_8826,N_8544,N_8693);
nand U8827 (N_8827,N_8397,N_8412);
nand U8828 (N_8828,N_8735,N_8450);
and U8829 (N_8829,N_8376,N_8473);
nand U8830 (N_8830,N_8246,N_8325);
nor U8831 (N_8831,N_8744,N_8135);
nor U8832 (N_8832,N_8275,N_8698);
xor U8833 (N_8833,N_8536,N_8574);
nand U8834 (N_8834,N_8723,N_8458);
nand U8835 (N_8835,N_8715,N_8583);
nand U8836 (N_8836,N_8348,N_8212);
nor U8837 (N_8837,N_8283,N_8696);
xor U8838 (N_8838,N_8385,N_8303);
xor U8839 (N_8839,N_8358,N_8452);
nor U8840 (N_8840,N_8227,N_8570);
nand U8841 (N_8841,N_8429,N_8386);
nor U8842 (N_8842,N_8333,N_8688);
and U8843 (N_8843,N_8577,N_8668);
nand U8844 (N_8844,N_8323,N_8464);
nor U8845 (N_8845,N_8188,N_8632);
and U8846 (N_8846,N_8169,N_8641);
nor U8847 (N_8847,N_8672,N_8713);
nor U8848 (N_8848,N_8274,N_8506);
nand U8849 (N_8849,N_8449,N_8502);
or U8850 (N_8850,N_8137,N_8253);
nor U8851 (N_8851,N_8237,N_8340);
xor U8852 (N_8852,N_8344,N_8533);
nor U8853 (N_8853,N_8479,N_8287);
and U8854 (N_8854,N_8232,N_8276);
xor U8855 (N_8855,N_8176,N_8315);
or U8856 (N_8856,N_8680,N_8192);
or U8857 (N_8857,N_8480,N_8620);
nand U8858 (N_8858,N_8299,N_8571);
and U8859 (N_8859,N_8503,N_8651);
and U8860 (N_8860,N_8327,N_8392);
or U8861 (N_8861,N_8168,N_8528);
nand U8862 (N_8862,N_8546,N_8181);
and U8863 (N_8863,N_8587,N_8659);
nor U8864 (N_8864,N_8592,N_8451);
xnor U8865 (N_8865,N_8530,N_8578);
nor U8866 (N_8866,N_8318,N_8439);
or U8867 (N_8867,N_8162,N_8509);
xor U8868 (N_8868,N_8601,N_8466);
and U8869 (N_8869,N_8567,N_8599);
nand U8870 (N_8870,N_8606,N_8552);
nand U8871 (N_8871,N_8646,N_8401);
or U8872 (N_8872,N_8684,N_8372);
nand U8873 (N_8873,N_8304,N_8510);
and U8874 (N_8874,N_8718,N_8633);
xor U8875 (N_8875,N_8500,N_8424);
or U8876 (N_8876,N_8204,N_8558);
nand U8877 (N_8877,N_8637,N_8384);
nand U8878 (N_8878,N_8127,N_8360);
nand U8879 (N_8879,N_8295,N_8526);
xor U8880 (N_8880,N_8444,N_8731);
or U8881 (N_8881,N_8476,N_8347);
xnor U8882 (N_8882,N_8497,N_8482);
and U8883 (N_8883,N_8322,N_8539);
nand U8884 (N_8884,N_8547,N_8736);
xor U8885 (N_8885,N_8655,N_8317);
nand U8886 (N_8886,N_8313,N_8368);
nand U8887 (N_8887,N_8435,N_8235);
or U8888 (N_8888,N_8387,N_8468);
or U8889 (N_8889,N_8336,N_8341);
and U8890 (N_8890,N_8610,N_8427);
nor U8891 (N_8891,N_8743,N_8156);
or U8892 (N_8892,N_8584,N_8614);
and U8893 (N_8893,N_8280,N_8515);
nand U8894 (N_8894,N_8209,N_8626);
nand U8895 (N_8895,N_8576,N_8602);
and U8896 (N_8896,N_8582,N_8186);
nand U8897 (N_8897,N_8406,N_8231);
xor U8898 (N_8898,N_8191,N_8228);
nand U8899 (N_8899,N_8475,N_8271);
and U8900 (N_8900,N_8351,N_8189);
xnor U8901 (N_8901,N_8363,N_8428);
and U8902 (N_8902,N_8580,N_8648);
xnor U8903 (N_8903,N_8588,N_8562);
and U8904 (N_8904,N_8408,N_8747);
and U8905 (N_8905,N_8241,N_8575);
and U8906 (N_8906,N_8226,N_8709);
xor U8907 (N_8907,N_8499,N_8369);
or U8908 (N_8908,N_8615,N_8540);
nor U8909 (N_8909,N_8200,N_8495);
xnor U8910 (N_8910,N_8170,N_8726);
xor U8911 (N_8911,N_8631,N_8213);
nor U8912 (N_8912,N_8417,N_8230);
or U8913 (N_8913,N_8538,N_8238);
or U8914 (N_8914,N_8354,N_8148);
and U8915 (N_8915,N_8206,N_8297);
xor U8916 (N_8916,N_8404,N_8682);
nand U8917 (N_8917,N_8339,N_8513);
and U8918 (N_8918,N_8425,N_8390);
xor U8919 (N_8919,N_8221,N_8233);
xor U8920 (N_8920,N_8294,N_8470);
xor U8921 (N_8921,N_8182,N_8416);
or U8922 (N_8922,N_8284,N_8525);
or U8923 (N_8923,N_8312,N_8249);
nor U8924 (N_8924,N_8657,N_8355);
nand U8925 (N_8925,N_8678,N_8618);
and U8926 (N_8926,N_8738,N_8374);
and U8927 (N_8927,N_8281,N_8258);
and U8928 (N_8928,N_8395,N_8512);
and U8929 (N_8929,N_8409,N_8411);
nand U8930 (N_8930,N_8332,N_8716);
and U8931 (N_8931,N_8268,N_8493);
xor U8932 (N_8932,N_8172,N_8658);
and U8933 (N_8933,N_8517,N_8504);
nand U8934 (N_8934,N_8413,N_8669);
nor U8935 (N_8935,N_8670,N_8455);
xnor U8936 (N_8936,N_8663,N_8519);
or U8937 (N_8937,N_8154,N_8153);
xor U8938 (N_8938,N_8467,N_8555);
or U8939 (N_8939,N_8277,N_8289);
nand U8940 (N_8940,N_8446,N_8234);
xor U8941 (N_8941,N_8647,N_8243);
or U8942 (N_8942,N_8342,N_8639);
or U8943 (N_8943,N_8679,N_8507);
xnor U8944 (N_8944,N_8349,N_8346);
xor U8945 (N_8945,N_8178,N_8165);
and U8946 (N_8946,N_8300,N_8256);
nor U8947 (N_8947,N_8543,N_8296);
and U8948 (N_8948,N_8700,N_8600);
nand U8949 (N_8949,N_8197,N_8640);
nand U8950 (N_8950,N_8535,N_8604);
nand U8951 (N_8951,N_8252,N_8704);
nor U8952 (N_8952,N_8133,N_8524);
nand U8953 (N_8953,N_8622,N_8155);
xnor U8954 (N_8954,N_8352,N_8381);
nor U8955 (N_8955,N_8740,N_8329);
nand U8956 (N_8956,N_8308,N_8216);
nor U8957 (N_8957,N_8453,N_8383);
and U8958 (N_8958,N_8666,N_8654);
nand U8959 (N_8959,N_8434,N_8724);
xnor U8960 (N_8960,N_8605,N_8142);
nand U8961 (N_8961,N_8566,N_8290);
and U8962 (N_8962,N_8661,N_8375);
and U8963 (N_8963,N_8465,N_8695);
and U8964 (N_8964,N_8361,N_8541);
and U8965 (N_8965,N_8702,N_8665);
nand U8966 (N_8966,N_8143,N_8591);
and U8967 (N_8967,N_8477,N_8309);
nand U8968 (N_8968,N_8185,N_8405);
xnor U8969 (N_8969,N_8527,N_8161);
xnor U8970 (N_8970,N_8711,N_8420);
nor U8971 (N_8971,N_8311,N_8343);
or U8972 (N_8972,N_8630,N_8202);
and U8973 (N_8973,N_8596,N_8548);
and U8974 (N_8974,N_8217,N_8586);
xnor U8975 (N_8975,N_8292,N_8272);
or U8976 (N_8976,N_8398,N_8291);
and U8977 (N_8977,N_8486,N_8180);
or U8978 (N_8978,N_8590,N_8328);
or U8979 (N_8979,N_8207,N_8211);
and U8980 (N_8980,N_8220,N_8373);
nand U8981 (N_8981,N_8326,N_8316);
xnor U8982 (N_8982,N_8471,N_8556);
or U8983 (N_8983,N_8742,N_8662);
nand U8984 (N_8984,N_8649,N_8334);
or U8985 (N_8985,N_8359,N_8203);
xnor U8986 (N_8986,N_8380,N_8643);
and U8987 (N_8987,N_8219,N_8144);
and U8988 (N_8988,N_8537,N_8490);
nand U8989 (N_8989,N_8251,N_8561);
or U8990 (N_8990,N_8701,N_8163);
xor U8991 (N_8991,N_8288,N_8488);
nor U8992 (N_8992,N_8708,N_8293);
nand U8993 (N_8993,N_8125,N_8491);
nand U8994 (N_8994,N_8158,N_8645);
and U8995 (N_8995,N_8694,N_8396);
and U8996 (N_8996,N_8516,N_8157);
nor U8997 (N_8997,N_8727,N_8721);
nand U8998 (N_8998,N_8609,N_8257);
or U8999 (N_8999,N_8729,N_8697);
nor U9000 (N_9000,N_8707,N_8593);
nor U9001 (N_9001,N_8690,N_8245);
nand U9002 (N_9002,N_8676,N_8739);
nor U9003 (N_9003,N_8565,N_8703);
and U9004 (N_9004,N_8254,N_8129);
or U9005 (N_9005,N_8402,N_8619);
and U9006 (N_9006,N_8607,N_8660);
xnor U9007 (N_9007,N_8644,N_8269);
and U9008 (N_9008,N_8377,N_8636);
nand U9009 (N_9009,N_8399,N_8414);
nor U9010 (N_9010,N_8394,N_8159);
xnor U9011 (N_9011,N_8734,N_8557);
nand U9012 (N_9012,N_8514,N_8136);
nor U9013 (N_9013,N_8681,N_8489);
or U9014 (N_9014,N_8314,N_8436);
xor U9015 (N_9015,N_8522,N_8306);
nor U9016 (N_9016,N_8568,N_8498);
nor U9017 (N_9017,N_8461,N_8307);
and U9018 (N_9018,N_8282,N_8262);
nor U9019 (N_9019,N_8222,N_8511);
and U9020 (N_9020,N_8706,N_8443);
nor U9021 (N_9021,N_8149,N_8147);
xor U9022 (N_9022,N_8603,N_8481);
or U9023 (N_9023,N_8175,N_8563);
nor U9024 (N_9024,N_8474,N_8302);
nor U9025 (N_9025,N_8247,N_8248);
nand U9026 (N_9026,N_8330,N_8508);
nor U9027 (N_9027,N_8687,N_8225);
or U9028 (N_9028,N_8564,N_8581);
xor U9029 (N_9029,N_8456,N_8671);
nor U9030 (N_9030,N_8585,N_8331);
and U9031 (N_9031,N_8177,N_8529);
nand U9032 (N_9032,N_8215,N_8494);
nand U9033 (N_9033,N_8173,N_8366);
nand U9034 (N_9034,N_8242,N_8447);
nor U9035 (N_9035,N_8266,N_8389);
or U9036 (N_9036,N_8370,N_8223);
nand U9037 (N_9037,N_8214,N_8430);
or U9038 (N_9038,N_8699,N_8193);
or U9039 (N_9039,N_8549,N_8559);
xnor U9040 (N_9040,N_8250,N_8305);
nand U9041 (N_9041,N_8683,N_8612);
nand U9042 (N_9042,N_8553,N_8260);
xnor U9043 (N_9043,N_8259,N_8218);
nand U9044 (N_9044,N_8572,N_8728);
nor U9045 (N_9045,N_8675,N_8705);
xnor U9046 (N_9046,N_8378,N_8717);
or U9047 (N_9047,N_8532,N_8410);
or U9048 (N_9048,N_8462,N_8279);
nand U9049 (N_9049,N_8419,N_8310);
nand U9050 (N_9050,N_8677,N_8531);
nor U9051 (N_9051,N_8440,N_8505);
or U9052 (N_9052,N_8201,N_8265);
xnor U9053 (N_9053,N_8391,N_8442);
xor U9054 (N_9054,N_8418,N_8745);
and U9055 (N_9055,N_8132,N_8448);
and U9056 (N_9056,N_8131,N_8613);
xor U9057 (N_9057,N_8379,N_8422);
xor U9058 (N_9058,N_8521,N_8128);
or U9059 (N_9059,N_8689,N_8264);
nand U9060 (N_9060,N_8198,N_8285);
nand U9061 (N_9061,N_8629,N_8421);
nor U9062 (N_9062,N_8594,N_8547);
nand U9063 (N_9063,N_8131,N_8708);
xnor U9064 (N_9064,N_8266,N_8485);
nand U9065 (N_9065,N_8277,N_8191);
nand U9066 (N_9066,N_8498,N_8245);
or U9067 (N_9067,N_8174,N_8675);
nor U9068 (N_9068,N_8663,N_8366);
nand U9069 (N_9069,N_8158,N_8467);
or U9070 (N_9070,N_8551,N_8178);
xnor U9071 (N_9071,N_8568,N_8554);
and U9072 (N_9072,N_8307,N_8252);
nand U9073 (N_9073,N_8198,N_8213);
nand U9074 (N_9074,N_8133,N_8612);
and U9075 (N_9075,N_8595,N_8334);
nor U9076 (N_9076,N_8441,N_8613);
xnor U9077 (N_9077,N_8135,N_8188);
and U9078 (N_9078,N_8188,N_8450);
xor U9079 (N_9079,N_8600,N_8388);
nor U9080 (N_9080,N_8207,N_8439);
xor U9081 (N_9081,N_8316,N_8276);
nor U9082 (N_9082,N_8660,N_8331);
nand U9083 (N_9083,N_8273,N_8407);
xor U9084 (N_9084,N_8446,N_8712);
nand U9085 (N_9085,N_8731,N_8446);
nor U9086 (N_9086,N_8145,N_8214);
and U9087 (N_9087,N_8266,N_8643);
xnor U9088 (N_9088,N_8551,N_8560);
xnor U9089 (N_9089,N_8476,N_8749);
and U9090 (N_9090,N_8385,N_8537);
or U9091 (N_9091,N_8710,N_8433);
or U9092 (N_9092,N_8312,N_8182);
or U9093 (N_9093,N_8176,N_8495);
xnor U9094 (N_9094,N_8254,N_8523);
xor U9095 (N_9095,N_8169,N_8383);
or U9096 (N_9096,N_8605,N_8525);
or U9097 (N_9097,N_8528,N_8196);
or U9098 (N_9098,N_8170,N_8153);
nand U9099 (N_9099,N_8143,N_8686);
or U9100 (N_9100,N_8477,N_8649);
and U9101 (N_9101,N_8651,N_8274);
nor U9102 (N_9102,N_8232,N_8332);
xnor U9103 (N_9103,N_8361,N_8349);
nand U9104 (N_9104,N_8203,N_8472);
and U9105 (N_9105,N_8503,N_8640);
nand U9106 (N_9106,N_8555,N_8576);
and U9107 (N_9107,N_8406,N_8441);
nor U9108 (N_9108,N_8374,N_8314);
or U9109 (N_9109,N_8648,N_8241);
xnor U9110 (N_9110,N_8293,N_8506);
nor U9111 (N_9111,N_8437,N_8226);
or U9112 (N_9112,N_8668,N_8268);
xor U9113 (N_9113,N_8220,N_8203);
xor U9114 (N_9114,N_8702,N_8366);
nor U9115 (N_9115,N_8356,N_8583);
xnor U9116 (N_9116,N_8572,N_8466);
nand U9117 (N_9117,N_8199,N_8203);
nand U9118 (N_9118,N_8335,N_8680);
xor U9119 (N_9119,N_8747,N_8660);
nor U9120 (N_9120,N_8702,N_8719);
and U9121 (N_9121,N_8485,N_8203);
and U9122 (N_9122,N_8343,N_8723);
nand U9123 (N_9123,N_8387,N_8401);
xor U9124 (N_9124,N_8698,N_8586);
xor U9125 (N_9125,N_8591,N_8513);
and U9126 (N_9126,N_8367,N_8296);
and U9127 (N_9127,N_8504,N_8721);
nand U9128 (N_9128,N_8742,N_8250);
and U9129 (N_9129,N_8399,N_8275);
xor U9130 (N_9130,N_8609,N_8313);
and U9131 (N_9131,N_8446,N_8405);
nor U9132 (N_9132,N_8289,N_8488);
xor U9133 (N_9133,N_8599,N_8161);
xor U9134 (N_9134,N_8248,N_8673);
and U9135 (N_9135,N_8733,N_8721);
and U9136 (N_9136,N_8175,N_8609);
or U9137 (N_9137,N_8158,N_8566);
and U9138 (N_9138,N_8218,N_8396);
nand U9139 (N_9139,N_8283,N_8290);
xnor U9140 (N_9140,N_8576,N_8448);
and U9141 (N_9141,N_8741,N_8438);
or U9142 (N_9142,N_8383,N_8553);
nor U9143 (N_9143,N_8544,N_8354);
nand U9144 (N_9144,N_8356,N_8216);
nand U9145 (N_9145,N_8363,N_8250);
xor U9146 (N_9146,N_8676,N_8413);
or U9147 (N_9147,N_8217,N_8383);
nand U9148 (N_9148,N_8258,N_8583);
and U9149 (N_9149,N_8353,N_8441);
xor U9150 (N_9150,N_8519,N_8200);
nand U9151 (N_9151,N_8437,N_8503);
nand U9152 (N_9152,N_8625,N_8418);
and U9153 (N_9153,N_8159,N_8645);
or U9154 (N_9154,N_8140,N_8235);
or U9155 (N_9155,N_8650,N_8475);
nand U9156 (N_9156,N_8702,N_8240);
and U9157 (N_9157,N_8507,N_8683);
xnor U9158 (N_9158,N_8343,N_8632);
or U9159 (N_9159,N_8465,N_8128);
xor U9160 (N_9160,N_8457,N_8433);
nand U9161 (N_9161,N_8498,N_8681);
nor U9162 (N_9162,N_8143,N_8543);
nor U9163 (N_9163,N_8520,N_8296);
and U9164 (N_9164,N_8263,N_8619);
and U9165 (N_9165,N_8502,N_8303);
and U9166 (N_9166,N_8265,N_8238);
and U9167 (N_9167,N_8473,N_8676);
xnor U9168 (N_9168,N_8367,N_8163);
or U9169 (N_9169,N_8146,N_8193);
nor U9170 (N_9170,N_8424,N_8490);
xor U9171 (N_9171,N_8700,N_8657);
nor U9172 (N_9172,N_8342,N_8457);
and U9173 (N_9173,N_8729,N_8468);
and U9174 (N_9174,N_8520,N_8295);
or U9175 (N_9175,N_8368,N_8746);
nor U9176 (N_9176,N_8257,N_8347);
or U9177 (N_9177,N_8586,N_8132);
nor U9178 (N_9178,N_8539,N_8320);
and U9179 (N_9179,N_8660,N_8273);
and U9180 (N_9180,N_8130,N_8499);
nor U9181 (N_9181,N_8598,N_8141);
and U9182 (N_9182,N_8684,N_8249);
nand U9183 (N_9183,N_8423,N_8394);
or U9184 (N_9184,N_8210,N_8628);
nand U9185 (N_9185,N_8271,N_8162);
or U9186 (N_9186,N_8198,N_8586);
xnor U9187 (N_9187,N_8134,N_8549);
or U9188 (N_9188,N_8186,N_8747);
or U9189 (N_9189,N_8247,N_8616);
nor U9190 (N_9190,N_8613,N_8239);
nand U9191 (N_9191,N_8660,N_8582);
nor U9192 (N_9192,N_8680,N_8570);
xnor U9193 (N_9193,N_8293,N_8358);
and U9194 (N_9194,N_8572,N_8287);
nor U9195 (N_9195,N_8733,N_8507);
or U9196 (N_9196,N_8250,N_8434);
nor U9197 (N_9197,N_8183,N_8432);
nor U9198 (N_9198,N_8211,N_8334);
xnor U9199 (N_9199,N_8237,N_8745);
or U9200 (N_9200,N_8129,N_8500);
nor U9201 (N_9201,N_8290,N_8206);
nand U9202 (N_9202,N_8332,N_8133);
xor U9203 (N_9203,N_8545,N_8338);
xnor U9204 (N_9204,N_8578,N_8711);
xnor U9205 (N_9205,N_8595,N_8376);
or U9206 (N_9206,N_8414,N_8303);
and U9207 (N_9207,N_8586,N_8134);
xor U9208 (N_9208,N_8190,N_8646);
nor U9209 (N_9209,N_8739,N_8146);
nor U9210 (N_9210,N_8322,N_8512);
or U9211 (N_9211,N_8552,N_8461);
xnor U9212 (N_9212,N_8570,N_8686);
or U9213 (N_9213,N_8468,N_8579);
and U9214 (N_9214,N_8263,N_8598);
or U9215 (N_9215,N_8583,N_8597);
xnor U9216 (N_9216,N_8187,N_8747);
or U9217 (N_9217,N_8263,N_8435);
nand U9218 (N_9218,N_8324,N_8130);
nor U9219 (N_9219,N_8153,N_8632);
and U9220 (N_9220,N_8400,N_8178);
nor U9221 (N_9221,N_8747,N_8451);
nand U9222 (N_9222,N_8614,N_8220);
xor U9223 (N_9223,N_8617,N_8692);
or U9224 (N_9224,N_8651,N_8728);
or U9225 (N_9225,N_8651,N_8613);
xor U9226 (N_9226,N_8632,N_8228);
nor U9227 (N_9227,N_8213,N_8411);
and U9228 (N_9228,N_8382,N_8468);
and U9229 (N_9229,N_8192,N_8195);
xnor U9230 (N_9230,N_8558,N_8358);
xnor U9231 (N_9231,N_8441,N_8177);
or U9232 (N_9232,N_8317,N_8479);
nand U9233 (N_9233,N_8465,N_8739);
nand U9234 (N_9234,N_8213,N_8163);
nand U9235 (N_9235,N_8529,N_8626);
xor U9236 (N_9236,N_8630,N_8352);
and U9237 (N_9237,N_8639,N_8519);
nor U9238 (N_9238,N_8309,N_8535);
nor U9239 (N_9239,N_8345,N_8555);
xnor U9240 (N_9240,N_8427,N_8225);
nand U9241 (N_9241,N_8182,N_8466);
xor U9242 (N_9242,N_8682,N_8742);
or U9243 (N_9243,N_8455,N_8233);
xnor U9244 (N_9244,N_8575,N_8685);
xor U9245 (N_9245,N_8645,N_8139);
or U9246 (N_9246,N_8266,N_8463);
or U9247 (N_9247,N_8254,N_8679);
xnor U9248 (N_9248,N_8512,N_8349);
and U9249 (N_9249,N_8574,N_8581);
nand U9250 (N_9250,N_8280,N_8420);
nand U9251 (N_9251,N_8296,N_8720);
nand U9252 (N_9252,N_8592,N_8225);
or U9253 (N_9253,N_8625,N_8556);
and U9254 (N_9254,N_8522,N_8462);
xnor U9255 (N_9255,N_8245,N_8528);
and U9256 (N_9256,N_8310,N_8349);
nor U9257 (N_9257,N_8274,N_8298);
nand U9258 (N_9258,N_8566,N_8509);
and U9259 (N_9259,N_8353,N_8268);
nand U9260 (N_9260,N_8524,N_8345);
nand U9261 (N_9261,N_8393,N_8587);
or U9262 (N_9262,N_8149,N_8169);
and U9263 (N_9263,N_8696,N_8338);
nand U9264 (N_9264,N_8264,N_8312);
or U9265 (N_9265,N_8734,N_8652);
and U9266 (N_9266,N_8703,N_8415);
xnor U9267 (N_9267,N_8176,N_8189);
or U9268 (N_9268,N_8222,N_8246);
xnor U9269 (N_9269,N_8223,N_8524);
nand U9270 (N_9270,N_8151,N_8417);
nand U9271 (N_9271,N_8261,N_8450);
nor U9272 (N_9272,N_8549,N_8357);
nor U9273 (N_9273,N_8726,N_8336);
xnor U9274 (N_9274,N_8553,N_8577);
xor U9275 (N_9275,N_8332,N_8499);
nor U9276 (N_9276,N_8653,N_8443);
xor U9277 (N_9277,N_8677,N_8273);
xnor U9278 (N_9278,N_8561,N_8270);
nand U9279 (N_9279,N_8685,N_8694);
nor U9280 (N_9280,N_8290,N_8225);
nor U9281 (N_9281,N_8694,N_8714);
and U9282 (N_9282,N_8552,N_8716);
xor U9283 (N_9283,N_8670,N_8724);
nor U9284 (N_9284,N_8321,N_8511);
xor U9285 (N_9285,N_8329,N_8519);
nor U9286 (N_9286,N_8418,N_8313);
xnor U9287 (N_9287,N_8209,N_8563);
xor U9288 (N_9288,N_8309,N_8640);
xnor U9289 (N_9289,N_8289,N_8284);
or U9290 (N_9290,N_8500,N_8607);
and U9291 (N_9291,N_8437,N_8154);
or U9292 (N_9292,N_8373,N_8566);
nor U9293 (N_9293,N_8656,N_8265);
xnor U9294 (N_9294,N_8293,N_8426);
xor U9295 (N_9295,N_8364,N_8243);
nand U9296 (N_9296,N_8658,N_8590);
nand U9297 (N_9297,N_8357,N_8476);
nor U9298 (N_9298,N_8408,N_8344);
or U9299 (N_9299,N_8700,N_8712);
nor U9300 (N_9300,N_8185,N_8346);
xor U9301 (N_9301,N_8692,N_8746);
or U9302 (N_9302,N_8147,N_8207);
xnor U9303 (N_9303,N_8716,N_8338);
nand U9304 (N_9304,N_8395,N_8716);
nor U9305 (N_9305,N_8271,N_8730);
or U9306 (N_9306,N_8185,N_8674);
xor U9307 (N_9307,N_8650,N_8654);
nor U9308 (N_9308,N_8677,N_8712);
and U9309 (N_9309,N_8209,N_8219);
nor U9310 (N_9310,N_8713,N_8589);
nor U9311 (N_9311,N_8425,N_8274);
xor U9312 (N_9312,N_8660,N_8670);
or U9313 (N_9313,N_8596,N_8299);
or U9314 (N_9314,N_8455,N_8364);
or U9315 (N_9315,N_8133,N_8684);
nor U9316 (N_9316,N_8302,N_8383);
and U9317 (N_9317,N_8195,N_8137);
nor U9318 (N_9318,N_8364,N_8299);
nand U9319 (N_9319,N_8588,N_8160);
nor U9320 (N_9320,N_8322,N_8362);
nor U9321 (N_9321,N_8176,N_8327);
nor U9322 (N_9322,N_8714,N_8130);
nor U9323 (N_9323,N_8268,N_8182);
xor U9324 (N_9324,N_8610,N_8346);
nand U9325 (N_9325,N_8293,N_8148);
or U9326 (N_9326,N_8670,N_8253);
or U9327 (N_9327,N_8347,N_8547);
nand U9328 (N_9328,N_8310,N_8245);
and U9329 (N_9329,N_8143,N_8740);
xor U9330 (N_9330,N_8409,N_8438);
nor U9331 (N_9331,N_8146,N_8469);
nor U9332 (N_9332,N_8201,N_8680);
and U9333 (N_9333,N_8467,N_8310);
or U9334 (N_9334,N_8260,N_8178);
or U9335 (N_9335,N_8499,N_8692);
xnor U9336 (N_9336,N_8389,N_8682);
or U9337 (N_9337,N_8195,N_8482);
nand U9338 (N_9338,N_8413,N_8518);
nor U9339 (N_9339,N_8251,N_8133);
and U9340 (N_9340,N_8224,N_8222);
or U9341 (N_9341,N_8393,N_8386);
and U9342 (N_9342,N_8389,N_8586);
nor U9343 (N_9343,N_8703,N_8277);
or U9344 (N_9344,N_8252,N_8136);
xor U9345 (N_9345,N_8639,N_8409);
xor U9346 (N_9346,N_8400,N_8238);
xor U9347 (N_9347,N_8425,N_8740);
xnor U9348 (N_9348,N_8288,N_8430);
or U9349 (N_9349,N_8514,N_8342);
or U9350 (N_9350,N_8431,N_8232);
nand U9351 (N_9351,N_8180,N_8396);
or U9352 (N_9352,N_8587,N_8261);
nor U9353 (N_9353,N_8580,N_8265);
xor U9354 (N_9354,N_8197,N_8538);
nand U9355 (N_9355,N_8665,N_8495);
nand U9356 (N_9356,N_8601,N_8276);
nand U9357 (N_9357,N_8453,N_8699);
nor U9358 (N_9358,N_8609,N_8606);
xor U9359 (N_9359,N_8293,N_8397);
and U9360 (N_9360,N_8261,N_8201);
nand U9361 (N_9361,N_8189,N_8620);
or U9362 (N_9362,N_8560,N_8297);
xor U9363 (N_9363,N_8704,N_8203);
xnor U9364 (N_9364,N_8607,N_8609);
nor U9365 (N_9365,N_8339,N_8310);
and U9366 (N_9366,N_8399,N_8472);
and U9367 (N_9367,N_8605,N_8655);
nor U9368 (N_9368,N_8456,N_8494);
and U9369 (N_9369,N_8430,N_8188);
nand U9370 (N_9370,N_8393,N_8242);
nor U9371 (N_9371,N_8257,N_8706);
nor U9372 (N_9372,N_8514,N_8133);
nand U9373 (N_9373,N_8702,N_8564);
xnor U9374 (N_9374,N_8148,N_8500);
or U9375 (N_9375,N_8936,N_8910);
nand U9376 (N_9376,N_9053,N_9091);
nand U9377 (N_9377,N_9116,N_8952);
nand U9378 (N_9378,N_9278,N_8822);
nand U9379 (N_9379,N_9035,N_8805);
or U9380 (N_9380,N_9284,N_9010);
and U9381 (N_9381,N_9130,N_8761);
and U9382 (N_9382,N_9121,N_8782);
nor U9383 (N_9383,N_8801,N_8827);
and U9384 (N_9384,N_8843,N_8996);
nor U9385 (N_9385,N_9242,N_9033);
nor U9386 (N_9386,N_9192,N_9215);
xor U9387 (N_9387,N_9084,N_9313);
xnor U9388 (N_9388,N_9235,N_9283);
and U9389 (N_9389,N_9339,N_8965);
or U9390 (N_9390,N_9341,N_9141);
xor U9391 (N_9391,N_9224,N_8988);
and U9392 (N_9392,N_8977,N_9005);
nand U9393 (N_9393,N_9251,N_9318);
nand U9394 (N_9394,N_9070,N_9365);
nor U9395 (N_9395,N_8750,N_8986);
or U9396 (N_9396,N_9300,N_8788);
nor U9397 (N_9397,N_8984,N_8922);
xor U9398 (N_9398,N_9234,N_9248);
xor U9399 (N_9399,N_9176,N_8828);
or U9400 (N_9400,N_8860,N_8757);
nand U9401 (N_9401,N_9250,N_9208);
and U9402 (N_9402,N_9098,N_8904);
xnor U9403 (N_9403,N_9100,N_8833);
and U9404 (N_9404,N_8769,N_9027);
nor U9405 (N_9405,N_9139,N_9069);
xnor U9406 (N_9406,N_9221,N_8932);
nand U9407 (N_9407,N_9281,N_9145);
xnor U9408 (N_9408,N_9132,N_8943);
xor U9409 (N_9409,N_8945,N_9326);
nand U9410 (N_9410,N_9324,N_8927);
xnor U9411 (N_9411,N_9340,N_9085);
nor U9412 (N_9412,N_8792,N_9233);
and U9413 (N_9413,N_9225,N_8851);
xnor U9414 (N_9414,N_8949,N_9052);
nor U9415 (N_9415,N_8781,N_9187);
nor U9416 (N_9416,N_8855,N_8919);
xnor U9417 (N_9417,N_9136,N_9325);
and U9418 (N_9418,N_9354,N_8902);
nand U9419 (N_9419,N_9018,N_8914);
nand U9420 (N_9420,N_9277,N_8925);
xor U9421 (N_9421,N_9209,N_9111);
or U9422 (N_9422,N_8989,N_8998);
and U9423 (N_9423,N_8928,N_9280);
nor U9424 (N_9424,N_8838,N_8960);
or U9425 (N_9425,N_9072,N_9152);
nor U9426 (N_9426,N_9282,N_9331);
xor U9427 (N_9427,N_9115,N_8853);
nor U9428 (N_9428,N_9368,N_8923);
xnor U9429 (N_9429,N_8979,N_8844);
and U9430 (N_9430,N_9008,N_9095);
or U9431 (N_9431,N_9007,N_8975);
nand U9432 (N_9432,N_9303,N_9046);
and U9433 (N_9433,N_9020,N_9129);
xor U9434 (N_9434,N_9106,N_9269);
and U9435 (N_9435,N_9011,N_9289);
and U9436 (N_9436,N_8888,N_9026);
or U9437 (N_9437,N_9237,N_8946);
and U9438 (N_9438,N_9147,N_9352);
and U9439 (N_9439,N_8909,N_9276);
or U9440 (N_9440,N_9193,N_9062);
and U9441 (N_9441,N_8883,N_9135);
nor U9442 (N_9442,N_9314,N_9217);
nand U9443 (N_9443,N_8839,N_8869);
and U9444 (N_9444,N_9342,N_9330);
or U9445 (N_9445,N_8818,N_8917);
nand U9446 (N_9446,N_8972,N_9185);
nor U9447 (N_9447,N_9291,N_9114);
nor U9448 (N_9448,N_8892,N_9143);
nand U9449 (N_9449,N_8825,N_8790);
xor U9450 (N_9450,N_9161,N_9370);
nand U9451 (N_9451,N_8956,N_8768);
nor U9452 (N_9452,N_9299,N_8845);
and U9453 (N_9453,N_8889,N_8884);
xor U9454 (N_9454,N_9174,N_9353);
nor U9455 (N_9455,N_9335,N_8955);
and U9456 (N_9456,N_8967,N_9261);
or U9457 (N_9457,N_8934,N_8803);
nor U9458 (N_9458,N_8906,N_9264);
xnor U9459 (N_9459,N_8879,N_8774);
nand U9460 (N_9460,N_9189,N_8873);
or U9461 (N_9461,N_9068,N_9078);
or U9462 (N_9462,N_8942,N_9076);
nor U9463 (N_9463,N_9037,N_8916);
nor U9464 (N_9464,N_8908,N_9241);
nor U9465 (N_9465,N_8793,N_8937);
or U9466 (N_9466,N_8765,N_9262);
nand U9467 (N_9467,N_8810,N_8890);
and U9468 (N_9468,N_9231,N_9265);
and U9469 (N_9469,N_9080,N_9323);
xor U9470 (N_9470,N_9322,N_9061);
xor U9471 (N_9471,N_9267,N_8852);
nor U9472 (N_9472,N_9126,N_8773);
nand U9473 (N_9473,N_8820,N_9140);
xor U9474 (N_9474,N_8775,N_8756);
and U9475 (N_9475,N_8866,N_8935);
or U9476 (N_9476,N_9124,N_9169);
xnor U9477 (N_9477,N_8870,N_9366);
nand U9478 (N_9478,N_8872,N_9023);
or U9479 (N_9479,N_9031,N_9311);
nor U9480 (N_9480,N_9109,N_8905);
nand U9481 (N_9481,N_9297,N_9119);
nor U9482 (N_9482,N_9266,N_8991);
and U9483 (N_9483,N_9239,N_8857);
and U9484 (N_9484,N_8858,N_9182);
nor U9485 (N_9485,N_9079,N_9160);
and U9486 (N_9486,N_9133,N_9216);
xnor U9487 (N_9487,N_9315,N_9252);
or U9488 (N_9488,N_9194,N_9117);
xnor U9489 (N_9489,N_8824,N_8913);
nor U9490 (N_9490,N_9017,N_8983);
xor U9491 (N_9491,N_9157,N_8950);
nor U9492 (N_9492,N_8924,N_9336);
nor U9493 (N_9493,N_9198,N_8899);
or U9494 (N_9494,N_8931,N_9083);
and U9495 (N_9495,N_9374,N_9088);
nor U9496 (N_9496,N_9190,N_8784);
nor U9497 (N_9497,N_9286,N_9293);
xnor U9498 (N_9498,N_8766,N_9044);
and U9499 (N_9499,N_8802,N_9038);
nand U9500 (N_9500,N_9155,N_9320);
or U9501 (N_9501,N_8830,N_9226);
nor U9502 (N_9502,N_8990,N_9148);
nor U9503 (N_9503,N_8835,N_8918);
and U9504 (N_9504,N_9271,N_8959);
and U9505 (N_9505,N_8846,N_9028);
or U9506 (N_9506,N_9244,N_9255);
and U9507 (N_9507,N_8886,N_8877);
nand U9508 (N_9508,N_9164,N_8817);
nand U9509 (N_9509,N_9362,N_8799);
xor U9510 (N_9510,N_9258,N_9099);
nand U9511 (N_9511,N_8981,N_9257);
nor U9512 (N_9512,N_8895,N_8786);
or U9513 (N_9513,N_8929,N_9372);
nand U9514 (N_9514,N_8896,N_9210);
nand U9515 (N_9515,N_8915,N_8856);
xnor U9516 (N_9516,N_9247,N_8785);
or U9517 (N_9517,N_9029,N_9249);
or U9518 (N_9518,N_9066,N_8767);
or U9519 (N_9519,N_8941,N_9361);
nor U9520 (N_9520,N_8814,N_9019);
nand U9521 (N_9521,N_8848,N_8821);
or U9522 (N_9522,N_8966,N_8962);
xor U9523 (N_9523,N_9165,N_8829);
nand U9524 (N_9524,N_9301,N_9230);
and U9525 (N_9525,N_9074,N_9367);
nand U9526 (N_9526,N_8787,N_9296);
xor U9527 (N_9527,N_8885,N_8847);
or U9528 (N_9528,N_8970,N_8926);
nor U9529 (N_9529,N_9067,N_9082);
nand U9530 (N_9530,N_9025,N_9347);
nand U9531 (N_9531,N_8974,N_9183);
xnor U9532 (N_9532,N_9071,N_8760);
nand U9533 (N_9533,N_9359,N_9142);
nor U9534 (N_9534,N_9039,N_9006);
nand U9535 (N_9535,N_8997,N_9127);
and U9536 (N_9536,N_9144,N_9150);
nor U9537 (N_9537,N_9309,N_8789);
or U9538 (N_9538,N_9118,N_8819);
xnor U9539 (N_9539,N_8854,N_8980);
nor U9540 (N_9540,N_8808,N_8809);
or U9541 (N_9541,N_8957,N_8815);
and U9542 (N_9542,N_9056,N_8812);
xor U9543 (N_9543,N_9223,N_8753);
xor U9544 (N_9544,N_9333,N_8794);
nor U9545 (N_9545,N_9212,N_9358);
and U9546 (N_9546,N_8944,N_9346);
nand U9547 (N_9547,N_8912,N_9290);
or U9548 (N_9548,N_8964,N_9087);
or U9549 (N_9549,N_9058,N_9338);
and U9550 (N_9550,N_8771,N_9064);
xnor U9551 (N_9551,N_9321,N_9319);
and U9552 (N_9552,N_9051,N_8796);
nor U9553 (N_9553,N_9077,N_9310);
xor U9554 (N_9554,N_9063,N_8903);
nand U9555 (N_9555,N_8762,N_9065);
and U9556 (N_9556,N_9181,N_9108);
and U9557 (N_9557,N_9360,N_9120);
and U9558 (N_9558,N_8759,N_8907);
xnor U9559 (N_9559,N_8807,N_9003);
or U9560 (N_9560,N_8841,N_8832);
or U9561 (N_9561,N_9016,N_8804);
nand U9562 (N_9562,N_9045,N_9200);
or U9563 (N_9563,N_8837,N_8995);
nor U9564 (N_9564,N_9214,N_9246);
and U9565 (N_9565,N_8940,N_8813);
xor U9566 (N_9566,N_8836,N_9171);
nor U9567 (N_9567,N_9213,N_9093);
and U9568 (N_9568,N_9287,N_9253);
xnor U9569 (N_9569,N_9199,N_8939);
nand U9570 (N_9570,N_9173,N_9256);
nor U9571 (N_9571,N_9103,N_9369);
or U9572 (N_9572,N_9306,N_8951);
and U9573 (N_9573,N_9096,N_8791);
xor U9574 (N_9574,N_9057,N_9112);
or U9575 (N_9575,N_8806,N_9328);
nand U9576 (N_9576,N_8850,N_9355);
nand U9577 (N_9577,N_8976,N_9337);
xnor U9578 (N_9578,N_9204,N_9288);
and U9579 (N_9579,N_9104,N_9364);
nand U9580 (N_9580,N_9123,N_9110);
and U9581 (N_9581,N_9081,N_8875);
xnor U9582 (N_9582,N_9030,N_8894);
nand U9583 (N_9583,N_8780,N_9363);
or U9584 (N_9584,N_9302,N_9285);
or U9585 (N_9585,N_9371,N_8987);
and U9586 (N_9586,N_9180,N_9222);
and U9587 (N_9587,N_8831,N_9050);
or U9588 (N_9588,N_9154,N_9240);
nand U9589 (N_9589,N_9205,N_9259);
nand U9590 (N_9590,N_9350,N_9015);
nand U9591 (N_9591,N_9149,N_9036);
nor U9592 (N_9592,N_8920,N_9356);
nor U9593 (N_9593,N_8994,N_8921);
nor U9594 (N_9594,N_8985,N_9166);
nor U9595 (N_9595,N_9270,N_9156);
or U9596 (N_9596,N_9263,N_8755);
and U9597 (N_9597,N_9024,N_8865);
nor U9598 (N_9598,N_8973,N_8823);
nand U9599 (N_9599,N_9307,N_9048);
nor U9600 (N_9600,N_8898,N_9305);
nand U9601 (N_9601,N_8783,N_9334);
and U9602 (N_9602,N_8758,N_9220);
xnor U9603 (N_9603,N_8953,N_9186);
nor U9604 (N_9604,N_8861,N_8897);
or U9605 (N_9605,N_8881,N_9295);
or U9606 (N_9606,N_8878,N_8840);
or U9607 (N_9607,N_8993,N_9040);
nor U9608 (N_9608,N_9268,N_8763);
nand U9609 (N_9609,N_9177,N_8752);
or U9610 (N_9610,N_9218,N_9279);
nand U9611 (N_9611,N_8864,N_8978);
nor U9612 (N_9612,N_9178,N_9043);
nand U9613 (N_9613,N_8963,N_9042);
nor U9614 (N_9614,N_8772,N_9349);
and U9615 (N_9615,N_9196,N_9245);
and U9616 (N_9616,N_9122,N_9184);
and U9617 (N_9617,N_9298,N_8862);
and U9618 (N_9618,N_8868,N_8893);
and U9619 (N_9619,N_9094,N_9107);
xor U9620 (N_9620,N_9001,N_9236);
nand U9621 (N_9621,N_9097,N_9228);
xnor U9622 (N_9622,N_8938,N_9002);
and U9623 (N_9623,N_9211,N_9332);
xnor U9624 (N_9624,N_8826,N_9312);
xnor U9625 (N_9625,N_9092,N_9075);
xor U9626 (N_9626,N_9229,N_9175);
or U9627 (N_9627,N_8954,N_9000);
nand U9628 (N_9628,N_9014,N_9275);
xor U9629 (N_9629,N_9195,N_8900);
or U9630 (N_9630,N_9012,N_8867);
and U9631 (N_9631,N_9134,N_9327);
or U9632 (N_9632,N_8834,N_9274);
or U9633 (N_9633,N_9238,N_9138);
xor U9634 (N_9634,N_8880,N_9032);
nor U9635 (N_9635,N_9034,N_9060);
and U9636 (N_9636,N_8797,N_9273);
xnor U9637 (N_9637,N_8947,N_9153);
or U9638 (N_9638,N_8958,N_9201);
xnor U9639 (N_9639,N_9089,N_9203);
and U9640 (N_9640,N_9013,N_8969);
or U9641 (N_9641,N_8842,N_9343);
nor U9642 (N_9642,N_8930,N_9049);
or U9643 (N_9643,N_8849,N_8798);
or U9644 (N_9644,N_9004,N_9022);
nand U9645 (N_9645,N_8933,N_9207);
or U9646 (N_9646,N_9373,N_9167);
or U9647 (N_9647,N_8777,N_9344);
nand U9648 (N_9648,N_9101,N_8882);
xor U9649 (N_9649,N_8982,N_9158);
or U9650 (N_9650,N_8971,N_9073);
nand U9651 (N_9651,N_8776,N_9170);
or U9652 (N_9652,N_8859,N_9054);
and U9653 (N_9653,N_9168,N_9009);
xor U9654 (N_9654,N_8901,N_8754);
and U9655 (N_9655,N_9086,N_9151);
nand U9656 (N_9656,N_9260,N_9125);
nor U9657 (N_9657,N_9172,N_8764);
nand U9658 (N_9658,N_9041,N_8816);
nand U9659 (N_9659,N_9090,N_8770);
xnor U9660 (N_9660,N_8779,N_9047);
nand U9661 (N_9661,N_9159,N_9219);
xnor U9662 (N_9662,N_9292,N_9113);
nor U9663 (N_9663,N_9317,N_8999);
xnor U9664 (N_9664,N_9131,N_9055);
nor U9665 (N_9665,N_8911,N_8992);
nand U9666 (N_9666,N_8871,N_8778);
nor U9667 (N_9667,N_9316,N_9146);
xnor U9668 (N_9668,N_9059,N_9272);
and U9669 (N_9669,N_9021,N_9163);
nand U9670 (N_9670,N_9102,N_8863);
xnor U9671 (N_9671,N_9254,N_8795);
and U9672 (N_9672,N_8811,N_9232);
or U9673 (N_9673,N_8891,N_9329);
or U9674 (N_9674,N_8887,N_9188);
nand U9675 (N_9675,N_8874,N_9294);
or U9676 (N_9676,N_9304,N_9308);
nand U9677 (N_9677,N_9345,N_8800);
xnor U9678 (N_9678,N_9351,N_8968);
nor U9679 (N_9679,N_9348,N_9105);
or U9680 (N_9680,N_8751,N_9197);
nor U9681 (N_9681,N_9227,N_9137);
and U9682 (N_9682,N_8948,N_9191);
nor U9683 (N_9683,N_8876,N_9357);
nand U9684 (N_9684,N_8961,N_9202);
and U9685 (N_9685,N_9162,N_9179);
nor U9686 (N_9686,N_9206,N_9128);
xor U9687 (N_9687,N_9243,N_8751);
or U9688 (N_9688,N_8825,N_9330);
nor U9689 (N_9689,N_8877,N_9341);
nand U9690 (N_9690,N_9109,N_9303);
nand U9691 (N_9691,N_9087,N_9203);
nor U9692 (N_9692,N_9054,N_9207);
xnor U9693 (N_9693,N_8829,N_9256);
nor U9694 (N_9694,N_9322,N_8864);
or U9695 (N_9695,N_9079,N_9292);
or U9696 (N_9696,N_8805,N_9115);
or U9697 (N_9697,N_8929,N_9075);
xnor U9698 (N_9698,N_9047,N_9315);
xor U9699 (N_9699,N_8904,N_9021);
or U9700 (N_9700,N_8763,N_8805);
and U9701 (N_9701,N_9207,N_9265);
xor U9702 (N_9702,N_8912,N_9094);
xnor U9703 (N_9703,N_8915,N_9147);
xor U9704 (N_9704,N_8931,N_9357);
and U9705 (N_9705,N_9278,N_9060);
or U9706 (N_9706,N_9115,N_9267);
or U9707 (N_9707,N_9366,N_9329);
or U9708 (N_9708,N_8929,N_9265);
or U9709 (N_9709,N_9299,N_8900);
nand U9710 (N_9710,N_8879,N_9176);
and U9711 (N_9711,N_9177,N_8801);
xnor U9712 (N_9712,N_8977,N_9076);
nor U9713 (N_9713,N_9102,N_8894);
nor U9714 (N_9714,N_8801,N_9211);
xnor U9715 (N_9715,N_9347,N_9326);
nor U9716 (N_9716,N_9116,N_9099);
nand U9717 (N_9717,N_9188,N_9165);
or U9718 (N_9718,N_9315,N_8913);
or U9719 (N_9719,N_9120,N_9242);
and U9720 (N_9720,N_9259,N_9059);
nor U9721 (N_9721,N_9288,N_8822);
nor U9722 (N_9722,N_9316,N_9307);
or U9723 (N_9723,N_9028,N_8935);
and U9724 (N_9724,N_9280,N_8988);
or U9725 (N_9725,N_9196,N_9097);
and U9726 (N_9726,N_9115,N_8943);
and U9727 (N_9727,N_8799,N_8915);
xnor U9728 (N_9728,N_9287,N_9348);
or U9729 (N_9729,N_9247,N_9312);
nand U9730 (N_9730,N_9060,N_8789);
or U9731 (N_9731,N_8948,N_8782);
nor U9732 (N_9732,N_9226,N_8868);
nand U9733 (N_9733,N_8759,N_9341);
xnor U9734 (N_9734,N_9283,N_8820);
or U9735 (N_9735,N_9146,N_9330);
nor U9736 (N_9736,N_9133,N_9319);
and U9737 (N_9737,N_9092,N_9232);
nand U9738 (N_9738,N_9215,N_8972);
or U9739 (N_9739,N_9298,N_9289);
or U9740 (N_9740,N_9094,N_9250);
nand U9741 (N_9741,N_8962,N_8945);
xor U9742 (N_9742,N_8774,N_9154);
or U9743 (N_9743,N_8762,N_9250);
xor U9744 (N_9744,N_8859,N_9374);
and U9745 (N_9745,N_9041,N_8761);
nor U9746 (N_9746,N_9158,N_8863);
xnor U9747 (N_9747,N_9017,N_9337);
nand U9748 (N_9748,N_8911,N_9072);
nor U9749 (N_9749,N_8971,N_8798);
xnor U9750 (N_9750,N_8969,N_9258);
nand U9751 (N_9751,N_9363,N_8771);
xnor U9752 (N_9752,N_9007,N_9259);
xor U9753 (N_9753,N_8915,N_8890);
nand U9754 (N_9754,N_8935,N_9009);
xor U9755 (N_9755,N_8848,N_8805);
nor U9756 (N_9756,N_9261,N_8916);
nand U9757 (N_9757,N_9122,N_9076);
xor U9758 (N_9758,N_9083,N_9119);
nand U9759 (N_9759,N_9089,N_8956);
xor U9760 (N_9760,N_9141,N_8875);
or U9761 (N_9761,N_8976,N_8849);
nand U9762 (N_9762,N_8895,N_8989);
or U9763 (N_9763,N_9305,N_8894);
nand U9764 (N_9764,N_8949,N_9261);
xor U9765 (N_9765,N_9240,N_9188);
xnor U9766 (N_9766,N_8844,N_8939);
xor U9767 (N_9767,N_9186,N_9255);
nand U9768 (N_9768,N_9241,N_9090);
and U9769 (N_9769,N_9246,N_9147);
nor U9770 (N_9770,N_9308,N_9250);
xor U9771 (N_9771,N_9260,N_9006);
xnor U9772 (N_9772,N_9055,N_8920);
or U9773 (N_9773,N_9143,N_9169);
nand U9774 (N_9774,N_9203,N_9000);
nor U9775 (N_9775,N_8779,N_8804);
nand U9776 (N_9776,N_8809,N_9108);
xnor U9777 (N_9777,N_8946,N_8893);
and U9778 (N_9778,N_9331,N_9018);
and U9779 (N_9779,N_9260,N_9033);
and U9780 (N_9780,N_9223,N_9256);
nor U9781 (N_9781,N_9332,N_9221);
nand U9782 (N_9782,N_8832,N_9286);
nand U9783 (N_9783,N_9333,N_9352);
nand U9784 (N_9784,N_9266,N_9029);
or U9785 (N_9785,N_8832,N_8992);
xor U9786 (N_9786,N_9005,N_8782);
nand U9787 (N_9787,N_8792,N_9004);
nand U9788 (N_9788,N_8927,N_9197);
or U9789 (N_9789,N_8829,N_9065);
or U9790 (N_9790,N_9099,N_9035);
nand U9791 (N_9791,N_8931,N_8771);
nand U9792 (N_9792,N_8815,N_9314);
nand U9793 (N_9793,N_8854,N_8934);
or U9794 (N_9794,N_8808,N_9352);
and U9795 (N_9795,N_8792,N_9121);
and U9796 (N_9796,N_8801,N_8892);
or U9797 (N_9797,N_8951,N_8844);
xnor U9798 (N_9798,N_8930,N_9281);
or U9799 (N_9799,N_9034,N_9265);
xnor U9800 (N_9800,N_9183,N_8904);
nor U9801 (N_9801,N_8919,N_9205);
nand U9802 (N_9802,N_9200,N_9254);
nor U9803 (N_9803,N_9253,N_9013);
nor U9804 (N_9804,N_9362,N_8879);
xor U9805 (N_9805,N_9204,N_8778);
or U9806 (N_9806,N_8808,N_9261);
nand U9807 (N_9807,N_8808,N_9229);
nand U9808 (N_9808,N_9265,N_8899);
or U9809 (N_9809,N_9150,N_9218);
or U9810 (N_9810,N_9343,N_8897);
nand U9811 (N_9811,N_8924,N_9043);
and U9812 (N_9812,N_9043,N_8996);
xnor U9813 (N_9813,N_8981,N_9093);
or U9814 (N_9814,N_9142,N_9067);
xor U9815 (N_9815,N_8995,N_8829);
nand U9816 (N_9816,N_9214,N_9241);
nand U9817 (N_9817,N_9043,N_9121);
or U9818 (N_9818,N_9296,N_8878);
xnor U9819 (N_9819,N_8927,N_8757);
and U9820 (N_9820,N_9140,N_8939);
xnor U9821 (N_9821,N_8987,N_9181);
nand U9822 (N_9822,N_9212,N_9063);
nand U9823 (N_9823,N_8796,N_8809);
nand U9824 (N_9824,N_8910,N_8947);
or U9825 (N_9825,N_9248,N_9138);
nor U9826 (N_9826,N_8945,N_9026);
nand U9827 (N_9827,N_9074,N_9163);
xor U9828 (N_9828,N_8899,N_8753);
and U9829 (N_9829,N_9205,N_8755);
or U9830 (N_9830,N_9280,N_9272);
nand U9831 (N_9831,N_9274,N_8874);
xor U9832 (N_9832,N_9098,N_8805);
nor U9833 (N_9833,N_8752,N_9171);
nand U9834 (N_9834,N_8867,N_9358);
nand U9835 (N_9835,N_8974,N_9301);
nor U9836 (N_9836,N_8952,N_9184);
nand U9837 (N_9837,N_9155,N_8939);
xor U9838 (N_9838,N_8867,N_9037);
or U9839 (N_9839,N_9179,N_8928);
or U9840 (N_9840,N_9021,N_8876);
nand U9841 (N_9841,N_9275,N_9120);
nand U9842 (N_9842,N_9102,N_8971);
nand U9843 (N_9843,N_9188,N_8787);
nor U9844 (N_9844,N_9177,N_9342);
nand U9845 (N_9845,N_9039,N_9022);
or U9846 (N_9846,N_8973,N_9245);
nor U9847 (N_9847,N_9363,N_8767);
or U9848 (N_9848,N_9171,N_8767);
nor U9849 (N_9849,N_9247,N_8871);
nor U9850 (N_9850,N_8896,N_9038);
xnor U9851 (N_9851,N_8865,N_9291);
xnor U9852 (N_9852,N_9326,N_9355);
or U9853 (N_9853,N_9194,N_8926);
nor U9854 (N_9854,N_8816,N_8837);
or U9855 (N_9855,N_8910,N_8956);
nand U9856 (N_9856,N_8904,N_8769);
and U9857 (N_9857,N_8821,N_9259);
or U9858 (N_9858,N_8831,N_9233);
nand U9859 (N_9859,N_9262,N_8986);
nor U9860 (N_9860,N_9031,N_8807);
or U9861 (N_9861,N_9367,N_9164);
xor U9862 (N_9862,N_9225,N_9197);
and U9863 (N_9863,N_9234,N_9330);
xnor U9864 (N_9864,N_8907,N_9279);
and U9865 (N_9865,N_9310,N_9165);
nand U9866 (N_9866,N_8781,N_9108);
xor U9867 (N_9867,N_9250,N_8760);
nand U9868 (N_9868,N_9225,N_8845);
xnor U9869 (N_9869,N_9326,N_8934);
and U9870 (N_9870,N_8884,N_9078);
and U9871 (N_9871,N_9036,N_9340);
xor U9872 (N_9872,N_9105,N_9064);
nor U9873 (N_9873,N_8876,N_8909);
or U9874 (N_9874,N_9001,N_9164);
and U9875 (N_9875,N_9230,N_8752);
nand U9876 (N_9876,N_9109,N_8947);
nand U9877 (N_9877,N_9319,N_8757);
xnor U9878 (N_9878,N_9188,N_9081);
nand U9879 (N_9879,N_9131,N_8752);
nor U9880 (N_9880,N_8795,N_9357);
or U9881 (N_9881,N_9361,N_8836);
and U9882 (N_9882,N_8777,N_9171);
or U9883 (N_9883,N_8972,N_9140);
and U9884 (N_9884,N_8953,N_9090);
nor U9885 (N_9885,N_9194,N_9323);
xnor U9886 (N_9886,N_9340,N_8971);
nand U9887 (N_9887,N_9017,N_9003);
nand U9888 (N_9888,N_9327,N_9359);
xnor U9889 (N_9889,N_8917,N_9024);
or U9890 (N_9890,N_8991,N_8752);
nand U9891 (N_9891,N_8857,N_9086);
xnor U9892 (N_9892,N_8799,N_8787);
nand U9893 (N_9893,N_9098,N_9346);
or U9894 (N_9894,N_9070,N_9242);
nor U9895 (N_9895,N_9257,N_9260);
nor U9896 (N_9896,N_8753,N_8809);
nand U9897 (N_9897,N_9272,N_9105);
and U9898 (N_9898,N_9056,N_9194);
nand U9899 (N_9899,N_9224,N_8892);
or U9900 (N_9900,N_9292,N_9160);
or U9901 (N_9901,N_9017,N_9011);
or U9902 (N_9902,N_9178,N_9172);
and U9903 (N_9903,N_8878,N_8872);
and U9904 (N_9904,N_9331,N_9152);
nand U9905 (N_9905,N_8907,N_9289);
and U9906 (N_9906,N_9106,N_9340);
nor U9907 (N_9907,N_8858,N_9314);
or U9908 (N_9908,N_8915,N_9364);
xnor U9909 (N_9909,N_8766,N_8886);
or U9910 (N_9910,N_9310,N_8786);
nand U9911 (N_9911,N_8881,N_9239);
xnor U9912 (N_9912,N_9187,N_9335);
and U9913 (N_9913,N_9017,N_8945);
nor U9914 (N_9914,N_9127,N_9059);
nand U9915 (N_9915,N_9185,N_9336);
nor U9916 (N_9916,N_8754,N_9342);
nor U9917 (N_9917,N_9063,N_9115);
nand U9918 (N_9918,N_8796,N_8758);
xor U9919 (N_9919,N_9310,N_9212);
nor U9920 (N_9920,N_8805,N_9066);
nand U9921 (N_9921,N_9052,N_8802);
nand U9922 (N_9922,N_8830,N_9107);
or U9923 (N_9923,N_9194,N_8939);
nor U9924 (N_9924,N_8764,N_8914);
and U9925 (N_9925,N_9154,N_9205);
or U9926 (N_9926,N_8868,N_8826);
xor U9927 (N_9927,N_9259,N_9364);
xor U9928 (N_9928,N_8852,N_9143);
nor U9929 (N_9929,N_9368,N_8827);
nand U9930 (N_9930,N_9165,N_9073);
and U9931 (N_9931,N_8958,N_8909);
and U9932 (N_9932,N_8809,N_8896);
or U9933 (N_9933,N_8816,N_9185);
or U9934 (N_9934,N_9253,N_9208);
nand U9935 (N_9935,N_8891,N_8986);
nand U9936 (N_9936,N_8911,N_8858);
and U9937 (N_9937,N_9370,N_8786);
and U9938 (N_9938,N_8971,N_8810);
or U9939 (N_9939,N_9330,N_9109);
nor U9940 (N_9940,N_9137,N_9150);
xnor U9941 (N_9941,N_8759,N_8936);
nand U9942 (N_9942,N_9061,N_9372);
or U9943 (N_9943,N_9059,N_8935);
or U9944 (N_9944,N_8993,N_8948);
nor U9945 (N_9945,N_8975,N_8837);
xnor U9946 (N_9946,N_8847,N_9133);
or U9947 (N_9947,N_8969,N_9289);
and U9948 (N_9948,N_9303,N_9250);
nand U9949 (N_9949,N_9351,N_9353);
or U9950 (N_9950,N_8935,N_8843);
nor U9951 (N_9951,N_8814,N_8917);
nor U9952 (N_9952,N_8809,N_9140);
xor U9953 (N_9953,N_8973,N_9144);
nand U9954 (N_9954,N_8839,N_9179);
nor U9955 (N_9955,N_9086,N_9303);
nand U9956 (N_9956,N_8926,N_9057);
xnor U9957 (N_9957,N_8987,N_9112);
nand U9958 (N_9958,N_9131,N_9244);
nor U9959 (N_9959,N_8842,N_8775);
or U9960 (N_9960,N_9335,N_8948);
xnor U9961 (N_9961,N_9209,N_8834);
nor U9962 (N_9962,N_9052,N_9108);
nor U9963 (N_9963,N_9295,N_8873);
nor U9964 (N_9964,N_9150,N_9175);
nand U9965 (N_9965,N_8886,N_9208);
nand U9966 (N_9966,N_9300,N_9218);
and U9967 (N_9967,N_8766,N_9013);
xor U9968 (N_9968,N_8753,N_8978);
nand U9969 (N_9969,N_9365,N_9164);
nor U9970 (N_9970,N_8976,N_8836);
and U9971 (N_9971,N_9226,N_8952);
nor U9972 (N_9972,N_9082,N_8871);
xor U9973 (N_9973,N_9002,N_8911);
or U9974 (N_9974,N_9033,N_9172);
nor U9975 (N_9975,N_9149,N_9257);
or U9976 (N_9976,N_8799,N_9373);
nor U9977 (N_9977,N_8866,N_8788);
or U9978 (N_9978,N_9250,N_9062);
xnor U9979 (N_9979,N_9216,N_9079);
nor U9980 (N_9980,N_9079,N_9319);
xnor U9981 (N_9981,N_9182,N_8945);
nand U9982 (N_9982,N_8876,N_9071);
xor U9983 (N_9983,N_9080,N_8936);
xor U9984 (N_9984,N_9150,N_9230);
xnor U9985 (N_9985,N_9343,N_9359);
and U9986 (N_9986,N_8762,N_9358);
nor U9987 (N_9987,N_9142,N_9208);
nor U9988 (N_9988,N_9120,N_8881);
xnor U9989 (N_9989,N_9317,N_9100);
or U9990 (N_9990,N_9357,N_8838);
xor U9991 (N_9991,N_9216,N_8845);
nor U9992 (N_9992,N_9143,N_8939);
nor U9993 (N_9993,N_8798,N_9235);
or U9994 (N_9994,N_8895,N_8899);
xnor U9995 (N_9995,N_8909,N_8881);
nand U9996 (N_9996,N_9133,N_9270);
or U9997 (N_9997,N_8960,N_9055);
and U9998 (N_9998,N_9372,N_9136);
and U9999 (N_9999,N_9237,N_9196);
or U10000 (N_10000,N_9965,N_9562);
nor U10001 (N_10001,N_9925,N_9733);
xor U10002 (N_10002,N_9608,N_9420);
nand U10003 (N_10003,N_9854,N_9823);
xor U10004 (N_10004,N_9503,N_9787);
nand U10005 (N_10005,N_9446,N_9576);
nand U10006 (N_10006,N_9809,N_9388);
nor U10007 (N_10007,N_9996,N_9794);
and U10008 (N_10008,N_9881,N_9546);
and U10009 (N_10009,N_9430,N_9805);
or U10010 (N_10010,N_9395,N_9880);
nor U10011 (N_10011,N_9398,N_9651);
or U10012 (N_10012,N_9400,N_9511);
nor U10013 (N_10013,N_9834,N_9859);
xnor U10014 (N_10014,N_9640,N_9720);
nand U10015 (N_10015,N_9500,N_9605);
or U10016 (N_10016,N_9862,N_9396);
nand U10017 (N_10017,N_9948,N_9833);
nand U10018 (N_10018,N_9957,N_9840);
nor U10019 (N_10019,N_9556,N_9930);
nand U10020 (N_10020,N_9981,N_9634);
xnor U10021 (N_10021,N_9413,N_9879);
nor U10022 (N_10022,N_9941,N_9693);
or U10023 (N_10023,N_9803,N_9642);
or U10024 (N_10024,N_9839,N_9628);
nor U10025 (N_10025,N_9766,N_9582);
or U10026 (N_10026,N_9997,N_9580);
or U10027 (N_10027,N_9968,N_9403);
xor U10028 (N_10028,N_9416,N_9598);
or U10029 (N_10029,N_9801,N_9380);
or U10030 (N_10030,N_9568,N_9650);
xor U10031 (N_10031,N_9566,N_9744);
or U10032 (N_10032,N_9414,N_9783);
xor U10033 (N_10033,N_9501,N_9928);
nor U10034 (N_10034,N_9807,N_9635);
nor U10035 (N_10035,N_9687,N_9603);
xnor U10036 (N_10036,N_9892,N_9683);
or U10037 (N_10037,N_9713,N_9481);
nand U10038 (N_10038,N_9726,N_9982);
and U10039 (N_10039,N_9675,N_9953);
or U10040 (N_10040,N_9999,N_9520);
nor U10041 (N_10041,N_9735,N_9983);
and U10042 (N_10042,N_9757,N_9742);
or U10043 (N_10043,N_9410,N_9577);
xnor U10044 (N_10044,N_9732,N_9902);
and U10045 (N_10045,N_9819,N_9602);
nor U10046 (N_10046,N_9775,N_9728);
or U10047 (N_10047,N_9377,N_9922);
nand U10048 (N_10048,N_9616,N_9774);
nand U10049 (N_10049,N_9574,N_9575);
and U10050 (N_10050,N_9518,N_9569);
and U10051 (N_10051,N_9588,N_9644);
xnor U10052 (N_10052,N_9561,N_9769);
or U10053 (N_10053,N_9952,N_9937);
and U10054 (N_10054,N_9549,N_9853);
nand U10055 (N_10055,N_9724,N_9496);
nand U10056 (N_10056,N_9986,N_9464);
xor U10057 (N_10057,N_9876,N_9466);
nand U10058 (N_10058,N_9652,N_9802);
or U10059 (N_10059,N_9459,N_9714);
and U10060 (N_10060,N_9495,N_9754);
nor U10061 (N_10061,N_9516,N_9538);
nor U10062 (N_10062,N_9393,N_9830);
nor U10063 (N_10063,N_9878,N_9895);
and U10064 (N_10064,N_9612,N_9804);
and U10065 (N_10065,N_9731,N_9931);
nor U10066 (N_10066,N_9792,N_9920);
or U10067 (N_10067,N_9747,N_9405);
xor U10068 (N_10068,N_9858,N_9715);
or U10069 (N_10069,N_9970,N_9703);
nand U10070 (N_10070,N_9739,N_9475);
nand U10071 (N_10071,N_9991,N_9601);
xnor U10072 (N_10072,N_9385,N_9445);
or U10073 (N_10073,N_9631,N_9505);
nor U10074 (N_10074,N_9844,N_9647);
nand U10075 (N_10075,N_9978,N_9686);
nor U10076 (N_10076,N_9589,N_9412);
and U10077 (N_10077,N_9725,N_9417);
or U10078 (N_10078,N_9756,N_9710);
nand U10079 (N_10079,N_9552,N_9852);
or U10080 (N_10080,N_9509,N_9523);
xor U10081 (N_10081,N_9818,N_9889);
nor U10082 (N_10082,N_9663,N_9531);
nor U10083 (N_10083,N_9565,N_9474);
and U10084 (N_10084,N_9623,N_9606);
xnor U10085 (N_10085,N_9404,N_9989);
and U10086 (N_10086,N_9846,N_9402);
and U10087 (N_10087,N_9488,N_9617);
xnor U10088 (N_10088,N_9419,N_9870);
and U10089 (N_10089,N_9966,N_9842);
nor U10090 (N_10090,N_9951,N_9528);
or U10091 (N_10091,N_9706,N_9873);
nor U10092 (N_10092,N_9450,N_9884);
or U10093 (N_10093,N_9944,N_9692);
xor U10094 (N_10094,N_9591,N_9529);
and U10095 (N_10095,N_9590,N_9824);
and U10096 (N_10096,N_9421,N_9378);
xnor U10097 (N_10097,N_9704,N_9699);
or U10098 (N_10098,N_9537,N_9613);
and U10099 (N_10099,N_9648,N_9843);
or U10100 (N_10100,N_9610,N_9817);
xnor U10101 (N_10101,N_9691,N_9776);
nor U10102 (N_10102,N_9814,N_9670);
nand U10103 (N_10103,N_9765,N_9424);
and U10104 (N_10104,N_9806,N_9502);
nor U10105 (N_10105,N_9442,N_9738);
xnor U10106 (N_10106,N_9826,N_9749);
xnor U10107 (N_10107,N_9780,N_9901);
nor U10108 (N_10108,N_9427,N_9479);
nor U10109 (N_10109,N_9536,N_9657);
or U10110 (N_10110,N_9519,N_9915);
nand U10111 (N_10111,N_9596,N_9480);
and U10112 (N_10112,N_9960,N_9764);
or U10113 (N_10113,N_9639,N_9964);
nand U10114 (N_10114,N_9468,N_9871);
xnor U10115 (N_10115,N_9521,N_9390);
or U10116 (N_10116,N_9541,N_9909);
nand U10117 (N_10117,N_9543,N_9719);
xnor U10118 (N_10118,N_9690,N_9389);
nor U10119 (N_10119,N_9907,N_9768);
or U10120 (N_10120,N_9912,N_9782);
and U10121 (N_10121,N_9674,N_9583);
and U10122 (N_10122,N_9935,N_9578);
xnor U10123 (N_10123,N_9685,N_9615);
nor U10124 (N_10124,N_9487,N_9882);
xnor U10125 (N_10125,N_9790,N_9632);
or U10126 (N_10126,N_9581,N_9856);
nor U10127 (N_10127,N_9600,N_9433);
and U10128 (N_10128,N_9471,N_9770);
xnor U10129 (N_10129,N_9810,N_9545);
xor U10130 (N_10130,N_9483,N_9553);
nor U10131 (N_10131,N_9406,N_9837);
and U10132 (N_10132,N_9684,N_9939);
nand U10133 (N_10133,N_9698,N_9513);
xnor U10134 (N_10134,N_9493,N_9701);
nand U10135 (N_10135,N_9694,N_9867);
or U10136 (N_10136,N_9463,N_9857);
or U10137 (N_10137,N_9666,N_9740);
and U10138 (N_10138,N_9485,N_9458);
and U10139 (N_10139,N_9932,N_9727);
or U10140 (N_10140,N_9750,N_9671);
or U10141 (N_10141,N_9921,N_9849);
or U10142 (N_10142,N_9426,N_9812);
and U10143 (N_10143,N_9383,N_9387);
nand U10144 (N_10144,N_9494,N_9702);
nand U10145 (N_10145,N_9517,N_9800);
and U10146 (N_10146,N_9891,N_9872);
nand U10147 (N_10147,N_9753,N_9641);
xnor U10148 (N_10148,N_9990,N_9579);
or U10149 (N_10149,N_9914,N_9447);
nor U10150 (N_10150,N_9936,N_9751);
nand U10151 (N_10151,N_9927,N_9435);
or U10152 (N_10152,N_9508,N_9415);
nand U10153 (N_10153,N_9969,N_9918);
or U10154 (N_10154,N_9938,N_9898);
or U10155 (N_10155,N_9993,N_9897);
and U10156 (N_10156,N_9662,N_9636);
or U10157 (N_10157,N_9504,N_9729);
nor U10158 (N_10158,N_9795,N_9955);
nand U10159 (N_10159,N_9786,N_9877);
nand U10160 (N_10160,N_9465,N_9900);
and U10161 (N_10161,N_9886,N_9919);
or U10162 (N_10162,N_9697,N_9721);
nand U10163 (N_10163,N_9676,N_9791);
xor U10164 (N_10164,N_9593,N_9954);
or U10165 (N_10165,N_9525,N_9988);
nor U10166 (N_10166,N_9376,N_9476);
or U10167 (N_10167,N_9530,N_9796);
nand U10168 (N_10168,N_9894,N_9618);
and U10169 (N_10169,N_9910,N_9599);
nand U10170 (N_10170,N_9484,N_9865);
nand U10171 (N_10171,N_9443,N_9512);
or U10172 (N_10172,N_9736,N_9841);
xor U10173 (N_10173,N_9680,N_9571);
nand U10174 (N_10174,N_9933,N_9831);
and U10175 (N_10175,N_9607,N_9779);
nand U10176 (N_10176,N_9646,N_9718);
and U10177 (N_10177,N_9401,N_9436);
nand U10178 (N_10178,N_9974,N_9498);
and U10179 (N_10179,N_9429,N_9557);
nand U10180 (N_10180,N_9861,N_9994);
nand U10181 (N_10181,N_9542,N_9559);
and U10182 (N_10182,N_9869,N_9967);
nand U10183 (N_10183,N_9755,N_9899);
and U10184 (N_10184,N_9864,N_9486);
xnor U10185 (N_10185,N_9949,N_9832);
xor U10186 (N_10186,N_9437,N_9460);
or U10187 (N_10187,N_9822,N_9630);
or U10188 (N_10188,N_9962,N_9771);
xnor U10189 (N_10189,N_9825,N_9958);
or U10190 (N_10190,N_9668,N_9422);
nor U10191 (N_10191,N_9375,N_9903);
and U10192 (N_10192,N_9813,N_9527);
xor U10193 (N_10193,N_9924,N_9976);
and U10194 (N_10194,N_9611,N_9828);
nor U10195 (N_10195,N_9868,N_9679);
xor U10196 (N_10196,N_9441,N_9708);
or U10197 (N_10197,N_9449,N_9712);
nor U10198 (N_10198,N_9885,N_9929);
nor U10199 (N_10199,N_9497,N_9626);
xor U10200 (N_10200,N_9391,N_9655);
and U10201 (N_10201,N_9461,N_9984);
and U10202 (N_10202,N_9619,N_9992);
or U10203 (N_10203,N_9477,N_9798);
and U10204 (N_10204,N_9956,N_9746);
nand U10205 (N_10205,N_9829,N_9482);
xnor U10206 (N_10206,N_9547,N_9643);
xor U10207 (N_10207,N_9673,N_9773);
nand U10208 (N_10208,N_9785,N_9473);
and U10209 (N_10209,N_9656,N_9467);
nand U10210 (N_10210,N_9908,N_9911);
and U10211 (N_10211,N_9896,N_9510);
nor U10212 (N_10212,N_9621,N_9462);
nand U10213 (N_10213,N_9609,N_9987);
nand U10214 (N_10214,N_9689,N_9455);
and U10215 (N_10215,N_9407,N_9638);
nand U10216 (N_10216,N_9558,N_9515);
and U10217 (N_10217,N_9478,N_9851);
and U10218 (N_10218,N_9863,N_9977);
xor U10219 (N_10219,N_9883,N_9848);
nor U10220 (N_10220,N_9550,N_9847);
nand U10221 (N_10221,N_9836,N_9444);
xnor U10222 (N_10222,N_9816,N_9972);
xor U10223 (N_10223,N_9532,N_9860);
or U10224 (N_10224,N_9408,N_9597);
xor U10225 (N_10225,N_9760,N_9758);
nor U10226 (N_10226,N_9397,N_9423);
or U10227 (N_10227,N_9709,N_9448);
nor U10228 (N_10228,N_9716,N_9425);
xnor U10229 (N_10229,N_9431,N_9667);
and U10230 (N_10230,N_9379,N_9490);
and U10231 (N_10231,N_9835,N_9548);
or U10232 (N_10232,N_9661,N_9917);
and U10233 (N_10233,N_9409,N_9434);
nand U10234 (N_10234,N_9700,N_9658);
xor U10235 (N_10235,N_9620,N_9604);
or U10236 (N_10236,N_9625,N_9454);
nor U10237 (N_10237,N_9722,N_9524);
xor U10238 (N_10238,N_9456,N_9554);
xor U10239 (N_10239,N_9586,N_9781);
nor U10240 (N_10240,N_9411,N_9797);
nor U10241 (N_10241,N_9905,N_9678);
nor U10242 (N_10242,N_9737,N_9560);
xnor U10243 (N_10243,N_9637,N_9633);
nor U10244 (N_10244,N_9904,N_9975);
and U10245 (N_10245,N_9752,N_9767);
or U10246 (N_10246,N_9855,N_9734);
xor U10247 (N_10247,N_9916,N_9695);
nand U10248 (N_10248,N_9971,N_9555);
or U10249 (N_10249,N_9492,N_9961);
xor U10250 (N_10250,N_9945,N_9614);
or U10251 (N_10251,N_9584,N_9784);
nand U10252 (N_10252,N_9453,N_9763);
xnor U10253 (N_10253,N_9748,N_9514);
and U10254 (N_10254,N_9942,N_9645);
or U10255 (N_10255,N_9808,N_9827);
or U10256 (N_10256,N_9688,N_9866);
xnor U10257 (N_10257,N_9723,N_9382);
nand U10258 (N_10258,N_9821,N_9522);
nor U10259 (N_10259,N_9696,N_9711);
nor U10260 (N_10260,N_9789,N_9499);
or U10261 (N_10261,N_9535,N_9567);
nand U10262 (N_10262,N_9533,N_9440);
nor U10263 (N_10263,N_9979,N_9381);
xor U10264 (N_10264,N_9624,N_9887);
xnor U10265 (N_10265,N_9980,N_9820);
and U10266 (N_10266,N_9946,N_9664);
and U10267 (N_10267,N_9963,N_9592);
xnor U10268 (N_10268,N_9392,N_9995);
and U10269 (N_10269,N_9595,N_9439);
or U10270 (N_10270,N_9838,N_9890);
nand U10271 (N_10271,N_9940,N_9428);
and U10272 (N_10272,N_9570,N_9759);
nor U10273 (N_10273,N_9660,N_9506);
nand U10274 (N_10274,N_9681,N_9394);
and U10275 (N_10275,N_9452,N_9888);
xor U10276 (N_10276,N_9893,N_9669);
or U10277 (N_10277,N_9418,N_9534);
or U10278 (N_10278,N_9665,N_9998);
nand U10279 (N_10279,N_9923,N_9741);
nor U10280 (N_10280,N_9438,N_9585);
nand U10281 (N_10281,N_9649,N_9654);
xor U10282 (N_10282,N_9622,N_9985);
nor U10283 (N_10283,N_9705,N_9850);
xnor U10284 (N_10284,N_9507,N_9573);
xor U10285 (N_10285,N_9913,N_9777);
and U10286 (N_10286,N_9762,N_9793);
nor U10287 (N_10287,N_9926,N_9544);
nor U10288 (N_10288,N_9627,N_9594);
nand U10289 (N_10289,N_9943,N_9778);
and U10290 (N_10290,N_9934,N_9815);
and U10291 (N_10291,N_9761,N_9906);
and U10292 (N_10292,N_9717,N_9659);
and U10293 (N_10293,N_9959,N_9587);
nor U10294 (N_10294,N_9551,N_9672);
xnor U10295 (N_10295,N_9526,N_9875);
nand U10296 (N_10296,N_9811,N_9629);
or U10297 (N_10297,N_9563,N_9743);
nor U10298 (N_10298,N_9432,N_9950);
xor U10299 (N_10299,N_9539,N_9384);
xor U10300 (N_10300,N_9572,N_9564);
nand U10301 (N_10301,N_9540,N_9386);
or U10302 (N_10302,N_9947,N_9799);
or U10303 (N_10303,N_9451,N_9677);
xor U10304 (N_10304,N_9682,N_9489);
or U10305 (N_10305,N_9874,N_9772);
xor U10306 (N_10306,N_9730,N_9707);
and U10307 (N_10307,N_9653,N_9469);
nand U10308 (N_10308,N_9845,N_9399);
and U10309 (N_10309,N_9788,N_9457);
or U10310 (N_10310,N_9973,N_9472);
nor U10311 (N_10311,N_9745,N_9470);
or U10312 (N_10312,N_9491,N_9376);
and U10313 (N_10313,N_9731,N_9836);
nand U10314 (N_10314,N_9681,N_9414);
or U10315 (N_10315,N_9665,N_9641);
xnor U10316 (N_10316,N_9964,N_9435);
xor U10317 (N_10317,N_9518,N_9744);
and U10318 (N_10318,N_9414,N_9996);
and U10319 (N_10319,N_9606,N_9673);
xor U10320 (N_10320,N_9993,N_9812);
xnor U10321 (N_10321,N_9862,N_9828);
nand U10322 (N_10322,N_9689,N_9605);
or U10323 (N_10323,N_9519,N_9436);
xnor U10324 (N_10324,N_9620,N_9980);
nand U10325 (N_10325,N_9693,N_9805);
xnor U10326 (N_10326,N_9896,N_9600);
nor U10327 (N_10327,N_9733,N_9441);
nand U10328 (N_10328,N_9915,N_9962);
or U10329 (N_10329,N_9615,N_9383);
and U10330 (N_10330,N_9934,N_9803);
nor U10331 (N_10331,N_9933,N_9761);
nor U10332 (N_10332,N_9508,N_9694);
xnor U10333 (N_10333,N_9724,N_9670);
xor U10334 (N_10334,N_9533,N_9458);
and U10335 (N_10335,N_9446,N_9811);
or U10336 (N_10336,N_9580,N_9828);
nor U10337 (N_10337,N_9924,N_9678);
nand U10338 (N_10338,N_9589,N_9552);
or U10339 (N_10339,N_9614,N_9712);
nand U10340 (N_10340,N_9841,N_9400);
xnor U10341 (N_10341,N_9432,N_9783);
nand U10342 (N_10342,N_9926,N_9641);
nand U10343 (N_10343,N_9962,N_9854);
nor U10344 (N_10344,N_9575,N_9838);
and U10345 (N_10345,N_9833,N_9784);
and U10346 (N_10346,N_9669,N_9795);
xnor U10347 (N_10347,N_9717,N_9406);
xor U10348 (N_10348,N_9553,N_9668);
nor U10349 (N_10349,N_9946,N_9464);
nand U10350 (N_10350,N_9441,N_9998);
and U10351 (N_10351,N_9685,N_9806);
nand U10352 (N_10352,N_9874,N_9536);
or U10353 (N_10353,N_9751,N_9760);
nand U10354 (N_10354,N_9946,N_9622);
and U10355 (N_10355,N_9910,N_9504);
and U10356 (N_10356,N_9700,N_9549);
nor U10357 (N_10357,N_9914,N_9609);
xnor U10358 (N_10358,N_9484,N_9465);
nor U10359 (N_10359,N_9736,N_9702);
nand U10360 (N_10360,N_9586,N_9953);
nand U10361 (N_10361,N_9710,N_9877);
and U10362 (N_10362,N_9729,N_9963);
or U10363 (N_10363,N_9722,N_9675);
and U10364 (N_10364,N_9460,N_9955);
and U10365 (N_10365,N_9496,N_9584);
and U10366 (N_10366,N_9454,N_9517);
and U10367 (N_10367,N_9705,N_9908);
nand U10368 (N_10368,N_9815,N_9640);
nor U10369 (N_10369,N_9655,N_9576);
xor U10370 (N_10370,N_9508,N_9577);
or U10371 (N_10371,N_9482,N_9824);
or U10372 (N_10372,N_9890,N_9615);
and U10373 (N_10373,N_9744,N_9849);
nand U10374 (N_10374,N_9607,N_9846);
nor U10375 (N_10375,N_9672,N_9864);
or U10376 (N_10376,N_9950,N_9528);
or U10377 (N_10377,N_9409,N_9624);
and U10378 (N_10378,N_9582,N_9604);
or U10379 (N_10379,N_9766,N_9597);
or U10380 (N_10380,N_9830,N_9906);
xnor U10381 (N_10381,N_9785,N_9548);
or U10382 (N_10382,N_9435,N_9952);
and U10383 (N_10383,N_9776,N_9995);
nand U10384 (N_10384,N_9513,N_9637);
xor U10385 (N_10385,N_9972,N_9484);
or U10386 (N_10386,N_9591,N_9612);
xnor U10387 (N_10387,N_9907,N_9440);
nor U10388 (N_10388,N_9797,N_9424);
nand U10389 (N_10389,N_9560,N_9446);
nor U10390 (N_10390,N_9990,N_9954);
xor U10391 (N_10391,N_9974,N_9641);
nand U10392 (N_10392,N_9980,N_9705);
xnor U10393 (N_10393,N_9895,N_9971);
xnor U10394 (N_10394,N_9423,N_9452);
xor U10395 (N_10395,N_9718,N_9456);
nor U10396 (N_10396,N_9910,N_9978);
nand U10397 (N_10397,N_9716,N_9880);
xor U10398 (N_10398,N_9903,N_9793);
or U10399 (N_10399,N_9705,N_9932);
nor U10400 (N_10400,N_9765,N_9444);
xor U10401 (N_10401,N_9687,N_9709);
nand U10402 (N_10402,N_9947,N_9582);
xor U10403 (N_10403,N_9520,N_9719);
xor U10404 (N_10404,N_9793,N_9922);
and U10405 (N_10405,N_9899,N_9717);
or U10406 (N_10406,N_9609,N_9638);
or U10407 (N_10407,N_9567,N_9613);
and U10408 (N_10408,N_9977,N_9998);
xor U10409 (N_10409,N_9830,N_9718);
nor U10410 (N_10410,N_9545,N_9825);
nand U10411 (N_10411,N_9837,N_9660);
xnor U10412 (N_10412,N_9592,N_9392);
nand U10413 (N_10413,N_9615,N_9456);
nand U10414 (N_10414,N_9634,N_9869);
nor U10415 (N_10415,N_9480,N_9883);
or U10416 (N_10416,N_9818,N_9756);
or U10417 (N_10417,N_9502,N_9980);
nor U10418 (N_10418,N_9479,N_9649);
or U10419 (N_10419,N_9453,N_9837);
nor U10420 (N_10420,N_9764,N_9424);
and U10421 (N_10421,N_9615,N_9682);
nor U10422 (N_10422,N_9963,N_9389);
or U10423 (N_10423,N_9553,N_9896);
xor U10424 (N_10424,N_9920,N_9680);
nand U10425 (N_10425,N_9613,N_9390);
xor U10426 (N_10426,N_9760,N_9757);
and U10427 (N_10427,N_9908,N_9443);
nand U10428 (N_10428,N_9907,N_9875);
xor U10429 (N_10429,N_9933,N_9572);
nand U10430 (N_10430,N_9558,N_9781);
xor U10431 (N_10431,N_9604,N_9824);
nor U10432 (N_10432,N_9641,N_9632);
xnor U10433 (N_10433,N_9564,N_9516);
xnor U10434 (N_10434,N_9697,N_9429);
or U10435 (N_10435,N_9888,N_9879);
xnor U10436 (N_10436,N_9951,N_9967);
or U10437 (N_10437,N_9487,N_9708);
nand U10438 (N_10438,N_9722,N_9624);
and U10439 (N_10439,N_9469,N_9425);
and U10440 (N_10440,N_9575,N_9790);
nand U10441 (N_10441,N_9866,N_9464);
nand U10442 (N_10442,N_9521,N_9738);
xnor U10443 (N_10443,N_9926,N_9543);
and U10444 (N_10444,N_9898,N_9560);
or U10445 (N_10445,N_9509,N_9959);
nor U10446 (N_10446,N_9642,N_9682);
xnor U10447 (N_10447,N_9725,N_9771);
xnor U10448 (N_10448,N_9728,N_9885);
and U10449 (N_10449,N_9942,N_9593);
nand U10450 (N_10450,N_9993,N_9810);
nor U10451 (N_10451,N_9478,N_9502);
nand U10452 (N_10452,N_9969,N_9530);
xnor U10453 (N_10453,N_9857,N_9813);
nand U10454 (N_10454,N_9898,N_9946);
nor U10455 (N_10455,N_9781,N_9929);
nor U10456 (N_10456,N_9816,N_9600);
nor U10457 (N_10457,N_9632,N_9875);
and U10458 (N_10458,N_9663,N_9570);
or U10459 (N_10459,N_9632,N_9452);
xor U10460 (N_10460,N_9662,N_9758);
xor U10461 (N_10461,N_9904,N_9900);
xnor U10462 (N_10462,N_9501,N_9721);
and U10463 (N_10463,N_9585,N_9898);
xnor U10464 (N_10464,N_9609,N_9712);
xor U10465 (N_10465,N_9378,N_9977);
nor U10466 (N_10466,N_9695,N_9864);
xor U10467 (N_10467,N_9947,N_9984);
and U10468 (N_10468,N_9712,N_9757);
xor U10469 (N_10469,N_9383,N_9890);
nor U10470 (N_10470,N_9739,N_9450);
or U10471 (N_10471,N_9840,N_9860);
xnor U10472 (N_10472,N_9524,N_9462);
nor U10473 (N_10473,N_9754,N_9686);
or U10474 (N_10474,N_9913,N_9878);
or U10475 (N_10475,N_9592,N_9443);
and U10476 (N_10476,N_9633,N_9524);
xor U10477 (N_10477,N_9894,N_9487);
nand U10478 (N_10478,N_9701,N_9509);
nor U10479 (N_10479,N_9619,N_9777);
or U10480 (N_10480,N_9912,N_9410);
and U10481 (N_10481,N_9554,N_9562);
nor U10482 (N_10482,N_9797,N_9532);
nand U10483 (N_10483,N_9845,N_9966);
nand U10484 (N_10484,N_9964,N_9618);
or U10485 (N_10485,N_9976,N_9719);
xnor U10486 (N_10486,N_9472,N_9587);
and U10487 (N_10487,N_9856,N_9936);
xor U10488 (N_10488,N_9587,N_9893);
and U10489 (N_10489,N_9899,N_9704);
nand U10490 (N_10490,N_9588,N_9786);
nand U10491 (N_10491,N_9746,N_9377);
and U10492 (N_10492,N_9395,N_9742);
nor U10493 (N_10493,N_9792,N_9785);
or U10494 (N_10494,N_9591,N_9633);
nand U10495 (N_10495,N_9987,N_9919);
and U10496 (N_10496,N_9686,N_9436);
nor U10497 (N_10497,N_9854,N_9417);
nor U10498 (N_10498,N_9945,N_9377);
and U10499 (N_10499,N_9537,N_9497);
nor U10500 (N_10500,N_9991,N_9393);
or U10501 (N_10501,N_9647,N_9632);
and U10502 (N_10502,N_9405,N_9696);
or U10503 (N_10503,N_9870,N_9549);
nor U10504 (N_10504,N_9984,N_9992);
xor U10505 (N_10505,N_9630,N_9440);
nor U10506 (N_10506,N_9710,N_9534);
nand U10507 (N_10507,N_9539,N_9653);
or U10508 (N_10508,N_9566,N_9427);
nand U10509 (N_10509,N_9915,N_9896);
nor U10510 (N_10510,N_9401,N_9678);
and U10511 (N_10511,N_9747,N_9380);
nand U10512 (N_10512,N_9956,N_9717);
xor U10513 (N_10513,N_9375,N_9442);
nor U10514 (N_10514,N_9812,N_9386);
nand U10515 (N_10515,N_9811,N_9991);
and U10516 (N_10516,N_9696,N_9655);
xnor U10517 (N_10517,N_9482,N_9774);
or U10518 (N_10518,N_9431,N_9844);
nand U10519 (N_10519,N_9440,N_9662);
xor U10520 (N_10520,N_9684,N_9993);
xnor U10521 (N_10521,N_9683,N_9772);
or U10522 (N_10522,N_9772,N_9477);
or U10523 (N_10523,N_9996,N_9497);
nor U10524 (N_10524,N_9644,N_9804);
or U10525 (N_10525,N_9894,N_9764);
nand U10526 (N_10526,N_9528,N_9594);
nor U10527 (N_10527,N_9474,N_9773);
or U10528 (N_10528,N_9679,N_9449);
or U10529 (N_10529,N_9904,N_9395);
nand U10530 (N_10530,N_9520,N_9706);
and U10531 (N_10531,N_9875,N_9498);
xnor U10532 (N_10532,N_9848,N_9841);
nor U10533 (N_10533,N_9721,N_9464);
nand U10534 (N_10534,N_9508,N_9928);
xnor U10535 (N_10535,N_9803,N_9741);
and U10536 (N_10536,N_9402,N_9760);
and U10537 (N_10537,N_9860,N_9996);
nand U10538 (N_10538,N_9577,N_9409);
nor U10539 (N_10539,N_9496,N_9846);
nor U10540 (N_10540,N_9670,N_9416);
or U10541 (N_10541,N_9793,N_9417);
and U10542 (N_10542,N_9725,N_9532);
nand U10543 (N_10543,N_9672,N_9490);
nor U10544 (N_10544,N_9880,N_9652);
and U10545 (N_10545,N_9434,N_9514);
nand U10546 (N_10546,N_9762,N_9696);
and U10547 (N_10547,N_9907,N_9446);
xor U10548 (N_10548,N_9992,N_9404);
and U10549 (N_10549,N_9896,N_9907);
nor U10550 (N_10550,N_9952,N_9860);
or U10551 (N_10551,N_9717,N_9442);
nand U10552 (N_10552,N_9712,N_9686);
xnor U10553 (N_10553,N_9386,N_9609);
nand U10554 (N_10554,N_9631,N_9457);
nor U10555 (N_10555,N_9577,N_9593);
nand U10556 (N_10556,N_9737,N_9596);
and U10557 (N_10557,N_9761,N_9778);
or U10558 (N_10558,N_9899,N_9724);
xnor U10559 (N_10559,N_9746,N_9882);
xor U10560 (N_10560,N_9689,N_9711);
nand U10561 (N_10561,N_9651,N_9510);
nor U10562 (N_10562,N_9648,N_9641);
and U10563 (N_10563,N_9578,N_9455);
and U10564 (N_10564,N_9943,N_9487);
or U10565 (N_10565,N_9747,N_9496);
nor U10566 (N_10566,N_9510,N_9491);
nand U10567 (N_10567,N_9620,N_9947);
nand U10568 (N_10568,N_9912,N_9648);
xnor U10569 (N_10569,N_9857,N_9517);
and U10570 (N_10570,N_9432,N_9450);
and U10571 (N_10571,N_9764,N_9469);
xor U10572 (N_10572,N_9571,N_9623);
and U10573 (N_10573,N_9802,N_9875);
or U10574 (N_10574,N_9605,N_9966);
or U10575 (N_10575,N_9956,N_9663);
nor U10576 (N_10576,N_9416,N_9457);
nor U10577 (N_10577,N_9403,N_9647);
and U10578 (N_10578,N_9768,N_9664);
xnor U10579 (N_10579,N_9556,N_9550);
xor U10580 (N_10580,N_9584,N_9622);
nor U10581 (N_10581,N_9843,N_9938);
and U10582 (N_10582,N_9548,N_9482);
nor U10583 (N_10583,N_9834,N_9803);
xnor U10584 (N_10584,N_9431,N_9780);
nand U10585 (N_10585,N_9831,N_9424);
nand U10586 (N_10586,N_9695,N_9783);
nand U10587 (N_10587,N_9443,N_9881);
and U10588 (N_10588,N_9405,N_9680);
nand U10589 (N_10589,N_9489,N_9549);
nand U10590 (N_10590,N_9877,N_9993);
or U10591 (N_10591,N_9800,N_9893);
nand U10592 (N_10592,N_9826,N_9780);
and U10593 (N_10593,N_9916,N_9557);
xor U10594 (N_10594,N_9738,N_9636);
and U10595 (N_10595,N_9948,N_9841);
xor U10596 (N_10596,N_9756,N_9812);
nor U10597 (N_10597,N_9421,N_9985);
nand U10598 (N_10598,N_9979,N_9927);
or U10599 (N_10599,N_9713,N_9403);
xnor U10600 (N_10600,N_9403,N_9609);
and U10601 (N_10601,N_9625,N_9473);
and U10602 (N_10602,N_9575,N_9624);
xor U10603 (N_10603,N_9456,N_9398);
and U10604 (N_10604,N_9820,N_9937);
nor U10605 (N_10605,N_9616,N_9657);
and U10606 (N_10606,N_9610,N_9456);
xnor U10607 (N_10607,N_9448,N_9735);
nor U10608 (N_10608,N_9528,N_9616);
and U10609 (N_10609,N_9458,N_9855);
or U10610 (N_10610,N_9614,N_9660);
nand U10611 (N_10611,N_9842,N_9817);
and U10612 (N_10612,N_9958,N_9861);
xnor U10613 (N_10613,N_9647,N_9532);
nand U10614 (N_10614,N_9678,N_9511);
nand U10615 (N_10615,N_9440,N_9577);
nand U10616 (N_10616,N_9655,N_9611);
nor U10617 (N_10617,N_9668,N_9900);
xnor U10618 (N_10618,N_9453,N_9760);
xnor U10619 (N_10619,N_9628,N_9656);
and U10620 (N_10620,N_9984,N_9843);
nand U10621 (N_10621,N_9589,N_9759);
or U10622 (N_10622,N_9937,N_9456);
xnor U10623 (N_10623,N_9414,N_9398);
nor U10624 (N_10624,N_9998,N_9521);
nor U10625 (N_10625,N_10020,N_10125);
and U10626 (N_10626,N_10417,N_10189);
nand U10627 (N_10627,N_10214,N_10498);
nand U10628 (N_10628,N_10314,N_10477);
nand U10629 (N_10629,N_10537,N_10600);
or U10630 (N_10630,N_10137,N_10155);
xnor U10631 (N_10631,N_10107,N_10004);
nor U10632 (N_10632,N_10355,N_10218);
nand U10633 (N_10633,N_10240,N_10006);
and U10634 (N_10634,N_10028,N_10396);
nor U10635 (N_10635,N_10301,N_10057);
xor U10636 (N_10636,N_10503,N_10543);
and U10637 (N_10637,N_10599,N_10444);
nand U10638 (N_10638,N_10463,N_10067);
nand U10639 (N_10639,N_10281,N_10465);
nor U10640 (N_10640,N_10063,N_10493);
xnor U10641 (N_10641,N_10364,N_10051);
or U10642 (N_10642,N_10603,N_10235);
or U10643 (N_10643,N_10297,N_10466);
and U10644 (N_10644,N_10306,N_10354);
nor U10645 (N_10645,N_10255,N_10391);
nor U10646 (N_10646,N_10030,N_10393);
nand U10647 (N_10647,N_10222,N_10581);
nand U10648 (N_10648,N_10487,N_10249);
nand U10649 (N_10649,N_10430,N_10367);
nor U10650 (N_10650,N_10029,N_10387);
or U10651 (N_10651,N_10315,N_10005);
nand U10652 (N_10652,N_10163,N_10259);
nor U10653 (N_10653,N_10335,N_10619);
or U10654 (N_10654,N_10494,N_10344);
or U10655 (N_10655,N_10054,N_10144);
xnor U10656 (N_10656,N_10188,N_10217);
and U10657 (N_10657,N_10021,N_10254);
nor U10658 (N_10658,N_10602,N_10452);
and U10659 (N_10659,N_10408,N_10076);
and U10660 (N_10660,N_10124,N_10224);
or U10661 (N_10661,N_10184,N_10010);
or U10662 (N_10662,N_10034,N_10129);
nand U10663 (N_10663,N_10490,N_10597);
nand U10664 (N_10664,N_10202,N_10071);
or U10665 (N_10665,N_10194,N_10516);
nor U10666 (N_10666,N_10548,N_10209);
xnor U10667 (N_10667,N_10100,N_10522);
xor U10668 (N_10668,N_10445,N_10571);
nor U10669 (N_10669,N_10366,N_10120);
and U10670 (N_10670,N_10081,N_10389);
or U10671 (N_10671,N_10577,N_10303);
xnor U10672 (N_10672,N_10458,N_10583);
xor U10673 (N_10673,N_10098,N_10165);
and U10674 (N_10674,N_10002,N_10008);
xnor U10675 (N_10675,N_10173,N_10433);
nor U10676 (N_10676,N_10461,N_10175);
and U10677 (N_10677,N_10261,N_10294);
nand U10678 (N_10678,N_10530,N_10378);
nand U10679 (N_10679,N_10312,N_10350);
nor U10680 (N_10680,N_10527,N_10183);
or U10681 (N_10681,N_10154,N_10035);
or U10682 (N_10682,N_10150,N_10251);
nand U10683 (N_10683,N_10171,N_10410);
nand U10684 (N_10684,N_10440,N_10455);
nor U10685 (N_10685,N_10232,N_10418);
xnor U10686 (N_10686,N_10404,N_10011);
nand U10687 (N_10687,N_10203,N_10561);
xor U10688 (N_10688,N_10308,N_10342);
or U10689 (N_10689,N_10015,N_10438);
nand U10690 (N_10690,N_10291,N_10346);
xnor U10691 (N_10691,N_10409,N_10595);
or U10692 (N_10692,N_10003,N_10095);
or U10693 (N_10693,N_10616,N_10206);
xnor U10694 (N_10694,N_10620,N_10453);
or U10695 (N_10695,N_10234,N_10450);
xor U10696 (N_10696,N_10119,N_10544);
nand U10697 (N_10697,N_10462,N_10106);
nor U10698 (N_10698,N_10267,N_10045);
xor U10699 (N_10699,N_10538,N_10307);
nand U10700 (N_10700,N_10041,N_10351);
and U10701 (N_10701,N_10193,N_10072);
and U10702 (N_10702,N_10093,N_10609);
nor U10703 (N_10703,N_10013,N_10488);
nand U10704 (N_10704,N_10509,N_10135);
xnor U10705 (N_10705,N_10186,N_10385);
xnor U10706 (N_10706,N_10166,N_10562);
nor U10707 (N_10707,N_10177,N_10241);
xnor U10708 (N_10708,N_10591,N_10607);
xor U10709 (N_10709,N_10078,N_10468);
nor U10710 (N_10710,N_10037,N_10141);
nand U10711 (N_10711,N_10176,N_10500);
or U10712 (N_10712,N_10549,N_10476);
or U10713 (N_10713,N_10428,N_10017);
or U10714 (N_10714,N_10330,N_10215);
or U10715 (N_10715,N_10457,N_10375);
xnor U10716 (N_10716,N_10127,N_10042);
or U10717 (N_10717,N_10533,N_10483);
nor U10718 (N_10718,N_10216,N_10091);
nor U10719 (N_10719,N_10180,N_10624);
nand U10720 (N_10720,N_10038,N_10491);
nand U10721 (N_10721,N_10399,N_10467);
nand U10722 (N_10722,N_10160,N_10394);
and U10723 (N_10723,N_10276,N_10134);
nor U10724 (N_10724,N_10511,N_10001);
nor U10725 (N_10725,N_10066,N_10575);
or U10726 (N_10726,N_10475,N_10579);
nor U10727 (N_10727,N_10074,N_10320);
nor U10728 (N_10728,N_10446,N_10227);
nand U10729 (N_10729,N_10372,N_10231);
nor U10730 (N_10730,N_10123,N_10473);
and U10731 (N_10731,N_10529,N_10300);
nand U10732 (N_10732,N_10429,N_10590);
nor U10733 (N_10733,N_10547,N_10223);
nor U10734 (N_10734,N_10401,N_10060);
nor U10735 (N_10735,N_10268,N_10299);
and U10736 (N_10736,N_10109,N_10586);
xnor U10737 (N_10737,N_10545,N_10053);
nand U10738 (N_10738,N_10061,N_10266);
nor U10739 (N_10739,N_10132,N_10158);
or U10740 (N_10740,N_10345,N_10079);
nand U10741 (N_10741,N_10258,N_10497);
xor U10742 (N_10742,N_10524,N_10392);
or U10743 (N_10743,N_10334,N_10148);
nor U10744 (N_10744,N_10432,N_10526);
xnor U10745 (N_10745,N_10534,N_10271);
xor U10746 (N_10746,N_10229,N_10088);
or U10747 (N_10747,N_10049,N_10610);
or U10748 (N_10748,N_10237,N_10230);
nor U10749 (N_10749,N_10523,N_10283);
and U10750 (N_10750,N_10167,N_10027);
nand U10751 (N_10751,N_10349,N_10402);
and U10752 (N_10752,N_10170,N_10302);
nand U10753 (N_10753,N_10421,N_10313);
nor U10754 (N_10754,N_10210,N_10605);
nand U10755 (N_10755,N_10289,N_10484);
xnor U10756 (N_10756,N_10515,N_10578);
nor U10757 (N_10757,N_10617,N_10564);
nand U10758 (N_10758,N_10133,N_10448);
xor U10759 (N_10759,N_10520,N_10069);
xnor U10760 (N_10760,N_10279,N_10309);
nor U10761 (N_10761,N_10540,N_10019);
nand U10762 (N_10762,N_10370,N_10192);
nor U10763 (N_10763,N_10437,N_10169);
or U10764 (N_10764,N_10039,N_10552);
and U10765 (N_10765,N_10615,N_10460);
nand U10766 (N_10766,N_10089,N_10513);
xnor U10767 (N_10767,N_10592,N_10598);
xor U10768 (N_10768,N_10246,N_10501);
and U10769 (N_10769,N_10032,N_10269);
xnor U10770 (N_10770,N_10555,N_10606);
nor U10771 (N_10771,N_10153,N_10566);
xnor U10772 (N_10772,N_10064,N_10338);
nor U10773 (N_10773,N_10225,N_10113);
xor U10774 (N_10774,N_10156,N_10521);
or U10775 (N_10775,N_10130,N_10442);
nor U10776 (N_10776,N_10360,N_10481);
nor U10777 (N_10777,N_10492,N_10587);
nand U10778 (N_10778,N_10226,N_10398);
nand U10779 (N_10779,N_10353,N_10018);
nor U10780 (N_10780,N_10556,N_10435);
and U10781 (N_10781,N_10146,N_10205);
and U10782 (N_10782,N_10256,N_10569);
nand U10783 (N_10783,N_10397,N_10085);
or U10784 (N_10784,N_10007,N_10075);
nor U10785 (N_10785,N_10142,N_10265);
and U10786 (N_10786,N_10567,N_10140);
xor U10787 (N_10787,N_10324,N_10425);
nand U10788 (N_10788,N_10196,N_10407);
or U10789 (N_10789,N_10439,N_10058);
xnor U10790 (N_10790,N_10187,N_10116);
xnor U10791 (N_10791,N_10377,N_10479);
or U10792 (N_10792,N_10369,N_10546);
and U10793 (N_10793,N_10292,N_10233);
and U10794 (N_10794,N_10036,N_10178);
nand U10795 (N_10795,N_10048,N_10162);
nand U10796 (N_10796,N_10025,N_10362);
xnor U10797 (N_10797,N_10204,N_10024);
nand U10798 (N_10798,N_10185,N_10449);
and U10799 (N_10799,N_10298,N_10097);
or U10800 (N_10800,N_10117,N_10244);
xor U10801 (N_10801,N_10560,N_10325);
nor U10802 (N_10802,N_10424,N_10043);
xor U10803 (N_10803,N_10262,N_10570);
xnor U10804 (N_10804,N_10273,N_10131);
nor U10805 (N_10805,N_10252,N_10339);
xnor U10806 (N_10806,N_10613,N_10584);
and U10807 (N_10807,N_10601,N_10427);
nand U10808 (N_10808,N_10031,N_10406);
or U10809 (N_10809,N_10507,N_10374);
nand U10810 (N_10810,N_10337,N_10373);
nor U10811 (N_10811,N_10363,N_10253);
nand U10812 (N_10812,N_10589,N_10441);
or U10813 (N_10813,N_10593,N_10506);
xor U10814 (N_10814,N_10248,N_10622);
nand U10815 (N_10815,N_10502,N_10270);
nand U10816 (N_10816,N_10508,N_10542);
nand U10817 (N_10817,N_10535,N_10104);
and U10818 (N_10818,N_10023,N_10618);
and U10819 (N_10819,N_10052,N_10086);
nor U10820 (N_10820,N_10247,N_10110);
xnor U10821 (N_10821,N_10288,N_10168);
xnor U10822 (N_10822,N_10604,N_10573);
or U10823 (N_10823,N_10000,N_10151);
and U10824 (N_10824,N_10574,N_10614);
xnor U10825 (N_10825,N_10212,N_10576);
nor U10826 (N_10826,N_10044,N_10356);
and U10827 (N_10827,N_10343,N_10105);
nand U10828 (N_10828,N_10138,N_10012);
nor U10829 (N_10829,N_10381,N_10147);
and U10830 (N_10830,N_10422,N_10191);
xnor U10831 (N_10831,N_10358,N_10594);
or U10832 (N_10832,N_10588,N_10321);
and U10833 (N_10833,N_10528,N_10263);
or U10834 (N_10834,N_10456,N_10318);
nand U10835 (N_10835,N_10236,N_10111);
and U10836 (N_10836,N_10347,N_10068);
and U10837 (N_10837,N_10277,N_10411);
and U10838 (N_10838,N_10272,N_10257);
nand U10839 (N_10839,N_10380,N_10447);
nor U10840 (N_10840,N_10046,N_10536);
and U10841 (N_10841,N_10050,N_10517);
nor U10842 (N_10842,N_10149,N_10357);
nor U10843 (N_10843,N_10388,N_10114);
xnor U10844 (N_10844,N_10532,N_10365);
nand U10845 (N_10845,N_10065,N_10416);
nand U10846 (N_10846,N_10621,N_10161);
or U10847 (N_10847,N_10096,N_10128);
or U10848 (N_10848,N_10480,N_10510);
or U10849 (N_10849,N_10403,N_10323);
xnor U10850 (N_10850,N_10239,N_10199);
or U10851 (N_10851,N_10296,N_10331);
xnor U10852 (N_10852,N_10379,N_10182);
nor U10853 (N_10853,N_10310,N_10539);
and U10854 (N_10854,N_10434,N_10181);
and U10855 (N_10855,N_10221,N_10126);
or U10856 (N_10856,N_10340,N_10612);
and U10857 (N_10857,N_10108,N_10213);
and U10858 (N_10858,N_10159,N_10368);
and U10859 (N_10859,N_10115,N_10541);
xor U10860 (N_10860,N_10080,N_10033);
or U10861 (N_10861,N_10073,N_10305);
or U10862 (N_10862,N_10197,N_10359);
nand U10863 (N_10863,N_10383,N_10101);
or U10864 (N_10864,N_10412,N_10563);
xnor U10865 (N_10865,N_10145,N_10519);
nand U10866 (N_10866,N_10431,N_10200);
xor U10867 (N_10867,N_10504,N_10022);
and U10868 (N_10868,N_10195,N_10495);
xnor U10869 (N_10869,N_10201,N_10486);
nor U10870 (N_10870,N_10489,N_10352);
nand U10871 (N_10871,N_10295,N_10623);
nand U10872 (N_10872,N_10557,N_10316);
xor U10873 (N_10873,N_10293,N_10290);
nor U10874 (N_10874,N_10414,N_10512);
or U10875 (N_10875,N_10275,N_10423);
xnor U10876 (N_10876,N_10384,N_10608);
or U10877 (N_10877,N_10284,N_10436);
and U10878 (N_10878,N_10568,N_10395);
xnor U10879 (N_10879,N_10443,N_10333);
xnor U10880 (N_10880,N_10471,N_10287);
xnor U10881 (N_10881,N_10611,N_10238);
or U10882 (N_10882,N_10092,N_10580);
nand U10883 (N_10883,N_10328,N_10157);
xnor U10884 (N_10884,N_10280,N_10152);
and U10885 (N_10885,N_10059,N_10274);
nor U10886 (N_10886,N_10582,N_10136);
nor U10887 (N_10887,N_10084,N_10220);
nand U10888 (N_10888,N_10371,N_10469);
xor U10889 (N_10889,N_10103,N_10329);
nand U10890 (N_10890,N_10099,N_10102);
and U10891 (N_10891,N_10317,N_10470);
nor U10892 (N_10892,N_10139,N_10174);
nand U10893 (N_10893,N_10122,N_10478);
nor U10894 (N_10894,N_10286,N_10327);
and U10895 (N_10895,N_10260,N_10454);
nor U10896 (N_10896,N_10550,N_10525);
nor U10897 (N_10897,N_10207,N_10070);
nor U10898 (N_10898,N_10243,N_10278);
or U10899 (N_10899,N_10083,N_10211);
xor U10900 (N_10900,N_10016,N_10499);
xnor U10901 (N_10901,N_10062,N_10558);
nand U10902 (N_10902,N_10172,N_10553);
xor U10903 (N_10903,N_10164,N_10348);
or U10904 (N_10904,N_10496,N_10426);
xor U10905 (N_10905,N_10040,N_10179);
and U10906 (N_10906,N_10474,N_10121);
nor U10907 (N_10907,N_10056,N_10319);
nor U10908 (N_10908,N_10245,N_10143);
or U10909 (N_10909,N_10219,N_10190);
and U10910 (N_10910,N_10400,N_10336);
and U10911 (N_10911,N_10326,N_10341);
and U10912 (N_10912,N_10118,N_10472);
nor U10913 (N_10913,N_10311,N_10596);
nand U10914 (N_10914,N_10282,N_10087);
and U10915 (N_10915,N_10228,N_10585);
and U10916 (N_10916,N_10112,N_10559);
or U10917 (N_10917,N_10415,N_10531);
nor U10918 (N_10918,N_10514,N_10208);
or U10919 (N_10919,N_10304,N_10451);
nor U10920 (N_10920,N_10026,N_10242);
and U10921 (N_10921,N_10382,N_10264);
nor U10922 (N_10922,N_10376,N_10485);
and U10923 (N_10923,N_10090,N_10014);
or U10924 (N_10924,N_10082,N_10482);
nor U10925 (N_10925,N_10077,N_10386);
xnor U10926 (N_10926,N_10551,N_10405);
nor U10927 (N_10927,N_10361,N_10572);
or U10928 (N_10928,N_10332,N_10250);
or U10929 (N_10929,N_10420,N_10554);
xor U10930 (N_10930,N_10390,N_10322);
xnor U10931 (N_10931,N_10419,N_10505);
nand U10932 (N_10932,N_10285,N_10094);
nor U10933 (N_10933,N_10055,N_10464);
or U10934 (N_10934,N_10413,N_10047);
nand U10935 (N_10935,N_10198,N_10459);
nor U10936 (N_10936,N_10565,N_10009);
xnor U10937 (N_10937,N_10518,N_10544);
and U10938 (N_10938,N_10550,N_10298);
nand U10939 (N_10939,N_10153,N_10550);
and U10940 (N_10940,N_10355,N_10624);
and U10941 (N_10941,N_10010,N_10311);
or U10942 (N_10942,N_10315,N_10402);
nor U10943 (N_10943,N_10210,N_10333);
and U10944 (N_10944,N_10565,N_10498);
nor U10945 (N_10945,N_10453,N_10427);
and U10946 (N_10946,N_10345,N_10439);
nor U10947 (N_10947,N_10352,N_10354);
or U10948 (N_10948,N_10277,N_10157);
or U10949 (N_10949,N_10536,N_10594);
nand U10950 (N_10950,N_10341,N_10284);
nor U10951 (N_10951,N_10581,N_10149);
nor U10952 (N_10952,N_10482,N_10581);
nor U10953 (N_10953,N_10228,N_10081);
nor U10954 (N_10954,N_10071,N_10431);
or U10955 (N_10955,N_10023,N_10006);
xor U10956 (N_10956,N_10022,N_10027);
xnor U10957 (N_10957,N_10619,N_10442);
or U10958 (N_10958,N_10584,N_10049);
and U10959 (N_10959,N_10605,N_10209);
nor U10960 (N_10960,N_10185,N_10409);
nand U10961 (N_10961,N_10197,N_10287);
nand U10962 (N_10962,N_10261,N_10559);
or U10963 (N_10963,N_10084,N_10502);
nor U10964 (N_10964,N_10525,N_10522);
or U10965 (N_10965,N_10610,N_10199);
xor U10966 (N_10966,N_10029,N_10007);
nor U10967 (N_10967,N_10456,N_10115);
nor U10968 (N_10968,N_10193,N_10010);
nor U10969 (N_10969,N_10458,N_10230);
or U10970 (N_10970,N_10091,N_10475);
and U10971 (N_10971,N_10322,N_10410);
xnor U10972 (N_10972,N_10533,N_10395);
xnor U10973 (N_10973,N_10334,N_10317);
or U10974 (N_10974,N_10481,N_10257);
or U10975 (N_10975,N_10607,N_10606);
or U10976 (N_10976,N_10420,N_10451);
nor U10977 (N_10977,N_10437,N_10151);
or U10978 (N_10978,N_10276,N_10390);
and U10979 (N_10979,N_10613,N_10376);
or U10980 (N_10980,N_10341,N_10026);
nor U10981 (N_10981,N_10359,N_10296);
nor U10982 (N_10982,N_10124,N_10364);
or U10983 (N_10983,N_10372,N_10085);
xnor U10984 (N_10984,N_10438,N_10148);
nor U10985 (N_10985,N_10082,N_10118);
nand U10986 (N_10986,N_10210,N_10094);
or U10987 (N_10987,N_10014,N_10306);
xnor U10988 (N_10988,N_10416,N_10171);
xor U10989 (N_10989,N_10099,N_10049);
nor U10990 (N_10990,N_10464,N_10098);
nand U10991 (N_10991,N_10127,N_10370);
xnor U10992 (N_10992,N_10152,N_10025);
nand U10993 (N_10993,N_10463,N_10167);
or U10994 (N_10994,N_10438,N_10312);
nor U10995 (N_10995,N_10263,N_10387);
xnor U10996 (N_10996,N_10290,N_10399);
nand U10997 (N_10997,N_10058,N_10030);
and U10998 (N_10998,N_10605,N_10112);
and U10999 (N_10999,N_10167,N_10016);
or U11000 (N_11000,N_10610,N_10245);
nor U11001 (N_11001,N_10336,N_10061);
xnor U11002 (N_11002,N_10119,N_10598);
or U11003 (N_11003,N_10208,N_10264);
and U11004 (N_11004,N_10449,N_10050);
nor U11005 (N_11005,N_10554,N_10244);
nor U11006 (N_11006,N_10502,N_10349);
or U11007 (N_11007,N_10061,N_10399);
nor U11008 (N_11008,N_10519,N_10188);
xor U11009 (N_11009,N_10372,N_10401);
nand U11010 (N_11010,N_10083,N_10402);
or U11011 (N_11011,N_10172,N_10556);
and U11012 (N_11012,N_10604,N_10495);
or U11013 (N_11013,N_10302,N_10213);
nor U11014 (N_11014,N_10394,N_10500);
and U11015 (N_11015,N_10481,N_10181);
nand U11016 (N_11016,N_10425,N_10553);
or U11017 (N_11017,N_10317,N_10125);
and U11018 (N_11018,N_10312,N_10365);
nor U11019 (N_11019,N_10586,N_10070);
xnor U11020 (N_11020,N_10416,N_10005);
nor U11021 (N_11021,N_10034,N_10548);
nand U11022 (N_11022,N_10332,N_10622);
or U11023 (N_11023,N_10082,N_10607);
or U11024 (N_11024,N_10112,N_10240);
nand U11025 (N_11025,N_10168,N_10020);
nor U11026 (N_11026,N_10284,N_10612);
xnor U11027 (N_11027,N_10066,N_10007);
and U11028 (N_11028,N_10067,N_10397);
nor U11029 (N_11029,N_10314,N_10195);
xnor U11030 (N_11030,N_10240,N_10115);
nand U11031 (N_11031,N_10455,N_10443);
and U11032 (N_11032,N_10119,N_10593);
nor U11033 (N_11033,N_10353,N_10504);
and U11034 (N_11034,N_10346,N_10608);
nor U11035 (N_11035,N_10193,N_10367);
or U11036 (N_11036,N_10467,N_10451);
nand U11037 (N_11037,N_10471,N_10098);
xnor U11038 (N_11038,N_10600,N_10281);
xor U11039 (N_11039,N_10098,N_10542);
nor U11040 (N_11040,N_10228,N_10468);
nand U11041 (N_11041,N_10526,N_10384);
or U11042 (N_11042,N_10561,N_10053);
nand U11043 (N_11043,N_10182,N_10161);
and U11044 (N_11044,N_10032,N_10408);
or U11045 (N_11045,N_10602,N_10181);
and U11046 (N_11046,N_10602,N_10148);
or U11047 (N_11047,N_10094,N_10032);
or U11048 (N_11048,N_10414,N_10493);
nand U11049 (N_11049,N_10234,N_10062);
xor U11050 (N_11050,N_10345,N_10413);
or U11051 (N_11051,N_10117,N_10095);
or U11052 (N_11052,N_10289,N_10546);
and U11053 (N_11053,N_10195,N_10373);
nand U11054 (N_11054,N_10041,N_10563);
nand U11055 (N_11055,N_10566,N_10344);
xor U11056 (N_11056,N_10613,N_10127);
nor U11057 (N_11057,N_10183,N_10424);
nand U11058 (N_11058,N_10123,N_10421);
or U11059 (N_11059,N_10319,N_10281);
nor U11060 (N_11060,N_10140,N_10094);
and U11061 (N_11061,N_10390,N_10573);
or U11062 (N_11062,N_10461,N_10394);
and U11063 (N_11063,N_10063,N_10255);
nand U11064 (N_11064,N_10603,N_10204);
or U11065 (N_11065,N_10475,N_10102);
nor U11066 (N_11066,N_10504,N_10208);
or U11067 (N_11067,N_10145,N_10446);
or U11068 (N_11068,N_10573,N_10302);
and U11069 (N_11069,N_10404,N_10005);
nand U11070 (N_11070,N_10232,N_10343);
and U11071 (N_11071,N_10260,N_10576);
or U11072 (N_11072,N_10085,N_10457);
nand U11073 (N_11073,N_10157,N_10339);
or U11074 (N_11074,N_10239,N_10201);
xor U11075 (N_11075,N_10167,N_10610);
nand U11076 (N_11076,N_10174,N_10225);
and U11077 (N_11077,N_10464,N_10146);
xor U11078 (N_11078,N_10405,N_10030);
or U11079 (N_11079,N_10256,N_10090);
or U11080 (N_11080,N_10568,N_10560);
nand U11081 (N_11081,N_10013,N_10374);
and U11082 (N_11082,N_10070,N_10568);
xor U11083 (N_11083,N_10246,N_10499);
or U11084 (N_11084,N_10234,N_10469);
and U11085 (N_11085,N_10504,N_10062);
and U11086 (N_11086,N_10406,N_10410);
xnor U11087 (N_11087,N_10430,N_10211);
or U11088 (N_11088,N_10338,N_10264);
nor U11089 (N_11089,N_10547,N_10244);
and U11090 (N_11090,N_10405,N_10075);
or U11091 (N_11091,N_10384,N_10531);
and U11092 (N_11092,N_10059,N_10082);
and U11093 (N_11093,N_10304,N_10386);
and U11094 (N_11094,N_10448,N_10461);
nor U11095 (N_11095,N_10312,N_10047);
nand U11096 (N_11096,N_10489,N_10223);
xnor U11097 (N_11097,N_10222,N_10451);
xor U11098 (N_11098,N_10022,N_10025);
xnor U11099 (N_11099,N_10310,N_10207);
nand U11100 (N_11100,N_10211,N_10259);
nor U11101 (N_11101,N_10475,N_10223);
nand U11102 (N_11102,N_10041,N_10583);
xor U11103 (N_11103,N_10041,N_10096);
nand U11104 (N_11104,N_10447,N_10544);
and U11105 (N_11105,N_10267,N_10534);
nand U11106 (N_11106,N_10529,N_10421);
nor U11107 (N_11107,N_10448,N_10364);
or U11108 (N_11108,N_10268,N_10082);
xor U11109 (N_11109,N_10290,N_10326);
nor U11110 (N_11110,N_10009,N_10410);
nand U11111 (N_11111,N_10315,N_10301);
or U11112 (N_11112,N_10002,N_10262);
nand U11113 (N_11113,N_10407,N_10162);
nor U11114 (N_11114,N_10280,N_10144);
nor U11115 (N_11115,N_10156,N_10133);
nor U11116 (N_11116,N_10511,N_10436);
nand U11117 (N_11117,N_10231,N_10164);
nand U11118 (N_11118,N_10126,N_10150);
nand U11119 (N_11119,N_10026,N_10397);
xor U11120 (N_11120,N_10144,N_10523);
nand U11121 (N_11121,N_10412,N_10203);
and U11122 (N_11122,N_10337,N_10176);
and U11123 (N_11123,N_10371,N_10162);
or U11124 (N_11124,N_10472,N_10288);
nand U11125 (N_11125,N_10341,N_10539);
or U11126 (N_11126,N_10537,N_10189);
nor U11127 (N_11127,N_10540,N_10534);
and U11128 (N_11128,N_10133,N_10341);
nor U11129 (N_11129,N_10466,N_10251);
and U11130 (N_11130,N_10058,N_10172);
nand U11131 (N_11131,N_10352,N_10104);
xnor U11132 (N_11132,N_10455,N_10422);
nand U11133 (N_11133,N_10162,N_10368);
nand U11134 (N_11134,N_10051,N_10485);
and U11135 (N_11135,N_10541,N_10252);
xor U11136 (N_11136,N_10321,N_10503);
or U11137 (N_11137,N_10327,N_10363);
nor U11138 (N_11138,N_10464,N_10290);
xor U11139 (N_11139,N_10486,N_10187);
nor U11140 (N_11140,N_10482,N_10510);
or U11141 (N_11141,N_10067,N_10241);
and U11142 (N_11142,N_10250,N_10530);
nand U11143 (N_11143,N_10523,N_10596);
or U11144 (N_11144,N_10520,N_10501);
or U11145 (N_11145,N_10083,N_10503);
nand U11146 (N_11146,N_10419,N_10451);
and U11147 (N_11147,N_10143,N_10180);
nand U11148 (N_11148,N_10458,N_10035);
nor U11149 (N_11149,N_10218,N_10539);
nor U11150 (N_11150,N_10067,N_10331);
and U11151 (N_11151,N_10178,N_10134);
and U11152 (N_11152,N_10230,N_10527);
or U11153 (N_11153,N_10018,N_10508);
nor U11154 (N_11154,N_10333,N_10389);
xnor U11155 (N_11155,N_10416,N_10128);
and U11156 (N_11156,N_10484,N_10477);
or U11157 (N_11157,N_10022,N_10365);
nor U11158 (N_11158,N_10217,N_10371);
and U11159 (N_11159,N_10009,N_10364);
nand U11160 (N_11160,N_10106,N_10378);
or U11161 (N_11161,N_10299,N_10535);
xor U11162 (N_11162,N_10485,N_10453);
nor U11163 (N_11163,N_10003,N_10157);
nand U11164 (N_11164,N_10459,N_10167);
xnor U11165 (N_11165,N_10021,N_10279);
xnor U11166 (N_11166,N_10525,N_10419);
and U11167 (N_11167,N_10150,N_10278);
or U11168 (N_11168,N_10542,N_10615);
and U11169 (N_11169,N_10351,N_10329);
nand U11170 (N_11170,N_10023,N_10571);
nor U11171 (N_11171,N_10167,N_10188);
xnor U11172 (N_11172,N_10589,N_10255);
and U11173 (N_11173,N_10202,N_10137);
and U11174 (N_11174,N_10027,N_10074);
and U11175 (N_11175,N_10284,N_10414);
nand U11176 (N_11176,N_10596,N_10050);
and U11177 (N_11177,N_10409,N_10280);
nor U11178 (N_11178,N_10295,N_10305);
nor U11179 (N_11179,N_10134,N_10157);
nor U11180 (N_11180,N_10192,N_10473);
nand U11181 (N_11181,N_10138,N_10039);
xnor U11182 (N_11182,N_10444,N_10371);
nor U11183 (N_11183,N_10388,N_10539);
nand U11184 (N_11184,N_10394,N_10426);
nand U11185 (N_11185,N_10207,N_10472);
nand U11186 (N_11186,N_10302,N_10249);
xor U11187 (N_11187,N_10286,N_10492);
nand U11188 (N_11188,N_10519,N_10312);
xnor U11189 (N_11189,N_10162,N_10411);
or U11190 (N_11190,N_10190,N_10057);
or U11191 (N_11191,N_10077,N_10287);
or U11192 (N_11192,N_10086,N_10320);
and U11193 (N_11193,N_10428,N_10081);
and U11194 (N_11194,N_10121,N_10278);
nor U11195 (N_11195,N_10222,N_10617);
or U11196 (N_11196,N_10482,N_10433);
nand U11197 (N_11197,N_10485,N_10424);
xor U11198 (N_11198,N_10062,N_10403);
or U11199 (N_11199,N_10029,N_10244);
or U11200 (N_11200,N_10067,N_10324);
nor U11201 (N_11201,N_10376,N_10594);
nor U11202 (N_11202,N_10060,N_10366);
and U11203 (N_11203,N_10517,N_10306);
and U11204 (N_11204,N_10191,N_10592);
or U11205 (N_11205,N_10552,N_10212);
nor U11206 (N_11206,N_10241,N_10506);
nor U11207 (N_11207,N_10198,N_10082);
or U11208 (N_11208,N_10546,N_10526);
xnor U11209 (N_11209,N_10309,N_10126);
xor U11210 (N_11210,N_10090,N_10502);
and U11211 (N_11211,N_10035,N_10405);
or U11212 (N_11212,N_10092,N_10300);
nor U11213 (N_11213,N_10465,N_10052);
and U11214 (N_11214,N_10518,N_10197);
nor U11215 (N_11215,N_10211,N_10623);
and U11216 (N_11216,N_10557,N_10544);
or U11217 (N_11217,N_10037,N_10408);
xnor U11218 (N_11218,N_10392,N_10190);
or U11219 (N_11219,N_10412,N_10020);
xor U11220 (N_11220,N_10005,N_10165);
xnor U11221 (N_11221,N_10489,N_10006);
nor U11222 (N_11222,N_10246,N_10261);
and U11223 (N_11223,N_10285,N_10248);
xnor U11224 (N_11224,N_10575,N_10582);
nand U11225 (N_11225,N_10171,N_10567);
xnor U11226 (N_11226,N_10570,N_10019);
nor U11227 (N_11227,N_10168,N_10604);
and U11228 (N_11228,N_10235,N_10443);
or U11229 (N_11229,N_10160,N_10269);
or U11230 (N_11230,N_10085,N_10389);
xnor U11231 (N_11231,N_10063,N_10360);
and U11232 (N_11232,N_10567,N_10620);
and U11233 (N_11233,N_10614,N_10254);
xnor U11234 (N_11234,N_10318,N_10168);
nand U11235 (N_11235,N_10347,N_10367);
or U11236 (N_11236,N_10540,N_10380);
xor U11237 (N_11237,N_10113,N_10062);
xnor U11238 (N_11238,N_10136,N_10440);
nor U11239 (N_11239,N_10210,N_10474);
and U11240 (N_11240,N_10271,N_10337);
or U11241 (N_11241,N_10272,N_10427);
xor U11242 (N_11242,N_10332,N_10583);
nor U11243 (N_11243,N_10503,N_10553);
nor U11244 (N_11244,N_10348,N_10352);
or U11245 (N_11245,N_10554,N_10391);
and U11246 (N_11246,N_10298,N_10135);
or U11247 (N_11247,N_10372,N_10361);
nand U11248 (N_11248,N_10326,N_10383);
or U11249 (N_11249,N_10208,N_10525);
nand U11250 (N_11250,N_10676,N_10722);
and U11251 (N_11251,N_10988,N_10778);
xor U11252 (N_11252,N_10886,N_10963);
xnor U11253 (N_11253,N_11122,N_10652);
nor U11254 (N_11254,N_11058,N_11129);
nand U11255 (N_11255,N_11148,N_11013);
and U11256 (N_11256,N_11157,N_10893);
nor U11257 (N_11257,N_10701,N_11040);
and U11258 (N_11258,N_11047,N_11233);
and U11259 (N_11259,N_10929,N_10744);
or U11260 (N_11260,N_10944,N_10838);
nand U11261 (N_11261,N_10877,N_11135);
and U11262 (N_11262,N_10712,N_11017);
and U11263 (N_11263,N_11239,N_11195);
nand U11264 (N_11264,N_10834,N_11089);
and U11265 (N_11265,N_10991,N_11043);
nand U11266 (N_11266,N_11042,N_10885);
and U11267 (N_11267,N_10897,N_10949);
xor U11268 (N_11268,N_11073,N_10969);
xnor U11269 (N_11269,N_11224,N_10688);
nand U11270 (N_11270,N_10696,N_10842);
xor U11271 (N_11271,N_10642,N_10999);
nand U11272 (N_11272,N_10715,N_11082);
and U11273 (N_11273,N_10937,N_10862);
nand U11274 (N_11274,N_10864,N_11235);
nor U11275 (N_11275,N_10729,N_10987);
or U11276 (N_11276,N_11211,N_10972);
nor U11277 (N_11277,N_10917,N_11039);
and U11278 (N_11278,N_10665,N_11117);
nand U11279 (N_11279,N_10779,N_11010);
nor U11280 (N_11280,N_10690,N_10694);
and U11281 (N_11281,N_11190,N_10835);
xor U11282 (N_11282,N_10967,N_10793);
xor U11283 (N_11283,N_10852,N_11203);
and U11284 (N_11284,N_10750,N_10892);
nand U11285 (N_11285,N_10713,N_10824);
and U11286 (N_11286,N_10931,N_11174);
or U11287 (N_11287,N_11212,N_11034);
xnor U11288 (N_11288,N_10792,N_10662);
and U11289 (N_11289,N_10751,N_10871);
nand U11290 (N_11290,N_10936,N_10961);
and U11291 (N_11291,N_11238,N_10640);
nor U11292 (N_11292,N_11092,N_11242);
nand U11293 (N_11293,N_10724,N_10818);
or U11294 (N_11294,N_10958,N_10723);
and U11295 (N_11295,N_10634,N_11020);
and U11296 (N_11296,N_10669,N_11151);
and U11297 (N_11297,N_11119,N_11103);
xor U11298 (N_11298,N_11121,N_11231);
nor U11299 (N_11299,N_11230,N_10785);
xor U11300 (N_11300,N_10799,N_11142);
or U11301 (N_11301,N_10819,N_10625);
nand U11302 (N_11302,N_11194,N_10664);
xor U11303 (N_11303,N_10757,N_11139);
xor U11304 (N_11304,N_10687,N_10795);
xor U11305 (N_11305,N_11182,N_11169);
nand U11306 (N_11306,N_11220,N_10776);
and U11307 (N_11307,N_10794,N_10764);
nor U11308 (N_11308,N_10780,N_11120);
and U11309 (N_11309,N_11002,N_10727);
nor U11310 (N_11310,N_10800,N_11023);
or U11311 (N_11311,N_10895,N_11018);
or U11312 (N_11312,N_10741,N_10813);
and U11313 (N_11313,N_10959,N_11009);
nor U11314 (N_11314,N_11199,N_11068);
or U11315 (N_11315,N_11214,N_10925);
nor U11316 (N_11316,N_10884,N_11116);
and U11317 (N_11317,N_10636,N_10889);
nand U11318 (N_11318,N_10883,N_11081);
nand U11319 (N_11319,N_10839,N_10657);
nor U11320 (N_11320,N_10859,N_10675);
or U11321 (N_11321,N_10769,N_10922);
xor U11322 (N_11322,N_11221,N_10890);
or U11323 (N_11323,N_10853,N_11037);
xor U11324 (N_11324,N_11038,N_10844);
or U11325 (N_11325,N_10704,N_10858);
or U11326 (N_11326,N_10945,N_10656);
or U11327 (N_11327,N_11031,N_10771);
nand U11328 (N_11328,N_11210,N_10777);
and U11329 (N_11329,N_10627,N_11246);
nand U11330 (N_11330,N_10783,N_11025);
nand U11331 (N_11331,N_10789,N_11229);
nand U11332 (N_11332,N_11111,N_10717);
xor U11333 (N_11333,N_11140,N_11163);
and U11334 (N_11334,N_10797,N_11022);
nand U11335 (N_11335,N_11207,N_10882);
nand U11336 (N_11336,N_10948,N_10737);
nand U11337 (N_11337,N_10887,N_10721);
or U11338 (N_11338,N_11057,N_10957);
nand U11339 (N_11339,N_11027,N_10847);
and U11340 (N_11340,N_10697,N_10649);
xnor U11341 (N_11341,N_10924,N_10683);
or U11342 (N_11342,N_10720,N_10784);
or U11343 (N_11343,N_10740,N_10881);
xor U11344 (N_11344,N_11007,N_11192);
and U11345 (N_11345,N_10909,N_10989);
xor U11346 (N_11346,N_10761,N_10896);
nand U11347 (N_11347,N_11044,N_10747);
or U11348 (N_11348,N_11014,N_11079);
xnor U11349 (N_11349,N_11130,N_11209);
nand U11350 (N_11350,N_11005,N_10663);
nand U11351 (N_11351,N_11074,N_10731);
xnor U11352 (N_11352,N_10906,N_10666);
and U11353 (N_11353,N_11184,N_10983);
xnor U11354 (N_11354,N_10860,N_11241);
nor U11355 (N_11355,N_10770,N_10742);
xnor U11356 (N_11356,N_11024,N_10933);
or U11357 (N_11357,N_10997,N_11217);
xor U11358 (N_11358,N_11205,N_11249);
or U11359 (N_11359,N_10708,N_10833);
nand U11360 (N_11360,N_10910,N_11201);
nand U11361 (N_11361,N_11064,N_10828);
nor U11362 (N_11362,N_10935,N_10996);
xor U11363 (N_11363,N_10667,N_11104);
and U11364 (N_11364,N_11091,N_10756);
nor U11365 (N_11365,N_10826,N_10848);
xor U11366 (N_11366,N_10695,N_11245);
nor U11367 (N_11367,N_10661,N_10982);
nand U11368 (N_11368,N_11223,N_11186);
xor U11369 (N_11369,N_10953,N_10758);
nor U11370 (N_11370,N_11158,N_10643);
nor U11371 (N_11371,N_10907,N_10686);
nand U11372 (N_11372,N_11200,N_10787);
xor U11373 (N_11373,N_10861,N_10814);
xnor U11374 (N_11374,N_10626,N_10802);
and U11375 (N_11375,N_11088,N_11152);
and U11376 (N_11376,N_10926,N_11016);
nor U11377 (N_11377,N_10843,N_11054);
and U11378 (N_11378,N_10692,N_10762);
and U11379 (N_11379,N_10766,N_11164);
nand U11380 (N_11380,N_11096,N_10812);
nor U11381 (N_11381,N_11180,N_11226);
and U11382 (N_11382,N_10680,N_10898);
and U11383 (N_11383,N_10702,N_11030);
and U11384 (N_11384,N_10808,N_11049);
and U11385 (N_11385,N_11065,N_10806);
nor U11386 (N_11386,N_10811,N_10816);
or U11387 (N_11387,N_11185,N_10798);
nand U11388 (N_11388,N_11066,N_10920);
or U11389 (N_11389,N_10921,N_10790);
nor U11390 (N_11390,N_11087,N_11227);
nor U11391 (N_11391,N_11133,N_11021);
xnor U11392 (N_11392,N_10714,N_10960);
or U11393 (N_11393,N_10829,N_10857);
nor U11394 (N_11394,N_11015,N_10706);
or U11395 (N_11395,N_11166,N_11095);
xor U11396 (N_11396,N_10955,N_10934);
nand U11397 (N_11397,N_11191,N_11171);
or U11398 (N_11398,N_10840,N_10781);
nand U11399 (N_11399,N_10685,N_10942);
nand U11400 (N_11400,N_11046,N_10699);
xnor U11401 (N_11401,N_10850,N_10810);
and U11402 (N_11402,N_10651,N_10730);
or U11403 (N_11403,N_10950,N_10817);
or U11404 (N_11404,N_11181,N_10980);
xor U11405 (N_11405,N_10995,N_11094);
nor U11406 (N_11406,N_10752,N_10974);
and U11407 (N_11407,N_11189,N_11067);
or U11408 (N_11408,N_11100,N_11056);
or U11409 (N_11409,N_10658,N_10733);
nor U11410 (N_11410,N_10947,N_10849);
nand U11411 (N_11411,N_10970,N_10872);
or U11412 (N_11412,N_11032,N_10998);
xor U11413 (N_11413,N_11219,N_10992);
or U11414 (N_11414,N_10773,N_11041);
xor U11415 (N_11415,N_11055,N_10875);
and U11416 (N_11416,N_10763,N_10964);
and U11417 (N_11417,N_11161,N_10807);
and U11418 (N_11418,N_10728,N_10707);
and U11419 (N_11419,N_11247,N_11216);
nor U11420 (N_11420,N_10648,N_11126);
and U11421 (N_11421,N_11108,N_10775);
nor U11422 (N_11422,N_10759,N_10670);
nor U11423 (N_11423,N_10628,N_11144);
and U11424 (N_11424,N_11237,N_10919);
nor U11425 (N_11425,N_11143,N_10888);
xnor U11426 (N_11426,N_10845,N_10954);
nor U11427 (N_11427,N_11213,N_11125);
xnor U11428 (N_11428,N_10638,N_11076);
and U11429 (N_11429,N_11150,N_11168);
nor U11430 (N_11430,N_10746,N_10951);
nor U11431 (N_11431,N_11138,N_10673);
and U11432 (N_11432,N_10805,N_10856);
or U11433 (N_11433,N_11036,N_11167);
nand U11434 (N_11434,N_11061,N_10975);
and U11435 (N_11435,N_10841,N_10674);
xor U11436 (N_11436,N_11072,N_10863);
xnor U11437 (N_11437,N_10901,N_10635);
xnor U11438 (N_11438,N_11175,N_10946);
nor U11439 (N_11439,N_10985,N_10976);
nor U11440 (N_11440,N_10705,N_10911);
nor U11441 (N_11441,N_11053,N_10956);
and U11442 (N_11442,N_10788,N_11083);
nand U11443 (N_11443,N_10679,N_10718);
and U11444 (N_11444,N_11170,N_11172);
xor U11445 (N_11445,N_10908,N_11202);
xnor U11446 (N_11446,N_11136,N_11177);
xnor U11447 (N_11447,N_10873,N_10905);
nand U11448 (N_11448,N_10732,N_11196);
nor U11449 (N_11449,N_10938,N_10912);
nor U11450 (N_11450,N_11156,N_10827);
xor U11451 (N_11451,N_11098,N_10943);
and U11452 (N_11452,N_10637,N_10903);
or U11453 (N_11453,N_11085,N_11198);
nor U11454 (N_11454,N_11244,N_10641);
nor U11455 (N_11455,N_10820,N_11029);
nor U11456 (N_11456,N_10854,N_11075);
xor U11457 (N_11457,N_10772,N_10880);
nor U11458 (N_11458,N_11033,N_10633);
xor U11459 (N_11459,N_11028,N_10866);
or U11460 (N_11460,N_11128,N_10681);
and U11461 (N_11461,N_10966,N_10973);
xnor U11462 (N_11462,N_11124,N_11187);
xor U11463 (N_11463,N_11131,N_11109);
and U11464 (N_11464,N_11110,N_11078);
xnor U11465 (N_11465,N_10739,N_11162);
nand U11466 (N_11466,N_11069,N_11147);
nand U11467 (N_11467,N_10639,N_10913);
nor U11468 (N_11468,N_10825,N_11101);
xor U11469 (N_11469,N_10902,N_10647);
nor U11470 (N_11470,N_10869,N_10914);
or U11471 (N_11471,N_10804,N_11063);
nand U11472 (N_11472,N_10801,N_11232);
xor U11473 (N_11473,N_10918,N_10753);
xor U11474 (N_11474,N_10791,N_11060);
and U11475 (N_11475,N_11225,N_11149);
and U11476 (N_11476,N_11178,N_10645);
xor U11477 (N_11477,N_11008,N_10711);
or U11478 (N_11478,N_10928,N_11146);
or U11479 (N_11479,N_10900,N_11160);
and U11480 (N_11480,N_11080,N_10962);
nor U11481 (N_11481,N_10644,N_11222);
xor U11482 (N_11482,N_10735,N_10968);
xor U11483 (N_11483,N_11003,N_10993);
or U11484 (N_11484,N_11099,N_11011);
and U11485 (N_11485,N_11004,N_11102);
or U11486 (N_11486,N_10868,N_10655);
or U11487 (N_11487,N_11000,N_11123);
or U11488 (N_11488,N_10894,N_10650);
or U11489 (N_11489,N_10932,N_10930);
xnor U11490 (N_11490,N_11026,N_10803);
nand U11491 (N_11491,N_10977,N_11093);
nor U11492 (N_11492,N_10749,N_11153);
or U11493 (N_11493,N_11204,N_10703);
or U11494 (N_11494,N_10738,N_11206);
nor U11495 (N_11495,N_10981,N_10952);
and U11496 (N_11496,N_10986,N_10874);
and U11497 (N_11497,N_11070,N_11215);
or U11498 (N_11498,N_11112,N_11208);
or U11499 (N_11499,N_10755,N_10836);
or U11500 (N_11500,N_10831,N_11165);
nand U11501 (N_11501,N_10725,N_11107);
nor U11502 (N_11502,N_10629,N_10677);
xor U11503 (N_11503,N_11154,N_10672);
nor U11504 (N_11504,N_10754,N_10767);
nor U11505 (N_11505,N_10878,N_10984);
nand U11506 (N_11506,N_10646,N_10979);
nand U11507 (N_11507,N_10865,N_10891);
xnor U11508 (N_11508,N_11248,N_10734);
nand U11509 (N_11509,N_10855,N_10668);
xnor U11510 (N_11510,N_11141,N_11243);
and U11511 (N_11511,N_11137,N_11114);
or U11512 (N_11512,N_11086,N_10823);
nor U11513 (N_11513,N_10916,N_10927);
or U11514 (N_11514,N_10786,N_11228);
nor U11515 (N_11515,N_10700,N_11234);
nand U11516 (N_11516,N_10631,N_10830);
and U11517 (N_11517,N_10870,N_11045);
xor U11518 (N_11518,N_10815,N_11012);
xnor U11519 (N_11519,N_11240,N_11097);
and U11520 (N_11520,N_11183,N_10923);
nor U11521 (N_11521,N_11059,N_11132);
and U11522 (N_11522,N_10796,N_10904);
xor U11523 (N_11523,N_10748,N_11084);
nand U11524 (N_11524,N_11127,N_10994);
or U11525 (N_11525,N_11155,N_11113);
and U11526 (N_11526,N_10678,N_11236);
and U11527 (N_11527,N_10736,N_10971);
nand U11528 (N_11528,N_11115,N_10990);
and U11529 (N_11529,N_10709,N_10716);
xor U11530 (N_11530,N_10743,N_11188);
xor U11531 (N_11531,N_10654,N_11105);
nand U11532 (N_11532,N_10745,N_11106);
nor U11533 (N_11533,N_10939,N_11173);
nor U11534 (N_11534,N_10660,N_10821);
nor U11535 (N_11535,N_11179,N_10698);
nor U11536 (N_11536,N_10978,N_10632);
and U11537 (N_11537,N_10689,N_11218);
nor U11538 (N_11538,N_10682,N_10768);
or U11539 (N_11539,N_10832,N_10837);
nor U11540 (N_11540,N_11145,N_11071);
or U11541 (N_11541,N_10899,N_10940);
xnor U11542 (N_11542,N_11090,N_10876);
or U11543 (N_11543,N_10630,N_10851);
nor U11544 (N_11544,N_10760,N_10879);
and U11545 (N_11545,N_11134,N_11118);
nor U11546 (N_11546,N_11197,N_10659);
and U11547 (N_11547,N_10710,N_10765);
or U11548 (N_11548,N_11050,N_11052);
nand U11549 (N_11549,N_10691,N_11006);
or U11550 (N_11550,N_10782,N_10965);
or U11551 (N_11551,N_11019,N_10693);
nand U11552 (N_11552,N_11159,N_10774);
nand U11553 (N_11553,N_10915,N_11001);
or U11554 (N_11554,N_10846,N_10822);
nor U11555 (N_11555,N_10867,N_10671);
xor U11556 (N_11556,N_10653,N_11051);
nand U11557 (N_11557,N_10809,N_10719);
xnor U11558 (N_11558,N_10684,N_10941);
xor U11559 (N_11559,N_11035,N_11048);
nor U11560 (N_11560,N_11193,N_11077);
and U11561 (N_11561,N_10726,N_11062);
and U11562 (N_11562,N_11176,N_11211);
nand U11563 (N_11563,N_11092,N_10942);
and U11564 (N_11564,N_10775,N_11088);
and U11565 (N_11565,N_11104,N_10637);
nor U11566 (N_11566,N_10701,N_10866);
xor U11567 (N_11567,N_10701,N_11191);
or U11568 (N_11568,N_10973,N_10718);
and U11569 (N_11569,N_10726,N_10974);
nor U11570 (N_11570,N_11171,N_10816);
and U11571 (N_11571,N_11168,N_10885);
and U11572 (N_11572,N_11072,N_10784);
and U11573 (N_11573,N_10904,N_11127);
nand U11574 (N_11574,N_10864,N_10877);
nor U11575 (N_11575,N_10672,N_10665);
nand U11576 (N_11576,N_11099,N_11246);
nor U11577 (N_11577,N_10798,N_10806);
and U11578 (N_11578,N_11082,N_11118);
nand U11579 (N_11579,N_11243,N_10722);
and U11580 (N_11580,N_10719,N_10871);
nor U11581 (N_11581,N_10631,N_10810);
nor U11582 (N_11582,N_10983,N_10625);
and U11583 (N_11583,N_10755,N_10754);
or U11584 (N_11584,N_10799,N_11218);
xnor U11585 (N_11585,N_10896,N_10850);
nand U11586 (N_11586,N_11229,N_11243);
nor U11587 (N_11587,N_10865,N_10912);
nor U11588 (N_11588,N_10868,N_11224);
nand U11589 (N_11589,N_10885,N_10915);
nand U11590 (N_11590,N_10985,N_10913);
or U11591 (N_11591,N_11225,N_10881);
or U11592 (N_11592,N_10938,N_11115);
or U11593 (N_11593,N_10696,N_11044);
nand U11594 (N_11594,N_10870,N_10731);
xor U11595 (N_11595,N_11200,N_10781);
nor U11596 (N_11596,N_11009,N_11195);
or U11597 (N_11597,N_10909,N_10668);
and U11598 (N_11598,N_10864,N_11117);
or U11599 (N_11599,N_11156,N_10641);
xnor U11600 (N_11600,N_10993,N_11140);
nand U11601 (N_11601,N_10661,N_11176);
xor U11602 (N_11602,N_10687,N_11175);
and U11603 (N_11603,N_10739,N_10818);
nand U11604 (N_11604,N_10922,N_10979);
nor U11605 (N_11605,N_10775,N_10820);
xnor U11606 (N_11606,N_10963,N_10762);
nand U11607 (N_11607,N_10627,N_10975);
nand U11608 (N_11608,N_11031,N_10701);
or U11609 (N_11609,N_11240,N_10679);
or U11610 (N_11610,N_11215,N_10690);
or U11611 (N_11611,N_10830,N_11207);
and U11612 (N_11612,N_10925,N_10868);
and U11613 (N_11613,N_11142,N_10851);
or U11614 (N_11614,N_11151,N_10833);
and U11615 (N_11615,N_10970,N_11126);
nor U11616 (N_11616,N_11061,N_11059);
xnor U11617 (N_11617,N_10762,N_10694);
xor U11618 (N_11618,N_11026,N_10923);
or U11619 (N_11619,N_11186,N_10759);
nor U11620 (N_11620,N_10699,N_11017);
xnor U11621 (N_11621,N_10865,N_11037);
xor U11622 (N_11622,N_11148,N_11112);
or U11623 (N_11623,N_10765,N_10933);
nand U11624 (N_11624,N_11097,N_11235);
nand U11625 (N_11625,N_11125,N_10659);
xnor U11626 (N_11626,N_10818,N_11208);
xor U11627 (N_11627,N_10761,N_10644);
xnor U11628 (N_11628,N_10916,N_11030);
xnor U11629 (N_11629,N_11154,N_11233);
or U11630 (N_11630,N_10922,N_10757);
nor U11631 (N_11631,N_11232,N_10861);
xnor U11632 (N_11632,N_10724,N_10863);
xor U11633 (N_11633,N_11142,N_11017);
xor U11634 (N_11634,N_11131,N_11064);
and U11635 (N_11635,N_10915,N_10707);
nor U11636 (N_11636,N_11192,N_10873);
and U11637 (N_11637,N_11181,N_11077);
or U11638 (N_11638,N_11178,N_11190);
and U11639 (N_11639,N_10742,N_10971);
nand U11640 (N_11640,N_11105,N_10735);
and U11641 (N_11641,N_10645,N_11035);
nor U11642 (N_11642,N_10627,N_10829);
nand U11643 (N_11643,N_11226,N_10892);
nand U11644 (N_11644,N_11181,N_10842);
xnor U11645 (N_11645,N_11181,N_10647);
and U11646 (N_11646,N_10774,N_10836);
nor U11647 (N_11647,N_10841,N_11125);
nor U11648 (N_11648,N_11171,N_10679);
or U11649 (N_11649,N_10941,N_11048);
or U11650 (N_11650,N_10856,N_11024);
nor U11651 (N_11651,N_10759,N_10991);
or U11652 (N_11652,N_10957,N_11012);
nand U11653 (N_11653,N_10804,N_11178);
or U11654 (N_11654,N_10846,N_11240);
or U11655 (N_11655,N_11246,N_11142);
or U11656 (N_11656,N_10956,N_11177);
and U11657 (N_11657,N_10811,N_11194);
xor U11658 (N_11658,N_11215,N_10969);
nand U11659 (N_11659,N_10953,N_10817);
and U11660 (N_11660,N_10939,N_10645);
xnor U11661 (N_11661,N_11228,N_11000);
nand U11662 (N_11662,N_10968,N_10880);
xor U11663 (N_11663,N_10893,N_11105);
or U11664 (N_11664,N_10960,N_10938);
nor U11665 (N_11665,N_10906,N_10792);
nand U11666 (N_11666,N_10837,N_11203);
or U11667 (N_11667,N_11062,N_10952);
nand U11668 (N_11668,N_10923,N_11156);
xor U11669 (N_11669,N_10894,N_10746);
xnor U11670 (N_11670,N_11107,N_10789);
xnor U11671 (N_11671,N_10994,N_11045);
and U11672 (N_11672,N_10861,N_10832);
nand U11673 (N_11673,N_10996,N_10856);
nor U11674 (N_11674,N_11247,N_10853);
or U11675 (N_11675,N_10828,N_10839);
xor U11676 (N_11676,N_10757,N_10740);
nand U11677 (N_11677,N_10787,N_10991);
and U11678 (N_11678,N_11190,N_11236);
and U11679 (N_11679,N_10651,N_11152);
and U11680 (N_11680,N_10948,N_10996);
and U11681 (N_11681,N_10729,N_11228);
nand U11682 (N_11682,N_10767,N_10974);
xnor U11683 (N_11683,N_11238,N_10973);
and U11684 (N_11684,N_11086,N_11197);
nor U11685 (N_11685,N_10891,N_10923);
xor U11686 (N_11686,N_10834,N_10677);
or U11687 (N_11687,N_10743,N_10866);
or U11688 (N_11688,N_10884,N_10948);
or U11689 (N_11689,N_10790,N_10719);
and U11690 (N_11690,N_10777,N_10764);
xor U11691 (N_11691,N_11090,N_10747);
xor U11692 (N_11692,N_10905,N_10879);
or U11693 (N_11693,N_10909,N_11221);
nand U11694 (N_11694,N_11004,N_11086);
nand U11695 (N_11695,N_11046,N_10891);
and U11696 (N_11696,N_10807,N_11153);
nand U11697 (N_11697,N_11201,N_10946);
nand U11698 (N_11698,N_10981,N_11199);
or U11699 (N_11699,N_10978,N_10640);
nor U11700 (N_11700,N_10797,N_10731);
or U11701 (N_11701,N_10770,N_10720);
xnor U11702 (N_11702,N_11075,N_11030);
or U11703 (N_11703,N_10778,N_11229);
nand U11704 (N_11704,N_10650,N_11143);
nor U11705 (N_11705,N_10919,N_10688);
nor U11706 (N_11706,N_10641,N_11062);
nand U11707 (N_11707,N_10751,N_10737);
and U11708 (N_11708,N_10850,N_11230);
or U11709 (N_11709,N_10929,N_11161);
or U11710 (N_11710,N_11164,N_10889);
nor U11711 (N_11711,N_10801,N_11157);
nand U11712 (N_11712,N_10784,N_10660);
or U11713 (N_11713,N_10722,N_10735);
or U11714 (N_11714,N_10658,N_10852);
or U11715 (N_11715,N_11240,N_11092);
xor U11716 (N_11716,N_10690,N_11196);
or U11717 (N_11717,N_10838,N_11220);
or U11718 (N_11718,N_11130,N_10854);
and U11719 (N_11719,N_10788,N_10837);
or U11720 (N_11720,N_11010,N_10873);
xor U11721 (N_11721,N_11134,N_10948);
nand U11722 (N_11722,N_10699,N_10926);
nand U11723 (N_11723,N_10824,N_11035);
xnor U11724 (N_11724,N_10658,N_10684);
nor U11725 (N_11725,N_10867,N_10801);
nand U11726 (N_11726,N_10790,N_11006);
and U11727 (N_11727,N_10721,N_10889);
xnor U11728 (N_11728,N_11127,N_11024);
and U11729 (N_11729,N_10977,N_10750);
nor U11730 (N_11730,N_10876,N_10681);
nand U11731 (N_11731,N_11241,N_10692);
nand U11732 (N_11732,N_10634,N_10925);
nor U11733 (N_11733,N_11164,N_10967);
nand U11734 (N_11734,N_10970,N_11097);
or U11735 (N_11735,N_10846,N_11024);
and U11736 (N_11736,N_11126,N_10978);
or U11737 (N_11737,N_10806,N_10876);
xor U11738 (N_11738,N_10691,N_10814);
and U11739 (N_11739,N_11049,N_10910);
xnor U11740 (N_11740,N_10963,N_10846);
or U11741 (N_11741,N_10649,N_10915);
and U11742 (N_11742,N_11186,N_10791);
nand U11743 (N_11743,N_10779,N_10671);
nor U11744 (N_11744,N_10762,N_11073);
or U11745 (N_11745,N_10821,N_10942);
nand U11746 (N_11746,N_10815,N_10878);
nand U11747 (N_11747,N_10655,N_11005);
xor U11748 (N_11748,N_10952,N_10670);
nor U11749 (N_11749,N_11094,N_10625);
nor U11750 (N_11750,N_10746,N_10928);
and U11751 (N_11751,N_10929,N_10782);
and U11752 (N_11752,N_10782,N_11079);
or U11753 (N_11753,N_11047,N_10996);
xnor U11754 (N_11754,N_11026,N_10731);
and U11755 (N_11755,N_11221,N_11012);
and U11756 (N_11756,N_10687,N_11075);
nand U11757 (N_11757,N_10632,N_11059);
xor U11758 (N_11758,N_10859,N_11110);
xnor U11759 (N_11759,N_10954,N_10949);
nand U11760 (N_11760,N_10677,N_10849);
xor U11761 (N_11761,N_10889,N_10694);
xor U11762 (N_11762,N_11249,N_10886);
xnor U11763 (N_11763,N_11063,N_11125);
or U11764 (N_11764,N_10744,N_11168);
nand U11765 (N_11765,N_10789,N_10953);
nand U11766 (N_11766,N_10998,N_11045);
or U11767 (N_11767,N_11166,N_10893);
or U11768 (N_11768,N_10727,N_10969);
nand U11769 (N_11769,N_11168,N_10653);
nor U11770 (N_11770,N_10739,N_10681);
and U11771 (N_11771,N_10717,N_10762);
nor U11772 (N_11772,N_10815,N_10635);
nor U11773 (N_11773,N_10705,N_11034);
xnor U11774 (N_11774,N_10723,N_10694);
nor U11775 (N_11775,N_10660,N_11112);
xor U11776 (N_11776,N_11021,N_10885);
and U11777 (N_11777,N_10655,N_10710);
or U11778 (N_11778,N_11058,N_10740);
or U11779 (N_11779,N_10776,N_10700);
or U11780 (N_11780,N_11140,N_11228);
xor U11781 (N_11781,N_10746,N_11100);
nor U11782 (N_11782,N_10981,N_11052);
or U11783 (N_11783,N_11031,N_10816);
xnor U11784 (N_11784,N_10725,N_10777);
or U11785 (N_11785,N_11151,N_11217);
xnor U11786 (N_11786,N_10990,N_10985);
and U11787 (N_11787,N_10973,N_11195);
xnor U11788 (N_11788,N_10859,N_11028);
xnor U11789 (N_11789,N_11004,N_10656);
and U11790 (N_11790,N_10823,N_10826);
nor U11791 (N_11791,N_11042,N_10672);
nor U11792 (N_11792,N_11156,N_10694);
and U11793 (N_11793,N_10847,N_11062);
or U11794 (N_11794,N_10934,N_11036);
or U11795 (N_11795,N_11038,N_11221);
xor U11796 (N_11796,N_10957,N_11145);
or U11797 (N_11797,N_10860,N_11060);
or U11798 (N_11798,N_11088,N_11094);
and U11799 (N_11799,N_10674,N_11038);
nand U11800 (N_11800,N_10754,N_11248);
and U11801 (N_11801,N_11002,N_10805);
nand U11802 (N_11802,N_11245,N_10662);
and U11803 (N_11803,N_10982,N_10909);
and U11804 (N_11804,N_10805,N_11235);
nand U11805 (N_11805,N_10855,N_10811);
or U11806 (N_11806,N_10866,N_10630);
nor U11807 (N_11807,N_10882,N_10998);
nand U11808 (N_11808,N_10922,N_10744);
or U11809 (N_11809,N_10726,N_10907);
nor U11810 (N_11810,N_11169,N_10912);
nand U11811 (N_11811,N_10772,N_10800);
nor U11812 (N_11812,N_10756,N_11025);
and U11813 (N_11813,N_10681,N_10841);
nand U11814 (N_11814,N_10673,N_11097);
xor U11815 (N_11815,N_10958,N_10816);
or U11816 (N_11816,N_10827,N_10821);
and U11817 (N_11817,N_10643,N_11023);
xnor U11818 (N_11818,N_10684,N_10806);
and U11819 (N_11819,N_10745,N_10860);
xor U11820 (N_11820,N_11096,N_11094);
nor U11821 (N_11821,N_10664,N_10715);
and U11822 (N_11822,N_11077,N_10765);
or U11823 (N_11823,N_10939,N_10945);
or U11824 (N_11824,N_10687,N_11076);
nor U11825 (N_11825,N_11117,N_10961);
xnor U11826 (N_11826,N_10646,N_10809);
and U11827 (N_11827,N_11189,N_11111);
or U11828 (N_11828,N_10643,N_10999);
or U11829 (N_11829,N_10787,N_10982);
or U11830 (N_11830,N_10912,N_10952);
and U11831 (N_11831,N_10924,N_10633);
nand U11832 (N_11832,N_11242,N_10871);
nor U11833 (N_11833,N_11166,N_11245);
nor U11834 (N_11834,N_10625,N_10746);
nor U11835 (N_11835,N_10633,N_11072);
nand U11836 (N_11836,N_10994,N_11200);
xor U11837 (N_11837,N_10834,N_11118);
or U11838 (N_11838,N_11126,N_10995);
xnor U11839 (N_11839,N_11033,N_11110);
or U11840 (N_11840,N_10683,N_10866);
nand U11841 (N_11841,N_11182,N_10871);
nor U11842 (N_11842,N_10918,N_10632);
and U11843 (N_11843,N_10966,N_11094);
nand U11844 (N_11844,N_10736,N_10877);
xor U11845 (N_11845,N_10806,N_10909);
nand U11846 (N_11846,N_10839,N_11159);
or U11847 (N_11847,N_11075,N_10953);
nor U11848 (N_11848,N_10809,N_11162);
nor U11849 (N_11849,N_10913,N_10908);
xor U11850 (N_11850,N_10887,N_10934);
and U11851 (N_11851,N_11067,N_10809);
nor U11852 (N_11852,N_10868,N_10989);
nand U11853 (N_11853,N_11162,N_10785);
nor U11854 (N_11854,N_10927,N_11040);
or U11855 (N_11855,N_11085,N_10803);
xnor U11856 (N_11856,N_10805,N_11031);
nand U11857 (N_11857,N_10839,N_10769);
nor U11858 (N_11858,N_10863,N_11232);
nor U11859 (N_11859,N_10763,N_10683);
nor U11860 (N_11860,N_10980,N_11096);
or U11861 (N_11861,N_10835,N_11062);
nor U11862 (N_11862,N_10827,N_11015);
nand U11863 (N_11863,N_10760,N_10647);
or U11864 (N_11864,N_10820,N_11161);
xor U11865 (N_11865,N_10905,N_10952);
nand U11866 (N_11866,N_10665,N_11165);
and U11867 (N_11867,N_10745,N_10905);
or U11868 (N_11868,N_10838,N_11043);
nand U11869 (N_11869,N_11024,N_10748);
and U11870 (N_11870,N_11065,N_10660);
or U11871 (N_11871,N_11158,N_11159);
xor U11872 (N_11872,N_10818,N_10976);
or U11873 (N_11873,N_11133,N_11239);
and U11874 (N_11874,N_10738,N_11148);
nand U11875 (N_11875,N_11430,N_11505);
and U11876 (N_11876,N_11283,N_11780);
and U11877 (N_11877,N_11758,N_11294);
nand U11878 (N_11878,N_11831,N_11607);
nor U11879 (N_11879,N_11458,N_11477);
nand U11880 (N_11880,N_11502,N_11318);
or U11881 (N_11881,N_11545,N_11394);
nand U11882 (N_11882,N_11753,N_11614);
and U11883 (N_11883,N_11671,N_11496);
nand U11884 (N_11884,N_11290,N_11714);
xor U11885 (N_11885,N_11587,N_11651);
nand U11886 (N_11886,N_11300,N_11795);
nor U11887 (N_11887,N_11360,N_11588);
or U11888 (N_11888,N_11484,N_11821);
nand U11889 (N_11889,N_11736,N_11703);
xor U11890 (N_11890,N_11303,N_11514);
xnor U11891 (N_11891,N_11422,N_11779);
and U11892 (N_11892,N_11532,N_11759);
or U11893 (N_11893,N_11688,N_11486);
and U11894 (N_11894,N_11834,N_11464);
or U11895 (N_11895,N_11629,N_11811);
xnor U11896 (N_11896,N_11694,N_11278);
nand U11897 (N_11897,N_11507,N_11251);
nor U11898 (N_11898,N_11510,N_11563);
xnor U11899 (N_11899,N_11579,N_11827);
or U11900 (N_11900,N_11730,N_11570);
and U11901 (N_11901,N_11874,N_11566);
xnor U11902 (N_11902,N_11280,N_11552);
nand U11903 (N_11903,N_11462,N_11749);
or U11904 (N_11904,N_11351,N_11538);
and U11905 (N_11905,N_11645,N_11344);
or U11906 (N_11906,N_11818,N_11358);
xor U11907 (N_11907,N_11723,N_11312);
and U11908 (N_11908,N_11316,N_11633);
nor U11909 (N_11909,N_11812,N_11619);
nor U11910 (N_11910,N_11508,N_11757);
or U11911 (N_11911,N_11698,N_11289);
nand U11912 (N_11912,N_11425,N_11589);
and U11913 (N_11913,N_11867,N_11324);
nor U11914 (N_11914,N_11338,N_11838);
nand U11915 (N_11915,N_11768,N_11426);
nand U11916 (N_11916,N_11597,N_11382);
or U11917 (N_11917,N_11761,N_11481);
nor U11918 (N_11918,N_11847,N_11330);
xnor U11919 (N_11919,N_11729,N_11727);
nor U11920 (N_11920,N_11349,N_11849);
nor U11921 (N_11921,N_11371,N_11606);
nor U11922 (N_11922,N_11769,N_11770);
xor U11923 (N_11923,N_11465,N_11431);
and U11924 (N_11924,N_11712,N_11334);
or U11925 (N_11925,N_11355,N_11257);
xnor U11926 (N_11926,N_11561,N_11540);
nand U11927 (N_11927,N_11390,N_11495);
xor U11928 (N_11928,N_11569,N_11443);
nor U11929 (N_11929,N_11754,N_11807);
nand U11930 (N_11930,N_11678,N_11436);
nor U11931 (N_11931,N_11347,N_11695);
xnor U11932 (N_11932,N_11262,N_11663);
nor U11933 (N_11933,N_11775,N_11644);
nor U11934 (N_11934,N_11685,N_11476);
and U11935 (N_11935,N_11268,N_11771);
xor U11936 (N_11936,N_11764,N_11562);
or U11937 (N_11937,N_11529,N_11622);
nand U11938 (N_11938,N_11583,N_11466);
xnor U11939 (N_11939,N_11853,N_11500);
nand U11940 (N_11940,N_11591,N_11252);
or U11941 (N_11941,N_11325,N_11517);
nand U11942 (N_11942,N_11845,N_11787);
and U11943 (N_11943,N_11846,N_11533);
and U11944 (N_11944,N_11367,N_11593);
and U11945 (N_11945,N_11391,N_11718);
nand U11946 (N_11946,N_11317,N_11469);
xnor U11947 (N_11947,N_11420,N_11634);
nand U11948 (N_11948,N_11839,N_11599);
nor U11949 (N_11949,N_11667,N_11813);
and U11950 (N_11950,N_11711,N_11253);
nand U11951 (N_11951,N_11863,N_11261);
xor U11952 (N_11952,N_11616,N_11442);
xnor U11953 (N_11953,N_11642,N_11379);
nand U11954 (N_11954,N_11281,N_11407);
nor U11955 (N_11955,N_11833,N_11474);
nand U11956 (N_11956,N_11320,N_11499);
xnor U11957 (N_11957,N_11470,N_11661);
nand U11958 (N_11958,N_11781,N_11554);
and U11959 (N_11959,N_11665,N_11692);
nor U11960 (N_11960,N_11456,N_11733);
xnor U11961 (N_11961,N_11372,N_11441);
and U11962 (N_11962,N_11814,N_11708);
nor U11963 (N_11963,N_11704,N_11725);
xor U11964 (N_11964,N_11269,N_11746);
or U11965 (N_11965,N_11806,N_11447);
nor U11966 (N_11966,N_11732,N_11259);
and U11967 (N_11967,N_11669,N_11864);
or U11968 (N_11968,N_11670,N_11788);
or U11969 (N_11969,N_11717,N_11817);
and U11970 (N_11970,N_11627,N_11679);
nand U11971 (N_11971,N_11326,N_11673);
nor U11972 (N_11972,N_11415,N_11339);
xor U11973 (N_11973,N_11307,N_11329);
xnor U11974 (N_11974,N_11478,N_11271);
xor U11975 (N_11975,N_11286,N_11859);
or U11976 (N_11976,N_11352,N_11672);
or U11977 (N_11977,N_11328,N_11416);
nand U11978 (N_11978,N_11292,N_11792);
nand U11979 (N_11979,N_11560,N_11624);
or U11980 (N_11980,N_11632,N_11410);
xor U11981 (N_11981,N_11745,N_11653);
and U11982 (N_11982,N_11590,N_11751);
xnor U11983 (N_11983,N_11636,N_11686);
nand U11984 (N_11984,N_11424,N_11585);
or U11985 (N_11985,N_11374,N_11423);
nor U11986 (N_11986,N_11274,N_11648);
or U11987 (N_11987,N_11345,N_11835);
and U11988 (N_11988,N_11767,N_11612);
and U11989 (N_11989,N_11401,N_11809);
or U11990 (N_11990,N_11870,N_11828);
xnor U11991 (N_11991,N_11641,N_11494);
or U11992 (N_11992,N_11558,N_11542);
nor U11993 (N_11993,N_11309,N_11368);
xor U11994 (N_11994,N_11518,N_11819);
nor U11995 (N_11995,N_11836,N_11799);
nor U11996 (N_11996,N_11432,N_11284);
or U11997 (N_11997,N_11473,N_11549);
nor U11998 (N_11998,N_11305,N_11592);
xnor U11999 (N_11999,N_11315,N_11868);
xor U12000 (N_12000,N_11709,N_11618);
and U12001 (N_12001,N_11735,N_11264);
or U12002 (N_12002,N_11652,N_11387);
nor U12003 (N_12003,N_11706,N_11501);
and U12004 (N_12004,N_11630,N_11408);
xnor U12005 (N_12005,N_11567,N_11263);
or U12006 (N_12006,N_11395,N_11800);
or U12007 (N_12007,N_11364,N_11854);
or U12008 (N_12008,N_11375,N_11705);
and U12009 (N_12009,N_11490,N_11621);
xnor U12010 (N_12010,N_11454,N_11635);
nand U12011 (N_12011,N_11646,N_11666);
and U12012 (N_12012,N_11815,N_11580);
nand U12013 (N_12013,N_11689,N_11471);
nor U12014 (N_12014,N_11610,N_11675);
and U12015 (N_12015,N_11722,N_11656);
or U12016 (N_12016,N_11600,N_11536);
xor U12017 (N_12017,N_11460,N_11392);
nor U12018 (N_12018,N_11611,N_11457);
or U12019 (N_12019,N_11791,N_11412);
nor U12020 (N_12020,N_11535,N_11413);
or U12021 (N_12021,N_11522,N_11363);
xnor U12022 (N_12022,N_11340,N_11438);
or U12023 (N_12023,N_11620,N_11448);
nand U12024 (N_12024,N_11523,N_11657);
or U12025 (N_12025,N_11664,N_11285);
xnor U12026 (N_12026,N_11393,N_11322);
nand U12027 (N_12027,N_11304,N_11643);
xnor U12028 (N_12028,N_11556,N_11575);
nand U12029 (N_12029,N_11451,N_11265);
or U12030 (N_12030,N_11683,N_11343);
or U12031 (N_12031,N_11615,N_11639);
or U12032 (N_12032,N_11276,N_11681);
nand U12033 (N_12033,N_11760,N_11427);
xor U12034 (N_12034,N_11707,N_11319);
nand U12035 (N_12035,N_11737,N_11728);
and U12036 (N_12036,N_11796,N_11342);
or U12037 (N_12037,N_11862,N_11258);
xor U12038 (N_12038,N_11842,N_11539);
and U12039 (N_12039,N_11783,N_11295);
nor U12040 (N_12040,N_11802,N_11527);
nand U12041 (N_12041,N_11810,N_11720);
nand U12042 (N_12042,N_11871,N_11804);
nand U12043 (N_12043,N_11491,N_11411);
nand U12044 (N_12044,N_11713,N_11386);
or U12045 (N_12045,N_11861,N_11437);
nand U12046 (N_12046,N_11526,N_11385);
xor U12047 (N_12047,N_11816,N_11548);
xnor U12048 (N_12048,N_11452,N_11359);
nor U12049 (N_12049,N_11298,N_11299);
or U12050 (N_12050,N_11805,N_11521);
and U12051 (N_12051,N_11376,N_11366);
and U12052 (N_12052,N_11837,N_11254);
and U12053 (N_12053,N_11266,N_11346);
or U12054 (N_12054,N_11773,N_11841);
nor U12055 (N_12055,N_11640,N_11668);
or U12056 (N_12056,N_11399,N_11658);
xnor U12057 (N_12057,N_11763,N_11798);
xnor U12058 (N_12058,N_11573,N_11260);
and U12059 (N_12059,N_11335,N_11357);
or U12060 (N_12060,N_11701,N_11513);
xor U12061 (N_12061,N_11699,N_11564);
xor U12062 (N_12062,N_11855,N_11848);
xnor U12063 (N_12063,N_11414,N_11336);
nand U12064 (N_12064,N_11604,N_11647);
xor U12065 (N_12065,N_11479,N_11482);
or U12066 (N_12066,N_11444,N_11492);
or U12067 (N_12067,N_11608,N_11716);
xor U12068 (N_12068,N_11865,N_11524);
nor U12069 (N_12069,N_11744,N_11421);
nor U12070 (N_12070,N_11696,N_11302);
nand U12071 (N_12071,N_11565,N_11279);
xor U12072 (N_12072,N_11520,N_11715);
nand U12073 (N_12073,N_11777,N_11310);
nor U12074 (N_12074,N_11288,N_11786);
nand U12075 (N_12075,N_11512,N_11577);
or U12076 (N_12076,N_11361,N_11748);
nor U12077 (N_12077,N_11404,N_11445);
or U12078 (N_12078,N_11772,N_11388);
xor U12079 (N_12079,N_11553,N_11740);
and U12080 (N_12080,N_11406,N_11778);
nand U12081 (N_12081,N_11369,N_11873);
and U12082 (N_12082,N_11762,N_11398);
nor U12083 (N_12083,N_11596,N_11480);
and U12084 (N_12084,N_11793,N_11581);
xor U12085 (N_12085,N_11256,N_11409);
nor U12086 (N_12086,N_11691,N_11468);
and U12087 (N_12087,N_11774,N_11851);
and U12088 (N_12088,N_11497,N_11544);
nor U12089 (N_12089,N_11626,N_11852);
xnor U12090 (N_12090,N_11293,N_11439);
nand U12091 (N_12091,N_11595,N_11353);
nand U12092 (N_12092,N_11377,N_11726);
or U12093 (N_12093,N_11296,N_11677);
xnor U12094 (N_12094,N_11825,N_11693);
and U12095 (N_12095,N_11598,N_11383);
xnor U12096 (N_12096,N_11586,N_11537);
nand U12097 (N_12097,N_11820,N_11623);
xnor U12098 (N_12098,N_11282,N_11272);
and U12099 (N_12099,N_11857,N_11824);
and U12100 (N_12100,N_11277,N_11333);
nor U12101 (N_12101,N_11273,N_11493);
xnor U12102 (N_12102,N_11850,N_11337);
or U12103 (N_12103,N_11547,N_11455);
xor U12104 (N_12104,N_11250,N_11475);
or U12105 (N_12105,N_11756,N_11743);
nor U12106 (N_12106,N_11790,N_11826);
nand U12107 (N_12107,N_11637,N_11840);
or U12108 (N_12108,N_11797,N_11378);
xor U12109 (N_12109,N_11301,N_11662);
nor U12110 (N_12110,N_11690,N_11823);
xor U12111 (N_12111,N_11741,N_11435);
or U12112 (N_12112,N_11747,N_11434);
nand U12113 (N_12113,N_11739,N_11559);
nor U12114 (N_12114,N_11396,N_11801);
xor U12115 (N_12115,N_11543,N_11323);
nor U12116 (N_12116,N_11356,N_11511);
nand U12117 (N_12117,N_11384,N_11461);
or U12118 (N_12118,N_11546,N_11789);
and U12119 (N_12119,N_11370,N_11467);
or U12120 (N_12120,N_11687,N_11676);
and U12121 (N_12121,N_11794,N_11785);
nor U12122 (N_12122,N_11287,N_11638);
nor U12123 (N_12123,N_11381,N_11843);
and U12124 (N_12124,N_11306,N_11625);
or U12125 (N_12125,N_11530,N_11446);
and U12126 (N_12126,N_11700,N_11734);
nand U12127 (N_12127,N_11682,N_11459);
nand U12128 (N_12128,N_11551,N_11750);
xnor U12129 (N_12129,N_11555,N_11489);
and U12130 (N_12130,N_11308,N_11869);
xor U12131 (N_12131,N_11354,N_11582);
nor U12132 (N_12132,N_11568,N_11397);
or U12133 (N_12133,N_11605,N_11534);
and U12134 (N_12134,N_11291,N_11576);
and U12135 (N_12135,N_11418,N_11327);
nand U12136 (N_12136,N_11365,N_11649);
or U12137 (N_12137,N_11341,N_11516);
or U12138 (N_12138,N_11557,N_11731);
or U12139 (N_12139,N_11659,N_11485);
and U12140 (N_12140,N_11483,N_11449);
nand U12141 (N_12141,N_11509,N_11602);
nand U12142 (N_12142,N_11525,N_11405);
xnor U12143 (N_12143,N_11830,N_11419);
and U12144 (N_12144,N_11601,N_11721);
nor U12145 (N_12145,N_11428,N_11710);
nand U12146 (N_12146,N_11541,N_11631);
nand U12147 (N_12147,N_11680,N_11572);
or U12148 (N_12148,N_11498,N_11650);
nand U12149 (N_12149,N_11275,N_11584);
nand U12150 (N_12150,N_11782,N_11402);
xor U12151 (N_12151,N_11684,N_11311);
nor U12152 (N_12152,N_11488,N_11255);
nor U12153 (N_12153,N_11822,N_11550);
nand U12154 (N_12154,N_11429,N_11858);
xnor U12155 (N_12155,N_11674,N_11350);
nand U12156 (N_12156,N_11844,N_11503);
nor U12157 (N_12157,N_11531,N_11578);
xor U12158 (N_12158,N_11702,N_11784);
xor U12159 (N_12159,N_11872,N_11463);
nand U12160 (N_12160,N_11603,N_11380);
nand U12161 (N_12161,N_11755,N_11832);
xnor U12162 (N_12162,N_11313,N_11719);
xnor U12163 (N_12163,N_11504,N_11609);
nor U12164 (N_12164,N_11808,N_11403);
xor U12165 (N_12165,N_11297,N_11472);
nand U12166 (N_12166,N_11628,N_11417);
or U12167 (N_12167,N_11594,N_11321);
or U12168 (N_12168,N_11450,N_11766);
and U12169 (N_12169,N_11515,N_11613);
xor U12170 (N_12170,N_11571,N_11487);
xor U12171 (N_12171,N_11803,N_11506);
xnor U12172 (N_12172,N_11829,N_11738);
or U12173 (N_12173,N_11866,N_11574);
nand U12174 (N_12174,N_11314,N_11270);
or U12175 (N_12175,N_11528,N_11519);
nand U12176 (N_12176,N_11752,N_11856);
nand U12177 (N_12177,N_11697,N_11724);
and U12178 (N_12178,N_11860,N_11362);
nor U12179 (N_12179,N_11331,N_11332);
and U12180 (N_12180,N_11742,N_11440);
nand U12181 (N_12181,N_11453,N_11267);
xnor U12182 (N_12182,N_11433,N_11373);
nor U12183 (N_12183,N_11654,N_11348);
xor U12184 (N_12184,N_11660,N_11617);
and U12185 (N_12185,N_11776,N_11655);
and U12186 (N_12186,N_11389,N_11400);
and U12187 (N_12187,N_11765,N_11582);
xnor U12188 (N_12188,N_11556,N_11782);
nor U12189 (N_12189,N_11256,N_11331);
and U12190 (N_12190,N_11636,N_11622);
nand U12191 (N_12191,N_11461,N_11638);
xor U12192 (N_12192,N_11624,N_11860);
nor U12193 (N_12193,N_11499,N_11384);
or U12194 (N_12194,N_11790,N_11685);
nor U12195 (N_12195,N_11451,N_11493);
or U12196 (N_12196,N_11461,N_11559);
and U12197 (N_12197,N_11778,N_11838);
nor U12198 (N_12198,N_11639,N_11349);
and U12199 (N_12199,N_11421,N_11652);
xor U12200 (N_12200,N_11576,N_11698);
or U12201 (N_12201,N_11667,N_11466);
nor U12202 (N_12202,N_11278,N_11517);
or U12203 (N_12203,N_11657,N_11393);
xor U12204 (N_12204,N_11483,N_11366);
nand U12205 (N_12205,N_11498,N_11600);
or U12206 (N_12206,N_11808,N_11617);
and U12207 (N_12207,N_11826,N_11682);
nor U12208 (N_12208,N_11669,N_11705);
xnor U12209 (N_12209,N_11462,N_11437);
nor U12210 (N_12210,N_11741,N_11662);
nand U12211 (N_12211,N_11628,N_11767);
nand U12212 (N_12212,N_11383,N_11434);
xnor U12213 (N_12213,N_11409,N_11637);
nor U12214 (N_12214,N_11500,N_11509);
nand U12215 (N_12215,N_11867,N_11844);
and U12216 (N_12216,N_11412,N_11786);
nand U12217 (N_12217,N_11702,N_11521);
and U12218 (N_12218,N_11737,N_11369);
xnor U12219 (N_12219,N_11448,N_11284);
xnor U12220 (N_12220,N_11741,N_11432);
and U12221 (N_12221,N_11688,N_11550);
nor U12222 (N_12222,N_11735,N_11762);
xor U12223 (N_12223,N_11823,N_11541);
and U12224 (N_12224,N_11845,N_11516);
nand U12225 (N_12225,N_11786,N_11872);
nand U12226 (N_12226,N_11615,N_11412);
and U12227 (N_12227,N_11630,N_11825);
xnor U12228 (N_12228,N_11504,N_11309);
nand U12229 (N_12229,N_11456,N_11792);
xnor U12230 (N_12230,N_11828,N_11289);
nor U12231 (N_12231,N_11315,N_11693);
or U12232 (N_12232,N_11474,N_11764);
nor U12233 (N_12233,N_11389,N_11688);
or U12234 (N_12234,N_11471,N_11645);
and U12235 (N_12235,N_11368,N_11871);
nand U12236 (N_12236,N_11673,N_11683);
xnor U12237 (N_12237,N_11641,N_11565);
nor U12238 (N_12238,N_11388,N_11685);
or U12239 (N_12239,N_11452,N_11631);
nor U12240 (N_12240,N_11635,N_11646);
and U12241 (N_12241,N_11817,N_11417);
xnor U12242 (N_12242,N_11588,N_11526);
and U12243 (N_12243,N_11818,N_11611);
nand U12244 (N_12244,N_11341,N_11278);
and U12245 (N_12245,N_11670,N_11297);
or U12246 (N_12246,N_11603,N_11274);
nand U12247 (N_12247,N_11544,N_11385);
or U12248 (N_12248,N_11349,N_11722);
and U12249 (N_12249,N_11419,N_11340);
or U12250 (N_12250,N_11585,N_11349);
nand U12251 (N_12251,N_11491,N_11443);
nand U12252 (N_12252,N_11260,N_11450);
nand U12253 (N_12253,N_11478,N_11766);
or U12254 (N_12254,N_11574,N_11414);
nor U12255 (N_12255,N_11672,N_11874);
or U12256 (N_12256,N_11870,N_11450);
nand U12257 (N_12257,N_11649,N_11279);
or U12258 (N_12258,N_11490,N_11763);
nor U12259 (N_12259,N_11646,N_11582);
xnor U12260 (N_12260,N_11795,N_11469);
nor U12261 (N_12261,N_11841,N_11801);
xnor U12262 (N_12262,N_11420,N_11520);
nor U12263 (N_12263,N_11544,N_11680);
nand U12264 (N_12264,N_11468,N_11580);
nand U12265 (N_12265,N_11701,N_11804);
xnor U12266 (N_12266,N_11805,N_11708);
nor U12267 (N_12267,N_11637,N_11848);
and U12268 (N_12268,N_11355,N_11565);
nor U12269 (N_12269,N_11851,N_11443);
and U12270 (N_12270,N_11495,N_11285);
nand U12271 (N_12271,N_11846,N_11852);
or U12272 (N_12272,N_11657,N_11411);
nor U12273 (N_12273,N_11868,N_11293);
nor U12274 (N_12274,N_11599,N_11699);
xnor U12275 (N_12275,N_11399,N_11550);
xor U12276 (N_12276,N_11466,N_11403);
and U12277 (N_12277,N_11636,N_11646);
and U12278 (N_12278,N_11366,N_11859);
and U12279 (N_12279,N_11643,N_11588);
nor U12280 (N_12280,N_11688,N_11579);
xnor U12281 (N_12281,N_11490,N_11442);
nand U12282 (N_12282,N_11368,N_11747);
nand U12283 (N_12283,N_11777,N_11610);
nand U12284 (N_12284,N_11781,N_11461);
and U12285 (N_12285,N_11510,N_11273);
xor U12286 (N_12286,N_11310,N_11556);
and U12287 (N_12287,N_11742,N_11556);
nand U12288 (N_12288,N_11872,N_11541);
or U12289 (N_12289,N_11303,N_11816);
nand U12290 (N_12290,N_11487,N_11251);
and U12291 (N_12291,N_11409,N_11596);
nand U12292 (N_12292,N_11465,N_11540);
nand U12293 (N_12293,N_11472,N_11825);
and U12294 (N_12294,N_11739,N_11541);
or U12295 (N_12295,N_11428,N_11830);
nor U12296 (N_12296,N_11384,N_11526);
or U12297 (N_12297,N_11359,N_11317);
or U12298 (N_12298,N_11808,N_11341);
or U12299 (N_12299,N_11643,N_11626);
and U12300 (N_12300,N_11746,N_11422);
or U12301 (N_12301,N_11311,N_11524);
xor U12302 (N_12302,N_11613,N_11271);
xnor U12303 (N_12303,N_11731,N_11824);
xor U12304 (N_12304,N_11499,N_11699);
xor U12305 (N_12305,N_11400,N_11562);
xor U12306 (N_12306,N_11589,N_11453);
and U12307 (N_12307,N_11278,N_11378);
xnor U12308 (N_12308,N_11565,N_11683);
or U12309 (N_12309,N_11454,N_11577);
nand U12310 (N_12310,N_11610,N_11540);
nor U12311 (N_12311,N_11520,N_11614);
nand U12312 (N_12312,N_11391,N_11512);
nand U12313 (N_12313,N_11335,N_11373);
nand U12314 (N_12314,N_11748,N_11417);
xor U12315 (N_12315,N_11738,N_11661);
or U12316 (N_12316,N_11738,N_11692);
or U12317 (N_12317,N_11511,N_11279);
and U12318 (N_12318,N_11329,N_11524);
nand U12319 (N_12319,N_11522,N_11618);
and U12320 (N_12320,N_11423,N_11458);
xor U12321 (N_12321,N_11568,N_11521);
nor U12322 (N_12322,N_11720,N_11444);
nor U12323 (N_12323,N_11382,N_11577);
xnor U12324 (N_12324,N_11644,N_11343);
nor U12325 (N_12325,N_11670,N_11797);
or U12326 (N_12326,N_11475,N_11790);
xor U12327 (N_12327,N_11504,N_11460);
xnor U12328 (N_12328,N_11286,N_11474);
or U12329 (N_12329,N_11311,N_11345);
or U12330 (N_12330,N_11268,N_11569);
or U12331 (N_12331,N_11619,N_11341);
and U12332 (N_12332,N_11547,N_11714);
nand U12333 (N_12333,N_11704,N_11818);
xnor U12334 (N_12334,N_11517,N_11264);
xor U12335 (N_12335,N_11269,N_11387);
xnor U12336 (N_12336,N_11429,N_11760);
xnor U12337 (N_12337,N_11748,N_11446);
or U12338 (N_12338,N_11407,N_11624);
nand U12339 (N_12339,N_11521,N_11811);
nand U12340 (N_12340,N_11460,N_11463);
nand U12341 (N_12341,N_11386,N_11701);
or U12342 (N_12342,N_11713,N_11535);
or U12343 (N_12343,N_11766,N_11311);
nor U12344 (N_12344,N_11828,N_11263);
xnor U12345 (N_12345,N_11622,N_11274);
or U12346 (N_12346,N_11679,N_11470);
and U12347 (N_12347,N_11590,N_11441);
xnor U12348 (N_12348,N_11320,N_11536);
nor U12349 (N_12349,N_11446,N_11700);
nand U12350 (N_12350,N_11652,N_11681);
or U12351 (N_12351,N_11861,N_11290);
nand U12352 (N_12352,N_11600,N_11372);
and U12353 (N_12353,N_11505,N_11476);
nand U12354 (N_12354,N_11586,N_11780);
nand U12355 (N_12355,N_11566,N_11525);
xnor U12356 (N_12356,N_11340,N_11684);
or U12357 (N_12357,N_11801,N_11549);
and U12358 (N_12358,N_11750,N_11294);
nor U12359 (N_12359,N_11636,N_11695);
nand U12360 (N_12360,N_11800,N_11499);
nor U12361 (N_12361,N_11299,N_11531);
or U12362 (N_12362,N_11687,N_11392);
nor U12363 (N_12363,N_11834,N_11645);
and U12364 (N_12364,N_11691,N_11286);
nand U12365 (N_12365,N_11487,N_11320);
or U12366 (N_12366,N_11689,N_11417);
nand U12367 (N_12367,N_11745,N_11652);
nand U12368 (N_12368,N_11583,N_11342);
xor U12369 (N_12369,N_11534,N_11499);
or U12370 (N_12370,N_11391,N_11586);
nand U12371 (N_12371,N_11498,N_11606);
and U12372 (N_12372,N_11357,N_11856);
and U12373 (N_12373,N_11780,N_11862);
nand U12374 (N_12374,N_11815,N_11315);
nand U12375 (N_12375,N_11566,N_11582);
or U12376 (N_12376,N_11717,N_11301);
nand U12377 (N_12377,N_11345,N_11419);
or U12378 (N_12378,N_11758,N_11392);
or U12379 (N_12379,N_11431,N_11362);
nand U12380 (N_12380,N_11657,N_11374);
nor U12381 (N_12381,N_11532,N_11264);
xor U12382 (N_12382,N_11599,N_11355);
xnor U12383 (N_12383,N_11478,N_11291);
nor U12384 (N_12384,N_11288,N_11363);
xnor U12385 (N_12385,N_11462,N_11594);
xnor U12386 (N_12386,N_11867,N_11675);
nor U12387 (N_12387,N_11805,N_11807);
nand U12388 (N_12388,N_11418,N_11582);
xnor U12389 (N_12389,N_11499,N_11702);
and U12390 (N_12390,N_11415,N_11625);
or U12391 (N_12391,N_11561,N_11553);
nand U12392 (N_12392,N_11769,N_11570);
xor U12393 (N_12393,N_11596,N_11565);
xnor U12394 (N_12394,N_11410,N_11342);
xor U12395 (N_12395,N_11851,N_11287);
xnor U12396 (N_12396,N_11752,N_11341);
nor U12397 (N_12397,N_11745,N_11297);
and U12398 (N_12398,N_11664,N_11354);
and U12399 (N_12399,N_11584,N_11514);
or U12400 (N_12400,N_11699,N_11792);
nand U12401 (N_12401,N_11452,N_11834);
and U12402 (N_12402,N_11339,N_11456);
and U12403 (N_12403,N_11283,N_11744);
and U12404 (N_12404,N_11692,N_11304);
or U12405 (N_12405,N_11452,N_11425);
or U12406 (N_12406,N_11775,N_11588);
or U12407 (N_12407,N_11847,N_11556);
or U12408 (N_12408,N_11808,N_11631);
and U12409 (N_12409,N_11485,N_11801);
xnor U12410 (N_12410,N_11775,N_11474);
or U12411 (N_12411,N_11315,N_11817);
nand U12412 (N_12412,N_11757,N_11758);
nand U12413 (N_12413,N_11751,N_11633);
xor U12414 (N_12414,N_11772,N_11565);
xnor U12415 (N_12415,N_11607,N_11810);
or U12416 (N_12416,N_11562,N_11544);
and U12417 (N_12417,N_11464,N_11472);
nand U12418 (N_12418,N_11750,N_11598);
or U12419 (N_12419,N_11651,N_11784);
nand U12420 (N_12420,N_11539,N_11342);
or U12421 (N_12421,N_11608,N_11681);
nand U12422 (N_12422,N_11553,N_11510);
or U12423 (N_12423,N_11537,N_11354);
xor U12424 (N_12424,N_11870,N_11726);
nor U12425 (N_12425,N_11840,N_11553);
and U12426 (N_12426,N_11790,N_11745);
nand U12427 (N_12427,N_11337,N_11455);
nor U12428 (N_12428,N_11616,N_11844);
and U12429 (N_12429,N_11712,N_11540);
xnor U12430 (N_12430,N_11693,N_11866);
nand U12431 (N_12431,N_11410,N_11773);
nand U12432 (N_12432,N_11607,N_11742);
xnor U12433 (N_12433,N_11755,N_11662);
nand U12434 (N_12434,N_11705,N_11287);
xnor U12435 (N_12435,N_11394,N_11810);
or U12436 (N_12436,N_11418,N_11415);
or U12437 (N_12437,N_11688,N_11702);
or U12438 (N_12438,N_11345,N_11471);
or U12439 (N_12439,N_11811,N_11869);
or U12440 (N_12440,N_11351,N_11252);
nand U12441 (N_12441,N_11310,N_11684);
xnor U12442 (N_12442,N_11742,N_11274);
nand U12443 (N_12443,N_11318,N_11526);
or U12444 (N_12444,N_11453,N_11834);
xor U12445 (N_12445,N_11274,N_11564);
nor U12446 (N_12446,N_11442,N_11790);
nor U12447 (N_12447,N_11760,N_11828);
nor U12448 (N_12448,N_11504,N_11838);
nor U12449 (N_12449,N_11430,N_11313);
xor U12450 (N_12450,N_11420,N_11396);
and U12451 (N_12451,N_11296,N_11553);
nor U12452 (N_12452,N_11685,N_11312);
xnor U12453 (N_12453,N_11293,N_11283);
or U12454 (N_12454,N_11324,N_11753);
or U12455 (N_12455,N_11549,N_11509);
nand U12456 (N_12456,N_11252,N_11813);
xor U12457 (N_12457,N_11855,N_11374);
xnor U12458 (N_12458,N_11540,N_11673);
or U12459 (N_12459,N_11767,N_11572);
nor U12460 (N_12460,N_11372,N_11260);
or U12461 (N_12461,N_11860,N_11744);
xnor U12462 (N_12462,N_11416,N_11387);
or U12463 (N_12463,N_11688,N_11392);
and U12464 (N_12464,N_11585,N_11704);
nor U12465 (N_12465,N_11367,N_11740);
nand U12466 (N_12466,N_11486,N_11731);
xnor U12467 (N_12467,N_11756,N_11619);
nor U12468 (N_12468,N_11593,N_11355);
or U12469 (N_12469,N_11469,N_11799);
xor U12470 (N_12470,N_11770,N_11707);
xor U12471 (N_12471,N_11412,N_11482);
nand U12472 (N_12472,N_11740,N_11499);
nand U12473 (N_12473,N_11503,N_11469);
xor U12474 (N_12474,N_11670,N_11454);
nand U12475 (N_12475,N_11653,N_11480);
and U12476 (N_12476,N_11265,N_11554);
nand U12477 (N_12477,N_11690,N_11688);
and U12478 (N_12478,N_11665,N_11873);
or U12479 (N_12479,N_11475,N_11367);
xnor U12480 (N_12480,N_11405,N_11271);
nand U12481 (N_12481,N_11440,N_11543);
xnor U12482 (N_12482,N_11820,N_11614);
nand U12483 (N_12483,N_11482,N_11642);
nor U12484 (N_12484,N_11841,N_11611);
or U12485 (N_12485,N_11674,N_11788);
nand U12486 (N_12486,N_11261,N_11368);
xor U12487 (N_12487,N_11314,N_11642);
nand U12488 (N_12488,N_11392,N_11453);
xnor U12489 (N_12489,N_11541,N_11793);
or U12490 (N_12490,N_11656,N_11649);
nand U12491 (N_12491,N_11642,N_11342);
xnor U12492 (N_12492,N_11839,N_11852);
nor U12493 (N_12493,N_11465,N_11368);
nand U12494 (N_12494,N_11425,N_11556);
or U12495 (N_12495,N_11539,N_11485);
nor U12496 (N_12496,N_11660,N_11401);
nor U12497 (N_12497,N_11842,N_11777);
nor U12498 (N_12498,N_11419,N_11666);
nor U12499 (N_12499,N_11774,N_11553);
xor U12500 (N_12500,N_11930,N_12326);
and U12501 (N_12501,N_12309,N_12392);
nor U12502 (N_12502,N_12185,N_12340);
or U12503 (N_12503,N_12412,N_12076);
xor U12504 (N_12504,N_12409,N_12208);
xnor U12505 (N_12505,N_12329,N_12367);
nor U12506 (N_12506,N_12160,N_12399);
nor U12507 (N_12507,N_11959,N_12445);
nor U12508 (N_12508,N_12460,N_12043);
and U12509 (N_12509,N_12389,N_12463);
and U12510 (N_12510,N_12005,N_12475);
nand U12511 (N_12511,N_12453,N_11895);
xor U12512 (N_12512,N_12238,N_12250);
or U12513 (N_12513,N_12297,N_12162);
and U12514 (N_12514,N_11898,N_12133);
nor U12515 (N_12515,N_12210,N_12440);
and U12516 (N_12516,N_12322,N_11931);
xnor U12517 (N_12517,N_12016,N_12056);
xnor U12518 (N_12518,N_12293,N_12361);
xor U12519 (N_12519,N_12013,N_12189);
nand U12520 (N_12520,N_12469,N_12142);
xor U12521 (N_12521,N_11958,N_12441);
and U12522 (N_12522,N_12251,N_12486);
nor U12523 (N_12523,N_12490,N_11976);
and U12524 (N_12524,N_12258,N_12489);
nor U12525 (N_12525,N_11903,N_12304);
xor U12526 (N_12526,N_12324,N_12285);
or U12527 (N_12527,N_12333,N_12278);
and U12528 (N_12528,N_12176,N_12051);
nor U12529 (N_12529,N_12430,N_12194);
or U12530 (N_12530,N_12008,N_12306);
and U12531 (N_12531,N_12478,N_11975);
xnor U12532 (N_12532,N_12020,N_11884);
and U12533 (N_12533,N_12145,N_12281);
nand U12534 (N_12534,N_12003,N_11894);
or U12535 (N_12535,N_12091,N_11908);
xor U12536 (N_12536,N_12168,N_11902);
or U12537 (N_12537,N_12077,N_11955);
xor U12538 (N_12538,N_11879,N_12380);
and U12539 (N_12539,N_12066,N_11901);
or U12540 (N_12540,N_12071,N_12098);
nand U12541 (N_12541,N_12064,N_12063);
nand U12542 (N_12542,N_12332,N_12411);
xor U12543 (N_12543,N_12419,N_12230);
nor U12544 (N_12544,N_11915,N_12022);
xnor U12545 (N_12545,N_12213,N_12223);
xnor U12546 (N_12546,N_12196,N_12228);
nor U12547 (N_12547,N_12122,N_12180);
nand U12548 (N_12548,N_12347,N_12291);
nor U12549 (N_12549,N_12368,N_12294);
nand U12550 (N_12550,N_12439,N_12045);
xnor U12551 (N_12551,N_12165,N_12225);
or U12552 (N_12552,N_12061,N_12421);
and U12553 (N_12553,N_12334,N_12471);
xor U12554 (N_12554,N_11980,N_11921);
and U12555 (N_12555,N_12323,N_11998);
or U12556 (N_12556,N_11989,N_12179);
xnor U12557 (N_12557,N_12244,N_12277);
and U12558 (N_12558,N_11953,N_12127);
nor U12559 (N_12559,N_11964,N_12148);
or U12560 (N_12560,N_12204,N_12100);
nor U12561 (N_12561,N_12104,N_12152);
nand U12562 (N_12562,N_12195,N_12082);
xnor U12563 (N_12563,N_12090,N_12376);
nor U12564 (N_12564,N_12328,N_11887);
xor U12565 (N_12565,N_11918,N_12397);
xor U12566 (N_12566,N_12391,N_11912);
and U12567 (N_12567,N_12318,N_11994);
nor U12568 (N_12568,N_12079,N_12119);
xnor U12569 (N_12569,N_12164,N_12424);
nand U12570 (N_12570,N_12102,N_11897);
or U12571 (N_12571,N_12237,N_12470);
and U12572 (N_12572,N_11907,N_11965);
nand U12573 (N_12573,N_12214,N_12167);
nor U12574 (N_12574,N_12175,N_12089);
nor U12575 (N_12575,N_12492,N_12143);
or U12576 (N_12576,N_12386,N_12414);
and U12577 (N_12577,N_12209,N_11904);
and U12578 (N_12578,N_12394,N_12452);
or U12579 (N_12579,N_12117,N_12370);
nand U12580 (N_12580,N_11936,N_12290);
nor U12581 (N_12581,N_12353,N_11987);
nand U12582 (N_12582,N_12080,N_12062);
and U12583 (N_12583,N_11882,N_12074);
and U12584 (N_12584,N_12484,N_12203);
xnor U12585 (N_12585,N_11893,N_12288);
xor U12586 (N_12586,N_12136,N_12343);
and U12587 (N_12587,N_12435,N_12479);
nand U12588 (N_12588,N_12377,N_12495);
or U12589 (N_12589,N_11888,N_12444);
or U12590 (N_12590,N_11926,N_11962);
nor U12591 (N_12591,N_12171,N_12366);
and U12592 (N_12592,N_12023,N_11877);
and U12593 (N_12593,N_11927,N_12432);
and U12594 (N_12594,N_12425,N_12029);
nor U12595 (N_12595,N_12400,N_11974);
xor U12596 (N_12596,N_12241,N_12032);
nand U12597 (N_12597,N_12434,N_12103);
or U12598 (N_12598,N_11875,N_11956);
or U12599 (N_12599,N_12395,N_12357);
xor U12600 (N_12600,N_12216,N_12097);
nor U12601 (N_12601,N_12321,N_12027);
nand U12602 (N_12602,N_12011,N_11957);
xor U12603 (N_12603,N_12197,N_12450);
and U12604 (N_12604,N_12417,N_12438);
xor U12605 (N_12605,N_12387,N_12052);
nor U12606 (N_12606,N_12193,N_12497);
nor U12607 (N_12607,N_12087,N_12499);
nand U12608 (N_12608,N_12106,N_12068);
or U12609 (N_12609,N_12351,N_12256);
nand U12610 (N_12610,N_12099,N_12401);
and U12611 (N_12611,N_12153,N_12075);
and U12612 (N_12612,N_12243,N_12111);
nor U12613 (N_12613,N_12385,N_12408);
nor U12614 (N_12614,N_12156,N_12289);
nand U12615 (N_12615,N_12259,N_12163);
or U12616 (N_12616,N_11970,N_12363);
nor U12617 (N_12617,N_11944,N_12382);
nand U12618 (N_12618,N_12418,N_11981);
or U12619 (N_12619,N_12038,N_11885);
or U12620 (N_12620,N_12067,N_11977);
nand U12621 (N_12621,N_12224,N_12078);
or U12622 (N_12622,N_12229,N_11979);
xor U12623 (N_12623,N_12166,N_12252);
or U12624 (N_12624,N_12120,N_12423);
and U12625 (N_12625,N_11942,N_11978);
and U12626 (N_12626,N_12436,N_12406);
nand U12627 (N_12627,N_12384,N_12096);
nand U12628 (N_12628,N_12192,N_12447);
nand U12629 (N_12629,N_12126,N_12182);
nand U12630 (N_12630,N_12398,N_11947);
nor U12631 (N_12631,N_12232,N_12257);
and U12632 (N_12632,N_11941,N_12069);
and U12633 (N_12633,N_12480,N_12477);
and U12634 (N_12634,N_12174,N_12010);
nor U12635 (N_12635,N_12118,N_12327);
nor U12636 (N_12636,N_12365,N_12039);
or U12637 (N_12637,N_12085,N_12300);
or U12638 (N_12638,N_12443,N_11929);
or U12639 (N_12639,N_12275,N_11937);
xor U12640 (N_12640,N_12302,N_12217);
and U12641 (N_12641,N_12428,N_12320);
xnor U12642 (N_12642,N_12147,N_12049);
nand U12643 (N_12643,N_12132,N_12072);
nor U12644 (N_12644,N_11971,N_12170);
and U12645 (N_12645,N_11952,N_11945);
or U12646 (N_12646,N_12157,N_12220);
and U12647 (N_12647,N_12172,N_11909);
xor U12648 (N_12648,N_12420,N_11982);
xnor U12649 (N_12649,N_12042,N_12242);
nand U12650 (N_12650,N_12169,N_11892);
xnor U12651 (N_12651,N_12253,N_11896);
or U12652 (N_12652,N_12219,N_12007);
xnor U12653 (N_12653,N_12065,N_11911);
or U12654 (N_12654,N_12025,N_12422);
or U12655 (N_12655,N_12084,N_12303);
and U12656 (N_12656,N_12044,N_12338);
or U12657 (N_12657,N_12205,N_12383);
and U12658 (N_12658,N_11997,N_12186);
or U12659 (N_12659,N_12151,N_12141);
and U12660 (N_12660,N_11948,N_12449);
and U12661 (N_12661,N_12462,N_12108);
xor U12662 (N_12662,N_12105,N_11996);
nor U12663 (N_12663,N_12040,N_12249);
xnor U12664 (N_12664,N_12466,N_12234);
nor U12665 (N_12665,N_12266,N_12112);
and U12666 (N_12666,N_12159,N_12375);
or U12667 (N_12667,N_12131,N_12002);
nor U12668 (N_12668,N_11932,N_12222);
or U12669 (N_12669,N_12355,N_12437);
or U12670 (N_12670,N_12009,N_12155);
nor U12671 (N_12671,N_12483,N_12041);
and U12672 (N_12672,N_11920,N_12206);
nor U12673 (N_12673,N_12198,N_11969);
and U12674 (N_12674,N_11933,N_12456);
and U12675 (N_12675,N_12487,N_11990);
and U12676 (N_12676,N_12083,N_12073);
nand U12677 (N_12677,N_12388,N_12239);
nand U12678 (N_12678,N_11986,N_12468);
xor U12679 (N_12679,N_12012,N_12476);
and U12680 (N_12680,N_12431,N_12033);
xor U12681 (N_12681,N_12272,N_12378);
nand U12682 (N_12682,N_12298,N_12339);
nand U12683 (N_12683,N_11943,N_12121);
nand U12684 (N_12684,N_12092,N_11935);
nor U12685 (N_12685,N_12372,N_12371);
and U12686 (N_12686,N_12183,N_12413);
nor U12687 (N_12687,N_12050,N_12358);
nand U12688 (N_12688,N_11949,N_12070);
nor U12689 (N_12689,N_12130,N_12233);
and U12690 (N_12690,N_11972,N_12265);
nand U12691 (N_12691,N_12279,N_12267);
xor U12692 (N_12692,N_12352,N_12458);
and U12693 (N_12693,N_12493,N_12190);
nor U12694 (N_12694,N_12301,N_11928);
nor U12695 (N_12695,N_12429,N_11881);
and U12696 (N_12696,N_12218,N_12396);
nor U12697 (N_12697,N_11924,N_12086);
nor U12698 (N_12698,N_12402,N_12260);
and U12699 (N_12699,N_11914,N_12240);
nand U12700 (N_12700,N_12114,N_12261);
xor U12701 (N_12701,N_12004,N_11954);
and U12702 (N_12702,N_12405,N_12331);
nand U12703 (N_12703,N_12247,N_12047);
nor U12704 (N_12704,N_12128,N_12015);
nand U12705 (N_12705,N_12416,N_12137);
nand U12706 (N_12706,N_12379,N_12173);
nor U12707 (N_12707,N_12482,N_12360);
and U12708 (N_12708,N_11922,N_12390);
xnor U12709 (N_12709,N_12348,N_11876);
nor U12710 (N_12710,N_11992,N_12124);
and U12711 (N_12711,N_12188,N_12088);
and U12712 (N_12712,N_11991,N_12054);
or U12713 (N_12713,N_12410,N_12354);
xnor U12714 (N_12714,N_12000,N_11984);
nor U12715 (N_12715,N_12433,N_12337);
and U12716 (N_12716,N_12280,N_12021);
or U12717 (N_12717,N_11913,N_12319);
nand U12718 (N_12718,N_12415,N_12427);
or U12719 (N_12719,N_12349,N_12317);
xor U12720 (N_12720,N_12274,N_12109);
or U12721 (N_12721,N_12307,N_12231);
nand U12722 (N_12722,N_12215,N_11999);
nor U12723 (N_12723,N_12123,N_12227);
or U12724 (N_12724,N_12393,N_12036);
or U12725 (N_12725,N_11917,N_12006);
xnor U12726 (N_12726,N_11940,N_12454);
nor U12727 (N_12727,N_12161,N_12212);
nand U12728 (N_12728,N_12053,N_12467);
nor U12729 (N_12729,N_11900,N_12094);
nor U12730 (N_12730,N_12113,N_12026);
and U12731 (N_12731,N_12017,N_12146);
or U12732 (N_12732,N_12191,N_12001);
and U12733 (N_12733,N_11899,N_12426);
nor U12734 (N_12734,N_12035,N_12364);
nand U12735 (N_12735,N_11938,N_11963);
or U12736 (N_12736,N_12150,N_11946);
xnor U12737 (N_12737,N_12181,N_12448);
nor U12738 (N_12738,N_12014,N_12060);
nor U12739 (N_12739,N_12115,N_12138);
and U12740 (N_12740,N_12403,N_11995);
and U12741 (N_12741,N_12407,N_12286);
nand U12742 (N_12742,N_12442,N_12313);
and U12743 (N_12743,N_12201,N_12095);
and U12744 (N_12744,N_12158,N_12135);
or U12745 (N_12745,N_12465,N_12451);
nand U12746 (N_12746,N_12263,N_11910);
and U12747 (N_12747,N_12494,N_11878);
nand U12748 (N_12748,N_11890,N_11906);
or U12749 (N_12749,N_12177,N_11916);
or U12750 (N_12750,N_12144,N_12236);
nor U12751 (N_12751,N_12312,N_12046);
and U12752 (N_12752,N_12374,N_12474);
nor U12753 (N_12753,N_12200,N_12129);
nor U12754 (N_12754,N_12211,N_11960);
nand U12755 (N_12755,N_12481,N_12305);
nand U12756 (N_12756,N_12140,N_12154);
or U12757 (N_12757,N_12316,N_11968);
and U12758 (N_12758,N_12270,N_11880);
nor U12759 (N_12759,N_11939,N_11891);
and U12760 (N_12760,N_11988,N_12283);
xor U12761 (N_12761,N_12292,N_12255);
and U12762 (N_12762,N_11889,N_12359);
or U12763 (N_12763,N_12055,N_12308);
xor U12764 (N_12764,N_12335,N_12264);
nor U12765 (N_12765,N_12187,N_12342);
nand U12766 (N_12766,N_12498,N_12110);
nand U12767 (N_12767,N_12221,N_12116);
nor U12768 (N_12768,N_12184,N_12245);
nand U12769 (N_12769,N_12296,N_11966);
or U12770 (N_12770,N_12101,N_12031);
and U12771 (N_12771,N_12282,N_12344);
nand U12772 (N_12772,N_12310,N_12457);
and U12773 (N_12773,N_11973,N_12488);
or U12774 (N_12774,N_12246,N_12341);
nand U12775 (N_12775,N_12134,N_12149);
xnor U12776 (N_12776,N_11886,N_12314);
and U12777 (N_12777,N_12273,N_12018);
or U12778 (N_12778,N_11983,N_12325);
xor U12779 (N_12779,N_12350,N_12464);
nand U12780 (N_12780,N_12081,N_12373);
xor U12781 (N_12781,N_12269,N_12330);
nand U12782 (N_12782,N_12235,N_12381);
nand U12783 (N_12783,N_12248,N_12485);
xnor U12784 (N_12784,N_12028,N_12139);
nor U12785 (N_12785,N_11993,N_12276);
xor U12786 (N_12786,N_12496,N_12059);
nand U12787 (N_12787,N_12207,N_11967);
nand U12788 (N_12788,N_12295,N_12346);
xor U12789 (N_12789,N_12315,N_12491);
nand U12790 (N_12790,N_12369,N_11985);
or U12791 (N_12791,N_12019,N_12362);
nor U12792 (N_12792,N_12459,N_12461);
or U12793 (N_12793,N_11961,N_12125);
nand U12794 (N_12794,N_11951,N_12345);
xor U12795 (N_12795,N_12446,N_11905);
and U12796 (N_12796,N_12178,N_12268);
or U12797 (N_12797,N_12254,N_12311);
and U12798 (N_12798,N_12262,N_12299);
nor U12799 (N_12799,N_12336,N_12226);
xnor U12800 (N_12800,N_12202,N_12024);
xor U12801 (N_12801,N_11883,N_12037);
or U12802 (N_12802,N_12455,N_11923);
and U12803 (N_12803,N_12271,N_11950);
nand U12804 (N_12804,N_12404,N_12093);
nor U12805 (N_12805,N_12057,N_12287);
nand U12806 (N_12806,N_12356,N_12058);
nor U12807 (N_12807,N_12472,N_11925);
xor U12808 (N_12808,N_12034,N_12284);
or U12809 (N_12809,N_12107,N_12030);
nand U12810 (N_12810,N_11934,N_11919);
xnor U12811 (N_12811,N_12048,N_12199);
nand U12812 (N_12812,N_12473,N_12030);
nor U12813 (N_12813,N_12102,N_12001);
and U12814 (N_12814,N_12155,N_12427);
nor U12815 (N_12815,N_11904,N_11907);
nand U12816 (N_12816,N_12111,N_11890);
nand U12817 (N_12817,N_12450,N_12393);
nand U12818 (N_12818,N_12124,N_12046);
nand U12819 (N_12819,N_12269,N_12215);
and U12820 (N_12820,N_12104,N_12012);
xnor U12821 (N_12821,N_12379,N_11922);
and U12822 (N_12822,N_11934,N_12277);
nand U12823 (N_12823,N_12438,N_11904);
or U12824 (N_12824,N_12071,N_11878);
xor U12825 (N_12825,N_11985,N_12321);
xnor U12826 (N_12826,N_12214,N_12215);
xor U12827 (N_12827,N_12437,N_12341);
and U12828 (N_12828,N_12271,N_12023);
and U12829 (N_12829,N_11986,N_12160);
or U12830 (N_12830,N_12222,N_11936);
nand U12831 (N_12831,N_12057,N_12168);
xnor U12832 (N_12832,N_11960,N_12486);
and U12833 (N_12833,N_11994,N_11885);
xnor U12834 (N_12834,N_12359,N_12097);
or U12835 (N_12835,N_12252,N_12083);
and U12836 (N_12836,N_12237,N_12212);
or U12837 (N_12837,N_12192,N_12345);
xor U12838 (N_12838,N_11950,N_12010);
or U12839 (N_12839,N_12135,N_11901);
xor U12840 (N_12840,N_12385,N_12047);
nand U12841 (N_12841,N_12116,N_12126);
and U12842 (N_12842,N_12455,N_12313);
nor U12843 (N_12843,N_12132,N_12091);
or U12844 (N_12844,N_12078,N_12368);
nand U12845 (N_12845,N_12387,N_12131);
nor U12846 (N_12846,N_11930,N_12418);
xnor U12847 (N_12847,N_11931,N_12381);
nand U12848 (N_12848,N_12425,N_12218);
xor U12849 (N_12849,N_12433,N_12469);
nand U12850 (N_12850,N_12421,N_12463);
nor U12851 (N_12851,N_12446,N_12250);
or U12852 (N_12852,N_12215,N_12302);
nor U12853 (N_12853,N_11887,N_12008);
xnor U12854 (N_12854,N_12487,N_12418);
or U12855 (N_12855,N_12038,N_11968);
and U12856 (N_12856,N_12104,N_12249);
nand U12857 (N_12857,N_12227,N_11905);
nor U12858 (N_12858,N_12037,N_12269);
xnor U12859 (N_12859,N_12463,N_12273);
xor U12860 (N_12860,N_12278,N_12499);
nor U12861 (N_12861,N_12036,N_12474);
or U12862 (N_12862,N_12383,N_12390);
or U12863 (N_12863,N_12479,N_11976);
and U12864 (N_12864,N_12323,N_12176);
and U12865 (N_12865,N_12195,N_12443);
nor U12866 (N_12866,N_11902,N_11946);
nand U12867 (N_12867,N_12289,N_11974);
xor U12868 (N_12868,N_12022,N_12438);
nor U12869 (N_12869,N_12114,N_12154);
and U12870 (N_12870,N_12201,N_12312);
nand U12871 (N_12871,N_12025,N_12031);
xor U12872 (N_12872,N_12093,N_12250);
nor U12873 (N_12873,N_12118,N_12344);
nor U12874 (N_12874,N_11927,N_12124);
nor U12875 (N_12875,N_12017,N_12108);
and U12876 (N_12876,N_11971,N_12338);
and U12877 (N_12877,N_12379,N_11994);
nor U12878 (N_12878,N_12226,N_11992);
nor U12879 (N_12879,N_11944,N_12170);
nor U12880 (N_12880,N_11921,N_11968);
nand U12881 (N_12881,N_12038,N_12143);
nand U12882 (N_12882,N_12192,N_12474);
nor U12883 (N_12883,N_12000,N_12454);
and U12884 (N_12884,N_12384,N_12360);
or U12885 (N_12885,N_12328,N_11962);
xor U12886 (N_12886,N_12491,N_12263);
or U12887 (N_12887,N_12187,N_12268);
nor U12888 (N_12888,N_11924,N_12478);
or U12889 (N_12889,N_11887,N_12091);
or U12890 (N_12890,N_12426,N_12383);
xor U12891 (N_12891,N_12099,N_12314);
nor U12892 (N_12892,N_12488,N_12293);
xor U12893 (N_12893,N_12157,N_12386);
nand U12894 (N_12894,N_12086,N_12417);
xor U12895 (N_12895,N_12374,N_12244);
nor U12896 (N_12896,N_12348,N_12094);
nor U12897 (N_12897,N_12246,N_12184);
nor U12898 (N_12898,N_12038,N_12127);
nand U12899 (N_12899,N_11890,N_11915);
nor U12900 (N_12900,N_12075,N_12474);
nand U12901 (N_12901,N_11997,N_12086);
or U12902 (N_12902,N_12305,N_12345);
xnor U12903 (N_12903,N_11878,N_12057);
and U12904 (N_12904,N_11912,N_12211);
nor U12905 (N_12905,N_11942,N_12001);
or U12906 (N_12906,N_12175,N_12342);
nor U12907 (N_12907,N_12110,N_11946);
nand U12908 (N_12908,N_12212,N_12479);
nor U12909 (N_12909,N_12211,N_12194);
or U12910 (N_12910,N_12022,N_12175);
and U12911 (N_12911,N_12121,N_12395);
nor U12912 (N_12912,N_12069,N_12363);
xnor U12913 (N_12913,N_12172,N_12146);
xnor U12914 (N_12914,N_12181,N_12280);
nor U12915 (N_12915,N_12325,N_12099);
xnor U12916 (N_12916,N_12469,N_12345);
or U12917 (N_12917,N_12156,N_11917);
nand U12918 (N_12918,N_12477,N_12145);
nor U12919 (N_12919,N_11887,N_12242);
or U12920 (N_12920,N_12089,N_11935);
or U12921 (N_12921,N_12278,N_12033);
or U12922 (N_12922,N_11991,N_11915);
and U12923 (N_12923,N_12140,N_11896);
nor U12924 (N_12924,N_12175,N_12158);
and U12925 (N_12925,N_12404,N_12248);
xor U12926 (N_12926,N_12220,N_12173);
or U12927 (N_12927,N_12208,N_12141);
nor U12928 (N_12928,N_11884,N_12402);
nand U12929 (N_12929,N_11965,N_12159);
and U12930 (N_12930,N_12091,N_11972);
nor U12931 (N_12931,N_12273,N_12361);
nand U12932 (N_12932,N_12134,N_12155);
nor U12933 (N_12933,N_12406,N_12084);
or U12934 (N_12934,N_11920,N_12421);
or U12935 (N_12935,N_12045,N_12237);
nor U12936 (N_12936,N_12216,N_12193);
nor U12937 (N_12937,N_12093,N_12201);
nand U12938 (N_12938,N_12001,N_12012);
nor U12939 (N_12939,N_11942,N_12143);
nand U12940 (N_12940,N_12080,N_12196);
nand U12941 (N_12941,N_12413,N_12485);
xnor U12942 (N_12942,N_12432,N_12358);
xor U12943 (N_12943,N_12302,N_12360);
nand U12944 (N_12944,N_11931,N_12404);
and U12945 (N_12945,N_12260,N_12361);
xnor U12946 (N_12946,N_12077,N_12165);
or U12947 (N_12947,N_11985,N_12015);
and U12948 (N_12948,N_12153,N_12027);
and U12949 (N_12949,N_12261,N_12162);
nand U12950 (N_12950,N_12286,N_11993);
xor U12951 (N_12951,N_12309,N_12084);
or U12952 (N_12952,N_12223,N_11939);
nand U12953 (N_12953,N_12227,N_12225);
or U12954 (N_12954,N_12112,N_12338);
and U12955 (N_12955,N_12105,N_12338);
and U12956 (N_12956,N_12391,N_11984);
or U12957 (N_12957,N_12367,N_12423);
nand U12958 (N_12958,N_11956,N_11982);
nor U12959 (N_12959,N_12320,N_12314);
xor U12960 (N_12960,N_12208,N_12385);
and U12961 (N_12961,N_12025,N_11996);
or U12962 (N_12962,N_12202,N_12463);
nor U12963 (N_12963,N_12432,N_12488);
xor U12964 (N_12964,N_11945,N_12495);
or U12965 (N_12965,N_11922,N_12248);
nand U12966 (N_12966,N_12332,N_12176);
nand U12967 (N_12967,N_11926,N_12409);
nor U12968 (N_12968,N_11912,N_11971);
xor U12969 (N_12969,N_12444,N_12170);
or U12970 (N_12970,N_12478,N_12424);
or U12971 (N_12971,N_11878,N_12400);
xor U12972 (N_12972,N_12420,N_12406);
nand U12973 (N_12973,N_12400,N_12061);
nor U12974 (N_12974,N_12340,N_12241);
and U12975 (N_12975,N_12494,N_12130);
and U12976 (N_12976,N_11988,N_12334);
nor U12977 (N_12977,N_12155,N_12441);
or U12978 (N_12978,N_12004,N_12086);
xor U12979 (N_12979,N_12003,N_12371);
nor U12980 (N_12980,N_12061,N_12166);
and U12981 (N_12981,N_12343,N_12032);
nor U12982 (N_12982,N_12187,N_12215);
and U12983 (N_12983,N_12406,N_11958);
or U12984 (N_12984,N_11932,N_12269);
or U12985 (N_12985,N_11951,N_11964);
xor U12986 (N_12986,N_12167,N_12324);
nor U12987 (N_12987,N_12009,N_11927);
and U12988 (N_12988,N_12244,N_12140);
nand U12989 (N_12989,N_12306,N_12072);
nor U12990 (N_12990,N_12406,N_11982);
nor U12991 (N_12991,N_12054,N_12092);
and U12992 (N_12992,N_12238,N_12171);
nor U12993 (N_12993,N_12418,N_12387);
nor U12994 (N_12994,N_11947,N_12396);
and U12995 (N_12995,N_11880,N_12129);
or U12996 (N_12996,N_12144,N_12189);
nand U12997 (N_12997,N_12101,N_12146);
xnor U12998 (N_12998,N_11964,N_12303);
or U12999 (N_12999,N_12049,N_12270);
nor U13000 (N_13000,N_12227,N_12264);
nor U13001 (N_13001,N_11929,N_12010);
nand U13002 (N_13002,N_12346,N_12261);
or U13003 (N_13003,N_12072,N_12163);
nand U13004 (N_13004,N_12459,N_12003);
xnor U13005 (N_13005,N_12103,N_12417);
nor U13006 (N_13006,N_12101,N_12166);
nand U13007 (N_13007,N_12053,N_12396);
and U13008 (N_13008,N_12273,N_12406);
nor U13009 (N_13009,N_12144,N_12475);
and U13010 (N_13010,N_12432,N_12163);
nor U13011 (N_13011,N_12254,N_12225);
and U13012 (N_13012,N_11886,N_12360);
and U13013 (N_13013,N_12231,N_12415);
or U13014 (N_13014,N_11969,N_12168);
xor U13015 (N_13015,N_11906,N_12358);
or U13016 (N_13016,N_12120,N_11935);
xor U13017 (N_13017,N_12173,N_12116);
nor U13018 (N_13018,N_12318,N_12391);
and U13019 (N_13019,N_12355,N_12221);
xnor U13020 (N_13020,N_12409,N_12077);
nand U13021 (N_13021,N_12046,N_11990);
and U13022 (N_13022,N_12257,N_12266);
or U13023 (N_13023,N_11982,N_11888);
nand U13024 (N_13024,N_12411,N_12242);
xor U13025 (N_13025,N_12081,N_11906);
nor U13026 (N_13026,N_12118,N_11994);
nand U13027 (N_13027,N_11917,N_12033);
xor U13028 (N_13028,N_12302,N_12179);
nor U13029 (N_13029,N_12171,N_11973);
or U13030 (N_13030,N_12045,N_11983);
xor U13031 (N_13031,N_12438,N_12157);
nor U13032 (N_13032,N_11966,N_11885);
xor U13033 (N_13033,N_12491,N_12049);
xor U13034 (N_13034,N_11954,N_12003);
nor U13035 (N_13035,N_12492,N_12443);
xor U13036 (N_13036,N_12499,N_12153);
nor U13037 (N_13037,N_12112,N_12193);
nor U13038 (N_13038,N_12149,N_12380);
xnor U13039 (N_13039,N_12162,N_12093);
and U13040 (N_13040,N_12037,N_11940);
nand U13041 (N_13041,N_11942,N_12197);
nand U13042 (N_13042,N_12121,N_12095);
or U13043 (N_13043,N_12198,N_11901);
and U13044 (N_13044,N_12304,N_12263);
nand U13045 (N_13045,N_12111,N_12266);
or U13046 (N_13046,N_12016,N_12229);
or U13047 (N_13047,N_11988,N_12256);
xnor U13048 (N_13048,N_12079,N_11978);
or U13049 (N_13049,N_11956,N_12084);
xnor U13050 (N_13050,N_12468,N_12160);
nand U13051 (N_13051,N_12168,N_12154);
nand U13052 (N_13052,N_12110,N_12182);
nor U13053 (N_13053,N_11949,N_12388);
nand U13054 (N_13054,N_12276,N_12173);
nor U13055 (N_13055,N_11915,N_12329);
or U13056 (N_13056,N_12333,N_12355);
and U13057 (N_13057,N_12339,N_12175);
nor U13058 (N_13058,N_12239,N_12123);
and U13059 (N_13059,N_12337,N_12115);
xnor U13060 (N_13060,N_12226,N_11995);
xor U13061 (N_13061,N_11897,N_11949);
or U13062 (N_13062,N_12108,N_12302);
and U13063 (N_13063,N_12364,N_12135);
nand U13064 (N_13064,N_12422,N_12355);
nand U13065 (N_13065,N_12249,N_12349);
or U13066 (N_13066,N_12054,N_12259);
or U13067 (N_13067,N_12081,N_12367);
or U13068 (N_13068,N_11879,N_11878);
nor U13069 (N_13069,N_12185,N_12320);
or U13070 (N_13070,N_12075,N_12364);
nor U13071 (N_13071,N_12151,N_12204);
nand U13072 (N_13072,N_12035,N_12399);
xnor U13073 (N_13073,N_12120,N_12069);
nor U13074 (N_13074,N_12441,N_11935);
nand U13075 (N_13075,N_12334,N_12220);
nand U13076 (N_13076,N_11884,N_12044);
or U13077 (N_13077,N_12320,N_12369);
xor U13078 (N_13078,N_12075,N_12289);
xnor U13079 (N_13079,N_12084,N_12447);
nor U13080 (N_13080,N_11904,N_12380);
or U13081 (N_13081,N_12420,N_11984);
xor U13082 (N_13082,N_12358,N_12308);
nand U13083 (N_13083,N_12162,N_11897);
or U13084 (N_13084,N_12452,N_12211);
and U13085 (N_13085,N_12196,N_12499);
or U13086 (N_13086,N_12399,N_12379);
or U13087 (N_13087,N_11917,N_12435);
nand U13088 (N_13088,N_12276,N_12091);
nand U13089 (N_13089,N_11895,N_12178);
and U13090 (N_13090,N_12311,N_12467);
and U13091 (N_13091,N_12099,N_12079);
xnor U13092 (N_13092,N_12339,N_12361);
and U13093 (N_13093,N_12176,N_12077);
nand U13094 (N_13094,N_12338,N_12089);
nor U13095 (N_13095,N_11977,N_12095);
and U13096 (N_13096,N_12492,N_12270);
xor U13097 (N_13097,N_12487,N_12261);
and U13098 (N_13098,N_12192,N_12454);
and U13099 (N_13099,N_12463,N_12013);
and U13100 (N_13100,N_12101,N_12412);
nand U13101 (N_13101,N_11982,N_12324);
nor U13102 (N_13102,N_12252,N_12114);
nor U13103 (N_13103,N_12165,N_11980);
and U13104 (N_13104,N_12236,N_11960);
nand U13105 (N_13105,N_12240,N_12393);
nand U13106 (N_13106,N_11975,N_12165);
nand U13107 (N_13107,N_12446,N_12268);
or U13108 (N_13108,N_12367,N_12364);
or U13109 (N_13109,N_12234,N_12345);
or U13110 (N_13110,N_12351,N_12426);
xor U13111 (N_13111,N_12258,N_11910);
nor U13112 (N_13112,N_12332,N_11991);
and U13113 (N_13113,N_12252,N_12289);
nand U13114 (N_13114,N_11895,N_12054);
and U13115 (N_13115,N_12276,N_12185);
and U13116 (N_13116,N_12239,N_12494);
or U13117 (N_13117,N_11943,N_12127);
xnor U13118 (N_13118,N_12033,N_12114);
nand U13119 (N_13119,N_12083,N_11911);
nor U13120 (N_13120,N_12217,N_12481);
or U13121 (N_13121,N_12319,N_12367);
and U13122 (N_13122,N_11980,N_11934);
nand U13123 (N_13123,N_12215,N_11981);
and U13124 (N_13124,N_12129,N_12274);
nand U13125 (N_13125,N_13025,N_12844);
or U13126 (N_13126,N_12803,N_12589);
xor U13127 (N_13127,N_12945,N_12779);
and U13128 (N_13128,N_13090,N_12969);
xnor U13129 (N_13129,N_12532,N_12656);
or U13130 (N_13130,N_13087,N_12591);
and U13131 (N_13131,N_13110,N_12903);
xnor U13132 (N_13132,N_12511,N_12713);
nor U13133 (N_13133,N_12520,N_12936);
nand U13134 (N_13134,N_13084,N_12916);
nand U13135 (N_13135,N_12515,N_13053);
xnor U13136 (N_13136,N_13014,N_12841);
or U13137 (N_13137,N_13062,N_12576);
and U13138 (N_13138,N_12724,N_12551);
and U13139 (N_13139,N_13052,N_12715);
nand U13140 (N_13140,N_12813,N_12788);
and U13141 (N_13141,N_12906,N_13109);
or U13142 (N_13142,N_12896,N_12653);
nor U13143 (N_13143,N_12765,N_12990);
xnor U13144 (N_13144,N_12766,N_12710);
nor U13145 (N_13145,N_13124,N_12840);
nor U13146 (N_13146,N_12633,N_12654);
nor U13147 (N_13147,N_12745,N_12519);
or U13148 (N_13148,N_13101,N_12821);
xnor U13149 (N_13149,N_13032,N_12899);
nand U13150 (N_13150,N_13107,N_12608);
or U13151 (N_13151,N_12791,N_12742);
nand U13152 (N_13152,N_13082,N_12802);
nor U13153 (N_13153,N_12577,N_12627);
nand U13154 (N_13154,N_12749,N_13008);
nor U13155 (N_13155,N_12826,N_13022);
xnor U13156 (N_13156,N_12734,N_13013);
xor U13157 (N_13157,N_12770,N_12865);
xnor U13158 (N_13158,N_12513,N_12685);
xor U13159 (N_13159,N_12946,N_12582);
xnor U13160 (N_13160,N_12890,N_12683);
xor U13161 (N_13161,N_12668,N_12951);
nor U13162 (N_13162,N_13113,N_13118);
xnor U13163 (N_13163,N_12509,N_13075);
nand U13164 (N_13164,N_13058,N_13065);
or U13165 (N_13165,N_12883,N_12535);
and U13166 (N_13166,N_12774,N_12988);
nand U13167 (N_13167,N_12763,N_12941);
nand U13168 (N_13168,N_12772,N_12508);
nand U13169 (N_13169,N_12722,N_12987);
or U13170 (N_13170,N_12950,N_12503);
and U13171 (N_13171,N_13044,N_12610);
nor U13172 (N_13172,N_12973,N_12557);
nand U13173 (N_13173,N_13046,N_12548);
or U13174 (N_13174,N_12614,N_12693);
nand U13175 (N_13175,N_12971,N_13059);
or U13176 (N_13176,N_13045,N_13070);
xor U13177 (N_13177,N_13097,N_12856);
or U13178 (N_13178,N_12561,N_12963);
nand U13179 (N_13179,N_12609,N_12905);
nor U13180 (N_13180,N_12790,N_12613);
or U13181 (N_13181,N_12599,N_13120);
nor U13182 (N_13182,N_12932,N_12898);
or U13183 (N_13183,N_13011,N_13068);
nor U13184 (N_13184,N_12706,N_12921);
xnor U13185 (N_13185,N_12611,N_12913);
nor U13186 (N_13186,N_12578,N_12678);
nand U13187 (N_13187,N_12984,N_12544);
or U13188 (N_13188,N_12825,N_12979);
and U13189 (N_13189,N_12965,N_12934);
or U13190 (N_13190,N_12670,N_12731);
and U13191 (N_13191,N_12564,N_12690);
nand U13192 (N_13192,N_13104,N_13081);
nand U13193 (N_13193,N_12838,N_12510);
nand U13194 (N_13194,N_12638,N_12581);
nand U13195 (N_13195,N_12721,N_12504);
and U13196 (N_13196,N_13023,N_12902);
or U13197 (N_13197,N_12618,N_12874);
or U13198 (N_13198,N_12789,N_12639);
nand U13199 (N_13199,N_13050,N_12809);
nor U13200 (N_13200,N_12775,N_12716);
nor U13201 (N_13201,N_13064,N_13095);
nor U13202 (N_13202,N_12933,N_12605);
xor U13203 (N_13203,N_12691,N_12681);
and U13204 (N_13204,N_12636,N_13092);
nand U13205 (N_13205,N_12637,N_12806);
xnor U13206 (N_13206,N_13063,N_12760);
or U13207 (N_13207,N_12632,N_12980);
xor U13208 (N_13208,N_12518,N_12938);
xor U13209 (N_13209,N_12918,N_12660);
and U13210 (N_13210,N_13005,N_12817);
nand U13211 (N_13211,N_12908,N_12620);
nor U13212 (N_13212,N_12995,N_12805);
and U13213 (N_13213,N_12640,N_12996);
or U13214 (N_13214,N_12960,N_12646);
or U13215 (N_13215,N_13004,N_12725);
and U13216 (N_13216,N_12781,N_12870);
and U13217 (N_13217,N_12617,N_12730);
nor U13218 (N_13218,N_12523,N_13091);
xnor U13219 (N_13219,N_12753,N_13074);
xor U13220 (N_13220,N_12924,N_12621);
nor U13221 (N_13221,N_12699,N_12642);
and U13222 (N_13222,N_12955,N_12850);
xnor U13223 (N_13223,N_12993,N_12502);
nor U13224 (N_13224,N_12616,N_12507);
nor U13225 (N_13225,N_12784,N_12815);
xor U13226 (N_13226,N_12956,N_13027);
or U13227 (N_13227,N_12748,N_12857);
and U13228 (N_13228,N_12831,N_12836);
or U13229 (N_13229,N_12859,N_12889);
nand U13230 (N_13230,N_12694,N_12601);
or U13231 (N_13231,N_12922,N_12628);
xor U13232 (N_13232,N_13105,N_12701);
nor U13233 (N_13233,N_12901,N_12667);
or U13234 (N_13234,N_13039,N_12600);
nor U13235 (N_13235,N_13057,N_12759);
nor U13236 (N_13236,N_13094,N_12580);
nand U13237 (N_13237,N_12675,N_12674);
nand U13238 (N_13238,N_13029,N_12568);
xnor U13239 (N_13239,N_13021,N_12992);
nand U13240 (N_13240,N_12529,N_12545);
xor U13241 (N_13241,N_12506,N_12500);
xor U13242 (N_13242,N_13038,N_12572);
and U13243 (N_13243,N_12538,N_12891);
nand U13244 (N_13244,N_12739,N_12727);
xor U13245 (N_13245,N_12937,N_12735);
and U13246 (N_13246,N_13069,N_12861);
nand U13247 (N_13247,N_12834,N_13028);
nor U13248 (N_13248,N_12782,N_12758);
nand U13249 (N_13249,N_12944,N_13106);
or U13250 (N_13250,N_12931,N_13103);
nor U13251 (N_13251,N_12798,N_13085);
nor U13252 (N_13252,N_12754,N_12909);
nor U13253 (N_13253,N_12968,N_12869);
nor U13254 (N_13254,N_12663,N_13119);
nor U13255 (N_13255,N_12530,N_12575);
or U13256 (N_13256,N_13009,N_12569);
nand U13257 (N_13257,N_12741,N_12839);
and U13258 (N_13258,N_12935,N_12652);
and U13259 (N_13259,N_12867,N_12875);
xnor U13260 (N_13260,N_13037,N_12723);
nand U13261 (N_13261,N_12705,N_12737);
nor U13262 (N_13262,N_12863,N_12573);
and U13263 (N_13263,N_12682,N_12594);
nor U13264 (N_13264,N_12787,N_12923);
or U13265 (N_13265,N_12837,N_12711);
nor U13266 (N_13266,N_12688,N_12743);
xor U13267 (N_13267,N_12738,N_12846);
or U13268 (N_13268,N_12647,N_12583);
and U13269 (N_13269,N_12952,N_13066);
nor U13270 (N_13270,N_12804,N_13010);
or U13271 (N_13271,N_12824,N_12720);
nor U13272 (N_13272,N_12943,N_13018);
nand U13273 (N_13273,N_12534,N_12827);
or U13274 (N_13274,N_12847,N_12851);
nor U13275 (N_13275,N_12686,N_12574);
and U13276 (N_13276,N_12989,N_12877);
xnor U13277 (N_13277,N_12894,N_12566);
nor U13278 (N_13278,N_12658,N_13076);
nand U13279 (N_13279,N_12907,N_13089);
nor U13280 (N_13280,N_12926,N_12887);
nand U13281 (N_13281,N_13048,N_12974);
or U13282 (N_13282,N_13002,N_12929);
or U13283 (N_13283,N_13054,N_12631);
nor U13284 (N_13284,N_12958,N_12517);
nand U13285 (N_13285,N_12829,N_13003);
or U13286 (N_13286,N_12832,N_13040);
xor U13287 (N_13287,N_12703,N_12830);
or U13288 (N_13288,N_12567,N_12536);
and U13289 (N_13289,N_13047,N_12732);
nor U13290 (N_13290,N_13121,N_12858);
and U13291 (N_13291,N_12910,N_12587);
or U13292 (N_13292,N_12957,N_12537);
nor U13293 (N_13293,N_12949,N_12860);
nand U13294 (N_13294,N_12904,N_12914);
xnor U13295 (N_13295,N_13100,N_12598);
nand U13296 (N_13296,N_12884,N_12679);
nand U13297 (N_13297,N_12501,N_12892);
xor U13298 (N_13298,N_13112,N_12786);
xor U13299 (N_13299,N_12991,N_13036);
and U13300 (N_13300,N_12533,N_12771);
and U13301 (N_13301,N_12967,N_13111);
nand U13302 (N_13302,N_12661,N_12927);
xor U13303 (N_13303,N_12842,N_12746);
or U13304 (N_13304,N_12553,N_12912);
nand U13305 (N_13305,N_12733,N_12764);
or U13306 (N_13306,N_12612,N_12543);
or U13307 (N_13307,N_12976,N_12666);
nor U13308 (N_13308,N_12843,N_13086);
xor U13309 (N_13309,N_12563,N_13051);
or U13310 (N_13310,N_12604,N_13080);
nor U13311 (N_13311,N_12982,N_12981);
or U13312 (N_13312,N_12560,N_12940);
nand U13313 (N_13313,N_12712,N_12635);
and U13314 (N_13314,N_12925,N_12552);
and U13315 (N_13315,N_12709,N_12665);
xor U13316 (N_13316,N_12778,N_12864);
or U13317 (N_13317,N_12876,N_12586);
xnor U13318 (N_13318,N_12895,N_13083);
nor U13319 (N_13319,N_12659,N_12871);
nand U13320 (N_13320,N_12729,N_12780);
nand U13321 (N_13321,N_12845,N_12897);
xor U13322 (N_13322,N_12579,N_13043);
nand U13323 (N_13323,N_12593,N_12920);
xor U13324 (N_13324,N_13072,N_12796);
nand U13325 (N_13325,N_13017,N_12671);
nor U13326 (N_13326,N_13122,N_12886);
or U13327 (N_13327,N_12736,N_12556);
xor U13328 (N_13328,N_12792,N_12873);
and U13329 (N_13329,N_12752,N_12769);
xor U13330 (N_13330,N_12624,N_13041);
nand U13331 (N_13331,N_13071,N_12546);
xor U13332 (N_13332,N_12602,N_12570);
nor U13333 (N_13333,N_13115,N_13000);
nand U13334 (N_13334,N_13055,N_12972);
and U13335 (N_13335,N_12880,N_12505);
nand U13336 (N_13336,N_12607,N_12626);
xor U13337 (N_13337,N_12645,N_12603);
and U13338 (N_13338,N_12630,N_12812);
or U13339 (N_13339,N_12983,N_12695);
xor U13340 (N_13340,N_12558,N_12585);
and U13341 (N_13341,N_12526,N_12740);
nand U13342 (N_13342,N_12999,N_13030);
xnor U13343 (N_13343,N_12588,N_12719);
or U13344 (N_13344,N_12978,N_13098);
or U13345 (N_13345,N_13108,N_13001);
xor U13346 (N_13346,N_12854,N_12820);
xor U13347 (N_13347,N_13096,N_12672);
nor U13348 (N_13348,N_12975,N_13088);
nand U13349 (N_13349,N_13033,N_12879);
nor U13350 (N_13350,N_12828,N_12649);
nor U13351 (N_13351,N_13026,N_12522);
and U13352 (N_13352,N_12814,N_12664);
or U13353 (N_13353,N_12997,N_12900);
nor U13354 (N_13354,N_12966,N_12868);
nor U13355 (N_13355,N_12888,N_13007);
xnor U13356 (N_13356,N_12964,N_12718);
nand U13357 (N_13357,N_12962,N_12862);
xnor U13358 (N_13358,N_12692,N_12986);
nor U13359 (N_13359,N_12751,N_12704);
xor U13360 (N_13360,N_13006,N_12625);
nand U13361 (N_13361,N_12762,N_12800);
or U13362 (N_13362,N_12702,N_13116);
xor U13363 (N_13363,N_12785,N_12644);
xnor U13364 (N_13364,N_12849,N_13042);
nor U13365 (N_13365,N_13016,N_13079);
and U13366 (N_13366,N_13102,N_12689);
nand U13367 (N_13367,N_12684,N_12595);
xor U13368 (N_13368,N_12606,N_12669);
or U13369 (N_13369,N_13049,N_12959);
nor U13370 (N_13370,N_12848,N_12756);
nand U13371 (N_13371,N_13061,N_12584);
and U13372 (N_13372,N_12833,N_12651);
and U13373 (N_13373,N_12590,N_12643);
and U13374 (N_13374,N_12717,N_12634);
xnor U13375 (N_13375,N_12714,N_12855);
or U13376 (N_13376,N_12539,N_13123);
nand U13377 (N_13377,N_12853,N_12559);
or U13378 (N_13378,N_12866,N_12977);
nor U13379 (N_13379,N_13020,N_12928);
and U13380 (N_13380,N_12676,N_12708);
or U13381 (N_13381,N_12767,N_12794);
nor U13382 (N_13382,N_12615,N_12961);
or U13383 (N_13383,N_12954,N_12540);
and U13384 (N_13384,N_12915,N_13012);
nor U13385 (N_13385,N_12680,N_12852);
nand U13386 (N_13386,N_12592,N_12985);
xor U13387 (N_13387,N_12521,N_12942);
and U13388 (N_13388,N_12677,N_12527);
and U13389 (N_13389,N_12911,N_13067);
nand U13390 (N_13390,N_12948,N_13034);
nand U13391 (N_13391,N_12747,N_12768);
nand U13392 (N_13392,N_12623,N_12650);
and U13393 (N_13393,N_12947,N_12516);
and U13394 (N_13394,N_12728,N_12619);
nand U13395 (N_13395,N_12822,N_12662);
or U13396 (N_13396,N_12554,N_12565);
or U13397 (N_13397,N_12872,N_12550);
or U13398 (N_13398,N_13035,N_12755);
nor U13399 (N_13399,N_12514,N_12597);
xnor U13400 (N_13400,N_12816,N_12801);
nor U13401 (N_13401,N_12970,N_12823);
xor U13402 (N_13402,N_13114,N_12761);
or U13403 (N_13403,N_13015,N_13078);
xnor U13404 (N_13404,N_13024,N_12882);
or U13405 (N_13405,N_12799,N_12528);
and U13406 (N_13406,N_12773,N_12524);
or U13407 (N_13407,N_13060,N_12697);
or U13408 (N_13408,N_12555,N_12783);
or U13409 (N_13409,N_12807,N_12641);
nand U13410 (N_13410,N_12797,N_12696);
or U13411 (N_13411,N_12698,N_12994);
xnor U13412 (N_13412,N_13093,N_12810);
xor U13413 (N_13413,N_13056,N_12687);
nand U13414 (N_13414,N_13019,N_12512);
nand U13415 (N_13415,N_12541,N_12531);
nor U13416 (N_13416,N_12819,N_12818);
xor U13417 (N_13417,N_12885,N_12750);
xnor U13418 (N_13418,N_12793,N_12648);
and U13419 (N_13419,N_12919,N_12776);
and U13420 (N_13420,N_12811,N_12547);
nor U13421 (N_13421,N_12525,N_12707);
nor U13422 (N_13422,N_13117,N_12562);
nand U13423 (N_13423,N_12673,N_12939);
xnor U13424 (N_13424,N_12757,N_12835);
or U13425 (N_13425,N_12878,N_12930);
nor U13426 (N_13426,N_12998,N_12795);
and U13427 (N_13427,N_12700,N_12542);
and U13428 (N_13428,N_12657,N_12881);
and U13429 (N_13429,N_12622,N_12549);
and U13430 (N_13430,N_12726,N_12596);
nor U13431 (N_13431,N_12777,N_12571);
nand U13432 (N_13432,N_12953,N_13099);
xor U13433 (N_13433,N_12917,N_13031);
and U13434 (N_13434,N_12744,N_12808);
and U13435 (N_13435,N_13077,N_12655);
xnor U13436 (N_13436,N_13073,N_12629);
or U13437 (N_13437,N_12893,N_12674);
xnor U13438 (N_13438,N_12710,N_12542);
nand U13439 (N_13439,N_12671,N_12786);
nand U13440 (N_13440,N_12586,N_12577);
nand U13441 (N_13441,N_12896,N_13064);
nand U13442 (N_13442,N_12768,N_12732);
xor U13443 (N_13443,N_12698,N_12797);
xor U13444 (N_13444,N_12835,N_12662);
nor U13445 (N_13445,N_12717,N_12738);
nand U13446 (N_13446,N_12581,N_13103);
or U13447 (N_13447,N_13103,N_12863);
nand U13448 (N_13448,N_12931,N_12671);
xnor U13449 (N_13449,N_12927,N_12891);
nand U13450 (N_13450,N_12933,N_12902);
xor U13451 (N_13451,N_12672,N_12907);
nand U13452 (N_13452,N_13028,N_12646);
xor U13453 (N_13453,N_12723,N_12977);
or U13454 (N_13454,N_12529,N_12872);
and U13455 (N_13455,N_12902,N_12842);
and U13456 (N_13456,N_12787,N_12939);
nor U13457 (N_13457,N_12567,N_12657);
nor U13458 (N_13458,N_12795,N_12620);
xnor U13459 (N_13459,N_13080,N_13079);
nand U13460 (N_13460,N_12745,N_12662);
xor U13461 (N_13461,N_12502,N_12936);
nand U13462 (N_13462,N_12706,N_12685);
xor U13463 (N_13463,N_13036,N_12882);
xnor U13464 (N_13464,N_13004,N_12736);
xnor U13465 (N_13465,N_12668,N_12874);
and U13466 (N_13466,N_12579,N_12665);
or U13467 (N_13467,N_12633,N_12935);
nand U13468 (N_13468,N_12874,N_12590);
or U13469 (N_13469,N_13061,N_12979);
xor U13470 (N_13470,N_12691,N_12543);
or U13471 (N_13471,N_12884,N_12872);
nor U13472 (N_13472,N_13030,N_13066);
and U13473 (N_13473,N_12827,N_12613);
nor U13474 (N_13474,N_12945,N_12960);
nand U13475 (N_13475,N_13104,N_13011);
and U13476 (N_13476,N_12839,N_12670);
and U13477 (N_13477,N_12973,N_12803);
or U13478 (N_13478,N_12837,N_12727);
and U13479 (N_13479,N_12594,N_12639);
nand U13480 (N_13480,N_12685,N_12698);
and U13481 (N_13481,N_12820,N_12589);
or U13482 (N_13482,N_12799,N_13000);
and U13483 (N_13483,N_12763,N_13059);
or U13484 (N_13484,N_12687,N_12686);
nor U13485 (N_13485,N_12586,N_13053);
nand U13486 (N_13486,N_13013,N_12882);
and U13487 (N_13487,N_12507,N_12727);
xnor U13488 (N_13488,N_12608,N_12534);
nor U13489 (N_13489,N_12877,N_12839);
nand U13490 (N_13490,N_12825,N_13010);
nor U13491 (N_13491,N_13057,N_12976);
or U13492 (N_13492,N_12797,N_13086);
xnor U13493 (N_13493,N_12640,N_12655);
nor U13494 (N_13494,N_12972,N_13102);
and U13495 (N_13495,N_12872,N_12599);
or U13496 (N_13496,N_12737,N_12775);
and U13497 (N_13497,N_12798,N_12547);
nand U13498 (N_13498,N_12564,N_12508);
nor U13499 (N_13499,N_12542,N_12563);
xnor U13500 (N_13500,N_12720,N_12945);
or U13501 (N_13501,N_12619,N_12709);
nor U13502 (N_13502,N_13003,N_13031);
nor U13503 (N_13503,N_12932,N_12960);
nand U13504 (N_13504,N_12775,N_12789);
xor U13505 (N_13505,N_12932,N_13029);
nand U13506 (N_13506,N_12582,N_12727);
and U13507 (N_13507,N_12744,N_12738);
or U13508 (N_13508,N_12745,N_13103);
or U13509 (N_13509,N_12599,N_13075);
xor U13510 (N_13510,N_13028,N_12891);
and U13511 (N_13511,N_12837,N_12668);
xnor U13512 (N_13512,N_12826,N_12524);
and U13513 (N_13513,N_12554,N_12947);
xnor U13514 (N_13514,N_12888,N_13061);
nand U13515 (N_13515,N_13003,N_12884);
nor U13516 (N_13516,N_12817,N_12505);
or U13517 (N_13517,N_13046,N_13031);
nor U13518 (N_13518,N_12786,N_12543);
or U13519 (N_13519,N_12637,N_12562);
nor U13520 (N_13520,N_12786,N_12738);
nand U13521 (N_13521,N_12782,N_12680);
and U13522 (N_13522,N_12631,N_12560);
nand U13523 (N_13523,N_13037,N_12706);
and U13524 (N_13524,N_12580,N_12592);
xnor U13525 (N_13525,N_12556,N_12569);
nand U13526 (N_13526,N_12566,N_12781);
or U13527 (N_13527,N_12878,N_12796);
xor U13528 (N_13528,N_12922,N_13116);
and U13529 (N_13529,N_12873,N_12931);
or U13530 (N_13530,N_12754,N_12733);
nor U13531 (N_13531,N_12822,N_12767);
nand U13532 (N_13532,N_12943,N_13069);
or U13533 (N_13533,N_12878,N_12936);
xor U13534 (N_13534,N_12569,N_12912);
nand U13535 (N_13535,N_12597,N_12886);
or U13536 (N_13536,N_12889,N_13012);
nor U13537 (N_13537,N_12573,N_12952);
nand U13538 (N_13538,N_12810,N_12996);
and U13539 (N_13539,N_12895,N_12620);
nand U13540 (N_13540,N_12655,N_12990);
nor U13541 (N_13541,N_12785,N_13049);
nor U13542 (N_13542,N_12899,N_12557);
and U13543 (N_13543,N_12595,N_12682);
xor U13544 (N_13544,N_12951,N_12940);
nand U13545 (N_13545,N_12818,N_12731);
nand U13546 (N_13546,N_12836,N_12781);
or U13547 (N_13547,N_12997,N_13066);
and U13548 (N_13548,N_13123,N_12667);
nand U13549 (N_13549,N_13063,N_13103);
or U13550 (N_13550,N_12685,N_12502);
nand U13551 (N_13551,N_12582,N_12624);
nor U13552 (N_13552,N_13083,N_13040);
xor U13553 (N_13553,N_12725,N_12526);
nand U13554 (N_13554,N_12508,N_12742);
nand U13555 (N_13555,N_12595,N_12703);
nor U13556 (N_13556,N_12528,N_12806);
or U13557 (N_13557,N_12837,N_12953);
nor U13558 (N_13558,N_12779,N_12614);
nor U13559 (N_13559,N_12567,N_12609);
nand U13560 (N_13560,N_13112,N_12931);
nor U13561 (N_13561,N_12946,N_12574);
xnor U13562 (N_13562,N_13115,N_12516);
or U13563 (N_13563,N_12818,N_12694);
nand U13564 (N_13564,N_12577,N_12926);
and U13565 (N_13565,N_12777,N_13028);
or U13566 (N_13566,N_13114,N_12742);
nand U13567 (N_13567,N_12890,N_12801);
nand U13568 (N_13568,N_12517,N_13030);
and U13569 (N_13569,N_12517,N_12597);
nor U13570 (N_13570,N_12641,N_12586);
nor U13571 (N_13571,N_12988,N_13077);
nand U13572 (N_13572,N_12803,N_12501);
xnor U13573 (N_13573,N_12839,N_12857);
xor U13574 (N_13574,N_12704,N_12858);
or U13575 (N_13575,N_12663,N_12865);
nor U13576 (N_13576,N_12918,N_12920);
nand U13577 (N_13577,N_12652,N_13104);
and U13578 (N_13578,N_13069,N_12652);
nand U13579 (N_13579,N_13012,N_12746);
nand U13580 (N_13580,N_12861,N_12822);
and U13581 (N_13581,N_12530,N_12510);
nand U13582 (N_13582,N_12642,N_12857);
and U13583 (N_13583,N_12598,N_13022);
nand U13584 (N_13584,N_12858,N_12694);
nor U13585 (N_13585,N_13016,N_12506);
xnor U13586 (N_13586,N_13118,N_12583);
and U13587 (N_13587,N_12698,N_12523);
xor U13588 (N_13588,N_12623,N_12625);
xnor U13589 (N_13589,N_12542,N_13105);
nor U13590 (N_13590,N_12512,N_13114);
and U13591 (N_13591,N_12800,N_12823);
and U13592 (N_13592,N_12752,N_13036);
nor U13593 (N_13593,N_12589,N_12719);
and U13594 (N_13594,N_12762,N_13011);
xnor U13595 (N_13595,N_12746,N_12856);
nand U13596 (N_13596,N_13037,N_13102);
nand U13597 (N_13597,N_12615,N_12915);
nor U13598 (N_13598,N_12936,N_12813);
xnor U13599 (N_13599,N_12910,N_12744);
or U13600 (N_13600,N_12619,N_12571);
or U13601 (N_13601,N_12850,N_12595);
nor U13602 (N_13602,N_12838,N_12871);
and U13603 (N_13603,N_12621,N_12655);
nor U13604 (N_13604,N_12627,N_12850);
nor U13605 (N_13605,N_12676,N_12576);
and U13606 (N_13606,N_12505,N_12588);
and U13607 (N_13607,N_12780,N_12820);
and U13608 (N_13608,N_12705,N_12955);
or U13609 (N_13609,N_13040,N_13068);
and U13610 (N_13610,N_12966,N_12677);
and U13611 (N_13611,N_12516,N_12861);
nand U13612 (N_13612,N_12776,N_13102);
and U13613 (N_13613,N_12873,N_12963);
xnor U13614 (N_13614,N_12561,N_13006);
or U13615 (N_13615,N_12680,N_12781);
xor U13616 (N_13616,N_12716,N_12978);
nor U13617 (N_13617,N_12563,N_12600);
xnor U13618 (N_13618,N_12994,N_12533);
nor U13619 (N_13619,N_12829,N_13050);
nand U13620 (N_13620,N_12677,N_12921);
or U13621 (N_13621,N_12821,N_12734);
nand U13622 (N_13622,N_12549,N_12941);
nand U13623 (N_13623,N_12705,N_12768);
xor U13624 (N_13624,N_12735,N_12507);
xor U13625 (N_13625,N_12827,N_12728);
nand U13626 (N_13626,N_13006,N_12606);
xnor U13627 (N_13627,N_12809,N_12611);
and U13628 (N_13628,N_13009,N_13044);
nor U13629 (N_13629,N_12682,N_13026);
and U13630 (N_13630,N_12808,N_12511);
and U13631 (N_13631,N_13115,N_12889);
or U13632 (N_13632,N_12607,N_12701);
and U13633 (N_13633,N_13012,N_12767);
xnor U13634 (N_13634,N_13025,N_12921);
nor U13635 (N_13635,N_12518,N_12787);
nand U13636 (N_13636,N_12759,N_12695);
xnor U13637 (N_13637,N_13024,N_13108);
nand U13638 (N_13638,N_13095,N_13120);
nor U13639 (N_13639,N_12910,N_12651);
nand U13640 (N_13640,N_12717,N_12917);
and U13641 (N_13641,N_12968,N_12938);
nand U13642 (N_13642,N_12637,N_12822);
or U13643 (N_13643,N_12937,N_12850);
xor U13644 (N_13644,N_12612,N_12675);
nor U13645 (N_13645,N_12571,N_12915);
nor U13646 (N_13646,N_12624,N_13081);
nand U13647 (N_13647,N_12973,N_12914);
nand U13648 (N_13648,N_12812,N_12667);
xor U13649 (N_13649,N_12786,N_12828);
xnor U13650 (N_13650,N_12908,N_13084);
or U13651 (N_13651,N_12767,N_12743);
and U13652 (N_13652,N_12969,N_12527);
or U13653 (N_13653,N_13079,N_12987);
or U13654 (N_13654,N_12665,N_12983);
or U13655 (N_13655,N_12706,N_12629);
or U13656 (N_13656,N_12750,N_12573);
nor U13657 (N_13657,N_12904,N_13077);
nand U13658 (N_13658,N_13116,N_12764);
or U13659 (N_13659,N_13051,N_12774);
xnor U13660 (N_13660,N_12732,N_13067);
or U13661 (N_13661,N_12796,N_12715);
nor U13662 (N_13662,N_12717,N_12706);
and U13663 (N_13663,N_12616,N_12770);
nand U13664 (N_13664,N_12632,N_12659);
and U13665 (N_13665,N_12736,N_12913);
nor U13666 (N_13666,N_12650,N_12529);
xor U13667 (N_13667,N_12892,N_12778);
nor U13668 (N_13668,N_12508,N_13072);
xnor U13669 (N_13669,N_12750,N_12592);
xor U13670 (N_13670,N_12828,N_12500);
nor U13671 (N_13671,N_12897,N_12825);
and U13672 (N_13672,N_12527,N_12512);
nor U13673 (N_13673,N_12758,N_12790);
nor U13674 (N_13674,N_12777,N_12845);
or U13675 (N_13675,N_12534,N_12748);
xnor U13676 (N_13676,N_12630,N_12793);
xor U13677 (N_13677,N_12855,N_12619);
nor U13678 (N_13678,N_12894,N_12957);
and U13679 (N_13679,N_12968,N_12889);
and U13680 (N_13680,N_12721,N_12964);
xnor U13681 (N_13681,N_13027,N_12846);
nand U13682 (N_13682,N_12969,N_13097);
and U13683 (N_13683,N_12707,N_12976);
and U13684 (N_13684,N_12939,N_13016);
xor U13685 (N_13685,N_13053,N_13006);
xor U13686 (N_13686,N_12712,N_12529);
nor U13687 (N_13687,N_12943,N_12587);
xor U13688 (N_13688,N_12905,N_12789);
and U13689 (N_13689,N_12999,N_12548);
and U13690 (N_13690,N_12655,N_12718);
nand U13691 (N_13691,N_12915,N_12871);
or U13692 (N_13692,N_12988,N_12747);
xor U13693 (N_13693,N_12547,N_12723);
nor U13694 (N_13694,N_12598,N_12789);
nand U13695 (N_13695,N_12571,N_12780);
and U13696 (N_13696,N_12935,N_12601);
xor U13697 (N_13697,N_12749,N_12787);
xnor U13698 (N_13698,N_12918,N_13082);
or U13699 (N_13699,N_12583,N_12867);
xor U13700 (N_13700,N_12670,N_12700);
nand U13701 (N_13701,N_12697,N_12528);
and U13702 (N_13702,N_12613,N_12505);
and U13703 (N_13703,N_12932,N_12836);
nand U13704 (N_13704,N_12576,N_12921);
nor U13705 (N_13705,N_12894,N_12728);
and U13706 (N_13706,N_12883,N_13002);
and U13707 (N_13707,N_13064,N_12768);
or U13708 (N_13708,N_13113,N_12693);
nor U13709 (N_13709,N_13077,N_13074);
nor U13710 (N_13710,N_13104,N_12780);
nor U13711 (N_13711,N_12692,N_13080);
nand U13712 (N_13712,N_12841,N_13108);
and U13713 (N_13713,N_12677,N_13028);
nand U13714 (N_13714,N_12902,N_12995);
nor U13715 (N_13715,N_12775,N_13054);
nor U13716 (N_13716,N_12547,N_12970);
xnor U13717 (N_13717,N_13032,N_12736);
nand U13718 (N_13718,N_12660,N_12579);
xnor U13719 (N_13719,N_13052,N_13038);
nor U13720 (N_13720,N_12872,N_12677);
and U13721 (N_13721,N_12958,N_12713);
xor U13722 (N_13722,N_13026,N_12568);
xor U13723 (N_13723,N_12511,N_12523);
xor U13724 (N_13724,N_12987,N_13102);
or U13725 (N_13725,N_12825,N_12999);
or U13726 (N_13726,N_12646,N_12881);
nor U13727 (N_13727,N_12621,N_12531);
nor U13728 (N_13728,N_12697,N_12848);
nor U13729 (N_13729,N_12555,N_12678);
and U13730 (N_13730,N_12651,N_13044);
or U13731 (N_13731,N_12601,N_13073);
nor U13732 (N_13732,N_12979,N_12650);
and U13733 (N_13733,N_12980,N_12985);
xor U13734 (N_13734,N_12989,N_13040);
and U13735 (N_13735,N_12605,N_13076);
and U13736 (N_13736,N_12587,N_13063);
nor U13737 (N_13737,N_12558,N_12508);
and U13738 (N_13738,N_12668,N_13083);
nand U13739 (N_13739,N_13027,N_12806);
and U13740 (N_13740,N_12531,N_12950);
nor U13741 (N_13741,N_12996,N_13035);
xor U13742 (N_13742,N_13064,N_12951);
or U13743 (N_13743,N_12540,N_12934);
nor U13744 (N_13744,N_12854,N_12920);
nand U13745 (N_13745,N_12547,N_12603);
nor U13746 (N_13746,N_12979,N_12869);
nand U13747 (N_13747,N_12770,N_13107);
nor U13748 (N_13748,N_12808,N_13009);
and U13749 (N_13749,N_12780,N_12939);
nand U13750 (N_13750,N_13415,N_13376);
or U13751 (N_13751,N_13486,N_13592);
nand U13752 (N_13752,N_13741,N_13568);
and U13753 (N_13753,N_13687,N_13314);
xor U13754 (N_13754,N_13626,N_13146);
and U13755 (N_13755,N_13522,N_13342);
or U13756 (N_13756,N_13419,N_13391);
nor U13757 (N_13757,N_13564,N_13251);
nand U13758 (N_13758,N_13427,N_13305);
nand U13759 (N_13759,N_13671,N_13240);
xor U13760 (N_13760,N_13683,N_13519);
or U13761 (N_13761,N_13622,N_13721);
xor U13762 (N_13762,N_13509,N_13563);
and U13763 (N_13763,N_13142,N_13295);
nor U13764 (N_13764,N_13565,N_13575);
nand U13765 (N_13765,N_13266,N_13432);
nand U13766 (N_13766,N_13647,N_13732);
and U13767 (N_13767,N_13663,N_13204);
nor U13768 (N_13768,N_13658,N_13170);
or U13769 (N_13769,N_13422,N_13218);
nand U13770 (N_13770,N_13746,N_13514);
nor U13771 (N_13771,N_13617,N_13479);
and U13772 (N_13772,N_13148,N_13413);
or U13773 (N_13773,N_13310,N_13225);
nand U13774 (N_13774,N_13337,N_13631);
nor U13775 (N_13775,N_13356,N_13395);
nand U13776 (N_13776,N_13580,N_13516);
nand U13777 (N_13777,N_13676,N_13633);
xor U13778 (N_13778,N_13484,N_13720);
nand U13779 (N_13779,N_13134,N_13618);
and U13780 (N_13780,N_13210,N_13181);
nand U13781 (N_13781,N_13616,N_13371);
xnor U13782 (N_13782,N_13169,N_13462);
nor U13783 (N_13783,N_13268,N_13137);
xor U13784 (N_13784,N_13284,N_13678);
nor U13785 (N_13785,N_13742,N_13696);
and U13786 (N_13786,N_13476,N_13151);
nand U13787 (N_13787,N_13641,N_13458);
xnor U13788 (N_13788,N_13452,N_13465);
nor U13789 (N_13789,N_13749,N_13457);
nand U13790 (N_13790,N_13220,N_13190);
nand U13791 (N_13791,N_13171,N_13283);
nor U13792 (N_13792,N_13144,N_13304);
nor U13793 (N_13793,N_13736,N_13277);
or U13794 (N_13794,N_13667,N_13232);
or U13795 (N_13795,N_13513,N_13420);
and U13796 (N_13796,N_13530,N_13377);
nor U13797 (N_13797,N_13497,N_13512);
and U13798 (N_13798,N_13672,N_13227);
nand U13799 (N_13799,N_13233,N_13609);
and U13800 (N_13800,N_13552,N_13161);
xor U13801 (N_13801,N_13689,N_13493);
and U13802 (N_13802,N_13318,N_13459);
nor U13803 (N_13803,N_13162,N_13650);
nand U13804 (N_13804,N_13273,N_13440);
and U13805 (N_13805,N_13136,N_13418);
or U13806 (N_13806,N_13322,N_13521);
nor U13807 (N_13807,N_13597,N_13475);
nand U13808 (N_13808,N_13333,N_13699);
or U13809 (N_13809,N_13383,N_13308);
nand U13810 (N_13810,N_13399,N_13525);
and U13811 (N_13811,N_13585,N_13397);
and U13812 (N_13812,N_13135,N_13620);
nand U13813 (N_13813,N_13213,N_13339);
or U13814 (N_13814,N_13272,N_13400);
nor U13815 (N_13815,N_13651,N_13348);
or U13816 (N_13816,N_13586,N_13589);
or U13817 (N_13817,N_13195,N_13186);
xnor U13818 (N_13818,N_13713,N_13487);
or U13819 (N_13819,N_13293,N_13401);
nand U13820 (N_13820,N_13707,N_13287);
and U13821 (N_13821,N_13133,N_13191);
xor U13822 (N_13822,N_13228,N_13574);
nand U13823 (N_13823,N_13543,N_13201);
or U13824 (N_13824,N_13526,N_13389);
or U13825 (N_13825,N_13163,N_13288);
nor U13826 (N_13826,N_13402,N_13498);
and U13827 (N_13827,N_13177,N_13692);
and U13828 (N_13828,N_13634,N_13435);
nand U13829 (N_13829,N_13143,N_13385);
and U13830 (N_13830,N_13159,N_13321);
and U13831 (N_13831,N_13700,N_13128);
and U13832 (N_13832,N_13278,N_13725);
nor U13833 (N_13833,N_13340,N_13551);
nand U13834 (N_13834,N_13320,N_13330);
nor U13835 (N_13835,N_13546,N_13361);
nor U13836 (N_13836,N_13200,N_13262);
or U13837 (N_13837,N_13734,N_13409);
and U13838 (N_13838,N_13194,N_13405);
xor U13839 (N_13839,N_13317,N_13613);
or U13840 (N_13840,N_13360,N_13203);
and U13841 (N_13841,N_13670,N_13160);
or U13842 (N_13842,N_13542,N_13224);
nand U13843 (N_13843,N_13545,N_13728);
or U13844 (N_13844,N_13346,N_13504);
nor U13845 (N_13845,N_13619,N_13444);
or U13846 (N_13846,N_13127,N_13534);
xor U13847 (N_13847,N_13433,N_13297);
and U13848 (N_13848,N_13198,N_13470);
and U13849 (N_13849,N_13209,N_13478);
and U13850 (N_13850,N_13403,N_13298);
nand U13851 (N_13851,N_13363,N_13247);
or U13852 (N_13852,N_13174,N_13446);
or U13853 (N_13853,N_13614,N_13294);
nand U13854 (N_13854,N_13531,N_13518);
nor U13855 (N_13855,N_13153,N_13680);
and U13856 (N_13856,N_13366,N_13515);
and U13857 (N_13857,N_13483,N_13147);
and U13858 (N_13858,N_13207,N_13248);
nor U13859 (N_13859,N_13410,N_13537);
nand U13860 (N_13860,N_13168,N_13390);
or U13861 (N_13861,N_13197,N_13566);
xnor U13862 (N_13862,N_13416,N_13276);
nand U13863 (N_13863,N_13445,N_13607);
nand U13864 (N_13864,N_13260,N_13747);
and U13865 (N_13865,N_13185,N_13659);
and U13866 (N_13866,N_13417,N_13702);
nand U13867 (N_13867,N_13471,N_13523);
and U13868 (N_13868,N_13508,N_13704);
or U13869 (N_13869,N_13660,N_13517);
nand U13870 (N_13870,N_13600,N_13398);
nor U13871 (N_13871,N_13381,N_13193);
and U13872 (N_13872,N_13735,N_13208);
nor U13873 (N_13873,N_13187,N_13296);
nor U13874 (N_13874,N_13219,N_13341);
nor U13875 (N_13875,N_13463,N_13610);
xnor U13876 (N_13876,N_13450,N_13679);
xnor U13877 (N_13877,N_13624,N_13500);
nand U13878 (N_13878,N_13349,N_13315);
and U13879 (N_13879,N_13718,N_13152);
nand U13880 (N_13880,N_13249,N_13584);
xnor U13881 (N_13881,N_13644,N_13733);
or U13882 (N_13882,N_13596,N_13234);
nand U13883 (N_13883,N_13214,N_13665);
nand U13884 (N_13884,N_13384,N_13673);
and U13885 (N_13885,N_13351,N_13290);
xor U13886 (N_13886,N_13691,N_13643);
nor U13887 (N_13887,N_13571,N_13374);
and U13888 (N_13888,N_13343,N_13263);
and U13889 (N_13889,N_13682,N_13538);
or U13890 (N_13890,N_13464,N_13173);
and U13891 (N_13891,N_13726,N_13695);
nor U13892 (N_13892,N_13140,N_13338);
nand U13893 (N_13893,N_13601,N_13473);
xor U13894 (N_13894,N_13434,N_13345);
or U13895 (N_13895,N_13453,N_13505);
or U13896 (N_13896,N_13697,N_13535);
nand U13897 (N_13897,N_13598,N_13307);
xnor U13898 (N_13898,N_13387,N_13611);
nand U13899 (N_13899,N_13274,N_13291);
and U13900 (N_13900,N_13594,N_13540);
and U13901 (N_13901,N_13369,N_13164);
or U13902 (N_13902,N_13235,N_13477);
nor U13903 (N_13903,N_13502,N_13547);
or U13904 (N_13904,N_13456,N_13533);
nand U13905 (N_13905,N_13559,N_13587);
and U13906 (N_13906,N_13335,N_13623);
xnor U13907 (N_13907,N_13602,N_13327);
nor U13908 (N_13908,N_13536,N_13373);
and U13909 (N_13909,N_13367,N_13629);
or U13910 (N_13910,N_13158,N_13271);
xor U13911 (N_13911,N_13724,N_13269);
and U13912 (N_13912,N_13183,N_13352);
and U13913 (N_13913,N_13549,N_13638);
xor U13914 (N_13914,N_13694,N_13380);
and U13915 (N_13915,N_13309,N_13489);
or U13916 (N_13916,N_13443,N_13496);
xor U13917 (N_13917,N_13583,N_13392);
xor U13918 (N_13918,N_13156,N_13336);
xnor U13919 (N_13919,N_13709,N_13328);
nand U13920 (N_13920,N_13529,N_13157);
xnor U13921 (N_13921,N_13421,N_13578);
or U13922 (N_13922,N_13241,N_13238);
xor U13923 (N_13923,N_13404,N_13179);
or U13924 (N_13924,N_13506,N_13226);
and U13925 (N_13925,N_13264,N_13582);
or U13926 (N_13926,N_13354,N_13690);
nor U13927 (N_13927,N_13524,N_13379);
nor U13928 (N_13928,N_13605,N_13180);
nand U13929 (N_13929,N_13576,N_13528);
nand U13930 (N_13930,N_13488,N_13606);
nor U13931 (N_13931,N_13729,N_13739);
nor U13932 (N_13932,N_13125,N_13581);
nor U13933 (N_13933,N_13579,N_13637);
nor U13934 (N_13934,N_13256,N_13282);
xor U13935 (N_13935,N_13635,N_13316);
xnor U13936 (N_13936,N_13603,N_13645);
or U13937 (N_13937,N_13299,N_13599);
and U13938 (N_13938,N_13743,N_13655);
nand U13939 (N_13939,N_13646,N_13737);
nor U13940 (N_13940,N_13292,N_13698);
and U13941 (N_13941,N_13710,N_13258);
and U13942 (N_13942,N_13372,N_13206);
and U13943 (N_13943,N_13431,N_13350);
and U13944 (N_13944,N_13550,N_13411);
or U13945 (N_13945,N_13244,N_13167);
nor U13946 (N_13946,N_13491,N_13306);
and U13947 (N_13947,N_13396,N_13166);
xor U13948 (N_13948,N_13362,N_13460);
xnor U13949 (N_13949,N_13242,N_13730);
xor U13950 (N_13950,N_13239,N_13378);
nand U13951 (N_13951,N_13357,N_13323);
and U13952 (N_13952,N_13731,N_13561);
nor U13953 (N_13953,N_13553,N_13359);
nand U13954 (N_13954,N_13253,N_13740);
or U13955 (N_13955,N_13325,N_13511);
xor U13956 (N_13956,N_13712,N_13236);
or U13957 (N_13957,N_13130,N_13237);
or U13958 (N_13958,N_13480,N_13567);
nor U13959 (N_13959,N_13532,N_13652);
and U13960 (N_13960,N_13714,N_13748);
xor U13961 (N_13961,N_13261,N_13715);
nand U13962 (N_13962,N_13243,N_13711);
and U13963 (N_13963,N_13628,N_13573);
nand U13964 (N_13964,N_13406,N_13621);
and U13965 (N_13965,N_13438,N_13331);
or U13966 (N_13966,N_13627,N_13324);
nand U13967 (N_13967,N_13745,N_13178);
nor U13968 (N_13968,N_13556,N_13329);
nor U13969 (N_13969,N_13469,N_13202);
nand U13970 (N_13970,N_13189,N_13615);
xor U13971 (N_13971,N_13590,N_13688);
and U13972 (N_13972,N_13286,N_13548);
nor U13973 (N_13973,N_13703,N_13426);
nand U13974 (N_13974,N_13192,N_13451);
xor U13975 (N_13975,N_13560,N_13216);
nand U13976 (N_13976,N_13708,N_13139);
xnor U13977 (N_13977,N_13557,N_13408);
and U13978 (N_13978,N_13149,N_13577);
nand U13979 (N_13979,N_13481,N_13722);
nand U13980 (N_13980,N_13215,N_13701);
nor U13981 (N_13981,N_13461,N_13686);
xnor U13982 (N_13982,N_13407,N_13437);
nor U13983 (N_13983,N_13544,N_13539);
nor U13984 (N_13984,N_13454,N_13270);
or U13985 (N_13985,N_13138,N_13661);
xnor U13986 (N_13986,N_13172,N_13222);
nand U13987 (N_13987,N_13555,N_13267);
nand U13988 (N_13988,N_13717,N_13259);
and U13989 (N_13989,N_13719,N_13612);
nand U13990 (N_13990,N_13448,N_13145);
xnor U13991 (N_13991,N_13668,N_13706);
nand U13992 (N_13992,N_13428,N_13669);
nor U13993 (N_13993,N_13693,N_13176);
nand U13994 (N_13994,N_13472,N_13591);
or U13995 (N_13995,N_13442,N_13312);
and U13996 (N_13996,N_13326,N_13265);
and U13997 (N_13997,N_13744,N_13188);
or U13998 (N_13998,N_13636,N_13510);
and U13999 (N_13999,N_13467,N_13595);
nor U14000 (N_14000,N_13570,N_13394);
or U14001 (N_14001,N_13449,N_13677);
xnor U14002 (N_14002,N_13370,N_13499);
and U14003 (N_14003,N_13501,N_13640);
or U14004 (N_14004,N_13572,N_13129);
or U14005 (N_14005,N_13664,N_13723);
nor U14006 (N_14006,N_13474,N_13141);
and U14007 (N_14007,N_13230,N_13250);
or U14008 (N_14008,N_13301,N_13334);
and U14009 (N_14009,N_13527,N_13344);
nand U14010 (N_14010,N_13439,N_13364);
nand U14011 (N_14011,N_13246,N_13554);
xnor U14012 (N_14012,N_13414,N_13468);
and U14013 (N_14013,N_13155,N_13593);
nand U14014 (N_14014,N_13727,N_13275);
xnor U14015 (N_14015,N_13495,N_13642);
xor U14016 (N_14016,N_13503,N_13441);
and U14017 (N_14017,N_13632,N_13520);
or U14018 (N_14018,N_13223,N_13199);
nand U14019 (N_14019,N_13436,N_13429);
nor U14020 (N_14020,N_13165,N_13205);
nor U14021 (N_14021,N_13355,N_13126);
nor U14022 (N_14022,N_13196,N_13393);
or U14023 (N_14023,N_13182,N_13684);
or U14024 (N_14024,N_13455,N_13666);
or U14025 (N_14025,N_13653,N_13662);
xor U14026 (N_14026,N_13388,N_13485);
nor U14027 (N_14027,N_13252,N_13657);
xor U14028 (N_14028,N_13300,N_13604);
nor U14029 (N_14029,N_13490,N_13211);
or U14030 (N_14030,N_13254,N_13302);
xor U14031 (N_14031,N_13630,N_13353);
nor U14032 (N_14032,N_13716,N_13303);
and U14033 (N_14033,N_13639,N_13150);
xor U14034 (N_14034,N_13358,N_13257);
and U14035 (N_14035,N_13131,N_13558);
nor U14036 (N_14036,N_13466,N_13507);
nand U14037 (N_14037,N_13705,N_13562);
or U14038 (N_14038,N_13674,N_13319);
or U14039 (N_14039,N_13386,N_13365);
nand U14040 (N_14040,N_13221,N_13347);
xnor U14041 (N_14041,N_13313,N_13281);
nor U14042 (N_14042,N_13482,N_13212);
xnor U14043 (N_14043,N_13625,N_13184);
and U14044 (N_14044,N_13425,N_13231);
or U14045 (N_14045,N_13649,N_13423);
xnor U14046 (N_14046,N_13382,N_13424);
nand U14047 (N_14047,N_13154,N_13245);
nor U14048 (N_14048,N_13311,N_13569);
nor U14049 (N_14049,N_13648,N_13656);
and U14050 (N_14050,N_13685,N_13412);
or U14051 (N_14051,N_13279,N_13255);
nand U14052 (N_14052,N_13229,N_13492);
or U14053 (N_14053,N_13175,N_13675);
nand U14054 (N_14054,N_13430,N_13368);
xor U14055 (N_14055,N_13289,N_13738);
nand U14056 (N_14056,N_13375,N_13588);
or U14057 (N_14057,N_13132,N_13681);
xor U14058 (N_14058,N_13217,N_13608);
nand U14059 (N_14059,N_13285,N_13280);
nor U14060 (N_14060,N_13494,N_13654);
nor U14061 (N_14061,N_13541,N_13447);
nor U14062 (N_14062,N_13332,N_13715);
or U14063 (N_14063,N_13179,N_13575);
and U14064 (N_14064,N_13700,N_13703);
or U14065 (N_14065,N_13595,N_13322);
nor U14066 (N_14066,N_13669,N_13398);
or U14067 (N_14067,N_13747,N_13635);
xnor U14068 (N_14068,N_13651,N_13576);
nor U14069 (N_14069,N_13167,N_13612);
nand U14070 (N_14070,N_13579,N_13589);
or U14071 (N_14071,N_13556,N_13171);
nor U14072 (N_14072,N_13615,N_13494);
or U14073 (N_14073,N_13699,N_13693);
or U14074 (N_14074,N_13161,N_13446);
nor U14075 (N_14075,N_13535,N_13366);
nand U14076 (N_14076,N_13456,N_13219);
and U14077 (N_14077,N_13574,N_13656);
or U14078 (N_14078,N_13538,N_13394);
or U14079 (N_14079,N_13658,N_13440);
nand U14080 (N_14080,N_13473,N_13650);
nor U14081 (N_14081,N_13536,N_13213);
nor U14082 (N_14082,N_13363,N_13678);
xnor U14083 (N_14083,N_13229,N_13362);
and U14084 (N_14084,N_13702,N_13378);
or U14085 (N_14085,N_13526,N_13547);
nand U14086 (N_14086,N_13600,N_13708);
or U14087 (N_14087,N_13548,N_13587);
or U14088 (N_14088,N_13339,N_13424);
xnor U14089 (N_14089,N_13183,N_13389);
nor U14090 (N_14090,N_13270,N_13645);
and U14091 (N_14091,N_13331,N_13478);
and U14092 (N_14092,N_13656,N_13542);
nor U14093 (N_14093,N_13274,N_13142);
xnor U14094 (N_14094,N_13409,N_13550);
or U14095 (N_14095,N_13462,N_13502);
nor U14096 (N_14096,N_13571,N_13378);
xnor U14097 (N_14097,N_13300,N_13192);
nor U14098 (N_14098,N_13533,N_13368);
and U14099 (N_14099,N_13188,N_13563);
xor U14100 (N_14100,N_13662,N_13563);
xor U14101 (N_14101,N_13668,N_13647);
nand U14102 (N_14102,N_13548,N_13139);
nand U14103 (N_14103,N_13205,N_13676);
and U14104 (N_14104,N_13277,N_13420);
or U14105 (N_14105,N_13363,N_13706);
and U14106 (N_14106,N_13582,N_13193);
and U14107 (N_14107,N_13151,N_13380);
or U14108 (N_14108,N_13493,N_13420);
or U14109 (N_14109,N_13429,N_13162);
xor U14110 (N_14110,N_13443,N_13403);
nand U14111 (N_14111,N_13500,N_13682);
nor U14112 (N_14112,N_13250,N_13419);
nor U14113 (N_14113,N_13452,N_13496);
nor U14114 (N_14114,N_13539,N_13678);
xor U14115 (N_14115,N_13293,N_13532);
or U14116 (N_14116,N_13434,N_13259);
nor U14117 (N_14117,N_13142,N_13263);
or U14118 (N_14118,N_13232,N_13278);
xnor U14119 (N_14119,N_13456,N_13717);
nand U14120 (N_14120,N_13406,N_13462);
or U14121 (N_14121,N_13205,N_13280);
nor U14122 (N_14122,N_13142,N_13680);
nand U14123 (N_14123,N_13289,N_13723);
or U14124 (N_14124,N_13700,N_13732);
nor U14125 (N_14125,N_13242,N_13744);
nor U14126 (N_14126,N_13392,N_13347);
xor U14127 (N_14127,N_13576,N_13331);
nand U14128 (N_14128,N_13684,N_13739);
and U14129 (N_14129,N_13344,N_13269);
nand U14130 (N_14130,N_13471,N_13153);
nand U14131 (N_14131,N_13705,N_13613);
xor U14132 (N_14132,N_13288,N_13521);
nor U14133 (N_14133,N_13402,N_13490);
or U14134 (N_14134,N_13533,N_13361);
nor U14135 (N_14135,N_13154,N_13671);
xor U14136 (N_14136,N_13450,N_13566);
nor U14137 (N_14137,N_13723,N_13673);
nand U14138 (N_14138,N_13318,N_13681);
and U14139 (N_14139,N_13485,N_13191);
or U14140 (N_14140,N_13489,N_13602);
nor U14141 (N_14141,N_13547,N_13305);
nor U14142 (N_14142,N_13350,N_13591);
nor U14143 (N_14143,N_13273,N_13731);
and U14144 (N_14144,N_13624,N_13549);
nand U14145 (N_14145,N_13407,N_13493);
nand U14146 (N_14146,N_13426,N_13566);
and U14147 (N_14147,N_13172,N_13506);
or U14148 (N_14148,N_13222,N_13151);
nand U14149 (N_14149,N_13175,N_13729);
or U14150 (N_14150,N_13332,N_13275);
or U14151 (N_14151,N_13703,N_13175);
and U14152 (N_14152,N_13581,N_13141);
or U14153 (N_14153,N_13693,N_13154);
or U14154 (N_14154,N_13394,N_13728);
xnor U14155 (N_14155,N_13476,N_13175);
or U14156 (N_14156,N_13412,N_13414);
xnor U14157 (N_14157,N_13685,N_13167);
or U14158 (N_14158,N_13603,N_13342);
and U14159 (N_14159,N_13692,N_13255);
nor U14160 (N_14160,N_13476,N_13254);
nand U14161 (N_14161,N_13401,N_13371);
nor U14162 (N_14162,N_13550,N_13281);
xnor U14163 (N_14163,N_13417,N_13324);
nor U14164 (N_14164,N_13303,N_13216);
xnor U14165 (N_14165,N_13144,N_13722);
or U14166 (N_14166,N_13749,N_13471);
xor U14167 (N_14167,N_13634,N_13588);
nand U14168 (N_14168,N_13159,N_13187);
xnor U14169 (N_14169,N_13216,N_13415);
or U14170 (N_14170,N_13589,N_13316);
and U14171 (N_14171,N_13689,N_13138);
or U14172 (N_14172,N_13374,N_13515);
xor U14173 (N_14173,N_13505,N_13708);
and U14174 (N_14174,N_13329,N_13194);
nand U14175 (N_14175,N_13552,N_13524);
and U14176 (N_14176,N_13611,N_13214);
nor U14177 (N_14177,N_13135,N_13125);
or U14178 (N_14178,N_13704,N_13562);
xor U14179 (N_14179,N_13487,N_13234);
nand U14180 (N_14180,N_13288,N_13353);
nor U14181 (N_14181,N_13595,N_13632);
nand U14182 (N_14182,N_13627,N_13657);
or U14183 (N_14183,N_13175,N_13601);
nor U14184 (N_14184,N_13281,N_13659);
or U14185 (N_14185,N_13239,N_13159);
nand U14186 (N_14186,N_13194,N_13513);
nor U14187 (N_14187,N_13210,N_13325);
nand U14188 (N_14188,N_13459,N_13533);
or U14189 (N_14189,N_13284,N_13677);
xor U14190 (N_14190,N_13495,N_13611);
nand U14191 (N_14191,N_13195,N_13668);
nor U14192 (N_14192,N_13325,N_13619);
xnor U14193 (N_14193,N_13517,N_13326);
xnor U14194 (N_14194,N_13372,N_13276);
and U14195 (N_14195,N_13714,N_13742);
nor U14196 (N_14196,N_13507,N_13459);
nand U14197 (N_14197,N_13142,N_13533);
and U14198 (N_14198,N_13592,N_13511);
nor U14199 (N_14199,N_13268,N_13590);
xnor U14200 (N_14200,N_13698,N_13241);
or U14201 (N_14201,N_13452,N_13371);
nor U14202 (N_14202,N_13656,N_13719);
or U14203 (N_14203,N_13663,N_13528);
and U14204 (N_14204,N_13417,N_13198);
or U14205 (N_14205,N_13279,N_13470);
nor U14206 (N_14206,N_13302,N_13409);
nor U14207 (N_14207,N_13679,N_13387);
xor U14208 (N_14208,N_13521,N_13158);
and U14209 (N_14209,N_13165,N_13336);
or U14210 (N_14210,N_13370,N_13333);
nand U14211 (N_14211,N_13615,N_13146);
and U14212 (N_14212,N_13494,N_13171);
and U14213 (N_14213,N_13182,N_13409);
nand U14214 (N_14214,N_13656,N_13626);
xnor U14215 (N_14215,N_13435,N_13474);
nor U14216 (N_14216,N_13272,N_13729);
nor U14217 (N_14217,N_13424,N_13607);
nand U14218 (N_14218,N_13315,N_13233);
and U14219 (N_14219,N_13616,N_13662);
xnor U14220 (N_14220,N_13444,N_13577);
nand U14221 (N_14221,N_13692,N_13325);
or U14222 (N_14222,N_13200,N_13246);
nand U14223 (N_14223,N_13713,N_13192);
xor U14224 (N_14224,N_13403,N_13460);
nor U14225 (N_14225,N_13552,N_13176);
nor U14226 (N_14226,N_13331,N_13268);
nor U14227 (N_14227,N_13412,N_13668);
xor U14228 (N_14228,N_13644,N_13410);
or U14229 (N_14229,N_13463,N_13674);
nor U14230 (N_14230,N_13293,N_13158);
xnor U14231 (N_14231,N_13128,N_13376);
and U14232 (N_14232,N_13420,N_13414);
nor U14233 (N_14233,N_13407,N_13512);
xor U14234 (N_14234,N_13288,N_13641);
nor U14235 (N_14235,N_13216,N_13344);
or U14236 (N_14236,N_13163,N_13509);
or U14237 (N_14237,N_13388,N_13328);
xnor U14238 (N_14238,N_13302,N_13280);
nor U14239 (N_14239,N_13344,N_13696);
nand U14240 (N_14240,N_13598,N_13377);
nor U14241 (N_14241,N_13138,N_13545);
and U14242 (N_14242,N_13552,N_13174);
or U14243 (N_14243,N_13532,N_13733);
or U14244 (N_14244,N_13521,N_13600);
nand U14245 (N_14245,N_13389,N_13699);
or U14246 (N_14246,N_13705,N_13283);
nor U14247 (N_14247,N_13312,N_13452);
xor U14248 (N_14248,N_13328,N_13743);
nor U14249 (N_14249,N_13236,N_13688);
or U14250 (N_14250,N_13547,N_13475);
nor U14251 (N_14251,N_13445,N_13494);
nor U14252 (N_14252,N_13157,N_13179);
or U14253 (N_14253,N_13429,N_13732);
xor U14254 (N_14254,N_13366,N_13370);
nor U14255 (N_14255,N_13500,N_13405);
xor U14256 (N_14256,N_13526,N_13689);
nor U14257 (N_14257,N_13357,N_13190);
nand U14258 (N_14258,N_13219,N_13135);
and U14259 (N_14259,N_13494,N_13725);
nand U14260 (N_14260,N_13744,N_13255);
or U14261 (N_14261,N_13622,N_13702);
or U14262 (N_14262,N_13461,N_13316);
nor U14263 (N_14263,N_13334,N_13716);
nor U14264 (N_14264,N_13184,N_13601);
nand U14265 (N_14265,N_13201,N_13668);
nand U14266 (N_14266,N_13608,N_13308);
or U14267 (N_14267,N_13548,N_13336);
or U14268 (N_14268,N_13512,N_13215);
and U14269 (N_14269,N_13213,N_13696);
xor U14270 (N_14270,N_13717,N_13684);
nand U14271 (N_14271,N_13642,N_13184);
or U14272 (N_14272,N_13474,N_13197);
and U14273 (N_14273,N_13613,N_13256);
and U14274 (N_14274,N_13248,N_13449);
and U14275 (N_14275,N_13264,N_13730);
xnor U14276 (N_14276,N_13553,N_13219);
nand U14277 (N_14277,N_13137,N_13634);
nor U14278 (N_14278,N_13420,N_13610);
and U14279 (N_14279,N_13653,N_13577);
and U14280 (N_14280,N_13437,N_13736);
nand U14281 (N_14281,N_13389,N_13497);
nor U14282 (N_14282,N_13246,N_13276);
or U14283 (N_14283,N_13660,N_13497);
or U14284 (N_14284,N_13504,N_13725);
or U14285 (N_14285,N_13202,N_13232);
xnor U14286 (N_14286,N_13640,N_13186);
xor U14287 (N_14287,N_13723,N_13707);
and U14288 (N_14288,N_13125,N_13539);
or U14289 (N_14289,N_13450,N_13556);
or U14290 (N_14290,N_13708,N_13478);
nor U14291 (N_14291,N_13299,N_13322);
xnor U14292 (N_14292,N_13126,N_13369);
xor U14293 (N_14293,N_13598,N_13343);
and U14294 (N_14294,N_13158,N_13301);
nand U14295 (N_14295,N_13640,N_13207);
xnor U14296 (N_14296,N_13537,N_13352);
xor U14297 (N_14297,N_13283,N_13355);
or U14298 (N_14298,N_13184,N_13497);
nand U14299 (N_14299,N_13637,N_13156);
nand U14300 (N_14300,N_13472,N_13592);
and U14301 (N_14301,N_13141,N_13397);
and U14302 (N_14302,N_13622,N_13711);
xnor U14303 (N_14303,N_13437,N_13360);
nand U14304 (N_14304,N_13199,N_13400);
nand U14305 (N_14305,N_13570,N_13200);
or U14306 (N_14306,N_13590,N_13727);
nand U14307 (N_14307,N_13200,N_13426);
nor U14308 (N_14308,N_13134,N_13450);
nor U14309 (N_14309,N_13422,N_13363);
nor U14310 (N_14310,N_13197,N_13491);
nor U14311 (N_14311,N_13417,N_13401);
or U14312 (N_14312,N_13231,N_13431);
or U14313 (N_14313,N_13334,N_13689);
nor U14314 (N_14314,N_13231,N_13636);
and U14315 (N_14315,N_13402,N_13186);
xor U14316 (N_14316,N_13317,N_13333);
nor U14317 (N_14317,N_13747,N_13529);
or U14318 (N_14318,N_13362,N_13632);
nor U14319 (N_14319,N_13590,N_13323);
nand U14320 (N_14320,N_13520,N_13484);
nand U14321 (N_14321,N_13640,N_13529);
nor U14322 (N_14322,N_13747,N_13347);
and U14323 (N_14323,N_13306,N_13432);
and U14324 (N_14324,N_13166,N_13185);
or U14325 (N_14325,N_13373,N_13275);
xor U14326 (N_14326,N_13717,N_13358);
nor U14327 (N_14327,N_13261,N_13337);
and U14328 (N_14328,N_13358,N_13572);
nand U14329 (N_14329,N_13223,N_13263);
and U14330 (N_14330,N_13594,N_13319);
nor U14331 (N_14331,N_13333,N_13707);
or U14332 (N_14332,N_13707,N_13372);
or U14333 (N_14333,N_13485,N_13256);
nor U14334 (N_14334,N_13449,N_13693);
or U14335 (N_14335,N_13306,N_13668);
nand U14336 (N_14336,N_13748,N_13252);
xor U14337 (N_14337,N_13406,N_13460);
xor U14338 (N_14338,N_13527,N_13725);
or U14339 (N_14339,N_13172,N_13270);
or U14340 (N_14340,N_13558,N_13292);
nand U14341 (N_14341,N_13523,N_13617);
and U14342 (N_14342,N_13482,N_13634);
nor U14343 (N_14343,N_13665,N_13498);
xnor U14344 (N_14344,N_13256,N_13210);
nor U14345 (N_14345,N_13336,N_13640);
nand U14346 (N_14346,N_13239,N_13525);
nor U14347 (N_14347,N_13732,N_13299);
and U14348 (N_14348,N_13565,N_13432);
xor U14349 (N_14349,N_13592,N_13676);
xnor U14350 (N_14350,N_13698,N_13290);
nor U14351 (N_14351,N_13558,N_13536);
xnor U14352 (N_14352,N_13319,N_13483);
xnor U14353 (N_14353,N_13257,N_13639);
and U14354 (N_14354,N_13598,N_13420);
nor U14355 (N_14355,N_13491,N_13507);
xnor U14356 (N_14356,N_13446,N_13674);
and U14357 (N_14357,N_13578,N_13693);
nand U14358 (N_14358,N_13634,N_13341);
xor U14359 (N_14359,N_13729,N_13428);
nor U14360 (N_14360,N_13577,N_13542);
and U14361 (N_14361,N_13646,N_13317);
xnor U14362 (N_14362,N_13654,N_13328);
nor U14363 (N_14363,N_13673,N_13160);
and U14364 (N_14364,N_13645,N_13589);
nand U14365 (N_14365,N_13412,N_13546);
or U14366 (N_14366,N_13726,N_13202);
or U14367 (N_14367,N_13136,N_13381);
or U14368 (N_14368,N_13161,N_13696);
xnor U14369 (N_14369,N_13511,N_13348);
xor U14370 (N_14370,N_13724,N_13179);
and U14371 (N_14371,N_13631,N_13222);
or U14372 (N_14372,N_13740,N_13206);
or U14373 (N_14373,N_13348,N_13431);
and U14374 (N_14374,N_13335,N_13505);
or U14375 (N_14375,N_13870,N_14359);
nor U14376 (N_14376,N_14239,N_14040);
xnor U14377 (N_14377,N_13966,N_13844);
xor U14378 (N_14378,N_14159,N_14278);
nor U14379 (N_14379,N_13779,N_14092);
and U14380 (N_14380,N_13893,N_14298);
nand U14381 (N_14381,N_14149,N_13774);
and U14382 (N_14382,N_14255,N_13760);
and U14383 (N_14383,N_13951,N_13808);
nand U14384 (N_14384,N_14083,N_14288);
nor U14385 (N_14385,N_14154,N_13936);
xnor U14386 (N_14386,N_14228,N_13801);
nor U14387 (N_14387,N_13830,N_13781);
nand U14388 (N_14388,N_13850,N_14105);
nor U14389 (N_14389,N_14273,N_13916);
nand U14390 (N_14390,N_14143,N_14155);
nor U14391 (N_14391,N_14370,N_13849);
nand U14392 (N_14392,N_14295,N_14342);
xnor U14393 (N_14393,N_14189,N_13755);
and U14394 (N_14394,N_14034,N_14281);
xor U14395 (N_14395,N_13923,N_13895);
nand U14396 (N_14396,N_14223,N_14249);
xor U14397 (N_14397,N_14080,N_14247);
nor U14398 (N_14398,N_13979,N_13836);
nand U14399 (N_14399,N_13820,N_14260);
or U14400 (N_14400,N_13778,N_13752);
nor U14401 (N_14401,N_13873,N_13941);
nand U14402 (N_14402,N_13823,N_14133);
nor U14403 (N_14403,N_14325,N_14332);
xor U14404 (N_14404,N_14055,N_13783);
nand U14405 (N_14405,N_14322,N_13840);
nand U14406 (N_14406,N_13964,N_14311);
and U14407 (N_14407,N_14290,N_13950);
nor U14408 (N_14408,N_14242,N_14213);
or U14409 (N_14409,N_14024,N_14183);
nand U14410 (N_14410,N_14196,N_13970);
nand U14411 (N_14411,N_14119,N_13975);
xnor U14412 (N_14412,N_14108,N_14349);
nor U14413 (N_14413,N_14137,N_14340);
nand U14414 (N_14414,N_14018,N_14266);
nand U14415 (N_14415,N_13766,N_13938);
or U14416 (N_14416,N_13793,N_13800);
and U14417 (N_14417,N_14127,N_14148);
or U14418 (N_14418,N_14160,N_13967);
nor U14419 (N_14419,N_14103,N_13998);
nor U14420 (N_14420,N_13999,N_14304);
xor U14421 (N_14421,N_13780,N_14136);
nand U14422 (N_14422,N_13829,N_13987);
nor U14423 (N_14423,N_14036,N_13764);
nor U14424 (N_14424,N_14333,N_14202);
xor U14425 (N_14425,N_13929,N_14263);
xor U14426 (N_14426,N_13955,N_13930);
or U14427 (N_14427,N_13882,N_14369);
and U14428 (N_14428,N_13933,N_13948);
nor U14429 (N_14429,N_14162,N_13856);
or U14430 (N_14430,N_13869,N_14361);
or U14431 (N_14431,N_13953,N_14363);
or U14432 (N_14432,N_13756,N_13985);
xnor U14433 (N_14433,N_14262,N_14256);
or U14434 (N_14434,N_14171,N_14274);
nor U14435 (N_14435,N_14368,N_13903);
nand U14436 (N_14436,N_13961,N_13906);
and U14437 (N_14437,N_14205,N_14043);
nor U14438 (N_14438,N_13937,N_13886);
or U14439 (N_14439,N_13837,N_14226);
and U14440 (N_14440,N_14229,N_13811);
nand U14441 (N_14441,N_14243,N_14111);
nor U14442 (N_14442,N_14151,N_14090);
or U14443 (N_14443,N_14087,N_14291);
and U14444 (N_14444,N_14033,N_14085);
nand U14445 (N_14445,N_13843,N_14195);
nand U14446 (N_14446,N_13911,N_14230);
nor U14447 (N_14447,N_14197,N_13891);
nand U14448 (N_14448,N_14314,N_14161);
and U14449 (N_14449,N_13879,N_14364);
or U14450 (N_14450,N_13822,N_14174);
and U14451 (N_14451,N_14209,N_14061);
nand U14452 (N_14452,N_13912,N_14072);
xnor U14453 (N_14453,N_13817,N_13928);
and U14454 (N_14454,N_13942,N_14177);
nand U14455 (N_14455,N_13786,N_14146);
nor U14456 (N_14456,N_14086,N_14147);
nand U14457 (N_14457,N_14032,N_14302);
and U14458 (N_14458,N_13839,N_14301);
nand U14459 (N_14459,N_14104,N_13806);
nor U14460 (N_14460,N_14144,N_14335);
or U14461 (N_14461,N_13784,N_14344);
and U14462 (N_14462,N_13924,N_14283);
nand U14463 (N_14463,N_14201,N_14084);
nor U14464 (N_14464,N_14128,N_14267);
xnor U14465 (N_14465,N_13842,N_14300);
or U14466 (N_14466,N_14020,N_14169);
xor U14467 (N_14467,N_14294,N_13767);
or U14468 (N_14468,N_13976,N_14096);
xnor U14469 (N_14469,N_13994,N_14038);
xor U14470 (N_14470,N_14269,N_13954);
or U14471 (N_14471,N_14270,N_14234);
xor U14472 (N_14472,N_13835,N_14303);
xor U14473 (N_14473,N_14088,N_13887);
nor U14474 (N_14474,N_13900,N_14132);
nand U14475 (N_14475,N_14225,N_14187);
nor U14476 (N_14476,N_13847,N_14012);
nand U14477 (N_14477,N_13914,N_14232);
or U14478 (N_14478,N_14045,N_14006);
or U14479 (N_14479,N_14318,N_14091);
nand U14480 (N_14480,N_14082,N_14221);
nor U14481 (N_14481,N_13771,N_13932);
and U14482 (N_14482,N_13946,N_14079);
xnor U14483 (N_14483,N_14337,N_14323);
nand U14484 (N_14484,N_14233,N_14317);
xnor U14485 (N_14485,N_13889,N_13880);
or U14486 (N_14486,N_14305,N_14178);
nand U14487 (N_14487,N_14078,N_13805);
xnor U14488 (N_14488,N_14007,N_14170);
nor U14489 (N_14489,N_14074,N_14003);
and U14490 (N_14490,N_14109,N_14194);
and U14491 (N_14491,N_14345,N_14009);
or U14492 (N_14492,N_13992,N_14004);
and U14493 (N_14493,N_14354,N_14126);
xnor U14494 (N_14494,N_13995,N_13958);
nand U14495 (N_14495,N_13753,N_14293);
xor U14496 (N_14496,N_14113,N_14060);
or U14497 (N_14497,N_13794,N_13819);
nor U14498 (N_14498,N_13990,N_14048);
xor U14499 (N_14499,N_13918,N_13775);
nor U14500 (N_14500,N_14210,N_13768);
nor U14501 (N_14501,N_14265,N_14041);
xnor U14502 (N_14502,N_14276,N_14238);
or U14503 (N_14503,N_14185,N_13861);
nor U14504 (N_14504,N_13845,N_14330);
nand U14505 (N_14505,N_14026,N_14331);
or U14506 (N_14506,N_14095,N_14106);
nand U14507 (N_14507,N_14181,N_13892);
nor U14508 (N_14508,N_14125,N_13792);
xor U14509 (N_14509,N_14164,N_13832);
and U14510 (N_14510,N_14219,N_14321);
nor U14511 (N_14511,N_14207,N_14039);
or U14512 (N_14512,N_13877,N_13790);
or U14513 (N_14513,N_13934,N_14044);
and U14514 (N_14514,N_14138,N_14114);
and U14515 (N_14515,N_14351,N_13859);
xor U14516 (N_14516,N_14237,N_14203);
or U14517 (N_14517,N_14051,N_14107);
xor U14518 (N_14518,N_14120,N_13831);
nor U14519 (N_14519,N_14259,N_14258);
or U14520 (N_14520,N_14081,N_13919);
xor U14521 (N_14521,N_14112,N_13782);
or U14522 (N_14522,N_14235,N_14002);
nor U14523 (N_14523,N_14328,N_14165);
and U14524 (N_14524,N_13864,N_14073);
and U14525 (N_14525,N_13988,N_14347);
xor U14526 (N_14526,N_14271,N_14116);
and U14527 (N_14527,N_14017,N_13812);
nand U14528 (N_14528,N_14299,N_14310);
or U14529 (N_14529,N_14182,N_14327);
xnor U14530 (N_14530,N_13815,N_14070);
nand U14531 (N_14531,N_13917,N_14215);
or U14532 (N_14532,N_14252,N_14275);
xnor U14533 (N_14533,N_13834,N_14062);
or U14534 (N_14534,N_13857,N_14069);
nor U14535 (N_14535,N_13980,N_14035);
and U14536 (N_14536,N_13876,N_13777);
nand U14537 (N_14537,N_14348,N_13810);
nor U14538 (N_14538,N_13972,N_13789);
and U14539 (N_14539,N_14218,N_14067);
xor U14540 (N_14540,N_13996,N_14150);
nor U14541 (N_14541,N_14102,N_14071);
and U14542 (N_14542,N_14157,N_14167);
nand U14543 (N_14543,N_13796,N_14287);
and U14544 (N_14544,N_13776,N_13982);
or U14545 (N_14545,N_14272,N_14145);
or U14546 (N_14546,N_14312,N_14118);
nor U14547 (N_14547,N_14190,N_14339);
nor U14548 (N_14548,N_14297,N_13909);
or U14549 (N_14549,N_14058,N_13927);
or U14550 (N_14550,N_14122,N_13825);
xnor U14551 (N_14551,N_13883,N_13787);
and U14552 (N_14552,N_13875,N_13904);
nand U14553 (N_14553,N_13798,N_14098);
nand U14554 (N_14554,N_14284,N_14204);
or U14555 (N_14555,N_13993,N_13974);
nand U14556 (N_14556,N_14176,N_13940);
nor U14557 (N_14557,N_13908,N_14306);
xnor U14558 (N_14558,N_14329,N_14357);
or U14559 (N_14559,N_14254,N_14101);
nand U14560 (N_14560,N_13898,N_13939);
nand U14561 (N_14561,N_14001,N_13751);
nor U14562 (N_14562,N_14343,N_13971);
nand U14563 (N_14563,N_13920,N_13865);
and U14564 (N_14564,N_13986,N_14015);
nand U14565 (N_14565,N_13969,N_14248);
nand U14566 (N_14566,N_13977,N_14000);
nor U14567 (N_14567,N_13788,N_14372);
xnor U14568 (N_14568,N_14246,N_14313);
nor U14569 (N_14569,N_13899,N_14139);
and U14570 (N_14570,N_14292,N_14030);
nor U14571 (N_14571,N_14053,N_14336);
nand U14572 (N_14572,N_13821,N_13943);
nand U14573 (N_14573,N_14175,N_14141);
nand U14574 (N_14574,N_13897,N_13769);
xnor U14575 (N_14575,N_14140,N_13905);
and U14576 (N_14576,N_14217,N_14153);
xor U14577 (N_14577,N_13824,N_13838);
xor U14578 (N_14578,N_13926,N_13795);
nor U14579 (N_14579,N_13809,N_14192);
nand U14580 (N_14580,N_13852,N_13956);
nor U14581 (N_14581,N_13791,N_13846);
and U14582 (N_14582,N_13848,N_13931);
or U14583 (N_14583,N_14059,N_14289);
nor U14584 (N_14584,N_14022,N_14050);
nand U14585 (N_14585,N_14063,N_14123);
and U14586 (N_14586,N_14367,N_14316);
xnor U14587 (N_14587,N_13758,N_14068);
nor U14588 (N_14588,N_13807,N_13759);
and U14589 (N_14589,N_14152,N_14186);
nand U14590 (N_14590,N_14191,N_14163);
or U14591 (N_14591,N_14200,N_13989);
xnor U14592 (N_14592,N_14031,N_14110);
nor U14593 (N_14593,N_14180,N_14064);
and U14594 (N_14594,N_14097,N_14326);
nand U14595 (N_14595,N_13827,N_14264);
xor U14596 (N_14596,N_14135,N_13997);
nor U14597 (N_14597,N_14168,N_13978);
nand U14598 (N_14598,N_13896,N_14014);
or U14599 (N_14599,N_13902,N_13773);
or U14600 (N_14600,N_14253,N_14371);
nor U14601 (N_14601,N_13858,N_14353);
and U14602 (N_14602,N_14358,N_14296);
xor U14603 (N_14603,N_14027,N_14241);
and U14604 (N_14604,N_13947,N_13890);
and U14605 (N_14605,N_13874,N_13866);
or U14606 (N_14606,N_13828,N_14016);
or U14607 (N_14607,N_13913,N_14057);
xnor U14608 (N_14608,N_14021,N_13944);
nand U14609 (N_14609,N_14356,N_14355);
and U14610 (N_14610,N_14240,N_14037);
nor U14611 (N_14611,N_14352,N_13772);
and U14612 (N_14612,N_14010,N_13885);
or U14613 (N_14613,N_14156,N_14268);
nor U14614 (N_14614,N_14320,N_14013);
nand U14615 (N_14615,N_14066,N_14220);
or U14616 (N_14616,N_13915,N_13816);
and U14617 (N_14617,N_13888,N_14334);
nor U14618 (N_14618,N_13762,N_14261);
or U14619 (N_14619,N_14236,N_14075);
and U14620 (N_14620,N_14172,N_14341);
nor U14621 (N_14621,N_14179,N_13826);
and U14622 (N_14622,N_14129,N_13963);
nand U14623 (N_14623,N_14028,N_14280);
or U14624 (N_14624,N_13814,N_13818);
and U14625 (N_14625,N_14224,N_14056);
xor U14626 (N_14626,N_13991,N_14042);
and U14627 (N_14627,N_14047,N_13854);
and U14628 (N_14628,N_14094,N_14115);
and U14629 (N_14629,N_13853,N_13871);
or U14630 (N_14630,N_13894,N_13922);
xnor U14631 (N_14631,N_14309,N_14023);
nor U14632 (N_14632,N_14319,N_14231);
or U14633 (N_14633,N_14245,N_14227);
xnor U14634 (N_14634,N_14025,N_14046);
or U14635 (N_14635,N_14124,N_14131);
nor U14636 (N_14636,N_13921,N_14099);
and U14637 (N_14637,N_13884,N_14208);
nand U14638 (N_14638,N_14360,N_14324);
nor U14639 (N_14639,N_13945,N_13878);
nand U14640 (N_14640,N_14166,N_14308);
nor U14641 (N_14641,N_13833,N_14049);
or U14642 (N_14642,N_14338,N_13925);
xnor U14643 (N_14643,N_14282,N_14285);
nand U14644 (N_14644,N_13962,N_13881);
and U14645 (N_14645,N_13959,N_14065);
or U14646 (N_14646,N_14011,N_13949);
xor U14647 (N_14647,N_14173,N_13804);
nor U14648 (N_14648,N_13935,N_14286);
xnor U14649 (N_14649,N_13797,N_13754);
xor U14650 (N_14650,N_13952,N_13770);
and U14651 (N_14651,N_13855,N_13867);
nand U14652 (N_14652,N_14193,N_13802);
nor U14653 (N_14653,N_13901,N_14257);
or U14654 (N_14654,N_13984,N_13860);
xor U14655 (N_14655,N_14093,N_14373);
xor U14656 (N_14656,N_14008,N_14222);
nand U14657 (N_14657,N_13813,N_14052);
and U14658 (N_14658,N_14198,N_14362);
or U14659 (N_14659,N_14250,N_14130);
and U14660 (N_14660,N_13960,N_13965);
or U14661 (N_14661,N_14346,N_14244);
nand U14662 (N_14662,N_13799,N_14100);
nor U14663 (N_14663,N_14214,N_13863);
and U14664 (N_14664,N_14350,N_13968);
xnor U14665 (N_14665,N_14206,N_13750);
xor U14666 (N_14666,N_14216,N_14117);
or U14667 (N_14667,N_13910,N_14315);
and U14668 (N_14668,N_13803,N_14251);
nand U14669 (N_14669,N_13957,N_13907);
xnor U14670 (N_14670,N_14029,N_14077);
xnor U14671 (N_14671,N_13851,N_13862);
nand U14672 (N_14672,N_14365,N_14279);
and U14673 (N_14673,N_13841,N_14005);
or U14674 (N_14674,N_14307,N_13983);
and U14675 (N_14675,N_14076,N_14211);
nor U14676 (N_14676,N_14366,N_14374);
nand U14677 (N_14677,N_13872,N_14134);
or U14678 (N_14678,N_14019,N_14121);
xnor U14679 (N_14679,N_13765,N_14277);
or U14680 (N_14680,N_13763,N_13785);
or U14681 (N_14681,N_13981,N_13761);
or U14682 (N_14682,N_14054,N_14158);
and U14683 (N_14683,N_14089,N_13868);
nand U14684 (N_14684,N_14199,N_14142);
xnor U14685 (N_14685,N_13757,N_14212);
xor U14686 (N_14686,N_14184,N_14188);
and U14687 (N_14687,N_13973,N_13764);
xnor U14688 (N_14688,N_13796,N_14113);
nand U14689 (N_14689,N_13877,N_14298);
and U14690 (N_14690,N_14038,N_13859);
or U14691 (N_14691,N_13920,N_13984);
or U14692 (N_14692,N_14158,N_14194);
xnor U14693 (N_14693,N_14084,N_14333);
nor U14694 (N_14694,N_14148,N_14361);
or U14695 (N_14695,N_13890,N_14254);
xor U14696 (N_14696,N_13806,N_14302);
or U14697 (N_14697,N_13927,N_13898);
and U14698 (N_14698,N_14242,N_14156);
xor U14699 (N_14699,N_14018,N_14109);
or U14700 (N_14700,N_13863,N_13950);
or U14701 (N_14701,N_14218,N_13884);
xor U14702 (N_14702,N_13773,N_14203);
and U14703 (N_14703,N_14182,N_14064);
xnor U14704 (N_14704,N_13881,N_13854);
nor U14705 (N_14705,N_14176,N_14341);
or U14706 (N_14706,N_13837,N_13961);
nor U14707 (N_14707,N_14237,N_13967);
nand U14708 (N_14708,N_13799,N_13797);
xnor U14709 (N_14709,N_14243,N_14361);
xnor U14710 (N_14710,N_13867,N_13866);
nor U14711 (N_14711,N_14168,N_13939);
nand U14712 (N_14712,N_13780,N_14249);
and U14713 (N_14713,N_14067,N_13802);
nand U14714 (N_14714,N_14361,N_14236);
nand U14715 (N_14715,N_14040,N_14269);
nor U14716 (N_14716,N_14230,N_14074);
and U14717 (N_14717,N_13966,N_14189);
xnor U14718 (N_14718,N_14049,N_14072);
or U14719 (N_14719,N_13802,N_14153);
and U14720 (N_14720,N_14014,N_13953);
and U14721 (N_14721,N_14199,N_14215);
and U14722 (N_14722,N_14018,N_13956);
nor U14723 (N_14723,N_14154,N_13802);
xnor U14724 (N_14724,N_14323,N_14310);
nor U14725 (N_14725,N_13922,N_13869);
and U14726 (N_14726,N_13926,N_13964);
xor U14727 (N_14727,N_13797,N_14198);
or U14728 (N_14728,N_14061,N_14269);
nand U14729 (N_14729,N_14253,N_14074);
xor U14730 (N_14730,N_14306,N_13993);
nor U14731 (N_14731,N_14372,N_14084);
xnor U14732 (N_14732,N_13837,N_13763);
and U14733 (N_14733,N_13917,N_13830);
xnor U14734 (N_14734,N_13854,N_14344);
nor U14735 (N_14735,N_13896,N_13917);
xor U14736 (N_14736,N_14173,N_14078);
nor U14737 (N_14737,N_14000,N_14001);
nand U14738 (N_14738,N_13977,N_14365);
nor U14739 (N_14739,N_14219,N_14216);
nand U14740 (N_14740,N_14067,N_14043);
xnor U14741 (N_14741,N_13774,N_13996);
nand U14742 (N_14742,N_14049,N_14088);
and U14743 (N_14743,N_14160,N_13783);
xnor U14744 (N_14744,N_13805,N_14361);
nand U14745 (N_14745,N_14163,N_14245);
nor U14746 (N_14746,N_14115,N_14206);
and U14747 (N_14747,N_13906,N_13960);
nor U14748 (N_14748,N_13831,N_14055);
nand U14749 (N_14749,N_14374,N_14302);
nand U14750 (N_14750,N_13870,N_13774);
nor U14751 (N_14751,N_13825,N_14094);
xor U14752 (N_14752,N_13901,N_14291);
nand U14753 (N_14753,N_14019,N_14115);
nand U14754 (N_14754,N_14355,N_13885);
nand U14755 (N_14755,N_14152,N_14089);
xor U14756 (N_14756,N_14302,N_14171);
and U14757 (N_14757,N_14132,N_14130);
or U14758 (N_14758,N_14089,N_14335);
xor U14759 (N_14759,N_14013,N_14367);
and U14760 (N_14760,N_14103,N_14301);
or U14761 (N_14761,N_13770,N_14031);
and U14762 (N_14762,N_13947,N_13907);
xnor U14763 (N_14763,N_13911,N_14319);
nand U14764 (N_14764,N_14208,N_14310);
and U14765 (N_14765,N_14156,N_14012);
xnor U14766 (N_14766,N_14165,N_14170);
nand U14767 (N_14767,N_14216,N_14249);
xor U14768 (N_14768,N_14057,N_14034);
or U14769 (N_14769,N_14348,N_14314);
nor U14770 (N_14770,N_13842,N_14338);
xnor U14771 (N_14771,N_13931,N_13775);
xor U14772 (N_14772,N_13978,N_14350);
nand U14773 (N_14773,N_13842,N_14099);
nand U14774 (N_14774,N_13820,N_14333);
nor U14775 (N_14775,N_14207,N_13764);
or U14776 (N_14776,N_14051,N_14055);
xnor U14777 (N_14777,N_14203,N_14011);
xnor U14778 (N_14778,N_14017,N_14082);
or U14779 (N_14779,N_14112,N_14301);
or U14780 (N_14780,N_13930,N_13877);
or U14781 (N_14781,N_13769,N_14306);
or U14782 (N_14782,N_13886,N_14062);
or U14783 (N_14783,N_14101,N_13809);
xnor U14784 (N_14784,N_13994,N_14370);
xor U14785 (N_14785,N_13768,N_14134);
nand U14786 (N_14786,N_14337,N_14028);
xor U14787 (N_14787,N_14269,N_14338);
xnor U14788 (N_14788,N_13771,N_13927);
nor U14789 (N_14789,N_14337,N_14228);
nor U14790 (N_14790,N_14342,N_13939);
nand U14791 (N_14791,N_13751,N_13929);
or U14792 (N_14792,N_13750,N_14358);
nor U14793 (N_14793,N_14367,N_14031);
nand U14794 (N_14794,N_14311,N_14167);
and U14795 (N_14795,N_13951,N_13800);
or U14796 (N_14796,N_14189,N_14001);
and U14797 (N_14797,N_14363,N_14305);
nor U14798 (N_14798,N_13813,N_14161);
nor U14799 (N_14799,N_14204,N_13989);
or U14800 (N_14800,N_14180,N_14254);
nand U14801 (N_14801,N_13935,N_14290);
and U14802 (N_14802,N_14263,N_14213);
xor U14803 (N_14803,N_13822,N_13891);
nand U14804 (N_14804,N_13930,N_13918);
xor U14805 (N_14805,N_13974,N_14328);
xor U14806 (N_14806,N_14354,N_13980);
nor U14807 (N_14807,N_13983,N_14185);
xor U14808 (N_14808,N_13779,N_14156);
and U14809 (N_14809,N_14226,N_14258);
or U14810 (N_14810,N_14007,N_14302);
xor U14811 (N_14811,N_13884,N_14117);
nand U14812 (N_14812,N_14008,N_13997);
nor U14813 (N_14813,N_14252,N_14360);
nand U14814 (N_14814,N_13806,N_14324);
nand U14815 (N_14815,N_14185,N_14209);
xor U14816 (N_14816,N_14229,N_14200);
nand U14817 (N_14817,N_14205,N_14282);
nor U14818 (N_14818,N_13817,N_13923);
nor U14819 (N_14819,N_14173,N_14213);
nand U14820 (N_14820,N_14036,N_13827);
and U14821 (N_14821,N_13844,N_14211);
and U14822 (N_14822,N_14257,N_13935);
or U14823 (N_14823,N_14212,N_13906);
xor U14824 (N_14824,N_14062,N_14159);
and U14825 (N_14825,N_14033,N_14147);
nand U14826 (N_14826,N_13988,N_13753);
nand U14827 (N_14827,N_14270,N_13773);
xor U14828 (N_14828,N_13993,N_13956);
nand U14829 (N_14829,N_14291,N_13898);
nor U14830 (N_14830,N_13864,N_14085);
nand U14831 (N_14831,N_14346,N_13793);
or U14832 (N_14832,N_14092,N_13861);
or U14833 (N_14833,N_13940,N_13760);
nor U14834 (N_14834,N_13880,N_14181);
and U14835 (N_14835,N_13828,N_14344);
nand U14836 (N_14836,N_14186,N_14333);
nand U14837 (N_14837,N_13827,N_14093);
and U14838 (N_14838,N_14208,N_14282);
and U14839 (N_14839,N_14050,N_14101);
nor U14840 (N_14840,N_14264,N_14017);
and U14841 (N_14841,N_14141,N_14096);
xnor U14842 (N_14842,N_14101,N_14323);
nor U14843 (N_14843,N_14060,N_14039);
nor U14844 (N_14844,N_14111,N_14312);
nand U14845 (N_14845,N_13836,N_13787);
and U14846 (N_14846,N_14248,N_14311);
or U14847 (N_14847,N_13751,N_13928);
nand U14848 (N_14848,N_13897,N_14321);
xnor U14849 (N_14849,N_14237,N_14319);
xor U14850 (N_14850,N_13925,N_13928);
or U14851 (N_14851,N_14273,N_13949);
or U14852 (N_14852,N_14268,N_13848);
nand U14853 (N_14853,N_14115,N_14044);
nand U14854 (N_14854,N_13834,N_14103);
xnor U14855 (N_14855,N_14273,N_13991);
nand U14856 (N_14856,N_13978,N_14149);
nand U14857 (N_14857,N_13900,N_14024);
nand U14858 (N_14858,N_13910,N_14222);
nor U14859 (N_14859,N_14370,N_14213);
xor U14860 (N_14860,N_14096,N_13964);
or U14861 (N_14861,N_13883,N_13825);
and U14862 (N_14862,N_13887,N_14154);
or U14863 (N_14863,N_14252,N_13933);
nor U14864 (N_14864,N_14195,N_13897);
xor U14865 (N_14865,N_13900,N_14142);
and U14866 (N_14866,N_14374,N_14206);
xnor U14867 (N_14867,N_14197,N_14203);
nor U14868 (N_14868,N_14309,N_14324);
nand U14869 (N_14869,N_14290,N_13967);
or U14870 (N_14870,N_14124,N_14286);
nor U14871 (N_14871,N_13835,N_13899);
or U14872 (N_14872,N_13750,N_14041);
and U14873 (N_14873,N_14199,N_13905);
and U14874 (N_14874,N_14363,N_14049);
nor U14875 (N_14875,N_14249,N_14232);
xnor U14876 (N_14876,N_13785,N_14319);
nor U14877 (N_14877,N_13949,N_13782);
nor U14878 (N_14878,N_14106,N_14013);
nor U14879 (N_14879,N_14159,N_13832);
nor U14880 (N_14880,N_13773,N_14275);
xor U14881 (N_14881,N_14329,N_14178);
nand U14882 (N_14882,N_13789,N_13943);
xor U14883 (N_14883,N_14150,N_13955);
nor U14884 (N_14884,N_14362,N_14317);
nor U14885 (N_14885,N_14316,N_14264);
and U14886 (N_14886,N_13807,N_14045);
or U14887 (N_14887,N_14108,N_14103);
or U14888 (N_14888,N_14354,N_14127);
nand U14889 (N_14889,N_13875,N_14011);
xor U14890 (N_14890,N_14208,N_14242);
nand U14891 (N_14891,N_13938,N_13926);
xor U14892 (N_14892,N_13867,N_13993);
nand U14893 (N_14893,N_13937,N_13764);
and U14894 (N_14894,N_14003,N_13837);
or U14895 (N_14895,N_14242,N_13967);
nor U14896 (N_14896,N_13984,N_13958);
xor U14897 (N_14897,N_14075,N_14273);
xnor U14898 (N_14898,N_14203,N_13844);
nand U14899 (N_14899,N_14101,N_13866);
xor U14900 (N_14900,N_13818,N_13994);
nor U14901 (N_14901,N_14131,N_14140);
nand U14902 (N_14902,N_14358,N_13916);
nand U14903 (N_14903,N_13790,N_13958);
or U14904 (N_14904,N_14140,N_14238);
and U14905 (N_14905,N_13960,N_13929);
nand U14906 (N_14906,N_13808,N_14173);
nor U14907 (N_14907,N_14100,N_14098);
nand U14908 (N_14908,N_14019,N_14108);
nor U14909 (N_14909,N_14204,N_14144);
xor U14910 (N_14910,N_14264,N_14120);
nand U14911 (N_14911,N_13839,N_13943);
or U14912 (N_14912,N_14237,N_14016);
nand U14913 (N_14913,N_14113,N_13770);
and U14914 (N_14914,N_14021,N_14049);
and U14915 (N_14915,N_14302,N_13785);
nor U14916 (N_14916,N_14182,N_13831);
nand U14917 (N_14917,N_13788,N_14178);
xnor U14918 (N_14918,N_14017,N_13866);
nor U14919 (N_14919,N_14239,N_14253);
nor U14920 (N_14920,N_13968,N_13796);
nor U14921 (N_14921,N_14077,N_13840);
and U14922 (N_14922,N_14008,N_14357);
nor U14923 (N_14923,N_14059,N_13793);
nor U14924 (N_14924,N_14131,N_13959);
nand U14925 (N_14925,N_14017,N_13762);
nor U14926 (N_14926,N_13941,N_14331);
xor U14927 (N_14927,N_13801,N_14210);
nand U14928 (N_14928,N_13984,N_13854);
nor U14929 (N_14929,N_13865,N_14055);
nand U14930 (N_14930,N_14015,N_13881);
nand U14931 (N_14931,N_14309,N_14164);
and U14932 (N_14932,N_14226,N_14199);
nand U14933 (N_14933,N_13802,N_14042);
or U14934 (N_14934,N_14260,N_14116);
and U14935 (N_14935,N_14237,N_13776);
and U14936 (N_14936,N_14141,N_14256);
and U14937 (N_14937,N_14347,N_14247);
nand U14938 (N_14938,N_14016,N_14104);
nand U14939 (N_14939,N_14350,N_13827);
xor U14940 (N_14940,N_14039,N_13963);
xor U14941 (N_14941,N_13892,N_13806);
or U14942 (N_14942,N_13915,N_14167);
nor U14943 (N_14943,N_13891,N_14038);
or U14944 (N_14944,N_13914,N_14363);
nor U14945 (N_14945,N_14225,N_14146);
or U14946 (N_14946,N_14319,N_14243);
nand U14947 (N_14947,N_13959,N_14128);
nor U14948 (N_14948,N_14327,N_14245);
nand U14949 (N_14949,N_14348,N_14252);
nand U14950 (N_14950,N_14358,N_14172);
nand U14951 (N_14951,N_14329,N_14313);
or U14952 (N_14952,N_13874,N_13938);
or U14953 (N_14953,N_14353,N_13965);
xor U14954 (N_14954,N_13781,N_13998);
xnor U14955 (N_14955,N_14067,N_14216);
and U14956 (N_14956,N_13760,N_13996);
or U14957 (N_14957,N_14182,N_14374);
or U14958 (N_14958,N_13946,N_13965);
and U14959 (N_14959,N_13885,N_13985);
nand U14960 (N_14960,N_13933,N_14126);
nand U14961 (N_14961,N_14002,N_13874);
and U14962 (N_14962,N_14045,N_14254);
and U14963 (N_14963,N_14167,N_14282);
xnor U14964 (N_14964,N_14270,N_13909);
nand U14965 (N_14965,N_14365,N_13882);
and U14966 (N_14966,N_13885,N_14135);
or U14967 (N_14967,N_13794,N_13956);
nand U14968 (N_14968,N_14206,N_13793);
xnor U14969 (N_14969,N_13829,N_14168);
xor U14970 (N_14970,N_14293,N_14145);
nand U14971 (N_14971,N_14317,N_14237);
xor U14972 (N_14972,N_13827,N_13953);
xor U14973 (N_14973,N_13929,N_14005);
and U14974 (N_14974,N_14166,N_14091);
xnor U14975 (N_14975,N_14203,N_13809);
or U14976 (N_14976,N_13911,N_14181);
or U14977 (N_14977,N_14001,N_14266);
nand U14978 (N_14978,N_13834,N_14045);
xnor U14979 (N_14979,N_13756,N_14243);
nor U14980 (N_14980,N_14215,N_14246);
nand U14981 (N_14981,N_13782,N_14118);
nor U14982 (N_14982,N_13751,N_13852);
nand U14983 (N_14983,N_13921,N_13944);
or U14984 (N_14984,N_14164,N_13792);
nand U14985 (N_14985,N_14281,N_13814);
nand U14986 (N_14986,N_14111,N_14295);
xor U14987 (N_14987,N_13797,N_13785);
and U14988 (N_14988,N_13999,N_14111);
and U14989 (N_14989,N_14114,N_13772);
or U14990 (N_14990,N_14156,N_13973);
nor U14991 (N_14991,N_14204,N_13792);
and U14992 (N_14992,N_13773,N_13952);
nand U14993 (N_14993,N_14335,N_14204);
xor U14994 (N_14994,N_13757,N_13899);
nor U14995 (N_14995,N_14371,N_13849);
or U14996 (N_14996,N_14062,N_13962);
and U14997 (N_14997,N_14309,N_14077);
xnor U14998 (N_14998,N_13987,N_14019);
xnor U14999 (N_14999,N_13778,N_14341);
nand U15000 (N_15000,N_14609,N_14516);
nor U15001 (N_15001,N_14753,N_14721);
and U15002 (N_15002,N_14934,N_14485);
and U15003 (N_15003,N_14462,N_14690);
or U15004 (N_15004,N_14428,N_14617);
nand U15005 (N_15005,N_14977,N_14730);
xnor U15006 (N_15006,N_14455,N_14954);
xnor U15007 (N_15007,N_14863,N_14830);
nand U15008 (N_15008,N_14917,N_14420);
xnor U15009 (N_15009,N_14435,N_14519);
or U15010 (N_15010,N_14590,N_14601);
or U15011 (N_15011,N_14566,N_14491);
nand U15012 (N_15012,N_14665,N_14377);
nand U15013 (N_15013,N_14962,N_14430);
nor U15014 (N_15014,N_14391,N_14952);
xnor U15015 (N_15015,N_14569,N_14828);
or U15016 (N_15016,N_14671,N_14771);
or U15017 (N_15017,N_14551,N_14549);
nand U15018 (N_15018,N_14965,N_14740);
and U15019 (N_15019,N_14788,N_14417);
and U15020 (N_15020,N_14759,N_14966);
nor U15021 (N_15021,N_14660,N_14736);
and U15022 (N_15022,N_14628,N_14638);
nor U15023 (N_15023,N_14780,N_14945);
and U15024 (N_15024,N_14472,N_14726);
xor U15025 (N_15025,N_14802,N_14614);
nand U15026 (N_15026,N_14879,N_14973);
and U15027 (N_15027,N_14513,N_14559);
or U15028 (N_15028,N_14826,N_14884);
nor U15029 (N_15029,N_14764,N_14910);
xor U15030 (N_15030,N_14637,N_14866);
or U15031 (N_15031,N_14935,N_14448);
and U15032 (N_15032,N_14747,N_14573);
nand U15033 (N_15033,N_14518,N_14475);
nor U15034 (N_15034,N_14508,N_14806);
or U15035 (N_15035,N_14631,N_14745);
nor U15036 (N_15036,N_14613,N_14693);
nand U15037 (N_15037,N_14615,N_14750);
or U15038 (N_15038,N_14585,N_14733);
or U15039 (N_15039,N_14798,N_14422);
or U15040 (N_15040,N_14525,N_14932);
xor U15041 (N_15041,N_14507,N_14488);
xnor U15042 (N_15042,N_14790,N_14535);
or U15043 (N_15043,N_14594,N_14844);
nor U15044 (N_15044,N_14816,N_14849);
nor U15045 (N_15045,N_14451,N_14714);
nor U15046 (N_15046,N_14527,N_14871);
or U15047 (N_15047,N_14443,N_14540);
and U15048 (N_15048,N_14689,N_14860);
nand U15049 (N_15049,N_14599,N_14602);
or U15050 (N_15050,N_14376,N_14592);
and U15051 (N_15051,N_14713,N_14735);
xnor U15052 (N_15052,N_14784,N_14562);
nor U15053 (N_15053,N_14738,N_14471);
xnor U15054 (N_15054,N_14496,N_14388);
xnor U15055 (N_15055,N_14839,N_14758);
xor U15056 (N_15056,N_14743,N_14916);
nor U15057 (N_15057,N_14545,N_14749);
and U15058 (N_15058,N_14792,N_14949);
nand U15059 (N_15059,N_14703,N_14897);
nor U15060 (N_15060,N_14850,N_14589);
or U15061 (N_15061,N_14990,N_14930);
and U15062 (N_15062,N_14940,N_14924);
xor U15063 (N_15063,N_14567,N_14554);
nor U15064 (N_15064,N_14546,N_14464);
nor U15065 (N_15065,N_14861,N_14881);
nor U15066 (N_15066,N_14395,N_14429);
or U15067 (N_15067,N_14803,N_14505);
xor U15068 (N_15068,N_14553,N_14494);
nand U15069 (N_15069,N_14538,N_14622);
xor U15070 (N_15070,N_14982,N_14819);
xor U15071 (N_15071,N_14958,N_14676);
nand U15072 (N_15072,N_14560,N_14704);
xor U15073 (N_15073,N_14920,N_14829);
or U15074 (N_15074,N_14517,N_14768);
nor U15075 (N_15075,N_14851,N_14423);
xnor U15076 (N_15076,N_14766,N_14441);
and U15077 (N_15077,N_14859,N_14805);
nand U15078 (N_15078,N_14978,N_14607);
and U15079 (N_15079,N_14827,N_14985);
xnor U15080 (N_15080,N_14765,N_14655);
nand U15081 (N_15081,N_14797,N_14993);
and U15082 (N_15082,N_14390,N_14754);
and U15083 (N_15083,N_14409,N_14720);
xor U15084 (N_15084,N_14571,N_14588);
xnor U15085 (N_15085,N_14634,N_14817);
and U15086 (N_15086,N_14999,N_14983);
or U15087 (N_15087,N_14731,N_14656);
nor U15088 (N_15088,N_14433,N_14465);
xnor U15089 (N_15089,N_14980,N_14652);
and U15090 (N_15090,N_14532,N_14635);
nand U15091 (N_15091,N_14431,N_14833);
xnor U15092 (N_15092,N_14523,N_14846);
and U15093 (N_15093,N_14490,N_14909);
nand U15094 (N_15094,N_14456,N_14555);
xor U15095 (N_15095,N_14639,N_14457);
nand U15096 (N_15096,N_14883,N_14436);
xnor U15097 (N_15097,N_14875,N_14831);
or U15098 (N_15098,N_14419,N_14579);
nor U15099 (N_15099,N_14936,N_14595);
and U15100 (N_15100,N_14823,N_14591);
nand U15101 (N_15101,N_14636,N_14653);
xor U15102 (N_15102,N_14610,N_14459);
xor U15103 (N_15103,N_14596,N_14537);
nor U15104 (N_15104,N_14862,N_14813);
and U15105 (N_15105,N_14915,N_14408);
nand U15106 (N_15106,N_14677,N_14556);
xnor U15107 (N_15107,N_14401,N_14892);
and U15108 (N_15108,N_14375,N_14629);
or U15109 (N_15109,N_14383,N_14520);
or U15110 (N_15110,N_14974,N_14927);
and U15111 (N_15111,N_14895,N_14522);
or U15112 (N_15112,N_14643,N_14509);
nor U15113 (N_15113,N_14761,N_14845);
and U15114 (N_15114,N_14841,N_14900);
and U15115 (N_15115,N_14769,N_14432);
xor U15116 (N_15116,N_14723,N_14427);
nor U15117 (N_15117,N_14529,N_14382);
nand U15118 (N_15118,N_14378,N_14387);
or U15119 (N_15119,N_14715,N_14548);
or U15120 (N_15120,N_14577,N_14558);
nor U15121 (N_15121,N_14698,N_14728);
nor U15122 (N_15122,N_14804,N_14692);
xor U15123 (N_15123,N_14458,N_14774);
and U15124 (N_15124,N_14604,N_14557);
nor U15125 (N_15125,N_14739,N_14444);
nand U15126 (N_15126,N_14493,N_14843);
xnor U15127 (N_15127,N_14953,N_14442);
nor U15128 (N_15128,N_14872,N_14778);
or U15129 (N_15129,N_14515,N_14770);
nor U15130 (N_15130,N_14623,N_14482);
or U15131 (N_15131,N_14822,N_14908);
and U15132 (N_15132,N_14938,N_14873);
nand U15133 (N_15133,N_14956,N_14729);
nand U15134 (N_15134,N_14572,N_14789);
nand U15135 (N_15135,N_14439,N_14886);
or U15136 (N_15136,N_14394,N_14959);
or U15137 (N_15137,N_14811,N_14600);
or U15138 (N_15138,N_14645,N_14521);
nand U15139 (N_15139,N_14800,N_14763);
xnor U15140 (N_15140,N_14412,N_14842);
xor U15141 (N_15141,N_14624,N_14466);
nor U15142 (N_15142,N_14732,N_14404);
and U15143 (N_15143,N_14975,N_14389);
nor U15144 (N_15144,N_14746,N_14552);
nand U15145 (N_15145,N_14603,N_14476);
or U15146 (N_15146,N_14406,N_14633);
and U15147 (N_15147,N_14669,N_14987);
nand U15148 (N_15148,N_14699,N_14434);
and U15149 (N_15149,N_14834,N_14744);
nor U15150 (N_15150,N_14481,N_14837);
nand U15151 (N_15151,N_14649,N_14384);
xor U15152 (N_15152,N_14898,N_14996);
and U15153 (N_15153,N_14461,N_14473);
or U15154 (N_15154,N_14812,N_14957);
xor U15155 (N_15155,N_14495,N_14685);
nor U15156 (N_15156,N_14727,N_14896);
or U15157 (N_15157,N_14581,N_14931);
nand U15158 (N_15158,N_14795,N_14870);
nor U15159 (N_15159,N_14809,N_14530);
nor U15160 (N_15160,N_14575,N_14818);
nand U15161 (N_15161,N_14963,N_14786);
and U15162 (N_15162,N_14869,N_14670);
nor U15163 (N_15163,N_14510,N_14994);
xor U15164 (N_15164,N_14854,N_14779);
and U15165 (N_15165,N_14752,N_14734);
xor U15166 (N_15166,N_14413,N_14791);
xor U15167 (N_15167,N_14719,N_14944);
xnor U15168 (N_15168,N_14664,N_14890);
and U15169 (N_15169,N_14947,N_14625);
xnor U15170 (N_15170,N_14756,N_14489);
and U15171 (N_15171,N_14832,N_14405);
nor U15172 (N_15172,N_14907,N_14626);
nand U15173 (N_15173,N_14899,N_14960);
xor U15174 (N_15174,N_14561,N_14741);
or U15175 (N_15175,N_14772,N_14673);
or U15176 (N_15176,N_14700,N_14825);
xor U15177 (N_15177,N_14528,N_14903);
xor U15178 (N_15178,N_14762,N_14407);
xor U15179 (N_15179,N_14820,N_14686);
nor U15180 (N_15180,N_14396,N_14503);
xnor U15181 (N_15181,N_14922,N_14650);
or U15182 (N_15182,N_14400,N_14492);
and U15183 (N_15183,N_14524,N_14782);
nor U15184 (N_15184,N_14705,N_14663);
and U15185 (N_15185,N_14570,N_14697);
nand U15186 (N_15186,N_14501,N_14445);
or U15187 (N_15187,N_14675,N_14526);
nor U15188 (N_15188,N_14647,N_14418);
nor U15189 (N_15189,N_14970,N_14381);
nand U15190 (N_15190,N_14512,N_14942);
nor U15191 (N_15191,N_14891,N_14937);
or U15192 (N_15192,N_14701,N_14799);
nor U15193 (N_15193,N_14696,N_14480);
xnor U15194 (N_15194,N_14808,N_14681);
or U15195 (N_15195,N_14576,N_14506);
nand U15196 (N_15196,N_14533,N_14868);
and U15197 (N_15197,N_14986,N_14787);
and U15198 (N_15198,N_14672,N_14662);
xnor U15199 (N_15199,N_14794,N_14776);
nor U15200 (N_15200,N_14880,N_14913);
nor U15201 (N_15201,N_14815,N_14687);
and U15202 (N_15202,N_14867,N_14995);
or U15203 (N_15203,N_14964,N_14393);
xnor U15204 (N_15204,N_14950,N_14991);
or U15205 (N_15205,N_14857,N_14646);
and U15206 (N_15206,N_14691,N_14684);
nor U15207 (N_15207,N_14642,N_14943);
nand U15208 (N_15208,N_14708,N_14580);
xor U15209 (N_15209,N_14925,N_14543);
or U15210 (N_15210,N_14416,N_14885);
or U15211 (N_15211,N_14534,N_14440);
and U15212 (N_15212,N_14933,N_14586);
and U15213 (N_15213,N_14454,N_14659);
nor U15214 (N_15214,N_14683,N_14853);
xnor U15215 (N_15215,N_14453,N_14775);
and U15216 (N_15216,N_14632,N_14619);
xor U15217 (N_15217,N_14550,N_14674);
nand U15218 (N_15218,N_14904,N_14666);
or U15219 (N_15219,N_14565,N_14814);
nor U15220 (N_15220,N_14469,N_14426);
nor U15221 (N_15221,N_14948,N_14478);
or U15222 (N_15222,N_14893,N_14468);
or U15223 (N_15223,N_14411,N_14608);
or U15224 (N_15224,N_14667,N_14497);
or U15225 (N_15225,N_14906,N_14547);
nor U15226 (N_15226,N_14644,N_14531);
nor U15227 (N_15227,N_14463,N_14997);
and U15228 (N_15228,N_14612,N_14998);
and U15229 (N_15229,N_14717,N_14386);
nand U15230 (N_15230,N_14611,N_14437);
xor U15231 (N_15231,N_14651,N_14410);
xor U15232 (N_15232,N_14971,N_14919);
xor U15233 (N_15233,N_14403,N_14564);
nor U15234 (N_15234,N_14598,N_14918);
and U15235 (N_15235,N_14709,N_14597);
nor U15236 (N_15236,N_14972,N_14855);
or U15237 (N_15237,N_14722,N_14486);
xor U15238 (N_15238,N_14658,N_14783);
nand U15239 (N_15239,N_14902,N_14976);
nor U15240 (N_15240,N_14452,N_14668);
xnor U15241 (N_15241,N_14888,N_14447);
xnor U15242 (N_15242,N_14923,N_14742);
and U15243 (N_15243,N_14620,N_14694);
nand U15244 (N_15244,N_14961,N_14912);
or U15245 (N_15245,N_14718,N_14716);
and U15246 (N_15246,N_14894,N_14967);
or U15247 (N_15247,N_14992,N_14583);
or U15248 (N_15248,N_14606,N_14882);
nor U15249 (N_15249,N_14711,N_14574);
nand U15250 (N_15250,N_14785,N_14712);
or U15251 (N_15251,N_14856,N_14836);
nand U15252 (N_15252,N_14605,N_14905);
nor U15253 (N_15253,N_14858,N_14499);
or U15254 (N_15254,N_14777,N_14641);
and U15255 (N_15255,N_14751,N_14467);
nand U15256 (N_15256,N_14946,N_14399);
nor U15257 (N_15257,N_14627,N_14511);
xnor U15258 (N_15258,N_14928,N_14767);
xor U15259 (N_15259,N_14379,N_14725);
and U15260 (N_15260,N_14385,N_14848);
and U15261 (N_15261,N_14706,N_14702);
nor U15262 (N_15262,N_14926,N_14661);
or U15263 (N_15263,N_14901,N_14648);
and U15264 (N_15264,N_14680,N_14911);
and U15265 (N_15265,N_14477,N_14415);
xor U15266 (N_15266,N_14724,N_14840);
and U15267 (N_15267,N_14536,N_14988);
nand U15268 (N_15268,N_14654,N_14449);
or U15269 (N_15269,N_14887,N_14929);
nor U15270 (N_15270,N_14397,N_14864);
nor U15271 (N_15271,N_14425,N_14498);
or U15272 (N_15272,N_14678,N_14593);
nor U15273 (N_15273,N_14748,N_14707);
or U15274 (N_15274,N_14474,N_14921);
xnor U15275 (N_15275,N_14539,N_14984);
nand U15276 (N_15276,N_14542,N_14757);
nand U15277 (N_15277,N_14487,N_14398);
nor U15278 (N_15278,N_14801,N_14969);
or U15279 (N_15279,N_14578,N_14951);
nand U15280 (N_15280,N_14450,N_14755);
or U15281 (N_15281,N_14438,N_14414);
xor U15282 (N_15282,N_14460,N_14852);
nand U15283 (N_15283,N_14989,N_14847);
xnor U15284 (N_15284,N_14479,N_14563);
xnor U15285 (N_15285,N_14796,N_14587);
xnor U15286 (N_15286,N_14483,N_14424);
or U15287 (N_15287,N_14688,N_14380);
nand U15288 (N_15288,N_14781,N_14979);
and U15289 (N_15289,N_14981,N_14941);
nor U15290 (N_15290,N_14914,N_14402);
nand U15291 (N_15291,N_14773,N_14968);
and U15292 (N_15292,N_14421,N_14760);
and U15293 (N_15293,N_14504,N_14679);
and U15294 (N_15294,N_14484,N_14392);
and U15295 (N_15295,N_14682,N_14710);
xor U15296 (N_15296,N_14876,N_14621);
nand U15297 (N_15297,N_14640,N_14470);
and U15298 (N_15298,N_14877,N_14618);
xor U15299 (N_15299,N_14657,N_14541);
or U15300 (N_15300,N_14544,N_14865);
nor U15301 (N_15301,N_14584,N_14821);
nand U15302 (N_15302,N_14616,N_14446);
and U15303 (N_15303,N_14874,N_14737);
xnor U15304 (N_15304,N_14838,N_14582);
or U15305 (N_15305,N_14695,N_14810);
and U15306 (N_15306,N_14502,N_14939);
nor U15307 (N_15307,N_14955,N_14889);
nand U15308 (N_15308,N_14835,N_14514);
or U15309 (N_15309,N_14793,N_14807);
and U15310 (N_15310,N_14500,N_14630);
and U15311 (N_15311,N_14568,N_14824);
and U15312 (N_15312,N_14878,N_14992);
and U15313 (N_15313,N_14451,N_14547);
or U15314 (N_15314,N_14604,N_14595);
nor U15315 (N_15315,N_14943,N_14634);
or U15316 (N_15316,N_14732,N_14473);
xor U15317 (N_15317,N_14504,N_14849);
and U15318 (N_15318,N_14888,N_14726);
or U15319 (N_15319,N_14487,N_14436);
nand U15320 (N_15320,N_14752,N_14679);
xnor U15321 (N_15321,N_14561,N_14375);
or U15322 (N_15322,N_14805,N_14460);
nor U15323 (N_15323,N_14949,N_14595);
xnor U15324 (N_15324,N_14591,N_14822);
nand U15325 (N_15325,N_14679,N_14465);
xnor U15326 (N_15326,N_14462,N_14546);
xor U15327 (N_15327,N_14808,N_14462);
and U15328 (N_15328,N_14690,N_14867);
or U15329 (N_15329,N_14445,N_14601);
nor U15330 (N_15330,N_14599,N_14466);
and U15331 (N_15331,N_14565,N_14651);
and U15332 (N_15332,N_14399,N_14477);
and U15333 (N_15333,N_14559,N_14890);
nand U15334 (N_15334,N_14952,N_14739);
or U15335 (N_15335,N_14424,N_14831);
and U15336 (N_15336,N_14382,N_14493);
and U15337 (N_15337,N_14521,N_14546);
nand U15338 (N_15338,N_14684,N_14444);
nand U15339 (N_15339,N_14501,N_14705);
and U15340 (N_15340,N_14746,N_14463);
nand U15341 (N_15341,N_14597,N_14383);
nand U15342 (N_15342,N_14789,N_14962);
and U15343 (N_15343,N_14724,N_14920);
or U15344 (N_15344,N_14605,N_14508);
xor U15345 (N_15345,N_14916,N_14575);
or U15346 (N_15346,N_14662,N_14821);
and U15347 (N_15347,N_14648,N_14424);
nand U15348 (N_15348,N_14821,N_14538);
xor U15349 (N_15349,N_14529,N_14716);
nor U15350 (N_15350,N_14529,N_14468);
nor U15351 (N_15351,N_14754,N_14474);
xnor U15352 (N_15352,N_14622,N_14474);
or U15353 (N_15353,N_14544,N_14803);
or U15354 (N_15354,N_14473,N_14460);
or U15355 (N_15355,N_14996,N_14912);
nand U15356 (N_15356,N_14837,N_14633);
nand U15357 (N_15357,N_14491,N_14570);
xnor U15358 (N_15358,N_14665,N_14808);
nand U15359 (N_15359,N_14699,N_14870);
and U15360 (N_15360,N_14837,N_14877);
nand U15361 (N_15361,N_14442,N_14452);
nor U15362 (N_15362,N_14489,N_14881);
and U15363 (N_15363,N_14380,N_14957);
and U15364 (N_15364,N_14851,N_14798);
and U15365 (N_15365,N_14503,N_14617);
and U15366 (N_15366,N_14687,N_14811);
xor U15367 (N_15367,N_14744,N_14946);
and U15368 (N_15368,N_14928,N_14568);
xnor U15369 (N_15369,N_14914,N_14567);
nand U15370 (N_15370,N_14400,N_14842);
xor U15371 (N_15371,N_14712,N_14849);
nand U15372 (N_15372,N_14451,N_14465);
and U15373 (N_15373,N_14982,N_14941);
or U15374 (N_15374,N_14569,N_14940);
nor U15375 (N_15375,N_14573,N_14492);
and U15376 (N_15376,N_14536,N_14946);
nor U15377 (N_15377,N_14656,N_14738);
and U15378 (N_15378,N_14699,N_14758);
or U15379 (N_15379,N_14418,N_14542);
nor U15380 (N_15380,N_14492,N_14412);
nor U15381 (N_15381,N_14666,N_14459);
nand U15382 (N_15382,N_14643,N_14451);
xor U15383 (N_15383,N_14743,N_14669);
nand U15384 (N_15384,N_14418,N_14968);
xor U15385 (N_15385,N_14528,N_14737);
xnor U15386 (N_15386,N_14607,N_14505);
nand U15387 (N_15387,N_14848,N_14448);
nor U15388 (N_15388,N_14497,N_14574);
and U15389 (N_15389,N_14552,N_14831);
and U15390 (N_15390,N_14500,N_14844);
or U15391 (N_15391,N_14784,N_14999);
xor U15392 (N_15392,N_14693,N_14448);
xor U15393 (N_15393,N_14650,N_14710);
xor U15394 (N_15394,N_14635,N_14737);
xnor U15395 (N_15395,N_14804,N_14578);
nand U15396 (N_15396,N_14726,N_14632);
xor U15397 (N_15397,N_14539,N_14497);
and U15398 (N_15398,N_14902,N_14547);
nand U15399 (N_15399,N_14842,N_14494);
nand U15400 (N_15400,N_14494,N_14956);
nor U15401 (N_15401,N_14619,N_14397);
and U15402 (N_15402,N_14623,N_14524);
nor U15403 (N_15403,N_14587,N_14436);
or U15404 (N_15404,N_14582,N_14647);
nor U15405 (N_15405,N_14984,N_14941);
nor U15406 (N_15406,N_14493,N_14603);
nor U15407 (N_15407,N_14590,N_14794);
nand U15408 (N_15408,N_14385,N_14995);
xnor U15409 (N_15409,N_14401,N_14670);
nand U15410 (N_15410,N_14583,N_14616);
xnor U15411 (N_15411,N_14802,N_14958);
xor U15412 (N_15412,N_14784,N_14494);
xor U15413 (N_15413,N_14949,N_14386);
or U15414 (N_15414,N_14699,N_14904);
xnor U15415 (N_15415,N_14525,N_14764);
nor U15416 (N_15416,N_14786,N_14571);
nand U15417 (N_15417,N_14522,N_14642);
or U15418 (N_15418,N_14887,N_14712);
nand U15419 (N_15419,N_14737,N_14658);
xnor U15420 (N_15420,N_14462,N_14784);
nand U15421 (N_15421,N_14676,N_14621);
and U15422 (N_15422,N_14384,N_14578);
xor U15423 (N_15423,N_14545,N_14954);
xnor U15424 (N_15424,N_14592,N_14568);
or U15425 (N_15425,N_14489,N_14510);
xor U15426 (N_15426,N_14638,N_14514);
nor U15427 (N_15427,N_14921,N_14893);
and U15428 (N_15428,N_14544,N_14936);
nand U15429 (N_15429,N_14913,N_14832);
xor U15430 (N_15430,N_14627,N_14663);
xor U15431 (N_15431,N_14890,N_14512);
nand U15432 (N_15432,N_14637,N_14871);
nor U15433 (N_15433,N_14669,N_14724);
nand U15434 (N_15434,N_14432,N_14859);
nor U15435 (N_15435,N_14778,N_14783);
xnor U15436 (N_15436,N_14926,N_14524);
nor U15437 (N_15437,N_14803,N_14892);
or U15438 (N_15438,N_14590,N_14733);
xnor U15439 (N_15439,N_14572,N_14931);
xor U15440 (N_15440,N_14835,N_14562);
nand U15441 (N_15441,N_14703,N_14622);
or U15442 (N_15442,N_14656,N_14384);
nor U15443 (N_15443,N_14836,N_14996);
xor U15444 (N_15444,N_14626,N_14418);
nand U15445 (N_15445,N_14514,N_14912);
nand U15446 (N_15446,N_14376,N_14578);
and U15447 (N_15447,N_14840,N_14837);
or U15448 (N_15448,N_14543,N_14772);
and U15449 (N_15449,N_14938,N_14481);
and U15450 (N_15450,N_14705,N_14589);
or U15451 (N_15451,N_14657,N_14655);
or U15452 (N_15452,N_14420,N_14822);
or U15453 (N_15453,N_14395,N_14379);
or U15454 (N_15454,N_14832,N_14840);
and U15455 (N_15455,N_14713,N_14398);
or U15456 (N_15456,N_14584,N_14430);
nor U15457 (N_15457,N_14903,N_14881);
or U15458 (N_15458,N_14565,N_14711);
nor U15459 (N_15459,N_14578,N_14998);
xnor U15460 (N_15460,N_14992,N_14648);
or U15461 (N_15461,N_14930,N_14726);
nand U15462 (N_15462,N_14967,N_14767);
xnor U15463 (N_15463,N_14716,N_14964);
xnor U15464 (N_15464,N_14608,N_14977);
nand U15465 (N_15465,N_14558,N_14537);
nor U15466 (N_15466,N_14672,N_14990);
nor U15467 (N_15467,N_14886,N_14974);
xnor U15468 (N_15468,N_14598,N_14428);
nor U15469 (N_15469,N_14491,N_14401);
and U15470 (N_15470,N_14479,N_14945);
or U15471 (N_15471,N_14491,N_14429);
xor U15472 (N_15472,N_14850,N_14965);
xor U15473 (N_15473,N_14975,N_14934);
and U15474 (N_15474,N_14997,N_14650);
xnor U15475 (N_15475,N_14946,N_14726);
nor U15476 (N_15476,N_14492,N_14649);
or U15477 (N_15477,N_14842,N_14810);
nor U15478 (N_15478,N_14748,N_14981);
xnor U15479 (N_15479,N_14383,N_14489);
nor U15480 (N_15480,N_14526,N_14991);
xnor U15481 (N_15481,N_14471,N_14894);
or U15482 (N_15482,N_14616,N_14947);
and U15483 (N_15483,N_14798,N_14726);
and U15484 (N_15484,N_14431,N_14408);
or U15485 (N_15485,N_14546,N_14960);
nand U15486 (N_15486,N_14385,N_14618);
nand U15487 (N_15487,N_14434,N_14509);
xor U15488 (N_15488,N_14861,N_14990);
nand U15489 (N_15489,N_14678,N_14505);
and U15490 (N_15490,N_14848,N_14866);
and U15491 (N_15491,N_14603,N_14907);
or U15492 (N_15492,N_14388,N_14562);
nand U15493 (N_15493,N_14731,N_14844);
nand U15494 (N_15494,N_14380,N_14819);
or U15495 (N_15495,N_14489,N_14676);
xor U15496 (N_15496,N_14395,N_14549);
nand U15497 (N_15497,N_14948,N_14682);
nor U15498 (N_15498,N_14656,N_14875);
nor U15499 (N_15499,N_14759,N_14662);
nand U15500 (N_15500,N_14853,N_14962);
nand U15501 (N_15501,N_14795,N_14583);
xor U15502 (N_15502,N_14849,N_14886);
and U15503 (N_15503,N_14410,N_14847);
nor U15504 (N_15504,N_14382,N_14904);
or U15505 (N_15505,N_14442,N_14706);
and U15506 (N_15506,N_14401,N_14488);
nand U15507 (N_15507,N_14884,N_14507);
or U15508 (N_15508,N_14896,N_14915);
xnor U15509 (N_15509,N_14909,N_14784);
or U15510 (N_15510,N_14973,N_14823);
or U15511 (N_15511,N_14654,N_14546);
xor U15512 (N_15512,N_14736,N_14935);
and U15513 (N_15513,N_14842,N_14682);
and U15514 (N_15514,N_14749,N_14813);
nor U15515 (N_15515,N_14574,N_14522);
nor U15516 (N_15516,N_14848,N_14489);
or U15517 (N_15517,N_14601,N_14843);
or U15518 (N_15518,N_14642,N_14394);
xor U15519 (N_15519,N_14518,N_14827);
xor U15520 (N_15520,N_14727,N_14908);
and U15521 (N_15521,N_14517,N_14657);
or U15522 (N_15522,N_14531,N_14646);
or U15523 (N_15523,N_14757,N_14759);
nor U15524 (N_15524,N_14458,N_14684);
xor U15525 (N_15525,N_14964,N_14758);
nor U15526 (N_15526,N_14514,N_14501);
or U15527 (N_15527,N_14449,N_14469);
nand U15528 (N_15528,N_14703,N_14440);
or U15529 (N_15529,N_14998,N_14746);
or U15530 (N_15530,N_14841,N_14477);
or U15531 (N_15531,N_14863,N_14611);
nor U15532 (N_15532,N_14517,N_14601);
and U15533 (N_15533,N_14991,N_14588);
xor U15534 (N_15534,N_14846,N_14679);
nand U15535 (N_15535,N_14430,N_14585);
and U15536 (N_15536,N_14553,N_14462);
and U15537 (N_15537,N_14401,N_14607);
and U15538 (N_15538,N_14776,N_14379);
nor U15539 (N_15539,N_14477,N_14710);
nor U15540 (N_15540,N_14920,N_14569);
and U15541 (N_15541,N_14703,N_14507);
xor U15542 (N_15542,N_14716,N_14651);
and U15543 (N_15543,N_14635,N_14741);
xnor U15544 (N_15544,N_14610,N_14930);
xor U15545 (N_15545,N_14973,N_14656);
nand U15546 (N_15546,N_14932,N_14996);
xor U15547 (N_15547,N_14879,N_14598);
and U15548 (N_15548,N_14805,N_14693);
nor U15549 (N_15549,N_14761,N_14957);
or U15550 (N_15550,N_14641,N_14870);
xnor U15551 (N_15551,N_14889,N_14424);
nor U15552 (N_15552,N_14422,N_14400);
and U15553 (N_15553,N_14634,N_14554);
or U15554 (N_15554,N_14926,N_14554);
and U15555 (N_15555,N_14755,N_14856);
or U15556 (N_15556,N_14759,N_14749);
nor U15557 (N_15557,N_14721,N_14620);
nor U15558 (N_15558,N_14781,N_14709);
or U15559 (N_15559,N_14804,N_14725);
or U15560 (N_15560,N_14893,N_14579);
nor U15561 (N_15561,N_14530,N_14715);
xor U15562 (N_15562,N_14565,N_14854);
or U15563 (N_15563,N_14793,N_14559);
xor U15564 (N_15564,N_14895,N_14881);
nand U15565 (N_15565,N_14815,N_14852);
nand U15566 (N_15566,N_14709,N_14656);
and U15567 (N_15567,N_14387,N_14894);
xnor U15568 (N_15568,N_14900,N_14724);
or U15569 (N_15569,N_14456,N_14761);
or U15570 (N_15570,N_14838,N_14477);
nand U15571 (N_15571,N_14413,N_14615);
and U15572 (N_15572,N_14881,N_14976);
nand U15573 (N_15573,N_14786,N_14707);
nor U15574 (N_15574,N_14445,N_14624);
or U15575 (N_15575,N_14889,N_14869);
xor U15576 (N_15576,N_14932,N_14526);
or U15577 (N_15577,N_14765,N_14394);
xnor U15578 (N_15578,N_14854,N_14457);
and U15579 (N_15579,N_14593,N_14798);
and U15580 (N_15580,N_14771,N_14775);
or U15581 (N_15581,N_14988,N_14562);
nand U15582 (N_15582,N_14537,N_14612);
nand U15583 (N_15583,N_14860,N_14381);
nand U15584 (N_15584,N_14616,N_14808);
or U15585 (N_15585,N_14694,N_14936);
or U15586 (N_15586,N_14548,N_14535);
nor U15587 (N_15587,N_14468,N_14655);
nor U15588 (N_15588,N_14378,N_14462);
nand U15589 (N_15589,N_14883,N_14639);
nand U15590 (N_15590,N_14411,N_14824);
or U15591 (N_15591,N_14489,N_14588);
nor U15592 (N_15592,N_14830,N_14760);
nand U15593 (N_15593,N_14706,N_14582);
and U15594 (N_15594,N_14545,N_14717);
nand U15595 (N_15595,N_14392,N_14748);
nor U15596 (N_15596,N_14954,N_14434);
nor U15597 (N_15597,N_14732,N_14731);
nor U15598 (N_15598,N_14908,N_14845);
xnor U15599 (N_15599,N_14693,N_14822);
nand U15600 (N_15600,N_14460,N_14959);
xnor U15601 (N_15601,N_14860,N_14385);
xor U15602 (N_15602,N_14558,N_14967);
nor U15603 (N_15603,N_14714,N_14640);
and U15604 (N_15604,N_14970,N_14481);
nor U15605 (N_15605,N_14730,N_14565);
nor U15606 (N_15606,N_14377,N_14597);
or U15607 (N_15607,N_14659,N_14633);
nand U15608 (N_15608,N_14447,N_14428);
xnor U15609 (N_15609,N_14519,N_14589);
nor U15610 (N_15610,N_14783,N_14429);
nor U15611 (N_15611,N_14436,N_14751);
nor U15612 (N_15612,N_14519,N_14693);
or U15613 (N_15613,N_14536,N_14947);
or U15614 (N_15614,N_14426,N_14526);
nor U15615 (N_15615,N_14617,N_14907);
or U15616 (N_15616,N_14450,N_14566);
nand U15617 (N_15617,N_14650,N_14807);
nor U15618 (N_15618,N_14543,N_14688);
nand U15619 (N_15619,N_14571,N_14980);
xor U15620 (N_15620,N_14928,N_14934);
xnor U15621 (N_15621,N_14879,N_14560);
xor U15622 (N_15622,N_14637,N_14801);
nand U15623 (N_15623,N_14832,N_14629);
or U15624 (N_15624,N_14451,N_14539);
xnor U15625 (N_15625,N_15461,N_15302);
nand U15626 (N_15626,N_15435,N_15209);
xnor U15627 (N_15627,N_15072,N_15450);
nor U15628 (N_15628,N_15032,N_15205);
nand U15629 (N_15629,N_15382,N_15419);
and U15630 (N_15630,N_15469,N_15191);
nor U15631 (N_15631,N_15414,N_15124);
or U15632 (N_15632,N_15423,N_15617);
xnor U15633 (N_15633,N_15091,N_15011);
nor U15634 (N_15634,N_15605,N_15543);
or U15635 (N_15635,N_15394,N_15041);
or U15636 (N_15636,N_15086,N_15075);
nand U15637 (N_15637,N_15022,N_15261);
xnor U15638 (N_15638,N_15189,N_15196);
nor U15639 (N_15639,N_15295,N_15030);
nor U15640 (N_15640,N_15380,N_15216);
nand U15641 (N_15641,N_15060,N_15584);
nor U15642 (N_15642,N_15095,N_15051);
and U15643 (N_15643,N_15146,N_15157);
nor U15644 (N_15644,N_15102,N_15468);
nand U15645 (N_15645,N_15046,N_15168);
and U15646 (N_15646,N_15043,N_15519);
and U15647 (N_15647,N_15203,N_15577);
xnor U15648 (N_15648,N_15156,N_15613);
or U15649 (N_15649,N_15400,N_15561);
xnor U15650 (N_15650,N_15565,N_15090);
nand U15651 (N_15651,N_15056,N_15366);
nand U15652 (N_15652,N_15129,N_15153);
nand U15653 (N_15653,N_15180,N_15276);
and U15654 (N_15654,N_15106,N_15337);
nand U15655 (N_15655,N_15356,N_15340);
and U15656 (N_15656,N_15431,N_15225);
nand U15657 (N_15657,N_15358,N_15334);
and U15658 (N_15658,N_15262,N_15004);
or U15659 (N_15659,N_15281,N_15158);
or U15660 (N_15660,N_15396,N_15512);
nor U15661 (N_15661,N_15019,N_15258);
nor U15662 (N_15662,N_15315,N_15260);
and U15663 (N_15663,N_15199,N_15525);
or U15664 (N_15664,N_15407,N_15593);
xnor U15665 (N_15665,N_15575,N_15355);
nand U15666 (N_15666,N_15006,N_15047);
and U15667 (N_15667,N_15485,N_15580);
nor U15668 (N_15668,N_15226,N_15067);
or U15669 (N_15669,N_15208,N_15193);
nand U15670 (N_15670,N_15327,N_15574);
xnor U15671 (N_15671,N_15369,N_15614);
xor U15672 (N_15672,N_15397,N_15351);
and U15673 (N_15673,N_15294,N_15456);
xnor U15674 (N_15674,N_15064,N_15161);
or U15675 (N_15675,N_15291,N_15378);
xnor U15676 (N_15676,N_15424,N_15109);
and U15677 (N_15677,N_15212,N_15445);
or U15678 (N_15678,N_15094,N_15235);
or U15679 (N_15679,N_15472,N_15087);
or U15680 (N_15680,N_15350,N_15105);
nor U15681 (N_15681,N_15421,N_15089);
nor U15682 (N_15682,N_15594,N_15304);
nand U15683 (N_15683,N_15365,N_15021);
nor U15684 (N_15684,N_15268,N_15517);
or U15685 (N_15685,N_15562,N_15504);
or U15686 (N_15686,N_15425,N_15462);
xor U15687 (N_15687,N_15240,N_15441);
nor U15688 (N_15688,N_15053,N_15368);
and U15689 (N_15689,N_15403,N_15275);
nor U15690 (N_15690,N_15583,N_15038);
nand U15691 (N_15691,N_15499,N_15406);
xor U15692 (N_15692,N_15353,N_15218);
and U15693 (N_15693,N_15540,N_15621);
nand U15694 (N_15694,N_15376,N_15470);
nand U15695 (N_15695,N_15137,N_15055);
or U15696 (N_15696,N_15411,N_15428);
nor U15697 (N_15697,N_15464,N_15392);
nor U15698 (N_15698,N_15172,N_15384);
nand U15699 (N_15699,N_15217,N_15017);
nor U15700 (N_15700,N_15541,N_15573);
or U15701 (N_15701,N_15306,N_15563);
nand U15702 (N_15702,N_15618,N_15555);
xnor U15703 (N_15703,N_15232,N_15404);
nand U15704 (N_15704,N_15220,N_15524);
and U15705 (N_15705,N_15219,N_15181);
nand U15706 (N_15706,N_15438,N_15164);
and U15707 (N_15707,N_15532,N_15527);
nand U15708 (N_15708,N_15549,N_15202);
and U15709 (N_15709,N_15045,N_15479);
and U15710 (N_15710,N_15393,N_15115);
xor U15711 (N_15711,N_15388,N_15552);
or U15712 (N_15712,N_15607,N_15098);
or U15713 (N_15713,N_15417,N_15033);
or U15714 (N_15714,N_15077,N_15223);
or U15715 (N_15715,N_15127,N_15572);
or U15716 (N_15716,N_15163,N_15429);
or U15717 (N_15717,N_15483,N_15335);
xnor U15718 (N_15718,N_15005,N_15332);
nand U15719 (N_15719,N_15453,N_15538);
nand U15720 (N_15720,N_15277,N_15426);
nor U15721 (N_15721,N_15269,N_15523);
or U15722 (N_15722,N_15195,N_15273);
or U15723 (N_15723,N_15535,N_15321);
or U15724 (N_15724,N_15314,N_15536);
nor U15725 (N_15725,N_15210,N_15062);
and U15726 (N_15726,N_15059,N_15263);
xnor U15727 (N_15727,N_15252,N_15074);
or U15728 (N_15728,N_15034,N_15344);
or U15729 (N_15729,N_15436,N_15080);
or U15730 (N_15730,N_15215,N_15514);
nand U15731 (N_15731,N_15134,N_15183);
nor U15732 (N_15732,N_15513,N_15178);
and U15733 (N_15733,N_15117,N_15248);
nand U15734 (N_15734,N_15526,N_15118);
or U15735 (N_15735,N_15012,N_15026);
and U15736 (N_15736,N_15130,N_15330);
or U15737 (N_15737,N_15606,N_15615);
xor U15738 (N_15738,N_15507,N_15323);
xor U15739 (N_15739,N_15307,N_15290);
nor U15740 (N_15740,N_15467,N_15151);
nor U15741 (N_15741,N_15126,N_15534);
nor U15742 (N_15742,N_15147,N_15624);
and U15743 (N_15743,N_15374,N_15265);
nor U15744 (N_15744,N_15296,N_15498);
and U15745 (N_15745,N_15297,N_15081);
nor U15746 (N_15746,N_15434,N_15533);
or U15747 (N_15747,N_15042,N_15206);
nand U15748 (N_15748,N_15010,N_15511);
nand U15749 (N_15749,N_15135,N_15009);
and U15750 (N_15750,N_15066,N_15385);
nand U15751 (N_15751,N_15610,N_15031);
nand U15752 (N_15752,N_15389,N_15515);
nor U15753 (N_15753,N_15559,N_15283);
and U15754 (N_15754,N_15308,N_15558);
nand U15755 (N_15755,N_15581,N_15027);
nor U15756 (N_15756,N_15174,N_15286);
xor U15757 (N_15757,N_15395,N_15326);
nand U15758 (N_15758,N_15182,N_15491);
and U15759 (N_15759,N_15586,N_15416);
nand U15760 (N_15760,N_15474,N_15224);
xnor U15761 (N_15761,N_15143,N_15221);
or U15762 (N_15762,N_15415,N_15054);
xor U15763 (N_15763,N_15370,N_15233);
and U15764 (N_15764,N_15255,N_15247);
or U15765 (N_15765,N_15363,N_15449);
nand U15766 (N_15766,N_15267,N_15239);
nand U15767 (N_15767,N_15371,N_15279);
xor U15768 (N_15768,N_15188,N_15387);
nand U15769 (N_15769,N_15443,N_15272);
and U15770 (N_15770,N_15390,N_15271);
nor U15771 (N_15771,N_15357,N_15024);
and U15772 (N_15772,N_15481,N_15037);
nor U15773 (N_15773,N_15016,N_15300);
nor U15774 (N_15774,N_15322,N_15061);
nor U15775 (N_15775,N_15142,N_15342);
nand U15776 (N_15776,N_15123,N_15293);
xnor U15777 (N_15777,N_15333,N_15571);
nor U15778 (N_15778,N_15166,N_15346);
nor U15779 (N_15779,N_15444,N_15508);
nand U15780 (N_15780,N_15254,N_15301);
xnor U15781 (N_15781,N_15207,N_15539);
or U15782 (N_15782,N_15408,N_15070);
and U15783 (N_15783,N_15317,N_15493);
nor U15784 (N_15784,N_15537,N_15497);
nand U15785 (N_15785,N_15299,N_15375);
and U15786 (N_15786,N_15201,N_15112);
xnor U15787 (N_15787,N_15484,N_15015);
or U15788 (N_15788,N_15457,N_15522);
nand U15789 (N_15789,N_15150,N_15092);
xor U15790 (N_15790,N_15554,N_15116);
or U15791 (N_15791,N_15413,N_15338);
or U15792 (N_15792,N_15602,N_15556);
or U15793 (N_15793,N_15285,N_15520);
nand U15794 (N_15794,N_15324,N_15176);
or U15795 (N_15795,N_15623,N_15597);
nor U15796 (N_15796,N_15229,N_15347);
xnor U15797 (N_15797,N_15132,N_15341);
xor U15798 (N_15798,N_15110,N_15590);
and U15799 (N_15799,N_15253,N_15148);
and U15800 (N_15800,N_15360,N_15402);
nor U15801 (N_15801,N_15320,N_15083);
nor U15802 (N_15802,N_15547,N_15364);
or U15803 (N_15803,N_15065,N_15236);
or U15804 (N_15804,N_15282,N_15138);
and U15805 (N_15805,N_15014,N_15251);
xor U15806 (N_15806,N_15104,N_15084);
nor U15807 (N_15807,N_15050,N_15437);
or U15808 (N_15808,N_15131,N_15412);
xnor U15809 (N_15809,N_15528,N_15440);
or U15810 (N_15810,N_15155,N_15319);
nand U15811 (N_15811,N_15316,N_15570);
and U15812 (N_15812,N_15608,N_15345);
or U15813 (N_15813,N_15177,N_15000);
or U15814 (N_15814,N_15093,N_15447);
and U15815 (N_15815,N_15367,N_15505);
nand U15816 (N_15816,N_15198,N_15008);
nand U15817 (N_15817,N_15100,N_15501);
nand U15818 (N_15818,N_15487,N_15194);
nor U15819 (N_15819,N_15566,N_15305);
and U15820 (N_15820,N_15274,N_15465);
xnor U15821 (N_15821,N_15001,N_15557);
nand U15822 (N_15822,N_15298,N_15489);
nand U15823 (N_15823,N_15318,N_15544);
nor U15824 (N_15824,N_15303,N_15230);
xnor U15825 (N_15825,N_15490,N_15482);
or U15826 (N_15826,N_15410,N_15187);
nor U15827 (N_15827,N_15107,N_15471);
and U15828 (N_15828,N_15496,N_15492);
nor U15829 (N_15829,N_15159,N_15057);
nor U15830 (N_15830,N_15312,N_15145);
nor U15831 (N_15831,N_15068,N_15582);
or U15832 (N_15832,N_15007,N_15500);
nand U15833 (N_15833,N_15354,N_15292);
nand U15834 (N_15834,N_15530,N_15099);
nor U15835 (N_15835,N_15204,N_15509);
and U15836 (N_15836,N_15518,N_15136);
nor U15837 (N_15837,N_15567,N_15133);
or U15838 (N_15838,N_15200,N_15144);
xnor U15839 (N_15839,N_15585,N_15542);
or U15840 (N_15840,N_15620,N_15044);
and U15841 (N_15841,N_15288,N_15329);
or U15842 (N_15842,N_15211,N_15601);
nand U15843 (N_15843,N_15560,N_15173);
nand U15844 (N_15844,N_15222,N_15197);
nor U15845 (N_15845,N_15439,N_15348);
xor U15846 (N_15846,N_15488,N_15241);
nor U15847 (N_15847,N_15113,N_15451);
nor U15848 (N_15848,N_15186,N_15448);
or U15849 (N_15849,N_15418,N_15069);
nor U15850 (N_15850,N_15103,N_15569);
and U15851 (N_15851,N_15386,N_15079);
nor U15852 (N_15852,N_15058,N_15463);
or U15853 (N_15853,N_15114,N_15568);
or U15854 (N_15854,N_15289,N_15078);
or U15855 (N_15855,N_15171,N_15170);
xor U15856 (N_15856,N_15578,N_15071);
or U15857 (N_15857,N_15139,N_15551);
nor U15858 (N_15858,N_15063,N_15002);
or U15859 (N_15859,N_15264,N_15029);
nor U15860 (N_15860,N_15190,N_15433);
or U15861 (N_15861,N_15082,N_15475);
or U15862 (N_15862,N_15160,N_15452);
xnor U15863 (N_15863,N_15266,N_15603);
xor U15864 (N_15864,N_15125,N_15227);
and U15865 (N_15865,N_15502,N_15284);
or U15866 (N_15866,N_15506,N_15154);
and U15867 (N_15867,N_15458,N_15018);
nor U15868 (N_15868,N_15588,N_15278);
or U15869 (N_15869,N_15473,N_15234);
nor U15870 (N_15870,N_15336,N_15013);
and U15871 (N_15871,N_15250,N_15399);
nand U15872 (N_15872,N_15422,N_15516);
nand U15873 (N_15873,N_15003,N_15256);
nor U15874 (N_15874,N_15373,N_15430);
nor U15875 (N_15875,N_15121,N_15361);
nand U15876 (N_15876,N_15432,N_15579);
nand U15877 (N_15877,N_15427,N_15480);
and U15878 (N_15878,N_15459,N_15245);
nand U15879 (N_15879,N_15587,N_15108);
xnor U15880 (N_15880,N_15119,N_15313);
xnor U15881 (N_15881,N_15372,N_15466);
xnor U15882 (N_15882,N_15494,N_15052);
xor U15883 (N_15883,N_15442,N_15049);
nand U15884 (N_15884,N_15162,N_15548);
and U15885 (N_15885,N_15595,N_15244);
xor U15886 (N_15886,N_15339,N_15179);
and U15887 (N_15887,N_15619,N_15242);
xnor U15888 (N_15888,N_15383,N_15401);
or U15889 (N_15889,N_15343,N_15510);
or U15890 (N_15890,N_15228,N_15391);
and U15891 (N_15891,N_15405,N_15454);
nor U15892 (N_15892,N_15149,N_15152);
and U15893 (N_15893,N_15280,N_15531);
xor U15894 (N_15894,N_15096,N_15611);
xor U15895 (N_15895,N_15328,N_15455);
or U15896 (N_15896,N_15352,N_15231);
or U15897 (N_15897,N_15048,N_15550);
xnor U15898 (N_15898,N_15599,N_15249);
xnor U15899 (N_15899,N_15545,N_15460);
nand U15900 (N_15900,N_15076,N_15025);
nand U15901 (N_15901,N_15287,N_15169);
nor U15902 (N_15902,N_15165,N_15379);
or U15903 (N_15903,N_15246,N_15311);
or U15904 (N_15904,N_15213,N_15546);
xor U15905 (N_15905,N_15167,N_15612);
and U15906 (N_15906,N_15622,N_15257);
or U15907 (N_15907,N_15141,N_15035);
nor U15908 (N_15908,N_15270,N_15598);
nand U15909 (N_15909,N_15097,N_15023);
nand U15910 (N_15910,N_15349,N_15592);
nand U15911 (N_15911,N_15085,N_15503);
nand U15912 (N_15912,N_15243,N_15039);
nand U15913 (N_15913,N_15521,N_15073);
nor U15914 (N_15914,N_15185,N_15028);
xor U15915 (N_15915,N_15604,N_15192);
nand U15916 (N_15916,N_15600,N_15564);
and U15917 (N_15917,N_15128,N_15120);
nor U15918 (N_15918,N_15101,N_15184);
and U15919 (N_15919,N_15576,N_15175);
xnor U15920 (N_15920,N_15331,N_15214);
and U15921 (N_15921,N_15529,N_15477);
xnor U15922 (N_15922,N_15362,N_15237);
or U15923 (N_15923,N_15420,N_15020);
nand U15924 (N_15924,N_15596,N_15553);
xor U15925 (N_15925,N_15111,N_15040);
xor U15926 (N_15926,N_15140,N_15359);
nor U15927 (N_15927,N_15476,N_15377);
and U15928 (N_15928,N_15591,N_15609);
xnor U15929 (N_15929,N_15495,N_15589);
xnor U15930 (N_15930,N_15122,N_15446);
or U15931 (N_15931,N_15309,N_15238);
xnor U15932 (N_15932,N_15325,N_15409);
or U15933 (N_15933,N_15398,N_15310);
or U15934 (N_15934,N_15088,N_15478);
xor U15935 (N_15935,N_15036,N_15381);
nand U15936 (N_15936,N_15616,N_15486);
xor U15937 (N_15937,N_15259,N_15272);
and U15938 (N_15938,N_15580,N_15278);
nand U15939 (N_15939,N_15363,N_15353);
nand U15940 (N_15940,N_15417,N_15084);
and U15941 (N_15941,N_15087,N_15431);
xnor U15942 (N_15942,N_15079,N_15620);
xor U15943 (N_15943,N_15324,N_15415);
nor U15944 (N_15944,N_15147,N_15260);
and U15945 (N_15945,N_15000,N_15574);
nand U15946 (N_15946,N_15261,N_15575);
nand U15947 (N_15947,N_15434,N_15249);
or U15948 (N_15948,N_15482,N_15212);
or U15949 (N_15949,N_15264,N_15034);
nand U15950 (N_15950,N_15184,N_15197);
nand U15951 (N_15951,N_15260,N_15279);
nand U15952 (N_15952,N_15274,N_15600);
nand U15953 (N_15953,N_15132,N_15286);
nand U15954 (N_15954,N_15369,N_15225);
xor U15955 (N_15955,N_15451,N_15472);
nand U15956 (N_15956,N_15159,N_15084);
and U15957 (N_15957,N_15185,N_15202);
or U15958 (N_15958,N_15125,N_15087);
nand U15959 (N_15959,N_15255,N_15389);
and U15960 (N_15960,N_15045,N_15225);
nand U15961 (N_15961,N_15042,N_15073);
nor U15962 (N_15962,N_15224,N_15131);
nand U15963 (N_15963,N_15532,N_15175);
nand U15964 (N_15964,N_15197,N_15145);
or U15965 (N_15965,N_15278,N_15357);
or U15966 (N_15966,N_15209,N_15164);
or U15967 (N_15967,N_15249,N_15590);
nand U15968 (N_15968,N_15389,N_15250);
or U15969 (N_15969,N_15410,N_15132);
nor U15970 (N_15970,N_15351,N_15307);
or U15971 (N_15971,N_15319,N_15254);
and U15972 (N_15972,N_15564,N_15451);
and U15973 (N_15973,N_15425,N_15351);
xnor U15974 (N_15974,N_15267,N_15342);
and U15975 (N_15975,N_15241,N_15283);
or U15976 (N_15976,N_15555,N_15121);
nor U15977 (N_15977,N_15127,N_15485);
xnor U15978 (N_15978,N_15578,N_15407);
nor U15979 (N_15979,N_15581,N_15106);
xnor U15980 (N_15980,N_15568,N_15169);
or U15981 (N_15981,N_15097,N_15426);
nor U15982 (N_15982,N_15265,N_15450);
or U15983 (N_15983,N_15044,N_15356);
nor U15984 (N_15984,N_15514,N_15609);
or U15985 (N_15985,N_15257,N_15051);
nand U15986 (N_15986,N_15451,N_15281);
or U15987 (N_15987,N_15156,N_15426);
xor U15988 (N_15988,N_15294,N_15019);
xnor U15989 (N_15989,N_15435,N_15065);
and U15990 (N_15990,N_15176,N_15025);
nand U15991 (N_15991,N_15070,N_15025);
xor U15992 (N_15992,N_15139,N_15425);
xnor U15993 (N_15993,N_15457,N_15337);
xor U15994 (N_15994,N_15441,N_15339);
or U15995 (N_15995,N_15209,N_15564);
or U15996 (N_15996,N_15355,N_15079);
xnor U15997 (N_15997,N_15247,N_15149);
nand U15998 (N_15998,N_15573,N_15129);
nand U15999 (N_15999,N_15038,N_15449);
and U16000 (N_16000,N_15068,N_15379);
nand U16001 (N_16001,N_15064,N_15039);
nand U16002 (N_16002,N_15032,N_15457);
nor U16003 (N_16003,N_15056,N_15355);
xor U16004 (N_16004,N_15166,N_15373);
and U16005 (N_16005,N_15504,N_15436);
nor U16006 (N_16006,N_15414,N_15422);
or U16007 (N_16007,N_15474,N_15596);
and U16008 (N_16008,N_15172,N_15326);
nor U16009 (N_16009,N_15343,N_15135);
nand U16010 (N_16010,N_15263,N_15490);
nand U16011 (N_16011,N_15338,N_15084);
nand U16012 (N_16012,N_15477,N_15027);
or U16013 (N_16013,N_15323,N_15041);
or U16014 (N_16014,N_15186,N_15144);
xor U16015 (N_16015,N_15216,N_15557);
xnor U16016 (N_16016,N_15002,N_15515);
nand U16017 (N_16017,N_15526,N_15067);
xnor U16018 (N_16018,N_15305,N_15265);
xor U16019 (N_16019,N_15585,N_15136);
and U16020 (N_16020,N_15446,N_15284);
nor U16021 (N_16021,N_15144,N_15606);
nand U16022 (N_16022,N_15423,N_15058);
nand U16023 (N_16023,N_15238,N_15386);
nand U16024 (N_16024,N_15053,N_15231);
or U16025 (N_16025,N_15361,N_15574);
nor U16026 (N_16026,N_15141,N_15191);
nor U16027 (N_16027,N_15544,N_15568);
or U16028 (N_16028,N_15228,N_15591);
and U16029 (N_16029,N_15194,N_15482);
and U16030 (N_16030,N_15303,N_15556);
or U16031 (N_16031,N_15168,N_15237);
xor U16032 (N_16032,N_15062,N_15253);
and U16033 (N_16033,N_15607,N_15599);
nor U16034 (N_16034,N_15314,N_15123);
and U16035 (N_16035,N_15575,N_15123);
nand U16036 (N_16036,N_15037,N_15421);
or U16037 (N_16037,N_15320,N_15512);
nand U16038 (N_16038,N_15301,N_15572);
and U16039 (N_16039,N_15467,N_15038);
nand U16040 (N_16040,N_15079,N_15613);
nand U16041 (N_16041,N_15269,N_15422);
or U16042 (N_16042,N_15155,N_15250);
or U16043 (N_16043,N_15502,N_15445);
or U16044 (N_16044,N_15029,N_15357);
xor U16045 (N_16045,N_15358,N_15174);
and U16046 (N_16046,N_15430,N_15068);
or U16047 (N_16047,N_15022,N_15453);
xnor U16048 (N_16048,N_15503,N_15173);
and U16049 (N_16049,N_15322,N_15057);
xor U16050 (N_16050,N_15560,N_15189);
or U16051 (N_16051,N_15279,N_15598);
nand U16052 (N_16052,N_15135,N_15569);
xor U16053 (N_16053,N_15477,N_15043);
nor U16054 (N_16054,N_15019,N_15318);
and U16055 (N_16055,N_15514,N_15401);
nor U16056 (N_16056,N_15039,N_15524);
nor U16057 (N_16057,N_15069,N_15586);
and U16058 (N_16058,N_15294,N_15193);
and U16059 (N_16059,N_15574,N_15463);
nor U16060 (N_16060,N_15494,N_15019);
and U16061 (N_16061,N_15482,N_15540);
and U16062 (N_16062,N_15291,N_15450);
xnor U16063 (N_16063,N_15315,N_15209);
or U16064 (N_16064,N_15230,N_15605);
or U16065 (N_16065,N_15290,N_15598);
and U16066 (N_16066,N_15336,N_15314);
xnor U16067 (N_16067,N_15372,N_15165);
nand U16068 (N_16068,N_15190,N_15232);
and U16069 (N_16069,N_15385,N_15045);
xnor U16070 (N_16070,N_15610,N_15374);
or U16071 (N_16071,N_15008,N_15285);
and U16072 (N_16072,N_15386,N_15545);
or U16073 (N_16073,N_15622,N_15480);
or U16074 (N_16074,N_15244,N_15067);
nand U16075 (N_16075,N_15353,N_15315);
nand U16076 (N_16076,N_15369,N_15498);
nor U16077 (N_16077,N_15064,N_15280);
nor U16078 (N_16078,N_15358,N_15262);
nand U16079 (N_16079,N_15474,N_15077);
xor U16080 (N_16080,N_15259,N_15478);
xor U16081 (N_16081,N_15414,N_15349);
nand U16082 (N_16082,N_15205,N_15604);
xnor U16083 (N_16083,N_15531,N_15077);
nor U16084 (N_16084,N_15506,N_15289);
nor U16085 (N_16085,N_15488,N_15034);
nor U16086 (N_16086,N_15281,N_15396);
nand U16087 (N_16087,N_15050,N_15327);
nor U16088 (N_16088,N_15446,N_15491);
xor U16089 (N_16089,N_15476,N_15175);
and U16090 (N_16090,N_15348,N_15349);
xnor U16091 (N_16091,N_15354,N_15477);
nand U16092 (N_16092,N_15221,N_15017);
xor U16093 (N_16093,N_15461,N_15297);
nand U16094 (N_16094,N_15272,N_15419);
nor U16095 (N_16095,N_15179,N_15601);
nand U16096 (N_16096,N_15321,N_15168);
nand U16097 (N_16097,N_15327,N_15082);
and U16098 (N_16098,N_15624,N_15393);
or U16099 (N_16099,N_15280,N_15302);
xor U16100 (N_16100,N_15523,N_15270);
or U16101 (N_16101,N_15057,N_15301);
or U16102 (N_16102,N_15423,N_15583);
nand U16103 (N_16103,N_15257,N_15176);
and U16104 (N_16104,N_15022,N_15343);
xor U16105 (N_16105,N_15508,N_15369);
or U16106 (N_16106,N_15313,N_15065);
nor U16107 (N_16107,N_15008,N_15225);
and U16108 (N_16108,N_15165,N_15128);
and U16109 (N_16109,N_15237,N_15543);
nand U16110 (N_16110,N_15569,N_15287);
or U16111 (N_16111,N_15338,N_15244);
nor U16112 (N_16112,N_15240,N_15513);
nor U16113 (N_16113,N_15183,N_15261);
xor U16114 (N_16114,N_15587,N_15010);
nor U16115 (N_16115,N_15606,N_15088);
nand U16116 (N_16116,N_15533,N_15512);
and U16117 (N_16117,N_15297,N_15310);
nor U16118 (N_16118,N_15081,N_15057);
xnor U16119 (N_16119,N_15100,N_15267);
and U16120 (N_16120,N_15423,N_15381);
and U16121 (N_16121,N_15267,N_15205);
xnor U16122 (N_16122,N_15414,N_15536);
or U16123 (N_16123,N_15583,N_15340);
xor U16124 (N_16124,N_15343,N_15511);
xor U16125 (N_16125,N_15249,N_15205);
nand U16126 (N_16126,N_15255,N_15095);
and U16127 (N_16127,N_15423,N_15138);
nand U16128 (N_16128,N_15242,N_15363);
and U16129 (N_16129,N_15173,N_15046);
or U16130 (N_16130,N_15275,N_15587);
nand U16131 (N_16131,N_15557,N_15552);
and U16132 (N_16132,N_15416,N_15384);
nand U16133 (N_16133,N_15158,N_15252);
xor U16134 (N_16134,N_15217,N_15104);
nand U16135 (N_16135,N_15523,N_15493);
or U16136 (N_16136,N_15425,N_15450);
and U16137 (N_16137,N_15326,N_15232);
nand U16138 (N_16138,N_15143,N_15613);
nor U16139 (N_16139,N_15318,N_15054);
nand U16140 (N_16140,N_15132,N_15258);
and U16141 (N_16141,N_15405,N_15047);
xnor U16142 (N_16142,N_15340,N_15487);
and U16143 (N_16143,N_15493,N_15122);
nand U16144 (N_16144,N_15277,N_15114);
or U16145 (N_16145,N_15215,N_15241);
xnor U16146 (N_16146,N_15493,N_15073);
nor U16147 (N_16147,N_15439,N_15156);
and U16148 (N_16148,N_15332,N_15125);
or U16149 (N_16149,N_15129,N_15408);
or U16150 (N_16150,N_15164,N_15074);
nor U16151 (N_16151,N_15246,N_15124);
nor U16152 (N_16152,N_15158,N_15058);
nor U16153 (N_16153,N_15187,N_15440);
xor U16154 (N_16154,N_15113,N_15442);
nor U16155 (N_16155,N_15136,N_15520);
and U16156 (N_16156,N_15515,N_15290);
xnor U16157 (N_16157,N_15509,N_15151);
or U16158 (N_16158,N_15356,N_15387);
nor U16159 (N_16159,N_15300,N_15293);
or U16160 (N_16160,N_15061,N_15020);
nand U16161 (N_16161,N_15019,N_15209);
xor U16162 (N_16162,N_15016,N_15490);
and U16163 (N_16163,N_15333,N_15440);
and U16164 (N_16164,N_15572,N_15186);
or U16165 (N_16165,N_15008,N_15372);
nor U16166 (N_16166,N_15620,N_15331);
and U16167 (N_16167,N_15575,N_15369);
and U16168 (N_16168,N_15461,N_15360);
and U16169 (N_16169,N_15447,N_15116);
or U16170 (N_16170,N_15108,N_15377);
nor U16171 (N_16171,N_15043,N_15530);
nor U16172 (N_16172,N_15519,N_15114);
nand U16173 (N_16173,N_15073,N_15263);
or U16174 (N_16174,N_15426,N_15354);
and U16175 (N_16175,N_15579,N_15490);
xnor U16176 (N_16176,N_15496,N_15264);
nor U16177 (N_16177,N_15505,N_15617);
and U16178 (N_16178,N_15551,N_15606);
nand U16179 (N_16179,N_15415,N_15240);
nor U16180 (N_16180,N_15617,N_15482);
and U16181 (N_16181,N_15578,N_15070);
or U16182 (N_16182,N_15211,N_15460);
nor U16183 (N_16183,N_15545,N_15397);
nor U16184 (N_16184,N_15267,N_15111);
or U16185 (N_16185,N_15405,N_15509);
or U16186 (N_16186,N_15216,N_15346);
or U16187 (N_16187,N_15093,N_15551);
xor U16188 (N_16188,N_15319,N_15343);
nor U16189 (N_16189,N_15386,N_15090);
and U16190 (N_16190,N_15481,N_15020);
xor U16191 (N_16191,N_15576,N_15241);
or U16192 (N_16192,N_15106,N_15332);
or U16193 (N_16193,N_15032,N_15065);
and U16194 (N_16194,N_15484,N_15621);
and U16195 (N_16195,N_15225,N_15433);
xor U16196 (N_16196,N_15510,N_15048);
or U16197 (N_16197,N_15403,N_15441);
and U16198 (N_16198,N_15596,N_15340);
nand U16199 (N_16199,N_15246,N_15025);
or U16200 (N_16200,N_15107,N_15621);
nor U16201 (N_16201,N_15384,N_15613);
and U16202 (N_16202,N_15505,N_15562);
or U16203 (N_16203,N_15337,N_15208);
or U16204 (N_16204,N_15326,N_15555);
nor U16205 (N_16205,N_15106,N_15482);
xnor U16206 (N_16206,N_15519,N_15289);
or U16207 (N_16207,N_15567,N_15471);
nand U16208 (N_16208,N_15485,N_15251);
nand U16209 (N_16209,N_15570,N_15114);
nor U16210 (N_16210,N_15004,N_15027);
or U16211 (N_16211,N_15372,N_15418);
or U16212 (N_16212,N_15023,N_15258);
or U16213 (N_16213,N_15287,N_15556);
nand U16214 (N_16214,N_15449,N_15134);
and U16215 (N_16215,N_15422,N_15328);
or U16216 (N_16216,N_15061,N_15277);
nor U16217 (N_16217,N_15394,N_15336);
xnor U16218 (N_16218,N_15033,N_15613);
or U16219 (N_16219,N_15573,N_15315);
xnor U16220 (N_16220,N_15342,N_15596);
and U16221 (N_16221,N_15245,N_15596);
nand U16222 (N_16222,N_15358,N_15534);
xor U16223 (N_16223,N_15193,N_15536);
and U16224 (N_16224,N_15094,N_15149);
or U16225 (N_16225,N_15480,N_15248);
and U16226 (N_16226,N_15435,N_15175);
nor U16227 (N_16227,N_15138,N_15578);
and U16228 (N_16228,N_15342,N_15139);
and U16229 (N_16229,N_15133,N_15056);
nor U16230 (N_16230,N_15089,N_15227);
and U16231 (N_16231,N_15578,N_15489);
xnor U16232 (N_16232,N_15389,N_15251);
nor U16233 (N_16233,N_15186,N_15583);
nor U16234 (N_16234,N_15455,N_15198);
nand U16235 (N_16235,N_15075,N_15515);
xor U16236 (N_16236,N_15622,N_15284);
xnor U16237 (N_16237,N_15088,N_15036);
or U16238 (N_16238,N_15519,N_15329);
and U16239 (N_16239,N_15619,N_15421);
and U16240 (N_16240,N_15259,N_15064);
nand U16241 (N_16241,N_15156,N_15106);
or U16242 (N_16242,N_15579,N_15552);
or U16243 (N_16243,N_15550,N_15527);
or U16244 (N_16244,N_15558,N_15462);
or U16245 (N_16245,N_15089,N_15238);
and U16246 (N_16246,N_15385,N_15451);
and U16247 (N_16247,N_15273,N_15192);
or U16248 (N_16248,N_15495,N_15211);
and U16249 (N_16249,N_15533,N_15540);
nand U16250 (N_16250,N_16134,N_15848);
nand U16251 (N_16251,N_15701,N_16054);
and U16252 (N_16252,N_15954,N_16114);
or U16253 (N_16253,N_16218,N_15722);
or U16254 (N_16254,N_16106,N_16100);
xor U16255 (N_16255,N_16008,N_16065);
and U16256 (N_16256,N_15869,N_15797);
xnor U16257 (N_16257,N_15929,N_16188);
and U16258 (N_16258,N_16240,N_15888);
or U16259 (N_16259,N_15827,N_15991);
nor U16260 (N_16260,N_15667,N_16174);
nor U16261 (N_16261,N_15661,N_16017);
and U16262 (N_16262,N_16050,N_16057);
nor U16263 (N_16263,N_16052,N_16047);
and U16264 (N_16264,N_15897,N_15750);
xor U16265 (N_16265,N_15939,N_15863);
nand U16266 (N_16266,N_16204,N_15705);
and U16267 (N_16267,N_15909,N_16150);
or U16268 (N_16268,N_15653,N_15889);
or U16269 (N_16269,N_15772,N_15833);
nor U16270 (N_16270,N_16042,N_16141);
and U16271 (N_16271,N_15799,N_15898);
and U16272 (N_16272,N_16233,N_16023);
nand U16273 (N_16273,N_16200,N_15912);
nand U16274 (N_16274,N_16142,N_15955);
and U16275 (N_16275,N_15710,N_15652);
or U16276 (N_16276,N_15822,N_15680);
nor U16277 (N_16277,N_15813,N_16128);
nor U16278 (N_16278,N_16104,N_15738);
or U16279 (N_16279,N_15695,N_15669);
nor U16280 (N_16280,N_16182,N_15875);
nor U16281 (N_16281,N_15636,N_16024);
nand U16282 (N_16282,N_15858,N_15974);
nor U16283 (N_16283,N_15989,N_16093);
nor U16284 (N_16284,N_15690,N_15730);
and U16285 (N_16285,N_16167,N_15966);
and U16286 (N_16286,N_15824,N_15718);
nand U16287 (N_16287,N_15994,N_15879);
and U16288 (N_16288,N_15693,N_16058);
nor U16289 (N_16289,N_15834,N_15656);
and U16290 (N_16290,N_15905,N_15812);
xor U16291 (N_16291,N_16078,N_15704);
xor U16292 (N_16292,N_15643,N_15684);
nand U16293 (N_16293,N_15655,N_16007);
nor U16294 (N_16294,N_15764,N_15628);
and U16295 (N_16295,N_16014,N_15745);
nor U16296 (N_16296,N_16116,N_16235);
nand U16297 (N_16297,N_15681,N_15884);
xor U16298 (N_16298,N_15950,N_15685);
nand U16299 (N_16299,N_16119,N_15658);
and U16300 (N_16300,N_15790,N_16028);
xor U16301 (N_16301,N_15860,N_15671);
nand U16302 (N_16302,N_15696,N_15990);
nand U16303 (N_16303,N_15765,N_15774);
and U16304 (N_16304,N_16232,N_16196);
xor U16305 (N_16305,N_16207,N_15675);
nand U16306 (N_16306,N_16230,N_15779);
and U16307 (N_16307,N_15885,N_15845);
xnor U16308 (N_16308,N_16103,N_16067);
xor U16309 (N_16309,N_15694,N_15717);
or U16310 (N_16310,N_16064,N_16153);
nor U16311 (N_16311,N_15677,N_16126);
nor U16312 (N_16312,N_15753,N_16236);
and U16313 (N_16313,N_16227,N_15712);
xnor U16314 (N_16314,N_15719,N_15944);
nor U16315 (N_16315,N_16055,N_15721);
or U16316 (N_16316,N_15956,N_15964);
xor U16317 (N_16317,N_16069,N_16178);
nand U16318 (N_16318,N_15793,N_16031);
or U16319 (N_16319,N_15842,N_15791);
or U16320 (N_16320,N_15855,N_15933);
or U16321 (N_16321,N_15672,N_15787);
and U16322 (N_16322,N_16193,N_15780);
nor U16323 (N_16323,N_15940,N_16076);
nor U16324 (N_16324,N_15917,N_16094);
nor U16325 (N_16325,N_16185,N_16013);
and U16326 (N_16326,N_16090,N_15918);
nand U16327 (N_16327,N_16181,N_16091);
and U16328 (N_16328,N_15843,N_15647);
nor U16329 (N_16329,N_15882,N_15640);
and U16330 (N_16330,N_15706,N_16086);
nor U16331 (N_16331,N_15851,N_16155);
nand U16332 (N_16332,N_16077,N_16049);
xor U16333 (N_16333,N_16095,N_15691);
or U16334 (N_16334,N_15818,N_15747);
xnor U16335 (N_16335,N_15945,N_16175);
xnor U16336 (N_16336,N_15935,N_15692);
xor U16337 (N_16337,N_15883,N_16140);
or U16338 (N_16338,N_16165,N_16187);
or U16339 (N_16339,N_16074,N_15659);
nand U16340 (N_16340,N_15798,N_16189);
and U16341 (N_16341,N_15642,N_15686);
or U16342 (N_16342,N_16039,N_15626);
or U16343 (N_16343,N_15911,N_15902);
nor U16344 (N_16344,N_16044,N_16159);
xor U16345 (N_16345,N_15679,N_15714);
nor U16346 (N_16346,N_15825,N_16118);
nand U16347 (N_16347,N_15984,N_15631);
nand U16348 (N_16348,N_16161,N_15922);
and U16349 (N_16349,N_15896,N_15689);
or U16350 (N_16350,N_15708,N_15648);
nand U16351 (N_16351,N_15998,N_15887);
or U16352 (N_16352,N_15785,N_16063);
nand U16353 (N_16353,N_15716,N_15763);
nand U16354 (N_16354,N_15670,N_15811);
and U16355 (N_16355,N_16152,N_16136);
nor U16356 (N_16356,N_15914,N_16247);
or U16357 (N_16357,N_15709,N_15934);
and U16358 (N_16358,N_16062,N_15649);
nand U16359 (N_16359,N_15816,N_16168);
nor U16360 (N_16360,N_15947,N_16171);
nand U16361 (N_16361,N_16190,N_16244);
nor U16362 (N_16362,N_15711,N_15891);
xor U16363 (N_16363,N_15949,N_16221);
xnor U16364 (N_16364,N_16032,N_15776);
or U16365 (N_16365,N_16217,N_16110);
nand U16366 (N_16366,N_15923,N_15702);
xnor U16367 (N_16367,N_15938,N_15996);
and U16368 (N_16368,N_15838,N_15641);
nand U16369 (N_16369,N_16082,N_16004);
nand U16370 (N_16370,N_15899,N_16087);
nor U16371 (N_16371,N_15874,N_16170);
xor U16372 (N_16372,N_15846,N_15856);
nor U16373 (N_16373,N_16071,N_15729);
xor U16374 (N_16374,N_15751,N_15726);
nand U16375 (N_16375,N_15740,N_15778);
and U16376 (N_16376,N_15660,N_15830);
nand U16377 (N_16377,N_15847,N_16143);
or U16378 (N_16378,N_16010,N_16029);
nor U16379 (N_16379,N_15928,N_16210);
xor U16380 (N_16380,N_16000,N_15635);
and U16381 (N_16381,N_15639,N_15756);
nand U16382 (N_16382,N_16117,N_16092);
nor U16383 (N_16383,N_16160,N_15937);
nand U16384 (N_16384,N_15892,N_16009);
and U16385 (N_16385,N_15971,N_16098);
nor U16386 (N_16386,N_15650,N_15881);
nand U16387 (N_16387,N_15699,N_16121);
nor U16388 (N_16388,N_16146,N_16149);
and U16389 (N_16389,N_15979,N_16172);
or U16390 (N_16390,N_15826,N_15796);
nor U16391 (N_16391,N_15724,N_16154);
nand U16392 (N_16392,N_16073,N_15900);
or U16393 (N_16393,N_15703,N_15895);
nand U16394 (N_16394,N_16113,N_16075);
or U16395 (N_16395,N_15638,N_16022);
or U16396 (N_16396,N_16249,N_15735);
nand U16397 (N_16397,N_15977,N_16206);
or U16398 (N_16398,N_15807,N_15629);
xor U16399 (N_16399,N_16016,N_16176);
xor U16400 (N_16400,N_15644,N_16226);
nor U16401 (N_16401,N_15829,N_15844);
nor U16402 (N_16402,N_16043,N_15821);
nand U16403 (N_16403,N_15697,N_15853);
or U16404 (N_16404,N_16215,N_16105);
nor U16405 (N_16405,N_15678,N_16056);
and U16406 (N_16406,N_16068,N_15803);
or U16407 (N_16407,N_15687,N_15982);
nor U16408 (N_16408,N_16179,N_15840);
or U16409 (N_16409,N_16132,N_16151);
or U16410 (N_16410,N_15878,N_15809);
nor U16411 (N_16411,N_16133,N_15698);
nand U16412 (N_16412,N_15806,N_15866);
or U16413 (N_16413,N_16184,N_15828);
and U16414 (N_16414,N_15664,N_16197);
and U16415 (N_16415,N_16231,N_15668);
nand U16416 (N_16416,N_15713,N_15849);
xor U16417 (N_16417,N_15666,N_16015);
or U16418 (N_16418,N_16245,N_16194);
xor U16419 (N_16419,N_15645,N_15980);
or U16420 (N_16420,N_15688,N_15960);
and U16421 (N_16421,N_15962,N_15771);
nor U16422 (N_16422,N_15737,N_15748);
nor U16423 (N_16423,N_16001,N_15723);
or U16424 (N_16424,N_16080,N_16101);
or U16425 (N_16425,N_15983,N_15852);
and U16426 (N_16426,N_15800,N_15720);
and U16427 (N_16427,N_16137,N_15676);
or U16428 (N_16428,N_16222,N_15894);
nor U16429 (N_16429,N_16239,N_15854);
nor U16430 (N_16430,N_16124,N_15728);
and U16431 (N_16431,N_15924,N_16180);
xnor U16432 (N_16432,N_15963,N_16243);
xor U16433 (N_16433,N_15981,N_15864);
and U16434 (N_16434,N_15744,N_15759);
or U16435 (N_16435,N_16059,N_15732);
or U16436 (N_16436,N_16003,N_15646);
or U16437 (N_16437,N_15760,N_15915);
or U16438 (N_16438,N_16212,N_15657);
nor U16439 (N_16439,N_15755,N_15727);
nand U16440 (N_16440,N_16051,N_15767);
xor U16441 (N_16441,N_15992,N_15739);
or U16442 (N_16442,N_16241,N_15943);
or U16443 (N_16443,N_15741,N_15865);
nand U16444 (N_16444,N_15967,N_15777);
xor U16445 (N_16445,N_16237,N_15769);
nand U16446 (N_16446,N_15784,N_15919);
xor U16447 (N_16447,N_16108,N_16025);
xor U16448 (N_16448,N_16203,N_16242);
nand U16449 (N_16449,N_16061,N_15682);
xor U16450 (N_16450,N_15789,N_15832);
nor U16451 (N_16451,N_15987,N_16053);
nor U16452 (N_16452,N_16102,N_16085);
nor U16453 (N_16453,N_15758,N_15958);
or U16454 (N_16454,N_16035,N_15975);
or U16455 (N_16455,N_16209,N_16041);
nand U16456 (N_16456,N_16070,N_15819);
and U16457 (N_16457,N_16202,N_16169);
or U16458 (N_16458,N_15988,N_16107);
and U16459 (N_16459,N_16211,N_15948);
nor U16460 (N_16460,N_15859,N_16198);
and U16461 (N_16461,N_16139,N_16224);
and U16462 (N_16462,N_16125,N_15903);
and U16463 (N_16463,N_15795,N_15872);
nand U16464 (N_16464,N_16219,N_16138);
and U16465 (N_16465,N_15862,N_15927);
nand U16466 (N_16466,N_16112,N_15941);
nor U16467 (N_16467,N_15986,N_16157);
nor U16468 (N_16468,N_15876,N_16123);
or U16469 (N_16469,N_15880,N_16177);
and U16470 (N_16470,N_16213,N_16191);
and U16471 (N_16471,N_15766,N_15742);
xnor U16472 (N_16472,N_15831,N_15993);
xnor U16473 (N_16473,N_15930,N_16163);
and U16474 (N_16474,N_15707,N_16156);
nand U16475 (N_16475,N_16248,N_15634);
and U16476 (N_16476,N_15932,N_16046);
nand U16477 (N_16477,N_16173,N_16034);
nor U16478 (N_16478,N_16081,N_15752);
xnor U16479 (N_16479,N_15886,N_15976);
nor U16480 (N_16480,N_15841,N_15632);
xnor U16481 (N_16481,N_15873,N_16109);
nor U16482 (N_16482,N_16223,N_15999);
xnor U16483 (N_16483,N_15957,N_15953);
or U16484 (N_16484,N_15916,N_15861);
and U16485 (N_16485,N_16205,N_15651);
xor U16486 (N_16486,N_15749,N_15823);
xnor U16487 (N_16487,N_16111,N_15970);
nand U16488 (N_16488,N_16164,N_15768);
xor U16489 (N_16489,N_15673,N_15820);
or U16490 (N_16490,N_16208,N_16115);
xor U16491 (N_16491,N_15817,N_15805);
xnor U16492 (N_16492,N_15835,N_15997);
nand U16493 (N_16493,N_16238,N_16036);
nor U16494 (N_16494,N_16089,N_15978);
and U16495 (N_16495,N_16225,N_16018);
or U16496 (N_16496,N_15951,N_16229);
and U16497 (N_16497,N_16038,N_16020);
nor U16498 (N_16498,N_15746,N_15973);
and U16499 (N_16499,N_15783,N_15715);
or U16500 (N_16500,N_15952,N_15877);
nand U16501 (N_16501,N_15788,N_15782);
nor U16502 (N_16502,N_16084,N_15910);
nor U16503 (N_16503,N_15870,N_16033);
nand U16504 (N_16504,N_15808,N_15674);
nor U16505 (N_16505,N_16002,N_16129);
and U16506 (N_16506,N_15810,N_16088);
or U16507 (N_16507,N_15662,N_15867);
xnor U16508 (N_16508,N_16048,N_15901);
xnor U16509 (N_16509,N_16214,N_16006);
or U16510 (N_16510,N_16019,N_16079);
xor U16511 (N_16511,N_16097,N_15627);
and U16512 (N_16512,N_15804,N_16027);
nand U16513 (N_16513,N_16045,N_16216);
nor U16514 (N_16514,N_15936,N_16145);
xor U16515 (N_16515,N_15743,N_16099);
nor U16516 (N_16516,N_16122,N_15761);
nand U16517 (N_16517,N_15754,N_15700);
xnor U16518 (N_16518,N_15815,N_15942);
nand U16519 (N_16519,N_16192,N_15762);
or U16520 (N_16520,N_16148,N_15931);
or U16521 (N_16521,N_15654,N_15961);
nor U16522 (N_16522,N_15733,N_16158);
and U16523 (N_16523,N_15965,N_15868);
and U16524 (N_16524,N_16060,N_15959);
or U16525 (N_16525,N_16072,N_16147);
nor U16526 (N_16526,N_16037,N_15890);
and U16527 (N_16527,N_15906,N_16012);
and U16528 (N_16528,N_15801,N_16228);
or U16529 (N_16529,N_15857,N_16120);
or U16530 (N_16530,N_15781,N_16166);
and U16531 (N_16531,N_15972,N_15968);
and U16532 (N_16532,N_16131,N_15871);
and U16533 (N_16533,N_16096,N_15839);
or U16534 (N_16534,N_16005,N_15637);
xor U16535 (N_16535,N_16183,N_15625);
nor U16536 (N_16536,N_15770,N_16021);
nor U16537 (N_16537,N_15850,N_16246);
nand U16538 (N_16538,N_16083,N_15921);
or U16539 (N_16539,N_16186,N_15913);
and U16540 (N_16540,N_15665,N_15893);
xor U16541 (N_16541,N_15907,N_15925);
and U16542 (N_16542,N_15731,N_15836);
and U16543 (N_16543,N_16011,N_15926);
and U16544 (N_16544,N_15794,N_15630);
or U16545 (N_16545,N_15837,N_15663);
nor U16546 (N_16546,N_16199,N_16040);
nand U16547 (N_16547,N_15904,N_16127);
and U16548 (N_16548,N_15908,N_15946);
nor U16549 (N_16549,N_16162,N_16201);
xor U16550 (N_16550,N_15757,N_15775);
nor U16551 (N_16551,N_15736,N_16026);
xor U16552 (N_16552,N_15683,N_15633);
and U16553 (N_16553,N_16130,N_16030);
nor U16554 (N_16554,N_15773,N_15786);
nor U16555 (N_16555,N_15802,N_16220);
xnor U16556 (N_16556,N_15814,N_16066);
nand U16557 (N_16557,N_16144,N_15792);
and U16558 (N_16558,N_15985,N_15995);
or U16559 (N_16559,N_16195,N_15725);
nor U16560 (N_16560,N_15734,N_15920);
nand U16561 (N_16561,N_16234,N_15969);
xor U16562 (N_16562,N_16135,N_16003);
nand U16563 (N_16563,N_15762,N_16133);
and U16564 (N_16564,N_15920,N_16103);
or U16565 (N_16565,N_16248,N_16192);
nor U16566 (N_16566,N_15862,N_16225);
xnor U16567 (N_16567,N_15817,N_15978);
nor U16568 (N_16568,N_15721,N_15711);
nand U16569 (N_16569,N_15869,N_16214);
xnor U16570 (N_16570,N_15890,N_16099);
and U16571 (N_16571,N_16067,N_15655);
and U16572 (N_16572,N_16029,N_15980);
or U16573 (N_16573,N_16168,N_16179);
xor U16574 (N_16574,N_15797,N_15705);
xor U16575 (N_16575,N_16161,N_15774);
nor U16576 (N_16576,N_15802,N_16071);
nor U16577 (N_16577,N_15725,N_16098);
or U16578 (N_16578,N_16215,N_15903);
nand U16579 (N_16579,N_16082,N_15988);
xnor U16580 (N_16580,N_16119,N_16026);
xor U16581 (N_16581,N_16025,N_15860);
nor U16582 (N_16582,N_16036,N_15980);
nor U16583 (N_16583,N_16212,N_15761);
nor U16584 (N_16584,N_15682,N_15642);
or U16585 (N_16585,N_15760,N_15633);
nand U16586 (N_16586,N_16173,N_16027);
and U16587 (N_16587,N_15975,N_15825);
and U16588 (N_16588,N_16126,N_16003);
xnor U16589 (N_16589,N_15723,N_15652);
or U16590 (N_16590,N_15816,N_16127);
nor U16591 (N_16591,N_15896,N_15634);
xnor U16592 (N_16592,N_15970,N_16085);
and U16593 (N_16593,N_15893,N_15748);
xor U16594 (N_16594,N_16024,N_16208);
nand U16595 (N_16595,N_15736,N_16121);
nand U16596 (N_16596,N_16125,N_15964);
nand U16597 (N_16597,N_15898,N_15676);
or U16598 (N_16598,N_15707,N_16225);
and U16599 (N_16599,N_16025,N_15698);
nor U16600 (N_16600,N_15759,N_15827);
or U16601 (N_16601,N_16108,N_16022);
nand U16602 (N_16602,N_16134,N_16244);
xor U16603 (N_16603,N_15802,N_15823);
nor U16604 (N_16604,N_15711,N_15850);
and U16605 (N_16605,N_15645,N_15794);
nand U16606 (N_16606,N_16150,N_16017);
xor U16607 (N_16607,N_15900,N_15711);
or U16608 (N_16608,N_15780,N_15849);
nor U16609 (N_16609,N_15710,N_16092);
xnor U16610 (N_16610,N_15687,N_15862);
or U16611 (N_16611,N_15798,N_16165);
xor U16612 (N_16612,N_15663,N_15732);
nand U16613 (N_16613,N_15961,N_16073);
nand U16614 (N_16614,N_15810,N_16129);
and U16615 (N_16615,N_15915,N_15852);
xnor U16616 (N_16616,N_15874,N_15731);
xor U16617 (N_16617,N_15821,N_15737);
or U16618 (N_16618,N_16039,N_16031);
nand U16619 (N_16619,N_15673,N_15632);
or U16620 (N_16620,N_15723,N_15864);
and U16621 (N_16621,N_15905,N_15764);
nor U16622 (N_16622,N_15645,N_16098);
xor U16623 (N_16623,N_15686,N_15712);
nor U16624 (N_16624,N_15799,N_16133);
and U16625 (N_16625,N_15865,N_15998);
xnor U16626 (N_16626,N_15974,N_16159);
or U16627 (N_16627,N_16178,N_16009);
nor U16628 (N_16628,N_16152,N_16143);
xnor U16629 (N_16629,N_15680,N_15932);
or U16630 (N_16630,N_15639,N_16165);
xor U16631 (N_16631,N_16142,N_16132);
or U16632 (N_16632,N_15749,N_16112);
or U16633 (N_16633,N_15692,N_15775);
xor U16634 (N_16634,N_15912,N_16105);
xor U16635 (N_16635,N_16144,N_16049);
nor U16636 (N_16636,N_16045,N_15726);
xor U16637 (N_16637,N_16105,N_16210);
or U16638 (N_16638,N_16218,N_15757);
or U16639 (N_16639,N_16137,N_16014);
or U16640 (N_16640,N_16164,N_15933);
and U16641 (N_16641,N_15811,N_15676);
nor U16642 (N_16642,N_16073,N_16025);
nor U16643 (N_16643,N_16013,N_16160);
and U16644 (N_16644,N_15762,N_15914);
xnor U16645 (N_16645,N_15626,N_16185);
xor U16646 (N_16646,N_16130,N_16064);
and U16647 (N_16647,N_15681,N_16071);
nand U16648 (N_16648,N_16003,N_16037);
xnor U16649 (N_16649,N_16098,N_15749);
xnor U16650 (N_16650,N_15911,N_15839);
or U16651 (N_16651,N_16143,N_15697);
nor U16652 (N_16652,N_16201,N_15782);
and U16653 (N_16653,N_15837,N_16108);
and U16654 (N_16654,N_16248,N_15814);
nand U16655 (N_16655,N_16244,N_15942);
nor U16656 (N_16656,N_16091,N_16178);
or U16657 (N_16657,N_16211,N_16217);
nor U16658 (N_16658,N_15849,N_15942);
nor U16659 (N_16659,N_15844,N_15781);
nand U16660 (N_16660,N_16109,N_15929);
or U16661 (N_16661,N_16203,N_16012);
nor U16662 (N_16662,N_15804,N_15991);
or U16663 (N_16663,N_15864,N_15857);
nor U16664 (N_16664,N_15932,N_15927);
xnor U16665 (N_16665,N_15829,N_15910);
and U16666 (N_16666,N_15820,N_15868);
and U16667 (N_16667,N_15726,N_16032);
nor U16668 (N_16668,N_16042,N_16232);
nor U16669 (N_16669,N_15838,N_16050);
and U16670 (N_16670,N_15679,N_15979);
nor U16671 (N_16671,N_15674,N_15750);
nor U16672 (N_16672,N_15773,N_15646);
and U16673 (N_16673,N_16227,N_15884);
and U16674 (N_16674,N_15628,N_16006);
or U16675 (N_16675,N_16163,N_15923);
nor U16676 (N_16676,N_16173,N_15894);
and U16677 (N_16677,N_16107,N_15945);
nor U16678 (N_16678,N_15787,N_15683);
and U16679 (N_16679,N_15742,N_15888);
xnor U16680 (N_16680,N_15924,N_16204);
nor U16681 (N_16681,N_15932,N_15672);
and U16682 (N_16682,N_15888,N_15921);
nor U16683 (N_16683,N_15893,N_15664);
or U16684 (N_16684,N_15785,N_16080);
or U16685 (N_16685,N_16064,N_15628);
nand U16686 (N_16686,N_16045,N_15732);
and U16687 (N_16687,N_15904,N_16107);
or U16688 (N_16688,N_15862,N_16079);
nand U16689 (N_16689,N_15992,N_16034);
nor U16690 (N_16690,N_16123,N_15789);
or U16691 (N_16691,N_16055,N_16205);
and U16692 (N_16692,N_15840,N_15763);
xor U16693 (N_16693,N_16223,N_16207);
xnor U16694 (N_16694,N_15746,N_16087);
nand U16695 (N_16695,N_15926,N_15712);
or U16696 (N_16696,N_16153,N_15829);
nor U16697 (N_16697,N_15994,N_15888);
or U16698 (N_16698,N_15870,N_16050);
or U16699 (N_16699,N_16021,N_16165);
xor U16700 (N_16700,N_15980,N_16027);
and U16701 (N_16701,N_15926,N_15715);
nor U16702 (N_16702,N_16201,N_15844);
nand U16703 (N_16703,N_15730,N_15665);
and U16704 (N_16704,N_15712,N_15935);
nand U16705 (N_16705,N_15692,N_15909);
and U16706 (N_16706,N_15693,N_16234);
xor U16707 (N_16707,N_15914,N_16182);
and U16708 (N_16708,N_16243,N_16137);
and U16709 (N_16709,N_15791,N_15935);
nor U16710 (N_16710,N_15656,N_16144);
nor U16711 (N_16711,N_15765,N_15633);
and U16712 (N_16712,N_16247,N_16025);
nand U16713 (N_16713,N_15995,N_15772);
nor U16714 (N_16714,N_15866,N_15751);
and U16715 (N_16715,N_15962,N_15843);
nor U16716 (N_16716,N_16215,N_15739);
and U16717 (N_16717,N_15912,N_15877);
and U16718 (N_16718,N_15775,N_15680);
or U16719 (N_16719,N_15849,N_16112);
nand U16720 (N_16720,N_15967,N_16240);
or U16721 (N_16721,N_15950,N_15779);
xor U16722 (N_16722,N_15746,N_15979);
nor U16723 (N_16723,N_16069,N_15844);
or U16724 (N_16724,N_15961,N_15664);
and U16725 (N_16725,N_15667,N_15827);
or U16726 (N_16726,N_15813,N_16113);
xnor U16727 (N_16727,N_15832,N_15962);
nor U16728 (N_16728,N_16107,N_15814);
nand U16729 (N_16729,N_15778,N_15703);
nand U16730 (N_16730,N_15981,N_15747);
xnor U16731 (N_16731,N_15837,N_16141);
nand U16732 (N_16732,N_16061,N_16119);
and U16733 (N_16733,N_15965,N_15802);
xor U16734 (N_16734,N_15856,N_15727);
nor U16735 (N_16735,N_15636,N_16244);
and U16736 (N_16736,N_15904,N_15694);
xor U16737 (N_16737,N_15711,N_15855);
nand U16738 (N_16738,N_15948,N_15874);
or U16739 (N_16739,N_15755,N_16198);
nand U16740 (N_16740,N_15831,N_15912);
or U16741 (N_16741,N_15760,N_15673);
or U16742 (N_16742,N_16075,N_15722);
nor U16743 (N_16743,N_15837,N_15757);
and U16744 (N_16744,N_15702,N_15928);
xnor U16745 (N_16745,N_16067,N_16249);
and U16746 (N_16746,N_16027,N_16202);
xnor U16747 (N_16747,N_15841,N_16165);
nand U16748 (N_16748,N_15752,N_16181);
nand U16749 (N_16749,N_15894,N_15944);
nor U16750 (N_16750,N_16140,N_16049);
xor U16751 (N_16751,N_16096,N_16007);
and U16752 (N_16752,N_16177,N_16226);
nand U16753 (N_16753,N_15907,N_15803);
or U16754 (N_16754,N_15883,N_16211);
nor U16755 (N_16755,N_16061,N_15778);
or U16756 (N_16756,N_15746,N_16150);
or U16757 (N_16757,N_16146,N_16047);
xnor U16758 (N_16758,N_16010,N_16094);
nor U16759 (N_16759,N_15658,N_15794);
and U16760 (N_16760,N_15912,N_15981);
or U16761 (N_16761,N_16202,N_15685);
nor U16762 (N_16762,N_16166,N_15638);
xor U16763 (N_16763,N_15689,N_16026);
nor U16764 (N_16764,N_15841,N_15700);
xor U16765 (N_16765,N_16154,N_15880);
xor U16766 (N_16766,N_15774,N_16011);
and U16767 (N_16767,N_16100,N_15722);
and U16768 (N_16768,N_15727,N_15752);
nor U16769 (N_16769,N_15742,N_15755);
nor U16770 (N_16770,N_15770,N_15812);
and U16771 (N_16771,N_16045,N_15799);
nand U16772 (N_16772,N_15719,N_15936);
or U16773 (N_16773,N_15904,N_15916);
nor U16774 (N_16774,N_15990,N_15847);
nand U16775 (N_16775,N_16021,N_15773);
and U16776 (N_16776,N_15943,N_15688);
xor U16777 (N_16777,N_15804,N_16128);
and U16778 (N_16778,N_16082,N_15773);
nor U16779 (N_16779,N_15927,N_15777);
nand U16780 (N_16780,N_15917,N_16131);
or U16781 (N_16781,N_15902,N_15644);
nand U16782 (N_16782,N_15743,N_16228);
nand U16783 (N_16783,N_15839,N_16174);
nor U16784 (N_16784,N_15844,N_15950);
nor U16785 (N_16785,N_15725,N_15635);
or U16786 (N_16786,N_15897,N_16008);
xnor U16787 (N_16787,N_15673,N_15738);
or U16788 (N_16788,N_16171,N_15867);
and U16789 (N_16789,N_16221,N_15675);
nand U16790 (N_16790,N_15884,N_16245);
or U16791 (N_16791,N_16054,N_15958);
xnor U16792 (N_16792,N_15995,N_15911);
nor U16793 (N_16793,N_15625,N_15955);
and U16794 (N_16794,N_16025,N_15911);
nor U16795 (N_16795,N_15940,N_15686);
nand U16796 (N_16796,N_15991,N_15643);
nand U16797 (N_16797,N_15662,N_15638);
and U16798 (N_16798,N_16172,N_16109);
or U16799 (N_16799,N_15639,N_15880);
and U16800 (N_16800,N_15868,N_16041);
nor U16801 (N_16801,N_16209,N_15943);
and U16802 (N_16802,N_16074,N_15804);
nand U16803 (N_16803,N_15763,N_15822);
and U16804 (N_16804,N_16058,N_16167);
or U16805 (N_16805,N_16048,N_15928);
nor U16806 (N_16806,N_16102,N_16088);
xnor U16807 (N_16807,N_15893,N_15798);
and U16808 (N_16808,N_15630,N_16164);
nand U16809 (N_16809,N_15709,N_15646);
nor U16810 (N_16810,N_16246,N_16140);
and U16811 (N_16811,N_16189,N_16154);
and U16812 (N_16812,N_15911,N_16145);
xor U16813 (N_16813,N_15641,N_15726);
or U16814 (N_16814,N_15779,N_15631);
xnor U16815 (N_16815,N_16097,N_16178);
xor U16816 (N_16816,N_15626,N_15937);
or U16817 (N_16817,N_15662,N_15635);
and U16818 (N_16818,N_15795,N_15863);
nand U16819 (N_16819,N_16035,N_15646);
xnor U16820 (N_16820,N_15876,N_16001);
xnor U16821 (N_16821,N_15937,N_15922);
and U16822 (N_16822,N_15858,N_15989);
nand U16823 (N_16823,N_16000,N_15983);
xor U16824 (N_16824,N_16225,N_16030);
or U16825 (N_16825,N_16120,N_15968);
nand U16826 (N_16826,N_15860,N_16062);
nand U16827 (N_16827,N_16202,N_15753);
nand U16828 (N_16828,N_15811,N_16199);
nand U16829 (N_16829,N_15731,N_15781);
or U16830 (N_16830,N_15956,N_16131);
nand U16831 (N_16831,N_15938,N_15870);
or U16832 (N_16832,N_16112,N_16086);
xor U16833 (N_16833,N_15705,N_16190);
xnor U16834 (N_16834,N_16162,N_16164);
nor U16835 (N_16835,N_15688,N_15961);
or U16836 (N_16836,N_15933,N_15982);
and U16837 (N_16837,N_16046,N_15983);
or U16838 (N_16838,N_15859,N_15677);
nor U16839 (N_16839,N_15904,N_16064);
or U16840 (N_16840,N_16009,N_16066);
or U16841 (N_16841,N_16127,N_15989);
and U16842 (N_16842,N_15965,N_16193);
and U16843 (N_16843,N_15707,N_16211);
nor U16844 (N_16844,N_15931,N_15711);
nand U16845 (N_16845,N_16143,N_16247);
and U16846 (N_16846,N_15727,N_15724);
and U16847 (N_16847,N_15815,N_16215);
nand U16848 (N_16848,N_15955,N_15900);
nand U16849 (N_16849,N_16197,N_15684);
or U16850 (N_16850,N_15711,N_15703);
xor U16851 (N_16851,N_16057,N_15932);
xor U16852 (N_16852,N_16190,N_16017);
or U16853 (N_16853,N_15698,N_16032);
or U16854 (N_16854,N_15739,N_16212);
nand U16855 (N_16855,N_15849,N_15950);
nand U16856 (N_16856,N_16003,N_15976);
xnor U16857 (N_16857,N_15748,N_15915);
or U16858 (N_16858,N_15729,N_16039);
and U16859 (N_16859,N_15764,N_15934);
xnor U16860 (N_16860,N_15652,N_16226);
nand U16861 (N_16861,N_15789,N_16034);
nand U16862 (N_16862,N_16133,N_16075);
nand U16863 (N_16863,N_15630,N_15971);
and U16864 (N_16864,N_15883,N_16214);
nand U16865 (N_16865,N_16206,N_15753);
nor U16866 (N_16866,N_16029,N_15826);
nand U16867 (N_16867,N_15750,N_15912);
and U16868 (N_16868,N_15870,N_15676);
and U16869 (N_16869,N_15678,N_15959);
or U16870 (N_16870,N_15728,N_15661);
and U16871 (N_16871,N_16166,N_15643);
or U16872 (N_16872,N_16172,N_16208);
xor U16873 (N_16873,N_15718,N_15653);
nand U16874 (N_16874,N_15751,N_16051);
or U16875 (N_16875,N_16848,N_16429);
nor U16876 (N_16876,N_16324,N_16763);
nor U16877 (N_16877,N_16451,N_16369);
nor U16878 (N_16878,N_16635,N_16803);
nand U16879 (N_16879,N_16439,N_16604);
xor U16880 (N_16880,N_16378,N_16660);
nand U16881 (N_16881,N_16301,N_16488);
and U16882 (N_16882,N_16323,N_16820);
xnor U16883 (N_16883,N_16550,N_16257);
xor U16884 (N_16884,N_16606,N_16628);
nor U16885 (N_16885,N_16362,N_16713);
or U16886 (N_16886,N_16574,N_16581);
or U16887 (N_16887,N_16529,N_16793);
or U16888 (N_16888,N_16302,N_16769);
nand U16889 (N_16889,N_16464,N_16477);
and U16890 (N_16890,N_16814,N_16521);
nor U16891 (N_16891,N_16554,N_16570);
nand U16892 (N_16892,N_16475,N_16780);
nor U16893 (N_16893,N_16449,N_16588);
xor U16894 (N_16894,N_16856,N_16473);
xor U16895 (N_16895,N_16357,N_16519);
xor U16896 (N_16896,N_16263,N_16250);
and U16897 (N_16897,N_16458,N_16617);
xnor U16898 (N_16898,N_16664,N_16643);
xor U16899 (N_16899,N_16440,N_16613);
nand U16900 (N_16900,N_16657,N_16382);
xnor U16901 (N_16901,N_16869,N_16747);
xor U16902 (N_16902,N_16602,N_16497);
nand U16903 (N_16903,N_16825,N_16322);
or U16904 (N_16904,N_16865,N_16446);
nand U16905 (N_16905,N_16259,N_16751);
or U16906 (N_16906,N_16867,N_16400);
or U16907 (N_16907,N_16425,N_16536);
nor U16908 (N_16908,N_16376,N_16444);
or U16909 (N_16909,N_16471,N_16494);
nor U16910 (N_16910,N_16873,N_16334);
and U16911 (N_16911,N_16579,N_16796);
or U16912 (N_16912,N_16538,N_16804);
and U16913 (N_16913,N_16505,N_16864);
nor U16914 (N_16914,N_16359,N_16491);
nand U16915 (N_16915,N_16732,N_16459);
xor U16916 (N_16916,N_16725,N_16789);
nor U16917 (N_16917,N_16582,N_16781);
xnor U16918 (N_16918,N_16540,N_16517);
or U16919 (N_16919,N_16450,N_16474);
and U16920 (N_16920,N_16799,N_16253);
nor U16921 (N_16921,N_16437,N_16347);
nor U16922 (N_16922,N_16590,N_16832);
xnor U16923 (N_16923,N_16808,N_16516);
nand U16924 (N_16924,N_16443,N_16315);
xor U16925 (N_16925,N_16397,N_16310);
xor U16926 (N_16926,N_16460,N_16702);
xnor U16927 (N_16927,N_16598,N_16348);
or U16928 (N_16928,N_16453,N_16679);
or U16929 (N_16929,N_16341,N_16871);
or U16930 (N_16930,N_16801,N_16828);
or U16931 (N_16931,N_16767,N_16276);
or U16932 (N_16932,N_16577,N_16327);
xor U16933 (N_16933,N_16578,N_16823);
or U16934 (N_16934,N_16407,N_16622);
or U16935 (N_16935,N_16788,N_16774);
and U16936 (N_16936,N_16470,N_16268);
nand U16937 (N_16937,N_16812,N_16618);
and U16938 (N_16938,N_16546,N_16467);
or U16939 (N_16939,N_16375,N_16696);
or U16940 (N_16940,N_16827,N_16409);
nor U16941 (N_16941,N_16633,N_16740);
or U16942 (N_16942,N_16686,N_16523);
nand U16943 (N_16943,N_16699,N_16843);
or U16944 (N_16944,N_16370,N_16851);
nor U16945 (N_16945,N_16379,N_16462);
nor U16946 (N_16946,N_16487,N_16743);
nor U16947 (N_16947,N_16594,N_16313);
nor U16948 (N_16948,N_16829,N_16668);
nor U16949 (N_16949,N_16316,N_16526);
nor U16950 (N_16950,N_16279,N_16716);
xor U16951 (N_16951,N_16291,N_16353);
nor U16952 (N_16952,N_16564,N_16714);
or U16953 (N_16953,N_16727,N_16768);
nand U16954 (N_16954,N_16294,N_16807);
nand U16955 (N_16955,N_16469,N_16481);
or U16956 (N_16956,N_16455,N_16508);
or U16957 (N_16957,N_16500,N_16720);
or U16958 (N_16958,N_16545,N_16662);
xor U16959 (N_16959,N_16326,N_16790);
or U16960 (N_16960,N_16398,N_16736);
nand U16961 (N_16961,N_16352,N_16297);
or U16962 (N_16962,N_16547,N_16433);
xnor U16963 (N_16963,N_16447,N_16381);
or U16964 (N_16964,N_16566,N_16778);
nor U16965 (N_16965,N_16558,N_16647);
xor U16966 (N_16966,N_16872,N_16603);
nand U16967 (N_16967,N_16553,N_16418);
nand U16968 (N_16968,N_16507,N_16849);
nor U16969 (N_16969,N_16625,N_16576);
nand U16970 (N_16970,N_16452,N_16358);
nor U16971 (N_16971,N_16300,N_16483);
nor U16972 (N_16972,N_16719,N_16534);
nor U16973 (N_16973,N_16824,N_16840);
nand U16974 (N_16974,N_16859,N_16502);
or U16975 (N_16975,N_16866,N_16401);
xnor U16976 (N_16976,N_16771,N_16614);
and U16977 (N_16977,N_16757,N_16766);
nand U16978 (N_16978,N_16626,N_16688);
nor U16979 (N_16979,N_16274,N_16621);
and U16980 (N_16980,N_16669,N_16412);
and U16981 (N_16981,N_16730,N_16798);
or U16982 (N_16982,N_16465,N_16676);
nor U16983 (N_16983,N_16645,N_16265);
or U16984 (N_16984,N_16785,N_16705);
nor U16985 (N_16985,N_16482,N_16329);
xnor U16986 (N_16986,N_16456,N_16853);
or U16987 (N_16987,N_16748,N_16372);
xnor U16988 (N_16988,N_16510,N_16434);
and U16989 (N_16989,N_16749,N_16765);
nand U16990 (N_16990,N_16531,N_16403);
nand U16991 (N_16991,N_16269,N_16844);
nand U16992 (N_16992,N_16742,N_16683);
nand U16993 (N_16993,N_16343,N_16770);
xor U16994 (N_16994,N_16394,N_16426);
nor U16995 (N_16995,N_16338,N_16410);
or U16996 (N_16996,N_16722,N_16364);
and U16997 (N_16997,N_16308,N_16415);
nor U16998 (N_16998,N_16288,N_16718);
nor U16999 (N_16999,N_16395,N_16834);
xnor U17000 (N_17000,N_16298,N_16320);
nand U17001 (N_17001,N_16646,N_16597);
nor U17002 (N_17002,N_16399,N_16680);
and U17003 (N_17003,N_16380,N_16396);
xnor U17004 (N_17004,N_16640,N_16729);
xor U17005 (N_17005,N_16721,N_16490);
nor U17006 (N_17006,N_16656,N_16802);
and U17007 (N_17007,N_16837,N_16572);
xor U17008 (N_17008,N_16653,N_16605);
or U17009 (N_17009,N_16822,N_16833);
nor U17010 (N_17010,N_16331,N_16484);
or U17011 (N_17011,N_16431,N_16511);
nor U17012 (N_17012,N_16363,N_16711);
nor U17013 (N_17013,N_16423,N_16715);
xnor U17014 (N_17014,N_16271,N_16651);
nor U17015 (N_17015,N_16411,N_16817);
and U17016 (N_17016,N_16659,N_16593);
nor U17017 (N_17017,N_16377,N_16775);
nor U17018 (N_17018,N_16667,N_16811);
or U17019 (N_17019,N_16607,N_16285);
or U17020 (N_17020,N_16518,N_16571);
nand U17021 (N_17021,N_16454,N_16750);
nand U17022 (N_17022,N_16530,N_16368);
or U17023 (N_17023,N_16586,N_16753);
xnor U17024 (N_17024,N_16361,N_16627);
and U17025 (N_17025,N_16670,N_16762);
or U17026 (N_17026,N_16524,N_16321);
xor U17027 (N_17027,N_16847,N_16623);
xnor U17028 (N_17028,N_16726,N_16280);
nand U17029 (N_17029,N_16461,N_16290);
xnor U17030 (N_17030,N_16703,N_16776);
xnor U17031 (N_17031,N_16665,N_16489);
xor U17032 (N_17032,N_16644,N_16346);
or U17033 (N_17033,N_16309,N_16786);
nand U17034 (N_17034,N_16835,N_16591);
nand U17035 (N_17035,N_16637,N_16528);
nand U17036 (N_17036,N_16655,N_16850);
nand U17037 (N_17037,N_16542,N_16330);
or U17038 (N_17038,N_16795,N_16266);
nor U17039 (N_17039,N_16739,N_16332);
xor U17040 (N_17040,N_16445,N_16791);
xor U17041 (N_17041,N_16701,N_16438);
nor U17042 (N_17042,N_16562,N_16286);
and U17043 (N_17043,N_16734,N_16556);
nor U17044 (N_17044,N_16709,N_16761);
and U17045 (N_17045,N_16335,N_16754);
and U17046 (N_17046,N_16312,N_16855);
xor U17047 (N_17047,N_16839,N_16800);
nor U17048 (N_17048,N_16432,N_16599);
nand U17049 (N_17049,N_16354,N_16846);
xor U17050 (N_17050,N_16672,N_16277);
or U17051 (N_17051,N_16583,N_16260);
or U17052 (N_17052,N_16784,N_16629);
nor U17053 (N_17053,N_16601,N_16503);
or U17054 (N_17054,N_16745,N_16671);
and U17055 (N_17055,N_16589,N_16402);
or U17056 (N_17056,N_16557,N_16619);
nor U17057 (N_17057,N_16306,N_16682);
xnor U17058 (N_17058,N_16374,N_16442);
nand U17059 (N_17059,N_16498,N_16448);
nor U17060 (N_17060,N_16392,N_16616);
and U17061 (N_17061,N_16311,N_16630);
or U17062 (N_17062,N_16819,N_16666);
and U17063 (N_17063,N_16319,N_16275);
and U17064 (N_17064,N_16695,N_16611);
and U17065 (N_17065,N_16639,N_16485);
nor U17066 (N_17066,N_16548,N_16794);
nand U17067 (N_17067,N_16661,N_16560);
and U17068 (N_17068,N_16854,N_16373);
and U17069 (N_17069,N_16525,N_16408);
nor U17070 (N_17070,N_16756,N_16631);
xor U17071 (N_17071,N_16841,N_16698);
xor U17072 (N_17072,N_16501,N_16813);
nand U17073 (N_17073,N_16638,N_16636);
nor U17074 (N_17074,N_16486,N_16870);
or U17075 (N_17075,N_16615,N_16388);
nor U17076 (N_17076,N_16413,N_16304);
nor U17077 (N_17077,N_16634,N_16317);
xnor U17078 (N_17078,N_16677,N_16340);
nand U17079 (N_17079,N_16584,N_16568);
xnor U17080 (N_17080,N_16648,N_16818);
nor U17081 (N_17081,N_16267,N_16385);
xnor U17082 (N_17082,N_16552,N_16792);
or U17083 (N_17083,N_16632,N_16281);
and U17084 (N_17084,N_16585,N_16532);
and U17085 (N_17085,N_16254,N_16384);
or U17086 (N_17086,N_16307,N_16731);
nand U17087 (N_17087,N_16520,N_16293);
or U17088 (N_17088,N_16805,N_16779);
or U17089 (N_17089,N_16262,N_16515);
or U17090 (N_17090,N_16251,N_16685);
and U17091 (N_17091,N_16522,N_16738);
nand U17092 (N_17092,N_16350,N_16624);
xor U17093 (N_17093,N_16816,N_16342);
and U17094 (N_17094,N_16608,N_16441);
xor U17095 (N_17095,N_16783,N_16499);
nor U17096 (N_17096,N_16472,N_16708);
nand U17097 (N_17097,N_16264,N_16533);
nand U17098 (N_17098,N_16328,N_16492);
nor U17099 (N_17099,N_16325,N_16777);
xnor U17100 (N_17100,N_16838,N_16351);
nor U17101 (N_17101,N_16365,N_16422);
xor U17102 (N_17102,N_16544,N_16305);
and U17103 (N_17103,N_16863,N_16436);
xnor U17104 (N_17104,N_16758,N_16314);
or U17105 (N_17105,N_16821,N_16504);
or U17106 (N_17106,N_16842,N_16543);
xor U17107 (N_17107,N_16691,N_16333);
nor U17108 (N_17108,N_16580,N_16512);
and U17109 (N_17109,N_16858,N_16417);
nor U17110 (N_17110,N_16383,N_16694);
or U17111 (N_17111,N_16673,N_16710);
nand U17112 (N_17112,N_16723,N_16692);
or U17113 (N_17113,N_16706,N_16687);
nand U17114 (N_17114,N_16569,N_16555);
and U17115 (N_17115,N_16336,N_16463);
nor U17116 (N_17116,N_16419,N_16700);
and U17117 (N_17117,N_16513,N_16697);
nor U17118 (N_17118,N_16292,N_16337);
nor U17119 (N_17119,N_16741,N_16712);
or U17120 (N_17120,N_16424,N_16826);
nor U17121 (N_17121,N_16421,N_16416);
nand U17122 (N_17122,N_16428,N_16296);
xnor U17123 (N_17123,N_16689,N_16600);
or U17124 (N_17124,N_16836,N_16735);
nand U17125 (N_17125,N_16693,N_16344);
xor U17126 (N_17126,N_16480,N_16874);
nand U17127 (N_17127,N_16349,N_16760);
or U17128 (N_17128,N_16371,N_16746);
xor U17129 (N_17129,N_16278,N_16420);
nand U17130 (N_17130,N_16609,N_16704);
nand U17131 (N_17131,N_16356,N_16567);
xnor U17132 (N_17132,N_16559,N_16283);
nand U17133 (N_17133,N_16389,N_16809);
and U17134 (N_17134,N_16284,N_16393);
or U17135 (N_17135,N_16258,N_16724);
xor U17136 (N_17136,N_16675,N_16592);
xor U17137 (N_17137,N_16535,N_16468);
and U17138 (N_17138,N_16537,N_16797);
or U17139 (N_17139,N_16595,N_16830);
nand U17140 (N_17140,N_16707,N_16355);
or U17141 (N_17141,N_16587,N_16642);
or U17142 (N_17142,N_16658,N_16386);
or U17143 (N_17143,N_16815,N_16541);
and U17144 (N_17144,N_16764,N_16733);
nand U17145 (N_17145,N_16345,N_16252);
or U17146 (N_17146,N_16861,N_16476);
xor U17147 (N_17147,N_16717,N_16782);
xor U17148 (N_17148,N_16360,N_16690);
and U17149 (N_17149,N_16684,N_16404);
and U17150 (N_17150,N_16272,N_16427);
or U17151 (N_17151,N_16366,N_16810);
xor U17152 (N_17152,N_16406,N_16405);
or U17153 (N_17153,N_16573,N_16561);
and U17154 (N_17154,N_16575,N_16565);
and U17155 (N_17155,N_16852,N_16457);
or U17156 (N_17156,N_16496,N_16650);
nand U17157 (N_17157,N_16787,N_16728);
nand U17158 (N_17158,N_16509,N_16549);
nor U17159 (N_17159,N_16478,N_16527);
or U17160 (N_17160,N_16282,N_16652);
or U17161 (N_17161,N_16414,N_16610);
or U17162 (N_17162,N_16430,N_16387);
xor U17163 (N_17163,N_16773,N_16752);
and U17164 (N_17164,N_16654,N_16596);
xor U17165 (N_17165,N_16506,N_16868);
or U17166 (N_17166,N_16772,N_16287);
or U17167 (N_17167,N_16295,N_16681);
and U17168 (N_17168,N_16339,N_16674);
and U17169 (N_17169,N_16303,N_16367);
or U17170 (N_17170,N_16759,N_16391);
and U17171 (N_17171,N_16860,N_16649);
xnor U17172 (N_17172,N_16493,N_16744);
and U17173 (N_17173,N_16806,N_16831);
nor U17174 (N_17174,N_16563,N_16289);
nand U17175 (N_17175,N_16318,N_16256);
or U17176 (N_17176,N_16479,N_16261);
and U17177 (N_17177,N_16299,N_16737);
nor U17178 (N_17178,N_16539,N_16641);
and U17179 (N_17179,N_16862,N_16255);
and U17180 (N_17180,N_16390,N_16845);
nor U17181 (N_17181,N_16435,N_16514);
xor U17182 (N_17182,N_16620,N_16551);
nand U17183 (N_17183,N_16857,N_16495);
nor U17184 (N_17184,N_16273,N_16466);
or U17185 (N_17185,N_16663,N_16270);
nor U17186 (N_17186,N_16612,N_16755);
or U17187 (N_17187,N_16678,N_16404);
nand U17188 (N_17188,N_16439,N_16588);
xor U17189 (N_17189,N_16797,N_16585);
xor U17190 (N_17190,N_16739,N_16659);
or U17191 (N_17191,N_16554,N_16697);
and U17192 (N_17192,N_16513,N_16698);
and U17193 (N_17193,N_16525,N_16437);
xnor U17194 (N_17194,N_16866,N_16411);
nor U17195 (N_17195,N_16281,N_16522);
nand U17196 (N_17196,N_16633,N_16718);
xnor U17197 (N_17197,N_16691,N_16866);
xnor U17198 (N_17198,N_16792,N_16821);
xnor U17199 (N_17199,N_16255,N_16685);
xor U17200 (N_17200,N_16405,N_16660);
nand U17201 (N_17201,N_16486,N_16753);
nor U17202 (N_17202,N_16549,N_16545);
nand U17203 (N_17203,N_16807,N_16856);
or U17204 (N_17204,N_16490,N_16621);
or U17205 (N_17205,N_16513,N_16768);
and U17206 (N_17206,N_16831,N_16652);
or U17207 (N_17207,N_16722,N_16344);
nor U17208 (N_17208,N_16542,N_16401);
or U17209 (N_17209,N_16463,N_16380);
nand U17210 (N_17210,N_16594,N_16687);
or U17211 (N_17211,N_16689,N_16594);
and U17212 (N_17212,N_16462,N_16456);
or U17213 (N_17213,N_16490,N_16447);
xnor U17214 (N_17214,N_16607,N_16315);
or U17215 (N_17215,N_16339,N_16490);
xor U17216 (N_17216,N_16778,N_16711);
nor U17217 (N_17217,N_16455,N_16847);
or U17218 (N_17218,N_16467,N_16311);
or U17219 (N_17219,N_16774,N_16719);
nor U17220 (N_17220,N_16399,N_16518);
or U17221 (N_17221,N_16462,N_16642);
and U17222 (N_17222,N_16621,N_16730);
nand U17223 (N_17223,N_16748,N_16625);
xor U17224 (N_17224,N_16658,N_16592);
and U17225 (N_17225,N_16632,N_16443);
nand U17226 (N_17226,N_16634,N_16320);
and U17227 (N_17227,N_16571,N_16463);
nand U17228 (N_17228,N_16404,N_16719);
or U17229 (N_17229,N_16800,N_16540);
nand U17230 (N_17230,N_16254,N_16530);
nand U17231 (N_17231,N_16603,N_16810);
nor U17232 (N_17232,N_16334,N_16314);
nand U17233 (N_17233,N_16472,N_16578);
nor U17234 (N_17234,N_16610,N_16864);
and U17235 (N_17235,N_16657,N_16622);
or U17236 (N_17236,N_16842,N_16370);
and U17237 (N_17237,N_16533,N_16305);
and U17238 (N_17238,N_16342,N_16831);
nand U17239 (N_17239,N_16665,N_16330);
nand U17240 (N_17240,N_16378,N_16350);
and U17241 (N_17241,N_16616,N_16444);
nor U17242 (N_17242,N_16441,N_16781);
nor U17243 (N_17243,N_16783,N_16521);
nand U17244 (N_17244,N_16841,N_16622);
nor U17245 (N_17245,N_16764,N_16864);
nand U17246 (N_17246,N_16419,N_16465);
or U17247 (N_17247,N_16590,N_16546);
nand U17248 (N_17248,N_16430,N_16313);
and U17249 (N_17249,N_16714,N_16322);
nand U17250 (N_17250,N_16453,N_16372);
nand U17251 (N_17251,N_16826,N_16386);
or U17252 (N_17252,N_16749,N_16488);
nand U17253 (N_17253,N_16447,N_16433);
xnor U17254 (N_17254,N_16376,N_16559);
nor U17255 (N_17255,N_16367,N_16775);
xnor U17256 (N_17256,N_16812,N_16283);
nand U17257 (N_17257,N_16614,N_16701);
nor U17258 (N_17258,N_16252,N_16408);
nand U17259 (N_17259,N_16371,N_16398);
and U17260 (N_17260,N_16850,N_16844);
xor U17261 (N_17261,N_16748,N_16643);
and U17262 (N_17262,N_16838,N_16278);
nand U17263 (N_17263,N_16567,N_16693);
nor U17264 (N_17264,N_16766,N_16562);
nor U17265 (N_17265,N_16614,N_16443);
nand U17266 (N_17266,N_16368,N_16433);
xor U17267 (N_17267,N_16374,N_16485);
nand U17268 (N_17268,N_16316,N_16252);
nor U17269 (N_17269,N_16780,N_16455);
xor U17270 (N_17270,N_16824,N_16343);
nand U17271 (N_17271,N_16677,N_16260);
and U17272 (N_17272,N_16691,N_16380);
xor U17273 (N_17273,N_16851,N_16541);
and U17274 (N_17274,N_16527,N_16804);
nand U17275 (N_17275,N_16836,N_16568);
nand U17276 (N_17276,N_16314,N_16648);
xor U17277 (N_17277,N_16637,N_16577);
xnor U17278 (N_17278,N_16784,N_16343);
nand U17279 (N_17279,N_16409,N_16828);
nand U17280 (N_17280,N_16722,N_16325);
or U17281 (N_17281,N_16359,N_16276);
nand U17282 (N_17282,N_16487,N_16520);
or U17283 (N_17283,N_16786,N_16702);
xnor U17284 (N_17284,N_16576,N_16846);
nand U17285 (N_17285,N_16400,N_16655);
xor U17286 (N_17286,N_16390,N_16473);
nor U17287 (N_17287,N_16285,N_16770);
xor U17288 (N_17288,N_16356,N_16646);
and U17289 (N_17289,N_16615,N_16760);
nand U17290 (N_17290,N_16336,N_16256);
xor U17291 (N_17291,N_16631,N_16291);
nor U17292 (N_17292,N_16256,N_16407);
nand U17293 (N_17293,N_16707,N_16752);
and U17294 (N_17294,N_16705,N_16255);
nand U17295 (N_17295,N_16372,N_16545);
nand U17296 (N_17296,N_16290,N_16623);
nand U17297 (N_17297,N_16463,N_16526);
and U17298 (N_17298,N_16316,N_16369);
nand U17299 (N_17299,N_16412,N_16687);
or U17300 (N_17300,N_16617,N_16431);
nor U17301 (N_17301,N_16468,N_16848);
and U17302 (N_17302,N_16450,N_16780);
xor U17303 (N_17303,N_16262,N_16830);
and U17304 (N_17304,N_16798,N_16863);
xnor U17305 (N_17305,N_16503,N_16696);
or U17306 (N_17306,N_16798,N_16825);
nor U17307 (N_17307,N_16315,N_16748);
nor U17308 (N_17308,N_16339,N_16850);
or U17309 (N_17309,N_16402,N_16461);
nor U17310 (N_17310,N_16512,N_16491);
nand U17311 (N_17311,N_16437,N_16871);
and U17312 (N_17312,N_16303,N_16396);
or U17313 (N_17313,N_16613,N_16859);
and U17314 (N_17314,N_16645,N_16459);
or U17315 (N_17315,N_16307,N_16800);
and U17316 (N_17316,N_16401,N_16869);
nand U17317 (N_17317,N_16476,N_16438);
nor U17318 (N_17318,N_16774,N_16854);
nor U17319 (N_17319,N_16726,N_16286);
nor U17320 (N_17320,N_16384,N_16547);
nand U17321 (N_17321,N_16756,N_16458);
and U17322 (N_17322,N_16583,N_16842);
xnor U17323 (N_17323,N_16792,N_16434);
nor U17324 (N_17324,N_16750,N_16564);
xor U17325 (N_17325,N_16642,N_16553);
nand U17326 (N_17326,N_16739,N_16717);
nor U17327 (N_17327,N_16703,N_16808);
nand U17328 (N_17328,N_16525,N_16564);
and U17329 (N_17329,N_16647,N_16439);
and U17330 (N_17330,N_16511,N_16322);
nor U17331 (N_17331,N_16724,N_16286);
nor U17332 (N_17332,N_16432,N_16508);
xnor U17333 (N_17333,N_16723,N_16479);
xnor U17334 (N_17334,N_16415,N_16262);
xor U17335 (N_17335,N_16295,N_16797);
or U17336 (N_17336,N_16447,N_16475);
and U17337 (N_17337,N_16535,N_16385);
xor U17338 (N_17338,N_16281,N_16653);
nor U17339 (N_17339,N_16295,N_16572);
xnor U17340 (N_17340,N_16585,N_16293);
and U17341 (N_17341,N_16570,N_16489);
nand U17342 (N_17342,N_16288,N_16269);
and U17343 (N_17343,N_16769,N_16258);
xnor U17344 (N_17344,N_16688,N_16837);
and U17345 (N_17345,N_16721,N_16633);
or U17346 (N_17346,N_16653,N_16492);
xor U17347 (N_17347,N_16765,N_16869);
or U17348 (N_17348,N_16573,N_16572);
and U17349 (N_17349,N_16612,N_16592);
and U17350 (N_17350,N_16375,N_16358);
nor U17351 (N_17351,N_16828,N_16499);
or U17352 (N_17352,N_16690,N_16273);
nor U17353 (N_17353,N_16356,N_16765);
xnor U17354 (N_17354,N_16406,N_16251);
nor U17355 (N_17355,N_16252,N_16445);
xor U17356 (N_17356,N_16564,N_16575);
nand U17357 (N_17357,N_16664,N_16765);
nor U17358 (N_17358,N_16420,N_16259);
or U17359 (N_17359,N_16868,N_16586);
nand U17360 (N_17360,N_16760,N_16414);
xor U17361 (N_17361,N_16470,N_16866);
and U17362 (N_17362,N_16687,N_16737);
nor U17363 (N_17363,N_16264,N_16498);
nand U17364 (N_17364,N_16674,N_16394);
and U17365 (N_17365,N_16271,N_16747);
nor U17366 (N_17366,N_16510,N_16273);
xor U17367 (N_17367,N_16531,N_16752);
and U17368 (N_17368,N_16812,N_16862);
nand U17369 (N_17369,N_16597,N_16347);
or U17370 (N_17370,N_16631,N_16524);
nor U17371 (N_17371,N_16772,N_16680);
nor U17372 (N_17372,N_16765,N_16393);
and U17373 (N_17373,N_16352,N_16458);
nand U17374 (N_17374,N_16304,N_16591);
or U17375 (N_17375,N_16785,N_16573);
xnor U17376 (N_17376,N_16476,N_16819);
xnor U17377 (N_17377,N_16558,N_16419);
or U17378 (N_17378,N_16631,N_16310);
nand U17379 (N_17379,N_16818,N_16569);
nor U17380 (N_17380,N_16533,N_16513);
xnor U17381 (N_17381,N_16520,N_16644);
nor U17382 (N_17382,N_16578,N_16400);
nand U17383 (N_17383,N_16847,N_16364);
nand U17384 (N_17384,N_16519,N_16820);
xnor U17385 (N_17385,N_16430,N_16615);
or U17386 (N_17386,N_16449,N_16696);
nor U17387 (N_17387,N_16352,N_16774);
or U17388 (N_17388,N_16435,N_16379);
nor U17389 (N_17389,N_16699,N_16271);
nor U17390 (N_17390,N_16408,N_16405);
or U17391 (N_17391,N_16508,N_16568);
or U17392 (N_17392,N_16532,N_16558);
or U17393 (N_17393,N_16633,N_16553);
xor U17394 (N_17394,N_16442,N_16355);
nand U17395 (N_17395,N_16317,N_16516);
nand U17396 (N_17396,N_16777,N_16519);
and U17397 (N_17397,N_16250,N_16328);
nand U17398 (N_17398,N_16400,N_16663);
xnor U17399 (N_17399,N_16414,N_16726);
nor U17400 (N_17400,N_16636,N_16351);
and U17401 (N_17401,N_16790,N_16328);
and U17402 (N_17402,N_16466,N_16804);
nand U17403 (N_17403,N_16635,N_16292);
and U17404 (N_17404,N_16510,N_16386);
nor U17405 (N_17405,N_16672,N_16754);
or U17406 (N_17406,N_16805,N_16724);
or U17407 (N_17407,N_16846,N_16267);
xnor U17408 (N_17408,N_16598,N_16426);
and U17409 (N_17409,N_16376,N_16617);
and U17410 (N_17410,N_16619,N_16874);
nand U17411 (N_17411,N_16464,N_16582);
and U17412 (N_17412,N_16258,N_16314);
xor U17413 (N_17413,N_16821,N_16596);
nor U17414 (N_17414,N_16548,N_16359);
nand U17415 (N_17415,N_16696,N_16779);
nand U17416 (N_17416,N_16281,N_16766);
xnor U17417 (N_17417,N_16396,N_16405);
nand U17418 (N_17418,N_16420,N_16637);
xor U17419 (N_17419,N_16591,N_16743);
and U17420 (N_17420,N_16341,N_16303);
or U17421 (N_17421,N_16443,N_16645);
xor U17422 (N_17422,N_16670,N_16783);
and U17423 (N_17423,N_16344,N_16620);
and U17424 (N_17424,N_16831,N_16625);
nor U17425 (N_17425,N_16525,N_16490);
or U17426 (N_17426,N_16252,N_16507);
nand U17427 (N_17427,N_16719,N_16694);
nand U17428 (N_17428,N_16359,N_16305);
nand U17429 (N_17429,N_16484,N_16258);
nor U17430 (N_17430,N_16482,N_16490);
nand U17431 (N_17431,N_16410,N_16372);
xnor U17432 (N_17432,N_16368,N_16639);
xnor U17433 (N_17433,N_16853,N_16752);
nand U17434 (N_17434,N_16345,N_16751);
nor U17435 (N_17435,N_16413,N_16865);
xor U17436 (N_17436,N_16867,N_16649);
and U17437 (N_17437,N_16280,N_16725);
and U17438 (N_17438,N_16783,N_16448);
nand U17439 (N_17439,N_16688,N_16470);
xor U17440 (N_17440,N_16819,N_16294);
xor U17441 (N_17441,N_16861,N_16399);
and U17442 (N_17442,N_16316,N_16370);
xnor U17443 (N_17443,N_16405,N_16767);
nor U17444 (N_17444,N_16413,N_16520);
xnor U17445 (N_17445,N_16735,N_16862);
nand U17446 (N_17446,N_16713,N_16418);
nor U17447 (N_17447,N_16799,N_16488);
and U17448 (N_17448,N_16417,N_16450);
or U17449 (N_17449,N_16399,N_16279);
nand U17450 (N_17450,N_16578,N_16821);
or U17451 (N_17451,N_16630,N_16771);
xor U17452 (N_17452,N_16724,N_16638);
and U17453 (N_17453,N_16845,N_16727);
xor U17454 (N_17454,N_16873,N_16312);
or U17455 (N_17455,N_16428,N_16322);
or U17456 (N_17456,N_16780,N_16578);
nor U17457 (N_17457,N_16723,N_16415);
xnor U17458 (N_17458,N_16766,N_16627);
or U17459 (N_17459,N_16751,N_16333);
nand U17460 (N_17460,N_16801,N_16813);
nand U17461 (N_17461,N_16870,N_16670);
nand U17462 (N_17462,N_16596,N_16383);
nor U17463 (N_17463,N_16407,N_16312);
nand U17464 (N_17464,N_16766,N_16414);
xor U17465 (N_17465,N_16597,N_16296);
or U17466 (N_17466,N_16383,N_16550);
xor U17467 (N_17467,N_16752,N_16508);
nand U17468 (N_17468,N_16479,N_16506);
nor U17469 (N_17469,N_16687,N_16378);
or U17470 (N_17470,N_16667,N_16654);
xnor U17471 (N_17471,N_16262,N_16407);
nor U17472 (N_17472,N_16321,N_16265);
and U17473 (N_17473,N_16580,N_16589);
nor U17474 (N_17474,N_16324,N_16759);
xor U17475 (N_17475,N_16422,N_16504);
nand U17476 (N_17476,N_16731,N_16672);
and U17477 (N_17477,N_16461,N_16775);
nand U17478 (N_17478,N_16358,N_16820);
and U17479 (N_17479,N_16284,N_16743);
and U17480 (N_17480,N_16420,N_16275);
and U17481 (N_17481,N_16584,N_16541);
and U17482 (N_17482,N_16766,N_16665);
nand U17483 (N_17483,N_16822,N_16797);
nor U17484 (N_17484,N_16529,N_16634);
nand U17485 (N_17485,N_16269,N_16444);
nand U17486 (N_17486,N_16772,N_16595);
and U17487 (N_17487,N_16398,N_16334);
and U17488 (N_17488,N_16806,N_16632);
nand U17489 (N_17489,N_16750,N_16771);
or U17490 (N_17490,N_16342,N_16722);
and U17491 (N_17491,N_16309,N_16737);
nor U17492 (N_17492,N_16429,N_16335);
nor U17493 (N_17493,N_16547,N_16620);
and U17494 (N_17494,N_16409,N_16817);
or U17495 (N_17495,N_16492,N_16693);
or U17496 (N_17496,N_16400,N_16648);
xor U17497 (N_17497,N_16484,N_16869);
or U17498 (N_17498,N_16443,N_16286);
nor U17499 (N_17499,N_16822,N_16608);
nor U17500 (N_17500,N_17018,N_17100);
or U17501 (N_17501,N_17446,N_16906);
nand U17502 (N_17502,N_16946,N_17229);
xor U17503 (N_17503,N_17287,N_16908);
nor U17504 (N_17504,N_17341,N_17241);
or U17505 (N_17505,N_16943,N_17261);
nand U17506 (N_17506,N_17468,N_17159);
and U17507 (N_17507,N_17364,N_16879);
or U17508 (N_17508,N_16902,N_17211);
nor U17509 (N_17509,N_17431,N_16982);
nand U17510 (N_17510,N_16942,N_17388);
xor U17511 (N_17511,N_17133,N_17228);
nand U17512 (N_17512,N_17420,N_17437);
nand U17513 (N_17513,N_16952,N_17371);
nor U17514 (N_17514,N_17224,N_17423);
nand U17515 (N_17515,N_16905,N_17308);
or U17516 (N_17516,N_17422,N_17059);
or U17517 (N_17517,N_17315,N_17326);
and U17518 (N_17518,N_16989,N_17263);
and U17519 (N_17519,N_17328,N_17413);
xnor U17520 (N_17520,N_16993,N_17017);
or U17521 (N_17521,N_17398,N_17268);
xnor U17522 (N_17522,N_17343,N_17373);
nor U17523 (N_17523,N_17362,N_17390);
or U17524 (N_17524,N_17406,N_16975);
or U17525 (N_17525,N_17411,N_16901);
xor U17526 (N_17526,N_17173,N_16882);
or U17527 (N_17527,N_16983,N_17276);
and U17528 (N_17528,N_17027,N_16985);
nand U17529 (N_17529,N_17128,N_17238);
or U17530 (N_17530,N_17160,N_17144);
xor U17531 (N_17531,N_17424,N_17338);
nand U17532 (N_17532,N_17119,N_17322);
xor U17533 (N_17533,N_17472,N_17037);
xnor U17534 (N_17534,N_17029,N_17384);
and U17535 (N_17535,N_17008,N_16962);
or U17536 (N_17536,N_17028,N_16877);
nand U17537 (N_17537,N_17433,N_17108);
xnor U17538 (N_17538,N_17414,N_17093);
and U17539 (N_17539,N_16964,N_16998);
or U17540 (N_17540,N_16984,N_17488);
xnor U17541 (N_17541,N_16893,N_17340);
and U17542 (N_17542,N_17215,N_17400);
and U17543 (N_17543,N_17448,N_17049);
nand U17544 (N_17544,N_17044,N_17478);
nand U17545 (N_17545,N_17091,N_17382);
and U17546 (N_17546,N_17239,N_16914);
nor U17547 (N_17547,N_17102,N_17447);
or U17548 (N_17548,N_17034,N_17054);
and U17549 (N_17549,N_16947,N_17242);
xor U17550 (N_17550,N_17376,N_17012);
or U17551 (N_17551,N_17244,N_17186);
nor U17552 (N_17552,N_17026,N_16969);
or U17553 (N_17553,N_17112,N_17461);
and U17554 (N_17554,N_17477,N_17097);
xor U17555 (N_17555,N_16996,N_17077);
or U17556 (N_17556,N_17220,N_17252);
nand U17557 (N_17557,N_17115,N_16967);
or U17558 (N_17558,N_16959,N_16890);
xnor U17559 (N_17559,N_17465,N_16940);
xnor U17560 (N_17560,N_17479,N_17493);
nand U17561 (N_17561,N_17174,N_17496);
nor U17562 (N_17562,N_17297,N_17069);
and U17563 (N_17563,N_17061,N_17006);
nand U17564 (N_17564,N_17421,N_17248);
nand U17565 (N_17565,N_16917,N_17455);
or U17566 (N_17566,N_17194,N_17264);
and U17567 (N_17567,N_17419,N_17016);
nor U17568 (N_17568,N_17052,N_17450);
and U17569 (N_17569,N_16912,N_17440);
nand U17570 (N_17570,N_17314,N_17349);
and U17571 (N_17571,N_16892,N_17139);
and U17572 (N_17572,N_16885,N_17272);
nand U17573 (N_17573,N_17429,N_16925);
nor U17574 (N_17574,N_17157,N_17381);
nor U17575 (N_17575,N_17356,N_17039);
xnor U17576 (N_17576,N_17366,N_16972);
nor U17577 (N_17577,N_17149,N_17432);
xor U17578 (N_17578,N_17222,N_17363);
and U17579 (N_17579,N_16971,N_17348);
nand U17580 (N_17580,N_17439,N_17487);
nand U17581 (N_17581,N_16979,N_17323);
or U17582 (N_17582,N_17058,N_17076);
nor U17583 (N_17583,N_17023,N_17473);
nand U17584 (N_17584,N_17416,N_17481);
and U17585 (N_17585,N_16988,N_16981);
xor U17586 (N_17586,N_17292,N_17075);
or U17587 (N_17587,N_17378,N_16991);
nor U17588 (N_17588,N_17060,N_17218);
nand U17589 (N_17589,N_16995,N_17131);
nand U17590 (N_17590,N_17457,N_17010);
nand U17591 (N_17591,N_17168,N_17275);
or U17592 (N_17592,N_17435,N_17083);
and U17593 (N_17593,N_17466,N_17281);
or U17594 (N_17594,N_16965,N_16910);
xnor U17595 (N_17595,N_17310,N_17033);
and U17596 (N_17596,N_17360,N_17246);
xnor U17597 (N_17597,N_17035,N_17143);
nor U17598 (N_17598,N_17367,N_16907);
nor U17599 (N_17599,N_17274,N_17452);
nand U17600 (N_17600,N_17085,N_17000);
xor U17601 (N_17601,N_17068,N_17319);
and U17602 (N_17602,N_17155,N_17464);
or U17603 (N_17603,N_17182,N_17205);
nor U17604 (N_17604,N_17480,N_17277);
or U17605 (N_17605,N_17257,N_17383);
xnor U17606 (N_17606,N_17483,N_17165);
or U17607 (N_17607,N_17207,N_17024);
or U17608 (N_17608,N_17270,N_17247);
nor U17609 (N_17609,N_17453,N_17331);
or U17610 (N_17610,N_17495,N_17064);
nand U17611 (N_17611,N_17237,N_17395);
xor U17612 (N_17612,N_17436,N_16957);
or U17613 (N_17613,N_17219,N_17041);
nor U17614 (N_17614,N_17369,N_17084);
nand U17615 (N_17615,N_17232,N_17181);
and U17616 (N_17616,N_17154,N_17193);
xor U17617 (N_17617,N_17305,N_17072);
nand U17618 (N_17618,N_16909,N_16898);
and U17619 (N_17619,N_17409,N_17463);
or U17620 (N_17620,N_17408,N_17405);
or U17621 (N_17621,N_17407,N_17474);
xnor U17622 (N_17622,N_17088,N_17210);
nor U17623 (N_17623,N_17001,N_17444);
xor U17624 (N_17624,N_17226,N_16896);
and U17625 (N_17625,N_17467,N_16935);
and U17626 (N_17626,N_17183,N_17179);
nand U17627 (N_17627,N_16973,N_17166);
xnor U17628 (N_17628,N_17005,N_17354);
nor U17629 (N_17629,N_17476,N_17158);
nor U17630 (N_17630,N_16949,N_17333);
nor U17631 (N_17631,N_17404,N_17445);
nor U17632 (N_17632,N_16970,N_17329);
nand U17633 (N_17633,N_17372,N_17336);
and U17634 (N_17634,N_17081,N_17002);
xnor U17635 (N_17635,N_17047,N_16963);
or U17636 (N_17636,N_17428,N_17441);
and U17637 (N_17637,N_16924,N_17073);
xnor U17638 (N_17638,N_17200,N_17212);
or U17639 (N_17639,N_17148,N_16883);
nor U17640 (N_17640,N_16980,N_17104);
nand U17641 (N_17641,N_17126,N_17391);
or U17642 (N_17642,N_16976,N_17282);
nand U17643 (N_17643,N_17462,N_17202);
and U17644 (N_17644,N_17418,N_17361);
and U17645 (N_17645,N_17350,N_17386);
or U17646 (N_17646,N_16968,N_17278);
and U17647 (N_17647,N_17048,N_17351);
xor U17648 (N_17648,N_16930,N_17399);
nor U17649 (N_17649,N_17055,N_17080);
or U17650 (N_17650,N_16931,N_17046);
and U17651 (N_17651,N_17298,N_16961);
xnor U17652 (N_17652,N_17011,N_17199);
xor U17653 (N_17653,N_17291,N_17164);
nor U17654 (N_17654,N_17067,N_17417);
or U17655 (N_17655,N_17306,N_17389);
xnor U17656 (N_17656,N_17095,N_17203);
nor U17657 (N_17657,N_16903,N_17189);
xnor U17658 (N_17658,N_16916,N_17188);
and U17659 (N_17659,N_17225,N_17260);
or U17660 (N_17660,N_17216,N_16951);
xor U17661 (N_17661,N_17051,N_16977);
xor U17662 (N_17662,N_17116,N_17107);
nand U17663 (N_17663,N_17254,N_16894);
and U17664 (N_17664,N_17290,N_16876);
or U17665 (N_17665,N_17233,N_17053);
xnor U17666 (N_17666,N_17153,N_17176);
and U17667 (N_17667,N_17134,N_17063);
or U17668 (N_17668,N_16919,N_17151);
nor U17669 (N_17669,N_17482,N_17357);
or U17670 (N_17670,N_17138,N_16881);
nor U17671 (N_17671,N_17316,N_17070);
and U17672 (N_17672,N_17125,N_17043);
xnor U17673 (N_17673,N_17230,N_17007);
xnor U17674 (N_17674,N_17489,N_16978);
or U17675 (N_17675,N_17271,N_17004);
xnor U17676 (N_17676,N_16904,N_17427);
or U17677 (N_17677,N_17380,N_16929);
xnor U17678 (N_17678,N_17377,N_17206);
and U17679 (N_17679,N_16880,N_17294);
and U17680 (N_17680,N_17344,N_17358);
and U17681 (N_17681,N_17201,N_17103);
and U17682 (N_17682,N_17045,N_17300);
xnor U17683 (N_17683,N_17145,N_17096);
nor U17684 (N_17684,N_17339,N_16927);
xor U17685 (N_17685,N_17471,N_17147);
or U17686 (N_17686,N_17332,N_16887);
xor U17687 (N_17687,N_17375,N_17460);
nand U17688 (N_17688,N_17137,N_17335);
or U17689 (N_17689,N_17256,N_17130);
or U17690 (N_17690,N_17296,N_17370);
and U17691 (N_17691,N_17135,N_17318);
xnor U17692 (N_17692,N_17236,N_17280);
and U17693 (N_17693,N_17227,N_17498);
nor U17694 (N_17694,N_17255,N_16948);
xor U17695 (N_17695,N_17123,N_17243);
or U17696 (N_17696,N_16937,N_17013);
nand U17697 (N_17697,N_17180,N_17214);
nor U17698 (N_17698,N_17410,N_17056);
xor U17699 (N_17699,N_17114,N_16997);
nand U17700 (N_17700,N_17320,N_16958);
nor U17701 (N_17701,N_17221,N_17295);
xnor U17702 (N_17702,N_17387,N_17451);
or U17703 (N_17703,N_17346,N_16918);
xnor U17704 (N_17704,N_17491,N_16923);
nor U17705 (N_17705,N_16934,N_17197);
or U17706 (N_17706,N_17022,N_16891);
or U17707 (N_17707,N_17309,N_17334);
nor U17708 (N_17708,N_17265,N_16913);
nor U17709 (N_17709,N_16889,N_17454);
and U17710 (N_17710,N_16932,N_17089);
nor U17711 (N_17711,N_17449,N_16878);
or U17712 (N_17712,N_16920,N_17311);
nand U17713 (N_17713,N_17190,N_17122);
xnor U17714 (N_17714,N_16884,N_17124);
and U17715 (N_17715,N_17178,N_16895);
nand U17716 (N_17716,N_17312,N_16994);
nor U17717 (N_17717,N_16953,N_16922);
nand U17718 (N_17718,N_17267,N_17142);
and U17719 (N_17719,N_17121,N_17438);
nand U17720 (N_17720,N_17032,N_17065);
and U17721 (N_17721,N_17099,N_17019);
and U17722 (N_17722,N_17394,N_17385);
nor U17723 (N_17723,N_17111,N_17110);
xor U17724 (N_17724,N_17475,N_17066);
nand U17725 (N_17725,N_17393,N_17402);
xor U17726 (N_17726,N_16875,N_17175);
xor U17727 (N_17727,N_17499,N_17020);
xor U17728 (N_17728,N_16954,N_17177);
or U17729 (N_17729,N_17266,N_16936);
nand U17730 (N_17730,N_17038,N_16897);
nand U17731 (N_17731,N_16933,N_16974);
or U17732 (N_17732,N_17379,N_17208);
xnor U17733 (N_17733,N_17458,N_17425);
nand U17734 (N_17734,N_17141,N_17184);
or U17735 (N_17735,N_17485,N_17231);
xor U17736 (N_17736,N_17434,N_17325);
or U17737 (N_17737,N_17250,N_17187);
or U17738 (N_17738,N_17127,N_16986);
nand U17739 (N_17739,N_17279,N_17087);
nand U17740 (N_17740,N_16941,N_17223);
xnor U17741 (N_17741,N_16928,N_17259);
or U17742 (N_17742,N_17162,N_17025);
nand U17743 (N_17743,N_16886,N_17330);
nor U17744 (N_17744,N_17050,N_17430);
and U17745 (N_17745,N_16960,N_17082);
nor U17746 (N_17746,N_16990,N_17490);
or U17747 (N_17747,N_17120,N_17217);
or U17748 (N_17748,N_16899,N_17106);
or U17749 (N_17749,N_17302,N_17273);
nor U17750 (N_17750,N_17003,N_17426);
nor U17751 (N_17751,N_17021,N_16999);
and U17752 (N_17752,N_17307,N_17062);
xnor U17753 (N_17753,N_16921,N_17132);
and U17754 (N_17754,N_16911,N_17342);
and U17755 (N_17755,N_17352,N_17078);
and U17756 (N_17756,N_17074,N_17172);
nor U17757 (N_17757,N_17345,N_16945);
nand U17758 (N_17758,N_17031,N_17253);
and U17759 (N_17759,N_17286,N_17057);
or U17760 (N_17760,N_17258,N_17015);
xor U17761 (N_17761,N_17470,N_17359);
nand U17762 (N_17762,N_17185,N_17105);
xor U17763 (N_17763,N_17443,N_17269);
nand U17764 (N_17764,N_17156,N_17484);
nor U17765 (N_17765,N_17456,N_17191);
nor U17766 (N_17766,N_17204,N_16987);
xnor U17767 (N_17767,N_17071,N_17192);
nor U17768 (N_17768,N_17494,N_17152);
and U17769 (N_17769,N_17289,N_17397);
nand U17770 (N_17770,N_17401,N_17396);
nand U17771 (N_17771,N_16900,N_17497);
nand U17772 (N_17772,N_17235,N_17234);
or U17773 (N_17773,N_17304,N_17288);
nand U17774 (N_17774,N_17150,N_17459);
nand U17775 (N_17775,N_17301,N_17392);
nor U17776 (N_17776,N_17140,N_17196);
xor U17777 (N_17777,N_17492,N_17040);
xnor U17778 (N_17778,N_16992,N_17324);
nand U17779 (N_17779,N_16944,N_16938);
nor U17780 (N_17780,N_17347,N_17118);
and U17781 (N_17781,N_17198,N_17365);
xor U17782 (N_17782,N_17213,N_17136);
nand U17783 (N_17783,N_17169,N_17353);
nand U17784 (N_17784,N_17469,N_17412);
xor U17785 (N_17785,N_17313,N_17161);
and U17786 (N_17786,N_17245,N_17368);
nor U17787 (N_17787,N_17337,N_17209);
and U17788 (N_17788,N_17101,N_17030);
or U17789 (N_17789,N_17098,N_16888);
nand U17790 (N_17790,N_16956,N_17283);
nand U17791 (N_17791,N_17170,N_17014);
nor U17792 (N_17792,N_17317,N_17171);
nand U17793 (N_17793,N_17086,N_17284);
nor U17794 (N_17794,N_17090,N_16955);
nor U17795 (N_17795,N_17374,N_17167);
nor U17796 (N_17796,N_17251,N_17009);
xnor U17797 (N_17797,N_17442,N_16915);
nor U17798 (N_17798,N_17240,N_17321);
or U17799 (N_17799,N_17117,N_17094);
or U17800 (N_17800,N_17146,N_16939);
nand U17801 (N_17801,N_17415,N_17109);
nor U17802 (N_17802,N_17163,N_16966);
xnor U17803 (N_17803,N_17299,N_17403);
and U17804 (N_17804,N_17079,N_17195);
nand U17805 (N_17805,N_17293,N_17355);
nand U17806 (N_17806,N_17303,N_17042);
xor U17807 (N_17807,N_17327,N_17285);
or U17808 (N_17808,N_17262,N_17113);
nand U17809 (N_17809,N_17129,N_17249);
or U17810 (N_17810,N_16950,N_17036);
nor U17811 (N_17811,N_16926,N_17092);
xor U17812 (N_17812,N_17486,N_17105);
xnor U17813 (N_17813,N_17387,N_17040);
or U17814 (N_17814,N_17408,N_17009);
and U17815 (N_17815,N_17003,N_17089);
nor U17816 (N_17816,N_17055,N_16985);
nor U17817 (N_17817,N_17210,N_17282);
xnor U17818 (N_17818,N_16891,N_17075);
nor U17819 (N_17819,N_17092,N_16971);
nand U17820 (N_17820,N_17075,N_17065);
nand U17821 (N_17821,N_17072,N_17288);
nand U17822 (N_17822,N_16906,N_17127);
nand U17823 (N_17823,N_17244,N_16969);
xnor U17824 (N_17824,N_17240,N_17218);
xnor U17825 (N_17825,N_17323,N_17462);
nand U17826 (N_17826,N_16909,N_17477);
nor U17827 (N_17827,N_17007,N_17220);
xnor U17828 (N_17828,N_17308,N_17314);
or U17829 (N_17829,N_17415,N_17467);
nor U17830 (N_17830,N_17388,N_17032);
and U17831 (N_17831,N_17288,N_16930);
nand U17832 (N_17832,N_17478,N_17382);
nand U17833 (N_17833,N_17322,N_17228);
nand U17834 (N_17834,N_17247,N_16983);
nand U17835 (N_17835,N_17066,N_17465);
or U17836 (N_17836,N_16950,N_17231);
nor U17837 (N_17837,N_17021,N_17399);
and U17838 (N_17838,N_17105,N_16877);
or U17839 (N_17839,N_17395,N_17430);
xor U17840 (N_17840,N_17340,N_17188);
xnor U17841 (N_17841,N_17235,N_17266);
nor U17842 (N_17842,N_16971,N_17382);
nor U17843 (N_17843,N_17202,N_17313);
nor U17844 (N_17844,N_17265,N_16954);
nor U17845 (N_17845,N_17433,N_17334);
or U17846 (N_17846,N_16992,N_17321);
nand U17847 (N_17847,N_16951,N_17150);
nor U17848 (N_17848,N_17285,N_17228);
xor U17849 (N_17849,N_16911,N_16943);
nor U17850 (N_17850,N_17195,N_17051);
xor U17851 (N_17851,N_17097,N_17348);
nand U17852 (N_17852,N_17027,N_17045);
or U17853 (N_17853,N_17263,N_17253);
and U17854 (N_17854,N_17483,N_17399);
nand U17855 (N_17855,N_17444,N_17439);
nor U17856 (N_17856,N_17232,N_17307);
or U17857 (N_17857,N_17481,N_16953);
or U17858 (N_17858,N_17129,N_17263);
nor U17859 (N_17859,N_17196,N_17006);
and U17860 (N_17860,N_17219,N_17373);
and U17861 (N_17861,N_17126,N_17001);
nand U17862 (N_17862,N_16962,N_17075);
nand U17863 (N_17863,N_17177,N_17123);
and U17864 (N_17864,N_17239,N_17345);
or U17865 (N_17865,N_17078,N_17321);
or U17866 (N_17866,N_17133,N_17219);
nand U17867 (N_17867,N_16931,N_17262);
nor U17868 (N_17868,N_16968,N_17168);
and U17869 (N_17869,N_17068,N_16925);
nor U17870 (N_17870,N_17258,N_17131);
nor U17871 (N_17871,N_17240,N_17227);
and U17872 (N_17872,N_17056,N_17407);
nor U17873 (N_17873,N_17394,N_17179);
xor U17874 (N_17874,N_16895,N_17117);
and U17875 (N_17875,N_17343,N_17079);
nor U17876 (N_17876,N_16931,N_17094);
nor U17877 (N_17877,N_17279,N_17261);
or U17878 (N_17878,N_17338,N_17213);
nand U17879 (N_17879,N_16978,N_17400);
xor U17880 (N_17880,N_17153,N_17243);
xor U17881 (N_17881,N_17000,N_17453);
nor U17882 (N_17882,N_17084,N_17298);
nand U17883 (N_17883,N_17165,N_17403);
and U17884 (N_17884,N_17321,N_17224);
nand U17885 (N_17885,N_17463,N_17275);
and U17886 (N_17886,N_17349,N_17018);
nor U17887 (N_17887,N_16903,N_17195);
nand U17888 (N_17888,N_16940,N_17044);
nor U17889 (N_17889,N_17262,N_16943);
nand U17890 (N_17890,N_17481,N_17143);
or U17891 (N_17891,N_17475,N_17311);
nand U17892 (N_17892,N_17189,N_17298);
and U17893 (N_17893,N_16907,N_17151);
nand U17894 (N_17894,N_16950,N_17298);
nand U17895 (N_17895,N_17100,N_17073);
xor U17896 (N_17896,N_16988,N_16928);
nand U17897 (N_17897,N_17251,N_17265);
xnor U17898 (N_17898,N_16895,N_17104);
nor U17899 (N_17899,N_17393,N_17082);
xnor U17900 (N_17900,N_17426,N_17311);
and U17901 (N_17901,N_17435,N_17145);
and U17902 (N_17902,N_17370,N_17067);
nor U17903 (N_17903,N_17082,N_17039);
nor U17904 (N_17904,N_17384,N_16881);
nand U17905 (N_17905,N_17042,N_17188);
and U17906 (N_17906,N_17044,N_17334);
nor U17907 (N_17907,N_16903,N_17076);
nand U17908 (N_17908,N_16996,N_17084);
xor U17909 (N_17909,N_17435,N_17290);
nor U17910 (N_17910,N_17373,N_17208);
and U17911 (N_17911,N_17483,N_16887);
nand U17912 (N_17912,N_17130,N_17164);
nor U17913 (N_17913,N_17030,N_17473);
xnor U17914 (N_17914,N_17383,N_17482);
nand U17915 (N_17915,N_17049,N_17463);
xnor U17916 (N_17916,N_17108,N_17173);
nor U17917 (N_17917,N_16892,N_17281);
xnor U17918 (N_17918,N_17095,N_17268);
xor U17919 (N_17919,N_17394,N_17333);
nand U17920 (N_17920,N_17343,N_16899);
xor U17921 (N_17921,N_17397,N_17222);
and U17922 (N_17922,N_17051,N_17197);
nor U17923 (N_17923,N_16995,N_17293);
or U17924 (N_17924,N_17428,N_17018);
nor U17925 (N_17925,N_16940,N_17391);
and U17926 (N_17926,N_17022,N_17162);
xor U17927 (N_17927,N_17127,N_17415);
nor U17928 (N_17928,N_17124,N_17059);
nand U17929 (N_17929,N_17432,N_17345);
xor U17930 (N_17930,N_17403,N_17203);
or U17931 (N_17931,N_17048,N_17292);
nand U17932 (N_17932,N_17127,N_17345);
or U17933 (N_17933,N_17400,N_16892);
nand U17934 (N_17934,N_17197,N_17046);
xor U17935 (N_17935,N_17271,N_17373);
nand U17936 (N_17936,N_17091,N_17243);
xor U17937 (N_17937,N_17118,N_17485);
xnor U17938 (N_17938,N_17358,N_17471);
nand U17939 (N_17939,N_17092,N_17400);
nor U17940 (N_17940,N_17264,N_16912);
or U17941 (N_17941,N_17302,N_16875);
nand U17942 (N_17942,N_17095,N_17395);
nand U17943 (N_17943,N_16911,N_17182);
and U17944 (N_17944,N_16994,N_17150);
nor U17945 (N_17945,N_16895,N_17446);
and U17946 (N_17946,N_16945,N_17054);
nand U17947 (N_17947,N_17140,N_17407);
nor U17948 (N_17948,N_17250,N_17120);
nand U17949 (N_17949,N_17339,N_17314);
xor U17950 (N_17950,N_16878,N_17396);
nor U17951 (N_17951,N_17250,N_17145);
or U17952 (N_17952,N_17008,N_17479);
nor U17953 (N_17953,N_17435,N_16932);
or U17954 (N_17954,N_17094,N_17441);
and U17955 (N_17955,N_17165,N_17371);
and U17956 (N_17956,N_17089,N_17133);
nor U17957 (N_17957,N_16892,N_17435);
xnor U17958 (N_17958,N_16953,N_16973);
nor U17959 (N_17959,N_17357,N_17318);
xnor U17960 (N_17960,N_17412,N_17389);
nand U17961 (N_17961,N_16920,N_17475);
or U17962 (N_17962,N_16962,N_17215);
nor U17963 (N_17963,N_16897,N_16914);
xnor U17964 (N_17964,N_17120,N_17400);
nor U17965 (N_17965,N_17288,N_17291);
and U17966 (N_17966,N_17278,N_17045);
nand U17967 (N_17967,N_16883,N_17468);
xor U17968 (N_17968,N_17334,N_17213);
xnor U17969 (N_17969,N_17323,N_16985);
or U17970 (N_17970,N_17124,N_17232);
or U17971 (N_17971,N_17262,N_17036);
nor U17972 (N_17972,N_17069,N_16991);
nand U17973 (N_17973,N_17074,N_17428);
or U17974 (N_17974,N_17451,N_17320);
nor U17975 (N_17975,N_17278,N_17357);
nand U17976 (N_17976,N_17112,N_17240);
or U17977 (N_17977,N_16967,N_17079);
nand U17978 (N_17978,N_17435,N_17220);
xnor U17979 (N_17979,N_17012,N_17322);
nand U17980 (N_17980,N_17340,N_17414);
or U17981 (N_17981,N_17001,N_17244);
xnor U17982 (N_17982,N_17110,N_16941);
or U17983 (N_17983,N_17485,N_17377);
xor U17984 (N_17984,N_17358,N_17469);
nor U17985 (N_17985,N_16895,N_17061);
or U17986 (N_17986,N_17307,N_17114);
nor U17987 (N_17987,N_17254,N_17414);
nor U17988 (N_17988,N_17365,N_17090);
or U17989 (N_17989,N_16966,N_17437);
xnor U17990 (N_17990,N_17238,N_16927);
or U17991 (N_17991,N_17437,N_17336);
or U17992 (N_17992,N_17372,N_17450);
or U17993 (N_17993,N_17251,N_16916);
xor U17994 (N_17994,N_17099,N_17456);
nor U17995 (N_17995,N_17099,N_16965);
and U17996 (N_17996,N_17446,N_16916);
nand U17997 (N_17997,N_17296,N_17126);
and U17998 (N_17998,N_17416,N_17358);
or U17999 (N_17999,N_16969,N_17283);
nor U18000 (N_18000,N_17486,N_17290);
nand U18001 (N_18001,N_17267,N_17177);
nand U18002 (N_18002,N_17462,N_17058);
nor U18003 (N_18003,N_17285,N_17334);
xnor U18004 (N_18004,N_17171,N_17316);
xor U18005 (N_18005,N_17363,N_17498);
or U18006 (N_18006,N_16886,N_17122);
or U18007 (N_18007,N_17487,N_17062);
and U18008 (N_18008,N_17461,N_17153);
xor U18009 (N_18009,N_16890,N_16966);
nor U18010 (N_18010,N_17030,N_17401);
nor U18011 (N_18011,N_16946,N_16981);
nand U18012 (N_18012,N_17402,N_17457);
and U18013 (N_18013,N_16908,N_17278);
and U18014 (N_18014,N_17383,N_17006);
and U18015 (N_18015,N_17429,N_17085);
and U18016 (N_18016,N_16917,N_17081);
nor U18017 (N_18017,N_17343,N_16883);
and U18018 (N_18018,N_17227,N_17444);
xor U18019 (N_18019,N_17485,N_17474);
and U18020 (N_18020,N_17201,N_17434);
nand U18021 (N_18021,N_17204,N_17077);
xnor U18022 (N_18022,N_17132,N_17181);
or U18023 (N_18023,N_17171,N_17023);
nor U18024 (N_18024,N_17200,N_17170);
xor U18025 (N_18025,N_17278,N_16969);
or U18026 (N_18026,N_17137,N_16994);
nand U18027 (N_18027,N_17427,N_17188);
nand U18028 (N_18028,N_17486,N_16961);
and U18029 (N_18029,N_17047,N_17403);
nor U18030 (N_18030,N_17262,N_16897);
and U18031 (N_18031,N_16918,N_17380);
or U18032 (N_18032,N_17313,N_17457);
nor U18033 (N_18033,N_17478,N_17163);
nand U18034 (N_18034,N_17080,N_17109);
or U18035 (N_18035,N_17178,N_17080);
and U18036 (N_18036,N_17417,N_17082);
or U18037 (N_18037,N_17210,N_17310);
nand U18038 (N_18038,N_17277,N_17375);
or U18039 (N_18039,N_17298,N_17249);
nand U18040 (N_18040,N_17274,N_17139);
or U18041 (N_18041,N_17334,N_16942);
or U18042 (N_18042,N_17175,N_17260);
nand U18043 (N_18043,N_17475,N_17033);
and U18044 (N_18044,N_17146,N_16880);
and U18045 (N_18045,N_17222,N_17438);
xor U18046 (N_18046,N_17433,N_17488);
xor U18047 (N_18047,N_17348,N_17397);
xnor U18048 (N_18048,N_17357,N_16911);
and U18049 (N_18049,N_16936,N_17481);
or U18050 (N_18050,N_17194,N_17337);
nand U18051 (N_18051,N_16882,N_17424);
nand U18052 (N_18052,N_16914,N_16993);
and U18053 (N_18053,N_16979,N_17166);
or U18054 (N_18054,N_17408,N_17433);
nand U18055 (N_18055,N_17103,N_16922);
xnor U18056 (N_18056,N_17348,N_17327);
and U18057 (N_18057,N_16958,N_17480);
or U18058 (N_18058,N_17340,N_17364);
or U18059 (N_18059,N_16944,N_16908);
nand U18060 (N_18060,N_17376,N_17205);
nand U18061 (N_18061,N_17091,N_16914);
and U18062 (N_18062,N_17373,N_17194);
nor U18063 (N_18063,N_17234,N_17082);
nand U18064 (N_18064,N_17147,N_17234);
nor U18065 (N_18065,N_17302,N_16893);
and U18066 (N_18066,N_16935,N_17058);
xnor U18067 (N_18067,N_17346,N_16887);
or U18068 (N_18068,N_16875,N_17284);
and U18069 (N_18069,N_17082,N_17236);
xor U18070 (N_18070,N_17212,N_17394);
or U18071 (N_18071,N_17219,N_17182);
or U18072 (N_18072,N_16978,N_17246);
nor U18073 (N_18073,N_17045,N_16991);
nor U18074 (N_18074,N_16969,N_17038);
xnor U18075 (N_18075,N_16960,N_17163);
and U18076 (N_18076,N_17300,N_17400);
xor U18077 (N_18077,N_17469,N_17387);
or U18078 (N_18078,N_17228,N_17386);
and U18079 (N_18079,N_17077,N_17037);
xor U18080 (N_18080,N_17334,N_16952);
and U18081 (N_18081,N_17494,N_17201);
and U18082 (N_18082,N_17003,N_16976);
nand U18083 (N_18083,N_17190,N_17369);
xor U18084 (N_18084,N_17064,N_16985);
nor U18085 (N_18085,N_16954,N_17443);
or U18086 (N_18086,N_17104,N_17316);
and U18087 (N_18087,N_16988,N_17191);
xor U18088 (N_18088,N_17401,N_16923);
nor U18089 (N_18089,N_16996,N_17246);
or U18090 (N_18090,N_17221,N_17263);
or U18091 (N_18091,N_17395,N_16971);
or U18092 (N_18092,N_16974,N_17117);
and U18093 (N_18093,N_17000,N_17297);
nand U18094 (N_18094,N_17331,N_17330);
or U18095 (N_18095,N_17497,N_17415);
xor U18096 (N_18096,N_16892,N_17274);
and U18097 (N_18097,N_16908,N_17093);
xnor U18098 (N_18098,N_17431,N_17133);
or U18099 (N_18099,N_17212,N_17160);
nor U18100 (N_18100,N_16996,N_17286);
and U18101 (N_18101,N_17278,N_17443);
and U18102 (N_18102,N_17096,N_17167);
or U18103 (N_18103,N_16915,N_16950);
xnor U18104 (N_18104,N_17259,N_17403);
or U18105 (N_18105,N_16905,N_17022);
and U18106 (N_18106,N_17368,N_16941);
xor U18107 (N_18107,N_17274,N_17368);
or U18108 (N_18108,N_17130,N_16980);
nor U18109 (N_18109,N_17185,N_17385);
or U18110 (N_18110,N_17477,N_17209);
nand U18111 (N_18111,N_16885,N_17283);
nand U18112 (N_18112,N_17450,N_16955);
nand U18113 (N_18113,N_17241,N_17301);
nor U18114 (N_18114,N_17038,N_17043);
and U18115 (N_18115,N_17429,N_17222);
xnor U18116 (N_18116,N_17092,N_16927);
nor U18117 (N_18117,N_17333,N_17397);
nor U18118 (N_18118,N_17357,N_17149);
or U18119 (N_18119,N_17260,N_17017);
or U18120 (N_18120,N_17389,N_17294);
and U18121 (N_18121,N_17144,N_17468);
nor U18122 (N_18122,N_16992,N_16985);
xor U18123 (N_18123,N_17438,N_16927);
nor U18124 (N_18124,N_17113,N_17076);
and U18125 (N_18125,N_18011,N_18112);
or U18126 (N_18126,N_17707,N_18109);
nor U18127 (N_18127,N_18118,N_17551);
nand U18128 (N_18128,N_17695,N_17878);
and U18129 (N_18129,N_17815,N_18059);
and U18130 (N_18130,N_17563,N_17895);
xor U18131 (N_18131,N_17715,N_18088);
nand U18132 (N_18132,N_17581,N_17961);
or U18133 (N_18133,N_17748,N_17831);
and U18134 (N_18134,N_18123,N_17663);
xor U18135 (N_18135,N_17540,N_17960);
nor U18136 (N_18136,N_17650,N_17717);
xnor U18137 (N_18137,N_18046,N_17951);
or U18138 (N_18138,N_17582,N_17810);
and U18139 (N_18139,N_17891,N_17693);
and U18140 (N_18140,N_17993,N_18095);
xnor U18141 (N_18141,N_17524,N_17728);
nor U18142 (N_18142,N_17845,N_17883);
nand U18143 (N_18143,N_17894,N_17791);
xor U18144 (N_18144,N_17697,N_17839);
xnor U18145 (N_18145,N_17516,N_17900);
or U18146 (N_18146,N_18001,N_17514);
xnor U18147 (N_18147,N_17572,N_17692);
nand U18148 (N_18148,N_17916,N_18013);
or U18149 (N_18149,N_17836,N_17701);
or U18150 (N_18150,N_17566,N_17610);
or U18151 (N_18151,N_17804,N_17884);
nand U18152 (N_18152,N_17953,N_17621);
nor U18153 (N_18153,N_17691,N_17532);
xor U18154 (N_18154,N_18116,N_17962);
xnor U18155 (N_18155,N_18077,N_18022);
nor U18156 (N_18156,N_17988,N_17665);
and U18157 (N_18157,N_17746,N_17786);
nor U18158 (N_18158,N_18043,N_17575);
or U18159 (N_18159,N_17535,N_18039);
and U18160 (N_18160,N_18049,N_17772);
and U18161 (N_18161,N_18082,N_17764);
and U18162 (N_18162,N_17600,N_18093);
nand U18163 (N_18163,N_17569,N_17817);
nand U18164 (N_18164,N_17677,N_18094);
or U18165 (N_18165,N_17596,N_17879);
nand U18166 (N_18166,N_17999,N_17979);
nand U18167 (N_18167,N_17741,N_17943);
or U18168 (N_18168,N_17763,N_18075);
or U18169 (N_18169,N_17808,N_17777);
or U18170 (N_18170,N_17866,N_18072);
xor U18171 (N_18171,N_18068,N_17842);
and U18172 (N_18172,N_18021,N_17548);
nand U18173 (N_18173,N_17814,N_17787);
xnor U18174 (N_18174,N_17850,N_17513);
nor U18175 (N_18175,N_17576,N_18105);
xnor U18176 (N_18176,N_17699,N_17694);
nand U18177 (N_18177,N_17729,N_18019);
and U18178 (N_18178,N_17966,N_17552);
xor U18179 (N_18179,N_17826,N_17615);
nor U18180 (N_18180,N_17867,N_18106);
nor U18181 (N_18181,N_17843,N_18121);
nand U18182 (N_18182,N_18099,N_17529);
nand U18183 (N_18183,N_17543,N_17823);
xor U18184 (N_18184,N_17958,N_17747);
nand U18185 (N_18185,N_17507,N_17557);
xnor U18186 (N_18186,N_18074,N_18045);
nor U18187 (N_18187,N_18030,N_17664);
nor U18188 (N_18188,N_17509,N_17944);
nand U18189 (N_18189,N_17604,N_17775);
or U18190 (N_18190,N_17760,N_17758);
and U18191 (N_18191,N_17969,N_18108);
or U18192 (N_18192,N_17964,N_17683);
and U18193 (N_18193,N_18124,N_17649);
nor U18194 (N_18194,N_18101,N_17530);
xnor U18195 (N_18195,N_17825,N_17835);
xor U18196 (N_18196,N_17594,N_17911);
nand U18197 (N_18197,N_17636,N_17934);
xnor U18198 (N_18198,N_17611,N_17505);
xor U18199 (N_18199,N_18023,N_17788);
nand U18200 (N_18200,N_17635,N_17613);
nand U18201 (N_18201,N_17560,N_17721);
nand U18202 (N_18202,N_17802,N_17720);
xnor U18203 (N_18203,N_17639,N_17725);
nand U18204 (N_18204,N_17501,N_17573);
or U18205 (N_18205,N_17863,N_17619);
xor U18206 (N_18206,N_17726,N_17756);
nor U18207 (N_18207,N_17738,N_18009);
or U18208 (N_18208,N_18063,N_17698);
and U18209 (N_18209,N_17869,N_17813);
xnor U18210 (N_18210,N_17938,N_17739);
and U18211 (N_18211,N_17660,N_17754);
nor U18212 (N_18212,N_17897,N_17538);
or U18213 (N_18213,N_17812,N_17965);
nor U18214 (N_18214,N_17877,N_17919);
nand U18215 (N_18215,N_18096,N_18110);
xor U18216 (N_18216,N_17983,N_17743);
and U18217 (N_18217,N_17702,N_17651);
nor U18218 (N_18218,N_17861,N_17912);
nand U18219 (N_18219,N_17931,N_17875);
xnor U18220 (N_18220,N_17771,N_17920);
nor U18221 (N_18221,N_17727,N_18026);
and U18222 (N_18222,N_17840,N_17527);
nor U18223 (N_18223,N_17722,N_17918);
nand U18224 (N_18224,N_17544,N_18073);
nor U18225 (N_18225,N_17656,N_17565);
nor U18226 (N_18226,N_17902,N_17984);
xnor U18227 (N_18227,N_17888,N_17941);
or U18228 (N_18228,N_17622,N_17982);
or U18229 (N_18229,N_18065,N_17967);
and U18230 (N_18230,N_17689,N_17704);
and U18231 (N_18231,N_17930,N_17935);
and U18232 (N_18232,N_17640,N_18057);
nor U18233 (N_18233,N_17906,N_17886);
and U18234 (N_18234,N_17686,N_18007);
nor U18235 (N_18235,N_17830,N_17751);
and U18236 (N_18236,N_18107,N_17921);
nand U18237 (N_18237,N_17924,N_18064);
and U18238 (N_18238,N_17968,N_17546);
and U18239 (N_18239,N_17745,N_17898);
nor U18240 (N_18240,N_18056,N_17809);
and U18241 (N_18241,N_17607,N_17506);
nand U18242 (N_18242,N_18047,N_17837);
nand U18243 (N_18243,N_18058,N_17948);
or U18244 (N_18244,N_17956,N_17774);
nor U18245 (N_18245,N_17871,N_17652);
xnor U18246 (N_18246,N_17922,N_18050);
and U18247 (N_18247,N_17688,N_17519);
xor U18248 (N_18248,N_17932,N_18015);
xnor U18249 (N_18249,N_17940,N_17757);
or U18250 (N_18250,N_17868,N_17537);
xor U18251 (N_18251,N_17627,N_17798);
nand U18252 (N_18252,N_17703,N_17954);
xnor U18253 (N_18253,N_17592,N_18041);
nor U18254 (N_18254,N_18115,N_18036);
and U18255 (N_18255,N_18066,N_17986);
nand U18256 (N_18256,N_17997,N_17915);
and U18257 (N_18257,N_17641,N_17862);
or U18258 (N_18258,N_17542,N_17976);
nor U18259 (N_18259,N_17851,N_17890);
nand U18260 (N_18260,N_17668,N_17770);
and U18261 (N_18261,N_17829,N_17602);
or U18262 (N_18262,N_17520,N_17970);
nand U18263 (N_18263,N_18067,N_17925);
and U18264 (N_18264,N_17980,N_18083);
xnor U18265 (N_18265,N_17939,N_17857);
or U18266 (N_18266,N_17515,N_17859);
nand U18267 (N_18267,N_17806,N_18120);
nand U18268 (N_18268,N_17526,N_17833);
nor U18269 (N_18269,N_17882,N_17679);
or U18270 (N_18270,N_17591,N_18025);
nor U18271 (N_18271,N_18003,N_18071);
nand U18272 (N_18272,N_18055,N_17755);
nand U18273 (N_18273,N_18061,N_17750);
xnor U18274 (N_18274,N_18037,N_17657);
or U18275 (N_18275,N_18069,N_17511);
nor U18276 (N_18276,N_17778,N_17603);
and U18277 (N_18277,N_17630,N_17658);
or U18278 (N_18278,N_18018,N_17647);
xnor U18279 (N_18279,N_17709,N_18012);
xor U18280 (N_18280,N_17846,N_18020);
and U18281 (N_18281,N_17854,N_17531);
and U18282 (N_18282,N_18052,N_17723);
nand U18283 (N_18283,N_17852,N_17533);
nand U18284 (N_18284,N_18048,N_17881);
xor U18285 (N_18285,N_17779,N_17669);
xnor U18286 (N_18286,N_17598,N_17644);
or U18287 (N_18287,N_17634,N_17662);
xor U18288 (N_18288,N_17684,N_17579);
and U18289 (N_18289,N_18119,N_17690);
nor U18290 (N_18290,N_17642,N_18122);
and U18291 (N_18291,N_17730,N_17927);
or U18292 (N_18292,N_18070,N_17666);
nor U18293 (N_18293,N_17913,N_18032);
nand U18294 (N_18294,N_18062,N_17625);
xnor U18295 (N_18295,N_17856,N_17549);
nor U18296 (N_18296,N_17670,N_17903);
nor U18297 (N_18297,N_17780,N_17672);
xor U18298 (N_18298,N_17737,N_17752);
xnor U18299 (N_18299,N_17795,N_17847);
and U18300 (N_18300,N_18079,N_17765);
xor U18301 (N_18301,N_17629,N_17525);
xor U18302 (N_18302,N_17517,N_17844);
and U18303 (N_18303,N_18091,N_17637);
nand U18304 (N_18304,N_17929,N_17998);
nand U18305 (N_18305,N_18031,N_17899);
or U18306 (N_18306,N_17908,N_17872);
nor U18307 (N_18307,N_17710,N_17949);
or U18308 (N_18308,N_17567,N_17818);
or U18309 (N_18309,N_17571,N_17586);
and U18310 (N_18310,N_17648,N_18092);
nor U18311 (N_18311,N_17564,N_18006);
nor U18312 (N_18312,N_18060,N_17952);
and U18313 (N_18313,N_17626,N_17901);
nand U18314 (N_18314,N_17676,N_17696);
nor U18315 (N_18315,N_18029,N_18010);
or U18316 (N_18316,N_18104,N_17945);
nand U18317 (N_18317,N_18117,N_17880);
or U18318 (N_18318,N_17711,N_17821);
and U18319 (N_18319,N_17887,N_17974);
or U18320 (N_18320,N_17645,N_18080);
and U18321 (N_18321,N_17820,N_17646);
or U18322 (N_18322,N_17554,N_17536);
or U18323 (N_18323,N_18035,N_17585);
nand U18324 (N_18324,N_17946,N_18017);
or U18325 (N_18325,N_17904,N_17675);
or U18326 (N_18326,N_17767,N_17827);
and U18327 (N_18327,N_17989,N_18097);
xnor U18328 (N_18328,N_17828,N_17589);
or U18329 (N_18329,N_17700,N_17947);
nand U18330 (N_18330,N_17759,N_17528);
and U18331 (N_18331,N_17807,N_17800);
xor U18332 (N_18332,N_17612,N_17678);
xor U18333 (N_18333,N_17601,N_17959);
nor U18334 (N_18334,N_18034,N_17504);
nor U18335 (N_18335,N_17975,N_17973);
nand U18336 (N_18336,N_17936,N_17991);
and U18337 (N_18337,N_18100,N_17796);
xnor U18338 (N_18338,N_17824,N_17628);
xor U18339 (N_18339,N_17855,N_17510);
nand U18340 (N_18340,N_17783,N_18054);
nand U18341 (N_18341,N_18113,N_17803);
nor U18342 (N_18342,N_17500,N_17910);
nand U18343 (N_18343,N_17805,N_17933);
nor U18344 (N_18344,N_17706,N_17508);
nor U18345 (N_18345,N_17896,N_17620);
and U18346 (N_18346,N_17761,N_17950);
xnor U18347 (N_18347,N_17577,N_17914);
and U18348 (N_18348,N_18084,N_17618);
nand U18349 (N_18349,N_17865,N_17718);
nor U18350 (N_18350,N_18040,N_17781);
nor U18351 (N_18351,N_17789,N_17539);
xor U18352 (N_18352,N_17978,N_17905);
nor U18353 (N_18353,N_17990,N_17608);
or U18354 (N_18354,N_17580,N_17981);
and U18355 (N_18355,N_17928,N_17860);
nand U18356 (N_18356,N_17885,N_17794);
nor U18357 (N_18357,N_17957,N_18016);
nor U18358 (N_18358,N_17735,N_17977);
or U18359 (N_18359,N_17588,N_18076);
or U18360 (N_18360,N_17578,N_17864);
nor U18361 (N_18361,N_17558,N_17616);
nor U18362 (N_18362,N_17655,N_17785);
nand U18363 (N_18363,N_17661,N_18078);
or U18364 (N_18364,N_17889,N_17838);
nor U18365 (N_18365,N_17744,N_17992);
nand U18366 (N_18366,N_17768,N_17907);
nand U18367 (N_18367,N_17556,N_17617);
and U18368 (N_18368,N_17955,N_17545);
or U18369 (N_18369,N_17849,N_17503);
xor U18370 (N_18370,N_18051,N_17633);
and U18371 (N_18371,N_17534,N_18114);
or U18372 (N_18372,N_17605,N_17512);
or U18373 (N_18373,N_17874,N_17547);
or U18374 (N_18374,N_17731,N_17832);
and U18375 (N_18375,N_17816,N_17797);
or U18376 (N_18376,N_18004,N_17873);
nor U18377 (N_18377,N_17740,N_18042);
nand U18378 (N_18378,N_17801,N_18033);
xnor U18379 (N_18379,N_17623,N_17631);
xor U18380 (N_18380,N_17659,N_17923);
xnor U18381 (N_18381,N_17521,N_17687);
nand U18382 (N_18382,N_17926,N_17587);
and U18383 (N_18383,N_17773,N_18102);
xor U18384 (N_18384,N_17892,N_17713);
nand U18385 (N_18385,N_17736,N_18005);
or U18386 (N_18386,N_17590,N_17673);
or U18387 (N_18387,N_17766,N_18086);
xnor U18388 (N_18388,N_17985,N_17716);
nor U18389 (N_18389,N_17541,N_18089);
nand U18390 (N_18390,N_17799,N_17681);
or U18391 (N_18391,N_18000,N_18038);
nand U18392 (N_18392,N_17555,N_17712);
and U18393 (N_18393,N_17553,N_17667);
and U18394 (N_18394,N_17599,N_17963);
or U18395 (N_18395,N_17685,N_17559);
or U18396 (N_18396,N_18085,N_17518);
xor U18397 (N_18397,N_17609,N_17732);
and U18398 (N_18398,N_18111,N_17834);
xnor U18399 (N_18399,N_17870,N_17654);
or U18400 (N_18400,N_17822,N_17909);
and U18401 (N_18401,N_18098,N_17742);
or U18402 (N_18402,N_17562,N_18053);
and U18403 (N_18403,N_17972,N_17994);
nand U18404 (N_18404,N_17942,N_17597);
nor U18405 (N_18405,N_17574,N_17853);
or U18406 (N_18406,N_17734,N_17753);
nor U18407 (N_18407,N_17762,N_17776);
xnor U18408 (N_18408,N_17653,N_17584);
nor U18409 (N_18409,N_17550,N_17841);
nand U18410 (N_18410,N_17523,N_17568);
and U18411 (N_18411,N_18081,N_17749);
and U18412 (N_18412,N_17793,N_17583);
nor U18413 (N_18413,N_17561,N_17671);
and U18414 (N_18414,N_17682,N_17593);
xor U18415 (N_18415,N_17782,N_17570);
or U18416 (N_18416,N_17595,N_17792);
nor U18417 (N_18417,N_17917,N_17680);
xor U18418 (N_18418,N_17876,N_17733);
xor U18419 (N_18419,N_17819,N_17606);
or U18420 (N_18420,N_18008,N_17674);
xnor U18421 (N_18421,N_17632,N_17987);
and U18422 (N_18422,N_17893,N_17769);
xnor U18423 (N_18423,N_17708,N_17522);
nor U18424 (N_18424,N_17614,N_17724);
nor U18425 (N_18425,N_18028,N_18087);
nand U18426 (N_18426,N_17848,N_18044);
nand U18427 (N_18427,N_17811,N_17624);
or U18428 (N_18428,N_17858,N_18103);
and U18429 (N_18429,N_18024,N_17790);
or U18430 (N_18430,N_17705,N_17937);
nand U18431 (N_18431,N_17638,N_17502);
nand U18432 (N_18432,N_17971,N_17719);
or U18433 (N_18433,N_18090,N_18002);
and U18434 (N_18434,N_17714,N_17784);
or U18435 (N_18435,N_17643,N_18027);
nand U18436 (N_18436,N_18014,N_17996);
and U18437 (N_18437,N_17995,N_17568);
nor U18438 (N_18438,N_17998,N_17846);
and U18439 (N_18439,N_17789,N_17590);
and U18440 (N_18440,N_17693,N_17908);
and U18441 (N_18441,N_17978,N_17961);
or U18442 (N_18442,N_18121,N_18106);
and U18443 (N_18443,N_17607,N_18022);
nand U18444 (N_18444,N_17723,N_17580);
nor U18445 (N_18445,N_17911,N_18019);
nand U18446 (N_18446,N_17756,N_17838);
xor U18447 (N_18447,N_17875,N_17712);
nand U18448 (N_18448,N_17856,N_17555);
nor U18449 (N_18449,N_17727,N_17504);
or U18450 (N_18450,N_17630,N_17538);
nor U18451 (N_18451,N_17707,N_18081);
nor U18452 (N_18452,N_17556,N_17580);
nand U18453 (N_18453,N_17735,N_17827);
and U18454 (N_18454,N_18034,N_17690);
xnor U18455 (N_18455,N_17880,N_18121);
nor U18456 (N_18456,N_17925,N_17989);
nor U18457 (N_18457,N_17765,N_17783);
and U18458 (N_18458,N_17500,N_17737);
nand U18459 (N_18459,N_17598,N_17652);
and U18460 (N_18460,N_17959,N_17934);
nand U18461 (N_18461,N_17979,N_17719);
and U18462 (N_18462,N_17709,N_17978);
and U18463 (N_18463,N_17714,N_17597);
nand U18464 (N_18464,N_17827,N_17967);
and U18465 (N_18465,N_17597,N_17722);
or U18466 (N_18466,N_17519,N_17578);
nand U18467 (N_18467,N_17560,N_17581);
nor U18468 (N_18468,N_17573,N_17645);
xnor U18469 (N_18469,N_18013,N_17933);
xor U18470 (N_18470,N_17967,N_17668);
and U18471 (N_18471,N_17978,N_18100);
or U18472 (N_18472,N_17565,N_17540);
and U18473 (N_18473,N_18006,N_17843);
nor U18474 (N_18474,N_17815,N_17553);
and U18475 (N_18475,N_17978,N_17963);
xnor U18476 (N_18476,N_17788,N_17805);
or U18477 (N_18477,N_17690,N_18124);
and U18478 (N_18478,N_17607,N_17554);
xor U18479 (N_18479,N_18069,N_18004);
nand U18480 (N_18480,N_17522,N_17786);
and U18481 (N_18481,N_17575,N_18089);
nor U18482 (N_18482,N_18091,N_17997);
and U18483 (N_18483,N_17520,N_17992);
or U18484 (N_18484,N_18111,N_17961);
and U18485 (N_18485,N_17745,N_17868);
or U18486 (N_18486,N_17753,N_17662);
xnor U18487 (N_18487,N_17527,N_17723);
nand U18488 (N_18488,N_17717,N_18062);
nor U18489 (N_18489,N_17961,N_17790);
nand U18490 (N_18490,N_18078,N_17895);
nor U18491 (N_18491,N_17839,N_18007);
xor U18492 (N_18492,N_17957,N_17532);
or U18493 (N_18493,N_17727,N_17992);
nor U18494 (N_18494,N_17636,N_17860);
and U18495 (N_18495,N_17676,N_17551);
nor U18496 (N_18496,N_17620,N_17862);
and U18497 (N_18497,N_18021,N_18081);
nand U18498 (N_18498,N_17676,N_17918);
xor U18499 (N_18499,N_17673,N_17688);
and U18500 (N_18500,N_17636,N_17643);
and U18501 (N_18501,N_17847,N_17740);
nor U18502 (N_18502,N_17624,N_18047);
or U18503 (N_18503,N_17562,N_17651);
nor U18504 (N_18504,N_18000,N_17807);
or U18505 (N_18505,N_17680,N_17949);
nand U18506 (N_18506,N_17670,N_18064);
or U18507 (N_18507,N_17551,N_17856);
or U18508 (N_18508,N_17636,N_17999);
nand U18509 (N_18509,N_17883,N_18044);
and U18510 (N_18510,N_17969,N_17875);
nand U18511 (N_18511,N_17828,N_17729);
or U18512 (N_18512,N_18045,N_18095);
nor U18513 (N_18513,N_17960,N_17927);
and U18514 (N_18514,N_17638,N_17947);
and U18515 (N_18515,N_18045,N_17543);
nor U18516 (N_18516,N_17944,N_18114);
xnor U18517 (N_18517,N_17604,N_17862);
or U18518 (N_18518,N_17557,N_17589);
nand U18519 (N_18519,N_18119,N_17895);
xor U18520 (N_18520,N_17502,N_17775);
and U18521 (N_18521,N_17649,N_17785);
nand U18522 (N_18522,N_17884,N_18021);
and U18523 (N_18523,N_17861,N_17544);
and U18524 (N_18524,N_17979,N_17635);
nand U18525 (N_18525,N_18075,N_17968);
xnor U18526 (N_18526,N_17767,N_17888);
xnor U18527 (N_18527,N_17752,N_18123);
xnor U18528 (N_18528,N_17984,N_17634);
and U18529 (N_18529,N_17985,N_18124);
nand U18530 (N_18530,N_17582,N_17920);
nor U18531 (N_18531,N_18095,N_17729);
and U18532 (N_18532,N_17807,N_18043);
xor U18533 (N_18533,N_18001,N_17526);
xnor U18534 (N_18534,N_17674,N_17527);
nor U18535 (N_18535,N_17847,N_17661);
or U18536 (N_18536,N_17949,N_17601);
or U18537 (N_18537,N_17586,N_17847);
xor U18538 (N_18538,N_17581,N_17645);
or U18539 (N_18539,N_17889,N_18038);
or U18540 (N_18540,N_17547,N_17628);
nand U18541 (N_18541,N_17668,N_18051);
nor U18542 (N_18542,N_17698,N_17732);
xor U18543 (N_18543,N_17834,N_17643);
nor U18544 (N_18544,N_17704,N_18122);
and U18545 (N_18545,N_17558,N_17508);
xnor U18546 (N_18546,N_17841,N_17675);
nor U18547 (N_18547,N_17854,N_18022);
and U18548 (N_18548,N_17883,N_17555);
and U18549 (N_18549,N_18026,N_18021);
nor U18550 (N_18550,N_17982,N_17731);
xor U18551 (N_18551,N_17613,N_17996);
xnor U18552 (N_18552,N_17919,N_17622);
xor U18553 (N_18553,N_17599,N_18123);
nor U18554 (N_18554,N_17926,N_17882);
xnor U18555 (N_18555,N_18035,N_17955);
or U18556 (N_18556,N_18044,N_18078);
nor U18557 (N_18557,N_17508,N_17982);
nor U18558 (N_18558,N_17803,N_17523);
nand U18559 (N_18559,N_17910,N_17573);
or U18560 (N_18560,N_18046,N_17815);
and U18561 (N_18561,N_17900,N_17607);
or U18562 (N_18562,N_17595,N_18082);
nor U18563 (N_18563,N_18004,N_17869);
nand U18564 (N_18564,N_17832,N_17600);
xor U18565 (N_18565,N_17948,N_17956);
nand U18566 (N_18566,N_17830,N_18063);
nand U18567 (N_18567,N_17641,N_17671);
or U18568 (N_18568,N_17658,N_17757);
nand U18569 (N_18569,N_17917,N_17843);
xor U18570 (N_18570,N_17922,N_17606);
nor U18571 (N_18571,N_17797,N_17778);
nand U18572 (N_18572,N_18076,N_18122);
xnor U18573 (N_18573,N_17874,N_17957);
xor U18574 (N_18574,N_17649,N_17851);
and U18575 (N_18575,N_17660,N_17795);
or U18576 (N_18576,N_17914,N_17590);
xnor U18577 (N_18577,N_17813,N_17903);
and U18578 (N_18578,N_17740,N_17706);
nand U18579 (N_18579,N_17674,N_17925);
xnor U18580 (N_18580,N_17864,N_17758);
xnor U18581 (N_18581,N_17772,N_17758);
nor U18582 (N_18582,N_17755,N_17889);
nor U18583 (N_18583,N_17821,N_17542);
xor U18584 (N_18584,N_17946,N_17897);
and U18585 (N_18585,N_17744,N_18051);
xnor U18586 (N_18586,N_18009,N_17903);
xor U18587 (N_18587,N_17681,N_17501);
or U18588 (N_18588,N_17623,N_17830);
nand U18589 (N_18589,N_17645,N_18112);
and U18590 (N_18590,N_17566,N_17616);
or U18591 (N_18591,N_18083,N_18076);
or U18592 (N_18592,N_17625,N_17940);
xor U18593 (N_18593,N_17850,N_18054);
nand U18594 (N_18594,N_17629,N_18065);
and U18595 (N_18595,N_17739,N_17863);
nand U18596 (N_18596,N_17507,N_17758);
or U18597 (N_18597,N_17517,N_17705);
nand U18598 (N_18598,N_18060,N_17971);
or U18599 (N_18599,N_18058,N_17855);
or U18600 (N_18600,N_17508,N_17814);
nor U18601 (N_18601,N_17942,N_17561);
and U18602 (N_18602,N_18078,N_17890);
and U18603 (N_18603,N_18065,N_17595);
xor U18604 (N_18604,N_17891,N_17569);
nor U18605 (N_18605,N_18088,N_17915);
or U18606 (N_18606,N_17537,N_17529);
xnor U18607 (N_18607,N_17949,N_17920);
nand U18608 (N_18608,N_17646,N_17706);
xnor U18609 (N_18609,N_17900,N_17517);
nor U18610 (N_18610,N_17768,N_17561);
and U18611 (N_18611,N_17767,N_17506);
nor U18612 (N_18612,N_17834,N_17912);
xor U18613 (N_18613,N_17853,N_17832);
nor U18614 (N_18614,N_17524,N_17811);
or U18615 (N_18615,N_17682,N_17538);
nor U18616 (N_18616,N_17679,N_17853);
and U18617 (N_18617,N_18085,N_17657);
nor U18618 (N_18618,N_17717,N_17922);
xnor U18619 (N_18619,N_17726,N_17695);
or U18620 (N_18620,N_17534,N_17565);
nor U18621 (N_18621,N_17696,N_17818);
nand U18622 (N_18622,N_18073,N_17841);
nor U18623 (N_18623,N_17899,N_17926);
and U18624 (N_18624,N_17987,N_17559);
nor U18625 (N_18625,N_17724,N_17530);
nor U18626 (N_18626,N_17853,N_17883);
and U18627 (N_18627,N_17811,N_17663);
xnor U18628 (N_18628,N_18116,N_18072);
xnor U18629 (N_18629,N_17834,N_17961);
xor U18630 (N_18630,N_17666,N_17794);
nand U18631 (N_18631,N_18070,N_18004);
nand U18632 (N_18632,N_17842,N_17650);
or U18633 (N_18633,N_17974,N_17509);
xnor U18634 (N_18634,N_17794,N_17772);
and U18635 (N_18635,N_17566,N_17650);
nand U18636 (N_18636,N_18007,N_17628);
or U18637 (N_18637,N_17523,N_17951);
or U18638 (N_18638,N_17682,N_18124);
or U18639 (N_18639,N_18097,N_17969);
nand U18640 (N_18640,N_17708,N_17696);
nor U18641 (N_18641,N_17832,N_17855);
nand U18642 (N_18642,N_17896,N_18045);
nand U18643 (N_18643,N_17862,N_17502);
nand U18644 (N_18644,N_18113,N_17613);
xor U18645 (N_18645,N_17643,N_17536);
xor U18646 (N_18646,N_18077,N_17561);
and U18647 (N_18647,N_18049,N_17728);
nand U18648 (N_18648,N_17515,N_17630);
xnor U18649 (N_18649,N_17818,N_17922);
nand U18650 (N_18650,N_17898,N_17920);
nand U18651 (N_18651,N_17894,N_17589);
or U18652 (N_18652,N_17521,N_18029);
or U18653 (N_18653,N_17641,N_17821);
and U18654 (N_18654,N_18018,N_17778);
or U18655 (N_18655,N_17732,N_17896);
or U18656 (N_18656,N_17903,N_17590);
and U18657 (N_18657,N_17769,N_17882);
nor U18658 (N_18658,N_18092,N_18018);
or U18659 (N_18659,N_17845,N_17864);
nor U18660 (N_18660,N_18061,N_18051);
xor U18661 (N_18661,N_17743,N_17720);
nor U18662 (N_18662,N_18064,N_18098);
nand U18663 (N_18663,N_17639,N_17957);
or U18664 (N_18664,N_17746,N_17906);
or U18665 (N_18665,N_17890,N_17535);
nor U18666 (N_18666,N_17792,N_17628);
or U18667 (N_18667,N_17530,N_17920);
and U18668 (N_18668,N_17912,N_18057);
nor U18669 (N_18669,N_17968,N_17610);
nor U18670 (N_18670,N_17899,N_17873);
xnor U18671 (N_18671,N_17775,N_17841);
or U18672 (N_18672,N_18068,N_17690);
nand U18673 (N_18673,N_17800,N_17863);
nand U18674 (N_18674,N_17926,N_17721);
nand U18675 (N_18675,N_17994,N_17500);
xor U18676 (N_18676,N_17810,N_17970);
nand U18677 (N_18677,N_17792,N_17901);
nand U18678 (N_18678,N_18021,N_17512);
and U18679 (N_18679,N_17729,N_17984);
or U18680 (N_18680,N_17556,N_17872);
or U18681 (N_18681,N_18006,N_17845);
and U18682 (N_18682,N_17572,N_18007);
or U18683 (N_18683,N_17962,N_18048);
and U18684 (N_18684,N_17826,N_18117);
nand U18685 (N_18685,N_17506,N_17574);
nand U18686 (N_18686,N_17766,N_17897);
or U18687 (N_18687,N_17961,N_17887);
and U18688 (N_18688,N_17600,N_17951);
nand U18689 (N_18689,N_17786,N_17902);
nand U18690 (N_18690,N_17613,N_17585);
nor U18691 (N_18691,N_18002,N_17686);
nor U18692 (N_18692,N_17711,N_17749);
xnor U18693 (N_18693,N_17593,N_17776);
xnor U18694 (N_18694,N_17554,N_17636);
nor U18695 (N_18695,N_18098,N_18045);
and U18696 (N_18696,N_17828,N_17619);
or U18697 (N_18697,N_17984,N_17873);
or U18698 (N_18698,N_17754,N_17652);
xnor U18699 (N_18699,N_17959,N_18054);
nand U18700 (N_18700,N_17807,N_17935);
nand U18701 (N_18701,N_17683,N_18119);
and U18702 (N_18702,N_17921,N_17644);
or U18703 (N_18703,N_17768,N_17650);
nor U18704 (N_18704,N_17652,N_17555);
nor U18705 (N_18705,N_17927,N_17972);
or U18706 (N_18706,N_17754,N_17569);
and U18707 (N_18707,N_18065,N_17918);
xor U18708 (N_18708,N_18097,N_17611);
and U18709 (N_18709,N_17604,N_17539);
or U18710 (N_18710,N_17740,N_17970);
nor U18711 (N_18711,N_17571,N_17882);
and U18712 (N_18712,N_17792,N_17878);
nand U18713 (N_18713,N_18044,N_18026);
and U18714 (N_18714,N_17830,N_18050);
nand U18715 (N_18715,N_17745,N_17991);
or U18716 (N_18716,N_17776,N_17574);
nor U18717 (N_18717,N_17710,N_17763);
nand U18718 (N_18718,N_17998,N_17745);
xnor U18719 (N_18719,N_17684,N_17635);
xor U18720 (N_18720,N_17650,N_17725);
nor U18721 (N_18721,N_17753,N_17754);
and U18722 (N_18722,N_18094,N_18014);
xor U18723 (N_18723,N_17806,N_17666);
nor U18724 (N_18724,N_17518,N_17520);
nor U18725 (N_18725,N_18024,N_17689);
or U18726 (N_18726,N_17844,N_17776);
nand U18727 (N_18727,N_17536,N_17925);
or U18728 (N_18728,N_18028,N_18085);
or U18729 (N_18729,N_17810,N_17790);
nor U18730 (N_18730,N_17674,N_17684);
nor U18731 (N_18731,N_17903,N_17615);
xnor U18732 (N_18732,N_17838,N_17975);
nand U18733 (N_18733,N_17665,N_18087);
nand U18734 (N_18734,N_17518,N_17857);
xor U18735 (N_18735,N_17726,N_17755);
and U18736 (N_18736,N_17847,N_17555);
and U18737 (N_18737,N_17987,N_18025);
nand U18738 (N_18738,N_17864,N_17613);
nor U18739 (N_18739,N_17563,N_17984);
and U18740 (N_18740,N_18073,N_17885);
or U18741 (N_18741,N_17865,N_17584);
or U18742 (N_18742,N_17805,N_17895);
and U18743 (N_18743,N_17562,N_17641);
or U18744 (N_18744,N_17792,N_18118);
or U18745 (N_18745,N_17950,N_17863);
nand U18746 (N_18746,N_18007,N_17795);
xor U18747 (N_18747,N_17572,N_18011);
xnor U18748 (N_18748,N_17950,N_17546);
xor U18749 (N_18749,N_17742,N_17568);
nand U18750 (N_18750,N_18218,N_18181);
xnor U18751 (N_18751,N_18205,N_18402);
and U18752 (N_18752,N_18687,N_18485);
and U18753 (N_18753,N_18264,N_18329);
xor U18754 (N_18754,N_18738,N_18158);
nand U18755 (N_18755,N_18502,N_18410);
nor U18756 (N_18756,N_18184,N_18471);
xnor U18757 (N_18757,N_18440,N_18345);
nor U18758 (N_18758,N_18257,N_18373);
and U18759 (N_18759,N_18347,N_18621);
or U18760 (N_18760,N_18454,N_18192);
or U18761 (N_18761,N_18146,N_18693);
nand U18762 (N_18762,N_18625,N_18370);
nor U18763 (N_18763,N_18371,N_18749);
nand U18764 (N_18764,N_18432,N_18281);
or U18765 (N_18765,N_18706,N_18518);
and U18766 (N_18766,N_18219,N_18479);
and U18767 (N_18767,N_18716,N_18187);
nor U18768 (N_18768,N_18611,N_18601);
or U18769 (N_18769,N_18211,N_18666);
nand U18770 (N_18770,N_18407,N_18164);
nand U18771 (N_18771,N_18126,N_18230);
nor U18772 (N_18772,N_18554,N_18378);
or U18773 (N_18773,N_18487,N_18623);
nand U18774 (N_18774,N_18435,N_18640);
nand U18775 (N_18775,N_18536,N_18385);
nand U18776 (N_18776,N_18201,N_18384);
or U18777 (N_18777,N_18542,N_18481);
nand U18778 (N_18778,N_18237,N_18178);
or U18779 (N_18779,N_18221,N_18141);
nor U18780 (N_18780,N_18392,N_18367);
xnor U18781 (N_18781,N_18494,N_18694);
xnor U18782 (N_18782,N_18550,N_18654);
and U18783 (N_18783,N_18317,N_18522);
and U18784 (N_18784,N_18683,N_18579);
nor U18785 (N_18785,N_18697,N_18599);
nand U18786 (N_18786,N_18584,N_18263);
or U18787 (N_18787,N_18353,N_18707);
or U18788 (N_18788,N_18595,N_18498);
nand U18789 (N_18789,N_18583,N_18632);
xor U18790 (N_18790,N_18429,N_18638);
xor U18791 (N_18791,N_18552,N_18288);
nand U18792 (N_18792,N_18280,N_18388);
nor U18793 (N_18793,N_18170,N_18728);
nand U18794 (N_18794,N_18301,N_18658);
xnor U18795 (N_18795,N_18349,N_18127);
nor U18796 (N_18796,N_18566,N_18417);
or U18797 (N_18797,N_18659,N_18437);
and U18798 (N_18798,N_18701,N_18745);
and U18799 (N_18799,N_18719,N_18161);
or U18800 (N_18800,N_18387,N_18334);
and U18801 (N_18801,N_18461,N_18664);
nor U18802 (N_18802,N_18656,N_18634);
nor U18803 (N_18803,N_18294,N_18453);
nor U18804 (N_18804,N_18155,N_18238);
xor U18805 (N_18805,N_18711,N_18403);
and U18806 (N_18806,N_18534,N_18555);
and U18807 (N_18807,N_18355,N_18190);
nand U18808 (N_18808,N_18436,N_18460);
and U18809 (N_18809,N_18273,N_18490);
nor U18810 (N_18810,N_18480,N_18400);
nand U18811 (N_18811,N_18330,N_18635);
nor U18812 (N_18812,N_18596,N_18176);
nand U18813 (N_18813,N_18434,N_18572);
xnor U18814 (N_18814,N_18246,N_18692);
or U18815 (N_18815,N_18136,N_18525);
nand U18816 (N_18816,N_18217,N_18653);
nand U18817 (N_18817,N_18447,N_18445);
and U18818 (N_18818,N_18142,N_18171);
and U18819 (N_18819,N_18382,N_18497);
xor U18820 (N_18820,N_18698,N_18274);
nor U18821 (N_18821,N_18501,N_18468);
xnor U18822 (N_18822,N_18473,N_18215);
nor U18823 (N_18823,N_18277,N_18372);
xnor U18824 (N_18824,N_18303,N_18651);
nand U18825 (N_18825,N_18637,N_18254);
xor U18826 (N_18826,N_18316,N_18450);
and U18827 (N_18827,N_18641,N_18517);
and U18828 (N_18828,N_18358,N_18448);
nor U18829 (N_18829,N_18681,N_18524);
nor U18830 (N_18830,N_18615,N_18655);
and U18831 (N_18831,N_18231,N_18673);
nor U18832 (N_18832,N_18463,N_18185);
nand U18833 (N_18833,N_18132,N_18243);
xnor U18834 (N_18834,N_18495,N_18741);
or U18835 (N_18835,N_18172,N_18269);
nand U18836 (N_18836,N_18203,N_18671);
nor U18837 (N_18837,N_18174,N_18175);
and U18838 (N_18838,N_18343,N_18685);
nand U18839 (N_18839,N_18169,N_18302);
and U18840 (N_18840,N_18527,N_18356);
nand U18841 (N_18841,N_18529,N_18369);
and U18842 (N_18842,N_18742,N_18399);
or U18843 (N_18843,N_18474,N_18475);
or U18844 (N_18844,N_18167,N_18374);
and U18845 (N_18845,N_18259,N_18298);
xor U18846 (N_18846,N_18415,N_18732);
and U18847 (N_18847,N_18558,N_18222);
or U18848 (N_18848,N_18245,N_18228);
or U18849 (N_18849,N_18723,N_18404);
and U18850 (N_18850,N_18156,N_18346);
or U18851 (N_18851,N_18613,N_18359);
nand U18852 (N_18852,N_18188,N_18262);
or U18853 (N_18853,N_18409,N_18278);
nand U18854 (N_18854,N_18260,N_18290);
and U18855 (N_18855,N_18748,N_18418);
or U18856 (N_18856,N_18512,N_18725);
nand U18857 (N_18857,N_18157,N_18179);
nor U18858 (N_18858,N_18325,N_18433);
and U18859 (N_18859,N_18457,N_18602);
nor U18860 (N_18860,N_18730,N_18444);
xor U18861 (N_18861,N_18139,N_18578);
xor U18862 (N_18862,N_18390,N_18150);
nor U18863 (N_18863,N_18248,N_18570);
xor U18864 (N_18864,N_18442,N_18605);
or U18865 (N_18865,N_18668,N_18735);
nand U18866 (N_18866,N_18213,N_18309);
xnor U18867 (N_18867,N_18603,N_18265);
or U18868 (N_18868,N_18267,N_18214);
nor U18869 (N_18869,N_18401,N_18282);
or U18870 (N_18870,N_18168,N_18191);
or U18871 (N_18871,N_18574,N_18670);
nor U18872 (N_18872,N_18530,N_18633);
and U18873 (N_18873,N_18207,N_18478);
and U18874 (N_18874,N_18580,N_18261);
nand U18875 (N_18875,N_18438,N_18675);
nand U18876 (N_18876,N_18331,N_18315);
nor U18877 (N_18877,N_18227,N_18567);
nand U18878 (N_18878,N_18624,N_18297);
or U18879 (N_18879,N_18128,N_18667);
or U18880 (N_18880,N_18287,N_18573);
nand U18881 (N_18881,N_18408,N_18339);
nand U18882 (N_18882,N_18272,N_18590);
nand U18883 (N_18883,N_18166,N_18712);
and U18884 (N_18884,N_18587,N_18456);
nor U18885 (N_18885,N_18266,N_18352);
nand U18886 (N_18886,N_18476,N_18513);
xnor U18887 (N_18887,N_18398,N_18559);
xnor U18888 (N_18888,N_18342,N_18690);
xnor U18889 (N_18889,N_18295,N_18427);
nand U18890 (N_18890,N_18677,N_18616);
or U18891 (N_18891,N_18720,N_18341);
xnor U18892 (N_18892,N_18628,N_18413);
nand U18893 (N_18893,N_18710,N_18242);
xnor U18894 (N_18894,N_18650,N_18240);
xor U18895 (N_18895,N_18321,N_18380);
nor U18896 (N_18896,N_18715,N_18147);
nor U18897 (N_18897,N_18645,N_18505);
and U18898 (N_18898,N_18199,N_18208);
nand U18899 (N_18899,N_18546,N_18465);
xor U18900 (N_18900,N_18506,N_18610);
nand U18901 (N_18901,N_18731,N_18581);
and U18902 (N_18902,N_18134,N_18593);
or U18903 (N_18903,N_18545,N_18285);
and U18904 (N_18904,N_18526,N_18129);
xor U18905 (N_18905,N_18704,N_18607);
and U18906 (N_18906,N_18152,N_18662);
or U18907 (N_18907,N_18443,N_18521);
xnor U18908 (N_18908,N_18577,N_18721);
nor U18909 (N_18909,N_18283,N_18140);
nor U18910 (N_18910,N_18575,N_18660);
nor U18911 (N_18911,N_18391,N_18130);
xnor U18912 (N_18912,N_18411,N_18647);
or U18913 (N_18913,N_18477,N_18705);
xor U18914 (N_18914,N_18699,N_18669);
nor U18915 (N_18915,N_18493,N_18318);
or U18916 (N_18916,N_18300,N_18676);
and U18917 (N_18917,N_18643,N_18430);
and U18918 (N_18918,N_18428,N_18617);
xor U18919 (N_18919,N_18733,N_18256);
nand U18920 (N_18920,N_18594,N_18486);
and U18921 (N_18921,N_18143,N_18520);
xor U18922 (N_18922,N_18173,N_18459);
nor U18923 (N_18923,N_18503,N_18600);
nor U18924 (N_18924,N_18162,N_18472);
nand U18925 (N_18925,N_18423,N_18271);
or U18926 (N_18926,N_18340,N_18193);
nor U18927 (N_18927,N_18560,N_18537);
xor U18928 (N_18928,N_18516,N_18551);
and U18929 (N_18929,N_18696,N_18586);
nand U18930 (N_18930,N_18186,N_18556);
nand U18931 (N_18931,N_18133,N_18612);
xnor U18932 (N_18932,N_18268,N_18135);
nor U18933 (N_18933,N_18609,N_18233);
nand U18934 (N_18934,N_18606,N_18622);
nand U18935 (N_18935,N_18636,N_18296);
or U18936 (N_18936,N_18684,N_18483);
nand U18937 (N_18937,N_18196,N_18239);
nor U18938 (N_18938,N_18327,N_18255);
nor U18939 (N_18939,N_18703,N_18700);
or U18940 (N_18940,N_18313,N_18293);
nand U18941 (N_18941,N_18197,N_18189);
nor U18942 (N_18942,N_18324,N_18348);
xor U18943 (N_18943,N_18743,N_18234);
nor U18944 (N_18944,N_18679,N_18252);
and U18945 (N_18945,N_18464,N_18326);
or U18946 (N_18946,N_18241,N_18709);
nor U18947 (N_18947,N_18236,N_18389);
nand U18948 (N_18948,N_18569,N_18449);
nand U18949 (N_18949,N_18539,N_18286);
and U18950 (N_18950,N_18717,N_18306);
or U18951 (N_18951,N_18200,N_18426);
nor U18952 (N_18952,N_18292,N_18466);
and U18953 (N_18953,N_18311,N_18561);
and U18954 (N_18954,N_18538,N_18496);
or U18955 (N_18955,N_18310,N_18304);
or U18956 (N_18956,N_18319,N_18504);
nor U18957 (N_18957,N_18220,N_18320);
nand U18958 (N_18958,N_18224,N_18629);
xor U18959 (N_18959,N_18365,N_18180);
and U18960 (N_18960,N_18350,N_18543);
nor U18961 (N_18961,N_18312,N_18469);
nor U18962 (N_18962,N_18713,N_18336);
nand U18963 (N_18963,N_18232,N_18729);
nand U18964 (N_18964,N_18665,N_18446);
nand U18965 (N_18965,N_18571,N_18531);
and U18966 (N_18966,N_18194,N_18682);
and U18967 (N_18967,N_18279,N_18289);
and U18968 (N_18968,N_18431,N_18702);
xnor U18969 (N_18969,N_18740,N_18395);
xor U18970 (N_18970,N_18565,N_18183);
nor U18971 (N_18971,N_18657,N_18618);
nor U18972 (N_18972,N_18416,N_18646);
and U18973 (N_18973,N_18363,N_18614);
nand U18974 (N_18974,N_18337,N_18535);
and U18975 (N_18975,N_18131,N_18332);
or U18976 (N_18976,N_18680,N_18598);
and U18977 (N_18977,N_18138,N_18620);
nand U18978 (N_18978,N_18182,N_18592);
nor U18979 (N_18979,N_18165,N_18689);
and U18980 (N_18980,N_18145,N_18159);
nor U18981 (N_18981,N_18379,N_18489);
xor U18982 (N_18982,N_18137,N_18549);
nor U18983 (N_18983,N_18314,N_18557);
or U18984 (N_18984,N_18674,N_18396);
xnor U18985 (N_18985,N_18688,N_18375);
nand U18986 (N_18986,N_18381,N_18344);
or U18987 (N_18987,N_18695,N_18376);
xnor U18988 (N_18988,N_18362,N_18307);
xor U18989 (N_18989,N_18360,N_18727);
or U18990 (N_18990,N_18533,N_18736);
and U18991 (N_18991,N_18528,N_18455);
or U18992 (N_18992,N_18508,N_18216);
or U18993 (N_18993,N_18523,N_18275);
nand U18994 (N_18994,N_18652,N_18644);
or U18995 (N_18995,N_18462,N_18467);
and U18996 (N_18996,N_18488,N_18414);
or U18997 (N_18997,N_18661,N_18510);
nand U18998 (N_18998,N_18582,N_18425);
nand U18999 (N_18999,N_18354,N_18626);
and U19000 (N_19000,N_18678,N_18335);
xor U19001 (N_19001,N_18509,N_18564);
nor U19002 (N_19002,N_18631,N_18225);
xnor U19003 (N_19003,N_18419,N_18722);
and U19004 (N_19004,N_18500,N_18125);
nor U19005 (N_19005,N_18212,N_18532);
or U19006 (N_19006,N_18515,N_18177);
or U19007 (N_19007,N_18144,N_18686);
nand U19008 (N_19008,N_18284,N_18734);
and U19009 (N_19009,N_18258,N_18420);
nand U19010 (N_19010,N_18149,N_18639);
and U19011 (N_19011,N_18393,N_18308);
xnor U19012 (N_19012,N_18323,N_18597);
nand U19013 (N_19013,N_18648,N_18250);
and U19014 (N_19014,N_18160,N_18451);
xor U19015 (N_19015,N_18195,N_18251);
and U19016 (N_19016,N_18470,N_18333);
nor U19017 (N_19017,N_18198,N_18441);
and U19018 (N_19018,N_18405,N_18351);
or U19019 (N_19019,N_18507,N_18591);
xnor U19020 (N_19020,N_18364,N_18724);
nand U19021 (N_19021,N_18739,N_18484);
nor U19022 (N_19022,N_18210,N_18383);
nor U19023 (N_19023,N_18714,N_18338);
or U19024 (N_19024,N_18397,N_18305);
xor U19025 (N_19025,N_18492,N_18366);
xor U19026 (N_19026,N_18163,N_18421);
xnor U19027 (N_19027,N_18604,N_18744);
or U19028 (N_19028,N_18544,N_18589);
nor U19029 (N_19029,N_18514,N_18202);
and U19030 (N_19030,N_18737,N_18642);
xnor U19031 (N_19031,N_18747,N_18540);
xnor U19032 (N_19032,N_18553,N_18209);
nor U19033 (N_19033,N_18458,N_18204);
xnor U19034 (N_19034,N_18424,N_18235);
nand U19035 (N_19035,N_18357,N_18563);
xnor U19036 (N_19036,N_18547,N_18627);
nand U19037 (N_19037,N_18226,N_18649);
and U19038 (N_19038,N_18153,N_18708);
or U19039 (N_19039,N_18244,N_18361);
nand U19040 (N_19040,N_18541,N_18328);
xor U19041 (N_19041,N_18718,N_18276);
and U19042 (N_19042,N_18247,N_18511);
nor U19043 (N_19043,N_18630,N_18151);
nand U19044 (N_19044,N_18422,N_18585);
nand U19045 (N_19045,N_18439,N_18412);
xor U19046 (N_19046,N_18548,N_18672);
xnor U19047 (N_19047,N_18386,N_18482);
nor U19048 (N_19048,N_18249,N_18619);
xnor U19049 (N_19049,N_18588,N_18148);
and U19050 (N_19050,N_18406,N_18576);
nor U19051 (N_19051,N_18377,N_18568);
xnor U19052 (N_19052,N_18253,N_18299);
nand U19053 (N_19053,N_18691,N_18519);
nor U19054 (N_19054,N_18452,N_18562);
nand U19055 (N_19055,N_18154,N_18491);
xor U19056 (N_19056,N_18394,N_18229);
nor U19057 (N_19057,N_18270,N_18746);
or U19058 (N_19058,N_18291,N_18368);
nor U19059 (N_19059,N_18322,N_18223);
nor U19060 (N_19060,N_18608,N_18206);
nand U19061 (N_19061,N_18499,N_18663);
and U19062 (N_19062,N_18726,N_18672);
xor U19063 (N_19063,N_18723,N_18320);
nor U19064 (N_19064,N_18623,N_18515);
and U19065 (N_19065,N_18519,N_18735);
xnor U19066 (N_19066,N_18285,N_18379);
and U19067 (N_19067,N_18526,N_18618);
xnor U19068 (N_19068,N_18273,N_18241);
or U19069 (N_19069,N_18622,N_18727);
or U19070 (N_19070,N_18426,N_18166);
nor U19071 (N_19071,N_18138,N_18355);
nand U19072 (N_19072,N_18264,N_18291);
or U19073 (N_19073,N_18162,N_18184);
and U19074 (N_19074,N_18278,N_18448);
xor U19075 (N_19075,N_18339,N_18587);
nor U19076 (N_19076,N_18574,N_18219);
or U19077 (N_19077,N_18618,N_18450);
and U19078 (N_19078,N_18226,N_18217);
or U19079 (N_19079,N_18411,N_18439);
nand U19080 (N_19080,N_18495,N_18592);
nor U19081 (N_19081,N_18701,N_18161);
and U19082 (N_19082,N_18180,N_18634);
xor U19083 (N_19083,N_18432,N_18498);
and U19084 (N_19084,N_18418,N_18607);
or U19085 (N_19085,N_18707,N_18142);
nor U19086 (N_19086,N_18501,N_18296);
nand U19087 (N_19087,N_18325,N_18244);
or U19088 (N_19088,N_18356,N_18666);
nor U19089 (N_19089,N_18533,N_18711);
and U19090 (N_19090,N_18208,N_18560);
and U19091 (N_19091,N_18465,N_18311);
and U19092 (N_19092,N_18276,N_18127);
and U19093 (N_19093,N_18182,N_18262);
and U19094 (N_19094,N_18264,N_18171);
and U19095 (N_19095,N_18569,N_18537);
nor U19096 (N_19096,N_18585,N_18235);
or U19097 (N_19097,N_18566,N_18434);
nand U19098 (N_19098,N_18722,N_18323);
or U19099 (N_19099,N_18346,N_18719);
nor U19100 (N_19100,N_18683,N_18570);
and U19101 (N_19101,N_18630,N_18331);
nor U19102 (N_19102,N_18295,N_18374);
nand U19103 (N_19103,N_18243,N_18488);
nand U19104 (N_19104,N_18383,N_18678);
and U19105 (N_19105,N_18516,N_18262);
nand U19106 (N_19106,N_18561,N_18515);
or U19107 (N_19107,N_18360,N_18610);
nand U19108 (N_19108,N_18215,N_18267);
and U19109 (N_19109,N_18155,N_18335);
and U19110 (N_19110,N_18491,N_18323);
nor U19111 (N_19111,N_18508,N_18643);
nor U19112 (N_19112,N_18549,N_18401);
and U19113 (N_19113,N_18580,N_18170);
xor U19114 (N_19114,N_18607,N_18195);
nand U19115 (N_19115,N_18529,N_18549);
xor U19116 (N_19116,N_18223,N_18208);
nor U19117 (N_19117,N_18135,N_18558);
nor U19118 (N_19118,N_18459,N_18636);
nand U19119 (N_19119,N_18511,N_18603);
xor U19120 (N_19120,N_18253,N_18678);
xnor U19121 (N_19121,N_18174,N_18143);
or U19122 (N_19122,N_18734,N_18610);
nor U19123 (N_19123,N_18341,N_18391);
nor U19124 (N_19124,N_18693,N_18681);
nor U19125 (N_19125,N_18264,N_18309);
and U19126 (N_19126,N_18219,N_18225);
and U19127 (N_19127,N_18419,N_18199);
xor U19128 (N_19128,N_18184,N_18338);
nand U19129 (N_19129,N_18551,N_18684);
xor U19130 (N_19130,N_18551,N_18440);
xor U19131 (N_19131,N_18142,N_18534);
or U19132 (N_19132,N_18290,N_18372);
nor U19133 (N_19133,N_18444,N_18162);
xor U19134 (N_19134,N_18393,N_18428);
and U19135 (N_19135,N_18617,N_18158);
and U19136 (N_19136,N_18436,N_18654);
nor U19137 (N_19137,N_18725,N_18595);
nor U19138 (N_19138,N_18396,N_18282);
xnor U19139 (N_19139,N_18220,N_18677);
and U19140 (N_19140,N_18353,N_18208);
xnor U19141 (N_19141,N_18128,N_18701);
nor U19142 (N_19142,N_18175,N_18471);
or U19143 (N_19143,N_18473,N_18706);
nor U19144 (N_19144,N_18196,N_18172);
xnor U19145 (N_19145,N_18641,N_18304);
nor U19146 (N_19146,N_18354,N_18273);
xor U19147 (N_19147,N_18506,N_18491);
nor U19148 (N_19148,N_18228,N_18436);
or U19149 (N_19149,N_18316,N_18384);
or U19150 (N_19150,N_18711,N_18430);
nor U19151 (N_19151,N_18425,N_18718);
xnor U19152 (N_19152,N_18252,N_18272);
nand U19153 (N_19153,N_18430,N_18373);
nor U19154 (N_19154,N_18343,N_18250);
and U19155 (N_19155,N_18685,N_18182);
nand U19156 (N_19156,N_18566,N_18272);
nor U19157 (N_19157,N_18475,N_18490);
or U19158 (N_19158,N_18142,N_18568);
or U19159 (N_19159,N_18579,N_18203);
xnor U19160 (N_19160,N_18372,N_18338);
or U19161 (N_19161,N_18487,N_18640);
and U19162 (N_19162,N_18424,N_18748);
nor U19163 (N_19163,N_18358,N_18300);
xor U19164 (N_19164,N_18303,N_18345);
nand U19165 (N_19165,N_18593,N_18306);
or U19166 (N_19166,N_18640,N_18177);
xnor U19167 (N_19167,N_18278,N_18323);
and U19168 (N_19168,N_18503,N_18265);
nand U19169 (N_19169,N_18308,N_18285);
nand U19170 (N_19170,N_18498,N_18408);
or U19171 (N_19171,N_18404,N_18355);
nor U19172 (N_19172,N_18194,N_18377);
and U19173 (N_19173,N_18324,N_18141);
or U19174 (N_19174,N_18184,N_18144);
xnor U19175 (N_19175,N_18156,N_18522);
nand U19176 (N_19176,N_18428,N_18580);
and U19177 (N_19177,N_18408,N_18293);
xor U19178 (N_19178,N_18598,N_18236);
and U19179 (N_19179,N_18524,N_18724);
xor U19180 (N_19180,N_18682,N_18322);
nor U19181 (N_19181,N_18456,N_18464);
nor U19182 (N_19182,N_18268,N_18562);
or U19183 (N_19183,N_18524,N_18423);
and U19184 (N_19184,N_18386,N_18346);
or U19185 (N_19185,N_18707,N_18600);
and U19186 (N_19186,N_18269,N_18271);
nor U19187 (N_19187,N_18152,N_18258);
or U19188 (N_19188,N_18548,N_18356);
and U19189 (N_19189,N_18488,N_18476);
nand U19190 (N_19190,N_18233,N_18299);
and U19191 (N_19191,N_18599,N_18714);
and U19192 (N_19192,N_18545,N_18250);
and U19193 (N_19193,N_18698,N_18556);
and U19194 (N_19194,N_18273,N_18194);
xor U19195 (N_19195,N_18556,N_18253);
nor U19196 (N_19196,N_18222,N_18192);
nand U19197 (N_19197,N_18496,N_18689);
nand U19198 (N_19198,N_18143,N_18399);
and U19199 (N_19199,N_18305,N_18653);
and U19200 (N_19200,N_18526,N_18604);
nand U19201 (N_19201,N_18374,N_18623);
and U19202 (N_19202,N_18523,N_18181);
xor U19203 (N_19203,N_18587,N_18331);
xnor U19204 (N_19204,N_18380,N_18355);
nor U19205 (N_19205,N_18595,N_18502);
or U19206 (N_19206,N_18666,N_18479);
nand U19207 (N_19207,N_18199,N_18714);
or U19208 (N_19208,N_18429,N_18424);
xor U19209 (N_19209,N_18655,N_18589);
and U19210 (N_19210,N_18292,N_18604);
and U19211 (N_19211,N_18134,N_18728);
and U19212 (N_19212,N_18288,N_18407);
or U19213 (N_19213,N_18308,N_18295);
nor U19214 (N_19214,N_18541,N_18665);
nor U19215 (N_19215,N_18592,N_18155);
or U19216 (N_19216,N_18431,N_18475);
xnor U19217 (N_19217,N_18564,N_18221);
or U19218 (N_19218,N_18343,N_18687);
or U19219 (N_19219,N_18423,N_18147);
xor U19220 (N_19220,N_18640,N_18131);
or U19221 (N_19221,N_18214,N_18484);
and U19222 (N_19222,N_18469,N_18147);
and U19223 (N_19223,N_18215,N_18147);
nand U19224 (N_19224,N_18501,N_18642);
or U19225 (N_19225,N_18522,N_18248);
xor U19226 (N_19226,N_18692,N_18571);
xor U19227 (N_19227,N_18566,N_18273);
nor U19228 (N_19228,N_18615,N_18221);
nand U19229 (N_19229,N_18664,N_18294);
nor U19230 (N_19230,N_18326,N_18318);
or U19231 (N_19231,N_18377,N_18272);
nor U19232 (N_19232,N_18238,N_18343);
and U19233 (N_19233,N_18339,N_18436);
nor U19234 (N_19234,N_18617,N_18403);
xor U19235 (N_19235,N_18625,N_18685);
nand U19236 (N_19236,N_18412,N_18278);
and U19237 (N_19237,N_18613,N_18584);
or U19238 (N_19238,N_18560,N_18159);
and U19239 (N_19239,N_18168,N_18673);
or U19240 (N_19240,N_18133,N_18517);
and U19241 (N_19241,N_18533,N_18138);
nor U19242 (N_19242,N_18711,N_18283);
xor U19243 (N_19243,N_18264,N_18497);
nor U19244 (N_19244,N_18704,N_18316);
xnor U19245 (N_19245,N_18374,N_18581);
nand U19246 (N_19246,N_18156,N_18359);
or U19247 (N_19247,N_18359,N_18685);
nand U19248 (N_19248,N_18303,N_18590);
or U19249 (N_19249,N_18511,N_18740);
and U19250 (N_19250,N_18239,N_18586);
nor U19251 (N_19251,N_18468,N_18621);
nor U19252 (N_19252,N_18552,N_18666);
or U19253 (N_19253,N_18722,N_18230);
nor U19254 (N_19254,N_18542,N_18632);
or U19255 (N_19255,N_18598,N_18567);
nand U19256 (N_19256,N_18641,N_18554);
or U19257 (N_19257,N_18382,N_18695);
and U19258 (N_19258,N_18626,N_18549);
nor U19259 (N_19259,N_18522,N_18315);
nand U19260 (N_19260,N_18147,N_18647);
or U19261 (N_19261,N_18297,N_18730);
nand U19262 (N_19262,N_18287,N_18170);
xor U19263 (N_19263,N_18316,N_18223);
and U19264 (N_19264,N_18478,N_18265);
and U19265 (N_19265,N_18531,N_18310);
and U19266 (N_19266,N_18567,N_18684);
nor U19267 (N_19267,N_18219,N_18737);
nor U19268 (N_19268,N_18630,N_18659);
nor U19269 (N_19269,N_18129,N_18180);
nor U19270 (N_19270,N_18648,N_18269);
and U19271 (N_19271,N_18261,N_18197);
nand U19272 (N_19272,N_18351,N_18373);
or U19273 (N_19273,N_18377,N_18579);
xnor U19274 (N_19274,N_18385,N_18380);
xnor U19275 (N_19275,N_18165,N_18617);
nor U19276 (N_19276,N_18126,N_18252);
nor U19277 (N_19277,N_18652,N_18159);
nor U19278 (N_19278,N_18261,N_18560);
and U19279 (N_19279,N_18477,N_18565);
nand U19280 (N_19280,N_18452,N_18457);
nand U19281 (N_19281,N_18433,N_18435);
nor U19282 (N_19282,N_18214,N_18736);
nand U19283 (N_19283,N_18264,N_18656);
nor U19284 (N_19284,N_18359,N_18527);
nor U19285 (N_19285,N_18616,N_18602);
nor U19286 (N_19286,N_18592,N_18146);
xor U19287 (N_19287,N_18339,N_18257);
or U19288 (N_19288,N_18572,N_18649);
xor U19289 (N_19289,N_18348,N_18298);
or U19290 (N_19290,N_18127,N_18633);
nor U19291 (N_19291,N_18573,N_18602);
or U19292 (N_19292,N_18446,N_18741);
nand U19293 (N_19293,N_18172,N_18268);
nand U19294 (N_19294,N_18310,N_18138);
and U19295 (N_19295,N_18535,N_18727);
nor U19296 (N_19296,N_18292,N_18671);
and U19297 (N_19297,N_18280,N_18520);
and U19298 (N_19298,N_18216,N_18646);
nor U19299 (N_19299,N_18382,N_18301);
or U19300 (N_19300,N_18297,N_18464);
xnor U19301 (N_19301,N_18577,N_18615);
or U19302 (N_19302,N_18323,N_18389);
nor U19303 (N_19303,N_18139,N_18612);
xor U19304 (N_19304,N_18164,N_18704);
and U19305 (N_19305,N_18259,N_18216);
nand U19306 (N_19306,N_18563,N_18559);
nand U19307 (N_19307,N_18195,N_18376);
nor U19308 (N_19308,N_18254,N_18170);
xnor U19309 (N_19309,N_18610,N_18490);
or U19310 (N_19310,N_18728,N_18671);
xnor U19311 (N_19311,N_18316,N_18649);
or U19312 (N_19312,N_18280,N_18475);
and U19313 (N_19313,N_18125,N_18196);
nor U19314 (N_19314,N_18533,N_18152);
xnor U19315 (N_19315,N_18262,N_18556);
nor U19316 (N_19316,N_18227,N_18410);
or U19317 (N_19317,N_18541,N_18197);
nor U19318 (N_19318,N_18363,N_18548);
xor U19319 (N_19319,N_18551,N_18478);
nand U19320 (N_19320,N_18230,N_18202);
xnor U19321 (N_19321,N_18502,N_18232);
xnor U19322 (N_19322,N_18140,N_18440);
xor U19323 (N_19323,N_18651,N_18361);
or U19324 (N_19324,N_18451,N_18673);
and U19325 (N_19325,N_18411,N_18503);
xor U19326 (N_19326,N_18166,N_18537);
nor U19327 (N_19327,N_18265,N_18636);
and U19328 (N_19328,N_18414,N_18630);
or U19329 (N_19329,N_18415,N_18265);
or U19330 (N_19330,N_18381,N_18682);
and U19331 (N_19331,N_18705,N_18433);
and U19332 (N_19332,N_18434,N_18480);
nand U19333 (N_19333,N_18378,N_18480);
xnor U19334 (N_19334,N_18432,N_18683);
or U19335 (N_19335,N_18134,N_18226);
or U19336 (N_19336,N_18341,N_18460);
nand U19337 (N_19337,N_18393,N_18551);
and U19338 (N_19338,N_18275,N_18291);
nand U19339 (N_19339,N_18271,N_18536);
or U19340 (N_19340,N_18207,N_18203);
or U19341 (N_19341,N_18413,N_18578);
and U19342 (N_19342,N_18640,N_18432);
nor U19343 (N_19343,N_18199,N_18716);
nand U19344 (N_19344,N_18665,N_18722);
or U19345 (N_19345,N_18636,N_18345);
nor U19346 (N_19346,N_18701,N_18259);
nand U19347 (N_19347,N_18155,N_18526);
or U19348 (N_19348,N_18310,N_18317);
xnor U19349 (N_19349,N_18515,N_18707);
xnor U19350 (N_19350,N_18528,N_18714);
nor U19351 (N_19351,N_18179,N_18279);
and U19352 (N_19352,N_18658,N_18219);
or U19353 (N_19353,N_18662,N_18229);
nor U19354 (N_19354,N_18560,N_18735);
or U19355 (N_19355,N_18471,N_18304);
nor U19356 (N_19356,N_18340,N_18254);
or U19357 (N_19357,N_18692,N_18455);
nor U19358 (N_19358,N_18606,N_18134);
or U19359 (N_19359,N_18381,N_18400);
or U19360 (N_19360,N_18728,N_18173);
xnor U19361 (N_19361,N_18540,N_18441);
nand U19362 (N_19362,N_18439,N_18161);
nor U19363 (N_19363,N_18447,N_18546);
xor U19364 (N_19364,N_18246,N_18677);
nor U19365 (N_19365,N_18610,N_18694);
and U19366 (N_19366,N_18403,N_18721);
and U19367 (N_19367,N_18510,N_18172);
nor U19368 (N_19368,N_18283,N_18235);
xnor U19369 (N_19369,N_18212,N_18279);
and U19370 (N_19370,N_18266,N_18621);
xor U19371 (N_19371,N_18197,N_18308);
or U19372 (N_19372,N_18173,N_18502);
or U19373 (N_19373,N_18327,N_18187);
xor U19374 (N_19374,N_18744,N_18125);
and U19375 (N_19375,N_18970,N_18990);
nand U19376 (N_19376,N_18938,N_19096);
nor U19377 (N_19377,N_19020,N_19332);
nand U19378 (N_19378,N_18948,N_19256);
nor U19379 (N_19379,N_18822,N_18855);
and U19380 (N_19380,N_18965,N_19040);
and U19381 (N_19381,N_18977,N_19154);
nor U19382 (N_19382,N_19266,N_19341);
or U19383 (N_19383,N_19172,N_19369);
or U19384 (N_19384,N_18945,N_19112);
and U19385 (N_19385,N_19336,N_18987);
nor U19386 (N_19386,N_18845,N_19026);
and U19387 (N_19387,N_19145,N_18810);
nor U19388 (N_19388,N_18867,N_18930);
and U19389 (N_19389,N_18826,N_19165);
xor U19390 (N_19390,N_18964,N_18903);
and U19391 (N_19391,N_19102,N_18849);
nand U19392 (N_19392,N_18901,N_18842);
nor U19393 (N_19393,N_19058,N_19185);
nor U19394 (N_19394,N_18952,N_18991);
nand U19395 (N_19395,N_19150,N_19033);
nor U19396 (N_19396,N_19351,N_19297);
xor U19397 (N_19397,N_19121,N_19328);
or U19398 (N_19398,N_18992,N_18864);
nor U19399 (N_19399,N_19092,N_19244);
or U19400 (N_19400,N_19246,N_19180);
nor U19401 (N_19401,N_18973,N_19048);
or U19402 (N_19402,N_19002,N_19343);
nand U19403 (N_19403,N_19074,N_18981);
and U19404 (N_19404,N_19116,N_18914);
or U19405 (N_19405,N_19182,N_19089);
nand U19406 (N_19406,N_19070,N_18881);
or U19407 (N_19407,N_19198,N_19207);
and U19408 (N_19408,N_19294,N_19114);
xor U19409 (N_19409,N_19255,N_19273);
nand U19410 (N_19410,N_19326,N_19071);
and U19411 (N_19411,N_19196,N_19358);
or U19412 (N_19412,N_19300,N_19005);
xor U19413 (N_19413,N_18850,N_18913);
nor U19414 (N_19414,N_19288,N_18820);
or U19415 (N_19415,N_18900,N_19023);
nand U19416 (N_19416,N_19100,N_18971);
xor U19417 (N_19417,N_18969,N_18986);
or U19418 (N_19418,N_19143,N_19148);
and U19419 (N_19419,N_19193,N_19238);
nor U19420 (N_19420,N_19069,N_18931);
or U19421 (N_19421,N_19038,N_19280);
and U19422 (N_19422,N_19050,N_19313);
or U19423 (N_19423,N_19331,N_19211);
xor U19424 (N_19424,N_19134,N_18804);
or U19425 (N_19425,N_18829,N_18780);
nand U19426 (N_19426,N_18768,N_19159);
or U19427 (N_19427,N_19021,N_19093);
nand U19428 (N_19428,N_19153,N_19212);
or U19429 (N_19429,N_18787,N_19208);
or U19430 (N_19430,N_19122,N_19022);
nand U19431 (N_19431,N_18925,N_19200);
nand U19432 (N_19432,N_19278,N_19029);
and U19433 (N_19433,N_18805,N_19129);
nand U19434 (N_19434,N_18764,N_19242);
nand U19435 (N_19435,N_19373,N_18801);
and U19436 (N_19436,N_19146,N_18889);
nand U19437 (N_19437,N_19101,N_18825);
and U19438 (N_19438,N_19276,N_18834);
nand U19439 (N_19439,N_18890,N_19220);
nand U19440 (N_19440,N_18766,N_19085);
xor U19441 (N_19441,N_19035,N_19016);
nand U19442 (N_19442,N_18891,N_19285);
or U19443 (N_19443,N_18781,N_19107);
nor U19444 (N_19444,N_19282,N_19299);
and U19445 (N_19445,N_18885,N_19304);
nand U19446 (N_19446,N_18773,N_18754);
and U19447 (N_19447,N_18934,N_19361);
xor U19448 (N_19448,N_18921,N_18776);
and U19449 (N_19449,N_19357,N_19311);
or U19450 (N_19450,N_18816,N_19229);
nand U19451 (N_19451,N_19362,N_19367);
nand U19452 (N_19452,N_19059,N_19004);
xor U19453 (N_19453,N_18908,N_19296);
nor U19454 (N_19454,N_19152,N_19133);
xor U19455 (N_19455,N_18761,N_19157);
xnor U19456 (N_19456,N_19090,N_18847);
xor U19457 (N_19457,N_19213,N_19291);
and U19458 (N_19458,N_19302,N_19234);
xnor U19459 (N_19459,N_19334,N_18767);
xor U19460 (N_19460,N_19352,N_18916);
or U19461 (N_19461,N_18750,N_19014);
or U19462 (N_19462,N_19173,N_19345);
xnor U19463 (N_19463,N_19252,N_19015);
nor U19464 (N_19464,N_19118,N_18996);
or U19465 (N_19465,N_19062,N_19295);
xnor U19466 (N_19466,N_18865,N_19272);
nor U19467 (N_19467,N_19161,N_19019);
and U19468 (N_19468,N_19123,N_19043);
nor U19469 (N_19469,N_19241,N_18836);
nor U19470 (N_19470,N_19080,N_19258);
xor U19471 (N_19471,N_18888,N_19077);
nand U19472 (N_19472,N_18868,N_19309);
or U19473 (N_19473,N_19222,N_19030);
xor U19474 (N_19474,N_19009,N_18758);
nor U19475 (N_19475,N_19247,N_19110);
and U19476 (N_19476,N_18994,N_19171);
or U19477 (N_19477,N_19265,N_19149);
xor U19478 (N_19478,N_18823,N_18751);
and U19479 (N_19479,N_18924,N_19250);
nand U19480 (N_19480,N_19012,N_19219);
and U19481 (N_19481,N_19327,N_19235);
nand U19482 (N_19482,N_19187,N_19174);
or U19483 (N_19483,N_18929,N_19271);
and U19484 (N_19484,N_18935,N_19053);
or U19485 (N_19485,N_19314,N_19191);
and U19486 (N_19486,N_19308,N_19216);
and U19487 (N_19487,N_18809,N_18880);
and U19488 (N_19488,N_19087,N_19274);
nand U19489 (N_19489,N_19210,N_19371);
and U19490 (N_19490,N_19163,N_19042);
nand U19491 (N_19491,N_18910,N_18875);
nor U19492 (N_19492,N_19061,N_19228);
nor U19493 (N_19493,N_19136,N_18897);
nor U19494 (N_19494,N_19318,N_19108);
xnor U19495 (N_19495,N_19325,N_19287);
and U19496 (N_19496,N_19013,N_19137);
and U19497 (N_19497,N_19164,N_19037);
xnor U19498 (N_19498,N_19056,N_18874);
xor U19499 (N_19499,N_19218,N_19183);
and U19500 (N_19500,N_18869,N_19227);
or U19501 (N_19501,N_19088,N_19011);
xnor U19502 (N_19502,N_18879,N_19251);
nor U19503 (N_19503,N_19073,N_18846);
xor U19504 (N_19504,N_18794,N_19094);
xor U19505 (N_19505,N_18968,N_19225);
nand U19506 (N_19506,N_19168,N_18976);
nor U19507 (N_19507,N_18792,N_18852);
nand U19508 (N_19508,N_19141,N_19259);
or U19509 (N_19509,N_19203,N_19236);
nand U19510 (N_19510,N_19270,N_19018);
xnor U19511 (N_19511,N_19349,N_19201);
xnor U19512 (N_19512,N_19156,N_18831);
or U19513 (N_19513,N_19105,N_18827);
xnor U19514 (N_19514,N_19374,N_18830);
xor U19515 (N_19515,N_19097,N_18843);
and U19516 (N_19516,N_18799,N_18815);
xor U19517 (N_19517,N_19158,N_19214);
or U19518 (N_19518,N_18797,N_19065);
nor U19519 (N_19519,N_18927,N_19209);
xor U19520 (N_19520,N_19269,N_19360);
or U19521 (N_19521,N_19281,N_18771);
or U19522 (N_19522,N_18893,N_18942);
nor U19523 (N_19523,N_19315,N_19032);
and U19524 (N_19524,N_19151,N_19139);
nand U19525 (N_19525,N_18756,N_18886);
or U19526 (N_19526,N_19338,N_18922);
and U19527 (N_19527,N_18943,N_19322);
nor U19528 (N_19528,N_19243,N_18819);
or U19529 (N_19529,N_19249,N_18993);
nor U19530 (N_19530,N_18769,N_19205);
nor U19531 (N_19531,N_18800,N_19135);
or U19532 (N_19532,N_19106,N_18862);
xnor U19533 (N_19533,N_19066,N_18998);
nor U19534 (N_19534,N_18839,N_19081);
or U19535 (N_19535,N_19292,N_19197);
xnor U19536 (N_19536,N_18923,N_19041);
nor U19537 (N_19537,N_18783,N_19082);
nor U19538 (N_19538,N_19025,N_18803);
and U19539 (N_19539,N_19231,N_19142);
nand U19540 (N_19540,N_18848,N_18940);
or U19541 (N_19541,N_19335,N_19047);
and U19542 (N_19542,N_19060,N_18902);
nor U19543 (N_19543,N_19323,N_19293);
and U19544 (N_19544,N_19348,N_19199);
and U19545 (N_19545,N_19124,N_19086);
nor U19546 (N_19546,N_19181,N_18956);
nand U19547 (N_19547,N_19028,N_19290);
nand U19548 (N_19548,N_18904,N_19232);
nor U19549 (N_19549,N_18953,N_19103);
xnor U19550 (N_19550,N_19359,N_18877);
xnor U19551 (N_19551,N_19039,N_18966);
nand U19552 (N_19552,N_19289,N_18790);
or U19553 (N_19553,N_19075,N_19329);
and U19554 (N_19554,N_18866,N_19303);
nand U19555 (N_19555,N_19054,N_18860);
nand U19556 (N_19556,N_18906,N_18912);
or U19557 (N_19557,N_19253,N_18932);
xor U19558 (N_19558,N_19277,N_19223);
xnor U19559 (N_19559,N_19179,N_19319);
nor U19560 (N_19560,N_18917,N_19144);
nor U19561 (N_19561,N_19215,N_19279);
nor U19562 (N_19562,N_19049,N_19057);
and U19563 (N_19563,N_19366,N_19119);
or U19564 (N_19564,N_19027,N_19340);
nand U19565 (N_19565,N_19160,N_19128);
and U19566 (N_19566,N_19125,N_19192);
xor U19567 (N_19567,N_19339,N_19068);
xor U19568 (N_19568,N_18833,N_19147);
or U19569 (N_19569,N_18988,N_18757);
xnor U19570 (N_19570,N_19190,N_19344);
and U19571 (N_19571,N_19007,N_18961);
nand U19572 (N_19572,N_18895,N_19240);
nand U19573 (N_19573,N_19298,N_18928);
or U19574 (N_19574,N_18944,N_19230);
xnor U19575 (N_19575,N_19372,N_18907);
or U19576 (N_19576,N_19310,N_19237);
nand U19577 (N_19577,N_19051,N_18853);
xnor U19578 (N_19578,N_19368,N_19098);
xor U19579 (N_19579,N_19120,N_19226);
and U19580 (N_19580,N_18979,N_18920);
nand U19581 (N_19581,N_19084,N_18808);
xor U19582 (N_19582,N_19010,N_19127);
or U19583 (N_19583,N_18898,N_19354);
nor U19584 (N_19584,N_19260,N_18974);
nor U19585 (N_19585,N_18775,N_18892);
or U19586 (N_19586,N_19003,N_18765);
nor U19587 (N_19587,N_19111,N_19166);
or U19588 (N_19588,N_18854,N_19370);
xor U19589 (N_19589,N_19130,N_18814);
and U19590 (N_19590,N_18997,N_18975);
nand U19591 (N_19591,N_19264,N_19320);
and U19592 (N_19592,N_19275,N_18995);
xnor U19593 (N_19593,N_18899,N_19099);
nand U19594 (N_19594,N_18789,N_19178);
or U19595 (N_19595,N_19248,N_19365);
nor U19596 (N_19596,N_19184,N_19064);
nand U19597 (N_19597,N_19044,N_18777);
or U19598 (N_19598,N_19346,N_18963);
xor U19599 (N_19599,N_19353,N_18989);
xor U19600 (N_19600,N_18958,N_19189);
nor U19601 (N_19601,N_18872,N_19206);
nand U19602 (N_19602,N_18779,N_18796);
and U19603 (N_19603,N_18985,N_19063);
xor U19604 (N_19604,N_19202,N_19046);
xor U19605 (N_19605,N_18763,N_19176);
or U19606 (N_19606,N_18878,N_18905);
xor U19607 (N_19607,N_18844,N_19155);
nor U19608 (N_19608,N_18752,N_19113);
nor U19609 (N_19609,N_18762,N_19283);
and U19610 (N_19610,N_19350,N_18962);
nand U19611 (N_19611,N_19078,N_18936);
nor U19612 (N_19612,N_19217,N_18772);
or U19613 (N_19613,N_18955,N_19017);
or U19614 (N_19614,N_19194,N_19306);
nor U19615 (N_19615,N_19245,N_18785);
xor U19616 (N_19616,N_19006,N_18918);
xor U19617 (N_19617,N_19067,N_19036);
nor U19618 (N_19618,N_18926,N_18774);
and U19619 (N_19619,N_18947,N_19330);
and U19620 (N_19620,N_18798,N_18982);
nand U19621 (N_19621,N_19091,N_19104);
or U19622 (N_19622,N_18821,N_19008);
xor U19623 (N_19623,N_19177,N_18807);
and U19624 (N_19624,N_19186,N_18791);
nand U19625 (N_19625,N_19052,N_18951);
nand U19626 (N_19626,N_18851,N_18863);
or U19627 (N_19627,N_19239,N_19333);
nand U19628 (N_19628,N_19170,N_19363);
xor U19629 (N_19629,N_19162,N_19079);
nand U19630 (N_19630,N_18793,N_18784);
nor U19631 (N_19631,N_18795,N_18949);
xnor U19632 (N_19632,N_19072,N_18978);
nor U19633 (N_19633,N_18937,N_19312);
nor U19634 (N_19634,N_18841,N_19109);
and U19635 (N_19635,N_19316,N_18882);
nand U19636 (N_19636,N_18840,N_18946);
nand U19637 (N_19637,N_18813,N_18832);
or U19638 (N_19638,N_18753,N_19233);
xor U19639 (N_19639,N_18859,N_18883);
or U19640 (N_19640,N_18786,N_19342);
and U19641 (N_19641,N_18950,N_19263);
or U19642 (N_19642,N_18933,N_19131);
or U19643 (N_19643,N_18941,N_18909);
nor U19644 (N_19644,N_18972,N_18770);
nand U19645 (N_19645,N_19286,N_18957);
xnor U19646 (N_19646,N_19117,N_19355);
nand U19647 (N_19647,N_18788,N_18980);
or U19648 (N_19648,N_18999,N_18778);
and U19649 (N_19649,N_19115,N_18894);
and U19650 (N_19650,N_19305,N_19126);
nand U19651 (N_19651,N_18802,N_19001);
and U19652 (N_19652,N_18967,N_18755);
or U19653 (N_19653,N_19031,N_18817);
nand U19654 (N_19654,N_19055,N_19224);
or U19655 (N_19655,N_19167,N_18818);
and U19656 (N_19656,N_18782,N_19254);
xnor U19657 (N_19657,N_19321,N_19356);
nor U19658 (N_19658,N_18835,N_19317);
nor U19659 (N_19659,N_18915,N_18759);
nor U19660 (N_19660,N_19301,N_19095);
or U19661 (N_19661,N_19268,N_18812);
or U19662 (N_19662,N_18861,N_19261);
or U19663 (N_19663,N_18856,N_19169);
and U19664 (N_19664,N_18806,N_18960);
nand U19665 (N_19665,N_19324,N_18871);
xor U19666 (N_19666,N_19083,N_19284);
nand U19667 (N_19667,N_19034,N_19000);
nand U19668 (N_19668,N_18959,N_18811);
nand U19669 (N_19669,N_18760,N_18939);
nor U19670 (N_19670,N_18824,N_18858);
nand U19671 (N_19671,N_18828,N_19364);
nand U19672 (N_19672,N_19307,N_19347);
nand U19673 (N_19673,N_19175,N_19221);
nor U19674 (N_19674,N_19140,N_19024);
or U19675 (N_19675,N_18954,N_19257);
xor U19676 (N_19676,N_19267,N_19076);
xor U19677 (N_19677,N_19138,N_18887);
nand U19678 (N_19678,N_19045,N_18873);
nand U19679 (N_19679,N_19132,N_18919);
nor U19680 (N_19680,N_18884,N_18837);
xnor U19681 (N_19681,N_18857,N_18896);
and U19682 (N_19682,N_19188,N_18984);
nor U19683 (N_19683,N_18983,N_19262);
or U19684 (N_19684,N_18911,N_19195);
xnor U19685 (N_19685,N_18838,N_19204);
xnor U19686 (N_19686,N_18870,N_19337);
xor U19687 (N_19687,N_18876,N_18854);
and U19688 (N_19688,N_19245,N_18991);
or U19689 (N_19689,N_19104,N_19286);
and U19690 (N_19690,N_18818,N_19116);
nand U19691 (N_19691,N_19163,N_19232);
or U19692 (N_19692,N_19137,N_19360);
or U19693 (N_19693,N_19001,N_19280);
nand U19694 (N_19694,N_19212,N_18837);
nor U19695 (N_19695,N_18930,N_18827);
nand U19696 (N_19696,N_19036,N_18974);
nor U19697 (N_19697,N_18796,N_18954);
xnor U19698 (N_19698,N_19307,N_19103);
and U19699 (N_19699,N_19281,N_19274);
nand U19700 (N_19700,N_18895,N_19228);
and U19701 (N_19701,N_19224,N_19273);
nor U19702 (N_19702,N_18946,N_19069);
or U19703 (N_19703,N_18831,N_19135);
nor U19704 (N_19704,N_19287,N_19136);
nor U19705 (N_19705,N_18955,N_19300);
xnor U19706 (N_19706,N_18895,N_18860);
nand U19707 (N_19707,N_19132,N_19245);
xor U19708 (N_19708,N_19257,N_19265);
or U19709 (N_19709,N_19368,N_19197);
or U19710 (N_19710,N_19255,N_19178);
and U19711 (N_19711,N_19279,N_18914);
and U19712 (N_19712,N_19247,N_18987);
nor U19713 (N_19713,N_18791,N_19163);
xor U19714 (N_19714,N_18777,N_18810);
nand U19715 (N_19715,N_19158,N_19273);
and U19716 (N_19716,N_19358,N_19336);
nand U19717 (N_19717,N_19350,N_19281);
and U19718 (N_19718,N_19056,N_19149);
or U19719 (N_19719,N_18791,N_19250);
or U19720 (N_19720,N_19328,N_18925);
xnor U19721 (N_19721,N_19048,N_19312);
and U19722 (N_19722,N_18756,N_19056);
nor U19723 (N_19723,N_19134,N_18800);
xnor U19724 (N_19724,N_18928,N_19032);
and U19725 (N_19725,N_19298,N_19313);
or U19726 (N_19726,N_18792,N_19203);
and U19727 (N_19727,N_18960,N_18840);
nand U19728 (N_19728,N_19069,N_18968);
or U19729 (N_19729,N_19119,N_19355);
and U19730 (N_19730,N_19096,N_18974);
xor U19731 (N_19731,N_18793,N_19347);
xor U19732 (N_19732,N_19125,N_19328);
and U19733 (N_19733,N_19151,N_19316);
nor U19734 (N_19734,N_18907,N_19001);
nor U19735 (N_19735,N_19181,N_18989);
xor U19736 (N_19736,N_19372,N_18790);
nor U19737 (N_19737,N_19233,N_19015);
nor U19738 (N_19738,N_18949,N_19363);
xnor U19739 (N_19739,N_19324,N_18877);
and U19740 (N_19740,N_19081,N_19157);
or U19741 (N_19741,N_19004,N_19215);
nor U19742 (N_19742,N_19367,N_19327);
nand U19743 (N_19743,N_18869,N_19131);
nor U19744 (N_19744,N_19097,N_18958);
nand U19745 (N_19745,N_18951,N_19085);
xnor U19746 (N_19746,N_19145,N_19113);
nand U19747 (N_19747,N_18898,N_19309);
nor U19748 (N_19748,N_18892,N_19294);
nand U19749 (N_19749,N_19318,N_19252);
nor U19750 (N_19750,N_19120,N_18839);
nor U19751 (N_19751,N_18799,N_19272);
xor U19752 (N_19752,N_18881,N_19278);
or U19753 (N_19753,N_19269,N_19163);
nand U19754 (N_19754,N_18954,N_19222);
xor U19755 (N_19755,N_19004,N_19060);
nand U19756 (N_19756,N_18767,N_19222);
xor U19757 (N_19757,N_18870,N_19190);
nand U19758 (N_19758,N_19090,N_19244);
nand U19759 (N_19759,N_19228,N_19239);
or U19760 (N_19760,N_19296,N_18751);
nor U19761 (N_19761,N_19060,N_19020);
nand U19762 (N_19762,N_19219,N_19254);
or U19763 (N_19763,N_19190,N_18936);
nor U19764 (N_19764,N_19251,N_19181);
xor U19765 (N_19765,N_19142,N_18895);
nor U19766 (N_19766,N_19077,N_19020);
and U19767 (N_19767,N_19340,N_19092);
xnor U19768 (N_19768,N_18767,N_19288);
and U19769 (N_19769,N_19123,N_19057);
nand U19770 (N_19770,N_18868,N_19015);
nor U19771 (N_19771,N_19070,N_18924);
and U19772 (N_19772,N_19331,N_19340);
or U19773 (N_19773,N_18920,N_19193);
nand U19774 (N_19774,N_19151,N_18936);
nor U19775 (N_19775,N_18964,N_19019);
or U19776 (N_19776,N_19079,N_19150);
xor U19777 (N_19777,N_19367,N_18841);
and U19778 (N_19778,N_19101,N_19100);
nor U19779 (N_19779,N_18928,N_18865);
and U19780 (N_19780,N_18835,N_19048);
nor U19781 (N_19781,N_19133,N_18990);
nor U19782 (N_19782,N_19257,N_18843);
or U19783 (N_19783,N_19118,N_19135);
and U19784 (N_19784,N_19058,N_19010);
xnor U19785 (N_19785,N_18931,N_19085);
and U19786 (N_19786,N_19329,N_18767);
nor U19787 (N_19787,N_18912,N_19223);
nand U19788 (N_19788,N_19030,N_19227);
nor U19789 (N_19789,N_19227,N_18871);
nand U19790 (N_19790,N_18837,N_18898);
and U19791 (N_19791,N_19149,N_19043);
xor U19792 (N_19792,N_18849,N_19227);
and U19793 (N_19793,N_19224,N_19033);
or U19794 (N_19794,N_18989,N_18823);
and U19795 (N_19795,N_19173,N_19018);
or U19796 (N_19796,N_19125,N_19369);
nand U19797 (N_19797,N_18946,N_19030);
xnor U19798 (N_19798,N_19004,N_19280);
or U19799 (N_19799,N_19353,N_19159);
nor U19800 (N_19800,N_19315,N_18877);
or U19801 (N_19801,N_18890,N_18768);
or U19802 (N_19802,N_19197,N_19282);
nand U19803 (N_19803,N_19320,N_18883);
nor U19804 (N_19804,N_18790,N_19274);
or U19805 (N_19805,N_19345,N_19123);
or U19806 (N_19806,N_18833,N_18897);
nor U19807 (N_19807,N_19051,N_19296);
xnor U19808 (N_19808,N_19144,N_19335);
nand U19809 (N_19809,N_18799,N_18950);
nor U19810 (N_19810,N_19212,N_19039);
and U19811 (N_19811,N_19094,N_19154);
and U19812 (N_19812,N_19132,N_18822);
nor U19813 (N_19813,N_19283,N_18979);
xnor U19814 (N_19814,N_18958,N_19185);
nor U19815 (N_19815,N_19204,N_19273);
nor U19816 (N_19816,N_19194,N_19222);
or U19817 (N_19817,N_19212,N_18821);
nor U19818 (N_19818,N_19142,N_19335);
and U19819 (N_19819,N_18829,N_18958);
nand U19820 (N_19820,N_19014,N_18776);
and U19821 (N_19821,N_19207,N_18759);
or U19822 (N_19822,N_18885,N_19050);
nor U19823 (N_19823,N_19182,N_19186);
xnor U19824 (N_19824,N_18753,N_18871);
nor U19825 (N_19825,N_19361,N_19139);
nand U19826 (N_19826,N_19224,N_19188);
nor U19827 (N_19827,N_19143,N_19211);
and U19828 (N_19828,N_19252,N_18857);
and U19829 (N_19829,N_18886,N_18787);
and U19830 (N_19830,N_19301,N_19003);
and U19831 (N_19831,N_18939,N_18804);
nand U19832 (N_19832,N_19314,N_19284);
xnor U19833 (N_19833,N_18951,N_18928);
nor U19834 (N_19834,N_19163,N_19345);
or U19835 (N_19835,N_19354,N_18903);
nor U19836 (N_19836,N_18766,N_18854);
or U19837 (N_19837,N_19265,N_18825);
nor U19838 (N_19838,N_19110,N_19181);
and U19839 (N_19839,N_19117,N_19347);
and U19840 (N_19840,N_19355,N_18824);
xor U19841 (N_19841,N_19035,N_18858);
nand U19842 (N_19842,N_18889,N_19098);
and U19843 (N_19843,N_19116,N_19149);
xnor U19844 (N_19844,N_18841,N_19136);
or U19845 (N_19845,N_18999,N_18979);
or U19846 (N_19846,N_18885,N_19227);
nor U19847 (N_19847,N_19118,N_18885);
and U19848 (N_19848,N_19094,N_19044);
or U19849 (N_19849,N_19124,N_18867);
xor U19850 (N_19850,N_19051,N_19127);
and U19851 (N_19851,N_19354,N_19213);
nor U19852 (N_19852,N_18870,N_18904);
nand U19853 (N_19853,N_18848,N_18923);
nor U19854 (N_19854,N_18960,N_19322);
xnor U19855 (N_19855,N_19196,N_19237);
or U19856 (N_19856,N_19220,N_19286);
nor U19857 (N_19857,N_19053,N_18917);
nand U19858 (N_19858,N_19006,N_19355);
nor U19859 (N_19859,N_19348,N_19328);
nand U19860 (N_19860,N_19195,N_18865);
and U19861 (N_19861,N_18806,N_19217);
nor U19862 (N_19862,N_19275,N_18860);
or U19863 (N_19863,N_18866,N_19249);
or U19864 (N_19864,N_19367,N_19306);
nor U19865 (N_19865,N_18881,N_18775);
nand U19866 (N_19866,N_19361,N_19255);
nor U19867 (N_19867,N_19150,N_18779);
and U19868 (N_19868,N_18986,N_19149);
xor U19869 (N_19869,N_19119,N_18912);
nand U19870 (N_19870,N_18783,N_19243);
and U19871 (N_19871,N_18908,N_18859);
or U19872 (N_19872,N_18831,N_19341);
xor U19873 (N_19873,N_18953,N_18976);
nor U19874 (N_19874,N_19001,N_18860);
and U19875 (N_19875,N_19182,N_18844);
or U19876 (N_19876,N_19174,N_19345);
nor U19877 (N_19877,N_19277,N_19184);
and U19878 (N_19878,N_18770,N_18759);
nand U19879 (N_19879,N_19190,N_18776);
and U19880 (N_19880,N_18846,N_19362);
and U19881 (N_19881,N_18820,N_19062);
xor U19882 (N_19882,N_18931,N_19328);
nand U19883 (N_19883,N_18783,N_18977);
nand U19884 (N_19884,N_19078,N_19324);
nand U19885 (N_19885,N_18760,N_19241);
nor U19886 (N_19886,N_19233,N_19125);
and U19887 (N_19887,N_19161,N_19088);
nand U19888 (N_19888,N_19118,N_18896);
or U19889 (N_19889,N_18877,N_19073);
nor U19890 (N_19890,N_19155,N_18842);
and U19891 (N_19891,N_18874,N_19141);
and U19892 (N_19892,N_18830,N_19341);
and U19893 (N_19893,N_19155,N_18775);
xnor U19894 (N_19894,N_18932,N_19168);
nand U19895 (N_19895,N_18783,N_19199);
xnor U19896 (N_19896,N_19372,N_19243);
nor U19897 (N_19897,N_19311,N_19142);
xor U19898 (N_19898,N_18789,N_19024);
xor U19899 (N_19899,N_19103,N_19248);
nand U19900 (N_19900,N_19326,N_19010);
xnor U19901 (N_19901,N_18915,N_19284);
and U19902 (N_19902,N_19206,N_18884);
nand U19903 (N_19903,N_19111,N_19370);
nor U19904 (N_19904,N_19337,N_18967);
xor U19905 (N_19905,N_19156,N_19036);
and U19906 (N_19906,N_19203,N_18781);
nand U19907 (N_19907,N_19162,N_19275);
nand U19908 (N_19908,N_18990,N_18982);
xnor U19909 (N_19909,N_18993,N_19117);
nor U19910 (N_19910,N_18985,N_19013);
or U19911 (N_19911,N_19011,N_18910);
nand U19912 (N_19912,N_19321,N_18994);
and U19913 (N_19913,N_18758,N_19290);
nand U19914 (N_19914,N_18767,N_18774);
nand U19915 (N_19915,N_19143,N_19349);
nand U19916 (N_19916,N_18833,N_19156);
nand U19917 (N_19917,N_18976,N_18989);
and U19918 (N_19918,N_19363,N_19063);
or U19919 (N_19919,N_19133,N_19241);
xnor U19920 (N_19920,N_18917,N_18925);
nor U19921 (N_19921,N_19353,N_18840);
nand U19922 (N_19922,N_19107,N_18826);
nor U19923 (N_19923,N_19287,N_18769);
or U19924 (N_19924,N_19109,N_19212);
and U19925 (N_19925,N_19047,N_19194);
nor U19926 (N_19926,N_18869,N_18953);
xnor U19927 (N_19927,N_19115,N_19110);
nor U19928 (N_19928,N_19175,N_18897);
and U19929 (N_19929,N_18780,N_18801);
or U19930 (N_19930,N_19216,N_19136);
and U19931 (N_19931,N_19372,N_18866);
nor U19932 (N_19932,N_19185,N_19368);
or U19933 (N_19933,N_18957,N_19038);
nor U19934 (N_19934,N_18980,N_19221);
xor U19935 (N_19935,N_18826,N_18796);
nand U19936 (N_19936,N_18783,N_18921);
and U19937 (N_19937,N_18867,N_18841);
or U19938 (N_19938,N_18961,N_18969);
nand U19939 (N_19939,N_19218,N_18913);
and U19940 (N_19940,N_19300,N_19189);
or U19941 (N_19941,N_19184,N_18952);
xnor U19942 (N_19942,N_18839,N_18927);
and U19943 (N_19943,N_18922,N_19264);
or U19944 (N_19944,N_18916,N_19256);
xnor U19945 (N_19945,N_19131,N_19141);
or U19946 (N_19946,N_19361,N_18884);
nand U19947 (N_19947,N_19166,N_18899);
and U19948 (N_19948,N_19324,N_19218);
nand U19949 (N_19949,N_18923,N_19269);
nor U19950 (N_19950,N_19210,N_18843);
or U19951 (N_19951,N_19284,N_19288);
xnor U19952 (N_19952,N_19350,N_19089);
xnor U19953 (N_19953,N_19020,N_19294);
nand U19954 (N_19954,N_18808,N_19218);
nor U19955 (N_19955,N_19354,N_19283);
or U19956 (N_19956,N_19115,N_18779);
or U19957 (N_19957,N_19040,N_18789);
nor U19958 (N_19958,N_19154,N_18900);
or U19959 (N_19959,N_18995,N_19109);
xnor U19960 (N_19960,N_18779,N_18789);
nand U19961 (N_19961,N_18927,N_19085);
xnor U19962 (N_19962,N_19284,N_18840);
or U19963 (N_19963,N_18946,N_18802);
nor U19964 (N_19964,N_18919,N_18913);
or U19965 (N_19965,N_19011,N_19324);
nor U19966 (N_19966,N_19260,N_18918);
or U19967 (N_19967,N_19021,N_18924);
and U19968 (N_19968,N_18909,N_18802);
or U19969 (N_19969,N_18993,N_19283);
and U19970 (N_19970,N_19159,N_19069);
nand U19971 (N_19971,N_19333,N_18993);
nand U19972 (N_19972,N_19292,N_19187);
nor U19973 (N_19973,N_18942,N_19073);
nand U19974 (N_19974,N_19128,N_19102);
nand U19975 (N_19975,N_19283,N_19151);
and U19976 (N_19976,N_18897,N_19034);
or U19977 (N_19977,N_18826,N_19289);
xnor U19978 (N_19978,N_18878,N_19184);
nor U19979 (N_19979,N_19093,N_18783);
and U19980 (N_19980,N_18874,N_18933);
or U19981 (N_19981,N_19336,N_18884);
nor U19982 (N_19982,N_19313,N_19252);
nor U19983 (N_19983,N_19345,N_18843);
nor U19984 (N_19984,N_18828,N_19189);
xor U19985 (N_19985,N_19322,N_18802);
and U19986 (N_19986,N_18967,N_19022);
nand U19987 (N_19987,N_19344,N_19187);
nor U19988 (N_19988,N_18831,N_18963);
nand U19989 (N_19989,N_18798,N_18931);
nor U19990 (N_19990,N_18980,N_18848);
nor U19991 (N_19991,N_18771,N_19346);
and U19992 (N_19992,N_19184,N_19198);
xor U19993 (N_19993,N_18829,N_19134);
nor U19994 (N_19994,N_18941,N_19115);
or U19995 (N_19995,N_19003,N_19164);
and U19996 (N_19996,N_19350,N_18823);
xor U19997 (N_19997,N_19048,N_18934);
or U19998 (N_19998,N_18831,N_19312);
xor U19999 (N_19999,N_18751,N_19052);
nor U20000 (N_20000,N_19741,N_19436);
nand U20001 (N_20001,N_19554,N_19932);
or U20002 (N_20002,N_19731,N_19886);
and U20003 (N_20003,N_19530,N_19552);
or U20004 (N_20004,N_19508,N_19405);
nand U20005 (N_20005,N_19446,N_19671);
nand U20006 (N_20006,N_19846,N_19420);
and U20007 (N_20007,N_19912,N_19401);
xor U20008 (N_20008,N_19953,N_19520);
xor U20009 (N_20009,N_19510,N_19557);
nor U20010 (N_20010,N_19475,N_19945);
xnor U20011 (N_20011,N_19704,N_19667);
xor U20012 (N_20012,N_19744,N_19491);
and U20013 (N_20013,N_19639,N_19551);
nor U20014 (N_20014,N_19974,N_19860);
nor U20015 (N_20015,N_19455,N_19934);
nor U20016 (N_20016,N_19394,N_19440);
xor U20017 (N_20017,N_19655,N_19687);
and U20018 (N_20018,N_19740,N_19644);
nand U20019 (N_20019,N_19636,N_19747);
nand U20020 (N_20020,N_19688,N_19449);
nor U20021 (N_20021,N_19398,N_19765);
nor U20022 (N_20022,N_19409,N_19489);
nor U20023 (N_20023,N_19638,N_19656);
nor U20024 (N_20024,N_19493,N_19997);
nand U20025 (N_20025,N_19385,N_19916);
nor U20026 (N_20026,N_19940,N_19481);
nand U20027 (N_20027,N_19939,N_19597);
or U20028 (N_20028,N_19676,N_19534);
nand U20029 (N_20029,N_19710,N_19992);
nor U20030 (N_20030,N_19877,N_19894);
or U20031 (N_20031,N_19701,N_19715);
xor U20032 (N_20032,N_19790,N_19458);
xor U20033 (N_20033,N_19680,N_19730);
xor U20034 (N_20034,N_19463,N_19649);
xor U20035 (N_20035,N_19544,N_19852);
and U20036 (N_20036,N_19388,N_19505);
nor U20037 (N_20037,N_19907,N_19482);
and U20038 (N_20038,N_19926,N_19573);
nor U20039 (N_20039,N_19819,N_19439);
or U20040 (N_20040,N_19654,N_19660);
xnor U20041 (N_20041,N_19470,N_19466);
nor U20042 (N_20042,N_19393,N_19820);
nor U20043 (N_20043,N_19679,N_19626);
or U20044 (N_20044,N_19523,N_19836);
nand U20045 (N_20045,N_19959,N_19700);
and U20046 (N_20046,N_19615,N_19514);
nand U20047 (N_20047,N_19996,N_19539);
or U20048 (N_20048,N_19981,N_19706);
xnor U20049 (N_20049,N_19979,N_19998);
nand U20050 (N_20050,N_19961,N_19856);
nor U20051 (N_20051,N_19471,N_19522);
nor U20052 (N_20052,N_19631,N_19788);
or U20053 (N_20053,N_19578,N_19468);
nand U20054 (N_20054,N_19814,N_19910);
nand U20055 (N_20055,N_19770,N_19702);
or U20056 (N_20056,N_19418,N_19600);
and U20057 (N_20057,N_19492,N_19445);
xnor U20058 (N_20058,N_19991,N_19891);
or U20059 (N_20059,N_19579,N_19598);
and U20060 (N_20060,N_19397,N_19708);
nor U20061 (N_20061,N_19748,N_19768);
nand U20062 (N_20062,N_19457,N_19434);
nand U20063 (N_20063,N_19919,N_19947);
nand U20064 (N_20064,N_19927,N_19777);
xnor U20065 (N_20065,N_19794,N_19812);
nand U20066 (N_20066,N_19875,N_19461);
nand U20067 (N_20067,N_19750,N_19561);
nand U20068 (N_20068,N_19862,N_19586);
nor U20069 (N_20069,N_19432,N_19593);
xor U20070 (N_20070,N_19456,N_19414);
and U20071 (N_20071,N_19925,N_19601);
nor U20072 (N_20072,N_19735,N_19413);
and U20073 (N_20073,N_19901,N_19973);
nor U20074 (N_20074,N_19848,N_19538);
or U20075 (N_20075,N_19640,N_19835);
nor U20076 (N_20076,N_19724,N_19437);
xnor U20077 (N_20077,N_19435,N_19904);
xor U20078 (N_20078,N_19751,N_19664);
nor U20079 (N_20079,N_19576,N_19659);
nor U20080 (N_20080,N_19563,N_19646);
and U20081 (N_20081,N_19823,N_19892);
nor U20082 (N_20082,N_19698,N_19635);
nor U20083 (N_20083,N_19567,N_19876);
and U20084 (N_20084,N_19645,N_19592);
nor U20085 (N_20085,N_19525,N_19766);
and U20086 (N_20086,N_19696,N_19666);
nor U20087 (N_20087,N_19949,N_19427);
and U20088 (N_20088,N_19588,N_19911);
xnor U20089 (N_20089,N_19753,N_19757);
or U20090 (N_20090,N_19506,N_19462);
nor U20091 (N_20091,N_19728,N_19537);
xor U20092 (N_20092,N_19851,N_19982);
and U20093 (N_20093,N_19454,N_19569);
or U20094 (N_20094,N_19970,N_19617);
and U20095 (N_20095,N_19692,N_19411);
nor U20096 (N_20096,N_19827,N_19575);
or U20097 (N_20097,N_19408,N_19494);
xor U20098 (N_20098,N_19375,N_19758);
xor U20099 (N_20099,N_19989,N_19499);
xor U20100 (N_20100,N_19976,N_19995);
or U20101 (N_20101,N_19738,N_19853);
nor U20102 (N_20102,N_19786,N_19697);
or U20103 (N_20103,N_19783,N_19611);
nand U20104 (N_20104,N_19746,N_19968);
or U20105 (N_20105,N_19616,N_19389);
nor U20106 (N_20106,N_19477,N_19651);
and U20107 (N_20107,N_19769,N_19625);
xnor U20108 (N_20108,N_19521,N_19921);
or U20109 (N_20109,N_19450,N_19821);
and U20110 (N_20110,N_19899,N_19859);
or U20111 (N_20111,N_19464,N_19583);
and U20112 (N_20112,N_19906,N_19864);
xnor U20113 (N_20113,N_19969,N_19825);
nand U20114 (N_20114,N_19683,N_19942);
xnor U20115 (N_20115,N_19548,N_19716);
xnor U20116 (N_20116,N_19399,N_19718);
xnor U20117 (N_20117,N_19412,N_19599);
and U20118 (N_20118,N_19721,N_19516);
nor U20119 (N_20119,N_19867,N_19971);
xnor U20120 (N_20120,N_19960,N_19818);
xor U20121 (N_20121,N_19791,N_19884);
xnor U20122 (N_20122,N_19465,N_19422);
nand U20123 (N_20123,N_19668,N_19734);
and U20124 (N_20124,N_19869,N_19447);
nor U20125 (N_20125,N_19632,N_19605);
or U20126 (N_20126,N_19870,N_19778);
and U20127 (N_20127,N_19620,N_19882);
xor U20128 (N_20128,N_19382,N_19681);
or U20129 (N_20129,N_19580,N_19661);
nor U20130 (N_20130,N_19547,N_19784);
or U20131 (N_20131,N_19951,N_19518);
xor U20132 (N_20132,N_19496,N_19903);
or U20133 (N_20133,N_19533,N_19383);
nand U20134 (N_20134,N_19379,N_19603);
and U20135 (N_20135,N_19587,N_19444);
or U20136 (N_20136,N_19653,N_19406);
xor U20137 (N_20137,N_19801,N_19665);
nor U20138 (N_20138,N_19650,N_19866);
nand U20139 (N_20139,N_19880,N_19441);
nor U20140 (N_20140,N_19905,N_19936);
nor U20141 (N_20141,N_19829,N_19990);
and U20142 (N_20142,N_19381,N_19658);
or U20143 (N_20143,N_19817,N_19808);
nand U20144 (N_20144,N_19485,N_19871);
or U20145 (N_20145,N_19967,N_19419);
nor U20146 (N_20146,N_19570,N_19811);
nor U20147 (N_20147,N_19944,N_19752);
or U20148 (N_20148,N_19608,N_19924);
nand U20149 (N_20149,N_19923,N_19562);
nor U20150 (N_20150,N_19623,N_19781);
nor U20151 (N_20151,N_19429,N_19622);
nand U20152 (N_20152,N_19527,N_19602);
and U20153 (N_20153,N_19802,N_19725);
nand U20154 (N_20154,N_19670,N_19713);
nand U20155 (N_20155,N_19749,N_19805);
nor U20156 (N_20156,N_19994,N_19965);
and U20157 (N_20157,N_19930,N_19705);
xnor U20158 (N_20158,N_19931,N_19536);
nand U20159 (N_20159,N_19610,N_19678);
nor U20160 (N_20160,N_19415,N_19502);
nand U20161 (N_20161,N_19963,N_19540);
nor U20162 (N_20162,N_19943,N_19815);
xor U20163 (N_20163,N_19543,N_19722);
nor U20164 (N_20164,N_19596,N_19428);
and U20165 (N_20165,N_19984,N_19855);
xor U20166 (N_20166,N_19800,N_19488);
and U20167 (N_20167,N_19918,N_19684);
or U20168 (N_20168,N_19675,N_19776);
and U20169 (N_20169,N_19633,N_19643);
and U20170 (N_20170,N_19830,N_19797);
xnor U20171 (N_20171,N_19621,N_19542);
nand U20172 (N_20172,N_19377,N_19809);
or U20173 (N_20173,N_19822,N_19614);
nand U20174 (N_20174,N_19560,N_19535);
xor U20175 (N_20175,N_19619,N_19785);
nor U20176 (N_20176,N_19709,N_19759);
or U20177 (N_20177,N_19952,N_19396);
or U20178 (N_20178,N_19513,N_19630);
and U20179 (N_20179,N_19528,N_19555);
xnor U20180 (N_20180,N_19553,N_19495);
and U20181 (N_20181,N_19400,N_19452);
and U20182 (N_20182,N_19714,N_19885);
and U20183 (N_20183,N_19849,N_19736);
and U20184 (N_20184,N_19410,N_19694);
nor U20185 (N_20185,N_19648,N_19727);
nor U20186 (N_20186,N_19972,N_19693);
or U20187 (N_20187,N_19566,N_19854);
xnor U20188 (N_20188,N_19574,N_19423);
or U20189 (N_20189,N_19985,N_19908);
nor U20190 (N_20190,N_19469,N_19888);
nor U20191 (N_20191,N_19711,N_19386);
xor U20192 (N_20192,N_19690,N_19545);
xnor U20193 (N_20193,N_19629,N_19980);
xnor U20194 (N_20194,N_19799,N_19816);
nor U20195 (N_20195,N_19824,N_19472);
nor U20196 (N_20196,N_19798,N_19928);
xor U20197 (N_20197,N_19498,N_19568);
and U20198 (N_20198,N_19433,N_19913);
and U20199 (N_20199,N_19473,N_19417);
or U20200 (N_20200,N_19430,N_19954);
or U20201 (N_20201,N_19612,N_19425);
xnor U20202 (N_20202,N_19917,N_19662);
nor U20203 (N_20203,N_19890,N_19507);
or U20204 (N_20204,N_19938,N_19509);
and U20205 (N_20205,N_19685,N_19443);
nand U20206 (N_20206,N_19832,N_19390);
nor U20207 (N_20207,N_19958,N_19863);
nor U20208 (N_20208,N_19881,N_19448);
or U20209 (N_20209,N_19889,N_19564);
and U20210 (N_20210,N_19459,N_19873);
nor U20211 (N_20211,N_19618,N_19672);
nor U20212 (N_20212,N_19691,N_19789);
xnor U20213 (N_20213,N_19402,N_19395);
nor U20214 (N_20214,N_19519,N_19515);
and U20215 (N_20215,N_19837,N_19609);
nor U20216 (N_20216,N_19594,N_19460);
nor U20217 (N_20217,N_19500,N_19893);
and U20218 (N_20218,N_19966,N_19442);
nand U20219 (N_20219,N_19842,N_19754);
or U20220 (N_20220,N_19627,N_19843);
and U20221 (N_20221,N_19977,N_19577);
nor U20222 (N_20222,N_19703,N_19868);
and U20223 (N_20223,N_19673,N_19946);
xor U20224 (N_20224,N_19589,N_19421);
nand U20225 (N_20225,N_19792,N_19806);
nor U20226 (N_20226,N_19717,N_19733);
nor U20227 (N_20227,N_19787,N_19699);
and U20228 (N_20228,N_19529,N_19581);
nor U20229 (N_20229,N_19857,N_19807);
and U20230 (N_20230,N_19779,N_19773);
or U20231 (N_20231,N_19831,N_19501);
or U20232 (N_20232,N_19865,N_19915);
and U20233 (N_20233,N_19795,N_19376);
or U20234 (N_20234,N_19761,N_19490);
xnor U20235 (N_20235,N_19504,N_19745);
or U20236 (N_20236,N_19756,N_19771);
nand U20237 (N_20237,N_19426,N_19503);
nor U20238 (N_20238,N_19541,N_19935);
xnor U20239 (N_20239,N_19484,N_19767);
nand U20240 (N_20240,N_19511,N_19955);
nor U20241 (N_20241,N_19641,N_19604);
and U20242 (N_20242,N_19719,N_19378);
nand U20243 (N_20243,N_19556,N_19590);
nand U20244 (N_20244,N_19897,N_19483);
or U20245 (N_20245,N_19909,N_19652);
or U20246 (N_20246,N_19898,N_19760);
nand U20247 (N_20247,N_19978,N_19595);
and U20248 (N_20248,N_19833,N_19526);
xnor U20249 (N_20249,N_19391,N_19392);
xnor U20250 (N_20250,N_19531,N_19642);
nand U20251 (N_20251,N_19387,N_19956);
nor U20252 (N_20252,N_19780,N_19828);
xnor U20253 (N_20253,N_19613,N_19826);
nor U20254 (N_20254,N_19607,N_19571);
and U20255 (N_20255,N_19624,N_19732);
nor U20256 (N_20256,N_19764,N_19582);
nor U20257 (N_20257,N_19486,N_19565);
xor U20258 (N_20258,N_19872,N_19993);
nand U20259 (N_20259,N_19845,N_19637);
nor U20260 (N_20260,N_19686,N_19782);
nand U20261 (N_20261,N_19920,N_19878);
or U20262 (N_20262,N_19657,N_19712);
xnor U20263 (N_20263,N_19847,N_19663);
xor U20264 (N_20264,N_19737,N_19723);
or U20265 (N_20265,N_19585,N_19677);
xor U20266 (N_20266,N_19900,N_19839);
nand U20267 (N_20267,N_19743,N_19532);
and U20268 (N_20268,N_19850,N_19497);
xnor U20269 (N_20269,N_19838,N_19775);
nand U20270 (N_20270,N_19606,N_19480);
xnor U20271 (N_20271,N_19707,N_19810);
nor U20272 (N_20272,N_19479,N_19803);
nand U20273 (N_20273,N_19550,N_19695);
or U20274 (N_20274,N_19933,N_19524);
and U20275 (N_20275,N_19558,N_19742);
and U20276 (N_20276,N_19772,N_19902);
nand U20277 (N_20277,N_19813,N_19431);
nand U20278 (N_20278,N_19796,N_19755);
nor U20279 (N_20279,N_19975,N_19879);
or U20280 (N_20280,N_19762,N_19874);
nor U20281 (N_20281,N_19957,N_19986);
nand U20282 (N_20282,N_19929,N_19840);
nand U20283 (N_20283,N_19999,N_19720);
xor U20284 (N_20284,N_19467,N_19517);
xor U20285 (N_20285,N_19844,N_19962);
and U20286 (N_20286,N_19987,N_19669);
nor U20287 (N_20287,N_19407,N_19634);
and U20288 (N_20288,N_19937,N_19726);
xnor U20289 (N_20289,N_19559,N_19451);
or U20290 (N_20290,N_19438,N_19988);
nor U20291 (N_20291,N_19834,N_19883);
or U20292 (N_20292,N_19478,N_19964);
or U20293 (N_20293,N_19424,N_19549);
nand U20294 (N_20294,N_19922,N_19572);
nor U20295 (N_20295,N_19896,N_19841);
nor U20296 (N_20296,N_19948,N_19474);
xnor U20297 (N_20297,N_19941,N_19453);
nand U20298 (N_20298,N_19476,N_19380);
or U20299 (N_20299,N_19914,N_19682);
and U20300 (N_20300,N_19858,N_19416);
nor U20301 (N_20301,N_19861,N_19774);
and U20302 (N_20302,N_19403,N_19546);
and U20303 (N_20303,N_19674,N_19950);
nand U20304 (N_20304,N_19729,N_19887);
or U20305 (N_20305,N_19487,N_19628);
xor U20306 (N_20306,N_19584,N_19804);
xor U20307 (N_20307,N_19647,N_19512);
nor U20308 (N_20308,N_19384,N_19895);
nand U20309 (N_20309,N_19983,N_19404);
xnor U20310 (N_20310,N_19793,N_19763);
nor U20311 (N_20311,N_19591,N_19689);
and U20312 (N_20312,N_19739,N_19915);
nand U20313 (N_20313,N_19636,N_19384);
nand U20314 (N_20314,N_19686,N_19669);
nand U20315 (N_20315,N_19718,N_19407);
nor U20316 (N_20316,N_19575,N_19905);
or U20317 (N_20317,N_19966,N_19769);
nor U20318 (N_20318,N_19760,N_19922);
xor U20319 (N_20319,N_19476,N_19525);
nand U20320 (N_20320,N_19942,N_19633);
xor U20321 (N_20321,N_19503,N_19597);
or U20322 (N_20322,N_19693,N_19629);
xor U20323 (N_20323,N_19411,N_19834);
and U20324 (N_20324,N_19480,N_19464);
or U20325 (N_20325,N_19622,N_19402);
nand U20326 (N_20326,N_19902,N_19480);
and U20327 (N_20327,N_19817,N_19378);
or U20328 (N_20328,N_19956,N_19624);
or U20329 (N_20329,N_19615,N_19440);
nor U20330 (N_20330,N_19718,N_19834);
or U20331 (N_20331,N_19761,N_19469);
nand U20332 (N_20332,N_19424,N_19381);
and U20333 (N_20333,N_19460,N_19938);
nor U20334 (N_20334,N_19802,N_19439);
nand U20335 (N_20335,N_19882,N_19524);
nor U20336 (N_20336,N_19826,N_19649);
nor U20337 (N_20337,N_19457,N_19405);
nand U20338 (N_20338,N_19927,N_19976);
or U20339 (N_20339,N_19799,N_19423);
and U20340 (N_20340,N_19755,N_19764);
nor U20341 (N_20341,N_19759,N_19874);
nor U20342 (N_20342,N_19639,N_19676);
nand U20343 (N_20343,N_19992,N_19775);
or U20344 (N_20344,N_19579,N_19541);
and U20345 (N_20345,N_19677,N_19479);
nand U20346 (N_20346,N_19981,N_19805);
xor U20347 (N_20347,N_19895,N_19992);
and U20348 (N_20348,N_19917,N_19684);
nand U20349 (N_20349,N_19978,N_19791);
and U20350 (N_20350,N_19468,N_19908);
or U20351 (N_20351,N_19443,N_19835);
nor U20352 (N_20352,N_19944,N_19623);
xor U20353 (N_20353,N_19480,N_19776);
and U20354 (N_20354,N_19992,N_19973);
nand U20355 (N_20355,N_19703,N_19977);
or U20356 (N_20356,N_19591,N_19432);
or U20357 (N_20357,N_19804,N_19438);
xnor U20358 (N_20358,N_19633,N_19993);
or U20359 (N_20359,N_19703,N_19748);
xor U20360 (N_20360,N_19893,N_19918);
or U20361 (N_20361,N_19818,N_19718);
xnor U20362 (N_20362,N_19525,N_19986);
or U20363 (N_20363,N_19772,N_19578);
and U20364 (N_20364,N_19428,N_19535);
and U20365 (N_20365,N_19502,N_19776);
nor U20366 (N_20366,N_19758,N_19558);
xnor U20367 (N_20367,N_19935,N_19996);
or U20368 (N_20368,N_19951,N_19917);
nand U20369 (N_20369,N_19973,N_19938);
nor U20370 (N_20370,N_19990,N_19982);
or U20371 (N_20371,N_19406,N_19610);
nor U20372 (N_20372,N_19905,N_19705);
and U20373 (N_20373,N_19601,N_19693);
nor U20374 (N_20374,N_19603,N_19894);
xnor U20375 (N_20375,N_19934,N_19991);
and U20376 (N_20376,N_19461,N_19904);
and U20377 (N_20377,N_19393,N_19456);
nor U20378 (N_20378,N_19621,N_19619);
nor U20379 (N_20379,N_19583,N_19810);
nor U20380 (N_20380,N_19419,N_19534);
and U20381 (N_20381,N_19900,N_19652);
and U20382 (N_20382,N_19607,N_19715);
or U20383 (N_20383,N_19830,N_19507);
nand U20384 (N_20384,N_19641,N_19937);
xor U20385 (N_20385,N_19744,N_19702);
xor U20386 (N_20386,N_19385,N_19631);
and U20387 (N_20387,N_19846,N_19422);
and U20388 (N_20388,N_19551,N_19416);
nor U20389 (N_20389,N_19995,N_19503);
nand U20390 (N_20390,N_19981,N_19734);
and U20391 (N_20391,N_19985,N_19917);
or U20392 (N_20392,N_19687,N_19381);
and U20393 (N_20393,N_19445,N_19588);
and U20394 (N_20394,N_19548,N_19661);
or U20395 (N_20395,N_19784,N_19651);
xnor U20396 (N_20396,N_19435,N_19697);
and U20397 (N_20397,N_19485,N_19583);
nand U20398 (N_20398,N_19423,N_19835);
xor U20399 (N_20399,N_19559,N_19594);
nor U20400 (N_20400,N_19453,N_19875);
xnor U20401 (N_20401,N_19960,N_19388);
xor U20402 (N_20402,N_19632,N_19956);
xnor U20403 (N_20403,N_19556,N_19455);
nor U20404 (N_20404,N_19407,N_19440);
or U20405 (N_20405,N_19666,N_19760);
or U20406 (N_20406,N_19740,N_19689);
nand U20407 (N_20407,N_19966,N_19975);
xnor U20408 (N_20408,N_19503,N_19789);
and U20409 (N_20409,N_19696,N_19932);
nand U20410 (N_20410,N_19999,N_19519);
nand U20411 (N_20411,N_19399,N_19685);
or U20412 (N_20412,N_19427,N_19799);
xnor U20413 (N_20413,N_19771,N_19858);
and U20414 (N_20414,N_19488,N_19876);
and U20415 (N_20415,N_19638,N_19451);
nor U20416 (N_20416,N_19918,N_19872);
nand U20417 (N_20417,N_19881,N_19861);
nor U20418 (N_20418,N_19876,N_19746);
or U20419 (N_20419,N_19962,N_19389);
and U20420 (N_20420,N_19691,N_19867);
nor U20421 (N_20421,N_19432,N_19466);
or U20422 (N_20422,N_19521,N_19568);
nor U20423 (N_20423,N_19987,N_19481);
and U20424 (N_20424,N_19807,N_19930);
and U20425 (N_20425,N_19784,N_19729);
xor U20426 (N_20426,N_19375,N_19508);
xnor U20427 (N_20427,N_19575,N_19881);
and U20428 (N_20428,N_19909,N_19595);
xnor U20429 (N_20429,N_19805,N_19688);
or U20430 (N_20430,N_19422,N_19887);
or U20431 (N_20431,N_19594,N_19824);
nand U20432 (N_20432,N_19843,N_19857);
nand U20433 (N_20433,N_19734,N_19935);
xor U20434 (N_20434,N_19725,N_19428);
nor U20435 (N_20435,N_19483,N_19528);
nor U20436 (N_20436,N_19797,N_19527);
or U20437 (N_20437,N_19386,N_19501);
nor U20438 (N_20438,N_19867,N_19877);
nor U20439 (N_20439,N_19665,N_19435);
or U20440 (N_20440,N_19533,N_19617);
nand U20441 (N_20441,N_19611,N_19440);
and U20442 (N_20442,N_19648,N_19564);
and U20443 (N_20443,N_19770,N_19994);
and U20444 (N_20444,N_19999,N_19920);
nand U20445 (N_20445,N_19872,N_19543);
xnor U20446 (N_20446,N_19911,N_19908);
or U20447 (N_20447,N_19870,N_19481);
nor U20448 (N_20448,N_19417,N_19549);
or U20449 (N_20449,N_19727,N_19719);
or U20450 (N_20450,N_19475,N_19454);
and U20451 (N_20451,N_19431,N_19843);
nand U20452 (N_20452,N_19405,N_19487);
nand U20453 (N_20453,N_19516,N_19540);
nand U20454 (N_20454,N_19533,N_19817);
nand U20455 (N_20455,N_19946,N_19456);
nand U20456 (N_20456,N_19751,N_19818);
xnor U20457 (N_20457,N_19839,N_19462);
xor U20458 (N_20458,N_19441,N_19994);
xnor U20459 (N_20459,N_19689,N_19972);
and U20460 (N_20460,N_19376,N_19892);
nor U20461 (N_20461,N_19430,N_19730);
or U20462 (N_20462,N_19603,N_19948);
or U20463 (N_20463,N_19730,N_19581);
xor U20464 (N_20464,N_19559,N_19381);
xnor U20465 (N_20465,N_19573,N_19622);
xor U20466 (N_20466,N_19380,N_19784);
and U20467 (N_20467,N_19774,N_19710);
nor U20468 (N_20468,N_19995,N_19449);
or U20469 (N_20469,N_19494,N_19853);
and U20470 (N_20470,N_19845,N_19995);
and U20471 (N_20471,N_19446,N_19462);
or U20472 (N_20472,N_19727,N_19726);
and U20473 (N_20473,N_19681,N_19590);
and U20474 (N_20474,N_19897,N_19646);
xor U20475 (N_20475,N_19956,N_19527);
and U20476 (N_20476,N_19555,N_19393);
nor U20477 (N_20477,N_19391,N_19917);
xnor U20478 (N_20478,N_19624,N_19379);
nand U20479 (N_20479,N_19879,N_19961);
nor U20480 (N_20480,N_19376,N_19377);
xnor U20481 (N_20481,N_19792,N_19699);
nand U20482 (N_20482,N_19537,N_19414);
and U20483 (N_20483,N_19530,N_19541);
xnor U20484 (N_20484,N_19472,N_19389);
or U20485 (N_20485,N_19490,N_19558);
nor U20486 (N_20486,N_19939,N_19887);
and U20487 (N_20487,N_19394,N_19526);
nand U20488 (N_20488,N_19840,N_19789);
xor U20489 (N_20489,N_19986,N_19966);
nand U20490 (N_20490,N_19647,N_19978);
or U20491 (N_20491,N_19539,N_19955);
xor U20492 (N_20492,N_19728,N_19995);
nand U20493 (N_20493,N_19836,N_19725);
xnor U20494 (N_20494,N_19539,N_19741);
or U20495 (N_20495,N_19568,N_19914);
xor U20496 (N_20496,N_19589,N_19840);
nor U20497 (N_20497,N_19423,N_19849);
and U20498 (N_20498,N_19726,N_19614);
or U20499 (N_20499,N_19672,N_19732);
xnor U20500 (N_20500,N_19753,N_19878);
nor U20501 (N_20501,N_19729,N_19772);
and U20502 (N_20502,N_19938,N_19511);
nor U20503 (N_20503,N_19742,N_19884);
nor U20504 (N_20504,N_19689,N_19771);
xnor U20505 (N_20505,N_19745,N_19616);
xnor U20506 (N_20506,N_19806,N_19439);
nor U20507 (N_20507,N_19632,N_19999);
and U20508 (N_20508,N_19538,N_19656);
or U20509 (N_20509,N_19778,N_19968);
and U20510 (N_20510,N_19510,N_19804);
or U20511 (N_20511,N_19676,N_19454);
or U20512 (N_20512,N_19830,N_19836);
nand U20513 (N_20513,N_19695,N_19697);
or U20514 (N_20514,N_19659,N_19642);
and U20515 (N_20515,N_19966,N_19835);
nand U20516 (N_20516,N_19391,N_19545);
or U20517 (N_20517,N_19913,N_19579);
xor U20518 (N_20518,N_19761,N_19444);
nor U20519 (N_20519,N_19614,N_19908);
or U20520 (N_20520,N_19453,N_19765);
and U20521 (N_20521,N_19582,N_19881);
xor U20522 (N_20522,N_19947,N_19988);
or U20523 (N_20523,N_19595,N_19797);
nor U20524 (N_20524,N_19890,N_19727);
or U20525 (N_20525,N_19731,N_19821);
and U20526 (N_20526,N_19444,N_19855);
and U20527 (N_20527,N_19748,N_19977);
xor U20528 (N_20528,N_19856,N_19965);
xor U20529 (N_20529,N_19976,N_19837);
nor U20530 (N_20530,N_19461,N_19444);
or U20531 (N_20531,N_19786,N_19739);
or U20532 (N_20532,N_19830,N_19760);
and U20533 (N_20533,N_19589,N_19742);
nor U20534 (N_20534,N_19951,N_19433);
nor U20535 (N_20535,N_19382,N_19413);
or U20536 (N_20536,N_19552,N_19621);
and U20537 (N_20537,N_19921,N_19397);
or U20538 (N_20538,N_19699,N_19750);
nor U20539 (N_20539,N_19631,N_19617);
nor U20540 (N_20540,N_19716,N_19711);
and U20541 (N_20541,N_19892,N_19455);
or U20542 (N_20542,N_19816,N_19384);
or U20543 (N_20543,N_19674,N_19589);
xor U20544 (N_20544,N_19913,N_19986);
or U20545 (N_20545,N_19516,N_19393);
xor U20546 (N_20546,N_19621,N_19822);
and U20547 (N_20547,N_19516,N_19915);
or U20548 (N_20548,N_19757,N_19540);
xnor U20549 (N_20549,N_19929,N_19856);
nand U20550 (N_20550,N_19750,N_19868);
nand U20551 (N_20551,N_19907,N_19495);
or U20552 (N_20552,N_19954,N_19579);
nand U20553 (N_20553,N_19831,N_19448);
and U20554 (N_20554,N_19920,N_19540);
or U20555 (N_20555,N_19401,N_19965);
nor U20556 (N_20556,N_19554,N_19644);
or U20557 (N_20557,N_19470,N_19721);
nor U20558 (N_20558,N_19387,N_19889);
nand U20559 (N_20559,N_19497,N_19675);
xnor U20560 (N_20560,N_19616,N_19873);
or U20561 (N_20561,N_19633,N_19986);
or U20562 (N_20562,N_19988,N_19975);
nand U20563 (N_20563,N_19893,N_19981);
or U20564 (N_20564,N_19707,N_19722);
nand U20565 (N_20565,N_19846,N_19653);
nand U20566 (N_20566,N_19982,N_19931);
or U20567 (N_20567,N_19442,N_19659);
and U20568 (N_20568,N_19620,N_19879);
xor U20569 (N_20569,N_19772,N_19534);
or U20570 (N_20570,N_19470,N_19958);
nand U20571 (N_20571,N_19576,N_19727);
nand U20572 (N_20572,N_19885,N_19426);
nor U20573 (N_20573,N_19547,N_19378);
or U20574 (N_20574,N_19891,N_19382);
nand U20575 (N_20575,N_19496,N_19540);
or U20576 (N_20576,N_19543,N_19794);
xor U20577 (N_20577,N_19941,N_19552);
and U20578 (N_20578,N_19583,N_19698);
xor U20579 (N_20579,N_19771,N_19862);
and U20580 (N_20580,N_19702,N_19749);
xor U20581 (N_20581,N_19755,N_19424);
nor U20582 (N_20582,N_19680,N_19901);
nand U20583 (N_20583,N_19815,N_19669);
nand U20584 (N_20584,N_19733,N_19981);
and U20585 (N_20585,N_19446,N_19915);
xnor U20586 (N_20586,N_19714,N_19831);
nand U20587 (N_20587,N_19649,N_19823);
xnor U20588 (N_20588,N_19665,N_19666);
or U20589 (N_20589,N_19917,N_19603);
and U20590 (N_20590,N_19413,N_19550);
and U20591 (N_20591,N_19572,N_19754);
nor U20592 (N_20592,N_19872,N_19733);
or U20593 (N_20593,N_19969,N_19978);
or U20594 (N_20594,N_19860,N_19813);
xnor U20595 (N_20595,N_19810,N_19992);
and U20596 (N_20596,N_19577,N_19565);
xnor U20597 (N_20597,N_19982,N_19945);
xnor U20598 (N_20598,N_19552,N_19993);
or U20599 (N_20599,N_19715,N_19396);
nand U20600 (N_20600,N_19613,N_19677);
xor U20601 (N_20601,N_19610,N_19511);
nor U20602 (N_20602,N_19381,N_19573);
xnor U20603 (N_20603,N_19718,N_19535);
nor U20604 (N_20604,N_19733,N_19711);
and U20605 (N_20605,N_19710,N_19606);
xnor U20606 (N_20606,N_19956,N_19650);
nor U20607 (N_20607,N_19842,N_19684);
and U20608 (N_20608,N_19739,N_19812);
or U20609 (N_20609,N_19519,N_19486);
nand U20610 (N_20610,N_19405,N_19789);
or U20611 (N_20611,N_19785,N_19906);
and U20612 (N_20612,N_19936,N_19857);
or U20613 (N_20613,N_19534,N_19421);
nor U20614 (N_20614,N_19384,N_19965);
or U20615 (N_20615,N_19517,N_19848);
nand U20616 (N_20616,N_19652,N_19610);
nand U20617 (N_20617,N_19763,N_19719);
or U20618 (N_20618,N_19414,N_19640);
nand U20619 (N_20619,N_19852,N_19690);
or U20620 (N_20620,N_19635,N_19610);
xor U20621 (N_20621,N_19514,N_19436);
xor U20622 (N_20622,N_19775,N_19818);
nand U20623 (N_20623,N_19762,N_19916);
nand U20624 (N_20624,N_19666,N_19380);
xor U20625 (N_20625,N_20057,N_20392);
nand U20626 (N_20626,N_20036,N_20336);
and U20627 (N_20627,N_20220,N_20483);
nor U20628 (N_20628,N_20241,N_20591);
xor U20629 (N_20629,N_20531,N_20138);
xor U20630 (N_20630,N_20107,N_20040);
xor U20631 (N_20631,N_20553,N_20323);
nor U20632 (N_20632,N_20484,N_20304);
nor U20633 (N_20633,N_20270,N_20221);
nand U20634 (N_20634,N_20294,N_20544);
nand U20635 (N_20635,N_20124,N_20134);
or U20636 (N_20636,N_20455,N_20361);
nand U20637 (N_20637,N_20616,N_20197);
nor U20638 (N_20638,N_20318,N_20487);
nand U20639 (N_20639,N_20267,N_20133);
nand U20640 (N_20640,N_20449,N_20486);
and U20641 (N_20641,N_20493,N_20492);
xnor U20642 (N_20642,N_20309,N_20230);
and U20643 (N_20643,N_20590,N_20005);
or U20644 (N_20644,N_20268,N_20025);
nand U20645 (N_20645,N_20118,N_20100);
and U20646 (N_20646,N_20279,N_20578);
or U20647 (N_20647,N_20212,N_20381);
nand U20648 (N_20648,N_20296,N_20184);
nand U20649 (N_20649,N_20021,N_20605);
nand U20650 (N_20650,N_20060,N_20186);
or U20651 (N_20651,N_20265,N_20130);
or U20652 (N_20652,N_20528,N_20460);
nor U20653 (N_20653,N_20365,N_20041);
and U20654 (N_20654,N_20191,N_20613);
or U20655 (N_20655,N_20252,N_20462);
or U20656 (N_20656,N_20007,N_20328);
xnor U20657 (N_20657,N_20196,N_20214);
or U20658 (N_20658,N_20141,N_20083);
nor U20659 (N_20659,N_20213,N_20282);
and U20660 (N_20660,N_20384,N_20136);
xnor U20661 (N_20661,N_20335,N_20488);
nand U20662 (N_20662,N_20371,N_20307);
xor U20663 (N_20663,N_20038,N_20208);
or U20664 (N_20664,N_20034,N_20610);
nor U20665 (N_20665,N_20079,N_20413);
or U20666 (N_20666,N_20390,N_20437);
or U20667 (N_20667,N_20147,N_20288);
and U20668 (N_20668,N_20148,N_20073);
and U20669 (N_20669,N_20565,N_20573);
and U20670 (N_20670,N_20574,N_20317);
nand U20671 (N_20671,N_20319,N_20217);
nand U20672 (N_20672,N_20406,N_20026);
or U20673 (N_20673,N_20002,N_20400);
nor U20674 (N_20674,N_20132,N_20620);
nand U20675 (N_20675,N_20447,N_20539);
and U20676 (N_20676,N_20510,N_20280);
nor U20677 (N_20677,N_20234,N_20346);
nor U20678 (N_20678,N_20172,N_20181);
nand U20679 (N_20679,N_20205,N_20609);
nand U20680 (N_20680,N_20473,N_20287);
nand U20681 (N_20681,N_20071,N_20242);
or U20682 (N_20682,N_20325,N_20209);
xor U20683 (N_20683,N_20190,N_20433);
nor U20684 (N_20684,N_20491,N_20135);
and U20685 (N_20685,N_20017,N_20056);
nand U20686 (N_20686,N_20117,N_20291);
xor U20687 (N_20687,N_20074,N_20314);
xor U20688 (N_20688,N_20321,N_20383);
nand U20689 (N_20689,N_20183,N_20103);
or U20690 (N_20690,N_20373,N_20570);
nand U20691 (N_20691,N_20224,N_20254);
and U20692 (N_20692,N_20431,N_20192);
xnor U20693 (N_20693,N_20305,N_20085);
xor U20694 (N_20694,N_20350,N_20116);
or U20695 (N_20695,N_20066,N_20398);
and U20696 (N_20696,N_20558,N_20016);
or U20697 (N_20697,N_20408,N_20320);
or U20698 (N_20698,N_20370,N_20253);
or U20699 (N_20699,N_20272,N_20396);
or U20700 (N_20700,N_20436,N_20012);
nor U20701 (N_20701,N_20478,N_20228);
nor U20702 (N_20702,N_20087,N_20417);
or U20703 (N_20703,N_20474,N_20584);
and U20704 (N_20704,N_20356,N_20549);
nand U20705 (N_20705,N_20432,N_20334);
nor U20706 (N_20706,N_20247,N_20472);
nand U20707 (N_20707,N_20042,N_20621);
nand U20708 (N_20708,N_20589,N_20115);
and U20709 (N_20709,N_20511,N_20581);
nand U20710 (N_20710,N_20399,N_20457);
xor U20711 (N_20711,N_20586,N_20162);
nor U20712 (N_20712,N_20033,N_20157);
or U20713 (N_20713,N_20201,N_20615);
nand U20714 (N_20714,N_20092,N_20149);
xnor U20715 (N_20715,N_20563,N_20226);
xor U20716 (N_20716,N_20559,N_20515);
nand U20717 (N_20717,N_20232,N_20137);
nand U20718 (N_20718,N_20127,N_20182);
or U20719 (N_20719,N_20407,N_20010);
nand U20720 (N_20720,N_20504,N_20552);
and U20721 (N_20721,N_20331,N_20046);
nand U20722 (N_20722,N_20543,N_20029);
and U20723 (N_20723,N_20490,N_20379);
and U20724 (N_20724,N_20262,N_20532);
xor U20725 (N_20725,N_20179,N_20499);
and U20726 (N_20726,N_20146,N_20524);
nand U20727 (N_20727,N_20275,N_20047);
and U20728 (N_20728,N_20322,N_20290);
nor U20729 (N_20729,N_20372,N_20126);
nand U20730 (N_20730,N_20061,N_20311);
or U20731 (N_20731,N_20299,N_20077);
or U20732 (N_20732,N_20378,N_20516);
nand U20733 (N_20733,N_20055,N_20110);
or U20734 (N_20734,N_20095,N_20065);
nand U20735 (N_20735,N_20258,N_20386);
nor U20736 (N_20736,N_20301,N_20240);
or U20737 (N_20737,N_20113,N_20150);
nand U20738 (N_20738,N_20557,N_20194);
nor U20739 (N_20739,N_20517,N_20572);
nor U20740 (N_20740,N_20211,N_20271);
nand U20741 (N_20741,N_20170,N_20145);
or U20742 (N_20742,N_20054,N_20366);
nand U20743 (N_20743,N_20342,N_20536);
xnor U20744 (N_20744,N_20550,N_20588);
nand U20745 (N_20745,N_20530,N_20180);
nand U20746 (N_20746,N_20344,N_20359);
nor U20747 (N_20747,N_20104,N_20480);
nand U20748 (N_20748,N_20561,N_20345);
xnor U20749 (N_20749,N_20114,N_20210);
or U20750 (N_20750,N_20128,N_20445);
and U20751 (N_20751,N_20506,N_20514);
xor U20752 (N_20752,N_20256,N_20028);
nor U20753 (N_20753,N_20303,N_20161);
nor U20754 (N_20754,N_20585,N_20418);
and U20755 (N_20755,N_20278,N_20402);
xnor U20756 (N_20756,N_20596,N_20566);
nor U20757 (N_20757,N_20101,N_20423);
or U20758 (N_20758,N_20369,N_20091);
nand U20759 (N_20759,N_20102,N_20422);
xnor U20760 (N_20760,N_20249,N_20125);
nand U20761 (N_20761,N_20140,N_20097);
nor U20762 (N_20762,N_20058,N_20355);
or U20763 (N_20763,N_20261,N_20526);
nor U20764 (N_20764,N_20229,N_20072);
and U20765 (N_20765,N_20439,N_20389);
or U20766 (N_20766,N_20090,N_20599);
nand U20767 (N_20767,N_20219,N_20037);
nand U20768 (N_20768,N_20604,N_20341);
nand U20769 (N_20769,N_20380,N_20298);
and U20770 (N_20770,N_20603,N_20419);
or U20771 (N_20771,N_20218,N_20403);
or U20772 (N_20772,N_20571,N_20274);
or U20773 (N_20773,N_20030,N_20156);
nor U20774 (N_20774,N_20583,N_20143);
and U20775 (N_20775,N_20231,N_20368);
xor U20776 (N_20776,N_20502,N_20059);
nor U20777 (N_20777,N_20458,N_20353);
nand U20778 (N_20778,N_20592,N_20397);
or U20779 (N_20779,N_20442,N_20312);
nand U20780 (N_20780,N_20204,N_20300);
nor U20781 (N_20781,N_20052,N_20428);
or U20782 (N_20782,N_20098,N_20468);
or U20783 (N_20783,N_20154,N_20175);
and U20784 (N_20784,N_20080,N_20215);
nor U20785 (N_20785,N_20580,N_20306);
and U20786 (N_20786,N_20310,N_20501);
nor U20787 (N_20787,N_20505,N_20440);
nand U20788 (N_20788,N_20485,N_20546);
nand U20789 (N_20789,N_20248,N_20465);
or U20790 (N_20790,N_20452,N_20374);
nand U20791 (N_20791,N_20203,N_20131);
or U20792 (N_20792,N_20283,N_20551);
nor U20793 (N_20793,N_20111,N_20263);
xnor U20794 (N_20794,N_20367,N_20329);
xor U20795 (N_20795,N_20009,N_20001);
nand U20796 (N_20796,N_20520,N_20388);
nand U20797 (N_20797,N_20424,N_20416);
xnor U20798 (N_20798,N_20405,N_20284);
nand U20799 (N_20799,N_20463,N_20286);
xor U20800 (N_20800,N_20601,N_20023);
or U20801 (N_20801,N_20509,N_20622);
nand U20802 (N_20802,N_20562,N_20438);
and U20803 (N_20803,N_20160,N_20412);
nand U20804 (N_20804,N_20343,N_20174);
and U20805 (N_20805,N_20257,N_20554);
nand U20806 (N_20806,N_20534,N_20339);
nand U20807 (N_20807,N_20595,N_20008);
xor U20808 (N_20808,N_20618,N_20227);
nor U20809 (N_20809,N_20123,N_20541);
or U20810 (N_20810,N_20357,N_20450);
nand U20811 (N_20811,N_20513,N_20049);
xnor U20812 (N_20812,N_20223,N_20597);
nand U20813 (N_20813,N_20582,N_20302);
nand U20814 (N_20814,N_20611,N_20414);
nand U20815 (N_20815,N_20142,N_20082);
nand U20816 (N_20816,N_20426,N_20015);
nor U20817 (N_20817,N_20099,N_20375);
xnor U20818 (N_20818,N_20276,N_20164);
or U20819 (N_20819,N_20429,N_20189);
nand U20820 (N_20820,N_20144,N_20503);
xnor U20821 (N_20821,N_20260,N_20069);
nor U20822 (N_20822,N_20293,N_20421);
or U20823 (N_20823,N_20420,N_20266);
nand U20824 (N_20824,N_20614,N_20555);
xnor U20825 (N_20825,N_20239,N_20243);
nor U20826 (N_20826,N_20285,N_20612);
or U20827 (N_20827,N_20560,N_20094);
or U20828 (N_20828,N_20489,N_20165);
and U20829 (N_20829,N_20199,N_20163);
and U20830 (N_20830,N_20019,N_20188);
or U20831 (N_20831,N_20151,N_20236);
nor U20832 (N_20832,N_20575,N_20018);
xnor U20833 (N_20833,N_20545,N_20434);
or U20834 (N_20834,N_20394,N_20479);
and U20835 (N_20835,N_20577,N_20579);
and U20836 (N_20836,N_20569,N_20385);
nand U20837 (N_20837,N_20568,N_20525);
and U20838 (N_20838,N_20173,N_20382);
or U20839 (N_20839,N_20624,N_20477);
xnor U20840 (N_20840,N_20540,N_20443);
xor U20841 (N_20841,N_20354,N_20178);
xnor U20842 (N_20842,N_20251,N_20200);
xor U20843 (N_20843,N_20522,N_20177);
nand U20844 (N_20844,N_20348,N_20576);
or U20845 (N_20845,N_20376,N_20292);
nand U20846 (N_20846,N_20084,N_20004);
and U20847 (N_20847,N_20139,N_20297);
xnor U20848 (N_20848,N_20587,N_20410);
nand U20849 (N_20849,N_20623,N_20467);
nand U20850 (N_20850,N_20527,N_20441);
nand U20851 (N_20851,N_20507,N_20498);
and U20852 (N_20852,N_20351,N_20519);
xnor U20853 (N_20853,N_20593,N_20481);
nor U20854 (N_20854,N_20387,N_20259);
xor U20855 (N_20855,N_20043,N_20062);
nand U20856 (N_20856,N_20496,N_20129);
xor U20857 (N_20857,N_20393,N_20606);
and U20858 (N_20858,N_20245,N_20482);
nor U20859 (N_20859,N_20521,N_20153);
nor U20860 (N_20860,N_20237,N_20088);
nor U20861 (N_20861,N_20076,N_20330);
and U20862 (N_20862,N_20168,N_20542);
or U20863 (N_20863,N_20273,N_20535);
or U20864 (N_20864,N_20362,N_20289);
nor U20865 (N_20865,N_20363,N_20564);
nand U20866 (N_20866,N_20024,N_20411);
nor U20867 (N_20867,N_20364,N_20324);
xor U20868 (N_20868,N_20451,N_20547);
nor U20869 (N_20869,N_20401,N_20078);
xor U20870 (N_20870,N_20152,N_20207);
nor U20871 (N_20871,N_20316,N_20166);
xnor U20872 (N_20872,N_20171,N_20000);
nor U20873 (N_20873,N_20454,N_20315);
or U20874 (N_20874,N_20063,N_20337);
or U20875 (N_20875,N_20255,N_20050);
and U20876 (N_20876,N_20169,N_20529);
and U20877 (N_20877,N_20053,N_20158);
nor U20878 (N_20878,N_20459,N_20430);
xor U20879 (N_20879,N_20120,N_20122);
xnor U20880 (N_20880,N_20086,N_20011);
nor U20881 (N_20881,N_20202,N_20548);
xnor U20882 (N_20882,N_20108,N_20600);
nand U20883 (N_20883,N_20333,N_20193);
xnor U20884 (N_20884,N_20444,N_20067);
or U20885 (N_20885,N_20075,N_20475);
or U20886 (N_20886,N_20537,N_20045);
or U20887 (N_20887,N_20081,N_20377);
nor U20888 (N_20888,N_20195,N_20360);
nand U20889 (N_20889,N_20497,N_20556);
nor U20890 (N_20890,N_20466,N_20014);
or U20891 (N_20891,N_20464,N_20006);
nand U20892 (N_20892,N_20494,N_20617);
nand U20893 (N_20893,N_20340,N_20044);
nand U20894 (N_20894,N_20495,N_20216);
xnor U20895 (N_20895,N_20027,N_20250);
or U20896 (N_20896,N_20469,N_20313);
nor U20897 (N_20897,N_20446,N_20471);
or U20898 (N_20898,N_20238,N_20500);
or U20899 (N_20899,N_20089,N_20176);
or U20900 (N_20900,N_20352,N_20105);
xnor U20901 (N_20901,N_20244,N_20523);
nand U20902 (N_20902,N_20031,N_20198);
nor U20903 (N_20903,N_20096,N_20427);
nand U20904 (N_20904,N_20020,N_20159);
and U20905 (N_20905,N_20235,N_20119);
nand U20906 (N_20906,N_20222,N_20518);
nor U20907 (N_20907,N_20035,N_20264);
nor U20908 (N_20908,N_20308,N_20508);
or U20909 (N_20909,N_20358,N_20327);
xor U20910 (N_20910,N_20187,N_20453);
nand U20911 (N_20911,N_20048,N_20093);
and U20912 (N_20912,N_20233,N_20013);
and U20913 (N_20913,N_20456,N_20404);
xnor U20914 (N_20914,N_20448,N_20476);
nor U20915 (N_20915,N_20594,N_20022);
nor U20916 (N_20916,N_20281,N_20051);
or U20917 (N_20917,N_20349,N_20391);
nor U20918 (N_20918,N_20003,N_20409);
nand U20919 (N_20919,N_20338,N_20512);
and U20920 (N_20920,N_20246,N_20435);
nor U20921 (N_20921,N_20064,N_20070);
and U20922 (N_20922,N_20121,N_20567);
nor U20923 (N_20923,N_20347,N_20608);
or U20924 (N_20924,N_20461,N_20602);
xor U20925 (N_20925,N_20533,N_20425);
nor U20926 (N_20926,N_20068,N_20225);
nand U20927 (N_20927,N_20155,N_20470);
nor U20928 (N_20928,N_20185,N_20538);
nor U20929 (N_20929,N_20326,N_20607);
or U20930 (N_20930,N_20112,N_20032);
xnor U20931 (N_20931,N_20109,N_20619);
or U20932 (N_20932,N_20395,N_20039);
nor U20933 (N_20933,N_20167,N_20295);
or U20934 (N_20934,N_20106,N_20277);
nand U20935 (N_20935,N_20332,N_20206);
and U20936 (N_20936,N_20269,N_20598);
nor U20937 (N_20937,N_20415,N_20106);
and U20938 (N_20938,N_20419,N_20365);
xnor U20939 (N_20939,N_20289,N_20318);
xor U20940 (N_20940,N_20045,N_20250);
or U20941 (N_20941,N_20188,N_20390);
and U20942 (N_20942,N_20007,N_20623);
or U20943 (N_20943,N_20001,N_20467);
xor U20944 (N_20944,N_20223,N_20377);
xor U20945 (N_20945,N_20037,N_20221);
nor U20946 (N_20946,N_20106,N_20352);
nand U20947 (N_20947,N_20219,N_20384);
or U20948 (N_20948,N_20468,N_20162);
nor U20949 (N_20949,N_20554,N_20506);
and U20950 (N_20950,N_20272,N_20110);
nor U20951 (N_20951,N_20118,N_20164);
nor U20952 (N_20952,N_20094,N_20428);
xor U20953 (N_20953,N_20506,N_20126);
and U20954 (N_20954,N_20509,N_20258);
nand U20955 (N_20955,N_20473,N_20349);
and U20956 (N_20956,N_20309,N_20255);
nor U20957 (N_20957,N_20147,N_20071);
nand U20958 (N_20958,N_20281,N_20078);
and U20959 (N_20959,N_20223,N_20076);
or U20960 (N_20960,N_20309,N_20155);
nand U20961 (N_20961,N_20163,N_20051);
xor U20962 (N_20962,N_20397,N_20278);
nor U20963 (N_20963,N_20148,N_20397);
nand U20964 (N_20964,N_20039,N_20299);
xor U20965 (N_20965,N_20602,N_20134);
nand U20966 (N_20966,N_20120,N_20082);
nor U20967 (N_20967,N_20451,N_20602);
and U20968 (N_20968,N_20525,N_20104);
nor U20969 (N_20969,N_20515,N_20344);
or U20970 (N_20970,N_20349,N_20604);
nor U20971 (N_20971,N_20574,N_20123);
nor U20972 (N_20972,N_20191,N_20253);
or U20973 (N_20973,N_20363,N_20245);
or U20974 (N_20974,N_20516,N_20471);
xor U20975 (N_20975,N_20317,N_20266);
nand U20976 (N_20976,N_20121,N_20393);
nand U20977 (N_20977,N_20526,N_20573);
or U20978 (N_20978,N_20430,N_20241);
nand U20979 (N_20979,N_20411,N_20447);
or U20980 (N_20980,N_20568,N_20565);
and U20981 (N_20981,N_20456,N_20043);
and U20982 (N_20982,N_20202,N_20613);
or U20983 (N_20983,N_20468,N_20197);
or U20984 (N_20984,N_20175,N_20282);
nand U20985 (N_20985,N_20520,N_20531);
xor U20986 (N_20986,N_20401,N_20571);
or U20987 (N_20987,N_20304,N_20422);
and U20988 (N_20988,N_20035,N_20299);
nor U20989 (N_20989,N_20224,N_20319);
nand U20990 (N_20990,N_20086,N_20264);
and U20991 (N_20991,N_20369,N_20016);
xor U20992 (N_20992,N_20043,N_20470);
and U20993 (N_20993,N_20134,N_20570);
nand U20994 (N_20994,N_20514,N_20168);
nand U20995 (N_20995,N_20619,N_20516);
xnor U20996 (N_20996,N_20156,N_20247);
and U20997 (N_20997,N_20222,N_20115);
nor U20998 (N_20998,N_20601,N_20468);
or U20999 (N_20999,N_20068,N_20369);
nand U21000 (N_21000,N_20597,N_20132);
or U21001 (N_21001,N_20143,N_20255);
and U21002 (N_21002,N_20434,N_20496);
nand U21003 (N_21003,N_20523,N_20193);
nor U21004 (N_21004,N_20130,N_20520);
nor U21005 (N_21005,N_20242,N_20004);
and U21006 (N_21006,N_20368,N_20251);
and U21007 (N_21007,N_20307,N_20359);
and U21008 (N_21008,N_20060,N_20300);
and U21009 (N_21009,N_20461,N_20126);
and U21010 (N_21010,N_20489,N_20073);
xnor U21011 (N_21011,N_20193,N_20376);
or U21012 (N_21012,N_20404,N_20447);
xnor U21013 (N_21013,N_20244,N_20563);
and U21014 (N_21014,N_20521,N_20090);
xor U21015 (N_21015,N_20621,N_20454);
xnor U21016 (N_21016,N_20572,N_20372);
or U21017 (N_21017,N_20275,N_20165);
nand U21018 (N_21018,N_20064,N_20518);
nand U21019 (N_21019,N_20358,N_20088);
xor U21020 (N_21020,N_20076,N_20288);
or U21021 (N_21021,N_20195,N_20594);
or U21022 (N_21022,N_20119,N_20477);
xnor U21023 (N_21023,N_20358,N_20377);
xor U21024 (N_21024,N_20329,N_20332);
nand U21025 (N_21025,N_20022,N_20086);
or U21026 (N_21026,N_20291,N_20504);
or U21027 (N_21027,N_20450,N_20373);
nand U21028 (N_21028,N_20558,N_20051);
or U21029 (N_21029,N_20372,N_20490);
and U21030 (N_21030,N_20255,N_20603);
xor U21031 (N_21031,N_20137,N_20114);
and U21032 (N_21032,N_20082,N_20519);
and U21033 (N_21033,N_20373,N_20202);
nor U21034 (N_21034,N_20223,N_20292);
xnor U21035 (N_21035,N_20013,N_20242);
nor U21036 (N_21036,N_20432,N_20236);
nand U21037 (N_21037,N_20036,N_20401);
xnor U21038 (N_21038,N_20470,N_20473);
nand U21039 (N_21039,N_20342,N_20271);
xor U21040 (N_21040,N_20217,N_20358);
nand U21041 (N_21041,N_20399,N_20225);
nor U21042 (N_21042,N_20249,N_20431);
xor U21043 (N_21043,N_20598,N_20621);
xor U21044 (N_21044,N_20003,N_20196);
or U21045 (N_21045,N_20450,N_20094);
xnor U21046 (N_21046,N_20320,N_20139);
nor U21047 (N_21047,N_20412,N_20325);
nor U21048 (N_21048,N_20465,N_20356);
xor U21049 (N_21049,N_20432,N_20124);
or U21050 (N_21050,N_20358,N_20479);
nand U21051 (N_21051,N_20575,N_20398);
xor U21052 (N_21052,N_20335,N_20013);
nand U21053 (N_21053,N_20010,N_20001);
nand U21054 (N_21054,N_20567,N_20331);
and U21055 (N_21055,N_20495,N_20488);
or U21056 (N_21056,N_20200,N_20050);
xor U21057 (N_21057,N_20489,N_20386);
or U21058 (N_21058,N_20542,N_20373);
nand U21059 (N_21059,N_20536,N_20546);
nand U21060 (N_21060,N_20405,N_20496);
nand U21061 (N_21061,N_20168,N_20509);
and U21062 (N_21062,N_20443,N_20341);
nand U21063 (N_21063,N_20296,N_20260);
nor U21064 (N_21064,N_20592,N_20055);
nand U21065 (N_21065,N_20457,N_20016);
xor U21066 (N_21066,N_20552,N_20079);
and U21067 (N_21067,N_20027,N_20113);
nand U21068 (N_21068,N_20537,N_20604);
or U21069 (N_21069,N_20503,N_20265);
xor U21070 (N_21070,N_20305,N_20032);
nand U21071 (N_21071,N_20547,N_20070);
or U21072 (N_21072,N_20131,N_20175);
xor U21073 (N_21073,N_20249,N_20591);
and U21074 (N_21074,N_20504,N_20151);
or U21075 (N_21075,N_20186,N_20462);
xor U21076 (N_21076,N_20300,N_20348);
nand U21077 (N_21077,N_20203,N_20001);
nor U21078 (N_21078,N_20440,N_20360);
or U21079 (N_21079,N_20356,N_20380);
nand U21080 (N_21080,N_20565,N_20213);
nor U21081 (N_21081,N_20172,N_20059);
and U21082 (N_21082,N_20389,N_20146);
and U21083 (N_21083,N_20435,N_20464);
or U21084 (N_21084,N_20381,N_20452);
or U21085 (N_21085,N_20165,N_20128);
xnor U21086 (N_21086,N_20466,N_20599);
xnor U21087 (N_21087,N_20069,N_20154);
xor U21088 (N_21088,N_20479,N_20272);
nand U21089 (N_21089,N_20060,N_20410);
xor U21090 (N_21090,N_20276,N_20404);
xor U21091 (N_21091,N_20257,N_20499);
nand U21092 (N_21092,N_20110,N_20094);
nand U21093 (N_21093,N_20401,N_20370);
nor U21094 (N_21094,N_20128,N_20612);
and U21095 (N_21095,N_20486,N_20586);
or U21096 (N_21096,N_20160,N_20175);
or U21097 (N_21097,N_20001,N_20428);
and U21098 (N_21098,N_20255,N_20078);
xor U21099 (N_21099,N_20036,N_20209);
or U21100 (N_21100,N_20418,N_20480);
xor U21101 (N_21101,N_20048,N_20470);
and U21102 (N_21102,N_20236,N_20210);
xnor U21103 (N_21103,N_20014,N_20510);
xor U21104 (N_21104,N_20193,N_20114);
and U21105 (N_21105,N_20043,N_20182);
or U21106 (N_21106,N_20256,N_20288);
nor U21107 (N_21107,N_20228,N_20090);
nand U21108 (N_21108,N_20412,N_20321);
nand U21109 (N_21109,N_20450,N_20383);
and U21110 (N_21110,N_20443,N_20112);
xnor U21111 (N_21111,N_20370,N_20080);
and U21112 (N_21112,N_20287,N_20057);
xnor U21113 (N_21113,N_20104,N_20195);
or U21114 (N_21114,N_20189,N_20573);
or U21115 (N_21115,N_20379,N_20401);
nor U21116 (N_21116,N_20206,N_20344);
xor U21117 (N_21117,N_20145,N_20099);
nand U21118 (N_21118,N_20398,N_20012);
and U21119 (N_21119,N_20187,N_20224);
and U21120 (N_21120,N_20288,N_20297);
and U21121 (N_21121,N_20346,N_20306);
nor U21122 (N_21122,N_20201,N_20340);
and U21123 (N_21123,N_20605,N_20548);
or U21124 (N_21124,N_20362,N_20326);
nor U21125 (N_21125,N_20032,N_20321);
nand U21126 (N_21126,N_20195,N_20401);
nor U21127 (N_21127,N_20093,N_20332);
and U21128 (N_21128,N_20331,N_20299);
or U21129 (N_21129,N_20393,N_20283);
nand U21130 (N_21130,N_20589,N_20131);
xor U21131 (N_21131,N_20179,N_20044);
or U21132 (N_21132,N_20119,N_20250);
and U21133 (N_21133,N_20461,N_20113);
or U21134 (N_21134,N_20115,N_20462);
nand U21135 (N_21135,N_20515,N_20267);
nor U21136 (N_21136,N_20333,N_20234);
nor U21137 (N_21137,N_20147,N_20558);
or U21138 (N_21138,N_20238,N_20119);
xor U21139 (N_21139,N_20310,N_20213);
or U21140 (N_21140,N_20293,N_20509);
xnor U21141 (N_21141,N_20549,N_20061);
xor U21142 (N_21142,N_20327,N_20620);
xnor U21143 (N_21143,N_20281,N_20431);
and U21144 (N_21144,N_20047,N_20111);
xnor U21145 (N_21145,N_20479,N_20008);
nor U21146 (N_21146,N_20136,N_20069);
xor U21147 (N_21147,N_20559,N_20429);
xor U21148 (N_21148,N_20314,N_20450);
nand U21149 (N_21149,N_20419,N_20109);
and U21150 (N_21150,N_20534,N_20470);
xnor U21151 (N_21151,N_20399,N_20471);
nand U21152 (N_21152,N_20578,N_20209);
nand U21153 (N_21153,N_20335,N_20097);
nor U21154 (N_21154,N_20128,N_20337);
xor U21155 (N_21155,N_20087,N_20032);
nor U21156 (N_21156,N_20553,N_20616);
nor U21157 (N_21157,N_20227,N_20268);
and U21158 (N_21158,N_20187,N_20234);
nor U21159 (N_21159,N_20121,N_20227);
nor U21160 (N_21160,N_20114,N_20397);
nor U21161 (N_21161,N_20420,N_20366);
nand U21162 (N_21162,N_20031,N_20096);
xor U21163 (N_21163,N_20243,N_20529);
xnor U21164 (N_21164,N_20287,N_20470);
nand U21165 (N_21165,N_20279,N_20110);
or U21166 (N_21166,N_20391,N_20359);
xor U21167 (N_21167,N_20177,N_20110);
and U21168 (N_21168,N_20316,N_20483);
or U21169 (N_21169,N_20329,N_20176);
nor U21170 (N_21170,N_20197,N_20196);
nand U21171 (N_21171,N_20290,N_20127);
nor U21172 (N_21172,N_20172,N_20067);
and U21173 (N_21173,N_20116,N_20100);
and U21174 (N_21174,N_20579,N_20197);
nor U21175 (N_21175,N_20173,N_20186);
nor U21176 (N_21176,N_20065,N_20450);
xnor U21177 (N_21177,N_20183,N_20298);
nor U21178 (N_21178,N_20128,N_20415);
xor U21179 (N_21179,N_20296,N_20324);
nor U21180 (N_21180,N_20522,N_20238);
xor U21181 (N_21181,N_20323,N_20502);
nand U21182 (N_21182,N_20321,N_20391);
nand U21183 (N_21183,N_20362,N_20623);
nor U21184 (N_21184,N_20456,N_20020);
nand U21185 (N_21185,N_20265,N_20544);
or U21186 (N_21186,N_20131,N_20427);
and U21187 (N_21187,N_20578,N_20101);
or U21188 (N_21188,N_20229,N_20622);
nand U21189 (N_21189,N_20117,N_20356);
xnor U21190 (N_21190,N_20095,N_20459);
or U21191 (N_21191,N_20346,N_20035);
or U21192 (N_21192,N_20397,N_20543);
or U21193 (N_21193,N_20511,N_20031);
nor U21194 (N_21194,N_20363,N_20171);
or U21195 (N_21195,N_20387,N_20105);
and U21196 (N_21196,N_20469,N_20585);
and U21197 (N_21197,N_20181,N_20493);
and U21198 (N_21198,N_20313,N_20054);
or U21199 (N_21199,N_20597,N_20116);
and U21200 (N_21200,N_20028,N_20218);
and U21201 (N_21201,N_20077,N_20503);
or U21202 (N_21202,N_20341,N_20334);
or U21203 (N_21203,N_20172,N_20193);
and U21204 (N_21204,N_20041,N_20079);
xor U21205 (N_21205,N_20310,N_20273);
nand U21206 (N_21206,N_20023,N_20101);
xor U21207 (N_21207,N_20056,N_20042);
and U21208 (N_21208,N_20101,N_20264);
or U21209 (N_21209,N_20478,N_20492);
xnor U21210 (N_21210,N_20361,N_20181);
nand U21211 (N_21211,N_20279,N_20328);
xnor U21212 (N_21212,N_20265,N_20245);
xor U21213 (N_21213,N_20548,N_20573);
nand U21214 (N_21214,N_20471,N_20036);
nand U21215 (N_21215,N_20416,N_20348);
xor U21216 (N_21216,N_20508,N_20516);
or U21217 (N_21217,N_20430,N_20126);
and U21218 (N_21218,N_20073,N_20170);
xor U21219 (N_21219,N_20219,N_20549);
xnor U21220 (N_21220,N_20037,N_20043);
or U21221 (N_21221,N_20267,N_20574);
xor U21222 (N_21222,N_20240,N_20616);
nor U21223 (N_21223,N_20553,N_20125);
xnor U21224 (N_21224,N_20206,N_20618);
or U21225 (N_21225,N_20067,N_20552);
or U21226 (N_21226,N_20595,N_20579);
nor U21227 (N_21227,N_20623,N_20032);
and U21228 (N_21228,N_20482,N_20180);
or U21229 (N_21229,N_20139,N_20287);
nor U21230 (N_21230,N_20453,N_20463);
nor U21231 (N_21231,N_20060,N_20483);
xor U21232 (N_21232,N_20105,N_20527);
xnor U21233 (N_21233,N_20385,N_20595);
or U21234 (N_21234,N_20103,N_20122);
nor U21235 (N_21235,N_20219,N_20061);
and U21236 (N_21236,N_20048,N_20135);
nor U21237 (N_21237,N_20236,N_20003);
nand U21238 (N_21238,N_20143,N_20386);
and U21239 (N_21239,N_20076,N_20601);
nand U21240 (N_21240,N_20594,N_20348);
and U21241 (N_21241,N_20026,N_20223);
or U21242 (N_21242,N_20348,N_20212);
or U21243 (N_21243,N_20257,N_20172);
nand U21244 (N_21244,N_20313,N_20253);
nand U21245 (N_21245,N_20285,N_20222);
nand U21246 (N_21246,N_20576,N_20328);
nor U21247 (N_21247,N_20255,N_20358);
or U21248 (N_21248,N_20385,N_20432);
nand U21249 (N_21249,N_20317,N_20536);
xor U21250 (N_21250,N_20694,N_20698);
or U21251 (N_21251,N_21164,N_21019);
and U21252 (N_21252,N_20932,N_21025);
xor U21253 (N_21253,N_21087,N_20776);
or U21254 (N_21254,N_20761,N_20803);
xor U21255 (N_21255,N_21005,N_20830);
xor U21256 (N_21256,N_21221,N_21136);
or U21257 (N_21257,N_20762,N_21162);
nand U21258 (N_21258,N_21062,N_21125);
nor U21259 (N_21259,N_20753,N_20840);
xor U21260 (N_21260,N_21220,N_20855);
nand U21261 (N_21261,N_21031,N_20969);
or U21262 (N_21262,N_20664,N_20641);
nor U21263 (N_21263,N_21000,N_20673);
or U21264 (N_21264,N_21114,N_20936);
nand U21265 (N_21265,N_20997,N_20631);
nand U21266 (N_21266,N_20654,N_21168);
nand U21267 (N_21267,N_20721,N_20890);
xor U21268 (N_21268,N_21068,N_20957);
nand U21269 (N_21269,N_21243,N_21034);
nor U21270 (N_21270,N_21110,N_21093);
xor U21271 (N_21271,N_20649,N_21094);
and U21272 (N_21272,N_20905,N_20923);
xnor U21273 (N_21273,N_20914,N_20975);
xor U21274 (N_21274,N_20951,N_20976);
or U21275 (N_21275,N_20960,N_20966);
nor U21276 (N_21276,N_20736,N_21248);
and U21277 (N_21277,N_21035,N_21191);
or U21278 (N_21278,N_20972,N_20910);
nand U21279 (N_21279,N_21172,N_20748);
and U21280 (N_21280,N_20772,N_21127);
nor U21281 (N_21281,N_21170,N_20984);
nor U21282 (N_21282,N_20731,N_21232);
or U21283 (N_21283,N_20791,N_20719);
xor U21284 (N_21284,N_20864,N_20640);
or U21285 (N_21285,N_21119,N_20849);
or U21286 (N_21286,N_21237,N_20908);
nor U21287 (N_21287,N_21069,N_20800);
xor U21288 (N_21288,N_20667,N_21144);
xor U21289 (N_21289,N_21176,N_21222);
and U21290 (N_21290,N_21063,N_20869);
and U21291 (N_21291,N_20713,N_20931);
nand U21292 (N_21292,N_21196,N_20690);
or U21293 (N_21293,N_20741,N_20944);
nor U21294 (N_21294,N_21228,N_20685);
xor U21295 (N_21295,N_21043,N_21004);
nand U21296 (N_21296,N_21099,N_21174);
nand U21297 (N_21297,N_20684,N_21245);
or U21298 (N_21298,N_21122,N_21060);
and U21299 (N_21299,N_20819,N_21048);
xnor U21300 (N_21300,N_21002,N_21064);
or U21301 (N_21301,N_20987,N_21102);
nand U21302 (N_21302,N_20643,N_21215);
and U21303 (N_21303,N_21238,N_20739);
and U21304 (N_21304,N_21124,N_20766);
or U21305 (N_21305,N_20938,N_20839);
nand U21306 (N_21306,N_20977,N_20818);
nor U21307 (N_21307,N_20705,N_20981);
and U21308 (N_21308,N_21077,N_20876);
xor U21309 (N_21309,N_20747,N_20841);
nand U21310 (N_21310,N_20734,N_20982);
nor U21311 (N_21311,N_21246,N_20799);
nor U21312 (N_21312,N_20968,N_20699);
nor U21313 (N_21313,N_20750,N_20921);
and U21314 (N_21314,N_21173,N_20848);
nand U21315 (N_21315,N_20952,N_21189);
or U21316 (N_21316,N_20785,N_20733);
xor U21317 (N_21317,N_21109,N_20744);
and U21318 (N_21318,N_20823,N_21233);
nor U21319 (N_21319,N_20674,N_20689);
xor U21320 (N_21320,N_20949,N_20948);
xnor U21321 (N_21321,N_20806,N_20720);
or U21322 (N_21322,N_21079,N_21186);
nor U21323 (N_21323,N_20971,N_21080);
nand U21324 (N_21324,N_21135,N_20911);
and U21325 (N_21325,N_20870,N_20798);
or U21326 (N_21326,N_20730,N_20878);
and U21327 (N_21327,N_20912,N_20754);
and U21328 (N_21328,N_21015,N_21218);
xor U21329 (N_21329,N_21017,N_21070);
and U21330 (N_21330,N_21234,N_20947);
nor U21331 (N_21331,N_21078,N_21129);
nand U21332 (N_21332,N_20933,N_21138);
and U21333 (N_21333,N_21033,N_20757);
xnor U21334 (N_21334,N_20706,N_21244);
xnor U21335 (N_21335,N_20755,N_21029);
nor U21336 (N_21336,N_21150,N_20732);
nand U21337 (N_21337,N_20979,N_21216);
or U21338 (N_21338,N_21120,N_20666);
nand U21339 (N_21339,N_21123,N_20718);
or U21340 (N_21340,N_21104,N_21058);
nand U21341 (N_21341,N_21038,N_20659);
or U21342 (N_21342,N_20826,N_21030);
and U21343 (N_21343,N_21241,N_20710);
and U21344 (N_21344,N_20887,N_20860);
xnor U21345 (N_21345,N_21089,N_21113);
or U21346 (N_21346,N_21160,N_20662);
xnor U21347 (N_21347,N_20919,N_21032);
and U21348 (N_21348,N_21202,N_21203);
nand U21349 (N_21349,N_20817,N_21247);
nor U21350 (N_21350,N_20894,N_21197);
nor U21351 (N_21351,N_20632,N_21107);
nand U21352 (N_21352,N_20941,N_21026);
xor U21353 (N_21353,N_20751,N_21201);
or U21354 (N_21354,N_20629,N_20652);
or U21355 (N_21355,N_20668,N_21157);
or U21356 (N_21356,N_21112,N_20821);
and U21357 (N_21357,N_20637,N_20775);
nand U21358 (N_21358,N_21214,N_21236);
nor U21359 (N_21359,N_21020,N_21084);
xnor U21360 (N_21360,N_20712,N_20970);
or U21361 (N_21361,N_20625,N_20644);
nor U21362 (N_21362,N_20686,N_21106);
xnor U21363 (N_21363,N_20889,N_20871);
nand U21364 (N_21364,N_21010,N_21118);
and U21365 (N_21365,N_21249,N_20888);
nand U21366 (N_21366,N_20737,N_20852);
or U21367 (N_21367,N_21028,N_20700);
nand U21368 (N_21368,N_21178,N_20851);
and U21369 (N_21369,N_21166,N_21121);
and U21370 (N_21370,N_20950,N_20939);
or U21371 (N_21371,N_20788,N_21139);
or U21372 (N_21372,N_20935,N_20735);
xnor U21373 (N_21373,N_21155,N_20831);
nor U21374 (N_21374,N_20843,N_20880);
nand U21375 (N_21375,N_21042,N_20927);
or U21376 (N_21376,N_20943,N_20716);
nand U21377 (N_21377,N_20683,N_20863);
and U21378 (N_21378,N_21022,N_21108);
nor U21379 (N_21379,N_20787,N_20925);
and U21380 (N_21380,N_20915,N_21148);
nor U21381 (N_21381,N_20691,N_20867);
and U21382 (N_21382,N_20942,N_20985);
or U21383 (N_21383,N_20742,N_20930);
and U21384 (N_21384,N_21116,N_21046);
xor U21385 (N_21385,N_21023,N_20782);
nand U21386 (N_21386,N_20893,N_20760);
nor U21387 (N_21387,N_21053,N_20702);
nor U21388 (N_21388,N_20879,N_21047);
and U21389 (N_21389,N_21165,N_20940);
and U21390 (N_21390,N_20992,N_21184);
or U21391 (N_21391,N_20635,N_20630);
xnor U21392 (N_21392,N_20790,N_20675);
xnor U21393 (N_21393,N_20695,N_20795);
nand U21394 (N_21394,N_20913,N_20820);
xor U21395 (N_21395,N_21152,N_20655);
or U21396 (N_21396,N_20978,N_20872);
xor U21397 (N_21397,N_20900,N_21141);
xor U21398 (N_21398,N_20844,N_20907);
or U21399 (N_21399,N_20647,N_20687);
and U21400 (N_21400,N_20810,N_20801);
and U21401 (N_21401,N_21149,N_20922);
nor U21402 (N_21402,N_21146,N_20645);
xnor U21403 (N_21403,N_20858,N_21151);
and U21404 (N_21404,N_21006,N_20868);
nand U21405 (N_21405,N_21057,N_21003);
nor U21406 (N_21406,N_20846,N_20758);
nand U21407 (N_21407,N_21194,N_20784);
nand U21408 (N_21408,N_20715,N_21179);
xor U21409 (N_21409,N_21163,N_21061);
xor U21410 (N_21410,N_21018,N_21027);
nor U21411 (N_21411,N_20909,N_20838);
nor U21412 (N_21412,N_21115,N_20634);
xnor U21413 (N_21413,N_20740,N_21223);
nand U21414 (N_21414,N_20937,N_20729);
xnor U21415 (N_21415,N_20676,N_21154);
or U21416 (N_21416,N_20901,N_20986);
xnor U21417 (N_21417,N_20990,N_20873);
or U21418 (N_21418,N_20722,N_20881);
xor U21419 (N_21419,N_21235,N_20824);
nand U21420 (N_21420,N_20709,N_20924);
xnor U21421 (N_21421,N_21131,N_21182);
nand U21422 (N_21422,N_21207,N_20663);
xnor U21423 (N_21423,N_20945,N_20964);
and U21424 (N_21424,N_20822,N_21198);
nand U21425 (N_21425,N_21059,N_20770);
and U21426 (N_21426,N_20726,N_20764);
nor U21427 (N_21427,N_20771,N_21217);
and U21428 (N_21428,N_20682,N_21211);
or U21429 (N_21429,N_21024,N_21187);
nor U21430 (N_21430,N_21066,N_21225);
and U21431 (N_21431,N_21224,N_21156);
or U21432 (N_21432,N_21159,N_20959);
or U21433 (N_21433,N_21067,N_20693);
or U21434 (N_21434,N_20707,N_20902);
nand U21435 (N_21435,N_21161,N_20955);
nor U21436 (N_21436,N_20743,N_21193);
nor U21437 (N_21437,N_20989,N_21098);
nor U21438 (N_21438,N_21011,N_21052);
and U21439 (N_21439,N_21075,N_20883);
and U21440 (N_21440,N_20874,N_20804);
and U21441 (N_21441,N_21056,N_20837);
nor U21442 (N_21442,N_20738,N_20661);
nor U21443 (N_21443,N_21040,N_21111);
and U21444 (N_21444,N_20928,N_21007);
xnor U21445 (N_21445,N_21190,N_21137);
nor U21446 (N_21446,N_21076,N_20842);
nor U21447 (N_21447,N_20657,N_20875);
and U21448 (N_21448,N_20877,N_20660);
nand U21449 (N_21449,N_20917,N_20669);
and U21450 (N_21450,N_20833,N_21192);
nor U21451 (N_21451,N_21158,N_20897);
xor U21452 (N_21452,N_20899,N_21101);
nand U21453 (N_21453,N_21016,N_20789);
nand U21454 (N_21454,N_20965,N_20996);
nand U21455 (N_21455,N_21169,N_20639);
nand U21456 (N_21456,N_20885,N_20805);
nand U21457 (N_21457,N_21199,N_21153);
and U21458 (N_21458,N_21090,N_20920);
xor U21459 (N_21459,N_21117,N_21096);
and U21460 (N_21460,N_21086,N_20793);
nor U21461 (N_21461,N_20797,N_21095);
xor U21462 (N_21462,N_20973,N_21185);
and U21463 (N_21463,N_21001,N_20827);
xnor U21464 (N_21464,N_20856,N_20814);
or U21465 (N_21465,N_21219,N_20816);
or U21466 (N_21466,N_20845,N_21092);
nand U21467 (N_21467,N_20882,N_21171);
nand U21468 (N_21468,N_21036,N_20658);
and U21469 (N_21469,N_20642,N_21195);
nor U21470 (N_21470,N_20847,N_20854);
nand U21471 (N_21471,N_21051,N_20794);
and U21472 (N_21472,N_20752,N_20832);
nand U21473 (N_21473,N_20815,N_20679);
nor U21474 (N_21474,N_20688,N_21209);
nand U21475 (N_21475,N_21081,N_21226);
and U21476 (N_21476,N_20999,N_20866);
nand U21477 (N_21477,N_21049,N_20769);
nand U21478 (N_21478,N_20995,N_20865);
nor U21479 (N_21479,N_21073,N_21205);
xor U21480 (N_21480,N_20892,N_20678);
xnor U21481 (N_21481,N_20665,N_20850);
or U21482 (N_21482,N_21147,N_21213);
or U21483 (N_21483,N_20813,N_20777);
nand U21484 (N_21484,N_21082,N_20672);
nand U21485 (N_21485,N_21074,N_20802);
or U21486 (N_21486,N_21103,N_20891);
nor U21487 (N_21487,N_20714,N_20704);
nand U21488 (N_21488,N_20627,N_21008);
or U21489 (N_21489,N_21097,N_20895);
or U21490 (N_21490,N_21039,N_21012);
and U21491 (N_21491,N_21140,N_20779);
nand U21492 (N_21492,N_21055,N_20774);
nand U21493 (N_21493,N_21229,N_20773);
and U21494 (N_21494,N_20768,N_20763);
nand U21495 (N_21495,N_21083,N_20708);
nor U21496 (N_21496,N_20727,N_20745);
or U21497 (N_21497,N_21145,N_20916);
nand U21498 (N_21498,N_20651,N_20648);
xor U21499 (N_21499,N_20717,N_21037);
nand U21500 (N_21500,N_21188,N_20808);
nor U21501 (N_21501,N_20954,N_20956);
or U21502 (N_21502,N_20697,N_21132);
nor U21503 (N_21503,N_20836,N_20756);
or U21504 (N_21504,N_21208,N_20692);
or U21505 (N_21505,N_20946,N_20828);
nor U21506 (N_21506,N_20696,N_21085);
and U21507 (N_21507,N_21167,N_20650);
nand U21508 (N_21508,N_21045,N_20767);
xor U21509 (N_21509,N_20835,N_20626);
nor U21510 (N_21510,N_20898,N_20988);
nand U21511 (N_21511,N_20680,N_21013);
nand U21512 (N_21512,N_21050,N_20778);
nor U21513 (N_21513,N_20812,N_21128);
or U21514 (N_21514,N_21239,N_20809);
nand U21515 (N_21515,N_21180,N_20896);
xnor U21516 (N_21516,N_20681,N_20904);
or U21517 (N_21517,N_20953,N_21126);
or U21518 (N_21518,N_21206,N_21009);
or U21519 (N_21519,N_21130,N_21054);
or U21520 (N_21520,N_20991,N_20884);
and U21521 (N_21521,N_21204,N_20636);
nand U21522 (N_21522,N_21227,N_20765);
nand U21523 (N_21523,N_20811,N_20961);
or U21524 (N_21524,N_20834,N_21200);
nand U21525 (N_21525,N_21105,N_20859);
nor U21526 (N_21526,N_20906,N_21100);
and U21527 (N_21527,N_20998,N_20781);
xor U21528 (N_21528,N_20963,N_20633);
nor U21529 (N_21529,N_20677,N_20929);
and U21530 (N_21530,N_21072,N_21230);
or U21531 (N_21531,N_20967,N_21133);
and U21532 (N_21532,N_20628,N_20646);
and U21533 (N_21533,N_20993,N_20792);
or U21534 (N_21534,N_21091,N_20711);
xor U21535 (N_21535,N_21142,N_20724);
nand U21536 (N_21536,N_20983,N_20653);
and U21537 (N_21537,N_20701,N_20962);
xor U21538 (N_21538,N_20934,N_20857);
or U21539 (N_21539,N_21041,N_20783);
xnor U21540 (N_21540,N_20725,N_20807);
nand U21541 (N_21541,N_20638,N_20980);
nor U21542 (N_21542,N_20861,N_20918);
xor U21543 (N_21543,N_21175,N_20903);
and U21544 (N_21544,N_20670,N_20829);
nor U21545 (N_21545,N_21014,N_21231);
xor U21546 (N_21546,N_20780,N_20703);
or U21547 (N_21547,N_21088,N_20728);
and U21548 (N_21548,N_21240,N_21071);
xor U21549 (N_21549,N_20796,N_21210);
or U21550 (N_21550,N_20926,N_21177);
xnor U21551 (N_21551,N_20749,N_20786);
nor U21552 (N_21552,N_21134,N_20862);
xnor U21553 (N_21553,N_20656,N_20974);
xor U21554 (N_21554,N_20853,N_21181);
or U21555 (N_21555,N_21065,N_20723);
and U21556 (N_21556,N_20994,N_20671);
xnor U21557 (N_21557,N_21143,N_20759);
xor U21558 (N_21558,N_20746,N_20958);
xnor U21559 (N_21559,N_21212,N_20825);
nor U21560 (N_21560,N_21242,N_20886);
nand U21561 (N_21561,N_21044,N_21021);
nor U21562 (N_21562,N_21183,N_21049);
and U21563 (N_21563,N_20913,N_21037);
xor U21564 (N_21564,N_20925,N_20918);
or U21565 (N_21565,N_20816,N_20696);
or U21566 (N_21566,N_20841,N_20785);
or U21567 (N_21567,N_20684,N_21068);
nand U21568 (N_21568,N_20986,N_21011);
or U21569 (N_21569,N_21134,N_20836);
nand U21570 (N_21570,N_20788,N_20840);
and U21571 (N_21571,N_21020,N_20674);
or U21572 (N_21572,N_21043,N_21109);
nand U21573 (N_21573,N_21123,N_21173);
and U21574 (N_21574,N_21173,N_21006);
and U21575 (N_21575,N_20846,N_21043);
xor U21576 (N_21576,N_20672,N_20824);
xnor U21577 (N_21577,N_21106,N_20638);
nor U21578 (N_21578,N_21183,N_20774);
or U21579 (N_21579,N_20974,N_20890);
xor U21580 (N_21580,N_20980,N_20848);
nor U21581 (N_21581,N_20853,N_21191);
and U21582 (N_21582,N_20886,N_20991);
or U21583 (N_21583,N_20680,N_21069);
nand U21584 (N_21584,N_21090,N_21148);
xor U21585 (N_21585,N_20897,N_20807);
and U21586 (N_21586,N_20893,N_20914);
xnor U21587 (N_21587,N_21202,N_21036);
or U21588 (N_21588,N_20796,N_21224);
nor U21589 (N_21589,N_20852,N_20756);
and U21590 (N_21590,N_21197,N_20933);
xor U21591 (N_21591,N_20876,N_20702);
xnor U21592 (N_21592,N_21222,N_21107);
nand U21593 (N_21593,N_21018,N_20782);
and U21594 (N_21594,N_20632,N_20942);
xnor U21595 (N_21595,N_21199,N_21184);
and U21596 (N_21596,N_21132,N_21210);
and U21597 (N_21597,N_21215,N_21082);
nor U21598 (N_21598,N_20924,N_20926);
and U21599 (N_21599,N_20712,N_20824);
and U21600 (N_21600,N_20664,N_20934);
nand U21601 (N_21601,N_20728,N_20928);
xor U21602 (N_21602,N_20935,N_20679);
nor U21603 (N_21603,N_20723,N_20796);
or U21604 (N_21604,N_21165,N_20899);
nand U21605 (N_21605,N_21128,N_21011);
xnor U21606 (N_21606,N_21213,N_20785);
xor U21607 (N_21607,N_21233,N_20651);
nand U21608 (N_21608,N_20916,N_21101);
and U21609 (N_21609,N_21004,N_21058);
nor U21610 (N_21610,N_20791,N_20915);
or U21611 (N_21611,N_20904,N_20867);
nand U21612 (N_21612,N_21149,N_20886);
and U21613 (N_21613,N_21138,N_20998);
or U21614 (N_21614,N_20845,N_20835);
and U21615 (N_21615,N_20761,N_20981);
nand U21616 (N_21616,N_21169,N_20886);
nor U21617 (N_21617,N_20686,N_21081);
xor U21618 (N_21618,N_21032,N_21241);
and U21619 (N_21619,N_20760,N_20800);
nor U21620 (N_21620,N_20664,N_21184);
or U21621 (N_21621,N_21061,N_20904);
xor U21622 (N_21622,N_20705,N_20937);
nand U21623 (N_21623,N_20814,N_21099);
xor U21624 (N_21624,N_21226,N_20997);
nand U21625 (N_21625,N_20639,N_20895);
and U21626 (N_21626,N_20875,N_20897);
nand U21627 (N_21627,N_21071,N_21177);
xor U21628 (N_21628,N_20944,N_20725);
or U21629 (N_21629,N_20833,N_20787);
nor U21630 (N_21630,N_21229,N_20730);
and U21631 (N_21631,N_20979,N_21167);
and U21632 (N_21632,N_21064,N_20632);
nand U21633 (N_21633,N_20705,N_20754);
or U21634 (N_21634,N_20870,N_20765);
nor U21635 (N_21635,N_20915,N_21143);
and U21636 (N_21636,N_21026,N_20707);
nand U21637 (N_21637,N_21125,N_20634);
or U21638 (N_21638,N_20810,N_20850);
nor U21639 (N_21639,N_21121,N_21195);
and U21640 (N_21640,N_21033,N_21220);
or U21641 (N_21641,N_20850,N_20646);
and U21642 (N_21642,N_21211,N_20879);
or U21643 (N_21643,N_21175,N_20631);
nand U21644 (N_21644,N_21060,N_21117);
or U21645 (N_21645,N_20929,N_20889);
nand U21646 (N_21646,N_20634,N_20731);
and U21647 (N_21647,N_20937,N_21223);
or U21648 (N_21648,N_21151,N_20872);
nor U21649 (N_21649,N_20756,N_20933);
xnor U21650 (N_21650,N_21132,N_21035);
and U21651 (N_21651,N_21232,N_21144);
and U21652 (N_21652,N_21051,N_20695);
and U21653 (N_21653,N_21062,N_21028);
nor U21654 (N_21654,N_20826,N_21119);
and U21655 (N_21655,N_21194,N_20894);
or U21656 (N_21656,N_21099,N_21049);
nor U21657 (N_21657,N_21107,N_21220);
xor U21658 (N_21658,N_20702,N_20893);
nand U21659 (N_21659,N_21073,N_21240);
xor U21660 (N_21660,N_20954,N_20690);
xor U21661 (N_21661,N_21103,N_21214);
nor U21662 (N_21662,N_20810,N_21133);
or U21663 (N_21663,N_20636,N_20695);
nand U21664 (N_21664,N_20654,N_20823);
and U21665 (N_21665,N_20823,N_21124);
nor U21666 (N_21666,N_20883,N_21181);
nand U21667 (N_21667,N_20730,N_20770);
nor U21668 (N_21668,N_20813,N_20833);
nor U21669 (N_21669,N_20873,N_20763);
nand U21670 (N_21670,N_20738,N_20672);
and U21671 (N_21671,N_20678,N_21118);
or U21672 (N_21672,N_21051,N_20830);
nand U21673 (N_21673,N_21241,N_20896);
and U21674 (N_21674,N_21173,N_20983);
nor U21675 (N_21675,N_20989,N_21175);
nand U21676 (N_21676,N_21033,N_20764);
nand U21677 (N_21677,N_20951,N_21139);
xnor U21678 (N_21678,N_20681,N_20814);
nand U21679 (N_21679,N_21075,N_21229);
or U21680 (N_21680,N_21152,N_20882);
nand U21681 (N_21681,N_20947,N_21068);
xor U21682 (N_21682,N_20662,N_21005);
or U21683 (N_21683,N_21096,N_20911);
nand U21684 (N_21684,N_21077,N_20966);
xnor U21685 (N_21685,N_20970,N_20680);
nor U21686 (N_21686,N_21044,N_21039);
nand U21687 (N_21687,N_20900,N_20899);
nand U21688 (N_21688,N_20771,N_21146);
and U21689 (N_21689,N_20739,N_20991);
or U21690 (N_21690,N_21135,N_20817);
nor U21691 (N_21691,N_20736,N_21172);
nand U21692 (N_21692,N_21081,N_20927);
xnor U21693 (N_21693,N_21149,N_21201);
or U21694 (N_21694,N_21012,N_20923);
nand U21695 (N_21695,N_20964,N_21173);
nor U21696 (N_21696,N_21005,N_21234);
or U21697 (N_21697,N_20791,N_20700);
nand U21698 (N_21698,N_20979,N_21236);
or U21699 (N_21699,N_20890,N_21180);
nand U21700 (N_21700,N_21245,N_21124);
and U21701 (N_21701,N_21071,N_20736);
and U21702 (N_21702,N_20626,N_20709);
and U21703 (N_21703,N_20795,N_21006);
or U21704 (N_21704,N_21133,N_20973);
and U21705 (N_21705,N_21237,N_21022);
nor U21706 (N_21706,N_21213,N_20736);
or U21707 (N_21707,N_21109,N_20936);
nand U21708 (N_21708,N_21139,N_20967);
and U21709 (N_21709,N_20839,N_20738);
xor U21710 (N_21710,N_20982,N_20987);
nor U21711 (N_21711,N_21011,N_21054);
xor U21712 (N_21712,N_21063,N_20806);
nor U21713 (N_21713,N_21173,N_21047);
or U21714 (N_21714,N_21169,N_21153);
xor U21715 (N_21715,N_21091,N_20966);
xor U21716 (N_21716,N_21002,N_21083);
or U21717 (N_21717,N_20810,N_21033);
nor U21718 (N_21718,N_20702,N_20681);
nor U21719 (N_21719,N_21021,N_20849);
or U21720 (N_21720,N_21156,N_20996);
nor U21721 (N_21721,N_20765,N_21072);
nor U21722 (N_21722,N_20974,N_21207);
and U21723 (N_21723,N_21139,N_20914);
and U21724 (N_21724,N_21019,N_21163);
and U21725 (N_21725,N_21142,N_20794);
nand U21726 (N_21726,N_21115,N_20805);
and U21727 (N_21727,N_20983,N_20749);
or U21728 (N_21728,N_21160,N_20752);
nor U21729 (N_21729,N_21109,N_20763);
nand U21730 (N_21730,N_21007,N_21001);
nand U21731 (N_21731,N_20946,N_20922);
and U21732 (N_21732,N_20969,N_20702);
or U21733 (N_21733,N_20645,N_20859);
or U21734 (N_21734,N_21078,N_20699);
nor U21735 (N_21735,N_21232,N_20960);
nor U21736 (N_21736,N_21049,N_20634);
and U21737 (N_21737,N_21091,N_21246);
nor U21738 (N_21738,N_20843,N_21103);
and U21739 (N_21739,N_20979,N_21088);
and U21740 (N_21740,N_21045,N_21221);
nand U21741 (N_21741,N_20997,N_20667);
nor U21742 (N_21742,N_20843,N_20781);
nor U21743 (N_21743,N_20821,N_20869);
nor U21744 (N_21744,N_21241,N_21069);
and U21745 (N_21745,N_20701,N_20777);
xor U21746 (N_21746,N_20857,N_21134);
or U21747 (N_21747,N_20756,N_21237);
xnor U21748 (N_21748,N_20819,N_20739);
and U21749 (N_21749,N_21174,N_21171);
and U21750 (N_21750,N_20728,N_20640);
or U21751 (N_21751,N_21067,N_21118);
nand U21752 (N_21752,N_21175,N_20675);
and U21753 (N_21753,N_20723,N_21189);
nor U21754 (N_21754,N_20682,N_21003);
nand U21755 (N_21755,N_20914,N_20772);
or U21756 (N_21756,N_21018,N_21012);
nor U21757 (N_21757,N_20745,N_21059);
or U21758 (N_21758,N_20930,N_20680);
xnor U21759 (N_21759,N_20868,N_20903);
nand U21760 (N_21760,N_20959,N_20894);
or U21761 (N_21761,N_21093,N_20866);
nor U21762 (N_21762,N_20874,N_20783);
nor U21763 (N_21763,N_21121,N_20958);
nor U21764 (N_21764,N_20843,N_20980);
xor U21765 (N_21765,N_20971,N_20860);
and U21766 (N_21766,N_21039,N_20626);
nand U21767 (N_21767,N_21173,N_20662);
nor U21768 (N_21768,N_20814,N_20743);
xor U21769 (N_21769,N_21182,N_20933);
or U21770 (N_21770,N_21096,N_21007);
xnor U21771 (N_21771,N_20871,N_20741);
and U21772 (N_21772,N_21138,N_21088);
nand U21773 (N_21773,N_21048,N_21123);
nor U21774 (N_21774,N_20995,N_20687);
nor U21775 (N_21775,N_20955,N_20877);
nand U21776 (N_21776,N_20679,N_20798);
nand U21777 (N_21777,N_20733,N_21100);
and U21778 (N_21778,N_21094,N_20721);
xnor U21779 (N_21779,N_21151,N_20845);
or U21780 (N_21780,N_20698,N_20768);
xnor U21781 (N_21781,N_21192,N_21163);
xor U21782 (N_21782,N_20888,N_20942);
xor U21783 (N_21783,N_20647,N_20843);
and U21784 (N_21784,N_20931,N_20755);
nand U21785 (N_21785,N_20657,N_20834);
and U21786 (N_21786,N_20790,N_20732);
nor U21787 (N_21787,N_20675,N_20881);
or U21788 (N_21788,N_20927,N_20872);
nor U21789 (N_21789,N_20967,N_20745);
xnor U21790 (N_21790,N_20992,N_20965);
and U21791 (N_21791,N_21079,N_20899);
nor U21792 (N_21792,N_21084,N_20657);
nand U21793 (N_21793,N_20875,N_20819);
nor U21794 (N_21794,N_21136,N_20764);
and U21795 (N_21795,N_20660,N_21036);
or U21796 (N_21796,N_20637,N_21103);
or U21797 (N_21797,N_20764,N_21101);
nor U21798 (N_21798,N_21033,N_20875);
nor U21799 (N_21799,N_21043,N_20701);
xnor U21800 (N_21800,N_20834,N_21152);
and U21801 (N_21801,N_20876,N_20789);
xnor U21802 (N_21802,N_21043,N_20963);
nor U21803 (N_21803,N_21156,N_21080);
nor U21804 (N_21804,N_21017,N_21123);
nand U21805 (N_21805,N_20873,N_21216);
nand U21806 (N_21806,N_21143,N_20757);
nand U21807 (N_21807,N_20790,N_21104);
nor U21808 (N_21808,N_20727,N_21009);
and U21809 (N_21809,N_21135,N_20980);
and U21810 (N_21810,N_20911,N_21046);
or U21811 (N_21811,N_20793,N_20935);
xor U21812 (N_21812,N_20662,N_21025);
nand U21813 (N_21813,N_20732,N_20680);
and U21814 (N_21814,N_20961,N_20850);
xnor U21815 (N_21815,N_21242,N_21034);
nand U21816 (N_21816,N_21029,N_21009);
nand U21817 (N_21817,N_21128,N_20875);
xor U21818 (N_21818,N_21018,N_21021);
xor U21819 (N_21819,N_20870,N_20823);
or U21820 (N_21820,N_21048,N_21002);
nor U21821 (N_21821,N_20724,N_21043);
and U21822 (N_21822,N_21192,N_20831);
or U21823 (N_21823,N_20752,N_21018);
and U21824 (N_21824,N_21195,N_20959);
and U21825 (N_21825,N_21039,N_21189);
xnor U21826 (N_21826,N_20724,N_21003);
nand U21827 (N_21827,N_20653,N_20913);
nand U21828 (N_21828,N_21122,N_21044);
and U21829 (N_21829,N_21013,N_20833);
or U21830 (N_21830,N_20997,N_20913);
xnor U21831 (N_21831,N_20734,N_20627);
nand U21832 (N_21832,N_20820,N_21138);
or U21833 (N_21833,N_21168,N_21227);
and U21834 (N_21834,N_20646,N_21004);
nand U21835 (N_21835,N_20979,N_20707);
xor U21836 (N_21836,N_20677,N_21183);
or U21837 (N_21837,N_21149,N_20771);
or U21838 (N_21838,N_21189,N_21230);
or U21839 (N_21839,N_21022,N_20921);
and U21840 (N_21840,N_20650,N_20799);
nand U21841 (N_21841,N_20885,N_21081);
xnor U21842 (N_21842,N_20901,N_20687);
or U21843 (N_21843,N_21041,N_20898);
and U21844 (N_21844,N_20695,N_21238);
nor U21845 (N_21845,N_21092,N_21123);
nand U21846 (N_21846,N_21165,N_20844);
or U21847 (N_21847,N_21081,N_20914);
or U21848 (N_21848,N_21211,N_20752);
and U21849 (N_21849,N_20980,N_20764);
nand U21850 (N_21850,N_20874,N_20907);
or U21851 (N_21851,N_21004,N_21174);
or U21852 (N_21852,N_20657,N_20696);
and U21853 (N_21853,N_20760,N_20717);
nor U21854 (N_21854,N_21118,N_21068);
nand U21855 (N_21855,N_20636,N_21144);
xnor U21856 (N_21856,N_21150,N_20652);
nor U21857 (N_21857,N_20905,N_21177);
or U21858 (N_21858,N_20633,N_20859);
and U21859 (N_21859,N_20672,N_21223);
nor U21860 (N_21860,N_21110,N_20804);
nand U21861 (N_21861,N_21192,N_21132);
and U21862 (N_21862,N_21014,N_21237);
and U21863 (N_21863,N_21228,N_20905);
xor U21864 (N_21864,N_21207,N_21236);
and U21865 (N_21865,N_21106,N_21164);
or U21866 (N_21866,N_20710,N_20876);
nor U21867 (N_21867,N_20651,N_20767);
xor U21868 (N_21868,N_20649,N_21050);
xor U21869 (N_21869,N_20825,N_21026);
or U21870 (N_21870,N_20706,N_20670);
nand U21871 (N_21871,N_21229,N_20696);
or U21872 (N_21872,N_21108,N_21129);
xor U21873 (N_21873,N_20797,N_21241);
nor U21874 (N_21874,N_20768,N_20642);
nor U21875 (N_21875,N_21326,N_21733);
or U21876 (N_21876,N_21254,N_21533);
nand U21877 (N_21877,N_21306,N_21697);
xnor U21878 (N_21878,N_21857,N_21447);
nor U21879 (N_21879,N_21856,N_21292);
or U21880 (N_21880,N_21501,N_21524);
nor U21881 (N_21881,N_21453,N_21559);
xnor U21882 (N_21882,N_21390,N_21526);
or U21883 (N_21883,N_21513,N_21627);
and U21884 (N_21884,N_21342,N_21379);
and U21885 (N_21885,N_21839,N_21630);
and U21886 (N_21886,N_21621,N_21723);
nand U21887 (N_21887,N_21400,N_21451);
or U21888 (N_21888,N_21796,N_21869);
nand U21889 (N_21889,N_21589,N_21472);
xor U21890 (N_21890,N_21430,N_21754);
xnor U21891 (N_21891,N_21276,N_21541);
or U21892 (N_21892,N_21789,N_21392);
xor U21893 (N_21893,N_21583,N_21591);
nor U21894 (N_21894,N_21318,N_21574);
xor U21895 (N_21895,N_21721,N_21441);
nor U21896 (N_21896,N_21855,N_21578);
nor U21897 (N_21897,N_21684,N_21614);
xor U21898 (N_21898,N_21289,N_21452);
nand U21899 (N_21899,N_21340,N_21407);
or U21900 (N_21900,N_21562,N_21655);
and U21901 (N_21901,N_21656,N_21794);
and U21902 (N_21902,N_21525,N_21479);
xnor U21903 (N_21903,N_21710,N_21290);
and U21904 (N_21904,N_21553,N_21831);
and U21905 (N_21905,N_21601,N_21722);
nand U21906 (N_21906,N_21256,N_21275);
xor U21907 (N_21907,N_21293,N_21465);
nand U21908 (N_21908,N_21715,N_21409);
nor U21909 (N_21909,N_21671,N_21809);
nor U21910 (N_21910,N_21301,N_21686);
nor U21911 (N_21911,N_21416,N_21548);
and U21912 (N_21912,N_21299,N_21825);
xnor U21913 (N_21913,N_21489,N_21713);
and U21914 (N_21914,N_21724,N_21760);
and U21915 (N_21915,N_21637,N_21444);
nand U21916 (N_21916,N_21519,N_21755);
nor U21917 (N_21917,N_21615,N_21650);
xor U21918 (N_21918,N_21285,N_21620);
nand U21919 (N_21919,N_21450,N_21606);
and U21920 (N_21920,N_21780,N_21458);
and U21921 (N_21921,N_21531,N_21477);
and U21922 (N_21922,N_21257,N_21824);
nand U21923 (N_21923,N_21281,N_21821);
and U21924 (N_21924,N_21491,N_21396);
or U21925 (N_21925,N_21675,N_21813);
xnor U21926 (N_21926,N_21726,N_21467);
xor U21927 (N_21927,N_21797,N_21707);
nor U21928 (N_21928,N_21366,N_21865);
xnor U21929 (N_21929,N_21787,N_21528);
or U21930 (N_21930,N_21308,N_21381);
nor U21931 (N_21931,N_21644,N_21547);
or U21932 (N_21932,N_21349,N_21862);
nor U21933 (N_21933,N_21410,N_21818);
nand U21934 (N_21934,N_21527,N_21463);
xnor U21935 (N_21935,N_21434,N_21420);
nand U21936 (N_21936,N_21832,N_21749);
and U21937 (N_21937,N_21736,N_21339);
xor U21938 (N_21938,N_21763,N_21532);
and U21939 (N_21939,N_21623,N_21297);
xor U21940 (N_21940,N_21508,N_21429);
or U21941 (N_21941,N_21500,N_21629);
and U21942 (N_21942,N_21778,N_21624);
and U21943 (N_21943,N_21835,N_21597);
and U21944 (N_21944,N_21808,N_21584);
nor U21945 (N_21945,N_21350,N_21268);
or U21946 (N_21946,N_21816,N_21571);
xnor U21947 (N_21947,N_21344,N_21545);
and U21948 (N_21948,N_21445,N_21642);
nand U21949 (N_21949,N_21783,N_21505);
nand U21950 (N_21950,N_21555,N_21725);
and U21951 (N_21951,N_21874,N_21564);
nor U21952 (N_21952,N_21628,N_21517);
and U21953 (N_21953,N_21577,N_21674);
and U21954 (N_21954,N_21424,N_21823);
nor U21955 (N_21955,N_21767,N_21422);
or U21956 (N_21956,N_21343,N_21575);
xor U21957 (N_21957,N_21779,N_21556);
or U21958 (N_21958,N_21798,N_21338);
nor U21959 (N_21959,N_21785,N_21603);
xor U21960 (N_21960,N_21534,N_21253);
nor U21961 (N_21961,N_21305,N_21259);
or U21962 (N_21962,N_21827,N_21554);
or U21963 (N_21963,N_21858,N_21661);
nand U21964 (N_21964,N_21511,N_21786);
and U21965 (N_21965,N_21522,N_21427);
nand U21966 (N_21966,N_21323,N_21506);
xnor U21967 (N_21967,N_21481,N_21411);
nor U21968 (N_21968,N_21252,N_21817);
or U21969 (N_21969,N_21509,N_21735);
and U21970 (N_21970,N_21362,N_21595);
xnor U21971 (N_21971,N_21565,N_21593);
xor U21972 (N_21972,N_21746,N_21529);
xor U21973 (N_21973,N_21668,N_21380);
xnor U21974 (N_21974,N_21868,N_21853);
nor U21975 (N_21975,N_21446,N_21776);
xnor U21976 (N_21976,N_21523,N_21731);
nor U21977 (N_21977,N_21382,N_21425);
nor U21978 (N_21978,N_21261,N_21274);
nor U21979 (N_21979,N_21647,N_21829);
or U21980 (N_21980,N_21714,N_21371);
or U21981 (N_21981,N_21795,N_21582);
and U21982 (N_21982,N_21302,N_21499);
or U21983 (N_21983,N_21769,N_21790);
xnor U21984 (N_21984,N_21368,N_21833);
or U21985 (N_21985,N_21360,N_21354);
nor U21986 (N_21986,N_21608,N_21561);
xnor U21987 (N_21987,N_21645,N_21588);
and U21988 (N_21988,N_21557,N_21426);
nand U21989 (N_21989,N_21328,N_21264);
or U21990 (N_21990,N_21456,N_21849);
xor U21991 (N_21991,N_21535,N_21777);
and U21992 (N_21992,N_21581,N_21518);
xnor U21993 (N_21993,N_21639,N_21280);
nor U21994 (N_21994,N_21665,N_21572);
or U21995 (N_21995,N_21706,N_21466);
xnor U21996 (N_21996,N_21325,N_21376);
or U21997 (N_21997,N_21699,N_21311);
nand U21998 (N_21998,N_21596,N_21459);
nand U21999 (N_21999,N_21337,N_21493);
or U22000 (N_22000,N_21830,N_21826);
and U22001 (N_22001,N_21277,N_21842);
nand U22002 (N_22002,N_21544,N_21404);
nor U22003 (N_22003,N_21613,N_21861);
nand U22004 (N_22004,N_21770,N_21258);
xnor U22005 (N_22005,N_21449,N_21805);
or U22006 (N_22006,N_21364,N_21774);
xor U22007 (N_22007,N_21654,N_21345);
nand U22008 (N_22008,N_21841,N_21643);
nor U22009 (N_22009,N_21347,N_21619);
nand U22010 (N_22010,N_21652,N_21622);
or U22011 (N_22011,N_21631,N_21802);
xnor U22012 (N_22012,N_21370,N_21696);
or U22013 (N_22013,N_21440,N_21514);
nand U22014 (N_22014,N_21316,N_21678);
and U22015 (N_22015,N_21483,N_21747);
or U22016 (N_22016,N_21815,N_21346);
nand U22017 (N_22017,N_21719,N_21848);
nor U22018 (N_22018,N_21634,N_21616);
nand U22019 (N_22019,N_21867,N_21618);
nor U22020 (N_22020,N_21384,N_21413);
xnor U22021 (N_22021,N_21437,N_21367);
or U22022 (N_22022,N_21663,N_21375);
or U22023 (N_22023,N_21324,N_21859);
xnor U22024 (N_22024,N_21487,N_21579);
nor U22025 (N_22025,N_21373,N_21419);
nor U22026 (N_22026,N_21872,N_21516);
nor U22027 (N_22027,N_21502,N_21317);
nor U22028 (N_22028,N_21609,N_21695);
nor U22029 (N_22029,N_21845,N_21335);
xnor U22030 (N_22030,N_21611,N_21498);
nor U22031 (N_22031,N_21474,N_21469);
xnor U22032 (N_22032,N_21334,N_21700);
or U22033 (N_22033,N_21540,N_21667);
nor U22034 (N_22034,N_21729,N_21740);
xnor U22035 (N_22035,N_21438,N_21415);
xnor U22036 (N_22036,N_21843,N_21551);
xnor U22037 (N_22037,N_21745,N_21473);
and U22038 (N_22038,N_21846,N_21357);
xor U22039 (N_22039,N_21383,N_21727);
and U22040 (N_22040,N_21295,N_21587);
and U22041 (N_22041,N_21560,N_21333);
and U22042 (N_22042,N_21393,N_21310);
nand U22043 (N_22043,N_21432,N_21679);
xnor U22044 (N_22044,N_21685,N_21819);
or U22045 (N_22045,N_21309,N_21687);
or U22046 (N_22046,N_21454,N_21761);
or U22047 (N_22047,N_21286,N_21507);
or U22048 (N_22048,N_21395,N_21494);
nor U22049 (N_22049,N_21298,N_21646);
nor U22050 (N_22050,N_21369,N_21542);
and U22051 (N_22051,N_21475,N_21568);
or U22052 (N_22052,N_21476,N_21741);
nand U22053 (N_22053,N_21329,N_21462);
and U22054 (N_22054,N_21355,N_21436);
or U22055 (N_22055,N_21739,N_21756);
or U22056 (N_22056,N_21319,N_21864);
nand U22057 (N_22057,N_21401,N_21693);
and U22058 (N_22058,N_21510,N_21418);
nand U22059 (N_22059,N_21636,N_21635);
and U22060 (N_22060,N_21269,N_21402);
nand U22061 (N_22061,N_21417,N_21734);
and U22062 (N_22062,N_21870,N_21775);
and U22063 (N_22063,N_21492,N_21590);
xnor U22064 (N_22064,N_21536,N_21708);
nand U22065 (N_22065,N_21398,N_21773);
xnor U22066 (N_22066,N_21336,N_21657);
nor U22067 (N_22067,N_21464,N_21251);
nand U22068 (N_22068,N_21847,N_21496);
nor U22069 (N_22069,N_21300,N_21272);
or U22070 (N_22070,N_21680,N_21312);
nand U22071 (N_22071,N_21712,N_21352);
xor U22072 (N_22072,N_21852,N_21602);
nor U22073 (N_22073,N_21698,N_21651);
nor U22074 (N_22074,N_21677,N_21626);
nor U22075 (N_22075,N_21716,N_21653);
nand U22076 (N_22076,N_21828,N_21604);
nand U22077 (N_22077,N_21648,N_21358);
or U22078 (N_22078,N_21497,N_21666);
xnor U22079 (N_22079,N_21807,N_21543);
and U22080 (N_22080,N_21690,N_21353);
nand U22081 (N_22081,N_21361,N_21633);
nor U22082 (N_22082,N_21428,N_21530);
nand U22083 (N_22083,N_21388,N_21711);
xor U22084 (N_22084,N_21810,N_21662);
nand U22085 (N_22085,N_21279,N_21598);
nor U22086 (N_22086,N_21488,N_21546);
nand U22087 (N_22087,N_21801,N_21263);
xnor U22088 (N_22088,N_21372,N_21688);
or U22089 (N_22089,N_21737,N_21610);
nor U22090 (N_22090,N_21752,N_21750);
xnor U22091 (N_22091,N_21512,N_21822);
nor U22092 (N_22092,N_21768,N_21592);
nor U22093 (N_22093,N_21641,N_21757);
and U22094 (N_22094,N_21717,N_21423);
nor U22095 (N_22095,N_21470,N_21387);
or U22096 (N_22096,N_21580,N_21320);
or U22097 (N_22097,N_21649,N_21332);
nor U22098 (N_22098,N_21594,N_21266);
nand U22099 (N_22099,N_21386,N_21781);
or U22100 (N_22100,N_21408,N_21341);
xnor U22101 (N_22101,N_21632,N_21799);
or U22102 (N_22102,N_21573,N_21558);
or U22103 (N_22103,N_21330,N_21854);
nand U22104 (N_22104,N_21600,N_21442);
nand U22105 (N_22105,N_21322,N_21840);
xnor U22106 (N_22106,N_21265,N_21730);
xnor U22107 (N_22107,N_21471,N_21307);
nand U22108 (N_22108,N_21670,N_21457);
nor U22109 (N_22109,N_21267,N_21549);
nand U22110 (N_22110,N_21570,N_21503);
or U22111 (N_22111,N_21638,N_21435);
nand U22112 (N_22112,N_21394,N_21748);
and U22113 (N_22113,N_21566,N_21814);
xor U22114 (N_22114,N_21738,N_21296);
xor U22115 (N_22115,N_21758,N_21692);
or U22116 (N_22116,N_21836,N_21672);
nor U22117 (N_22117,N_21676,N_21625);
xor U22118 (N_22118,N_21351,N_21374);
and U22119 (N_22119,N_21837,N_21691);
and U22120 (N_22120,N_21270,N_21607);
xnor U22121 (N_22121,N_21703,N_21315);
nand U22122 (N_22122,N_21771,N_21460);
and U22123 (N_22123,N_21850,N_21260);
and U22124 (N_22124,N_21397,N_21385);
and U22125 (N_22125,N_21284,N_21569);
nand U22126 (N_22126,N_21294,N_21811);
nand U22127 (N_22127,N_21820,N_21673);
xnor U22128 (N_22128,N_21288,N_21521);
and U22129 (N_22129,N_21718,N_21433);
and U22130 (N_22130,N_21537,N_21478);
and U22131 (N_22131,N_21412,N_21389);
or U22132 (N_22132,N_21331,N_21448);
and U22133 (N_22133,N_21866,N_21403);
and U22134 (N_22134,N_21863,N_21782);
nand U22135 (N_22135,N_21273,N_21694);
nor U22136 (N_22136,N_21728,N_21791);
or U22137 (N_22137,N_21664,N_21439);
xor U22138 (N_22138,N_21250,N_21443);
xnor U22139 (N_22139,N_21313,N_21844);
nor U22140 (N_22140,N_21480,N_21490);
nand U22141 (N_22141,N_21406,N_21405);
and U22142 (N_22142,N_21262,N_21485);
or U22143 (N_22143,N_21359,N_21399);
xnor U22144 (N_22144,N_21431,N_21804);
or U22145 (N_22145,N_21486,N_21659);
or U22146 (N_22146,N_21793,N_21660);
or U22147 (N_22147,N_21303,N_21585);
nor U22148 (N_22148,N_21291,N_21378);
or U22149 (N_22149,N_21586,N_21538);
nor U22150 (N_22150,N_21468,N_21484);
nor U22151 (N_22151,N_21834,N_21658);
xnor U22152 (N_22152,N_21576,N_21742);
nor U22153 (N_22153,N_21806,N_21838);
xor U22154 (N_22154,N_21304,N_21744);
and U22155 (N_22155,N_21520,N_21873);
and U22156 (N_22156,N_21504,N_21515);
nor U22157 (N_22157,N_21683,N_21539);
or U22158 (N_22158,N_21640,N_21482);
nor U22159 (N_22159,N_21552,N_21803);
or U22160 (N_22160,N_21702,N_21377);
nor U22161 (N_22161,N_21414,N_21563);
nand U22162 (N_22162,N_21681,N_21321);
xnor U22163 (N_22163,N_21283,N_21709);
xor U22164 (N_22164,N_21759,N_21365);
xnor U22165 (N_22165,N_21788,N_21282);
xor U22166 (N_22166,N_21356,N_21766);
nand U22167 (N_22167,N_21753,N_21669);
nand U22168 (N_22168,N_21732,N_21287);
xnor U22169 (N_22169,N_21851,N_21762);
xor U22170 (N_22170,N_21772,N_21765);
or U22171 (N_22171,N_21455,N_21495);
nor U22172 (N_22172,N_21871,N_21599);
nand U22173 (N_22173,N_21461,N_21720);
nand U22174 (N_22174,N_21421,N_21800);
xnor U22175 (N_22175,N_21314,N_21704);
and U22176 (N_22176,N_21682,N_21705);
nand U22177 (N_22177,N_21278,N_21617);
nor U22178 (N_22178,N_21860,N_21751);
xor U22179 (N_22179,N_21764,N_21271);
or U22180 (N_22180,N_21792,N_21255);
xnor U22181 (N_22181,N_21743,N_21605);
or U22182 (N_22182,N_21348,N_21701);
nor U22183 (N_22183,N_21363,N_21391);
nor U22184 (N_22184,N_21784,N_21327);
or U22185 (N_22185,N_21567,N_21612);
and U22186 (N_22186,N_21550,N_21689);
nor U22187 (N_22187,N_21812,N_21329);
nor U22188 (N_22188,N_21424,N_21707);
xnor U22189 (N_22189,N_21851,N_21790);
nand U22190 (N_22190,N_21321,N_21480);
and U22191 (N_22191,N_21826,N_21350);
xor U22192 (N_22192,N_21443,N_21857);
xnor U22193 (N_22193,N_21682,N_21708);
nand U22194 (N_22194,N_21468,N_21322);
nand U22195 (N_22195,N_21848,N_21382);
nor U22196 (N_22196,N_21860,N_21667);
xnor U22197 (N_22197,N_21468,N_21828);
nor U22198 (N_22198,N_21761,N_21656);
or U22199 (N_22199,N_21394,N_21341);
nor U22200 (N_22200,N_21461,N_21713);
xnor U22201 (N_22201,N_21336,N_21844);
nand U22202 (N_22202,N_21844,N_21318);
nand U22203 (N_22203,N_21843,N_21620);
nor U22204 (N_22204,N_21606,N_21281);
or U22205 (N_22205,N_21296,N_21469);
nand U22206 (N_22206,N_21851,N_21524);
nor U22207 (N_22207,N_21850,N_21263);
or U22208 (N_22208,N_21265,N_21844);
nand U22209 (N_22209,N_21291,N_21711);
xnor U22210 (N_22210,N_21705,N_21557);
or U22211 (N_22211,N_21862,N_21611);
nor U22212 (N_22212,N_21714,N_21779);
nand U22213 (N_22213,N_21677,N_21523);
xnor U22214 (N_22214,N_21614,N_21674);
or U22215 (N_22215,N_21604,N_21563);
and U22216 (N_22216,N_21687,N_21496);
xor U22217 (N_22217,N_21259,N_21488);
or U22218 (N_22218,N_21758,N_21795);
and U22219 (N_22219,N_21677,N_21468);
nor U22220 (N_22220,N_21826,N_21748);
xnor U22221 (N_22221,N_21562,N_21280);
xor U22222 (N_22222,N_21350,N_21482);
nand U22223 (N_22223,N_21762,N_21613);
xnor U22224 (N_22224,N_21632,N_21503);
xnor U22225 (N_22225,N_21292,N_21644);
and U22226 (N_22226,N_21559,N_21409);
nor U22227 (N_22227,N_21558,N_21675);
nor U22228 (N_22228,N_21546,N_21521);
or U22229 (N_22229,N_21630,N_21358);
nor U22230 (N_22230,N_21283,N_21723);
nand U22231 (N_22231,N_21690,N_21363);
nor U22232 (N_22232,N_21268,N_21654);
nor U22233 (N_22233,N_21299,N_21705);
xnor U22234 (N_22234,N_21364,N_21450);
nand U22235 (N_22235,N_21480,N_21461);
xor U22236 (N_22236,N_21746,N_21539);
and U22237 (N_22237,N_21570,N_21455);
xor U22238 (N_22238,N_21687,N_21320);
or U22239 (N_22239,N_21301,N_21278);
nand U22240 (N_22240,N_21300,N_21655);
or U22241 (N_22241,N_21330,N_21361);
and U22242 (N_22242,N_21839,N_21349);
and U22243 (N_22243,N_21380,N_21275);
nor U22244 (N_22244,N_21329,N_21544);
and U22245 (N_22245,N_21600,N_21541);
and U22246 (N_22246,N_21427,N_21704);
xor U22247 (N_22247,N_21454,N_21569);
xnor U22248 (N_22248,N_21664,N_21298);
nor U22249 (N_22249,N_21610,N_21467);
nand U22250 (N_22250,N_21831,N_21378);
nor U22251 (N_22251,N_21661,N_21592);
and U22252 (N_22252,N_21587,N_21412);
and U22253 (N_22253,N_21366,N_21356);
nor U22254 (N_22254,N_21636,N_21334);
or U22255 (N_22255,N_21263,N_21613);
xnor U22256 (N_22256,N_21763,N_21787);
nor U22257 (N_22257,N_21374,N_21421);
xnor U22258 (N_22258,N_21357,N_21340);
xor U22259 (N_22259,N_21565,N_21546);
or U22260 (N_22260,N_21462,N_21803);
and U22261 (N_22261,N_21631,N_21508);
nand U22262 (N_22262,N_21252,N_21837);
and U22263 (N_22263,N_21816,N_21689);
nor U22264 (N_22264,N_21330,N_21749);
nor U22265 (N_22265,N_21627,N_21780);
or U22266 (N_22266,N_21420,N_21717);
or U22267 (N_22267,N_21309,N_21741);
and U22268 (N_22268,N_21266,N_21281);
nor U22269 (N_22269,N_21673,N_21345);
xnor U22270 (N_22270,N_21791,N_21619);
nand U22271 (N_22271,N_21454,N_21519);
nand U22272 (N_22272,N_21493,N_21314);
or U22273 (N_22273,N_21723,N_21659);
nor U22274 (N_22274,N_21450,N_21401);
or U22275 (N_22275,N_21477,N_21788);
nor U22276 (N_22276,N_21825,N_21284);
nand U22277 (N_22277,N_21277,N_21626);
and U22278 (N_22278,N_21315,N_21333);
or U22279 (N_22279,N_21766,N_21317);
nor U22280 (N_22280,N_21366,N_21851);
or U22281 (N_22281,N_21463,N_21757);
nor U22282 (N_22282,N_21383,N_21554);
nor U22283 (N_22283,N_21526,N_21336);
xor U22284 (N_22284,N_21558,N_21661);
and U22285 (N_22285,N_21370,N_21560);
xnor U22286 (N_22286,N_21393,N_21263);
xor U22287 (N_22287,N_21510,N_21809);
nand U22288 (N_22288,N_21852,N_21490);
and U22289 (N_22289,N_21718,N_21786);
and U22290 (N_22290,N_21787,N_21706);
nand U22291 (N_22291,N_21427,N_21273);
nand U22292 (N_22292,N_21594,N_21472);
xnor U22293 (N_22293,N_21774,N_21475);
nor U22294 (N_22294,N_21491,N_21455);
xor U22295 (N_22295,N_21770,N_21822);
and U22296 (N_22296,N_21802,N_21521);
or U22297 (N_22297,N_21254,N_21832);
nor U22298 (N_22298,N_21307,N_21856);
nand U22299 (N_22299,N_21529,N_21269);
or U22300 (N_22300,N_21457,N_21422);
and U22301 (N_22301,N_21375,N_21708);
nor U22302 (N_22302,N_21655,N_21347);
or U22303 (N_22303,N_21309,N_21684);
nor U22304 (N_22304,N_21643,N_21442);
xnor U22305 (N_22305,N_21287,N_21606);
nor U22306 (N_22306,N_21697,N_21405);
and U22307 (N_22307,N_21599,N_21553);
and U22308 (N_22308,N_21802,N_21257);
nand U22309 (N_22309,N_21673,N_21404);
nor U22310 (N_22310,N_21723,N_21791);
or U22311 (N_22311,N_21795,N_21464);
nor U22312 (N_22312,N_21864,N_21451);
or U22313 (N_22313,N_21612,N_21304);
nand U22314 (N_22314,N_21764,N_21479);
and U22315 (N_22315,N_21736,N_21707);
xor U22316 (N_22316,N_21626,N_21483);
or U22317 (N_22317,N_21646,N_21475);
xnor U22318 (N_22318,N_21434,N_21360);
and U22319 (N_22319,N_21584,N_21411);
or U22320 (N_22320,N_21615,N_21527);
xnor U22321 (N_22321,N_21548,N_21290);
nor U22322 (N_22322,N_21308,N_21857);
nor U22323 (N_22323,N_21772,N_21741);
nand U22324 (N_22324,N_21481,N_21793);
and U22325 (N_22325,N_21253,N_21345);
or U22326 (N_22326,N_21777,N_21829);
xnor U22327 (N_22327,N_21814,N_21874);
xnor U22328 (N_22328,N_21853,N_21860);
nand U22329 (N_22329,N_21373,N_21536);
xnor U22330 (N_22330,N_21341,N_21515);
nand U22331 (N_22331,N_21396,N_21401);
nor U22332 (N_22332,N_21367,N_21291);
xor U22333 (N_22333,N_21626,N_21865);
nor U22334 (N_22334,N_21259,N_21400);
or U22335 (N_22335,N_21463,N_21423);
xnor U22336 (N_22336,N_21761,N_21456);
or U22337 (N_22337,N_21645,N_21426);
or U22338 (N_22338,N_21659,N_21745);
nor U22339 (N_22339,N_21821,N_21671);
nand U22340 (N_22340,N_21835,N_21665);
xor U22341 (N_22341,N_21780,N_21471);
or U22342 (N_22342,N_21694,N_21553);
nor U22343 (N_22343,N_21790,N_21861);
and U22344 (N_22344,N_21720,N_21433);
nor U22345 (N_22345,N_21509,N_21254);
nor U22346 (N_22346,N_21517,N_21663);
and U22347 (N_22347,N_21250,N_21641);
nor U22348 (N_22348,N_21419,N_21606);
nand U22349 (N_22349,N_21396,N_21870);
nor U22350 (N_22350,N_21861,N_21606);
xor U22351 (N_22351,N_21643,N_21343);
and U22352 (N_22352,N_21327,N_21360);
nor U22353 (N_22353,N_21762,N_21284);
and U22354 (N_22354,N_21352,N_21658);
nor U22355 (N_22355,N_21784,N_21806);
and U22356 (N_22356,N_21843,N_21860);
and U22357 (N_22357,N_21332,N_21721);
and U22358 (N_22358,N_21617,N_21634);
nand U22359 (N_22359,N_21445,N_21314);
xor U22360 (N_22360,N_21495,N_21354);
xor U22361 (N_22361,N_21649,N_21450);
nand U22362 (N_22362,N_21688,N_21589);
nand U22363 (N_22363,N_21344,N_21281);
nand U22364 (N_22364,N_21490,N_21344);
and U22365 (N_22365,N_21854,N_21743);
or U22366 (N_22366,N_21294,N_21473);
xnor U22367 (N_22367,N_21637,N_21579);
xnor U22368 (N_22368,N_21516,N_21484);
xnor U22369 (N_22369,N_21559,N_21627);
or U22370 (N_22370,N_21813,N_21359);
or U22371 (N_22371,N_21355,N_21317);
or U22372 (N_22372,N_21600,N_21533);
nor U22373 (N_22373,N_21422,N_21315);
and U22374 (N_22374,N_21588,N_21378);
or U22375 (N_22375,N_21538,N_21867);
nor U22376 (N_22376,N_21792,N_21728);
and U22377 (N_22377,N_21405,N_21408);
nand U22378 (N_22378,N_21381,N_21598);
and U22379 (N_22379,N_21508,N_21848);
or U22380 (N_22380,N_21867,N_21781);
nand U22381 (N_22381,N_21522,N_21683);
or U22382 (N_22382,N_21429,N_21479);
and U22383 (N_22383,N_21352,N_21753);
xnor U22384 (N_22384,N_21777,N_21427);
nor U22385 (N_22385,N_21502,N_21472);
nand U22386 (N_22386,N_21406,N_21599);
nand U22387 (N_22387,N_21252,N_21360);
and U22388 (N_22388,N_21765,N_21468);
xor U22389 (N_22389,N_21525,N_21444);
or U22390 (N_22390,N_21260,N_21686);
xor U22391 (N_22391,N_21403,N_21395);
and U22392 (N_22392,N_21397,N_21564);
nor U22393 (N_22393,N_21347,N_21448);
xor U22394 (N_22394,N_21622,N_21557);
nand U22395 (N_22395,N_21601,N_21583);
nand U22396 (N_22396,N_21594,N_21602);
and U22397 (N_22397,N_21552,N_21588);
nor U22398 (N_22398,N_21517,N_21820);
nor U22399 (N_22399,N_21537,N_21540);
and U22400 (N_22400,N_21387,N_21805);
nor U22401 (N_22401,N_21516,N_21874);
xnor U22402 (N_22402,N_21558,N_21549);
or U22403 (N_22403,N_21832,N_21696);
nor U22404 (N_22404,N_21642,N_21779);
nand U22405 (N_22405,N_21361,N_21769);
or U22406 (N_22406,N_21317,N_21468);
xnor U22407 (N_22407,N_21502,N_21496);
or U22408 (N_22408,N_21416,N_21546);
and U22409 (N_22409,N_21627,N_21750);
nand U22410 (N_22410,N_21838,N_21534);
nor U22411 (N_22411,N_21838,N_21664);
nor U22412 (N_22412,N_21391,N_21488);
nand U22413 (N_22413,N_21686,N_21843);
nor U22414 (N_22414,N_21601,N_21580);
and U22415 (N_22415,N_21751,N_21431);
xor U22416 (N_22416,N_21615,N_21789);
or U22417 (N_22417,N_21704,N_21385);
and U22418 (N_22418,N_21425,N_21275);
nor U22419 (N_22419,N_21504,N_21715);
or U22420 (N_22420,N_21346,N_21794);
nand U22421 (N_22421,N_21808,N_21611);
or U22422 (N_22422,N_21686,N_21385);
and U22423 (N_22423,N_21752,N_21854);
nor U22424 (N_22424,N_21813,N_21394);
or U22425 (N_22425,N_21375,N_21634);
nand U22426 (N_22426,N_21562,N_21328);
nand U22427 (N_22427,N_21317,N_21586);
xor U22428 (N_22428,N_21525,N_21313);
xnor U22429 (N_22429,N_21760,N_21603);
xor U22430 (N_22430,N_21281,N_21507);
nor U22431 (N_22431,N_21801,N_21458);
and U22432 (N_22432,N_21422,N_21544);
nand U22433 (N_22433,N_21746,N_21600);
or U22434 (N_22434,N_21646,N_21649);
or U22435 (N_22435,N_21749,N_21421);
nor U22436 (N_22436,N_21617,N_21546);
and U22437 (N_22437,N_21717,N_21417);
nor U22438 (N_22438,N_21294,N_21349);
and U22439 (N_22439,N_21729,N_21631);
or U22440 (N_22440,N_21790,N_21365);
nor U22441 (N_22441,N_21863,N_21294);
nor U22442 (N_22442,N_21541,N_21396);
and U22443 (N_22443,N_21869,N_21790);
xor U22444 (N_22444,N_21347,N_21263);
or U22445 (N_22445,N_21275,N_21492);
nand U22446 (N_22446,N_21386,N_21570);
nor U22447 (N_22447,N_21641,N_21654);
nand U22448 (N_22448,N_21477,N_21573);
or U22449 (N_22449,N_21703,N_21351);
and U22450 (N_22450,N_21809,N_21662);
or U22451 (N_22451,N_21379,N_21540);
or U22452 (N_22452,N_21520,N_21603);
xor U22453 (N_22453,N_21419,N_21775);
nand U22454 (N_22454,N_21554,N_21570);
nor U22455 (N_22455,N_21726,N_21417);
or U22456 (N_22456,N_21848,N_21770);
and U22457 (N_22457,N_21736,N_21785);
and U22458 (N_22458,N_21387,N_21688);
nand U22459 (N_22459,N_21300,N_21804);
or U22460 (N_22460,N_21314,N_21786);
xor U22461 (N_22461,N_21331,N_21521);
nor U22462 (N_22462,N_21730,N_21583);
or U22463 (N_22463,N_21846,N_21550);
nor U22464 (N_22464,N_21416,N_21814);
or U22465 (N_22465,N_21427,N_21610);
xnor U22466 (N_22466,N_21733,N_21402);
nand U22467 (N_22467,N_21285,N_21858);
xnor U22468 (N_22468,N_21325,N_21576);
nand U22469 (N_22469,N_21492,N_21807);
nor U22470 (N_22470,N_21594,N_21827);
nor U22471 (N_22471,N_21448,N_21563);
and U22472 (N_22472,N_21754,N_21685);
nand U22473 (N_22473,N_21353,N_21709);
or U22474 (N_22474,N_21432,N_21348);
xor U22475 (N_22475,N_21411,N_21649);
xor U22476 (N_22476,N_21461,N_21583);
nand U22477 (N_22477,N_21839,N_21343);
or U22478 (N_22478,N_21610,N_21340);
xor U22479 (N_22479,N_21628,N_21510);
xnor U22480 (N_22480,N_21376,N_21634);
and U22481 (N_22481,N_21835,N_21463);
and U22482 (N_22482,N_21360,N_21297);
nor U22483 (N_22483,N_21781,N_21612);
xor U22484 (N_22484,N_21819,N_21347);
xor U22485 (N_22485,N_21788,N_21551);
xnor U22486 (N_22486,N_21801,N_21829);
nand U22487 (N_22487,N_21646,N_21644);
nand U22488 (N_22488,N_21624,N_21491);
and U22489 (N_22489,N_21470,N_21550);
nand U22490 (N_22490,N_21790,N_21404);
or U22491 (N_22491,N_21380,N_21737);
nand U22492 (N_22492,N_21345,N_21467);
or U22493 (N_22493,N_21741,N_21575);
xnor U22494 (N_22494,N_21435,N_21482);
xor U22495 (N_22495,N_21570,N_21311);
and U22496 (N_22496,N_21341,N_21840);
and U22497 (N_22497,N_21673,N_21504);
and U22498 (N_22498,N_21411,N_21560);
and U22499 (N_22499,N_21548,N_21328);
nor U22500 (N_22500,N_22097,N_22155);
or U22501 (N_22501,N_21932,N_22242);
nand U22502 (N_22502,N_22241,N_22380);
xor U22503 (N_22503,N_21901,N_21941);
or U22504 (N_22504,N_22281,N_22215);
xnor U22505 (N_22505,N_22039,N_22295);
and U22506 (N_22506,N_22230,N_22382);
nor U22507 (N_22507,N_22287,N_22182);
or U22508 (N_22508,N_22361,N_22290);
nor U22509 (N_22509,N_22465,N_22112);
and U22510 (N_22510,N_22359,N_22147);
and U22511 (N_22511,N_22001,N_22398);
and U22512 (N_22512,N_22036,N_22114);
and U22513 (N_22513,N_22096,N_22058);
or U22514 (N_22514,N_22332,N_21951);
and U22515 (N_22515,N_22404,N_22499);
or U22516 (N_22516,N_21948,N_22354);
or U22517 (N_22517,N_22303,N_21890);
nand U22518 (N_22518,N_22231,N_21883);
xnor U22519 (N_22519,N_21986,N_22308);
nor U22520 (N_22520,N_21905,N_22024);
and U22521 (N_22521,N_22268,N_22366);
and U22522 (N_22522,N_22098,N_22353);
xnor U22523 (N_22523,N_22105,N_21975);
nor U22524 (N_22524,N_21985,N_21997);
or U22525 (N_22525,N_21884,N_21909);
or U22526 (N_22526,N_22343,N_22048);
nand U22527 (N_22527,N_22015,N_21968);
nor U22528 (N_22528,N_22176,N_22408);
xnor U22529 (N_22529,N_22314,N_22468);
xor U22530 (N_22530,N_21919,N_22031);
nand U22531 (N_22531,N_22175,N_22012);
nand U22532 (N_22532,N_21913,N_22466);
xor U22533 (N_22533,N_21914,N_22306);
and U22534 (N_22534,N_21952,N_22104);
or U22535 (N_22535,N_22291,N_22209);
and U22536 (N_22536,N_22235,N_22134);
xor U22537 (N_22537,N_22208,N_22035);
or U22538 (N_22538,N_21878,N_22158);
xnor U22539 (N_22539,N_21895,N_21931);
nand U22540 (N_22540,N_22243,N_22463);
nand U22541 (N_22541,N_22055,N_22373);
and U22542 (N_22542,N_22128,N_22172);
and U22543 (N_22543,N_22467,N_22420);
or U22544 (N_22544,N_22334,N_22063);
or U22545 (N_22545,N_22103,N_22118);
or U22546 (N_22546,N_22294,N_21927);
or U22547 (N_22547,N_22119,N_22014);
nor U22548 (N_22548,N_22296,N_21904);
and U22549 (N_22549,N_22122,N_22411);
xor U22550 (N_22550,N_21908,N_22106);
nor U22551 (N_22551,N_21998,N_22086);
nor U22552 (N_22552,N_22304,N_22260);
or U22553 (N_22553,N_22137,N_22358);
nor U22554 (N_22554,N_21924,N_22427);
nor U22555 (N_22555,N_22405,N_22084);
nor U22556 (N_22556,N_22222,N_22418);
or U22557 (N_22557,N_22356,N_22444);
xor U22558 (N_22558,N_22335,N_22191);
or U22559 (N_22559,N_21911,N_22214);
or U22560 (N_22560,N_22037,N_22348);
xnor U22561 (N_22561,N_22102,N_22280);
nor U22562 (N_22562,N_22376,N_22384);
nand U22563 (N_22563,N_21921,N_21926);
or U22564 (N_22564,N_22328,N_22113);
nor U22565 (N_22565,N_22099,N_22350);
nor U22566 (N_22566,N_22141,N_22347);
nand U22567 (N_22567,N_22310,N_22254);
and U22568 (N_22568,N_21888,N_21950);
nor U22569 (N_22569,N_22056,N_22364);
nand U22570 (N_22570,N_22046,N_22370);
xnor U22571 (N_22571,N_22441,N_21945);
and U22572 (N_22572,N_22093,N_22041);
nand U22573 (N_22573,N_22388,N_22409);
xor U22574 (N_22574,N_22205,N_22477);
xor U22575 (N_22575,N_22018,N_21922);
or U22576 (N_22576,N_21896,N_22166);
nor U22577 (N_22577,N_22107,N_22026);
xor U22578 (N_22578,N_22283,N_22321);
xnor U22579 (N_22579,N_22188,N_22336);
and U22580 (N_22580,N_22395,N_22124);
or U22581 (N_22581,N_22292,N_22152);
or U22582 (N_22582,N_21936,N_22498);
nor U22583 (N_22583,N_22437,N_22481);
nand U22584 (N_22584,N_22238,N_22351);
or U22585 (N_22585,N_22169,N_22111);
nor U22586 (N_22586,N_22436,N_22045);
nand U22587 (N_22587,N_22144,N_22285);
xnor U22588 (N_22588,N_21987,N_22478);
and U22589 (N_22589,N_22157,N_22325);
and U22590 (N_22590,N_22331,N_22064);
nand U22591 (N_22591,N_22272,N_22253);
nand U22592 (N_22592,N_22192,N_22471);
or U22593 (N_22593,N_22479,N_21877);
nor U22594 (N_22594,N_22091,N_21967);
nand U22595 (N_22595,N_22233,N_22203);
xor U22596 (N_22596,N_22109,N_22488);
nand U22597 (N_22597,N_21899,N_22313);
or U22598 (N_22598,N_22360,N_22252);
nor U22599 (N_22599,N_22089,N_22057);
nand U22600 (N_22600,N_22108,N_21947);
and U22601 (N_22601,N_22078,N_22394);
nand U22602 (N_22602,N_22355,N_22088);
nand U22603 (N_22603,N_22151,N_22446);
or U22604 (N_22604,N_21897,N_22412);
or U22605 (N_22605,N_22062,N_22156);
or U22606 (N_22606,N_22339,N_22223);
nand U22607 (N_22607,N_21972,N_22456);
nand U22608 (N_22608,N_22297,N_22345);
nor U22609 (N_22609,N_22342,N_21958);
and U22610 (N_22610,N_22464,N_22369);
nor U22611 (N_22611,N_22403,N_22421);
or U22612 (N_22612,N_22324,N_22365);
nor U22613 (N_22613,N_22126,N_22161);
and U22614 (N_22614,N_22312,N_22116);
or U22615 (N_22615,N_22074,N_22495);
and U22616 (N_22616,N_22445,N_22249);
nand U22617 (N_22617,N_21886,N_22061);
and U22618 (N_22618,N_22385,N_22167);
xor U22619 (N_22619,N_22362,N_21961);
or U22620 (N_22620,N_22150,N_22338);
and U22621 (N_22621,N_22115,N_21981);
and U22622 (N_22622,N_22459,N_21973);
and U22623 (N_22623,N_22042,N_22025);
nor U22624 (N_22624,N_21938,N_22486);
xor U22625 (N_22625,N_21984,N_22087);
nor U22626 (N_22626,N_22234,N_21889);
nor U22627 (N_22627,N_22417,N_22322);
nand U22628 (N_22628,N_22146,N_22487);
xnor U22629 (N_22629,N_22181,N_22386);
nor U22630 (N_22630,N_22049,N_21916);
or U22631 (N_22631,N_21969,N_21946);
and U22632 (N_22632,N_22413,N_22038);
xnor U22633 (N_22633,N_22199,N_22337);
and U22634 (N_22634,N_22485,N_21885);
and U22635 (N_22635,N_22069,N_21982);
and U22636 (N_22636,N_21979,N_22400);
nand U22637 (N_22637,N_22300,N_22258);
xnor U22638 (N_22638,N_22451,N_22017);
or U22639 (N_22639,N_22316,N_22317);
nor U22640 (N_22640,N_21966,N_22289);
xor U22641 (N_22641,N_22430,N_22344);
or U22642 (N_22642,N_22067,N_22326);
and U22643 (N_22643,N_22407,N_21925);
nand U22644 (N_22644,N_22117,N_22299);
and U22645 (N_22645,N_22346,N_22442);
or U22646 (N_22646,N_22180,N_21935);
nand U22647 (N_22647,N_22135,N_22140);
or U22648 (N_22648,N_22457,N_22263);
nor U22649 (N_22649,N_22315,N_22469);
and U22650 (N_22650,N_22226,N_22494);
xnor U22651 (N_22651,N_22414,N_22256);
nor U22652 (N_22652,N_22301,N_22189);
nand U22653 (N_22653,N_22318,N_22250);
and U22654 (N_22654,N_22173,N_22387);
xnor U22655 (N_22655,N_21923,N_22027);
or U22656 (N_22656,N_21893,N_22251);
xor U22657 (N_22657,N_22179,N_22406);
and U22658 (N_22658,N_22123,N_22068);
and U22659 (N_22659,N_22032,N_22051);
and U22660 (N_22660,N_22433,N_21881);
nor U22661 (N_22661,N_22177,N_22083);
nor U22662 (N_22662,N_22029,N_22132);
nor U22663 (N_22663,N_21934,N_22206);
nand U22664 (N_22664,N_22429,N_22327);
nor U22665 (N_22665,N_22071,N_22080);
xor U22666 (N_22666,N_21959,N_21953);
nor U22667 (N_22667,N_22121,N_22271);
nand U22668 (N_22668,N_22397,N_22110);
xnor U22669 (N_22669,N_22474,N_22440);
and U22670 (N_22670,N_22183,N_22257);
nand U22671 (N_22671,N_21939,N_22278);
nor U22672 (N_22672,N_22264,N_22019);
nor U22673 (N_22673,N_22174,N_22368);
nor U22674 (N_22674,N_22333,N_21907);
nand U22675 (N_22675,N_22033,N_22239);
or U22676 (N_22676,N_22454,N_22016);
and U22677 (N_22677,N_21955,N_22127);
and U22678 (N_22678,N_22476,N_22432);
nor U22679 (N_22679,N_22262,N_22021);
nand U22680 (N_22680,N_22043,N_22307);
or U22681 (N_22681,N_22425,N_22232);
nor U22682 (N_22682,N_22244,N_22261);
nand U22683 (N_22683,N_21974,N_22216);
and U22684 (N_22684,N_21976,N_22076);
and U22685 (N_22685,N_22492,N_22396);
xnor U22686 (N_22686,N_21882,N_22138);
or U22687 (N_22687,N_22482,N_22044);
nand U22688 (N_22688,N_22423,N_22200);
or U22689 (N_22689,N_22094,N_22090);
nand U22690 (N_22690,N_22393,N_22371);
xnor U22691 (N_22691,N_22490,N_22323);
or U22692 (N_22692,N_22245,N_22023);
and U22693 (N_22693,N_21917,N_22475);
and U22694 (N_22694,N_21910,N_22145);
nor U22695 (N_22695,N_21894,N_22309);
nor U22696 (N_22696,N_22081,N_22212);
or U22697 (N_22697,N_22160,N_22293);
nor U22698 (N_22698,N_22419,N_22066);
nor U22699 (N_22699,N_22217,N_21996);
nor U22700 (N_22700,N_22075,N_22237);
nor U22701 (N_22701,N_21920,N_22006);
nor U22702 (N_22702,N_22391,N_22073);
and U22703 (N_22703,N_22053,N_22473);
xor U22704 (N_22704,N_22480,N_22139);
nand U22705 (N_22705,N_22170,N_22184);
or U22706 (N_22706,N_21965,N_22491);
nor U22707 (N_22707,N_22470,N_22286);
nor U22708 (N_22708,N_21929,N_22439);
and U22709 (N_22709,N_22320,N_21933);
nand U22710 (N_22710,N_22047,N_22305);
xor U22711 (N_22711,N_21875,N_22329);
xnor U22712 (N_22712,N_21928,N_22375);
nand U22713 (N_22713,N_22266,N_22207);
and U22714 (N_22714,N_22428,N_22460);
or U22715 (N_22715,N_22493,N_22224);
and U22716 (N_22716,N_22399,N_22022);
and U22717 (N_22717,N_22211,N_22052);
or U22718 (N_22718,N_22028,N_22218);
xnor U22719 (N_22719,N_21942,N_22143);
nor U22720 (N_22720,N_22004,N_22210);
and U22721 (N_22721,N_21949,N_22340);
nor U22722 (N_22722,N_21915,N_21880);
xor U22723 (N_22723,N_22447,N_22030);
or U22724 (N_22724,N_22282,N_22229);
or U22725 (N_22725,N_22060,N_21963);
or U22726 (N_22726,N_21876,N_22159);
and U22727 (N_22727,N_21977,N_22378);
and U22728 (N_22728,N_22330,N_22194);
nand U22729 (N_22729,N_22267,N_22072);
nor U22730 (N_22730,N_21898,N_22221);
or U22731 (N_22731,N_22201,N_21903);
nor U22732 (N_22732,N_22185,N_22228);
nor U22733 (N_22733,N_22302,N_22450);
nand U22734 (N_22734,N_22095,N_22367);
nand U22735 (N_22735,N_22374,N_22050);
and U22736 (N_22736,N_22009,N_22082);
and U22737 (N_22737,N_21993,N_22392);
nor U22738 (N_22738,N_22426,N_22435);
and U22739 (N_22739,N_21887,N_22204);
nor U22740 (N_22740,N_21930,N_21940);
nor U22741 (N_22741,N_22040,N_22186);
xor U22742 (N_22742,N_22011,N_22213);
xor U22743 (N_22743,N_22389,N_22240);
and U22744 (N_22744,N_22401,N_22120);
or U22745 (N_22745,N_22270,N_21992);
nor U22746 (N_22746,N_22288,N_21999);
and U22747 (N_22747,N_22402,N_22219);
nor U22748 (N_22748,N_22438,N_21937);
nand U22749 (N_22749,N_22383,N_21957);
nand U22750 (N_22750,N_21994,N_22220);
or U22751 (N_22751,N_22357,N_22100);
nand U22752 (N_22752,N_22455,N_22003);
or U22753 (N_22753,N_22171,N_22372);
nand U22754 (N_22754,N_21944,N_22153);
nor U22755 (N_22755,N_21954,N_22453);
and U22756 (N_22756,N_22130,N_22255);
nor U22757 (N_22757,N_22225,N_22381);
and U22758 (N_22758,N_22311,N_22070);
or U22759 (N_22759,N_22273,N_22065);
xnor U22760 (N_22760,N_22163,N_21906);
nor U22761 (N_22761,N_22275,N_21995);
or U22762 (N_22762,N_22462,N_22390);
or U22763 (N_22763,N_22000,N_22416);
or U22764 (N_22764,N_22133,N_22363);
or U22765 (N_22765,N_22269,N_22164);
and U22766 (N_22766,N_22148,N_21960);
nor U22767 (N_22767,N_22298,N_22190);
nand U22768 (N_22768,N_22422,N_21892);
or U22769 (N_22769,N_21956,N_22008);
xnor U22770 (N_22770,N_22458,N_22198);
or U22771 (N_22771,N_21891,N_22279);
xnor U22772 (N_22772,N_22142,N_22187);
nand U22773 (N_22773,N_22248,N_22431);
or U22774 (N_22774,N_22005,N_22489);
nand U22775 (N_22775,N_22079,N_22352);
and U22776 (N_22776,N_21988,N_22424);
or U22777 (N_22777,N_22034,N_22077);
nor U22778 (N_22778,N_22149,N_22259);
or U22779 (N_22779,N_22379,N_22154);
and U22780 (N_22780,N_22227,N_22236);
or U22781 (N_22781,N_22472,N_22092);
or U22782 (N_22782,N_22193,N_22054);
nor U22783 (N_22783,N_22168,N_22247);
or U22784 (N_22784,N_22449,N_22284);
nand U22785 (N_22785,N_22162,N_21990);
nor U22786 (N_22786,N_22415,N_21991);
or U22787 (N_22787,N_22483,N_21971);
or U22788 (N_22788,N_21978,N_22484);
xor U22789 (N_22789,N_22497,N_22002);
and U22790 (N_22790,N_22125,N_22496);
nand U22791 (N_22791,N_22274,N_22443);
and U22792 (N_22792,N_22010,N_21918);
nand U22793 (N_22793,N_22059,N_22349);
nor U22794 (N_22794,N_21912,N_21980);
or U22795 (N_22795,N_22265,N_22448);
xor U22796 (N_22796,N_21970,N_22007);
xor U22797 (N_22797,N_21943,N_22434);
or U22798 (N_22798,N_22276,N_22129);
nor U22799 (N_22799,N_22452,N_22178);
and U22800 (N_22800,N_21879,N_22410);
nor U22801 (N_22801,N_21964,N_22461);
and U22802 (N_22802,N_22131,N_22020);
nand U22803 (N_22803,N_22377,N_22165);
nor U22804 (N_22804,N_22136,N_22197);
xnor U22805 (N_22805,N_22013,N_21989);
xor U22806 (N_22806,N_21983,N_22341);
xor U22807 (N_22807,N_22085,N_22246);
xor U22808 (N_22808,N_22319,N_22195);
or U22809 (N_22809,N_22101,N_22277);
nor U22810 (N_22810,N_21900,N_22202);
nor U22811 (N_22811,N_21902,N_21962);
nor U22812 (N_22812,N_22196,N_22206);
or U22813 (N_22813,N_22204,N_21935);
nor U22814 (N_22814,N_22062,N_22253);
and U22815 (N_22815,N_21966,N_22156);
nand U22816 (N_22816,N_21896,N_21951);
nor U22817 (N_22817,N_22082,N_22261);
or U22818 (N_22818,N_22326,N_22474);
nand U22819 (N_22819,N_22007,N_22239);
or U22820 (N_22820,N_22442,N_22141);
or U22821 (N_22821,N_21957,N_22144);
and U22822 (N_22822,N_22259,N_22032);
nor U22823 (N_22823,N_22452,N_22358);
xnor U22824 (N_22824,N_22017,N_22031);
nor U22825 (N_22825,N_22203,N_22433);
or U22826 (N_22826,N_22111,N_21966);
and U22827 (N_22827,N_21957,N_22195);
nor U22828 (N_22828,N_21902,N_22056);
nand U22829 (N_22829,N_22203,N_21954);
or U22830 (N_22830,N_22493,N_22495);
xnor U22831 (N_22831,N_22014,N_21982);
xor U22832 (N_22832,N_22302,N_22227);
nand U22833 (N_22833,N_21947,N_22437);
nand U22834 (N_22834,N_22212,N_22110);
nor U22835 (N_22835,N_22439,N_22294);
and U22836 (N_22836,N_21943,N_22416);
or U22837 (N_22837,N_22109,N_22310);
xnor U22838 (N_22838,N_22443,N_22091);
or U22839 (N_22839,N_21970,N_22267);
and U22840 (N_22840,N_22487,N_22019);
xor U22841 (N_22841,N_22496,N_22376);
nand U22842 (N_22842,N_22400,N_22371);
nor U22843 (N_22843,N_22024,N_22213);
nand U22844 (N_22844,N_22159,N_22426);
nand U22845 (N_22845,N_22305,N_22242);
or U22846 (N_22846,N_22280,N_22165);
nand U22847 (N_22847,N_22066,N_22435);
and U22848 (N_22848,N_22445,N_22462);
xnor U22849 (N_22849,N_21970,N_22200);
and U22850 (N_22850,N_22470,N_22288);
or U22851 (N_22851,N_22418,N_21938);
nor U22852 (N_22852,N_22459,N_21997);
nor U22853 (N_22853,N_22491,N_21914);
or U22854 (N_22854,N_22283,N_21893);
nor U22855 (N_22855,N_22441,N_22203);
xor U22856 (N_22856,N_22234,N_22150);
or U22857 (N_22857,N_22463,N_22197);
or U22858 (N_22858,N_22328,N_21882);
xor U22859 (N_22859,N_22256,N_22374);
nand U22860 (N_22860,N_22057,N_22488);
nor U22861 (N_22861,N_22175,N_22251);
xor U22862 (N_22862,N_21902,N_22217);
or U22863 (N_22863,N_22307,N_22217);
nand U22864 (N_22864,N_22420,N_22082);
xnor U22865 (N_22865,N_22201,N_22232);
xor U22866 (N_22866,N_21991,N_22463);
or U22867 (N_22867,N_22267,N_21898);
nor U22868 (N_22868,N_22147,N_21959);
or U22869 (N_22869,N_21954,N_21932);
xnor U22870 (N_22870,N_22163,N_22178);
and U22871 (N_22871,N_22254,N_21991);
or U22872 (N_22872,N_22092,N_21922);
xnor U22873 (N_22873,N_21938,N_21999);
nand U22874 (N_22874,N_22319,N_22235);
xor U22875 (N_22875,N_22498,N_22199);
nand U22876 (N_22876,N_22123,N_22415);
and U22877 (N_22877,N_22123,N_22095);
nand U22878 (N_22878,N_21946,N_22197);
xnor U22879 (N_22879,N_21968,N_22439);
xor U22880 (N_22880,N_22449,N_22293);
and U22881 (N_22881,N_22003,N_22474);
and U22882 (N_22882,N_22221,N_22335);
xor U22883 (N_22883,N_22491,N_22094);
nand U22884 (N_22884,N_22151,N_22319);
xor U22885 (N_22885,N_22415,N_22061);
xor U22886 (N_22886,N_22307,N_22144);
or U22887 (N_22887,N_21969,N_21877);
nand U22888 (N_22888,N_22314,N_22262);
nand U22889 (N_22889,N_22059,N_21901);
nor U22890 (N_22890,N_22351,N_22305);
or U22891 (N_22891,N_22408,N_22382);
nor U22892 (N_22892,N_22303,N_21984);
nand U22893 (N_22893,N_22219,N_22378);
xnor U22894 (N_22894,N_22055,N_22101);
xor U22895 (N_22895,N_22172,N_21906);
and U22896 (N_22896,N_22464,N_22333);
nand U22897 (N_22897,N_22113,N_22122);
nor U22898 (N_22898,N_22487,N_22379);
nor U22899 (N_22899,N_22242,N_21950);
nand U22900 (N_22900,N_22373,N_22202);
nor U22901 (N_22901,N_22133,N_22006);
xor U22902 (N_22902,N_21986,N_22249);
and U22903 (N_22903,N_21918,N_21885);
nand U22904 (N_22904,N_21930,N_22330);
and U22905 (N_22905,N_22276,N_22450);
and U22906 (N_22906,N_22390,N_22072);
nor U22907 (N_22907,N_22304,N_22239);
and U22908 (N_22908,N_22351,N_22031);
and U22909 (N_22909,N_22200,N_22242);
nor U22910 (N_22910,N_22453,N_22089);
nand U22911 (N_22911,N_22439,N_22028);
and U22912 (N_22912,N_22017,N_21879);
and U22913 (N_22913,N_22014,N_22167);
nor U22914 (N_22914,N_22489,N_22206);
nand U22915 (N_22915,N_22006,N_22327);
nor U22916 (N_22916,N_22239,N_22079);
xnor U22917 (N_22917,N_22153,N_22076);
and U22918 (N_22918,N_21968,N_22487);
or U22919 (N_22919,N_22023,N_22486);
or U22920 (N_22920,N_22390,N_22475);
nand U22921 (N_22921,N_22410,N_22394);
xnor U22922 (N_22922,N_22468,N_21888);
or U22923 (N_22923,N_21909,N_22259);
xnor U22924 (N_22924,N_22253,N_22433);
or U22925 (N_22925,N_21967,N_22218);
xnor U22926 (N_22926,N_22126,N_22343);
or U22927 (N_22927,N_22260,N_22087);
or U22928 (N_22928,N_22122,N_22146);
nor U22929 (N_22929,N_22475,N_22019);
or U22930 (N_22930,N_22179,N_22024);
xnor U22931 (N_22931,N_22335,N_22352);
and U22932 (N_22932,N_22361,N_22129);
xor U22933 (N_22933,N_22196,N_22165);
and U22934 (N_22934,N_22428,N_22419);
nand U22935 (N_22935,N_22495,N_22171);
nor U22936 (N_22936,N_21914,N_21964);
nor U22937 (N_22937,N_21974,N_22189);
or U22938 (N_22938,N_22437,N_22033);
or U22939 (N_22939,N_22427,N_21937);
and U22940 (N_22940,N_22258,N_21900);
and U22941 (N_22941,N_21984,N_21934);
or U22942 (N_22942,N_22227,N_22073);
and U22943 (N_22943,N_22175,N_22102);
or U22944 (N_22944,N_22055,N_22126);
nor U22945 (N_22945,N_22026,N_21909);
nor U22946 (N_22946,N_22471,N_22171);
nand U22947 (N_22947,N_22193,N_21975);
nand U22948 (N_22948,N_21926,N_22458);
xnor U22949 (N_22949,N_22356,N_22106);
nor U22950 (N_22950,N_22269,N_22143);
and U22951 (N_22951,N_22428,N_22473);
and U22952 (N_22952,N_22333,N_22151);
and U22953 (N_22953,N_22049,N_21973);
nor U22954 (N_22954,N_22208,N_22079);
xnor U22955 (N_22955,N_22173,N_21935);
xnor U22956 (N_22956,N_21904,N_22339);
or U22957 (N_22957,N_22425,N_22302);
or U22958 (N_22958,N_21981,N_22190);
or U22959 (N_22959,N_22092,N_22222);
nor U22960 (N_22960,N_22062,N_22409);
nand U22961 (N_22961,N_22384,N_22060);
and U22962 (N_22962,N_21998,N_21926);
or U22963 (N_22963,N_22437,N_22146);
or U22964 (N_22964,N_22481,N_22362);
nand U22965 (N_22965,N_22466,N_22250);
or U22966 (N_22966,N_22250,N_22388);
xnor U22967 (N_22967,N_22233,N_22104);
xnor U22968 (N_22968,N_22499,N_22263);
xnor U22969 (N_22969,N_22373,N_22166);
nor U22970 (N_22970,N_21906,N_22022);
nor U22971 (N_22971,N_22228,N_22029);
and U22972 (N_22972,N_22491,N_22047);
and U22973 (N_22973,N_22402,N_22042);
xor U22974 (N_22974,N_22206,N_22365);
xor U22975 (N_22975,N_22454,N_22072);
nor U22976 (N_22976,N_21980,N_22209);
nand U22977 (N_22977,N_21912,N_22475);
nor U22978 (N_22978,N_22309,N_22117);
or U22979 (N_22979,N_22436,N_21999);
xor U22980 (N_22980,N_22195,N_22388);
xnor U22981 (N_22981,N_22364,N_22174);
nand U22982 (N_22982,N_21969,N_22193);
or U22983 (N_22983,N_21934,N_22124);
xnor U22984 (N_22984,N_22289,N_22189);
xnor U22985 (N_22985,N_22251,N_21922);
nand U22986 (N_22986,N_22379,N_22228);
nor U22987 (N_22987,N_21936,N_22303);
and U22988 (N_22988,N_22455,N_22316);
nand U22989 (N_22989,N_21900,N_22120);
or U22990 (N_22990,N_22221,N_22180);
nand U22991 (N_22991,N_22046,N_22336);
and U22992 (N_22992,N_21880,N_22014);
xor U22993 (N_22993,N_22356,N_21911);
nor U22994 (N_22994,N_22250,N_22024);
xnor U22995 (N_22995,N_22105,N_21964);
xnor U22996 (N_22996,N_22105,N_22280);
and U22997 (N_22997,N_22238,N_22377);
and U22998 (N_22998,N_22196,N_22162);
or U22999 (N_22999,N_22479,N_22496);
and U23000 (N_23000,N_22173,N_21898);
nor U23001 (N_23001,N_22360,N_22090);
and U23002 (N_23002,N_22057,N_22144);
nand U23003 (N_23003,N_22444,N_22104);
xnor U23004 (N_23004,N_22084,N_22203);
xnor U23005 (N_23005,N_22188,N_22217);
or U23006 (N_23006,N_21947,N_22164);
and U23007 (N_23007,N_22357,N_22053);
nor U23008 (N_23008,N_22020,N_22065);
and U23009 (N_23009,N_22484,N_22208);
and U23010 (N_23010,N_22288,N_22307);
and U23011 (N_23011,N_22202,N_22259);
xnor U23012 (N_23012,N_22035,N_22303);
nand U23013 (N_23013,N_22141,N_22322);
and U23014 (N_23014,N_22184,N_22398);
nand U23015 (N_23015,N_22270,N_22222);
nor U23016 (N_23016,N_21991,N_22395);
nand U23017 (N_23017,N_22365,N_22088);
nor U23018 (N_23018,N_21911,N_21998);
and U23019 (N_23019,N_22485,N_22342);
nand U23020 (N_23020,N_22277,N_22302);
nand U23021 (N_23021,N_22480,N_22006);
or U23022 (N_23022,N_22067,N_22064);
nand U23023 (N_23023,N_22463,N_22220);
and U23024 (N_23024,N_22170,N_21891);
nand U23025 (N_23025,N_22494,N_22075);
and U23026 (N_23026,N_21927,N_22473);
xnor U23027 (N_23027,N_22131,N_22350);
xor U23028 (N_23028,N_22489,N_22313);
nand U23029 (N_23029,N_21923,N_21937);
xnor U23030 (N_23030,N_22460,N_22107);
xor U23031 (N_23031,N_22321,N_22197);
xnor U23032 (N_23032,N_21894,N_22403);
xnor U23033 (N_23033,N_22150,N_22480);
nor U23034 (N_23034,N_21982,N_21985);
nand U23035 (N_23035,N_21931,N_22306);
nor U23036 (N_23036,N_22288,N_21965);
nor U23037 (N_23037,N_22250,N_22246);
nor U23038 (N_23038,N_22214,N_22138);
or U23039 (N_23039,N_22161,N_21888);
and U23040 (N_23040,N_21985,N_21963);
xor U23041 (N_23041,N_21966,N_21915);
and U23042 (N_23042,N_22381,N_22112);
nor U23043 (N_23043,N_22299,N_21901);
or U23044 (N_23044,N_22115,N_22337);
xor U23045 (N_23045,N_22179,N_22061);
nor U23046 (N_23046,N_22118,N_22476);
nand U23047 (N_23047,N_21915,N_22115);
or U23048 (N_23048,N_22313,N_22317);
or U23049 (N_23049,N_22166,N_22366);
and U23050 (N_23050,N_22411,N_22336);
or U23051 (N_23051,N_22383,N_21953);
xor U23052 (N_23052,N_22315,N_22160);
nand U23053 (N_23053,N_22178,N_22004);
nand U23054 (N_23054,N_22480,N_22351);
nand U23055 (N_23055,N_22455,N_21904);
xnor U23056 (N_23056,N_22374,N_22388);
nor U23057 (N_23057,N_21981,N_22205);
nor U23058 (N_23058,N_22173,N_22137);
and U23059 (N_23059,N_22318,N_22089);
and U23060 (N_23060,N_22447,N_22243);
nor U23061 (N_23061,N_22432,N_21902);
nor U23062 (N_23062,N_22452,N_22107);
or U23063 (N_23063,N_22488,N_22432);
xnor U23064 (N_23064,N_22088,N_21962);
nand U23065 (N_23065,N_22334,N_21903);
nor U23066 (N_23066,N_22208,N_22052);
or U23067 (N_23067,N_22301,N_22248);
nand U23068 (N_23068,N_21895,N_22130);
or U23069 (N_23069,N_22250,N_22363);
xor U23070 (N_23070,N_22448,N_22182);
and U23071 (N_23071,N_22225,N_22159);
nand U23072 (N_23072,N_21981,N_21919);
nor U23073 (N_23073,N_22041,N_22141);
xnor U23074 (N_23074,N_22163,N_22468);
nor U23075 (N_23075,N_21929,N_22097);
xnor U23076 (N_23076,N_22074,N_21983);
and U23077 (N_23077,N_22344,N_22450);
nor U23078 (N_23078,N_22184,N_22201);
or U23079 (N_23079,N_21949,N_21988);
and U23080 (N_23080,N_22322,N_22242);
and U23081 (N_23081,N_22289,N_21887);
nor U23082 (N_23082,N_22280,N_21880);
and U23083 (N_23083,N_22340,N_21879);
and U23084 (N_23084,N_22411,N_22488);
xnor U23085 (N_23085,N_22012,N_22346);
xor U23086 (N_23086,N_22037,N_22341);
xor U23087 (N_23087,N_22202,N_22437);
nor U23088 (N_23088,N_22204,N_22142);
nand U23089 (N_23089,N_22277,N_22353);
nor U23090 (N_23090,N_22358,N_22228);
nand U23091 (N_23091,N_22447,N_21965);
xnor U23092 (N_23092,N_22052,N_22284);
or U23093 (N_23093,N_22195,N_22472);
nand U23094 (N_23094,N_22016,N_22132);
nand U23095 (N_23095,N_22188,N_21877);
nand U23096 (N_23096,N_22447,N_21913);
nor U23097 (N_23097,N_22242,N_22389);
xnor U23098 (N_23098,N_22498,N_22315);
nor U23099 (N_23099,N_22029,N_22222);
or U23100 (N_23100,N_21907,N_22317);
nand U23101 (N_23101,N_22492,N_22465);
and U23102 (N_23102,N_22454,N_21903);
xnor U23103 (N_23103,N_22022,N_22326);
xor U23104 (N_23104,N_22076,N_22408);
and U23105 (N_23105,N_22386,N_22463);
nor U23106 (N_23106,N_22334,N_22498);
xor U23107 (N_23107,N_22344,N_22425);
nand U23108 (N_23108,N_22322,N_22168);
and U23109 (N_23109,N_21964,N_22486);
xnor U23110 (N_23110,N_22061,N_22285);
or U23111 (N_23111,N_22199,N_22344);
nor U23112 (N_23112,N_22133,N_22369);
or U23113 (N_23113,N_22089,N_21939);
or U23114 (N_23114,N_22196,N_22145);
or U23115 (N_23115,N_22076,N_22407);
or U23116 (N_23116,N_21969,N_22037);
nand U23117 (N_23117,N_21988,N_22168);
nand U23118 (N_23118,N_22068,N_21969);
xor U23119 (N_23119,N_21898,N_22408);
nand U23120 (N_23120,N_22267,N_21919);
nand U23121 (N_23121,N_22466,N_22484);
xnor U23122 (N_23122,N_22258,N_22195);
or U23123 (N_23123,N_21962,N_22192);
or U23124 (N_23124,N_22131,N_22416);
xnor U23125 (N_23125,N_23032,N_22815);
and U23126 (N_23126,N_22615,N_22842);
xnor U23127 (N_23127,N_22625,N_22580);
nor U23128 (N_23128,N_22880,N_22841);
or U23129 (N_23129,N_22720,N_22688);
and U23130 (N_23130,N_22549,N_22639);
xnor U23131 (N_23131,N_23062,N_23080);
and U23132 (N_23132,N_23071,N_22777);
nor U23133 (N_23133,N_22729,N_22871);
nand U23134 (N_23134,N_22678,N_23037);
and U23135 (N_23135,N_22622,N_22530);
nand U23136 (N_23136,N_22614,N_22783);
or U23137 (N_23137,N_22870,N_22578);
nor U23138 (N_23138,N_22938,N_22764);
and U23139 (N_23139,N_22686,N_22765);
or U23140 (N_23140,N_23029,N_23002);
nor U23141 (N_23141,N_22893,N_22752);
nor U23142 (N_23142,N_22927,N_22597);
xor U23143 (N_23143,N_22721,N_23003);
xor U23144 (N_23144,N_23072,N_22994);
nor U23145 (N_23145,N_22664,N_22659);
or U23146 (N_23146,N_23038,N_22576);
or U23147 (N_23147,N_23118,N_22836);
and U23148 (N_23148,N_22600,N_22537);
and U23149 (N_23149,N_22540,N_23091);
nand U23150 (N_23150,N_22991,N_22918);
nor U23151 (N_23151,N_22932,N_23011);
or U23152 (N_23152,N_22901,N_22692);
or U23153 (N_23153,N_22786,N_22564);
and U23154 (N_23154,N_22903,N_22575);
nor U23155 (N_23155,N_22737,N_22892);
nor U23156 (N_23156,N_22953,N_22518);
and U23157 (N_23157,N_23027,N_22684);
xor U23158 (N_23158,N_22663,N_22621);
xnor U23159 (N_23159,N_23036,N_22562);
xnor U23160 (N_23160,N_22669,N_22833);
nand U23161 (N_23161,N_22898,N_22539);
nand U23162 (N_23162,N_22652,N_23121);
nor U23163 (N_23163,N_22662,N_22941);
nor U23164 (N_23164,N_23065,N_22679);
nand U23165 (N_23165,N_22793,N_22822);
nor U23166 (N_23166,N_22887,N_22873);
nand U23167 (N_23167,N_23031,N_23087);
or U23168 (N_23168,N_23108,N_22508);
nor U23169 (N_23169,N_22795,N_23025);
and U23170 (N_23170,N_22753,N_22657);
or U23171 (N_23171,N_23058,N_22587);
or U23172 (N_23172,N_22974,N_22972);
and U23173 (N_23173,N_23056,N_22637);
nand U23174 (N_23174,N_23006,N_22816);
nand U23175 (N_23175,N_22904,N_22541);
and U23176 (N_23176,N_23124,N_22650);
and U23177 (N_23177,N_22709,N_22520);
or U23178 (N_23178,N_23020,N_22512);
nor U23179 (N_23179,N_22961,N_22609);
or U23180 (N_23180,N_23061,N_23059);
and U23181 (N_23181,N_22642,N_23088);
xnor U23182 (N_23182,N_22837,N_22784);
xor U23183 (N_23183,N_23077,N_22946);
and U23184 (N_23184,N_22633,N_22981);
nor U23185 (N_23185,N_23090,N_22750);
or U23186 (N_23186,N_22949,N_22733);
xnor U23187 (N_23187,N_23084,N_22919);
nand U23188 (N_23188,N_22547,N_23107);
or U23189 (N_23189,N_22533,N_22846);
nor U23190 (N_23190,N_22661,N_22695);
xnor U23191 (N_23191,N_22568,N_22844);
nor U23192 (N_23192,N_22862,N_23008);
nand U23193 (N_23193,N_22566,N_22649);
nor U23194 (N_23194,N_22970,N_23075);
and U23195 (N_23195,N_22761,N_22601);
and U23196 (N_23196,N_22589,N_22990);
xor U23197 (N_23197,N_22704,N_22591);
nand U23198 (N_23198,N_22999,N_22996);
nand U23199 (N_23199,N_22735,N_22643);
and U23200 (N_23200,N_22856,N_22671);
or U23201 (N_23201,N_22628,N_22725);
nor U23202 (N_23202,N_23070,N_22624);
or U23203 (N_23203,N_22567,N_22526);
and U23204 (N_23204,N_22888,N_22611);
nor U23205 (N_23205,N_22824,N_22993);
nor U23206 (N_23206,N_22574,N_22909);
xor U23207 (N_23207,N_23044,N_22976);
nand U23208 (N_23208,N_23082,N_22937);
nand U23209 (N_23209,N_22668,N_22950);
nor U23210 (N_23210,N_22654,N_22978);
nand U23211 (N_23211,N_22785,N_22971);
nand U23212 (N_23212,N_23099,N_22523);
nand U23213 (N_23213,N_22807,N_22636);
nand U23214 (N_23214,N_22641,N_22998);
nand U23215 (N_23215,N_22944,N_22595);
and U23216 (N_23216,N_22581,N_22845);
or U23217 (N_23217,N_22930,N_22811);
or U23218 (N_23218,N_22703,N_22516);
nor U23219 (N_23219,N_22556,N_22675);
xnor U23220 (N_23220,N_22719,N_22958);
xnor U23221 (N_23221,N_22832,N_22532);
xnor U23222 (N_23222,N_22812,N_22963);
nand U23223 (N_23223,N_22813,N_22739);
or U23224 (N_23224,N_23116,N_23010);
or U23225 (N_23225,N_22718,N_22790);
or U23226 (N_23226,N_22690,N_22890);
or U23227 (N_23227,N_23110,N_22724);
nor U23228 (N_23228,N_22706,N_22859);
or U23229 (N_23229,N_23093,N_22986);
or U23230 (N_23230,N_23081,N_23086);
nor U23231 (N_23231,N_22948,N_22912);
xnor U23232 (N_23232,N_22602,N_22634);
or U23233 (N_23233,N_22527,N_22623);
xnor U23234 (N_23234,N_23076,N_22559);
xor U23235 (N_23235,N_22814,N_22683);
xor U23236 (N_23236,N_22774,N_23114);
nand U23237 (N_23237,N_23046,N_22939);
or U23238 (N_23238,N_22665,N_23120);
or U23239 (N_23239,N_23095,N_23078);
nor U23240 (N_23240,N_22504,N_22913);
xor U23241 (N_23241,N_22980,N_22908);
or U23242 (N_23242,N_22584,N_22770);
or U23243 (N_23243,N_22917,N_22571);
or U23244 (N_23244,N_22962,N_22630);
nor U23245 (N_23245,N_23034,N_22693);
or U23246 (N_23246,N_22985,N_22676);
nand U23247 (N_23247,N_23101,N_22509);
nand U23248 (N_23248,N_22947,N_22742);
or U23249 (N_23249,N_22900,N_22960);
and U23250 (N_23250,N_22943,N_22557);
nor U23251 (N_23251,N_23019,N_23069);
nand U23252 (N_23252,N_22585,N_22992);
or U23253 (N_23253,N_22705,N_22872);
or U23254 (N_23254,N_22808,N_22572);
nand U23255 (N_23255,N_23000,N_22744);
and U23256 (N_23256,N_23100,N_22826);
and U23257 (N_23257,N_22715,N_22945);
and U23258 (N_23258,N_22843,N_22910);
nand U23259 (N_23259,N_22681,N_22866);
nor U23260 (N_23260,N_22687,N_22989);
or U23261 (N_23261,N_22685,N_22726);
and U23262 (N_23262,N_22928,N_22613);
nand U23263 (N_23263,N_22874,N_22513);
nor U23264 (N_23264,N_22529,N_22987);
and U23265 (N_23265,N_22698,N_22926);
or U23266 (N_23266,N_22902,N_22922);
nor U23267 (N_23267,N_22797,N_22593);
xor U23268 (N_23268,N_23035,N_22689);
nor U23269 (N_23269,N_22925,N_22629);
nor U23270 (N_23270,N_22984,N_22732);
nand U23271 (N_23271,N_22653,N_22966);
xnor U23272 (N_23272,N_22916,N_22579);
and U23273 (N_23273,N_22590,N_22635);
and U23274 (N_23274,N_22594,N_23063);
or U23275 (N_23275,N_22514,N_22755);
and U23276 (N_23276,N_23096,N_22697);
nand U23277 (N_23277,N_22760,N_22616);
nor U23278 (N_23278,N_22552,N_22858);
nand U23279 (N_23279,N_23045,N_22792);
or U23280 (N_23280,N_22857,N_23068);
nor U23281 (N_23281,N_22640,N_23030);
or U23282 (N_23282,N_23040,N_23094);
xnor U23283 (N_23283,N_22804,N_23103);
nor U23284 (N_23284,N_22831,N_22535);
nor U23285 (N_23285,N_22769,N_22775);
nor U23286 (N_23286,N_22895,N_22670);
xnor U23287 (N_23287,N_23119,N_22731);
or U23288 (N_23288,N_23054,N_22906);
or U23289 (N_23289,N_22881,N_22632);
or U23290 (N_23290,N_22700,N_22800);
and U23291 (N_23291,N_22710,N_22531);
and U23292 (N_23292,N_22538,N_22544);
nor U23293 (N_23293,N_22924,N_22608);
nand U23294 (N_23294,N_22779,N_23113);
nand U23295 (N_23295,N_22696,N_22524);
and U23296 (N_23296,N_22738,N_22713);
xnor U23297 (N_23297,N_22796,N_22542);
nor U23298 (N_23298,N_22507,N_22711);
nand U23299 (N_23299,N_22536,N_22596);
nand U23300 (N_23300,N_23079,N_22519);
or U23301 (N_23301,N_23013,N_22701);
or U23302 (N_23302,N_22799,N_22849);
nor U23303 (N_23303,N_22631,N_22734);
nand U23304 (N_23304,N_22933,N_22864);
nand U23305 (N_23305,N_23073,N_22951);
xnor U23306 (N_23306,N_22560,N_23064);
xor U23307 (N_23307,N_22680,N_22782);
and U23308 (N_23308,N_22860,N_22565);
and U23309 (N_23309,N_22920,N_22603);
or U23310 (N_23310,N_23052,N_22869);
nand U23311 (N_23311,N_22772,N_22847);
xor U23312 (N_23312,N_22911,N_22914);
and U23313 (N_23313,N_22714,N_22707);
and U23314 (N_23314,N_23060,N_22598);
nand U23315 (N_23315,N_22778,N_23066);
or U23316 (N_23316,N_22666,N_22510);
and U23317 (N_23317,N_22759,N_22551);
nand U23318 (N_23318,N_22867,N_22754);
or U23319 (N_23319,N_23028,N_22505);
nand U23320 (N_23320,N_22868,N_23053);
nor U23321 (N_23321,N_23115,N_22656);
and U23322 (N_23322,N_22776,N_22968);
nand U23323 (N_23323,N_23024,N_22626);
and U23324 (N_23324,N_22682,N_22702);
or U23325 (N_23325,N_22672,N_23111);
nor U23326 (N_23326,N_22522,N_22854);
nand U23327 (N_23327,N_22889,N_22757);
nor U23328 (N_23328,N_23042,N_22882);
and U23329 (N_23329,N_22569,N_22740);
xor U23330 (N_23330,N_23039,N_22967);
and U23331 (N_23331,N_22583,N_22691);
or U23332 (N_23332,N_23051,N_22570);
or U23333 (N_23333,N_23050,N_22545);
nand U23334 (N_23334,N_22699,N_22787);
xnor U23335 (N_23335,N_22879,N_22521);
xnor U23336 (N_23336,N_22929,N_22528);
nor U23337 (N_23337,N_22931,N_22977);
xor U23338 (N_23338,N_22801,N_22762);
and U23339 (N_23339,N_23043,N_23112);
xnor U23340 (N_23340,N_22975,N_22878);
nor U23341 (N_23341,N_23097,N_23067);
or U23342 (N_23342,N_22751,N_22500);
nor U23343 (N_23343,N_23022,N_22604);
nand U23344 (N_23344,N_23004,N_22658);
xnor U23345 (N_23345,N_22850,N_22788);
xor U23346 (N_23346,N_22756,N_22964);
nand U23347 (N_23347,N_23009,N_23041);
and U23348 (N_23348,N_22502,N_22618);
or U23349 (N_23349,N_22674,N_22781);
or U23350 (N_23350,N_23085,N_23109);
xnor U23351 (N_23351,N_22934,N_23055);
or U23352 (N_23352,N_22546,N_23098);
nand U23353 (N_23353,N_22840,N_22543);
and U23354 (N_23354,N_22561,N_22852);
and U23355 (N_23355,N_22853,N_22525);
xor U23356 (N_23356,N_23001,N_22766);
nor U23357 (N_23357,N_22716,N_23117);
or U23358 (N_23358,N_23033,N_23016);
or U23359 (N_23359,N_23105,N_22988);
and U23360 (N_23360,N_22883,N_22952);
or U23361 (N_23361,N_22517,N_22673);
or U23362 (N_23362,N_23092,N_22956);
and U23363 (N_23363,N_22942,N_22550);
xor U23364 (N_23364,N_22548,N_22646);
xnor U23365 (N_23365,N_22651,N_22749);
nand U23366 (N_23366,N_22727,N_22767);
and U23367 (N_23367,N_22973,N_22875);
xnor U23368 (N_23368,N_22921,N_22899);
or U23369 (N_23369,N_23057,N_22667);
nand U23370 (N_23370,N_22955,N_22896);
xor U23371 (N_23371,N_22728,N_22555);
and U23372 (N_23372,N_23047,N_22708);
xor U23373 (N_23373,N_22823,N_22897);
or U23374 (N_23374,N_22617,N_22592);
nand U23375 (N_23375,N_22503,N_22791);
nand U23376 (N_23376,N_22820,N_22794);
and U23377 (N_23377,N_22954,N_22923);
and U23378 (N_23378,N_22554,N_22768);
nor U23379 (N_23379,N_22627,N_23049);
or U23380 (N_23380,N_22619,N_22979);
nand U23381 (N_23381,N_22825,N_22717);
or U23382 (N_23382,N_22805,N_22838);
or U23383 (N_23383,N_22798,N_22694);
xor U23384 (N_23384,N_22803,N_22736);
nand U23385 (N_23385,N_22810,N_23106);
xnor U23386 (N_23386,N_22773,N_22915);
nor U23387 (N_23387,N_23026,N_22957);
and U23388 (N_23388,N_22599,N_22819);
and U23389 (N_23389,N_23048,N_22730);
xor U23390 (N_23390,N_22817,N_22620);
nor U23391 (N_23391,N_22834,N_22648);
and U23392 (N_23392,N_23018,N_23015);
xnor U23393 (N_23393,N_22863,N_22758);
and U23394 (N_23394,N_22563,N_22606);
nand U23395 (N_23395,N_22607,N_22884);
xor U23396 (N_23396,N_23017,N_22515);
nor U23397 (N_23397,N_22969,N_22936);
and U23398 (N_23398,N_22997,N_22645);
nand U23399 (N_23399,N_22582,N_22982);
and U23400 (N_23400,N_22983,N_22588);
nand U23401 (N_23401,N_22746,N_22780);
and U23402 (N_23402,N_22723,N_22806);
and U23403 (N_23403,N_22763,N_22677);
or U23404 (N_23404,N_22861,N_22818);
and U23405 (N_23405,N_22743,N_22586);
xor U23406 (N_23406,N_22835,N_22828);
xor U23407 (N_23407,N_22506,N_22747);
nand U23408 (N_23408,N_22647,N_22741);
or U23409 (N_23409,N_22855,N_22851);
or U23410 (N_23410,N_22748,N_22907);
or U23411 (N_23411,N_23123,N_22534);
and U23412 (N_23412,N_23074,N_22809);
and U23413 (N_23413,N_23021,N_22558);
nor U23414 (N_23414,N_22940,N_22995);
and U23415 (N_23415,N_22771,N_23005);
nand U23416 (N_23416,N_22829,N_22830);
and U23417 (N_23417,N_22802,N_22638);
or U23418 (N_23418,N_22511,N_22821);
nor U23419 (N_23419,N_22935,N_22894);
and U23420 (N_23420,N_23083,N_23089);
nand U23421 (N_23421,N_22553,N_22839);
nor U23422 (N_23422,N_23007,N_23122);
nand U23423 (N_23423,N_22905,N_22745);
and U23424 (N_23424,N_22885,N_22573);
and U23425 (N_23425,N_22655,N_22891);
nor U23426 (N_23426,N_23104,N_23102);
or U23427 (N_23427,N_22660,N_22789);
and U23428 (N_23428,N_22877,N_22965);
nand U23429 (N_23429,N_22712,N_23014);
and U23430 (N_23430,N_23012,N_22722);
nand U23431 (N_23431,N_22605,N_22848);
nor U23432 (N_23432,N_22644,N_22876);
or U23433 (N_23433,N_22827,N_22577);
and U23434 (N_23434,N_22610,N_22612);
xor U23435 (N_23435,N_22501,N_22865);
nor U23436 (N_23436,N_23023,N_22959);
nor U23437 (N_23437,N_22886,N_22961);
xor U23438 (N_23438,N_22796,N_22566);
nor U23439 (N_23439,N_22731,N_22593);
and U23440 (N_23440,N_22566,N_22910);
xor U23441 (N_23441,N_22813,N_22765);
nand U23442 (N_23442,N_22569,N_22820);
nor U23443 (N_23443,N_22831,N_22792);
and U23444 (N_23444,N_23018,N_22686);
nor U23445 (N_23445,N_22694,N_22826);
nand U23446 (N_23446,N_22737,N_22713);
nor U23447 (N_23447,N_22577,N_23034);
xor U23448 (N_23448,N_22775,N_22710);
or U23449 (N_23449,N_23092,N_23063);
nor U23450 (N_23450,N_22909,N_22856);
nand U23451 (N_23451,N_22618,N_23124);
and U23452 (N_23452,N_22558,N_22713);
nand U23453 (N_23453,N_22690,N_22790);
and U23454 (N_23454,N_23068,N_22665);
nor U23455 (N_23455,N_22708,N_22957);
or U23456 (N_23456,N_22555,N_22928);
and U23457 (N_23457,N_22943,N_22946);
nand U23458 (N_23458,N_22797,N_23060);
nand U23459 (N_23459,N_22593,N_22843);
or U23460 (N_23460,N_22517,N_22748);
xnor U23461 (N_23461,N_22621,N_22713);
xor U23462 (N_23462,N_22684,N_22953);
nand U23463 (N_23463,N_23025,N_22787);
nor U23464 (N_23464,N_22927,N_23013);
or U23465 (N_23465,N_22932,N_23112);
xnor U23466 (N_23466,N_22756,N_23089);
and U23467 (N_23467,N_22686,N_22788);
nor U23468 (N_23468,N_23068,N_22634);
and U23469 (N_23469,N_22814,N_22873);
nor U23470 (N_23470,N_22683,N_22893);
nand U23471 (N_23471,N_23096,N_22790);
and U23472 (N_23472,N_23053,N_22756);
or U23473 (N_23473,N_22800,N_22707);
and U23474 (N_23474,N_22547,N_22958);
and U23475 (N_23475,N_22662,N_22587);
and U23476 (N_23476,N_22878,N_22504);
or U23477 (N_23477,N_22807,N_22515);
nand U23478 (N_23478,N_22616,N_22504);
xor U23479 (N_23479,N_22677,N_22825);
nand U23480 (N_23480,N_23037,N_22935);
xnor U23481 (N_23481,N_22610,N_22578);
nor U23482 (N_23482,N_22541,N_22556);
nor U23483 (N_23483,N_22595,N_22557);
nor U23484 (N_23484,N_22851,N_22742);
xnor U23485 (N_23485,N_22636,N_22801);
or U23486 (N_23486,N_22672,N_23003);
xor U23487 (N_23487,N_22941,N_23051);
nand U23488 (N_23488,N_23097,N_22608);
xor U23489 (N_23489,N_22882,N_22892);
xor U23490 (N_23490,N_22680,N_23031);
nand U23491 (N_23491,N_22699,N_22931);
or U23492 (N_23492,N_23053,N_22736);
nor U23493 (N_23493,N_22563,N_22927);
xor U23494 (N_23494,N_22559,N_22663);
or U23495 (N_23495,N_23084,N_22928);
nor U23496 (N_23496,N_22519,N_22819);
and U23497 (N_23497,N_22751,N_22880);
and U23498 (N_23498,N_22883,N_22827);
and U23499 (N_23499,N_23031,N_22910);
or U23500 (N_23500,N_22538,N_22634);
and U23501 (N_23501,N_22986,N_22868);
nand U23502 (N_23502,N_22813,N_23099);
xor U23503 (N_23503,N_22706,N_22576);
xor U23504 (N_23504,N_22966,N_22550);
and U23505 (N_23505,N_22683,N_22509);
and U23506 (N_23506,N_23067,N_22502);
xor U23507 (N_23507,N_22744,N_23046);
xnor U23508 (N_23508,N_22517,N_22852);
and U23509 (N_23509,N_22507,N_22640);
nor U23510 (N_23510,N_23071,N_23105);
nand U23511 (N_23511,N_22558,N_22730);
and U23512 (N_23512,N_22861,N_22738);
xnor U23513 (N_23513,N_22994,N_23020);
and U23514 (N_23514,N_23092,N_22797);
and U23515 (N_23515,N_22680,N_23119);
xnor U23516 (N_23516,N_22902,N_22568);
xor U23517 (N_23517,N_22672,N_22989);
or U23518 (N_23518,N_22701,N_22933);
nor U23519 (N_23519,N_22960,N_22745);
nand U23520 (N_23520,N_22938,N_22936);
or U23521 (N_23521,N_22956,N_22930);
and U23522 (N_23522,N_22690,N_22772);
nor U23523 (N_23523,N_22654,N_22817);
nor U23524 (N_23524,N_22682,N_22971);
nand U23525 (N_23525,N_23090,N_22823);
and U23526 (N_23526,N_22942,N_22621);
xor U23527 (N_23527,N_22611,N_22858);
nor U23528 (N_23528,N_22814,N_22690);
nor U23529 (N_23529,N_22792,N_22586);
xnor U23530 (N_23530,N_22867,N_22724);
or U23531 (N_23531,N_23010,N_22831);
nor U23532 (N_23532,N_22795,N_22841);
nor U23533 (N_23533,N_22571,N_22893);
and U23534 (N_23534,N_22891,N_22671);
and U23535 (N_23535,N_22802,N_22539);
nand U23536 (N_23536,N_22825,N_22975);
xor U23537 (N_23537,N_22623,N_22955);
and U23538 (N_23538,N_22712,N_23118);
or U23539 (N_23539,N_23123,N_22678);
and U23540 (N_23540,N_23063,N_22634);
or U23541 (N_23541,N_22518,N_22800);
nand U23542 (N_23542,N_23047,N_22506);
xor U23543 (N_23543,N_22683,N_23050);
and U23544 (N_23544,N_22825,N_22779);
nor U23545 (N_23545,N_22703,N_22535);
or U23546 (N_23546,N_22565,N_22796);
nand U23547 (N_23547,N_22721,N_22968);
or U23548 (N_23548,N_22676,N_22689);
and U23549 (N_23549,N_22870,N_22973);
nand U23550 (N_23550,N_22629,N_22613);
nor U23551 (N_23551,N_22510,N_22836);
xnor U23552 (N_23552,N_22660,N_22568);
or U23553 (N_23553,N_22667,N_22954);
xor U23554 (N_23554,N_22804,N_22683);
xnor U23555 (N_23555,N_22706,N_22569);
xor U23556 (N_23556,N_22753,N_23058);
nand U23557 (N_23557,N_22821,N_22624);
and U23558 (N_23558,N_22542,N_22594);
and U23559 (N_23559,N_22551,N_23000);
xnor U23560 (N_23560,N_22937,N_22872);
or U23561 (N_23561,N_22979,N_22687);
xor U23562 (N_23562,N_22567,N_22979);
or U23563 (N_23563,N_22569,N_23095);
nor U23564 (N_23564,N_22530,N_22520);
and U23565 (N_23565,N_22544,N_23083);
xor U23566 (N_23566,N_22800,N_22734);
and U23567 (N_23567,N_22633,N_22794);
and U23568 (N_23568,N_22731,N_22664);
and U23569 (N_23569,N_22569,N_23097);
nor U23570 (N_23570,N_22606,N_22830);
and U23571 (N_23571,N_23056,N_23094);
nand U23572 (N_23572,N_22602,N_23021);
nand U23573 (N_23573,N_22824,N_23028);
nand U23574 (N_23574,N_22548,N_22591);
or U23575 (N_23575,N_23109,N_22773);
or U23576 (N_23576,N_22891,N_22867);
nand U23577 (N_23577,N_22604,N_23075);
or U23578 (N_23578,N_23062,N_22567);
nand U23579 (N_23579,N_22859,N_22728);
xnor U23580 (N_23580,N_22560,N_23040);
xnor U23581 (N_23581,N_22893,N_22601);
xor U23582 (N_23582,N_23017,N_23019);
and U23583 (N_23583,N_22927,N_22809);
and U23584 (N_23584,N_22513,N_22767);
and U23585 (N_23585,N_22587,N_22750);
or U23586 (N_23586,N_23112,N_22790);
xnor U23587 (N_23587,N_22866,N_22941);
nand U23588 (N_23588,N_22938,N_22719);
nand U23589 (N_23589,N_23047,N_23109);
nand U23590 (N_23590,N_22564,N_22699);
and U23591 (N_23591,N_22666,N_22750);
and U23592 (N_23592,N_22763,N_22783);
nor U23593 (N_23593,N_22528,N_22675);
xnor U23594 (N_23594,N_23050,N_23024);
nor U23595 (N_23595,N_23003,N_23116);
or U23596 (N_23596,N_22989,N_22998);
nand U23597 (N_23597,N_23103,N_23058);
nor U23598 (N_23598,N_22912,N_23006);
and U23599 (N_23599,N_22934,N_23094);
nor U23600 (N_23600,N_23013,N_23049);
nand U23601 (N_23601,N_22572,N_22949);
or U23602 (N_23602,N_22996,N_22956);
nand U23603 (N_23603,N_22606,N_22736);
and U23604 (N_23604,N_22668,N_22722);
and U23605 (N_23605,N_22767,N_22678);
nor U23606 (N_23606,N_22677,N_23057);
nor U23607 (N_23607,N_22732,N_22956);
nor U23608 (N_23608,N_22936,N_22682);
and U23609 (N_23609,N_23103,N_22529);
and U23610 (N_23610,N_23124,N_23094);
and U23611 (N_23611,N_22982,N_22834);
or U23612 (N_23612,N_22728,N_22512);
nand U23613 (N_23613,N_23064,N_23103);
nand U23614 (N_23614,N_22701,N_22621);
and U23615 (N_23615,N_22597,N_22811);
or U23616 (N_23616,N_22689,N_22924);
nand U23617 (N_23617,N_23098,N_22856);
xnor U23618 (N_23618,N_22554,N_22908);
nand U23619 (N_23619,N_22569,N_23076);
xnor U23620 (N_23620,N_22973,N_23057);
nor U23621 (N_23621,N_22682,N_22769);
and U23622 (N_23622,N_22843,N_22854);
nor U23623 (N_23623,N_22649,N_22836);
nor U23624 (N_23624,N_22549,N_22894);
nand U23625 (N_23625,N_22973,N_22979);
nand U23626 (N_23626,N_23078,N_22510);
and U23627 (N_23627,N_23009,N_22600);
and U23628 (N_23628,N_22868,N_22604);
or U23629 (N_23629,N_23017,N_22832);
xor U23630 (N_23630,N_22658,N_22574);
nor U23631 (N_23631,N_22923,N_22570);
nor U23632 (N_23632,N_23086,N_23013);
nand U23633 (N_23633,N_22794,N_22600);
nor U23634 (N_23634,N_22791,N_22852);
nor U23635 (N_23635,N_22998,N_22718);
and U23636 (N_23636,N_22967,N_22864);
xor U23637 (N_23637,N_22767,N_22572);
nor U23638 (N_23638,N_22761,N_23063);
nand U23639 (N_23639,N_22688,N_22630);
nor U23640 (N_23640,N_22541,N_22935);
or U23641 (N_23641,N_22542,N_22775);
nor U23642 (N_23642,N_22872,N_22612);
and U23643 (N_23643,N_22687,N_23108);
and U23644 (N_23644,N_22830,N_22598);
and U23645 (N_23645,N_22757,N_22838);
xnor U23646 (N_23646,N_22578,N_23089);
or U23647 (N_23647,N_22717,N_22890);
nor U23648 (N_23648,N_22787,N_22789);
or U23649 (N_23649,N_22533,N_22814);
or U23650 (N_23650,N_22945,N_22792);
xnor U23651 (N_23651,N_22723,N_22540);
nor U23652 (N_23652,N_22522,N_22616);
nand U23653 (N_23653,N_22872,N_22726);
or U23654 (N_23654,N_23060,N_22796);
nor U23655 (N_23655,N_22552,N_22839);
or U23656 (N_23656,N_22986,N_22574);
or U23657 (N_23657,N_22812,N_22930);
nor U23658 (N_23658,N_22803,N_22639);
and U23659 (N_23659,N_22765,N_22807);
nand U23660 (N_23660,N_22943,N_23050);
nand U23661 (N_23661,N_22890,N_22814);
and U23662 (N_23662,N_22607,N_22822);
nor U23663 (N_23663,N_23092,N_22909);
nand U23664 (N_23664,N_22684,N_22692);
or U23665 (N_23665,N_22750,N_22963);
xnor U23666 (N_23666,N_22927,N_22659);
nand U23667 (N_23667,N_22591,N_22612);
nand U23668 (N_23668,N_22854,N_23010);
xor U23669 (N_23669,N_22711,N_22514);
or U23670 (N_23670,N_22801,N_22885);
nor U23671 (N_23671,N_23013,N_22871);
or U23672 (N_23672,N_22837,N_22674);
xor U23673 (N_23673,N_22909,N_22564);
nor U23674 (N_23674,N_23038,N_23082);
xnor U23675 (N_23675,N_23110,N_22924);
xor U23676 (N_23676,N_23105,N_22936);
and U23677 (N_23677,N_22598,N_22601);
or U23678 (N_23678,N_22838,N_22530);
nor U23679 (N_23679,N_23106,N_22622);
nand U23680 (N_23680,N_22734,N_22950);
nor U23681 (N_23681,N_23040,N_22632);
or U23682 (N_23682,N_22642,N_22923);
or U23683 (N_23683,N_23095,N_23046);
nor U23684 (N_23684,N_22976,N_23018);
or U23685 (N_23685,N_22764,N_23085);
nor U23686 (N_23686,N_23092,N_22821);
or U23687 (N_23687,N_22713,N_22973);
or U23688 (N_23688,N_22911,N_22670);
and U23689 (N_23689,N_22806,N_22739);
xnor U23690 (N_23690,N_22916,N_22803);
and U23691 (N_23691,N_22850,N_22899);
nand U23692 (N_23692,N_22730,N_22507);
nor U23693 (N_23693,N_22754,N_23079);
xnor U23694 (N_23694,N_22691,N_22991);
nand U23695 (N_23695,N_22981,N_23025);
nor U23696 (N_23696,N_22756,N_22527);
nand U23697 (N_23697,N_22535,N_22714);
nor U23698 (N_23698,N_22978,N_23100);
nor U23699 (N_23699,N_22909,N_23061);
and U23700 (N_23700,N_22824,N_23009);
and U23701 (N_23701,N_22568,N_22991);
nand U23702 (N_23702,N_23083,N_22791);
or U23703 (N_23703,N_22877,N_22694);
or U23704 (N_23704,N_23071,N_22833);
nand U23705 (N_23705,N_22554,N_22508);
nor U23706 (N_23706,N_23082,N_22861);
nand U23707 (N_23707,N_23039,N_23014);
xor U23708 (N_23708,N_22593,N_23010);
nand U23709 (N_23709,N_23048,N_23116);
or U23710 (N_23710,N_22532,N_23020);
xor U23711 (N_23711,N_22626,N_23029);
or U23712 (N_23712,N_22776,N_22774);
nand U23713 (N_23713,N_23006,N_22605);
and U23714 (N_23714,N_23002,N_22913);
nor U23715 (N_23715,N_22590,N_22558);
nand U23716 (N_23716,N_22662,N_22780);
nor U23717 (N_23717,N_22907,N_22576);
xor U23718 (N_23718,N_22951,N_22843);
xnor U23719 (N_23719,N_22647,N_22931);
or U23720 (N_23720,N_23041,N_22805);
nor U23721 (N_23721,N_22955,N_22642);
nor U23722 (N_23722,N_22648,N_22962);
xor U23723 (N_23723,N_23079,N_22624);
and U23724 (N_23724,N_22570,N_22942);
xnor U23725 (N_23725,N_22639,N_22916);
and U23726 (N_23726,N_23004,N_22772);
xor U23727 (N_23727,N_22506,N_23006);
or U23728 (N_23728,N_22619,N_22623);
xnor U23729 (N_23729,N_22633,N_22742);
and U23730 (N_23730,N_22623,N_23044);
and U23731 (N_23731,N_22830,N_22918);
or U23732 (N_23732,N_22807,N_22793);
or U23733 (N_23733,N_22536,N_22656);
nor U23734 (N_23734,N_23111,N_22583);
xnor U23735 (N_23735,N_22825,N_22589);
nor U23736 (N_23736,N_22863,N_22760);
and U23737 (N_23737,N_23038,N_22833);
and U23738 (N_23738,N_22869,N_22544);
nand U23739 (N_23739,N_23033,N_22753);
or U23740 (N_23740,N_23066,N_22656);
nor U23741 (N_23741,N_22712,N_22509);
and U23742 (N_23742,N_22635,N_22970);
nor U23743 (N_23743,N_22810,N_22866);
or U23744 (N_23744,N_22605,N_22718);
nor U23745 (N_23745,N_22541,N_22892);
xnor U23746 (N_23746,N_23083,N_22574);
or U23747 (N_23747,N_22579,N_22559);
nor U23748 (N_23748,N_22715,N_22830);
nor U23749 (N_23749,N_22630,N_22795);
nand U23750 (N_23750,N_23172,N_23214);
nand U23751 (N_23751,N_23454,N_23663);
nand U23752 (N_23752,N_23370,N_23287);
xnor U23753 (N_23753,N_23677,N_23338);
nand U23754 (N_23754,N_23162,N_23192);
xor U23755 (N_23755,N_23247,N_23188);
xor U23756 (N_23756,N_23424,N_23455);
and U23757 (N_23757,N_23461,N_23489);
nand U23758 (N_23758,N_23505,N_23198);
xor U23759 (N_23759,N_23436,N_23584);
nor U23760 (N_23760,N_23518,N_23204);
or U23761 (N_23761,N_23342,N_23711);
nand U23762 (N_23762,N_23682,N_23709);
or U23763 (N_23763,N_23208,N_23405);
and U23764 (N_23764,N_23353,N_23136);
or U23765 (N_23765,N_23612,N_23327);
xor U23766 (N_23766,N_23235,N_23263);
and U23767 (N_23767,N_23652,N_23134);
nor U23768 (N_23768,N_23252,N_23474);
or U23769 (N_23769,N_23499,N_23240);
xor U23770 (N_23770,N_23175,N_23275);
nor U23771 (N_23771,N_23656,N_23444);
nand U23772 (N_23772,N_23440,N_23699);
and U23773 (N_23773,N_23435,N_23278);
nor U23774 (N_23774,N_23328,N_23325);
and U23775 (N_23775,N_23193,N_23725);
xnor U23776 (N_23776,N_23265,N_23271);
and U23777 (N_23777,N_23254,N_23651);
or U23778 (N_23778,N_23243,N_23485);
nor U23779 (N_23779,N_23641,N_23572);
nor U23780 (N_23780,N_23391,N_23167);
and U23781 (N_23781,N_23521,N_23256);
or U23782 (N_23782,N_23675,N_23698);
xor U23783 (N_23783,N_23481,N_23697);
and U23784 (N_23784,N_23385,N_23470);
and U23785 (N_23785,N_23422,N_23230);
nand U23786 (N_23786,N_23558,N_23257);
or U23787 (N_23787,N_23219,N_23330);
or U23788 (N_23788,N_23678,N_23222);
or U23789 (N_23789,N_23732,N_23463);
xor U23790 (N_23790,N_23127,N_23365);
nor U23791 (N_23791,N_23524,N_23626);
xnor U23792 (N_23792,N_23442,N_23429);
and U23793 (N_23793,N_23593,N_23234);
nor U23794 (N_23794,N_23592,N_23180);
xor U23795 (N_23795,N_23186,N_23722);
and U23796 (N_23796,N_23532,N_23418);
or U23797 (N_23797,N_23655,N_23588);
or U23798 (N_23798,N_23143,N_23272);
nor U23799 (N_23799,N_23415,N_23406);
and U23800 (N_23800,N_23540,N_23494);
xnor U23801 (N_23801,N_23289,N_23610);
xor U23802 (N_23802,N_23684,N_23246);
and U23803 (N_23803,N_23182,N_23479);
and U23804 (N_23804,N_23163,N_23207);
xor U23805 (N_23805,N_23467,N_23377);
and U23806 (N_23806,N_23210,N_23332);
xor U23807 (N_23807,N_23191,N_23431);
nor U23808 (N_23808,N_23720,N_23129);
or U23809 (N_23809,N_23335,N_23279);
and U23810 (N_23810,N_23323,N_23346);
nor U23811 (N_23811,N_23449,N_23183);
nand U23812 (N_23812,N_23233,N_23329);
xnor U23813 (N_23813,N_23413,N_23423);
nor U23814 (N_23814,N_23586,N_23748);
and U23815 (N_23815,N_23139,N_23595);
xnor U23816 (N_23816,N_23303,N_23645);
xnor U23817 (N_23817,N_23340,N_23273);
or U23818 (N_23818,N_23533,N_23383);
nor U23819 (N_23819,N_23157,N_23491);
and U23820 (N_23820,N_23648,N_23591);
nor U23821 (N_23821,N_23304,N_23511);
nand U23822 (N_23822,N_23637,N_23149);
xor U23823 (N_23823,N_23636,N_23417);
nand U23824 (N_23824,N_23669,N_23613);
nand U23825 (N_23825,N_23421,N_23553);
nand U23826 (N_23826,N_23199,N_23217);
nand U23827 (N_23827,N_23245,N_23556);
and U23828 (N_23828,N_23380,N_23409);
nor U23829 (N_23829,N_23313,N_23476);
and U23830 (N_23830,N_23439,N_23482);
nand U23831 (N_23831,N_23293,N_23715);
or U23832 (N_23832,N_23140,N_23466);
xnor U23833 (N_23833,N_23742,N_23384);
xnor U23834 (N_23834,N_23507,N_23402);
nor U23835 (N_23835,N_23220,N_23559);
and U23836 (N_23836,N_23181,N_23398);
and U23837 (N_23837,N_23635,N_23729);
nand U23838 (N_23838,N_23331,N_23687);
and U23839 (N_23839,N_23185,N_23269);
nand U23840 (N_23840,N_23412,N_23375);
or U23841 (N_23841,N_23622,N_23253);
nor U23842 (N_23842,N_23512,N_23548);
or U23843 (N_23843,N_23570,N_23483);
or U23844 (N_23844,N_23708,N_23583);
nor U23845 (N_23845,N_23379,N_23647);
xnor U23846 (N_23846,N_23710,N_23343);
nand U23847 (N_23847,N_23724,N_23236);
xor U23848 (N_23848,N_23561,N_23721);
nand U23849 (N_23849,N_23224,N_23676);
nor U23850 (N_23850,N_23665,N_23369);
nor U23851 (N_23851,N_23602,N_23258);
xor U23852 (N_23852,N_23696,N_23357);
nand U23853 (N_23853,N_23128,N_23427);
xnor U23854 (N_23854,N_23268,N_23250);
nor U23855 (N_23855,N_23196,N_23259);
xor U23856 (N_23856,N_23156,N_23226);
nand U23857 (N_23857,N_23336,N_23453);
and U23858 (N_23858,N_23373,N_23450);
or U23859 (N_23859,N_23350,N_23419);
xor U23860 (N_23860,N_23484,N_23414);
or U23861 (N_23861,N_23364,N_23568);
and U23862 (N_23862,N_23301,N_23577);
xor U23863 (N_23863,N_23351,N_23542);
nor U23864 (N_23864,N_23171,N_23194);
xnor U23865 (N_23865,N_23623,N_23437);
nand U23866 (N_23866,N_23155,N_23575);
xor U23867 (N_23867,N_23374,N_23501);
nand U23868 (N_23868,N_23206,N_23739);
and U23869 (N_23869,N_23529,N_23526);
xnor U23870 (N_23870,N_23667,N_23161);
or U23871 (N_23871,N_23598,N_23174);
or U23872 (N_23872,N_23281,N_23490);
and U23873 (N_23873,N_23352,N_23694);
nand U23874 (N_23874,N_23309,N_23160);
nor U23875 (N_23875,N_23165,N_23471);
nor U23876 (N_23876,N_23154,N_23270);
nor U23877 (N_23877,N_23541,N_23685);
and U23878 (N_23878,N_23337,N_23625);
nor U23879 (N_23879,N_23286,N_23606);
xnor U23880 (N_23880,N_23552,N_23177);
nand U23881 (N_23881,N_23680,N_23689);
and U23882 (N_23882,N_23496,N_23513);
xor U23883 (N_23883,N_23433,N_23312);
nor U23884 (N_23884,N_23514,N_23349);
nand U23885 (N_23885,N_23280,N_23639);
nor U23886 (N_23886,N_23447,N_23142);
and U23887 (N_23887,N_23438,N_23544);
nand U23888 (N_23888,N_23321,N_23173);
or U23889 (N_23889,N_23536,N_23305);
nor U23890 (N_23890,N_23363,N_23658);
nand U23891 (N_23891,N_23430,N_23679);
or U23892 (N_23892,N_23695,N_23747);
nand U23893 (N_23893,N_23441,N_23251);
xnor U23894 (N_23894,N_23649,N_23492);
xnor U23895 (N_23895,N_23152,N_23306);
nand U23896 (N_23896,N_23378,N_23469);
or U23897 (N_23897,N_23451,N_23371);
xnor U23898 (N_23898,N_23642,N_23345);
xnor U23899 (N_23899,N_23218,N_23672);
nand U23900 (N_23900,N_23630,N_23277);
or U23901 (N_23901,N_23712,N_23334);
or U23902 (N_23902,N_23509,N_23580);
and U23903 (N_23903,N_23459,N_23516);
xor U23904 (N_23904,N_23632,N_23617);
nand U23905 (N_23905,N_23315,N_23587);
nor U23906 (N_23906,N_23464,N_23493);
nor U23907 (N_23907,N_23566,N_23590);
or U23908 (N_23908,N_23594,N_23576);
nand U23909 (N_23909,N_23307,N_23569);
nor U23910 (N_23910,N_23388,N_23151);
nor U23911 (N_23911,N_23434,N_23426);
nand U23912 (N_23912,N_23504,N_23531);
nor U23913 (N_23913,N_23164,N_23394);
xor U23914 (N_23914,N_23241,N_23389);
and U23915 (N_23915,N_23189,N_23734);
nand U23916 (N_23916,N_23411,N_23551);
nand U23917 (N_23917,N_23457,N_23141);
or U23918 (N_23918,N_23387,N_23316);
nand U23919 (N_23919,N_23131,N_23700);
nor U23920 (N_23920,N_23452,N_23497);
nand U23921 (N_23921,N_23376,N_23508);
or U23922 (N_23922,N_23231,N_23582);
nor U23923 (N_23923,N_23298,N_23232);
nor U23924 (N_23924,N_23654,N_23537);
nor U23925 (N_23925,N_23618,N_23660);
and U23926 (N_23926,N_23264,N_23554);
nor U23927 (N_23927,N_23673,N_23187);
or U23928 (N_23928,N_23318,N_23360);
xnor U23929 (N_23929,N_23738,N_23624);
nor U23930 (N_23930,N_23611,N_23614);
nor U23931 (N_23931,N_23314,N_23130);
xnor U23932 (N_23932,N_23666,N_23714);
or U23933 (N_23933,N_23627,N_23239);
or U23934 (N_23934,N_23486,N_23659);
nand U23935 (N_23935,N_23215,N_23460);
nor U23936 (N_23936,N_23297,N_23302);
nor U23937 (N_23937,N_23539,N_23547);
nand U23938 (N_23938,N_23535,N_23705);
and U23939 (N_23939,N_23744,N_23179);
nor U23940 (N_23940,N_23503,N_23520);
nand U23941 (N_23941,N_23367,N_23135);
or U23942 (N_23942,N_23223,N_23657);
nor U23943 (N_23943,N_23213,N_23468);
and U23944 (N_23944,N_23132,N_23145);
or U23945 (N_23945,N_23604,N_23557);
nor U23946 (N_23946,N_23170,N_23634);
or U23947 (N_23947,N_23545,N_23150);
nand U23948 (N_23948,N_23153,N_23361);
or U23949 (N_23949,N_23344,N_23644);
nand U23950 (N_23950,N_23146,N_23740);
nor U23951 (N_23951,N_23144,N_23716);
nand U23952 (N_23952,N_23359,N_23176);
nand U23953 (N_23953,N_23727,N_23190);
or U23954 (N_23954,N_23299,N_23478);
and U23955 (N_23955,N_23502,N_23341);
xnor U23956 (N_23956,N_23530,N_23719);
nor U23957 (N_23957,N_23358,N_23643);
nor U23958 (N_23958,N_23605,N_23290);
nor U23959 (N_23959,N_23456,N_23515);
or U23960 (N_23960,N_23354,N_23650);
xnor U23961 (N_23961,N_23543,N_23601);
nor U23962 (N_23962,N_23211,N_23138);
nor U23963 (N_23963,N_23395,N_23731);
or U23964 (N_23964,N_23326,N_23683);
xor U23965 (N_23965,N_23619,N_23495);
and U23966 (N_23966,N_23368,N_23549);
and U23967 (N_23967,N_23283,N_23274);
xor U23968 (N_23968,N_23227,N_23184);
nand U23969 (N_23969,N_23525,N_23631);
or U23970 (N_23970,N_23229,N_23372);
or U23971 (N_23971,N_23599,N_23693);
nor U23972 (N_23972,N_23147,N_23465);
nor U23973 (N_23973,N_23473,N_23248);
nor U23974 (N_23974,N_23324,N_23362);
xor U23975 (N_23975,N_23500,N_23661);
nor U23976 (N_23976,N_23237,N_23596);
nor U23977 (N_23977,N_23261,N_23550);
nand U23978 (N_23978,N_23581,N_23565);
and U23979 (N_23979,N_23670,N_23446);
nand U23980 (N_23980,N_23589,N_23730);
and U23981 (N_23981,N_23242,N_23472);
or U23982 (N_23982,N_23646,N_23339);
and U23983 (N_23983,N_23311,N_23487);
and U23984 (N_23984,N_23203,N_23523);
or U23985 (N_23985,N_23212,N_23462);
nor U23986 (N_23986,N_23690,N_23717);
nor U23987 (N_23987,N_23458,N_23662);
and U23988 (N_23988,N_23638,N_23578);
nor U23989 (N_23989,N_23510,N_23169);
xor U23990 (N_23990,N_23713,N_23317);
nand U23991 (N_23991,N_23749,N_23585);
nand U23992 (N_23992,N_23333,N_23216);
xnor U23993 (N_23993,N_23195,N_23355);
and U23994 (N_23994,N_23126,N_23322);
nor U23995 (N_23995,N_23420,N_23228);
nor U23996 (N_23996,N_23607,N_23407);
nor U23997 (N_23997,N_23562,N_23498);
xor U23998 (N_23998,N_23528,N_23480);
and U23999 (N_23999,N_23291,N_23396);
and U24000 (N_24000,N_23621,N_23288);
nand U24001 (N_24001,N_23159,N_23506);
xnor U24002 (N_24002,N_23640,N_23178);
nand U24003 (N_24003,N_23600,N_23671);
and U24004 (N_24004,N_23428,N_23347);
xnor U24005 (N_24005,N_23267,N_23706);
nor U24006 (N_24006,N_23320,N_23704);
xnor U24007 (N_24007,N_23262,N_23382);
nand U24008 (N_24008,N_23201,N_23432);
nand U24009 (N_24009,N_23616,N_23633);
and U24010 (N_24010,N_23563,N_23205);
and U24011 (N_24011,N_23608,N_23366);
or U24012 (N_24012,N_23733,N_23445);
or U24013 (N_24013,N_23238,N_23282);
xor U24014 (N_24014,N_23443,N_23381);
or U24015 (N_24015,N_23688,N_23517);
nand U24016 (N_24016,N_23404,N_23166);
xor U24017 (N_24017,N_23403,N_23475);
nand U24018 (N_24018,N_23664,N_23628);
and U24019 (N_24019,N_23538,N_23284);
nor U24020 (N_24020,N_23276,N_23488);
and U24021 (N_24021,N_23133,N_23620);
or U24022 (N_24022,N_23410,N_23527);
nor U24023 (N_24023,N_23386,N_23702);
or U24024 (N_24024,N_23266,N_23597);
nor U24025 (N_24025,N_23200,N_23448);
and U24026 (N_24026,N_23158,N_23197);
or U24027 (N_24027,N_23701,N_23477);
xor U24028 (N_24028,N_23629,N_23723);
or U24029 (N_24029,N_23292,N_23209);
xnor U24030 (N_24030,N_23137,N_23728);
or U24031 (N_24031,N_23168,N_23603);
nand U24032 (N_24032,N_23310,N_23564);
or U24033 (N_24033,N_23609,N_23348);
xnor U24034 (N_24034,N_23686,N_23737);
nor U24035 (N_24035,N_23125,N_23703);
or U24036 (N_24036,N_23615,N_23285);
nor U24037 (N_24037,N_23393,N_23745);
nor U24038 (N_24038,N_23743,N_23244);
nor U24039 (N_24039,N_23319,N_23735);
xnor U24040 (N_24040,N_23397,N_23401);
xor U24041 (N_24041,N_23399,N_23408);
nor U24042 (N_24042,N_23392,N_23726);
or U24043 (N_24043,N_23560,N_23567);
nor U24044 (N_24044,N_23718,N_23300);
and U24045 (N_24045,N_23522,N_23546);
xor U24046 (N_24046,N_23579,N_23681);
or U24047 (N_24047,N_23221,N_23425);
or U24048 (N_24048,N_23653,N_23519);
or U24049 (N_24049,N_23707,N_23741);
nand U24050 (N_24050,N_23249,N_23296);
nand U24051 (N_24051,N_23416,N_23295);
xnor U24052 (N_24052,N_23534,N_23668);
nor U24053 (N_24053,N_23260,N_23308);
nor U24054 (N_24054,N_23356,N_23400);
nor U24055 (N_24055,N_23255,N_23574);
nor U24056 (N_24056,N_23571,N_23691);
xnor U24057 (N_24057,N_23746,N_23148);
nand U24058 (N_24058,N_23736,N_23390);
nand U24059 (N_24059,N_23692,N_23202);
nor U24060 (N_24060,N_23573,N_23555);
or U24061 (N_24061,N_23674,N_23225);
nor U24062 (N_24062,N_23294,N_23243);
xor U24063 (N_24063,N_23279,N_23221);
nor U24064 (N_24064,N_23593,N_23261);
xor U24065 (N_24065,N_23255,N_23693);
and U24066 (N_24066,N_23408,N_23664);
nand U24067 (N_24067,N_23521,N_23339);
or U24068 (N_24068,N_23730,N_23446);
nor U24069 (N_24069,N_23449,N_23323);
nand U24070 (N_24070,N_23556,N_23147);
and U24071 (N_24071,N_23270,N_23244);
or U24072 (N_24072,N_23146,N_23721);
xnor U24073 (N_24073,N_23462,N_23358);
xnor U24074 (N_24074,N_23220,N_23736);
xnor U24075 (N_24075,N_23615,N_23174);
nand U24076 (N_24076,N_23149,N_23397);
and U24077 (N_24077,N_23469,N_23406);
nor U24078 (N_24078,N_23368,N_23230);
xor U24079 (N_24079,N_23309,N_23195);
nand U24080 (N_24080,N_23316,N_23261);
and U24081 (N_24081,N_23134,N_23741);
or U24082 (N_24082,N_23211,N_23529);
nor U24083 (N_24083,N_23314,N_23437);
xor U24084 (N_24084,N_23150,N_23325);
and U24085 (N_24085,N_23572,N_23668);
and U24086 (N_24086,N_23525,N_23590);
and U24087 (N_24087,N_23700,N_23635);
or U24088 (N_24088,N_23449,N_23268);
and U24089 (N_24089,N_23672,N_23345);
xnor U24090 (N_24090,N_23495,N_23602);
nor U24091 (N_24091,N_23378,N_23698);
or U24092 (N_24092,N_23172,N_23133);
nor U24093 (N_24093,N_23228,N_23629);
xor U24094 (N_24094,N_23646,N_23404);
and U24095 (N_24095,N_23290,N_23500);
xor U24096 (N_24096,N_23732,N_23483);
and U24097 (N_24097,N_23524,N_23576);
nor U24098 (N_24098,N_23351,N_23487);
nor U24099 (N_24099,N_23629,N_23342);
nor U24100 (N_24100,N_23251,N_23506);
or U24101 (N_24101,N_23560,N_23485);
or U24102 (N_24102,N_23356,N_23564);
xnor U24103 (N_24103,N_23644,N_23321);
xor U24104 (N_24104,N_23141,N_23618);
nor U24105 (N_24105,N_23453,N_23725);
or U24106 (N_24106,N_23489,N_23631);
and U24107 (N_24107,N_23352,N_23482);
or U24108 (N_24108,N_23456,N_23229);
or U24109 (N_24109,N_23687,N_23521);
or U24110 (N_24110,N_23431,N_23472);
or U24111 (N_24111,N_23178,N_23526);
and U24112 (N_24112,N_23687,N_23370);
xor U24113 (N_24113,N_23498,N_23163);
xor U24114 (N_24114,N_23694,N_23364);
xnor U24115 (N_24115,N_23184,N_23138);
and U24116 (N_24116,N_23159,N_23372);
or U24117 (N_24117,N_23708,N_23475);
nand U24118 (N_24118,N_23736,N_23644);
or U24119 (N_24119,N_23507,N_23323);
and U24120 (N_24120,N_23361,N_23525);
or U24121 (N_24121,N_23245,N_23517);
nand U24122 (N_24122,N_23457,N_23514);
and U24123 (N_24123,N_23242,N_23396);
xnor U24124 (N_24124,N_23304,N_23137);
and U24125 (N_24125,N_23495,N_23605);
or U24126 (N_24126,N_23698,N_23561);
and U24127 (N_24127,N_23191,N_23276);
and U24128 (N_24128,N_23229,N_23708);
nor U24129 (N_24129,N_23192,N_23693);
or U24130 (N_24130,N_23712,N_23199);
or U24131 (N_24131,N_23209,N_23405);
xnor U24132 (N_24132,N_23344,N_23204);
nor U24133 (N_24133,N_23300,N_23229);
xnor U24134 (N_24134,N_23722,N_23641);
or U24135 (N_24135,N_23147,N_23694);
and U24136 (N_24136,N_23446,N_23372);
nor U24137 (N_24137,N_23322,N_23541);
xnor U24138 (N_24138,N_23271,N_23609);
and U24139 (N_24139,N_23160,N_23199);
or U24140 (N_24140,N_23225,N_23180);
or U24141 (N_24141,N_23604,N_23225);
nand U24142 (N_24142,N_23587,N_23359);
nor U24143 (N_24143,N_23351,N_23533);
xor U24144 (N_24144,N_23211,N_23550);
xnor U24145 (N_24145,N_23286,N_23586);
and U24146 (N_24146,N_23148,N_23397);
nand U24147 (N_24147,N_23548,N_23594);
or U24148 (N_24148,N_23314,N_23294);
nor U24149 (N_24149,N_23724,N_23141);
nor U24150 (N_24150,N_23706,N_23407);
or U24151 (N_24151,N_23221,N_23329);
nand U24152 (N_24152,N_23266,N_23530);
xor U24153 (N_24153,N_23665,N_23611);
or U24154 (N_24154,N_23291,N_23309);
or U24155 (N_24155,N_23580,N_23721);
nor U24156 (N_24156,N_23686,N_23521);
or U24157 (N_24157,N_23462,N_23605);
xor U24158 (N_24158,N_23280,N_23361);
xor U24159 (N_24159,N_23134,N_23558);
or U24160 (N_24160,N_23611,N_23327);
or U24161 (N_24161,N_23236,N_23501);
nor U24162 (N_24162,N_23280,N_23657);
nand U24163 (N_24163,N_23276,N_23151);
and U24164 (N_24164,N_23466,N_23740);
xnor U24165 (N_24165,N_23659,N_23537);
nand U24166 (N_24166,N_23300,N_23629);
nor U24167 (N_24167,N_23320,N_23631);
nor U24168 (N_24168,N_23645,N_23749);
or U24169 (N_24169,N_23275,N_23601);
xor U24170 (N_24170,N_23214,N_23675);
nand U24171 (N_24171,N_23609,N_23350);
nor U24172 (N_24172,N_23475,N_23198);
or U24173 (N_24173,N_23708,N_23603);
nand U24174 (N_24174,N_23239,N_23179);
nor U24175 (N_24175,N_23690,N_23173);
xnor U24176 (N_24176,N_23544,N_23561);
nor U24177 (N_24177,N_23409,N_23253);
or U24178 (N_24178,N_23540,N_23478);
or U24179 (N_24179,N_23449,N_23228);
and U24180 (N_24180,N_23737,N_23677);
and U24181 (N_24181,N_23345,N_23455);
nor U24182 (N_24182,N_23194,N_23284);
xnor U24183 (N_24183,N_23343,N_23564);
xnor U24184 (N_24184,N_23389,N_23749);
and U24185 (N_24185,N_23201,N_23148);
or U24186 (N_24186,N_23591,N_23474);
and U24187 (N_24187,N_23580,N_23731);
xnor U24188 (N_24188,N_23310,N_23331);
or U24189 (N_24189,N_23372,N_23732);
or U24190 (N_24190,N_23320,N_23218);
or U24191 (N_24191,N_23651,N_23203);
and U24192 (N_24192,N_23322,N_23151);
nor U24193 (N_24193,N_23628,N_23311);
nand U24194 (N_24194,N_23386,N_23495);
nor U24195 (N_24195,N_23351,N_23588);
xnor U24196 (N_24196,N_23420,N_23156);
xnor U24197 (N_24197,N_23167,N_23620);
and U24198 (N_24198,N_23343,N_23673);
xnor U24199 (N_24199,N_23348,N_23611);
xor U24200 (N_24200,N_23404,N_23302);
or U24201 (N_24201,N_23265,N_23365);
xnor U24202 (N_24202,N_23616,N_23586);
nor U24203 (N_24203,N_23372,N_23300);
and U24204 (N_24204,N_23408,N_23715);
and U24205 (N_24205,N_23721,N_23538);
xnor U24206 (N_24206,N_23670,N_23133);
nand U24207 (N_24207,N_23298,N_23643);
xor U24208 (N_24208,N_23448,N_23347);
or U24209 (N_24209,N_23691,N_23457);
or U24210 (N_24210,N_23211,N_23673);
or U24211 (N_24211,N_23232,N_23474);
or U24212 (N_24212,N_23192,N_23499);
xnor U24213 (N_24213,N_23369,N_23268);
or U24214 (N_24214,N_23401,N_23578);
or U24215 (N_24215,N_23729,N_23415);
or U24216 (N_24216,N_23484,N_23251);
xnor U24217 (N_24217,N_23426,N_23541);
nor U24218 (N_24218,N_23240,N_23415);
xor U24219 (N_24219,N_23580,N_23531);
or U24220 (N_24220,N_23510,N_23172);
and U24221 (N_24221,N_23637,N_23180);
xnor U24222 (N_24222,N_23321,N_23267);
nand U24223 (N_24223,N_23374,N_23435);
and U24224 (N_24224,N_23368,N_23446);
and U24225 (N_24225,N_23314,N_23155);
nand U24226 (N_24226,N_23613,N_23144);
nor U24227 (N_24227,N_23451,N_23656);
or U24228 (N_24228,N_23244,N_23653);
and U24229 (N_24229,N_23671,N_23655);
xor U24230 (N_24230,N_23636,N_23517);
or U24231 (N_24231,N_23484,N_23297);
xnor U24232 (N_24232,N_23675,N_23176);
and U24233 (N_24233,N_23250,N_23696);
or U24234 (N_24234,N_23654,N_23743);
xnor U24235 (N_24235,N_23629,N_23423);
nand U24236 (N_24236,N_23489,N_23335);
and U24237 (N_24237,N_23512,N_23145);
nor U24238 (N_24238,N_23149,N_23564);
xnor U24239 (N_24239,N_23221,N_23493);
and U24240 (N_24240,N_23203,N_23597);
and U24241 (N_24241,N_23266,N_23556);
xor U24242 (N_24242,N_23381,N_23535);
or U24243 (N_24243,N_23433,N_23646);
xnor U24244 (N_24244,N_23360,N_23526);
xor U24245 (N_24245,N_23740,N_23167);
xor U24246 (N_24246,N_23682,N_23183);
or U24247 (N_24247,N_23368,N_23377);
nor U24248 (N_24248,N_23223,N_23555);
nor U24249 (N_24249,N_23412,N_23607);
nand U24250 (N_24250,N_23295,N_23569);
or U24251 (N_24251,N_23377,N_23158);
xor U24252 (N_24252,N_23434,N_23307);
xnor U24253 (N_24253,N_23483,N_23724);
or U24254 (N_24254,N_23140,N_23162);
and U24255 (N_24255,N_23448,N_23188);
or U24256 (N_24256,N_23289,N_23682);
nor U24257 (N_24257,N_23167,N_23555);
and U24258 (N_24258,N_23337,N_23325);
or U24259 (N_24259,N_23434,N_23331);
or U24260 (N_24260,N_23688,N_23544);
or U24261 (N_24261,N_23747,N_23407);
xor U24262 (N_24262,N_23449,N_23634);
nand U24263 (N_24263,N_23501,N_23591);
nand U24264 (N_24264,N_23511,N_23694);
xor U24265 (N_24265,N_23395,N_23346);
xor U24266 (N_24266,N_23641,N_23510);
or U24267 (N_24267,N_23250,N_23708);
or U24268 (N_24268,N_23308,N_23183);
or U24269 (N_24269,N_23606,N_23348);
nand U24270 (N_24270,N_23260,N_23632);
xnor U24271 (N_24271,N_23667,N_23703);
xnor U24272 (N_24272,N_23379,N_23653);
and U24273 (N_24273,N_23511,N_23126);
and U24274 (N_24274,N_23281,N_23565);
xor U24275 (N_24275,N_23250,N_23506);
nand U24276 (N_24276,N_23525,N_23188);
or U24277 (N_24277,N_23458,N_23223);
nand U24278 (N_24278,N_23430,N_23489);
nor U24279 (N_24279,N_23284,N_23278);
nand U24280 (N_24280,N_23578,N_23521);
nor U24281 (N_24281,N_23421,N_23680);
or U24282 (N_24282,N_23489,N_23130);
or U24283 (N_24283,N_23670,N_23368);
nand U24284 (N_24284,N_23190,N_23278);
or U24285 (N_24285,N_23552,N_23256);
xor U24286 (N_24286,N_23400,N_23315);
nand U24287 (N_24287,N_23453,N_23624);
and U24288 (N_24288,N_23705,N_23719);
xnor U24289 (N_24289,N_23266,N_23382);
and U24290 (N_24290,N_23371,N_23178);
xnor U24291 (N_24291,N_23606,N_23373);
and U24292 (N_24292,N_23618,N_23392);
and U24293 (N_24293,N_23512,N_23592);
and U24294 (N_24294,N_23183,N_23382);
and U24295 (N_24295,N_23462,N_23553);
xnor U24296 (N_24296,N_23699,N_23299);
nor U24297 (N_24297,N_23321,N_23432);
xnor U24298 (N_24298,N_23349,N_23396);
and U24299 (N_24299,N_23680,N_23361);
nor U24300 (N_24300,N_23502,N_23307);
and U24301 (N_24301,N_23548,N_23284);
xnor U24302 (N_24302,N_23320,N_23250);
nor U24303 (N_24303,N_23177,N_23353);
nor U24304 (N_24304,N_23238,N_23444);
xnor U24305 (N_24305,N_23730,N_23542);
and U24306 (N_24306,N_23299,N_23644);
and U24307 (N_24307,N_23172,N_23396);
nor U24308 (N_24308,N_23729,N_23437);
nor U24309 (N_24309,N_23197,N_23534);
or U24310 (N_24310,N_23661,N_23550);
nand U24311 (N_24311,N_23698,N_23311);
xnor U24312 (N_24312,N_23469,N_23345);
xor U24313 (N_24313,N_23497,N_23646);
nand U24314 (N_24314,N_23730,N_23650);
or U24315 (N_24315,N_23512,N_23640);
nand U24316 (N_24316,N_23162,N_23132);
nor U24317 (N_24317,N_23358,N_23520);
nor U24318 (N_24318,N_23277,N_23422);
xnor U24319 (N_24319,N_23370,N_23696);
or U24320 (N_24320,N_23671,N_23129);
nand U24321 (N_24321,N_23226,N_23545);
xnor U24322 (N_24322,N_23180,N_23518);
or U24323 (N_24323,N_23393,N_23215);
and U24324 (N_24324,N_23731,N_23544);
nand U24325 (N_24325,N_23526,N_23139);
xor U24326 (N_24326,N_23479,N_23665);
xnor U24327 (N_24327,N_23619,N_23205);
nor U24328 (N_24328,N_23531,N_23585);
or U24329 (N_24329,N_23604,N_23541);
and U24330 (N_24330,N_23609,N_23145);
xor U24331 (N_24331,N_23138,N_23634);
or U24332 (N_24332,N_23537,N_23680);
nor U24333 (N_24333,N_23616,N_23200);
or U24334 (N_24334,N_23314,N_23215);
nand U24335 (N_24335,N_23498,N_23614);
or U24336 (N_24336,N_23282,N_23471);
xnor U24337 (N_24337,N_23181,N_23282);
nor U24338 (N_24338,N_23329,N_23569);
or U24339 (N_24339,N_23710,N_23727);
and U24340 (N_24340,N_23725,N_23354);
nand U24341 (N_24341,N_23281,N_23245);
nor U24342 (N_24342,N_23368,N_23480);
xnor U24343 (N_24343,N_23260,N_23658);
xor U24344 (N_24344,N_23203,N_23632);
or U24345 (N_24345,N_23252,N_23270);
nor U24346 (N_24346,N_23267,N_23187);
or U24347 (N_24347,N_23681,N_23660);
nand U24348 (N_24348,N_23723,N_23597);
and U24349 (N_24349,N_23222,N_23349);
nor U24350 (N_24350,N_23264,N_23696);
nand U24351 (N_24351,N_23185,N_23217);
xor U24352 (N_24352,N_23624,N_23174);
nand U24353 (N_24353,N_23741,N_23543);
nand U24354 (N_24354,N_23252,N_23629);
or U24355 (N_24355,N_23694,N_23388);
nand U24356 (N_24356,N_23354,N_23525);
and U24357 (N_24357,N_23266,N_23587);
and U24358 (N_24358,N_23135,N_23127);
nand U24359 (N_24359,N_23709,N_23680);
and U24360 (N_24360,N_23221,N_23222);
xnor U24361 (N_24361,N_23217,N_23143);
xor U24362 (N_24362,N_23432,N_23265);
and U24363 (N_24363,N_23560,N_23222);
nor U24364 (N_24364,N_23406,N_23433);
nor U24365 (N_24365,N_23604,N_23395);
nand U24366 (N_24366,N_23427,N_23569);
nor U24367 (N_24367,N_23347,N_23261);
and U24368 (N_24368,N_23413,N_23245);
nand U24369 (N_24369,N_23405,N_23496);
nor U24370 (N_24370,N_23275,N_23347);
xnor U24371 (N_24371,N_23179,N_23266);
or U24372 (N_24372,N_23511,N_23364);
nor U24373 (N_24373,N_23400,N_23208);
or U24374 (N_24374,N_23628,N_23281);
nand U24375 (N_24375,N_23762,N_24126);
nor U24376 (N_24376,N_23757,N_24035);
and U24377 (N_24377,N_24354,N_24303);
nor U24378 (N_24378,N_23928,N_23940);
nor U24379 (N_24379,N_23843,N_24249);
and U24380 (N_24380,N_24308,N_23759);
nand U24381 (N_24381,N_23805,N_23828);
or U24382 (N_24382,N_24369,N_24257);
or U24383 (N_24383,N_24025,N_24358);
nor U24384 (N_24384,N_24190,N_23989);
nor U24385 (N_24385,N_23827,N_24193);
and U24386 (N_24386,N_24020,N_23986);
or U24387 (N_24387,N_24058,N_24227);
and U24388 (N_24388,N_23778,N_23849);
nand U24389 (N_24389,N_23945,N_23900);
nor U24390 (N_24390,N_23995,N_23894);
nor U24391 (N_24391,N_23798,N_24317);
and U24392 (N_24392,N_24062,N_23887);
nor U24393 (N_24393,N_24066,N_23978);
or U24394 (N_24394,N_24269,N_24338);
nor U24395 (N_24395,N_24319,N_24228);
xor U24396 (N_24396,N_23876,N_23942);
or U24397 (N_24397,N_24294,N_24106);
xnor U24398 (N_24398,N_24001,N_23958);
or U24399 (N_24399,N_24263,N_23954);
or U24400 (N_24400,N_24359,N_24260);
nand U24401 (N_24401,N_23856,N_23803);
xnor U24402 (N_24402,N_24323,N_24324);
or U24403 (N_24403,N_23943,N_23907);
xor U24404 (N_24404,N_24095,N_24104);
xor U24405 (N_24405,N_23829,N_24156);
xor U24406 (N_24406,N_23835,N_23851);
nor U24407 (N_24407,N_24343,N_24159);
or U24408 (N_24408,N_23949,N_24117);
nor U24409 (N_24409,N_23922,N_24049);
xnor U24410 (N_24410,N_23775,N_24216);
xnor U24411 (N_24411,N_23796,N_24366);
or U24412 (N_24412,N_23818,N_24160);
nand U24413 (N_24413,N_24112,N_24231);
nor U24414 (N_24414,N_24026,N_24187);
and U24415 (N_24415,N_24230,N_24098);
or U24416 (N_24416,N_23853,N_24105);
and U24417 (N_24417,N_23842,N_24219);
nor U24418 (N_24418,N_24059,N_24166);
nand U24419 (N_24419,N_23788,N_24044);
or U24420 (N_24420,N_23938,N_24013);
nor U24421 (N_24421,N_23925,N_24347);
xnor U24422 (N_24422,N_23977,N_24270);
or U24423 (N_24423,N_24250,N_23831);
nand U24424 (N_24424,N_24128,N_24145);
and U24425 (N_24425,N_24329,N_24141);
nand U24426 (N_24426,N_24217,N_23812);
or U24427 (N_24427,N_24043,N_24364);
xnor U24428 (N_24428,N_24362,N_23869);
or U24429 (N_24429,N_23824,N_24248);
nor U24430 (N_24430,N_24088,N_24287);
xnor U24431 (N_24431,N_24351,N_24094);
and U24432 (N_24432,N_23927,N_23886);
xnor U24433 (N_24433,N_23839,N_23874);
xor U24434 (N_24434,N_23974,N_24307);
xor U24435 (N_24435,N_24348,N_24185);
nand U24436 (N_24436,N_23859,N_24169);
nor U24437 (N_24437,N_24284,N_24144);
nor U24438 (N_24438,N_23936,N_24125);
xor U24439 (N_24439,N_24337,N_23772);
xnor U24440 (N_24440,N_24073,N_23765);
xor U24441 (N_24441,N_23911,N_24111);
xor U24442 (N_24442,N_24071,N_23779);
xnor U24443 (N_24443,N_24291,N_24109);
xor U24444 (N_24444,N_24229,N_24283);
or U24445 (N_24445,N_23821,N_23959);
xor U24446 (N_24446,N_24309,N_23982);
nand U24447 (N_24447,N_24280,N_23797);
or U24448 (N_24448,N_23806,N_23916);
or U24449 (N_24449,N_24310,N_24300);
nor U24450 (N_24450,N_24076,N_23973);
or U24451 (N_24451,N_24130,N_24334);
and U24452 (N_24452,N_23955,N_23915);
nand U24453 (N_24453,N_24138,N_24012);
nor U24454 (N_24454,N_23926,N_24009);
and U24455 (N_24455,N_24246,N_23836);
and U24456 (N_24456,N_23763,N_23910);
or U24457 (N_24457,N_24197,N_24274);
xor U24458 (N_24458,N_24191,N_23820);
and U24459 (N_24459,N_23944,N_24149);
nor U24460 (N_24460,N_23850,N_23905);
nand U24461 (N_24461,N_23976,N_24242);
nor U24462 (N_24462,N_24202,N_23848);
or U24463 (N_24463,N_24153,N_24003);
nand U24464 (N_24464,N_23840,N_24245);
nand U24465 (N_24465,N_24275,N_23947);
xor U24466 (N_24466,N_24277,N_23979);
nand U24467 (N_24467,N_23847,N_24092);
xnor U24468 (N_24468,N_24355,N_23929);
xor U24469 (N_24469,N_24063,N_24306);
and U24470 (N_24470,N_23794,N_24154);
nand U24471 (N_24471,N_24080,N_24212);
nor U24472 (N_24472,N_24244,N_23787);
xnor U24473 (N_24473,N_24298,N_24083);
xor U24474 (N_24474,N_24093,N_23776);
xnor U24475 (N_24475,N_23879,N_24221);
nand U24476 (N_24476,N_23813,N_24137);
or U24477 (N_24477,N_24254,N_24040);
nor U24478 (N_24478,N_23902,N_24201);
or U24479 (N_24479,N_24206,N_24181);
nand U24480 (N_24480,N_24038,N_23953);
nand U24481 (N_24481,N_24215,N_24052);
or U24482 (N_24482,N_24016,N_24099);
or U24483 (N_24483,N_24171,N_23985);
nand U24484 (N_24484,N_23948,N_23823);
nand U24485 (N_24485,N_24042,N_24086);
nand U24486 (N_24486,N_24296,N_23987);
or U24487 (N_24487,N_23956,N_24142);
and U24488 (N_24488,N_24315,N_24139);
xnor U24489 (N_24489,N_24258,N_24252);
nor U24490 (N_24490,N_23923,N_24301);
xnor U24491 (N_24491,N_23819,N_24236);
nor U24492 (N_24492,N_23800,N_24295);
xnor U24493 (N_24493,N_23814,N_23845);
or U24494 (N_24494,N_24361,N_24061);
and U24495 (N_24495,N_23767,N_24007);
or U24496 (N_24496,N_24082,N_23862);
nand U24497 (N_24497,N_23785,N_24045);
and U24498 (N_24498,N_24259,N_24234);
and U24499 (N_24499,N_23766,N_24031);
nor U24500 (N_24500,N_24183,N_24365);
nor U24501 (N_24501,N_24178,N_24288);
xor U24502 (N_24502,N_23852,N_24176);
nor U24503 (N_24503,N_23918,N_24136);
xnor U24504 (N_24504,N_23770,N_23752);
or U24505 (N_24505,N_24021,N_24124);
nor U24506 (N_24506,N_24218,N_24024);
nor U24507 (N_24507,N_24240,N_23860);
and U24508 (N_24508,N_24180,N_24172);
nand U24509 (N_24509,N_24195,N_23793);
xnor U24510 (N_24510,N_24220,N_24091);
xor U24511 (N_24511,N_24339,N_24267);
and U24512 (N_24512,N_24325,N_23980);
nor U24513 (N_24513,N_23795,N_24004);
and U24514 (N_24514,N_24285,N_24194);
nand U24515 (N_24515,N_24320,N_23888);
and U24516 (N_24516,N_23931,N_23877);
nand U24517 (N_24517,N_24048,N_24133);
xor U24518 (N_24518,N_23833,N_23924);
xor U24519 (N_24519,N_24135,N_23826);
or U24520 (N_24520,N_24108,N_24037);
nor U24521 (N_24521,N_23875,N_23970);
nor U24522 (N_24522,N_24333,N_23846);
or U24523 (N_24523,N_23758,N_24030);
nor U24524 (N_24524,N_24344,N_24121);
and U24525 (N_24525,N_24034,N_23825);
nand U24526 (N_24526,N_24349,N_24293);
and U24527 (N_24527,N_24271,N_23904);
or U24528 (N_24528,N_24151,N_23967);
and U24529 (N_24529,N_23782,N_23975);
nand U24530 (N_24530,N_24078,N_24055);
nand U24531 (N_24531,N_24064,N_24018);
nor U24532 (N_24532,N_24162,N_23906);
xnor U24533 (N_24533,N_24345,N_23755);
nor U24534 (N_24534,N_24005,N_23961);
xnor U24535 (N_24535,N_24264,N_24170);
nor U24536 (N_24536,N_23921,N_24208);
nand U24537 (N_24537,N_23773,N_23939);
xnor U24538 (N_24538,N_23998,N_23802);
nand U24539 (N_24539,N_23783,N_24318);
and U24540 (N_24540,N_24158,N_23844);
xor U24541 (N_24541,N_24173,N_24367);
and U24542 (N_24542,N_24199,N_23996);
and U24543 (N_24543,N_23934,N_24281);
and U24544 (N_24544,N_24148,N_24286);
or U24545 (N_24545,N_24127,N_23932);
nand U24546 (N_24546,N_24265,N_23769);
nand U24547 (N_24547,N_23937,N_23774);
xor U24548 (N_24548,N_23901,N_24085);
nor U24549 (N_24549,N_23784,N_24205);
or U24550 (N_24550,N_24207,N_24165);
and U24551 (N_24551,N_24029,N_24168);
nand U24552 (N_24552,N_24213,N_24353);
xor U24553 (N_24553,N_24008,N_24243);
and U24554 (N_24554,N_23832,N_24074);
nor U24555 (N_24555,N_23790,N_24372);
nand U24556 (N_24556,N_24279,N_23863);
xor U24557 (N_24557,N_23801,N_23873);
and U24558 (N_24558,N_24262,N_24179);
or U24559 (N_24559,N_23789,N_24210);
nor U24560 (N_24560,N_23997,N_24247);
nand U24561 (N_24561,N_24273,N_24211);
and U24562 (N_24562,N_23861,N_24255);
and U24563 (N_24563,N_23838,N_24060);
or U24564 (N_24564,N_23891,N_24299);
or U24565 (N_24565,N_23753,N_24113);
and U24566 (N_24566,N_23913,N_24253);
xor U24567 (N_24567,N_24019,N_23809);
or U24568 (N_24568,N_24023,N_24328);
and U24569 (N_24569,N_24161,N_23754);
nand U24570 (N_24570,N_24235,N_24374);
nor U24571 (N_24571,N_23804,N_24090);
or U24572 (N_24572,N_23816,N_24278);
nand U24573 (N_24573,N_23807,N_23935);
xor U24574 (N_24574,N_24346,N_24047);
or U24575 (N_24575,N_24313,N_24330);
xnor U24576 (N_24576,N_24184,N_24041);
and U24577 (N_24577,N_23969,N_24373);
nand U24578 (N_24578,N_24110,N_23751);
nor U24579 (N_24579,N_24157,N_23893);
xor U24580 (N_24580,N_23992,N_24370);
and U24581 (N_24581,N_23768,N_24297);
nand U24582 (N_24582,N_23981,N_24341);
nor U24583 (N_24583,N_24120,N_24316);
nand U24584 (N_24584,N_24340,N_23882);
and U24585 (N_24585,N_24204,N_24140);
and U24586 (N_24586,N_23781,N_24084);
xor U24587 (N_24587,N_24302,N_24068);
and U24588 (N_24588,N_24174,N_24039);
and U24589 (N_24589,N_24056,N_24203);
nor U24590 (N_24590,N_23855,N_24336);
or U24591 (N_24591,N_24002,N_24036);
or U24592 (N_24592,N_24322,N_24118);
nand U24593 (N_24593,N_24053,N_24006);
xnor U24594 (N_24594,N_23750,N_23870);
or U24595 (N_24595,N_24356,N_24129);
nand U24596 (N_24596,N_23885,N_24057);
xnor U24597 (N_24597,N_24321,N_23858);
xnor U24598 (N_24598,N_24226,N_23971);
or U24599 (N_24599,N_24233,N_24352);
and U24600 (N_24600,N_23965,N_23898);
nor U24601 (N_24601,N_24272,N_24163);
xor U24602 (N_24602,N_24266,N_23792);
xor U24603 (N_24603,N_23960,N_24022);
or U24604 (N_24604,N_24268,N_24150);
and U24605 (N_24605,N_24225,N_23872);
and U24606 (N_24606,N_23993,N_24223);
nand U24607 (N_24607,N_23865,N_24103);
nand U24608 (N_24608,N_23822,N_23830);
nor U24609 (N_24609,N_23780,N_24000);
xnor U24610 (N_24610,N_24232,N_24311);
xnor U24611 (N_24611,N_24239,N_24011);
and U24612 (N_24612,N_24327,N_23881);
or U24613 (N_24613,N_24027,N_24331);
and U24614 (N_24614,N_24251,N_24182);
xnor U24615 (N_24615,N_23760,N_24175);
and U24616 (N_24616,N_24087,N_24065);
or U24617 (N_24617,N_23988,N_23817);
or U24618 (N_24618,N_23999,N_23880);
or U24619 (N_24619,N_23892,N_24081);
nor U24620 (N_24620,N_24050,N_24209);
or U24621 (N_24621,N_24115,N_23857);
or U24622 (N_24622,N_24368,N_24123);
or U24623 (N_24623,N_24069,N_24134);
nand U24624 (N_24624,N_24028,N_23867);
or U24625 (N_24625,N_23991,N_24100);
and U24626 (N_24626,N_24097,N_23764);
and U24627 (N_24627,N_24146,N_23899);
nand U24628 (N_24628,N_23962,N_24214);
nand U24629 (N_24629,N_24132,N_23903);
and U24630 (N_24630,N_24363,N_23799);
nor U24631 (N_24631,N_23878,N_23994);
xor U24632 (N_24632,N_24238,N_23854);
xor U24633 (N_24633,N_24152,N_24116);
or U24634 (N_24634,N_24014,N_23950);
nor U24635 (N_24635,N_23811,N_23941);
nand U24636 (N_24636,N_24304,N_24054);
xnor U24637 (N_24637,N_23864,N_23933);
nand U24638 (N_24638,N_23756,N_24342);
and U24639 (N_24639,N_23777,N_24102);
nor U24640 (N_24640,N_24350,N_24292);
xor U24641 (N_24641,N_23951,N_23815);
nand U24642 (N_24642,N_24282,N_23786);
or U24643 (N_24643,N_24017,N_24256);
and U24644 (N_24644,N_23966,N_24305);
nand U24645 (N_24645,N_24147,N_24155);
xnor U24646 (N_24646,N_23895,N_24261);
nand U24647 (N_24647,N_24032,N_24143);
xnor U24648 (N_24648,N_24312,N_23889);
xnor U24649 (N_24649,N_24290,N_24051);
nand U24650 (N_24650,N_24164,N_23791);
nand U24651 (N_24651,N_24276,N_24131);
nand U24652 (N_24652,N_23930,N_24077);
xnor U24653 (N_24653,N_24186,N_23912);
nand U24654 (N_24654,N_23761,N_24101);
nand U24655 (N_24655,N_23808,N_24075);
nand U24656 (N_24656,N_23952,N_23963);
nor U24657 (N_24657,N_24326,N_23964);
and U24658 (N_24658,N_23837,N_23897);
nand U24659 (N_24659,N_24196,N_24289);
nor U24660 (N_24660,N_24200,N_23841);
nor U24661 (N_24661,N_23909,N_24119);
xor U24662 (N_24662,N_24237,N_24241);
nand U24663 (N_24663,N_24371,N_24072);
or U24664 (N_24664,N_24357,N_23920);
xor U24665 (N_24665,N_24046,N_23990);
nand U24666 (N_24666,N_23866,N_24192);
and U24667 (N_24667,N_24096,N_23908);
and U24668 (N_24668,N_23834,N_23871);
nand U24669 (N_24669,N_24335,N_24114);
and U24670 (N_24670,N_23771,N_23946);
and U24671 (N_24671,N_23972,N_23896);
nor U24672 (N_24672,N_23883,N_24314);
nand U24673 (N_24673,N_24089,N_24015);
or U24674 (N_24674,N_23884,N_24010);
nor U24675 (N_24675,N_23917,N_24189);
nand U24676 (N_24676,N_23957,N_24360);
xor U24677 (N_24677,N_24070,N_24122);
and U24678 (N_24678,N_23968,N_24079);
nor U24679 (N_24679,N_24033,N_24188);
nor U24680 (N_24680,N_24067,N_23983);
nand U24681 (N_24681,N_23868,N_24107);
or U24682 (N_24682,N_23914,N_23890);
nand U24683 (N_24683,N_24167,N_24177);
xnor U24684 (N_24684,N_23919,N_24222);
nand U24685 (N_24685,N_23810,N_24332);
nand U24686 (N_24686,N_24224,N_24198);
or U24687 (N_24687,N_23984,N_24039);
and U24688 (N_24688,N_23869,N_23787);
or U24689 (N_24689,N_24235,N_24168);
or U24690 (N_24690,N_24028,N_24021);
nor U24691 (N_24691,N_23768,N_24124);
and U24692 (N_24692,N_23816,N_24012);
nand U24693 (N_24693,N_23898,N_23823);
xor U24694 (N_24694,N_23757,N_23855);
and U24695 (N_24695,N_23858,N_24222);
and U24696 (N_24696,N_24122,N_23787);
xnor U24697 (N_24697,N_23756,N_24268);
or U24698 (N_24698,N_23760,N_23994);
nand U24699 (N_24699,N_24311,N_24280);
and U24700 (N_24700,N_24172,N_23785);
and U24701 (N_24701,N_24291,N_24183);
nand U24702 (N_24702,N_24267,N_23902);
and U24703 (N_24703,N_23993,N_24110);
or U24704 (N_24704,N_24291,N_23868);
nand U24705 (N_24705,N_23778,N_23847);
nand U24706 (N_24706,N_24325,N_24138);
or U24707 (N_24707,N_23914,N_23808);
xnor U24708 (N_24708,N_24179,N_23956);
nand U24709 (N_24709,N_23763,N_23866);
nand U24710 (N_24710,N_24282,N_24041);
and U24711 (N_24711,N_23764,N_24357);
or U24712 (N_24712,N_24069,N_23831);
nor U24713 (N_24713,N_24024,N_24211);
or U24714 (N_24714,N_24319,N_24046);
or U24715 (N_24715,N_24246,N_24207);
nand U24716 (N_24716,N_24013,N_23959);
xor U24717 (N_24717,N_24238,N_24086);
and U24718 (N_24718,N_23899,N_24186);
nor U24719 (N_24719,N_23943,N_24250);
nand U24720 (N_24720,N_24292,N_24110);
nand U24721 (N_24721,N_24041,N_24129);
or U24722 (N_24722,N_23993,N_23888);
xor U24723 (N_24723,N_24371,N_24170);
nand U24724 (N_24724,N_24278,N_24359);
nand U24725 (N_24725,N_24213,N_24148);
xor U24726 (N_24726,N_24250,N_23880);
xor U24727 (N_24727,N_23973,N_24263);
or U24728 (N_24728,N_24016,N_24039);
and U24729 (N_24729,N_23857,N_23859);
xor U24730 (N_24730,N_24316,N_24336);
nor U24731 (N_24731,N_24270,N_24035);
nand U24732 (N_24732,N_24072,N_23762);
xnor U24733 (N_24733,N_23999,N_23871);
or U24734 (N_24734,N_23781,N_24353);
xor U24735 (N_24735,N_23890,N_24043);
nor U24736 (N_24736,N_24035,N_24078);
xor U24737 (N_24737,N_23956,N_23999);
or U24738 (N_24738,N_24299,N_23820);
xor U24739 (N_24739,N_23947,N_23907);
or U24740 (N_24740,N_23960,N_23903);
or U24741 (N_24741,N_23825,N_24286);
and U24742 (N_24742,N_24115,N_24153);
xor U24743 (N_24743,N_24007,N_23837);
nand U24744 (N_24744,N_24021,N_24284);
or U24745 (N_24745,N_23987,N_24162);
and U24746 (N_24746,N_24071,N_23804);
xnor U24747 (N_24747,N_24052,N_23896);
and U24748 (N_24748,N_23948,N_24297);
xnor U24749 (N_24749,N_24185,N_24190);
nand U24750 (N_24750,N_24202,N_23955);
or U24751 (N_24751,N_24210,N_23992);
nand U24752 (N_24752,N_23911,N_24147);
and U24753 (N_24753,N_23979,N_24293);
nand U24754 (N_24754,N_23940,N_24344);
and U24755 (N_24755,N_24145,N_23919);
nor U24756 (N_24756,N_23751,N_23980);
nor U24757 (N_24757,N_24025,N_24271);
nor U24758 (N_24758,N_24367,N_24366);
and U24759 (N_24759,N_24372,N_24040);
nor U24760 (N_24760,N_23954,N_23853);
nor U24761 (N_24761,N_24197,N_24061);
nand U24762 (N_24762,N_23890,N_24036);
xnor U24763 (N_24763,N_24315,N_23775);
or U24764 (N_24764,N_23868,N_24095);
nor U24765 (N_24765,N_23843,N_24263);
and U24766 (N_24766,N_24198,N_24276);
xor U24767 (N_24767,N_24174,N_23970);
and U24768 (N_24768,N_24180,N_23759);
or U24769 (N_24769,N_24230,N_24108);
xor U24770 (N_24770,N_23983,N_23773);
xnor U24771 (N_24771,N_24257,N_24072);
nor U24772 (N_24772,N_24156,N_24047);
nand U24773 (N_24773,N_23791,N_24233);
or U24774 (N_24774,N_24072,N_23823);
xnor U24775 (N_24775,N_23870,N_23932);
nor U24776 (N_24776,N_23972,N_23834);
xnor U24777 (N_24777,N_23780,N_23914);
or U24778 (N_24778,N_24187,N_23837);
and U24779 (N_24779,N_24023,N_24315);
xor U24780 (N_24780,N_23791,N_24041);
or U24781 (N_24781,N_24338,N_24030);
or U24782 (N_24782,N_24058,N_23952);
nor U24783 (N_24783,N_23972,N_23928);
xor U24784 (N_24784,N_24357,N_23892);
nand U24785 (N_24785,N_24045,N_24322);
nand U24786 (N_24786,N_24209,N_24255);
and U24787 (N_24787,N_24272,N_24210);
or U24788 (N_24788,N_24191,N_24022);
xor U24789 (N_24789,N_24232,N_23993);
or U24790 (N_24790,N_24069,N_24205);
nor U24791 (N_24791,N_24074,N_23805);
or U24792 (N_24792,N_23823,N_23902);
or U24793 (N_24793,N_23841,N_23883);
and U24794 (N_24794,N_24356,N_24122);
or U24795 (N_24795,N_23787,N_24360);
or U24796 (N_24796,N_23818,N_23872);
nor U24797 (N_24797,N_24021,N_24291);
or U24798 (N_24798,N_23843,N_24240);
and U24799 (N_24799,N_23944,N_23886);
xnor U24800 (N_24800,N_24190,N_23869);
xor U24801 (N_24801,N_24234,N_24216);
nor U24802 (N_24802,N_24175,N_24048);
nor U24803 (N_24803,N_24349,N_24087);
xor U24804 (N_24804,N_24252,N_24009);
xor U24805 (N_24805,N_23896,N_23948);
nor U24806 (N_24806,N_23916,N_23963);
nor U24807 (N_24807,N_24019,N_23763);
and U24808 (N_24808,N_24236,N_24116);
xor U24809 (N_24809,N_23930,N_24138);
xor U24810 (N_24810,N_24073,N_24060);
and U24811 (N_24811,N_24352,N_24018);
nand U24812 (N_24812,N_23852,N_24258);
nor U24813 (N_24813,N_24365,N_24096);
nand U24814 (N_24814,N_24235,N_23886);
nor U24815 (N_24815,N_23884,N_24007);
xor U24816 (N_24816,N_23932,N_23854);
or U24817 (N_24817,N_24262,N_24097);
and U24818 (N_24818,N_23868,N_23987);
nor U24819 (N_24819,N_24247,N_24210);
and U24820 (N_24820,N_24253,N_24296);
xnor U24821 (N_24821,N_24340,N_24059);
or U24822 (N_24822,N_24297,N_24050);
nor U24823 (N_24823,N_24290,N_23933);
xnor U24824 (N_24824,N_24166,N_23917);
xnor U24825 (N_24825,N_23846,N_23777);
or U24826 (N_24826,N_23979,N_24046);
xor U24827 (N_24827,N_24291,N_23859);
or U24828 (N_24828,N_23773,N_24055);
or U24829 (N_24829,N_24125,N_23770);
nand U24830 (N_24830,N_23876,N_24207);
or U24831 (N_24831,N_24007,N_24135);
or U24832 (N_24832,N_24240,N_24050);
or U24833 (N_24833,N_24071,N_24296);
xnor U24834 (N_24834,N_24324,N_23963);
xnor U24835 (N_24835,N_23927,N_24175);
or U24836 (N_24836,N_24078,N_24201);
nand U24837 (N_24837,N_23851,N_23979);
nor U24838 (N_24838,N_24299,N_24287);
nand U24839 (N_24839,N_24024,N_24268);
and U24840 (N_24840,N_23825,N_24009);
and U24841 (N_24841,N_24334,N_24326);
nand U24842 (N_24842,N_24329,N_23865);
nor U24843 (N_24843,N_23967,N_24148);
or U24844 (N_24844,N_23993,N_23957);
nor U24845 (N_24845,N_24292,N_24156);
nand U24846 (N_24846,N_24325,N_23756);
and U24847 (N_24847,N_24153,N_23789);
xnor U24848 (N_24848,N_24335,N_24077);
or U24849 (N_24849,N_24360,N_24141);
nand U24850 (N_24850,N_24234,N_23809);
nand U24851 (N_24851,N_24069,N_23755);
nand U24852 (N_24852,N_24373,N_24078);
or U24853 (N_24853,N_24274,N_24147);
xor U24854 (N_24854,N_23863,N_23973);
nand U24855 (N_24855,N_23778,N_24046);
xor U24856 (N_24856,N_24371,N_23813);
nand U24857 (N_24857,N_24050,N_24188);
or U24858 (N_24858,N_23773,N_24198);
nor U24859 (N_24859,N_23768,N_23857);
or U24860 (N_24860,N_24341,N_23808);
xor U24861 (N_24861,N_24296,N_24239);
nand U24862 (N_24862,N_24150,N_23814);
nand U24863 (N_24863,N_23816,N_24241);
xor U24864 (N_24864,N_24085,N_24034);
nand U24865 (N_24865,N_24118,N_24369);
or U24866 (N_24866,N_24057,N_24157);
or U24867 (N_24867,N_23820,N_23860);
nand U24868 (N_24868,N_24146,N_24229);
nor U24869 (N_24869,N_23963,N_24113);
nor U24870 (N_24870,N_24331,N_23806);
and U24871 (N_24871,N_24273,N_23945);
nand U24872 (N_24872,N_24337,N_23807);
nand U24873 (N_24873,N_23788,N_23902);
nor U24874 (N_24874,N_23881,N_24367);
nand U24875 (N_24875,N_23959,N_24124);
nand U24876 (N_24876,N_24052,N_24266);
nor U24877 (N_24877,N_23750,N_23992);
nand U24878 (N_24878,N_24151,N_23997);
nand U24879 (N_24879,N_24055,N_23778);
nand U24880 (N_24880,N_23915,N_23908);
nand U24881 (N_24881,N_24118,N_23960);
xnor U24882 (N_24882,N_23957,N_24156);
or U24883 (N_24883,N_24089,N_23871);
and U24884 (N_24884,N_23770,N_24039);
xor U24885 (N_24885,N_23889,N_24235);
nand U24886 (N_24886,N_24357,N_23778);
or U24887 (N_24887,N_24143,N_23765);
nand U24888 (N_24888,N_24023,N_23773);
or U24889 (N_24889,N_24246,N_24244);
nor U24890 (N_24890,N_24356,N_23846);
nand U24891 (N_24891,N_24308,N_23913);
nor U24892 (N_24892,N_23965,N_23809);
nor U24893 (N_24893,N_24328,N_23907);
nand U24894 (N_24894,N_24110,N_23932);
xnor U24895 (N_24895,N_24184,N_24267);
nand U24896 (N_24896,N_24108,N_23873);
and U24897 (N_24897,N_24180,N_24334);
nand U24898 (N_24898,N_23793,N_23889);
nand U24899 (N_24899,N_23805,N_24239);
and U24900 (N_24900,N_23853,N_24221);
nor U24901 (N_24901,N_24057,N_24238);
xnor U24902 (N_24902,N_23793,N_23958);
xor U24903 (N_24903,N_23883,N_24322);
xor U24904 (N_24904,N_24269,N_23855);
nand U24905 (N_24905,N_24079,N_24036);
or U24906 (N_24906,N_23896,N_24224);
nor U24907 (N_24907,N_23751,N_24065);
and U24908 (N_24908,N_23848,N_24038);
nand U24909 (N_24909,N_24180,N_23968);
nor U24910 (N_24910,N_23932,N_24199);
and U24911 (N_24911,N_23991,N_23839);
nand U24912 (N_24912,N_23901,N_23829);
or U24913 (N_24913,N_24289,N_23832);
nand U24914 (N_24914,N_24364,N_24306);
xnor U24915 (N_24915,N_24101,N_24184);
or U24916 (N_24916,N_24262,N_24195);
nand U24917 (N_24917,N_23913,N_23799);
nand U24918 (N_24918,N_24319,N_23856);
nor U24919 (N_24919,N_24308,N_24035);
and U24920 (N_24920,N_23784,N_23887);
and U24921 (N_24921,N_24093,N_24073);
xnor U24922 (N_24922,N_23846,N_24130);
nor U24923 (N_24923,N_23808,N_24364);
xnor U24924 (N_24924,N_24346,N_24348);
or U24925 (N_24925,N_24346,N_24041);
and U24926 (N_24926,N_24268,N_23841);
or U24927 (N_24927,N_24100,N_24313);
and U24928 (N_24928,N_23945,N_24222);
nor U24929 (N_24929,N_24091,N_24320);
xor U24930 (N_24930,N_23752,N_23818);
xnor U24931 (N_24931,N_24032,N_24228);
or U24932 (N_24932,N_24040,N_24320);
or U24933 (N_24933,N_23783,N_24309);
nor U24934 (N_24934,N_24226,N_23913);
nand U24935 (N_24935,N_23880,N_23881);
xnor U24936 (N_24936,N_23880,N_24227);
nand U24937 (N_24937,N_23963,N_23830);
and U24938 (N_24938,N_23792,N_24155);
or U24939 (N_24939,N_24056,N_23883);
nand U24940 (N_24940,N_23935,N_24179);
and U24941 (N_24941,N_24223,N_24111);
or U24942 (N_24942,N_24074,N_24148);
nand U24943 (N_24943,N_24230,N_23930);
nor U24944 (N_24944,N_23826,N_24084);
xor U24945 (N_24945,N_24305,N_23829);
or U24946 (N_24946,N_24276,N_23871);
or U24947 (N_24947,N_23819,N_24247);
nor U24948 (N_24948,N_23854,N_24168);
nor U24949 (N_24949,N_24103,N_24313);
xnor U24950 (N_24950,N_24200,N_24362);
or U24951 (N_24951,N_24107,N_24347);
xnor U24952 (N_24952,N_23787,N_23904);
nand U24953 (N_24953,N_23950,N_23891);
and U24954 (N_24954,N_24357,N_24251);
nor U24955 (N_24955,N_24341,N_23788);
and U24956 (N_24956,N_24159,N_24103);
nand U24957 (N_24957,N_23976,N_24112);
nor U24958 (N_24958,N_24136,N_24188);
nand U24959 (N_24959,N_24277,N_24275);
or U24960 (N_24960,N_23871,N_24184);
xnor U24961 (N_24961,N_23935,N_23879);
nand U24962 (N_24962,N_24344,N_24138);
or U24963 (N_24963,N_23780,N_23751);
nand U24964 (N_24964,N_24208,N_24166);
or U24965 (N_24965,N_24002,N_24272);
xor U24966 (N_24966,N_23869,N_24132);
xor U24967 (N_24967,N_24021,N_24157);
or U24968 (N_24968,N_23969,N_23919);
nand U24969 (N_24969,N_23968,N_23834);
nand U24970 (N_24970,N_23825,N_24020);
and U24971 (N_24971,N_24096,N_24321);
or U24972 (N_24972,N_24287,N_24335);
xnor U24973 (N_24973,N_24247,N_24061);
nor U24974 (N_24974,N_23879,N_23989);
or U24975 (N_24975,N_24268,N_23843);
nand U24976 (N_24976,N_24237,N_23997);
nand U24977 (N_24977,N_24124,N_24367);
and U24978 (N_24978,N_23963,N_24170);
and U24979 (N_24979,N_23792,N_24160);
nand U24980 (N_24980,N_23818,N_23829);
or U24981 (N_24981,N_24087,N_24078);
or U24982 (N_24982,N_24067,N_23922);
and U24983 (N_24983,N_24139,N_24205);
nand U24984 (N_24984,N_23812,N_24309);
and U24985 (N_24985,N_24023,N_24254);
or U24986 (N_24986,N_23887,N_24129);
nand U24987 (N_24987,N_23896,N_23783);
xor U24988 (N_24988,N_23973,N_23877);
nand U24989 (N_24989,N_23816,N_24191);
and U24990 (N_24990,N_24074,N_24257);
nand U24991 (N_24991,N_23798,N_23776);
nor U24992 (N_24992,N_23936,N_24137);
nor U24993 (N_24993,N_24074,N_24012);
nor U24994 (N_24994,N_24310,N_23816);
nand U24995 (N_24995,N_24244,N_23942);
nand U24996 (N_24996,N_23860,N_24041);
or U24997 (N_24997,N_23760,N_24126);
xnor U24998 (N_24998,N_23938,N_24103);
nand U24999 (N_24999,N_24166,N_24049);
nand UO_0 (O_0,N_24507,N_24913);
nor UO_1 (O_1,N_24720,N_24460);
nand UO_2 (O_2,N_24597,N_24682);
xor UO_3 (O_3,N_24877,N_24830);
and UO_4 (O_4,N_24499,N_24896);
xor UO_5 (O_5,N_24490,N_24807);
xnor UO_6 (O_6,N_24378,N_24848);
and UO_7 (O_7,N_24817,N_24582);
nor UO_8 (O_8,N_24448,N_24738);
nor UO_9 (O_9,N_24822,N_24764);
xor UO_10 (O_10,N_24850,N_24483);
nor UO_11 (O_11,N_24418,N_24867);
nor UO_12 (O_12,N_24730,N_24561);
nand UO_13 (O_13,N_24481,N_24417);
xor UO_14 (O_14,N_24668,N_24611);
and UO_15 (O_15,N_24821,N_24878);
xor UO_16 (O_16,N_24925,N_24853);
xnor UO_17 (O_17,N_24773,N_24622);
or UO_18 (O_18,N_24672,N_24991);
nor UO_19 (O_19,N_24526,N_24472);
xnor UO_20 (O_20,N_24737,N_24780);
xnor UO_21 (O_21,N_24843,N_24596);
nor UO_22 (O_22,N_24884,N_24916);
nand UO_23 (O_23,N_24735,N_24661);
xnor UO_24 (O_24,N_24944,N_24971);
nand UO_25 (O_25,N_24576,N_24524);
and UO_26 (O_26,N_24439,N_24427);
xor UO_27 (O_27,N_24808,N_24694);
xor UO_28 (O_28,N_24686,N_24643);
nor UO_29 (O_29,N_24533,N_24412);
and UO_30 (O_30,N_24401,N_24774);
xnor UO_31 (O_31,N_24458,N_24678);
or UO_32 (O_32,N_24468,N_24651);
xor UO_33 (O_33,N_24411,N_24710);
xor UO_34 (O_34,N_24933,N_24477);
nor UO_35 (O_35,N_24690,N_24794);
nor UO_36 (O_36,N_24656,N_24939);
or UO_37 (O_37,N_24566,N_24380);
or UO_38 (O_38,N_24441,N_24654);
nor UO_39 (O_39,N_24713,N_24508);
nor UO_40 (O_40,N_24506,N_24459);
and UO_41 (O_41,N_24389,N_24619);
and UO_42 (O_42,N_24658,N_24819);
nor UO_43 (O_43,N_24581,N_24791);
xor UO_44 (O_44,N_24856,N_24861);
xor UO_45 (O_45,N_24544,N_24482);
xor UO_46 (O_46,N_24930,N_24503);
nand UO_47 (O_47,N_24457,N_24613);
nand UO_48 (O_48,N_24492,N_24731);
xor UO_49 (O_49,N_24766,N_24521);
and UO_50 (O_50,N_24946,N_24631);
nor UO_51 (O_51,N_24430,N_24859);
and UO_52 (O_52,N_24601,N_24692);
or UO_53 (O_53,N_24719,N_24886);
and UO_54 (O_54,N_24625,N_24624);
nand UO_55 (O_55,N_24531,N_24956);
nor UO_56 (O_56,N_24724,N_24741);
xnor UO_57 (O_57,N_24620,N_24865);
nand UO_58 (O_58,N_24762,N_24558);
nor UO_59 (O_59,N_24899,N_24381);
or UO_60 (O_60,N_24437,N_24704);
nor UO_61 (O_61,N_24447,N_24465);
and UO_62 (O_62,N_24960,N_24665);
xnor UO_63 (O_63,N_24897,N_24422);
xor UO_64 (O_64,N_24759,N_24801);
or UO_65 (O_65,N_24924,N_24876);
or UO_66 (O_66,N_24679,N_24997);
or UO_67 (O_67,N_24723,N_24464);
nand UO_68 (O_68,N_24749,N_24627);
or UO_69 (O_69,N_24926,N_24758);
nand UO_70 (O_70,N_24927,N_24813);
and UO_71 (O_71,N_24747,N_24823);
nand UO_72 (O_72,N_24442,N_24902);
or UO_73 (O_73,N_24510,N_24868);
nor UO_74 (O_74,N_24384,N_24825);
nor UO_75 (O_75,N_24776,N_24645);
or UO_76 (O_76,N_24862,N_24547);
and UO_77 (O_77,N_24891,N_24502);
xor UO_78 (O_78,N_24768,N_24603);
nand UO_79 (O_79,N_24540,N_24388);
nor UO_80 (O_80,N_24838,N_24961);
nand UO_81 (O_81,N_24727,N_24739);
nand UO_82 (O_82,N_24449,N_24847);
nand UO_83 (O_83,N_24845,N_24573);
and UO_84 (O_84,N_24528,N_24443);
and UO_85 (O_85,N_24541,N_24874);
and UO_86 (O_86,N_24479,N_24901);
or UO_87 (O_87,N_24785,N_24792);
nand UO_88 (O_88,N_24833,N_24889);
nand UO_89 (O_89,N_24387,N_24428);
or UO_90 (O_90,N_24728,N_24685);
nor UO_91 (O_91,N_24599,N_24957);
or UO_92 (O_92,N_24455,N_24438);
or UO_93 (O_93,N_24935,N_24466);
nor UO_94 (O_94,N_24734,N_24446);
and UO_95 (O_95,N_24977,N_24397);
nand UO_96 (O_96,N_24501,N_24638);
nor UO_97 (O_97,N_24688,N_24700);
or UO_98 (O_98,N_24907,N_24662);
and UO_99 (O_99,N_24639,N_24765);
xor UO_100 (O_100,N_24952,N_24980);
nand UO_101 (O_101,N_24753,N_24669);
xnor UO_102 (O_102,N_24659,N_24636);
nor UO_103 (O_103,N_24904,N_24424);
and UO_104 (O_104,N_24574,N_24615);
nor UO_105 (O_105,N_24937,N_24549);
xor UO_106 (O_106,N_24403,N_24851);
and UO_107 (O_107,N_24379,N_24992);
xnor UO_108 (O_108,N_24725,N_24606);
xor UO_109 (O_109,N_24872,N_24905);
and UO_110 (O_110,N_24664,N_24707);
and UO_111 (O_111,N_24751,N_24382);
and UO_112 (O_112,N_24979,N_24536);
nand UO_113 (O_113,N_24909,N_24721);
nand UO_114 (O_114,N_24908,N_24898);
nand UO_115 (O_115,N_24820,N_24425);
nand UO_116 (O_116,N_24718,N_24607);
or UO_117 (O_117,N_24475,N_24949);
nand UO_118 (O_118,N_24929,N_24605);
xnor UO_119 (O_119,N_24628,N_24947);
nand UO_120 (O_120,N_24551,N_24932);
and UO_121 (O_121,N_24858,N_24534);
nand UO_122 (O_122,N_24855,N_24965);
nor UO_123 (O_123,N_24511,N_24667);
xnor UO_124 (O_124,N_24955,N_24696);
and UO_125 (O_125,N_24588,N_24630);
nor UO_126 (O_126,N_24978,N_24885);
nand UO_127 (O_127,N_24405,N_24670);
nor UO_128 (O_128,N_24637,N_24635);
nor UO_129 (O_129,N_24648,N_24419);
and UO_130 (O_130,N_24553,N_24777);
nand UO_131 (O_131,N_24921,N_24461);
xnor UO_132 (O_132,N_24911,N_24647);
and UO_133 (O_133,N_24910,N_24711);
and UO_134 (O_134,N_24831,N_24386);
and UO_135 (O_135,N_24612,N_24954);
nor UO_136 (O_136,N_24772,N_24600);
or UO_137 (O_137,N_24890,N_24784);
nand UO_138 (O_138,N_24879,N_24476);
nor UO_139 (O_139,N_24839,N_24660);
and UO_140 (O_140,N_24532,N_24832);
nor UO_141 (O_141,N_24462,N_24915);
and UO_142 (O_142,N_24812,N_24585);
nand UO_143 (O_143,N_24505,N_24809);
xnor UO_144 (O_144,N_24591,N_24618);
nor UO_145 (O_145,N_24577,N_24959);
nand UO_146 (O_146,N_24967,N_24568);
xor UO_147 (O_147,N_24999,N_24775);
xnor UO_148 (O_148,N_24706,N_24485);
nor UO_149 (O_149,N_24496,N_24673);
xor UO_150 (O_150,N_24882,N_24746);
and UO_151 (O_151,N_24409,N_24840);
nand UO_152 (O_152,N_24798,N_24486);
nand UO_153 (O_153,N_24474,N_24681);
or UO_154 (O_154,N_24683,N_24402);
or UO_155 (O_155,N_24860,N_24870);
nand UO_156 (O_156,N_24875,N_24557);
and UO_157 (O_157,N_24626,N_24836);
or UO_158 (O_158,N_24488,N_24828);
nand UO_159 (O_159,N_24844,N_24396);
nand UO_160 (O_160,N_24974,N_24796);
nand UO_161 (O_161,N_24849,N_24883);
xnor UO_162 (O_162,N_24752,N_24827);
and UO_163 (O_163,N_24560,N_24671);
nor UO_164 (O_164,N_24988,N_24985);
nor UO_165 (O_165,N_24604,N_24608);
or UO_166 (O_166,N_24399,N_24571);
or UO_167 (O_167,N_24783,N_24824);
xor UO_168 (O_168,N_24590,N_24699);
nand UO_169 (O_169,N_24575,N_24495);
xor UO_170 (O_170,N_24803,N_24770);
nand UO_171 (O_171,N_24994,N_24516);
nand UO_172 (O_172,N_24757,N_24513);
or UO_173 (O_173,N_24938,N_24787);
nand UO_174 (O_174,N_24489,N_24674);
or UO_175 (O_175,N_24703,N_24716);
and UO_176 (O_176,N_24609,N_24680);
xor UO_177 (O_177,N_24518,N_24816);
and UO_178 (O_178,N_24778,N_24953);
nor UO_179 (O_179,N_24923,N_24733);
or UO_180 (O_180,N_24701,N_24852);
and UO_181 (O_181,N_24987,N_24454);
nand UO_182 (O_182,N_24846,N_24546);
nand UO_183 (O_183,N_24640,N_24708);
or UO_184 (O_184,N_24826,N_24487);
or UO_185 (O_185,N_24842,N_24854);
nor UO_186 (O_186,N_24951,N_24771);
and UO_187 (O_187,N_24788,N_24527);
and UO_188 (O_188,N_24722,N_24407);
nor UO_189 (O_189,N_24395,N_24385);
and UO_190 (O_190,N_24769,N_24709);
xor UO_191 (O_191,N_24408,N_24400);
nand UO_192 (O_192,N_24726,N_24912);
and UO_193 (O_193,N_24548,N_24941);
nand UO_194 (O_194,N_24383,N_24542);
xor UO_195 (O_195,N_24413,N_24423);
or UO_196 (O_196,N_24687,N_24434);
nand UO_197 (O_197,N_24964,N_24969);
or UO_198 (O_198,N_24864,N_24748);
nor UO_199 (O_199,N_24750,N_24790);
xnor UO_200 (O_200,N_24406,N_24984);
nand UO_201 (O_201,N_24653,N_24881);
xnor UO_202 (O_202,N_24806,N_24520);
nor UO_203 (O_203,N_24632,N_24426);
nand UO_204 (O_204,N_24989,N_24983);
and UO_205 (O_205,N_24958,N_24435);
nor UO_206 (O_206,N_24761,N_24471);
xnor UO_207 (O_207,N_24415,N_24456);
xor UO_208 (O_208,N_24550,N_24610);
and UO_209 (O_209,N_24922,N_24444);
nor UO_210 (O_210,N_24779,N_24975);
nand UO_211 (O_211,N_24641,N_24970);
or UO_212 (O_212,N_24990,N_24579);
xor UO_213 (O_213,N_24500,N_24452);
xnor UO_214 (O_214,N_24391,N_24837);
and UO_215 (O_215,N_24940,N_24982);
or UO_216 (O_216,N_24906,N_24567);
xor UO_217 (O_217,N_24973,N_24517);
and UO_218 (O_218,N_24918,N_24410);
and UO_219 (O_219,N_24655,N_24740);
xnor UO_220 (O_220,N_24804,N_24789);
and UO_221 (O_221,N_24436,N_24377);
or UO_222 (O_222,N_24375,N_24556);
and UO_223 (O_223,N_24420,N_24811);
xnor UO_224 (O_224,N_24931,N_24697);
xor UO_225 (O_225,N_24497,N_24934);
or UO_226 (O_226,N_24594,N_24782);
nor UO_227 (O_227,N_24586,N_24565);
nor UO_228 (O_228,N_24966,N_24433);
nand UO_229 (O_229,N_24756,N_24440);
and UO_230 (O_230,N_24504,N_24943);
nand UO_231 (O_231,N_24512,N_24835);
or UO_232 (O_232,N_24621,N_24689);
xor UO_233 (O_233,N_24691,N_24545);
or UO_234 (O_234,N_24469,N_24416);
nand UO_235 (O_235,N_24445,N_24800);
or UO_236 (O_236,N_24525,N_24972);
or UO_237 (O_237,N_24572,N_24614);
nor UO_238 (O_238,N_24755,N_24888);
nand UO_239 (O_239,N_24453,N_24702);
nor UO_240 (O_240,N_24592,N_24633);
nand UO_241 (O_241,N_24563,N_24996);
and UO_242 (O_242,N_24616,N_24394);
or UO_243 (O_243,N_24543,N_24584);
and UO_244 (O_244,N_24494,N_24666);
xor UO_245 (O_245,N_24871,N_24863);
xor UO_246 (O_246,N_24745,N_24698);
nand UO_247 (O_247,N_24578,N_24484);
nor UO_248 (O_248,N_24432,N_24519);
nand UO_249 (O_249,N_24535,N_24392);
nor UO_250 (O_250,N_24623,N_24981);
or UO_251 (O_251,N_24644,N_24805);
nand UO_252 (O_252,N_24900,N_24583);
nand UO_253 (O_253,N_24602,N_24450);
nand UO_254 (O_254,N_24936,N_24451);
xnor UO_255 (O_255,N_24552,N_24393);
nand UO_256 (O_256,N_24398,N_24580);
and UO_257 (O_257,N_24652,N_24559);
and UO_258 (O_258,N_24754,N_24522);
nor UO_259 (O_259,N_24514,N_24463);
and UO_260 (O_260,N_24986,N_24799);
nor UO_261 (O_261,N_24646,N_24657);
nor UO_262 (O_262,N_24928,N_24887);
and UO_263 (O_263,N_24917,N_24993);
xnor UO_264 (O_264,N_24642,N_24467);
nand UO_265 (O_265,N_24570,N_24963);
xor UO_266 (O_266,N_24793,N_24431);
and UO_267 (O_267,N_24742,N_24480);
or UO_268 (O_268,N_24914,N_24714);
nor UO_269 (O_269,N_24473,N_24950);
or UO_270 (O_270,N_24523,N_24795);
nand UO_271 (O_271,N_24675,N_24797);
and UO_272 (O_272,N_24732,N_24919);
nor UO_273 (O_273,N_24598,N_24478);
xor UO_274 (O_274,N_24509,N_24744);
xnor UO_275 (O_275,N_24873,N_24593);
nand UO_276 (O_276,N_24695,N_24802);
nand UO_277 (O_277,N_24515,N_24529);
xnor UO_278 (O_278,N_24995,N_24895);
nor UO_279 (O_279,N_24537,N_24945);
or UO_280 (O_280,N_24866,N_24491);
and UO_281 (O_281,N_24903,N_24760);
and UO_282 (O_282,N_24893,N_24892);
nor UO_283 (O_283,N_24555,N_24715);
nor UO_284 (O_284,N_24650,N_24693);
nand UO_285 (O_285,N_24470,N_24763);
xnor UO_286 (O_286,N_24538,N_24841);
nor UO_287 (O_287,N_24493,N_24429);
nor UO_288 (O_288,N_24976,N_24818);
xor UO_289 (O_289,N_24564,N_24869);
or UO_290 (O_290,N_24498,N_24729);
nor UO_291 (O_291,N_24634,N_24810);
or UO_292 (O_292,N_24962,N_24530);
or UO_293 (O_293,N_24376,N_24649);
nand UO_294 (O_294,N_24421,N_24414);
nand UO_295 (O_295,N_24562,N_24677);
and UO_296 (O_296,N_24717,N_24595);
and UO_297 (O_297,N_24587,N_24894);
xor UO_298 (O_298,N_24781,N_24998);
and UO_299 (O_299,N_24589,N_24712);
and UO_300 (O_300,N_24880,N_24736);
or UO_301 (O_301,N_24815,N_24920);
nor UO_302 (O_302,N_24834,N_24539);
nand UO_303 (O_303,N_24857,N_24948);
nand UO_304 (O_304,N_24404,N_24968);
and UO_305 (O_305,N_24829,N_24554);
nor UO_306 (O_306,N_24743,N_24569);
or UO_307 (O_307,N_24786,N_24684);
xnor UO_308 (O_308,N_24676,N_24767);
nor UO_309 (O_309,N_24663,N_24390);
nor UO_310 (O_310,N_24617,N_24705);
nor UO_311 (O_311,N_24814,N_24942);
nand UO_312 (O_312,N_24629,N_24657);
and UO_313 (O_313,N_24413,N_24706);
nand UO_314 (O_314,N_24716,N_24572);
or UO_315 (O_315,N_24481,N_24595);
and UO_316 (O_316,N_24783,N_24741);
nor UO_317 (O_317,N_24400,N_24757);
nand UO_318 (O_318,N_24797,N_24409);
xor UO_319 (O_319,N_24687,N_24582);
xnor UO_320 (O_320,N_24500,N_24922);
xnor UO_321 (O_321,N_24662,N_24637);
nand UO_322 (O_322,N_24824,N_24660);
or UO_323 (O_323,N_24831,N_24956);
and UO_324 (O_324,N_24705,N_24919);
or UO_325 (O_325,N_24714,N_24611);
and UO_326 (O_326,N_24720,N_24942);
xor UO_327 (O_327,N_24583,N_24590);
or UO_328 (O_328,N_24736,N_24760);
nand UO_329 (O_329,N_24856,N_24690);
nand UO_330 (O_330,N_24834,N_24998);
and UO_331 (O_331,N_24390,N_24513);
or UO_332 (O_332,N_24918,N_24967);
nand UO_333 (O_333,N_24846,N_24947);
nor UO_334 (O_334,N_24665,N_24486);
and UO_335 (O_335,N_24864,N_24646);
nand UO_336 (O_336,N_24403,N_24638);
and UO_337 (O_337,N_24722,N_24505);
nor UO_338 (O_338,N_24610,N_24828);
nand UO_339 (O_339,N_24439,N_24705);
or UO_340 (O_340,N_24849,N_24786);
or UO_341 (O_341,N_24410,N_24897);
nand UO_342 (O_342,N_24427,N_24636);
nor UO_343 (O_343,N_24669,N_24670);
xor UO_344 (O_344,N_24773,N_24617);
or UO_345 (O_345,N_24634,N_24464);
nand UO_346 (O_346,N_24407,N_24554);
nand UO_347 (O_347,N_24773,N_24493);
nor UO_348 (O_348,N_24846,N_24435);
nand UO_349 (O_349,N_24749,N_24476);
nand UO_350 (O_350,N_24789,N_24429);
nand UO_351 (O_351,N_24683,N_24413);
and UO_352 (O_352,N_24871,N_24458);
and UO_353 (O_353,N_24885,N_24800);
or UO_354 (O_354,N_24549,N_24990);
nand UO_355 (O_355,N_24872,N_24459);
or UO_356 (O_356,N_24799,N_24955);
xor UO_357 (O_357,N_24411,N_24726);
and UO_358 (O_358,N_24965,N_24801);
or UO_359 (O_359,N_24666,N_24944);
nor UO_360 (O_360,N_24943,N_24503);
xor UO_361 (O_361,N_24860,N_24437);
nor UO_362 (O_362,N_24531,N_24472);
nand UO_363 (O_363,N_24822,N_24426);
and UO_364 (O_364,N_24527,N_24757);
nand UO_365 (O_365,N_24482,N_24993);
xnor UO_366 (O_366,N_24945,N_24450);
and UO_367 (O_367,N_24929,N_24905);
nand UO_368 (O_368,N_24949,N_24509);
nor UO_369 (O_369,N_24732,N_24687);
nand UO_370 (O_370,N_24600,N_24912);
or UO_371 (O_371,N_24442,N_24649);
xnor UO_372 (O_372,N_24642,N_24593);
xor UO_373 (O_373,N_24939,N_24415);
nor UO_374 (O_374,N_24722,N_24405);
nand UO_375 (O_375,N_24440,N_24802);
xor UO_376 (O_376,N_24796,N_24822);
nand UO_377 (O_377,N_24964,N_24688);
xnor UO_378 (O_378,N_24599,N_24567);
nand UO_379 (O_379,N_24689,N_24618);
xor UO_380 (O_380,N_24966,N_24789);
or UO_381 (O_381,N_24636,N_24918);
nand UO_382 (O_382,N_24716,N_24442);
nor UO_383 (O_383,N_24460,N_24758);
or UO_384 (O_384,N_24748,N_24568);
or UO_385 (O_385,N_24844,N_24879);
nor UO_386 (O_386,N_24750,N_24967);
and UO_387 (O_387,N_24481,N_24979);
nand UO_388 (O_388,N_24975,N_24715);
or UO_389 (O_389,N_24671,N_24596);
and UO_390 (O_390,N_24927,N_24942);
or UO_391 (O_391,N_24906,N_24457);
xor UO_392 (O_392,N_24759,N_24836);
xnor UO_393 (O_393,N_24720,N_24953);
xor UO_394 (O_394,N_24651,N_24618);
nor UO_395 (O_395,N_24407,N_24475);
and UO_396 (O_396,N_24436,N_24967);
and UO_397 (O_397,N_24483,N_24389);
and UO_398 (O_398,N_24625,N_24465);
nor UO_399 (O_399,N_24382,N_24744);
nand UO_400 (O_400,N_24404,N_24640);
and UO_401 (O_401,N_24510,N_24462);
nor UO_402 (O_402,N_24766,N_24406);
or UO_403 (O_403,N_24853,N_24680);
nor UO_404 (O_404,N_24885,N_24943);
or UO_405 (O_405,N_24816,N_24385);
nor UO_406 (O_406,N_24531,N_24647);
and UO_407 (O_407,N_24551,N_24404);
nand UO_408 (O_408,N_24757,N_24478);
nor UO_409 (O_409,N_24650,N_24797);
or UO_410 (O_410,N_24828,N_24534);
nand UO_411 (O_411,N_24809,N_24476);
and UO_412 (O_412,N_24563,N_24580);
nand UO_413 (O_413,N_24443,N_24642);
or UO_414 (O_414,N_24728,N_24701);
nand UO_415 (O_415,N_24418,N_24551);
and UO_416 (O_416,N_24556,N_24934);
and UO_417 (O_417,N_24493,N_24911);
nor UO_418 (O_418,N_24729,N_24637);
and UO_419 (O_419,N_24857,N_24886);
and UO_420 (O_420,N_24859,N_24700);
xnor UO_421 (O_421,N_24426,N_24470);
nor UO_422 (O_422,N_24618,N_24553);
and UO_423 (O_423,N_24650,N_24992);
xor UO_424 (O_424,N_24448,N_24381);
nand UO_425 (O_425,N_24695,N_24803);
nand UO_426 (O_426,N_24715,N_24560);
nor UO_427 (O_427,N_24891,N_24814);
and UO_428 (O_428,N_24842,N_24626);
nor UO_429 (O_429,N_24791,N_24835);
and UO_430 (O_430,N_24507,N_24595);
or UO_431 (O_431,N_24859,N_24997);
nand UO_432 (O_432,N_24579,N_24979);
xor UO_433 (O_433,N_24618,N_24596);
xor UO_434 (O_434,N_24731,N_24460);
nand UO_435 (O_435,N_24691,N_24454);
nand UO_436 (O_436,N_24842,N_24944);
xor UO_437 (O_437,N_24708,N_24988);
xor UO_438 (O_438,N_24796,N_24394);
nor UO_439 (O_439,N_24782,N_24801);
xnor UO_440 (O_440,N_24944,N_24425);
and UO_441 (O_441,N_24554,N_24861);
nand UO_442 (O_442,N_24846,N_24560);
xor UO_443 (O_443,N_24646,N_24865);
xor UO_444 (O_444,N_24678,N_24882);
and UO_445 (O_445,N_24872,N_24957);
nor UO_446 (O_446,N_24696,N_24417);
xor UO_447 (O_447,N_24793,N_24972);
and UO_448 (O_448,N_24443,N_24865);
or UO_449 (O_449,N_24493,N_24974);
xor UO_450 (O_450,N_24733,N_24435);
nor UO_451 (O_451,N_24418,N_24498);
nand UO_452 (O_452,N_24949,N_24492);
nor UO_453 (O_453,N_24762,N_24948);
nor UO_454 (O_454,N_24568,N_24727);
and UO_455 (O_455,N_24438,N_24609);
and UO_456 (O_456,N_24533,N_24788);
nor UO_457 (O_457,N_24821,N_24443);
and UO_458 (O_458,N_24669,N_24892);
or UO_459 (O_459,N_24670,N_24406);
nor UO_460 (O_460,N_24485,N_24890);
nand UO_461 (O_461,N_24985,N_24840);
xor UO_462 (O_462,N_24471,N_24825);
and UO_463 (O_463,N_24523,N_24639);
or UO_464 (O_464,N_24750,N_24661);
or UO_465 (O_465,N_24806,N_24845);
nand UO_466 (O_466,N_24754,N_24740);
nor UO_467 (O_467,N_24817,N_24981);
and UO_468 (O_468,N_24509,N_24755);
or UO_469 (O_469,N_24845,N_24914);
xor UO_470 (O_470,N_24736,N_24948);
and UO_471 (O_471,N_24850,N_24689);
and UO_472 (O_472,N_24954,N_24468);
nand UO_473 (O_473,N_24513,N_24900);
and UO_474 (O_474,N_24912,N_24993);
and UO_475 (O_475,N_24792,N_24509);
nor UO_476 (O_476,N_24960,N_24485);
nand UO_477 (O_477,N_24915,N_24429);
or UO_478 (O_478,N_24831,N_24597);
or UO_479 (O_479,N_24552,N_24937);
or UO_480 (O_480,N_24894,N_24476);
xnor UO_481 (O_481,N_24599,N_24638);
nor UO_482 (O_482,N_24509,N_24647);
or UO_483 (O_483,N_24687,N_24833);
or UO_484 (O_484,N_24839,N_24403);
nand UO_485 (O_485,N_24427,N_24703);
or UO_486 (O_486,N_24646,N_24952);
nor UO_487 (O_487,N_24898,N_24623);
and UO_488 (O_488,N_24867,N_24624);
nor UO_489 (O_489,N_24806,N_24890);
or UO_490 (O_490,N_24623,N_24924);
nand UO_491 (O_491,N_24379,N_24723);
or UO_492 (O_492,N_24832,N_24473);
or UO_493 (O_493,N_24853,N_24917);
nand UO_494 (O_494,N_24613,N_24637);
xnor UO_495 (O_495,N_24596,N_24954);
nand UO_496 (O_496,N_24724,N_24691);
xor UO_497 (O_497,N_24994,N_24979);
and UO_498 (O_498,N_24994,N_24426);
or UO_499 (O_499,N_24453,N_24828);
and UO_500 (O_500,N_24743,N_24880);
nor UO_501 (O_501,N_24902,N_24716);
nand UO_502 (O_502,N_24874,N_24458);
nand UO_503 (O_503,N_24634,N_24585);
or UO_504 (O_504,N_24416,N_24572);
xnor UO_505 (O_505,N_24921,N_24420);
and UO_506 (O_506,N_24441,N_24920);
nand UO_507 (O_507,N_24499,N_24952);
nor UO_508 (O_508,N_24473,N_24535);
nor UO_509 (O_509,N_24711,N_24792);
nor UO_510 (O_510,N_24678,N_24643);
nor UO_511 (O_511,N_24560,N_24645);
xnor UO_512 (O_512,N_24919,N_24382);
nor UO_513 (O_513,N_24797,N_24906);
xor UO_514 (O_514,N_24538,N_24640);
xnor UO_515 (O_515,N_24569,N_24588);
nor UO_516 (O_516,N_24820,N_24872);
xor UO_517 (O_517,N_24429,N_24688);
nor UO_518 (O_518,N_24627,N_24597);
or UO_519 (O_519,N_24846,N_24662);
or UO_520 (O_520,N_24756,N_24488);
and UO_521 (O_521,N_24928,N_24451);
nor UO_522 (O_522,N_24888,N_24393);
nand UO_523 (O_523,N_24421,N_24631);
xor UO_524 (O_524,N_24470,N_24852);
and UO_525 (O_525,N_24584,N_24525);
xor UO_526 (O_526,N_24395,N_24477);
xor UO_527 (O_527,N_24796,N_24860);
nand UO_528 (O_528,N_24620,N_24627);
nor UO_529 (O_529,N_24709,N_24932);
xnor UO_530 (O_530,N_24564,N_24865);
nor UO_531 (O_531,N_24471,N_24697);
or UO_532 (O_532,N_24505,N_24743);
xnor UO_533 (O_533,N_24431,N_24427);
and UO_534 (O_534,N_24632,N_24564);
nor UO_535 (O_535,N_24729,N_24560);
xnor UO_536 (O_536,N_24929,N_24402);
nor UO_537 (O_537,N_24721,N_24419);
xor UO_538 (O_538,N_24581,N_24875);
or UO_539 (O_539,N_24947,N_24890);
xor UO_540 (O_540,N_24534,N_24439);
nor UO_541 (O_541,N_24415,N_24569);
or UO_542 (O_542,N_24768,N_24390);
and UO_543 (O_543,N_24659,N_24748);
or UO_544 (O_544,N_24692,N_24961);
nor UO_545 (O_545,N_24475,N_24724);
and UO_546 (O_546,N_24634,N_24791);
xnor UO_547 (O_547,N_24376,N_24941);
and UO_548 (O_548,N_24652,N_24755);
and UO_549 (O_549,N_24587,N_24514);
nand UO_550 (O_550,N_24783,N_24959);
xor UO_551 (O_551,N_24810,N_24619);
and UO_552 (O_552,N_24473,N_24427);
nor UO_553 (O_553,N_24692,N_24787);
and UO_554 (O_554,N_24949,N_24868);
nor UO_555 (O_555,N_24889,N_24393);
xnor UO_556 (O_556,N_24663,N_24532);
nand UO_557 (O_557,N_24842,N_24863);
or UO_558 (O_558,N_24600,N_24848);
and UO_559 (O_559,N_24563,N_24791);
nor UO_560 (O_560,N_24516,N_24809);
and UO_561 (O_561,N_24523,N_24524);
nor UO_562 (O_562,N_24686,N_24746);
nor UO_563 (O_563,N_24884,N_24994);
xnor UO_564 (O_564,N_24576,N_24961);
xnor UO_565 (O_565,N_24462,N_24821);
xnor UO_566 (O_566,N_24643,N_24494);
nor UO_567 (O_567,N_24619,N_24840);
xnor UO_568 (O_568,N_24532,N_24946);
nor UO_569 (O_569,N_24840,N_24401);
xor UO_570 (O_570,N_24722,N_24454);
nand UO_571 (O_571,N_24547,N_24420);
and UO_572 (O_572,N_24689,N_24948);
xnor UO_573 (O_573,N_24420,N_24695);
xor UO_574 (O_574,N_24858,N_24838);
or UO_575 (O_575,N_24902,N_24868);
xor UO_576 (O_576,N_24948,N_24670);
or UO_577 (O_577,N_24649,N_24652);
nor UO_578 (O_578,N_24878,N_24605);
and UO_579 (O_579,N_24599,N_24477);
nand UO_580 (O_580,N_24770,N_24880);
or UO_581 (O_581,N_24853,N_24928);
or UO_582 (O_582,N_24651,N_24538);
nand UO_583 (O_583,N_24478,N_24686);
xnor UO_584 (O_584,N_24765,N_24609);
nor UO_585 (O_585,N_24865,N_24512);
xnor UO_586 (O_586,N_24978,N_24710);
and UO_587 (O_587,N_24640,N_24807);
nor UO_588 (O_588,N_24481,N_24436);
xnor UO_589 (O_589,N_24731,N_24564);
and UO_590 (O_590,N_24547,N_24563);
or UO_591 (O_591,N_24754,N_24445);
or UO_592 (O_592,N_24395,N_24894);
xnor UO_593 (O_593,N_24576,N_24889);
nor UO_594 (O_594,N_24570,N_24635);
and UO_595 (O_595,N_24989,N_24428);
nor UO_596 (O_596,N_24629,N_24460);
xnor UO_597 (O_597,N_24716,N_24875);
nand UO_598 (O_598,N_24827,N_24692);
or UO_599 (O_599,N_24928,N_24488);
or UO_600 (O_600,N_24545,N_24714);
nand UO_601 (O_601,N_24669,N_24749);
xor UO_602 (O_602,N_24724,N_24938);
nand UO_603 (O_603,N_24627,N_24679);
and UO_604 (O_604,N_24918,N_24802);
and UO_605 (O_605,N_24840,N_24422);
nand UO_606 (O_606,N_24454,N_24568);
xnor UO_607 (O_607,N_24641,N_24818);
and UO_608 (O_608,N_24560,N_24856);
nand UO_609 (O_609,N_24727,N_24767);
and UO_610 (O_610,N_24795,N_24482);
nand UO_611 (O_611,N_24536,N_24684);
or UO_612 (O_612,N_24790,N_24473);
and UO_613 (O_613,N_24873,N_24568);
or UO_614 (O_614,N_24909,N_24449);
nor UO_615 (O_615,N_24502,N_24444);
nor UO_616 (O_616,N_24977,N_24756);
nor UO_617 (O_617,N_24912,N_24742);
nand UO_618 (O_618,N_24790,N_24965);
nand UO_619 (O_619,N_24702,N_24382);
nand UO_620 (O_620,N_24557,N_24572);
and UO_621 (O_621,N_24540,N_24730);
xor UO_622 (O_622,N_24701,N_24599);
nand UO_623 (O_623,N_24381,N_24919);
or UO_624 (O_624,N_24819,N_24728);
nor UO_625 (O_625,N_24487,N_24738);
nand UO_626 (O_626,N_24696,N_24594);
xnor UO_627 (O_627,N_24726,N_24418);
nand UO_628 (O_628,N_24836,N_24914);
and UO_629 (O_629,N_24953,N_24902);
or UO_630 (O_630,N_24613,N_24529);
xor UO_631 (O_631,N_24824,N_24915);
or UO_632 (O_632,N_24631,N_24783);
and UO_633 (O_633,N_24752,N_24527);
xnor UO_634 (O_634,N_24967,N_24744);
xor UO_635 (O_635,N_24975,N_24768);
or UO_636 (O_636,N_24997,N_24910);
or UO_637 (O_637,N_24773,N_24924);
xor UO_638 (O_638,N_24553,N_24427);
and UO_639 (O_639,N_24764,N_24994);
or UO_640 (O_640,N_24762,N_24464);
nor UO_641 (O_641,N_24747,N_24677);
xnor UO_642 (O_642,N_24998,N_24859);
xor UO_643 (O_643,N_24677,N_24840);
and UO_644 (O_644,N_24696,N_24518);
and UO_645 (O_645,N_24524,N_24951);
xor UO_646 (O_646,N_24843,N_24921);
nand UO_647 (O_647,N_24550,N_24600);
xnor UO_648 (O_648,N_24485,N_24658);
and UO_649 (O_649,N_24770,N_24979);
nor UO_650 (O_650,N_24502,N_24792);
and UO_651 (O_651,N_24984,N_24799);
xnor UO_652 (O_652,N_24855,N_24665);
nor UO_653 (O_653,N_24879,N_24854);
nand UO_654 (O_654,N_24668,N_24458);
nor UO_655 (O_655,N_24688,N_24813);
xor UO_656 (O_656,N_24724,N_24707);
xor UO_657 (O_657,N_24981,N_24752);
or UO_658 (O_658,N_24878,N_24604);
nand UO_659 (O_659,N_24693,N_24827);
xor UO_660 (O_660,N_24800,N_24949);
nand UO_661 (O_661,N_24630,N_24714);
nand UO_662 (O_662,N_24942,N_24810);
nor UO_663 (O_663,N_24496,N_24594);
or UO_664 (O_664,N_24591,N_24978);
xor UO_665 (O_665,N_24561,N_24606);
nand UO_666 (O_666,N_24644,N_24459);
nand UO_667 (O_667,N_24572,N_24437);
nand UO_668 (O_668,N_24564,N_24935);
xnor UO_669 (O_669,N_24385,N_24397);
nand UO_670 (O_670,N_24428,N_24848);
or UO_671 (O_671,N_24747,N_24786);
and UO_672 (O_672,N_24692,N_24829);
xnor UO_673 (O_673,N_24475,N_24692);
or UO_674 (O_674,N_24522,N_24980);
or UO_675 (O_675,N_24642,N_24702);
nand UO_676 (O_676,N_24512,N_24937);
nand UO_677 (O_677,N_24770,N_24690);
nor UO_678 (O_678,N_24775,N_24482);
or UO_679 (O_679,N_24995,N_24872);
and UO_680 (O_680,N_24661,N_24602);
and UO_681 (O_681,N_24490,N_24759);
nand UO_682 (O_682,N_24603,N_24607);
and UO_683 (O_683,N_24693,N_24684);
xnor UO_684 (O_684,N_24460,N_24826);
and UO_685 (O_685,N_24547,N_24422);
or UO_686 (O_686,N_24747,N_24404);
and UO_687 (O_687,N_24741,N_24636);
or UO_688 (O_688,N_24914,N_24981);
xnor UO_689 (O_689,N_24588,N_24835);
xor UO_690 (O_690,N_24522,N_24548);
xor UO_691 (O_691,N_24567,N_24885);
nand UO_692 (O_692,N_24778,N_24507);
xor UO_693 (O_693,N_24642,N_24388);
or UO_694 (O_694,N_24668,N_24514);
xor UO_695 (O_695,N_24876,N_24548);
nor UO_696 (O_696,N_24628,N_24620);
or UO_697 (O_697,N_24705,N_24691);
and UO_698 (O_698,N_24528,N_24872);
nor UO_699 (O_699,N_24642,N_24525);
nand UO_700 (O_700,N_24736,N_24641);
and UO_701 (O_701,N_24389,N_24865);
and UO_702 (O_702,N_24789,N_24728);
nor UO_703 (O_703,N_24641,N_24698);
nor UO_704 (O_704,N_24401,N_24516);
nor UO_705 (O_705,N_24703,N_24401);
xor UO_706 (O_706,N_24939,N_24774);
or UO_707 (O_707,N_24999,N_24476);
xor UO_708 (O_708,N_24765,N_24404);
and UO_709 (O_709,N_24538,N_24492);
and UO_710 (O_710,N_24769,N_24623);
nand UO_711 (O_711,N_24465,N_24619);
nand UO_712 (O_712,N_24702,N_24807);
xor UO_713 (O_713,N_24512,N_24654);
and UO_714 (O_714,N_24521,N_24670);
and UO_715 (O_715,N_24941,N_24768);
and UO_716 (O_716,N_24873,N_24510);
and UO_717 (O_717,N_24846,N_24661);
nor UO_718 (O_718,N_24578,N_24615);
xor UO_719 (O_719,N_24709,N_24578);
nor UO_720 (O_720,N_24808,N_24450);
or UO_721 (O_721,N_24840,N_24595);
nand UO_722 (O_722,N_24682,N_24433);
and UO_723 (O_723,N_24985,N_24873);
nand UO_724 (O_724,N_24685,N_24489);
xor UO_725 (O_725,N_24618,N_24764);
or UO_726 (O_726,N_24961,N_24858);
nor UO_727 (O_727,N_24638,N_24710);
or UO_728 (O_728,N_24388,N_24685);
or UO_729 (O_729,N_24375,N_24704);
and UO_730 (O_730,N_24724,N_24464);
xnor UO_731 (O_731,N_24413,N_24651);
xor UO_732 (O_732,N_24771,N_24410);
and UO_733 (O_733,N_24406,N_24603);
and UO_734 (O_734,N_24394,N_24497);
or UO_735 (O_735,N_24844,N_24787);
xnor UO_736 (O_736,N_24419,N_24825);
nor UO_737 (O_737,N_24675,N_24629);
and UO_738 (O_738,N_24978,N_24741);
and UO_739 (O_739,N_24732,N_24829);
xor UO_740 (O_740,N_24815,N_24647);
or UO_741 (O_741,N_24603,N_24609);
and UO_742 (O_742,N_24548,N_24632);
nand UO_743 (O_743,N_24499,N_24598);
and UO_744 (O_744,N_24511,N_24999);
and UO_745 (O_745,N_24856,N_24896);
xor UO_746 (O_746,N_24592,N_24525);
nor UO_747 (O_747,N_24670,N_24529);
nor UO_748 (O_748,N_24723,N_24430);
nor UO_749 (O_749,N_24570,N_24860);
or UO_750 (O_750,N_24589,N_24429);
and UO_751 (O_751,N_24644,N_24897);
nor UO_752 (O_752,N_24705,N_24948);
or UO_753 (O_753,N_24624,N_24912);
nand UO_754 (O_754,N_24466,N_24781);
or UO_755 (O_755,N_24956,N_24895);
and UO_756 (O_756,N_24903,N_24661);
nand UO_757 (O_757,N_24817,N_24875);
or UO_758 (O_758,N_24660,N_24815);
xnor UO_759 (O_759,N_24587,N_24873);
xnor UO_760 (O_760,N_24819,N_24549);
and UO_761 (O_761,N_24586,N_24935);
or UO_762 (O_762,N_24737,N_24543);
or UO_763 (O_763,N_24663,N_24558);
or UO_764 (O_764,N_24841,N_24914);
and UO_765 (O_765,N_24517,N_24589);
nand UO_766 (O_766,N_24596,N_24474);
nand UO_767 (O_767,N_24825,N_24515);
or UO_768 (O_768,N_24513,N_24449);
xor UO_769 (O_769,N_24717,N_24518);
xnor UO_770 (O_770,N_24519,N_24663);
nand UO_771 (O_771,N_24931,N_24444);
and UO_772 (O_772,N_24607,N_24761);
nor UO_773 (O_773,N_24837,N_24833);
or UO_774 (O_774,N_24420,N_24487);
xor UO_775 (O_775,N_24968,N_24814);
nand UO_776 (O_776,N_24856,N_24954);
and UO_777 (O_777,N_24495,N_24604);
or UO_778 (O_778,N_24715,N_24601);
nand UO_779 (O_779,N_24773,N_24801);
nand UO_780 (O_780,N_24765,N_24719);
nor UO_781 (O_781,N_24713,N_24752);
nand UO_782 (O_782,N_24641,N_24743);
xor UO_783 (O_783,N_24408,N_24717);
or UO_784 (O_784,N_24720,N_24531);
xor UO_785 (O_785,N_24524,N_24797);
and UO_786 (O_786,N_24756,N_24600);
nor UO_787 (O_787,N_24645,N_24444);
xor UO_788 (O_788,N_24796,N_24652);
nor UO_789 (O_789,N_24689,N_24716);
xor UO_790 (O_790,N_24758,N_24633);
or UO_791 (O_791,N_24711,N_24549);
or UO_792 (O_792,N_24984,N_24588);
or UO_793 (O_793,N_24514,N_24941);
or UO_794 (O_794,N_24633,N_24628);
xor UO_795 (O_795,N_24911,N_24502);
xor UO_796 (O_796,N_24691,N_24402);
xor UO_797 (O_797,N_24428,N_24634);
nand UO_798 (O_798,N_24556,N_24381);
and UO_799 (O_799,N_24872,N_24979);
nand UO_800 (O_800,N_24695,N_24795);
or UO_801 (O_801,N_24883,N_24790);
and UO_802 (O_802,N_24515,N_24713);
and UO_803 (O_803,N_24730,N_24400);
nand UO_804 (O_804,N_24643,N_24570);
nand UO_805 (O_805,N_24486,N_24811);
nor UO_806 (O_806,N_24648,N_24969);
and UO_807 (O_807,N_24538,N_24602);
nor UO_808 (O_808,N_24850,N_24939);
and UO_809 (O_809,N_24680,N_24701);
xnor UO_810 (O_810,N_24623,N_24767);
xnor UO_811 (O_811,N_24904,N_24697);
nand UO_812 (O_812,N_24619,N_24395);
and UO_813 (O_813,N_24875,N_24977);
nand UO_814 (O_814,N_24419,N_24400);
and UO_815 (O_815,N_24621,N_24656);
nor UO_816 (O_816,N_24860,N_24880);
nand UO_817 (O_817,N_24788,N_24710);
nand UO_818 (O_818,N_24777,N_24474);
xnor UO_819 (O_819,N_24460,N_24644);
nor UO_820 (O_820,N_24633,N_24483);
and UO_821 (O_821,N_24644,N_24471);
xnor UO_822 (O_822,N_24479,N_24677);
or UO_823 (O_823,N_24872,N_24473);
nand UO_824 (O_824,N_24771,N_24932);
nand UO_825 (O_825,N_24764,N_24669);
nand UO_826 (O_826,N_24765,N_24955);
nand UO_827 (O_827,N_24646,N_24610);
nand UO_828 (O_828,N_24453,N_24952);
nor UO_829 (O_829,N_24786,N_24420);
xnor UO_830 (O_830,N_24576,N_24617);
xnor UO_831 (O_831,N_24532,N_24569);
and UO_832 (O_832,N_24785,N_24407);
nand UO_833 (O_833,N_24747,N_24968);
nor UO_834 (O_834,N_24624,N_24838);
xor UO_835 (O_835,N_24856,N_24573);
xnor UO_836 (O_836,N_24455,N_24911);
or UO_837 (O_837,N_24457,N_24802);
nand UO_838 (O_838,N_24716,N_24418);
nand UO_839 (O_839,N_24676,N_24449);
nand UO_840 (O_840,N_24613,N_24848);
nor UO_841 (O_841,N_24735,N_24392);
or UO_842 (O_842,N_24725,N_24745);
nand UO_843 (O_843,N_24523,N_24573);
nor UO_844 (O_844,N_24908,N_24976);
or UO_845 (O_845,N_24788,N_24692);
xor UO_846 (O_846,N_24413,N_24734);
nand UO_847 (O_847,N_24439,N_24536);
xnor UO_848 (O_848,N_24670,N_24810);
xor UO_849 (O_849,N_24425,N_24452);
nand UO_850 (O_850,N_24865,N_24973);
xor UO_851 (O_851,N_24587,N_24412);
xor UO_852 (O_852,N_24739,N_24781);
or UO_853 (O_853,N_24831,N_24401);
nor UO_854 (O_854,N_24999,N_24478);
nor UO_855 (O_855,N_24835,N_24498);
nand UO_856 (O_856,N_24399,N_24915);
nand UO_857 (O_857,N_24919,N_24570);
nand UO_858 (O_858,N_24792,N_24395);
nand UO_859 (O_859,N_24944,N_24599);
or UO_860 (O_860,N_24695,N_24947);
nand UO_861 (O_861,N_24481,N_24691);
nor UO_862 (O_862,N_24528,N_24994);
nor UO_863 (O_863,N_24407,N_24885);
nand UO_864 (O_864,N_24958,N_24972);
xnor UO_865 (O_865,N_24620,N_24581);
nor UO_866 (O_866,N_24700,N_24715);
xnor UO_867 (O_867,N_24714,N_24952);
and UO_868 (O_868,N_24547,N_24638);
or UO_869 (O_869,N_24825,N_24815);
nor UO_870 (O_870,N_24487,N_24867);
nor UO_871 (O_871,N_24430,N_24444);
nand UO_872 (O_872,N_24672,N_24920);
nor UO_873 (O_873,N_24888,N_24639);
nor UO_874 (O_874,N_24985,N_24391);
xnor UO_875 (O_875,N_24716,N_24654);
or UO_876 (O_876,N_24994,N_24716);
or UO_877 (O_877,N_24635,N_24757);
nor UO_878 (O_878,N_24814,N_24605);
and UO_879 (O_879,N_24832,N_24478);
nor UO_880 (O_880,N_24451,N_24577);
and UO_881 (O_881,N_24845,N_24744);
xor UO_882 (O_882,N_24586,N_24678);
or UO_883 (O_883,N_24955,N_24912);
or UO_884 (O_884,N_24567,N_24805);
xor UO_885 (O_885,N_24586,N_24566);
and UO_886 (O_886,N_24999,N_24619);
nand UO_887 (O_887,N_24391,N_24797);
nand UO_888 (O_888,N_24721,N_24464);
nand UO_889 (O_889,N_24490,N_24624);
nor UO_890 (O_890,N_24894,N_24543);
and UO_891 (O_891,N_24659,N_24634);
and UO_892 (O_892,N_24605,N_24998);
or UO_893 (O_893,N_24776,N_24718);
nor UO_894 (O_894,N_24677,N_24998);
nor UO_895 (O_895,N_24943,N_24951);
or UO_896 (O_896,N_24983,N_24807);
nor UO_897 (O_897,N_24668,N_24575);
nor UO_898 (O_898,N_24914,N_24378);
nor UO_899 (O_899,N_24904,N_24686);
or UO_900 (O_900,N_24767,N_24946);
and UO_901 (O_901,N_24576,N_24624);
nand UO_902 (O_902,N_24575,N_24709);
and UO_903 (O_903,N_24948,N_24826);
nor UO_904 (O_904,N_24881,N_24464);
xnor UO_905 (O_905,N_24724,N_24846);
or UO_906 (O_906,N_24967,N_24916);
nand UO_907 (O_907,N_24772,N_24410);
nor UO_908 (O_908,N_24405,N_24568);
xnor UO_909 (O_909,N_24705,N_24601);
nor UO_910 (O_910,N_24900,N_24857);
nor UO_911 (O_911,N_24884,N_24965);
and UO_912 (O_912,N_24552,N_24476);
nand UO_913 (O_913,N_24733,N_24417);
nand UO_914 (O_914,N_24666,N_24492);
nor UO_915 (O_915,N_24461,N_24867);
xnor UO_916 (O_916,N_24854,N_24553);
and UO_917 (O_917,N_24732,N_24873);
and UO_918 (O_918,N_24391,N_24636);
and UO_919 (O_919,N_24696,N_24842);
or UO_920 (O_920,N_24844,N_24746);
and UO_921 (O_921,N_24917,N_24447);
and UO_922 (O_922,N_24980,N_24493);
and UO_923 (O_923,N_24841,N_24649);
or UO_924 (O_924,N_24873,N_24616);
or UO_925 (O_925,N_24387,N_24454);
or UO_926 (O_926,N_24909,N_24384);
and UO_927 (O_927,N_24709,N_24445);
and UO_928 (O_928,N_24702,N_24413);
and UO_929 (O_929,N_24625,N_24749);
and UO_930 (O_930,N_24841,N_24784);
or UO_931 (O_931,N_24846,N_24905);
or UO_932 (O_932,N_24470,N_24672);
nor UO_933 (O_933,N_24894,N_24780);
and UO_934 (O_934,N_24680,N_24518);
nand UO_935 (O_935,N_24869,N_24589);
nor UO_936 (O_936,N_24497,N_24709);
nand UO_937 (O_937,N_24610,N_24484);
nor UO_938 (O_938,N_24427,N_24792);
or UO_939 (O_939,N_24959,N_24851);
and UO_940 (O_940,N_24463,N_24739);
or UO_941 (O_941,N_24575,N_24860);
or UO_942 (O_942,N_24483,N_24679);
xnor UO_943 (O_943,N_24978,N_24818);
and UO_944 (O_944,N_24758,N_24887);
nor UO_945 (O_945,N_24694,N_24416);
nand UO_946 (O_946,N_24384,N_24536);
xor UO_947 (O_947,N_24474,N_24895);
or UO_948 (O_948,N_24932,N_24793);
nand UO_949 (O_949,N_24960,N_24658);
xor UO_950 (O_950,N_24815,N_24848);
nor UO_951 (O_951,N_24670,N_24685);
xor UO_952 (O_952,N_24397,N_24884);
xor UO_953 (O_953,N_24739,N_24825);
and UO_954 (O_954,N_24802,N_24637);
or UO_955 (O_955,N_24479,N_24797);
xnor UO_956 (O_956,N_24720,N_24635);
or UO_957 (O_957,N_24687,N_24723);
xor UO_958 (O_958,N_24450,N_24500);
and UO_959 (O_959,N_24857,N_24972);
and UO_960 (O_960,N_24829,N_24835);
or UO_961 (O_961,N_24627,N_24465);
nor UO_962 (O_962,N_24429,N_24615);
xnor UO_963 (O_963,N_24819,N_24885);
nand UO_964 (O_964,N_24622,N_24386);
nand UO_965 (O_965,N_24915,N_24443);
nor UO_966 (O_966,N_24670,N_24874);
or UO_967 (O_967,N_24940,N_24558);
or UO_968 (O_968,N_24542,N_24643);
and UO_969 (O_969,N_24941,N_24616);
xnor UO_970 (O_970,N_24616,N_24500);
and UO_971 (O_971,N_24716,N_24722);
nor UO_972 (O_972,N_24405,N_24754);
nand UO_973 (O_973,N_24397,N_24469);
and UO_974 (O_974,N_24691,N_24472);
or UO_975 (O_975,N_24909,N_24503);
or UO_976 (O_976,N_24406,N_24628);
nor UO_977 (O_977,N_24966,N_24631);
nor UO_978 (O_978,N_24899,N_24810);
or UO_979 (O_979,N_24549,N_24560);
and UO_980 (O_980,N_24949,N_24383);
nand UO_981 (O_981,N_24660,N_24533);
nand UO_982 (O_982,N_24737,N_24661);
or UO_983 (O_983,N_24983,N_24457);
or UO_984 (O_984,N_24735,N_24801);
xnor UO_985 (O_985,N_24535,N_24570);
xnor UO_986 (O_986,N_24662,N_24920);
nor UO_987 (O_987,N_24882,N_24996);
xnor UO_988 (O_988,N_24660,N_24727);
and UO_989 (O_989,N_24442,N_24650);
nor UO_990 (O_990,N_24575,N_24517);
or UO_991 (O_991,N_24424,N_24731);
nor UO_992 (O_992,N_24421,N_24937);
nor UO_993 (O_993,N_24441,N_24827);
nand UO_994 (O_994,N_24968,N_24937);
nand UO_995 (O_995,N_24416,N_24967);
nand UO_996 (O_996,N_24652,N_24630);
or UO_997 (O_997,N_24760,N_24992);
xor UO_998 (O_998,N_24452,N_24535);
nor UO_999 (O_999,N_24513,N_24747);
nor UO_1000 (O_1000,N_24988,N_24734);
nor UO_1001 (O_1001,N_24809,N_24543);
nor UO_1002 (O_1002,N_24472,N_24380);
xor UO_1003 (O_1003,N_24977,N_24576);
and UO_1004 (O_1004,N_24894,N_24816);
and UO_1005 (O_1005,N_24976,N_24800);
nand UO_1006 (O_1006,N_24569,N_24459);
or UO_1007 (O_1007,N_24545,N_24613);
and UO_1008 (O_1008,N_24664,N_24387);
nor UO_1009 (O_1009,N_24528,N_24640);
or UO_1010 (O_1010,N_24394,N_24591);
xnor UO_1011 (O_1011,N_24441,N_24738);
or UO_1012 (O_1012,N_24538,N_24515);
nor UO_1013 (O_1013,N_24895,N_24751);
nand UO_1014 (O_1014,N_24993,N_24970);
nor UO_1015 (O_1015,N_24488,N_24577);
nor UO_1016 (O_1016,N_24525,N_24886);
or UO_1017 (O_1017,N_24587,N_24513);
nand UO_1018 (O_1018,N_24784,N_24425);
xor UO_1019 (O_1019,N_24774,N_24624);
or UO_1020 (O_1020,N_24799,N_24560);
xnor UO_1021 (O_1021,N_24940,N_24413);
nand UO_1022 (O_1022,N_24399,N_24867);
xor UO_1023 (O_1023,N_24799,N_24433);
xor UO_1024 (O_1024,N_24516,N_24694);
nor UO_1025 (O_1025,N_24377,N_24755);
xor UO_1026 (O_1026,N_24500,N_24927);
xnor UO_1027 (O_1027,N_24922,N_24651);
nand UO_1028 (O_1028,N_24847,N_24946);
and UO_1029 (O_1029,N_24426,N_24854);
nor UO_1030 (O_1030,N_24391,N_24531);
nand UO_1031 (O_1031,N_24411,N_24689);
and UO_1032 (O_1032,N_24402,N_24609);
nand UO_1033 (O_1033,N_24550,N_24982);
xnor UO_1034 (O_1034,N_24622,N_24403);
or UO_1035 (O_1035,N_24811,N_24810);
or UO_1036 (O_1036,N_24686,N_24955);
or UO_1037 (O_1037,N_24981,N_24650);
or UO_1038 (O_1038,N_24997,N_24526);
or UO_1039 (O_1039,N_24732,N_24678);
nand UO_1040 (O_1040,N_24803,N_24782);
xnor UO_1041 (O_1041,N_24877,N_24480);
or UO_1042 (O_1042,N_24942,N_24383);
or UO_1043 (O_1043,N_24612,N_24579);
or UO_1044 (O_1044,N_24903,N_24759);
and UO_1045 (O_1045,N_24697,N_24738);
xor UO_1046 (O_1046,N_24727,N_24741);
or UO_1047 (O_1047,N_24998,N_24493);
nand UO_1048 (O_1048,N_24401,N_24388);
xnor UO_1049 (O_1049,N_24997,N_24860);
nand UO_1050 (O_1050,N_24684,N_24443);
nor UO_1051 (O_1051,N_24562,N_24990);
xor UO_1052 (O_1052,N_24675,N_24744);
nand UO_1053 (O_1053,N_24541,N_24494);
and UO_1054 (O_1054,N_24852,N_24750);
nor UO_1055 (O_1055,N_24593,N_24818);
and UO_1056 (O_1056,N_24935,N_24892);
nand UO_1057 (O_1057,N_24994,N_24930);
xor UO_1058 (O_1058,N_24854,N_24978);
or UO_1059 (O_1059,N_24680,N_24583);
nor UO_1060 (O_1060,N_24675,N_24592);
or UO_1061 (O_1061,N_24903,N_24599);
and UO_1062 (O_1062,N_24828,N_24799);
and UO_1063 (O_1063,N_24597,N_24810);
nand UO_1064 (O_1064,N_24475,N_24431);
xor UO_1065 (O_1065,N_24862,N_24462);
or UO_1066 (O_1066,N_24842,N_24720);
nand UO_1067 (O_1067,N_24886,N_24385);
xor UO_1068 (O_1068,N_24759,N_24454);
nand UO_1069 (O_1069,N_24437,N_24685);
nor UO_1070 (O_1070,N_24751,N_24618);
and UO_1071 (O_1071,N_24487,N_24874);
and UO_1072 (O_1072,N_24472,N_24663);
nor UO_1073 (O_1073,N_24437,N_24490);
nor UO_1074 (O_1074,N_24803,N_24784);
xnor UO_1075 (O_1075,N_24456,N_24892);
xnor UO_1076 (O_1076,N_24965,N_24680);
and UO_1077 (O_1077,N_24553,N_24625);
or UO_1078 (O_1078,N_24500,N_24398);
nor UO_1079 (O_1079,N_24999,N_24920);
and UO_1080 (O_1080,N_24992,N_24395);
and UO_1081 (O_1081,N_24522,N_24636);
and UO_1082 (O_1082,N_24855,N_24948);
or UO_1083 (O_1083,N_24780,N_24420);
and UO_1084 (O_1084,N_24387,N_24487);
nand UO_1085 (O_1085,N_24436,N_24559);
and UO_1086 (O_1086,N_24846,N_24856);
xnor UO_1087 (O_1087,N_24603,N_24766);
and UO_1088 (O_1088,N_24891,N_24494);
nand UO_1089 (O_1089,N_24606,N_24773);
or UO_1090 (O_1090,N_24826,N_24411);
and UO_1091 (O_1091,N_24473,N_24698);
nor UO_1092 (O_1092,N_24489,N_24554);
and UO_1093 (O_1093,N_24729,N_24723);
or UO_1094 (O_1094,N_24401,N_24403);
and UO_1095 (O_1095,N_24826,N_24579);
and UO_1096 (O_1096,N_24621,N_24970);
nand UO_1097 (O_1097,N_24829,N_24611);
and UO_1098 (O_1098,N_24944,N_24477);
nand UO_1099 (O_1099,N_24628,N_24833);
nor UO_1100 (O_1100,N_24885,N_24733);
and UO_1101 (O_1101,N_24944,N_24396);
and UO_1102 (O_1102,N_24862,N_24888);
nand UO_1103 (O_1103,N_24697,N_24845);
xnor UO_1104 (O_1104,N_24711,N_24407);
and UO_1105 (O_1105,N_24436,N_24603);
nand UO_1106 (O_1106,N_24697,N_24652);
xor UO_1107 (O_1107,N_24530,N_24585);
xnor UO_1108 (O_1108,N_24577,N_24638);
nand UO_1109 (O_1109,N_24795,N_24395);
nand UO_1110 (O_1110,N_24612,N_24511);
nor UO_1111 (O_1111,N_24455,N_24834);
or UO_1112 (O_1112,N_24881,N_24612);
nand UO_1113 (O_1113,N_24821,N_24872);
or UO_1114 (O_1114,N_24411,N_24654);
xnor UO_1115 (O_1115,N_24842,N_24468);
nand UO_1116 (O_1116,N_24546,N_24640);
or UO_1117 (O_1117,N_24602,N_24558);
or UO_1118 (O_1118,N_24732,N_24594);
nor UO_1119 (O_1119,N_24651,N_24726);
or UO_1120 (O_1120,N_24828,N_24499);
xor UO_1121 (O_1121,N_24418,N_24459);
nand UO_1122 (O_1122,N_24581,N_24796);
and UO_1123 (O_1123,N_24971,N_24541);
or UO_1124 (O_1124,N_24388,N_24451);
and UO_1125 (O_1125,N_24385,N_24529);
xor UO_1126 (O_1126,N_24827,N_24880);
or UO_1127 (O_1127,N_24557,N_24788);
or UO_1128 (O_1128,N_24397,N_24414);
or UO_1129 (O_1129,N_24639,N_24876);
xor UO_1130 (O_1130,N_24828,N_24433);
xnor UO_1131 (O_1131,N_24459,N_24969);
nor UO_1132 (O_1132,N_24911,N_24447);
nand UO_1133 (O_1133,N_24463,N_24527);
nand UO_1134 (O_1134,N_24572,N_24900);
xnor UO_1135 (O_1135,N_24418,N_24715);
nand UO_1136 (O_1136,N_24525,N_24875);
xnor UO_1137 (O_1137,N_24477,N_24405);
nor UO_1138 (O_1138,N_24415,N_24568);
xnor UO_1139 (O_1139,N_24525,N_24711);
xor UO_1140 (O_1140,N_24987,N_24764);
or UO_1141 (O_1141,N_24618,N_24767);
xnor UO_1142 (O_1142,N_24375,N_24577);
or UO_1143 (O_1143,N_24950,N_24893);
xnor UO_1144 (O_1144,N_24634,N_24887);
and UO_1145 (O_1145,N_24396,N_24745);
or UO_1146 (O_1146,N_24816,N_24375);
or UO_1147 (O_1147,N_24746,N_24423);
nand UO_1148 (O_1148,N_24532,N_24493);
nor UO_1149 (O_1149,N_24566,N_24996);
nor UO_1150 (O_1150,N_24887,N_24990);
xnor UO_1151 (O_1151,N_24756,N_24694);
nand UO_1152 (O_1152,N_24655,N_24565);
and UO_1153 (O_1153,N_24430,N_24741);
nor UO_1154 (O_1154,N_24399,N_24614);
or UO_1155 (O_1155,N_24864,N_24921);
xor UO_1156 (O_1156,N_24922,N_24411);
nor UO_1157 (O_1157,N_24889,N_24642);
and UO_1158 (O_1158,N_24609,N_24415);
nand UO_1159 (O_1159,N_24526,N_24536);
nor UO_1160 (O_1160,N_24922,N_24976);
nor UO_1161 (O_1161,N_24487,N_24443);
xnor UO_1162 (O_1162,N_24623,N_24885);
nor UO_1163 (O_1163,N_24444,N_24831);
and UO_1164 (O_1164,N_24595,N_24436);
or UO_1165 (O_1165,N_24518,N_24707);
nand UO_1166 (O_1166,N_24737,N_24655);
and UO_1167 (O_1167,N_24855,N_24487);
nand UO_1168 (O_1168,N_24971,N_24532);
or UO_1169 (O_1169,N_24689,N_24486);
xnor UO_1170 (O_1170,N_24849,N_24573);
and UO_1171 (O_1171,N_24591,N_24557);
xnor UO_1172 (O_1172,N_24795,N_24518);
nand UO_1173 (O_1173,N_24682,N_24494);
nand UO_1174 (O_1174,N_24404,N_24812);
and UO_1175 (O_1175,N_24582,N_24980);
xnor UO_1176 (O_1176,N_24670,N_24811);
xor UO_1177 (O_1177,N_24624,N_24729);
nor UO_1178 (O_1178,N_24502,N_24710);
and UO_1179 (O_1179,N_24762,N_24775);
xor UO_1180 (O_1180,N_24776,N_24919);
nand UO_1181 (O_1181,N_24884,N_24485);
and UO_1182 (O_1182,N_24677,N_24510);
nand UO_1183 (O_1183,N_24964,N_24899);
nand UO_1184 (O_1184,N_24621,N_24427);
nand UO_1185 (O_1185,N_24876,N_24688);
xnor UO_1186 (O_1186,N_24673,N_24714);
and UO_1187 (O_1187,N_24400,N_24833);
nand UO_1188 (O_1188,N_24828,N_24529);
and UO_1189 (O_1189,N_24692,N_24660);
nor UO_1190 (O_1190,N_24888,N_24637);
nor UO_1191 (O_1191,N_24956,N_24475);
or UO_1192 (O_1192,N_24986,N_24574);
or UO_1193 (O_1193,N_24711,N_24757);
nor UO_1194 (O_1194,N_24401,N_24826);
or UO_1195 (O_1195,N_24821,N_24460);
nand UO_1196 (O_1196,N_24888,N_24426);
nor UO_1197 (O_1197,N_24983,N_24730);
nor UO_1198 (O_1198,N_24670,N_24913);
nor UO_1199 (O_1199,N_24768,N_24926);
or UO_1200 (O_1200,N_24481,N_24600);
xnor UO_1201 (O_1201,N_24765,N_24922);
and UO_1202 (O_1202,N_24453,N_24431);
and UO_1203 (O_1203,N_24989,N_24515);
nor UO_1204 (O_1204,N_24586,N_24845);
nor UO_1205 (O_1205,N_24850,N_24492);
xnor UO_1206 (O_1206,N_24852,N_24618);
nor UO_1207 (O_1207,N_24500,N_24414);
xor UO_1208 (O_1208,N_24614,N_24713);
nor UO_1209 (O_1209,N_24440,N_24705);
xor UO_1210 (O_1210,N_24582,N_24996);
xnor UO_1211 (O_1211,N_24442,N_24418);
or UO_1212 (O_1212,N_24540,N_24830);
and UO_1213 (O_1213,N_24762,N_24492);
nor UO_1214 (O_1214,N_24836,N_24597);
nor UO_1215 (O_1215,N_24718,N_24819);
xnor UO_1216 (O_1216,N_24515,N_24456);
xnor UO_1217 (O_1217,N_24393,N_24892);
and UO_1218 (O_1218,N_24658,N_24453);
or UO_1219 (O_1219,N_24730,N_24638);
xnor UO_1220 (O_1220,N_24546,N_24457);
xnor UO_1221 (O_1221,N_24926,N_24747);
or UO_1222 (O_1222,N_24568,N_24528);
nand UO_1223 (O_1223,N_24766,N_24884);
and UO_1224 (O_1224,N_24668,N_24833);
nor UO_1225 (O_1225,N_24604,N_24657);
nand UO_1226 (O_1226,N_24523,N_24396);
nor UO_1227 (O_1227,N_24430,N_24436);
nor UO_1228 (O_1228,N_24736,N_24739);
or UO_1229 (O_1229,N_24452,N_24761);
nand UO_1230 (O_1230,N_24976,N_24405);
or UO_1231 (O_1231,N_24607,N_24932);
nand UO_1232 (O_1232,N_24470,N_24682);
and UO_1233 (O_1233,N_24883,N_24561);
and UO_1234 (O_1234,N_24988,N_24908);
nand UO_1235 (O_1235,N_24851,N_24867);
or UO_1236 (O_1236,N_24624,N_24960);
and UO_1237 (O_1237,N_24649,N_24966);
or UO_1238 (O_1238,N_24771,N_24978);
nand UO_1239 (O_1239,N_24656,N_24702);
xor UO_1240 (O_1240,N_24531,N_24928);
nor UO_1241 (O_1241,N_24839,N_24992);
nor UO_1242 (O_1242,N_24642,N_24779);
xnor UO_1243 (O_1243,N_24537,N_24676);
nor UO_1244 (O_1244,N_24815,N_24609);
nand UO_1245 (O_1245,N_24976,N_24677);
nand UO_1246 (O_1246,N_24906,N_24744);
nand UO_1247 (O_1247,N_24847,N_24389);
xor UO_1248 (O_1248,N_24711,N_24859);
and UO_1249 (O_1249,N_24502,N_24790);
xor UO_1250 (O_1250,N_24884,N_24477);
nor UO_1251 (O_1251,N_24428,N_24747);
or UO_1252 (O_1252,N_24895,N_24472);
or UO_1253 (O_1253,N_24407,N_24846);
nor UO_1254 (O_1254,N_24849,N_24410);
and UO_1255 (O_1255,N_24617,N_24844);
and UO_1256 (O_1256,N_24389,N_24550);
nor UO_1257 (O_1257,N_24728,N_24731);
nor UO_1258 (O_1258,N_24865,N_24994);
nor UO_1259 (O_1259,N_24596,N_24910);
and UO_1260 (O_1260,N_24710,N_24408);
xnor UO_1261 (O_1261,N_24568,N_24895);
nor UO_1262 (O_1262,N_24983,N_24956);
or UO_1263 (O_1263,N_24763,N_24918);
nand UO_1264 (O_1264,N_24606,N_24717);
or UO_1265 (O_1265,N_24443,N_24931);
nor UO_1266 (O_1266,N_24520,N_24717);
nand UO_1267 (O_1267,N_24508,N_24782);
xor UO_1268 (O_1268,N_24951,N_24651);
and UO_1269 (O_1269,N_24722,N_24447);
xor UO_1270 (O_1270,N_24488,N_24859);
nand UO_1271 (O_1271,N_24493,N_24842);
xor UO_1272 (O_1272,N_24914,N_24804);
nand UO_1273 (O_1273,N_24872,N_24573);
or UO_1274 (O_1274,N_24509,N_24839);
or UO_1275 (O_1275,N_24562,N_24591);
or UO_1276 (O_1276,N_24678,N_24734);
and UO_1277 (O_1277,N_24582,N_24899);
nand UO_1278 (O_1278,N_24793,N_24592);
or UO_1279 (O_1279,N_24868,N_24801);
nand UO_1280 (O_1280,N_24450,N_24489);
nand UO_1281 (O_1281,N_24863,N_24766);
nand UO_1282 (O_1282,N_24868,N_24375);
nand UO_1283 (O_1283,N_24400,N_24562);
xor UO_1284 (O_1284,N_24671,N_24948);
xnor UO_1285 (O_1285,N_24481,N_24617);
nor UO_1286 (O_1286,N_24753,N_24723);
and UO_1287 (O_1287,N_24594,N_24483);
nor UO_1288 (O_1288,N_24932,N_24861);
nor UO_1289 (O_1289,N_24982,N_24699);
and UO_1290 (O_1290,N_24901,N_24711);
nor UO_1291 (O_1291,N_24816,N_24974);
or UO_1292 (O_1292,N_24891,N_24550);
and UO_1293 (O_1293,N_24964,N_24903);
xnor UO_1294 (O_1294,N_24918,N_24762);
and UO_1295 (O_1295,N_24653,N_24440);
nand UO_1296 (O_1296,N_24915,N_24437);
xnor UO_1297 (O_1297,N_24445,N_24772);
and UO_1298 (O_1298,N_24641,N_24539);
nand UO_1299 (O_1299,N_24679,N_24743);
xor UO_1300 (O_1300,N_24527,N_24808);
or UO_1301 (O_1301,N_24907,N_24755);
nor UO_1302 (O_1302,N_24516,N_24614);
and UO_1303 (O_1303,N_24926,N_24827);
nand UO_1304 (O_1304,N_24794,N_24976);
and UO_1305 (O_1305,N_24469,N_24486);
or UO_1306 (O_1306,N_24882,N_24724);
nand UO_1307 (O_1307,N_24508,N_24464);
and UO_1308 (O_1308,N_24981,N_24404);
xor UO_1309 (O_1309,N_24595,N_24969);
nand UO_1310 (O_1310,N_24955,N_24702);
nor UO_1311 (O_1311,N_24902,N_24810);
or UO_1312 (O_1312,N_24823,N_24850);
and UO_1313 (O_1313,N_24962,N_24812);
or UO_1314 (O_1314,N_24815,N_24521);
and UO_1315 (O_1315,N_24861,N_24730);
xor UO_1316 (O_1316,N_24450,N_24864);
or UO_1317 (O_1317,N_24875,N_24737);
and UO_1318 (O_1318,N_24780,N_24541);
and UO_1319 (O_1319,N_24713,N_24559);
nand UO_1320 (O_1320,N_24488,N_24912);
nor UO_1321 (O_1321,N_24538,N_24891);
and UO_1322 (O_1322,N_24806,N_24992);
nor UO_1323 (O_1323,N_24381,N_24417);
nand UO_1324 (O_1324,N_24506,N_24923);
or UO_1325 (O_1325,N_24959,N_24647);
nor UO_1326 (O_1326,N_24732,N_24441);
nand UO_1327 (O_1327,N_24427,N_24974);
xor UO_1328 (O_1328,N_24987,N_24543);
nand UO_1329 (O_1329,N_24378,N_24450);
and UO_1330 (O_1330,N_24953,N_24660);
or UO_1331 (O_1331,N_24424,N_24502);
nor UO_1332 (O_1332,N_24734,N_24924);
xor UO_1333 (O_1333,N_24933,N_24986);
and UO_1334 (O_1334,N_24932,N_24587);
xor UO_1335 (O_1335,N_24458,N_24935);
nor UO_1336 (O_1336,N_24550,N_24889);
nor UO_1337 (O_1337,N_24671,N_24480);
xnor UO_1338 (O_1338,N_24731,N_24888);
and UO_1339 (O_1339,N_24973,N_24540);
xor UO_1340 (O_1340,N_24711,N_24765);
and UO_1341 (O_1341,N_24785,N_24634);
xor UO_1342 (O_1342,N_24649,N_24934);
nor UO_1343 (O_1343,N_24445,N_24440);
nand UO_1344 (O_1344,N_24913,N_24881);
nor UO_1345 (O_1345,N_24563,N_24566);
nand UO_1346 (O_1346,N_24421,N_24698);
nand UO_1347 (O_1347,N_24515,N_24733);
and UO_1348 (O_1348,N_24452,N_24537);
nand UO_1349 (O_1349,N_24912,N_24552);
nand UO_1350 (O_1350,N_24456,N_24381);
nand UO_1351 (O_1351,N_24987,N_24931);
or UO_1352 (O_1352,N_24915,N_24431);
or UO_1353 (O_1353,N_24816,N_24389);
nor UO_1354 (O_1354,N_24410,N_24376);
nand UO_1355 (O_1355,N_24693,N_24879);
and UO_1356 (O_1356,N_24428,N_24413);
xor UO_1357 (O_1357,N_24614,N_24886);
nand UO_1358 (O_1358,N_24866,N_24982);
xor UO_1359 (O_1359,N_24928,N_24622);
and UO_1360 (O_1360,N_24467,N_24674);
or UO_1361 (O_1361,N_24496,N_24890);
and UO_1362 (O_1362,N_24498,N_24508);
or UO_1363 (O_1363,N_24745,N_24444);
nand UO_1364 (O_1364,N_24517,N_24886);
nand UO_1365 (O_1365,N_24375,N_24478);
nand UO_1366 (O_1366,N_24733,N_24574);
nor UO_1367 (O_1367,N_24740,N_24491);
and UO_1368 (O_1368,N_24716,N_24730);
xnor UO_1369 (O_1369,N_24792,N_24950);
xnor UO_1370 (O_1370,N_24853,N_24782);
and UO_1371 (O_1371,N_24632,N_24958);
nor UO_1372 (O_1372,N_24885,N_24849);
or UO_1373 (O_1373,N_24688,N_24953);
xor UO_1374 (O_1374,N_24676,N_24551);
or UO_1375 (O_1375,N_24994,N_24743);
and UO_1376 (O_1376,N_24716,N_24666);
nor UO_1377 (O_1377,N_24484,N_24901);
xor UO_1378 (O_1378,N_24857,N_24546);
xnor UO_1379 (O_1379,N_24650,N_24614);
and UO_1380 (O_1380,N_24705,N_24774);
nand UO_1381 (O_1381,N_24528,N_24630);
xnor UO_1382 (O_1382,N_24669,N_24934);
nor UO_1383 (O_1383,N_24393,N_24434);
nand UO_1384 (O_1384,N_24383,N_24509);
and UO_1385 (O_1385,N_24584,N_24871);
nand UO_1386 (O_1386,N_24851,N_24814);
or UO_1387 (O_1387,N_24650,N_24798);
or UO_1388 (O_1388,N_24811,N_24655);
nor UO_1389 (O_1389,N_24647,N_24493);
nor UO_1390 (O_1390,N_24891,N_24930);
and UO_1391 (O_1391,N_24817,N_24885);
or UO_1392 (O_1392,N_24390,N_24595);
xnor UO_1393 (O_1393,N_24410,N_24973);
nor UO_1394 (O_1394,N_24626,N_24927);
nor UO_1395 (O_1395,N_24776,N_24620);
xor UO_1396 (O_1396,N_24459,N_24507);
nor UO_1397 (O_1397,N_24796,N_24714);
xnor UO_1398 (O_1398,N_24409,N_24450);
xor UO_1399 (O_1399,N_24885,N_24423);
or UO_1400 (O_1400,N_24712,N_24504);
nor UO_1401 (O_1401,N_24745,N_24925);
nor UO_1402 (O_1402,N_24838,N_24817);
or UO_1403 (O_1403,N_24770,N_24629);
or UO_1404 (O_1404,N_24673,N_24384);
nand UO_1405 (O_1405,N_24939,N_24478);
nor UO_1406 (O_1406,N_24542,N_24629);
nand UO_1407 (O_1407,N_24420,N_24980);
xor UO_1408 (O_1408,N_24486,N_24928);
xnor UO_1409 (O_1409,N_24450,N_24675);
or UO_1410 (O_1410,N_24778,N_24891);
nor UO_1411 (O_1411,N_24681,N_24900);
nor UO_1412 (O_1412,N_24482,N_24856);
nand UO_1413 (O_1413,N_24911,N_24424);
and UO_1414 (O_1414,N_24977,N_24786);
nor UO_1415 (O_1415,N_24532,N_24862);
or UO_1416 (O_1416,N_24389,N_24960);
or UO_1417 (O_1417,N_24870,N_24750);
and UO_1418 (O_1418,N_24852,N_24709);
xnor UO_1419 (O_1419,N_24974,N_24945);
nand UO_1420 (O_1420,N_24377,N_24978);
nor UO_1421 (O_1421,N_24537,N_24395);
or UO_1422 (O_1422,N_24768,N_24632);
or UO_1423 (O_1423,N_24747,N_24885);
nor UO_1424 (O_1424,N_24722,N_24888);
nand UO_1425 (O_1425,N_24512,N_24656);
or UO_1426 (O_1426,N_24843,N_24937);
or UO_1427 (O_1427,N_24578,N_24762);
or UO_1428 (O_1428,N_24468,N_24808);
and UO_1429 (O_1429,N_24668,N_24966);
and UO_1430 (O_1430,N_24681,N_24691);
nor UO_1431 (O_1431,N_24795,N_24557);
and UO_1432 (O_1432,N_24486,N_24613);
nand UO_1433 (O_1433,N_24594,N_24668);
xnor UO_1434 (O_1434,N_24504,N_24379);
xnor UO_1435 (O_1435,N_24402,N_24866);
xor UO_1436 (O_1436,N_24721,N_24611);
nor UO_1437 (O_1437,N_24758,N_24677);
and UO_1438 (O_1438,N_24888,N_24705);
nand UO_1439 (O_1439,N_24596,N_24642);
nand UO_1440 (O_1440,N_24613,N_24887);
nor UO_1441 (O_1441,N_24629,N_24910);
and UO_1442 (O_1442,N_24859,N_24792);
xor UO_1443 (O_1443,N_24418,N_24630);
nand UO_1444 (O_1444,N_24443,N_24562);
xnor UO_1445 (O_1445,N_24927,N_24946);
and UO_1446 (O_1446,N_24700,N_24638);
and UO_1447 (O_1447,N_24730,N_24897);
xor UO_1448 (O_1448,N_24712,N_24755);
nor UO_1449 (O_1449,N_24751,N_24652);
or UO_1450 (O_1450,N_24777,N_24588);
nor UO_1451 (O_1451,N_24481,N_24737);
xnor UO_1452 (O_1452,N_24377,N_24404);
nand UO_1453 (O_1453,N_24861,N_24639);
nand UO_1454 (O_1454,N_24645,N_24638);
and UO_1455 (O_1455,N_24908,N_24566);
nand UO_1456 (O_1456,N_24725,N_24955);
nand UO_1457 (O_1457,N_24846,N_24816);
xor UO_1458 (O_1458,N_24589,N_24490);
nor UO_1459 (O_1459,N_24440,N_24655);
or UO_1460 (O_1460,N_24721,N_24835);
nor UO_1461 (O_1461,N_24542,N_24795);
xnor UO_1462 (O_1462,N_24739,N_24488);
or UO_1463 (O_1463,N_24519,N_24925);
and UO_1464 (O_1464,N_24571,N_24461);
and UO_1465 (O_1465,N_24407,N_24725);
or UO_1466 (O_1466,N_24595,N_24605);
or UO_1467 (O_1467,N_24465,N_24599);
or UO_1468 (O_1468,N_24532,N_24867);
nor UO_1469 (O_1469,N_24633,N_24834);
nand UO_1470 (O_1470,N_24947,N_24821);
nor UO_1471 (O_1471,N_24835,N_24589);
nand UO_1472 (O_1472,N_24753,N_24700);
or UO_1473 (O_1473,N_24548,N_24637);
xnor UO_1474 (O_1474,N_24617,N_24869);
xnor UO_1475 (O_1475,N_24876,N_24516);
or UO_1476 (O_1476,N_24854,N_24475);
nand UO_1477 (O_1477,N_24971,N_24485);
and UO_1478 (O_1478,N_24726,N_24444);
and UO_1479 (O_1479,N_24995,N_24696);
xnor UO_1480 (O_1480,N_24786,N_24842);
or UO_1481 (O_1481,N_24506,N_24981);
and UO_1482 (O_1482,N_24705,N_24887);
nand UO_1483 (O_1483,N_24556,N_24931);
and UO_1484 (O_1484,N_24912,N_24813);
xnor UO_1485 (O_1485,N_24703,N_24559);
xnor UO_1486 (O_1486,N_24950,N_24517);
nand UO_1487 (O_1487,N_24791,N_24924);
and UO_1488 (O_1488,N_24444,N_24414);
nand UO_1489 (O_1489,N_24875,N_24654);
or UO_1490 (O_1490,N_24793,N_24839);
or UO_1491 (O_1491,N_24736,N_24608);
nand UO_1492 (O_1492,N_24582,N_24730);
xnor UO_1493 (O_1493,N_24846,N_24420);
or UO_1494 (O_1494,N_24398,N_24619);
xor UO_1495 (O_1495,N_24846,N_24827);
nor UO_1496 (O_1496,N_24755,N_24881);
nand UO_1497 (O_1497,N_24581,N_24996);
nand UO_1498 (O_1498,N_24962,N_24660);
or UO_1499 (O_1499,N_24802,N_24738);
and UO_1500 (O_1500,N_24538,N_24504);
xnor UO_1501 (O_1501,N_24525,N_24554);
nand UO_1502 (O_1502,N_24436,N_24628);
xnor UO_1503 (O_1503,N_24969,N_24970);
or UO_1504 (O_1504,N_24727,N_24865);
xor UO_1505 (O_1505,N_24656,N_24394);
xnor UO_1506 (O_1506,N_24695,N_24428);
or UO_1507 (O_1507,N_24531,N_24536);
xnor UO_1508 (O_1508,N_24758,N_24697);
nor UO_1509 (O_1509,N_24648,N_24718);
nor UO_1510 (O_1510,N_24588,N_24986);
nand UO_1511 (O_1511,N_24394,N_24786);
xor UO_1512 (O_1512,N_24760,N_24902);
or UO_1513 (O_1513,N_24987,N_24403);
nor UO_1514 (O_1514,N_24709,N_24752);
and UO_1515 (O_1515,N_24727,N_24791);
nor UO_1516 (O_1516,N_24761,N_24786);
nand UO_1517 (O_1517,N_24880,N_24883);
nand UO_1518 (O_1518,N_24510,N_24414);
nand UO_1519 (O_1519,N_24517,N_24920);
and UO_1520 (O_1520,N_24710,N_24621);
nor UO_1521 (O_1521,N_24942,N_24995);
or UO_1522 (O_1522,N_24610,N_24466);
xor UO_1523 (O_1523,N_24512,N_24637);
xor UO_1524 (O_1524,N_24493,N_24979);
nor UO_1525 (O_1525,N_24403,N_24954);
or UO_1526 (O_1526,N_24428,N_24462);
xor UO_1527 (O_1527,N_24701,N_24394);
nand UO_1528 (O_1528,N_24431,N_24659);
or UO_1529 (O_1529,N_24489,N_24930);
and UO_1530 (O_1530,N_24674,N_24548);
nand UO_1531 (O_1531,N_24904,N_24759);
nand UO_1532 (O_1532,N_24662,N_24743);
or UO_1533 (O_1533,N_24871,N_24666);
and UO_1534 (O_1534,N_24510,N_24415);
xor UO_1535 (O_1535,N_24891,N_24841);
nor UO_1536 (O_1536,N_24615,N_24979);
xnor UO_1537 (O_1537,N_24935,N_24573);
or UO_1538 (O_1538,N_24800,N_24986);
or UO_1539 (O_1539,N_24418,N_24526);
nor UO_1540 (O_1540,N_24873,N_24922);
and UO_1541 (O_1541,N_24724,N_24903);
and UO_1542 (O_1542,N_24793,N_24407);
and UO_1543 (O_1543,N_24911,N_24404);
and UO_1544 (O_1544,N_24734,N_24917);
nand UO_1545 (O_1545,N_24992,N_24836);
and UO_1546 (O_1546,N_24776,N_24515);
nand UO_1547 (O_1547,N_24517,N_24453);
xor UO_1548 (O_1548,N_24458,N_24516);
or UO_1549 (O_1549,N_24593,N_24706);
nor UO_1550 (O_1550,N_24644,N_24648);
nor UO_1551 (O_1551,N_24519,N_24878);
nand UO_1552 (O_1552,N_24969,N_24615);
and UO_1553 (O_1553,N_24628,N_24746);
xor UO_1554 (O_1554,N_24642,N_24860);
or UO_1555 (O_1555,N_24834,N_24879);
and UO_1556 (O_1556,N_24956,N_24992);
nand UO_1557 (O_1557,N_24754,N_24994);
and UO_1558 (O_1558,N_24741,N_24586);
nor UO_1559 (O_1559,N_24872,N_24924);
and UO_1560 (O_1560,N_24990,N_24965);
nor UO_1561 (O_1561,N_24801,N_24938);
nor UO_1562 (O_1562,N_24940,N_24856);
and UO_1563 (O_1563,N_24761,N_24386);
nand UO_1564 (O_1564,N_24643,N_24528);
nor UO_1565 (O_1565,N_24546,N_24603);
and UO_1566 (O_1566,N_24812,N_24546);
nor UO_1567 (O_1567,N_24739,N_24846);
nor UO_1568 (O_1568,N_24850,N_24852);
nor UO_1569 (O_1569,N_24893,N_24606);
xor UO_1570 (O_1570,N_24917,N_24819);
and UO_1571 (O_1571,N_24797,N_24539);
nor UO_1572 (O_1572,N_24442,N_24973);
and UO_1573 (O_1573,N_24818,N_24811);
nor UO_1574 (O_1574,N_24664,N_24825);
xnor UO_1575 (O_1575,N_24517,N_24949);
xor UO_1576 (O_1576,N_24616,N_24994);
nand UO_1577 (O_1577,N_24439,N_24827);
and UO_1578 (O_1578,N_24476,N_24840);
nand UO_1579 (O_1579,N_24395,N_24966);
or UO_1580 (O_1580,N_24961,N_24905);
xnor UO_1581 (O_1581,N_24936,N_24724);
nand UO_1582 (O_1582,N_24819,N_24645);
or UO_1583 (O_1583,N_24737,N_24620);
or UO_1584 (O_1584,N_24857,N_24898);
nand UO_1585 (O_1585,N_24950,N_24866);
or UO_1586 (O_1586,N_24756,N_24690);
xor UO_1587 (O_1587,N_24422,N_24747);
nor UO_1588 (O_1588,N_24792,N_24660);
or UO_1589 (O_1589,N_24711,N_24382);
xnor UO_1590 (O_1590,N_24648,N_24894);
nor UO_1591 (O_1591,N_24732,N_24847);
xnor UO_1592 (O_1592,N_24573,N_24613);
nor UO_1593 (O_1593,N_24559,N_24758);
nand UO_1594 (O_1594,N_24854,N_24969);
xor UO_1595 (O_1595,N_24677,N_24989);
nor UO_1596 (O_1596,N_24884,N_24681);
xor UO_1597 (O_1597,N_24856,N_24765);
xor UO_1598 (O_1598,N_24634,N_24723);
nand UO_1599 (O_1599,N_24961,N_24409);
and UO_1600 (O_1600,N_24942,N_24997);
or UO_1601 (O_1601,N_24741,N_24594);
or UO_1602 (O_1602,N_24777,N_24941);
or UO_1603 (O_1603,N_24522,N_24377);
or UO_1604 (O_1604,N_24388,N_24690);
and UO_1605 (O_1605,N_24877,N_24813);
and UO_1606 (O_1606,N_24901,N_24392);
and UO_1607 (O_1607,N_24592,N_24625);
and UO_1608 (O_1608,N_24902,N_24796);
nand UO_1609 (O_1609,N_24745,N_24952);
nand UO_1610 (O_1610,N_24620,N_24818);
nand UO_1611 (O_1611,N_24753,N_24759);
xnor UO_1612 (O_1612,N_24906,N_24565);
and UO_1613 (O_1613,N_24569,N_24983);
and UO_1614 (O_1614,N_24827,N_24934);
xor UO_1615 (O_1615,N_24383,N_24561);
nand UO_1616 (O_1616,N_24527,N_24847);
and UO_1617 (O_1617,N_24672,N_24472);
nand UO_1618 (O_1618,N_24945,N_24560);
xnor UO_1619 (O_1619,N_24886,N_24931);
xor UO_1620 (O_1620,N_24606,N_24572);
or UO_1621 (O_1621,N_24440,N_24677);
nand UO_1622 (O_1622,N_24600,N_24943);
xor UO_1623 (O_1623,N_24935,N_24910);
xnor UO_1624 (O_1624,N_24642,N_24519);
xnor UO_1625 (O_1625,N_24680,N_24933);
and UO_1626 (O_1626,N_24462,N_24692);
or UO_1627 (O_1627,N_24734,N_24822);
nand UO_1628 (O_1628,N_24905,N_24930);
and UO_1629 (O_1629,N_24888,N_24473);
and UO_1630 (O_1630,N_24930,N_24512);
xor UO_1631 (O_1631,N_24626,N_24520);
or UO_1632 (O_1632,N_24735,N_24880);
xnor UO_1633 (O_1633,N_24907,N_24956);
and UO_1634 (O_1634,N_24790,N_24514);
and UO_1635 (O_1635,N_24514,N_24763);
and UO_1636 (O_1636,N_24703,N_24536);
or UO_1637 (O_1637,N_24539,N_24766);
nor UO_1638 (O_1638,N_24876,N_24420);
xnor UO_1639 (O_1639,N_24854,N_24664);
or UO_1640 (O_1640,N_24729,N_24437);
xnor UO_1641 (O_1641,N_24614,N_24632);
or UO_1642 (O_1642,N_24731,N_24811);
nor UO_1643 (O_1643,N_24806,N_24713);
nand UO_1644 (O_1644,N_24540,N_24511);
and UO_1645 (O_1645,N_24725,N_24957);
or UO_1646 (O_1646,N_24653,N_24828);
or UO_1647 (O_1647,N_24454,N_24798);
and UO_1648 (O_1648,N_24718,N_24713);
or UO_1649 (O_1649,N_24831,N_24703);
nand UO_1650 (O_1650,N_24596,N_24550);
and UO_1651 (O_1651,N_24982,N_24771);
nor UO_1652 (O_1652,N_24833,N_24724);
or UO_1653 (O_1653,N_24484,N_24911);
or UO_1654 (O_1654,N_24437,N_24691);
xor UO_1655 (O_1655,N_24881,N_24629);
nand UO_1656 (O_1656,N_24426,N_24941);
and UO_1657 (O_1657,N_24638,N_24803);
nor UO_1658 (O_1658,N_24556,N_24906);
nand UO_1659 (O_1659,N_24918,N_24998);
nand UO_1660 (O_1660,N_24434,N_24380);
nand UO_1661 (O_1661,N_24672,N_24715);
nand UO_1662 (O_1662,N_24935,N_24845);
and UO_1663 (O_1663,N_24677,N_24739);
or UO_1664 (O_1664,N_24942,N_24957);
nand UO_1665 (O_1665,N_24753,N_24591);
nor UO_1666 (O_1666,N_24724,N_24802);
and UO_1667 (O_1667,N_24704,N_24965);
or UO_1668 (O_1668,N_24813,N_24607);
and UO_1669 (O_1669,N_24410,N_24491);
or UO_1670 (O_1670,N_24402,N_24986);
nand UO_1671 (O_1671,N_24655,N_24577);
or UO_1672 (O_1672,N_24593,N_24988);
nor UO_1673 (O_1673,N_24668,N_24676);
and UO_1674 (O_1674,N_24854,N_24520);
and UO_1675 (O_1675,N_24656,N_24449);
xnor UO_1676 (O_1676,N_24501,N_24848);
or UO_1677 (O_1677,N_24757,N_24516);
or UO_1678 (O_1678,N_24492,N_24823);
nor UO_1679 (O_1679,N_24414,N_24569);
and UO_1680 (O_1680,N_24587,N_24441);
and UO_1681 (O_1681,N_24828,N_24790);
or UO_1682 (O_1682,N_24624,N_24420);
nand UO_1683 (O_1683,N_24553,N_24386);
nor UO_1684 (O_1684,N_24841,N_24687);
nor UO_1685 (O_1685,N_24753,N_24481);
nand UO_1686 (O_1686,N_24483,N_24573);
xor UO_1687 (O_1687,N_24424,N_24765);
xor UO_1688 (O_1688,N_24989,N_24606);
nor UO_1689 (O_1689,N_24650,N_24491);
or UO_1690 (O_1690,N_24474,N_24798);
nand UO_1691 (O_1691,N_24631,N_24545);
xor UO_1692 (O_1692,N_24520,N_24559);
and UO_1693 (O_1693,N_24679,N_24956);
xnor UO_1694 (O_1694,N_24831,N_24433);
nand UO_1695 (O_1695,N_24378,N_24866);
nand UO_1696 (O_1696,N_24390,N_24420);
or UO_1697 (O_1697,N_24524,N_24932);
nand UO_1698 (O_1698,N_24396,N_24735);
nor UO_1699 (O_1699,N_24609,N_24735);
nand UO_1700 (O_1700,N_24570,N_24965);
and UO_1701 (O_1701,N_24719,N_24381);
or UO_1702 (O_1702,N_24774,N_24379);
xnor UO_1703 (O_1703,N_24744,N_24598);
nand UO_1704 (O_1704,N_24874,N_24770);
xnor UO_1705 (O_1705,N_24813,N_24837);
and UO_1706 (O_1706,N_24479,N_24482);
or UO_1707 (O_1707,N_24860,N_24694);
nor UO_1708 (O_1708,N_24992,N_24667);
or UO_1709 (O_1709,N_24706,N_24554);
nand UO_1710 (O_1710,N_24837,N_24838);
nor UO_1711 (O_1711,N_24706,N_24674);
nand UO_1712 (O_1712,N_24479,N_24926);
and UO_1713 (O_1713,N_24756,N_24615);
or UO_1714 (O_1714,N_24378,N_24711);
xnor UO_1715 (O_1715,N_24752,N_24548);
nand UO_1716 (O_1716,N_24672,N_24570);
or UO_1717 (O_1717,N_24826,N_24586);
xor UO_1718 (O_1718,N_24525,N_24485);
and UO_1719 (O_1719,N_24786,N_24682);
nor UO_1720 (O_1720,N_24561,N_24947);
or UO_1721 (O_1721,N_24792,N_24469);
xnor UO_1722 (O_1722,N_24820,N_24827);
nand UO_1723 (O_1723,N_24760,N_24770);
xor UO_1724 (O_1724,N_24683,N_24810);
nor UO_1725 (O_1725,N_24702,N_24536);
nand UO_1726 (O_1726,N_24831,N_24414);
and UO_1727 (O_1727,N_24435,N_24520);
nor UO_1728 (O_1728,N_24670,N_24609);
nor UO_1729 (O_1729,N_24602,N_24554);
nor UO_1730 (O_1730,N_24871,N_24887);
and UO_1731 (O_1731,N_24881,N_24781);
and UO_1732 (O_1732,N_24977,N_24845);
and UO_1733 (O_1733,N_24681,N_24986);
nand UO_1734 (O_1734,N_24485,N_24640);
or UO_1735 (O_1735,N_24668,N_24809);
nor UO_1736 (O_1736,N_24943,N_24892);
or UO_1737 (O_1737,N_24706,N_24605);
nor UO_1738 (O_1738,N_24586,N_24708);
nand UO_1739 (O_1739,N_24484,N_24792);
xor UO_1740 (O_1740,N_24707,N_24506);
nand UO_1741 (O_1741,N_24626,N_24933);
nand UO_1742 (O_1742,N_24889,N_24429);
and UO_1743 (O_1743,N_24404,N_24819);
or UO_1744 (O_1744,N_24936,N_24795);
or UO_1745 (O_1745,N_24813,N_24829);
xor UO_1746 (O_1746,N_24785,N_24475);
or UO_1747 (O_1747,N_24872,N_24839);
nand UO_1748 (O_1748,N_24823,N_24917);
or UO_1749 (O_1749,N_24398,N_24795);
or UO_1750 (O_1750,N_24492,N_24570);
and UO_1751 (O_1751,N_24873,N_24496);
xor UO_1752 (O_1752,N_24863,N_24893);
nand UO_1753 (O_1753,N_24573,N_24836);
and UO_1754 (O_1754,N_24539,N_24531);
and UO_1755 (O_1755,N_24387,N_24724);
xnor UO_1756 (O_1756,N_24865,N_24640);
or UO_1757 (O_1757,N_24626,N_24962);
xor UO_1758 (O_1758,N_24641,N_24538);
nor UO_1759 (O_1759,N_24757,N_24865);
or UO_1760 (O_1760,N_24492,N_24790);
or UO_1761 (O_1761,N_24680,N_24983);
nor UO_1762 (O_1762,N_24807,N_24753);
xnor UO_1763 (O_1763,N_24905,N_24387);
or UO_1764 (O_1764,N_24691,N_24455);
and UO_1765 (O_1765,N_24565,N_24969);
nor UO_1766 (O_1766,N_24951,N_24416);
xnor UO_1767 (O_1767,N_24603,N_24993);
nand UO_1768 (O_1768,N_24586,N_24631);
nand UO_1769 (O_1769,N_24585,N_24831);
nor UO_1770 (O_1770,N_24722,N_24891);
nand UO_1771 (O_1771,N_24953,N_24625);
xor UO_1772 (O_1772,N_24455,N_24930);
nor UO_1773 (O_1773,N_24806,N_24546);
or UO_1774 (O_1774,N_24538,N_24757);
and UO_1775 (O_1775,N_24986,N_24806);
or UO_1776 (O_1776,N_24742,N_24769);
xnor UO_1777 (O_1777,N_24648,N_24697);
or UO_1778 (O_1778,N_24725,N_24722);
and UO_1779 (O_1779,N_24553,N_24963);
nand UO_1780 (O_1780,N_24767,N_24834);
nand UO_1781 (O_1781,N_24574,N_24762);
xor UO_1782 (O_1782,N_24389,N_24632);
nor UO_1783 (O_1783,N_24792,N_24655);
nand UO_1784 (O_1784,N_24425,N_24873);
nand UO_1785 (O_1785,N_24755,N_24502);
and UO_1786 (O_1786,N_24929,N_24703);
or UO_1787 (O_1787,N_24823,N_24639);
nand UO_1788 (O_1788,N_24903,N_24496);
or UO_1789 (O_1789,N_24609,N_24938);
nor UO_1790 (O_1790,N_24888,N_24537);
or UO_1791 (O_1791,N_24520,N_24605);
nand UO_1792 (O_1792,N_24544,N_24862);
nand UO_1793 (O_1793,N_24955,N_24426);
and UO_1794 (O_1794,N_24712,N_24631);
or UO_1795 (O_1795,N_24664,N_24843);
and UO_1796 (O_1796,N_24483,N_24890);
nor UO_1797 (O_1797,N_24757,N_24649);
xnor UO_1798 (O_1798,N_24398,N_24910);
and UO_1799 (O_1799,N_24859,N_24819);
or UO_1800 (O_1800,N_24615,N_24727);
or UO_1801 (O_1801,N_24887,N_24478);
xor UO_1802 (O_1802,N_24996,N_24458);
nand UO_1803 (O_1803,N_24987,N_24483);
nand UO_1804 (O_1804,N_24870,N_24826);
or UO_1805 (O_1805,N_24580,N_24590);
nand UO_1806 (O_1806,N_24427,N_24633);
xor UO_1807 (O_1807,N_24928,N_24554);
or UO_1808 (O_1808,N_24431,N_24545);
or UO_1809 (O_1809,N_24863,N_24617);
xnor UO_1810 (O_1810,N_24828,N_24958);
nand UO_1811 (O_1811,N_24964,N_24857);
xnor UO_1812 (O_1812,N_24567,N_24724);
nor UO_1813 (O_1813,N_24386,N_24895);
xnor UO_1814 (O_1814,N_24399,N_24698);
nor UO_1815 (O_1815,N_24642,N_24505);
or UO_1816 (O_1816,N_24747,N_24756);
or UO_1817 (O_1817,N_24880,N_24476);
and UO_1818 (O_1818,N_24888,N_24971);
xnor UO_1819 (O_1819,N_24452,N_24424);
xor UO_1820 (O_1820,N_24877,N_24792);
or UO_1821 (O_1821,N_24763,N_24635);
nand UO_1822 (O_1822,N_24417,N_24861);
and UO_1823 (O_1823,N_24564,N_24598);
nand UO_1824 (O_1824,N_24908,N_24965);
xor UO_1825 (O_1825,N_24909,N_24687);
xnor UO_1826 (O_1826,N_24657,N_24735);
or UO_1827 (O_1827,N_24607,N_24475);
xor UO_1828 (O_1828,N_24777,N_24694);
nand UO_1829 (O_1829,N_24782,N_24713);
nor UO_1830 (O_1830,N_24502,N_24950);
xor UO_1831 (O_1831,N_24512,N_24674);
and UO_1832 (O_1832,N_24545,N_24806);
nand UO_1833 (O_1833,N_24641,N_24605);
nor UO_1834 (O_1834,N_24735,N_24381);
xor UO_1835 (O_1835,N_24625,N_24701);
nand UO_1836 (O_1836,N_24745,N_24932);
nand UO_1837 (O_1837,N_24768,N_24973);
xor UO_1838 (O_1838,N_24376,N_24394);
and UO_1839 (O_1839,N_24585,N_24788);
nand UO_1840 (O_1840,N_24778,N_24903);
xor UO_1841 (O_1841,N_24835,N_24546);
or UO_1842 (O_1842,N_24798,N_24560);
and UO_1843 (O_1843,N_24569,N_24442);
nand UO_1844 (O_1844,N_24815,N_24398);
or UO_1845 (O_1845,N_24790,N_24762);
xor UO_1846 (O_1846,N_24736,N_24380);
or UO_1847 (O_1847,N_24513,N_24482);
or UO_1848 (O_1848,N_24657,N_24406);
nor UO_1849 (O_1849,N_24686,N_24717);
nor UO_1850 (O_1850,N_24878,N_24460);
nand UO_1851 (O_1851,N_24428,N_24650);
nor UO_1852 (O_1852,N_24952,N_24855);
xnor UO_1853 (O_1853,N_24390,N_24885);
xnor UO_1854 (O_1854,N_24415,N_24684);
xnor UO_1855 (O_1855,N_24920,N_24918);
or UO_1856 (O_1856,N_24735,N_24389);
or UO_1857 (O_1857,N_24886,N_24491);
nor UO_1858 (O_1858,N_24581,N_24908);
and UO_1859 (O_1859,N_24605,N_24512);
and UO_1860 (O_1860,N_24929,N_24967);
or UO_1861 (O_1861,N_24484,N_24836);
nand UO_1862 (O_1862,N_24672,N_24793);
and UO_1863 (O_1863,N_24476,N_24844);
or UO_1864 (O_1864,N_24541,N_24570);
or UO_1865 (O_1865,N_24853,N_24676);
xnor UO_1866 (O_1866,N_24548,N_24490);
nand UO_1867 (O_1867,N_24406,N_24745);
nand UO_1868 (O_1868,N_24453,N_24424);
and UO_1869 (O_1869,N_24681,N_24851);
xnor UO_1870 (O_1870,N_24483,N_24758);
nor UO_1871 (O_1871,N_24803,N_24643);
nand UO_1872 (O_1872,N_24937,N_24524);
nand UO_1873 (O_1873,N_24742,N_24786);
nand UO_1874 (O_1874,N_24864,N_24735);
nor UO_1875 (O_1875,N_24716,N_24933);
or UO_1876 (O_1876,N_24571,N_24784);
nor UO_1877 (O_1877,N_24487,N_24398);
or UO_1878 (O_1878,N_24616,N_24708);
nand UO_1879 (O_1879,N_24704,N_24801);
nand UO_1880 (O_1880,N_24772,N_24473);
xor UO_1881 (O_1881,N_24811,N_24737);
nand UO_1882 (O_1882,N_24817,N_24393);
or UO_1883 (O_1883,N_24980,N_24444);
and UO_1884 (O_1884,N_24634,N_24617);
and UO_1885 (O_1885,N_24605,N_24845);
or UO_1886 (O_1886,N_24806,N_24919);
xnor UO_1887 (O_1887,N_24885,N_24972);
xnor UO_1888 (O_1888,N_24630,N_24998);
nor UO_1889 (O_1889,N_24916,N_24834);
nand UO_1890 (O_1890,N_24861,N_24477);
nand UO_1891 (O_1891,N_24518,N_24461);
and UO_1892 (O_1892,N_24508,N_24872);
nor UO_1893 (O_1893,N_24778,N_24807);
or UO_1894 (O_1894,N_24878,N_24525);
xor UO_1895 (O_1895,N_24802,N_24885);
xnor UO_1896 (O_1896,N_24425,N_24976);
nor UO_1897 (O_1897,N_24846,N_24925);
xnor UO_1898 (O_1898,N_24771,N_24704);
or UO_1899 (O_1899,N_24973,N_24858);
nor UO_1900 (O_1900,N_24768,N_24700);
or UO_1901 (O_1901,N_24976,N_24541);
nor UO_1902 (O_1902,N_24457,N_24746);
nand UO_1903 (O_1903,N_24799,N_24937);
nor UO_1904 (O_1904,N_24668,N_24606);
xor UO_1905 (O_1905,N_24960,N_24823);
xor UO_1906 (O_1906,N_24501,N_24658);
xor UO_1907 (O_1907,N_24655,N_24843);
nor UO_1908 (O_1908,N_24853,N_24656);
nand UO_1909 (O_1909,N_24492,N_24937);
nand UO_1910 (O_1910,N_24458,N_24989);
nand UO_1911 (O_1911,N_24446,N_24739);
xor UO_1912 (O_1912,N_24537,N_24730);
nor UO_1913 (O_1913,N_24479,N_24646);
nand UO_1914 (O_1914,N_24464,N_24956);
xor UO_1915 (O_1915,N_24753,N_24905);
or UO_1916 (O_1916,N_24557,N_24688);
xnor UO_1917 (O_1917,N_24604,N_24911);
and UO_1918 (O_1918,N_24529,N_24783);
or UO_1919 (O_1919,N_24834,N_24467);
xnor UO_1920 (O_1920,N_24909,N_24523);
xnor UO_1921 (O_1921,N_24858,N_24623);
nor UO_1922 (O_1922,N_24675,N_24379);
or UO_1923 (O_1923,N_24438,N_24864);
nor UO_1924 (O_1924,N_24557,N_24988);
nand UO_1925 (O_1925,N_24713,N_24797);
and UO_1926 (O_1926,N_24377,N_24744);
nor UO_1927 (O_1927,N_24466,N_24708);
and UO_1928 (O_1928,N_24429,N_24541);
xnor UO_1929 (O_1929,N_24968,N_24916);
xor UO_1930 (O_1930,N_24806,N_24711);
xor UO_1931 (O_1931,N_24850,N_24922);
nand UO_1932 (O_1932,N_24553,N_24581);
xnor UO_1933 (O_1933,N_24530,N_24500);
nand UO_1934 (O_1934,N_24517,N_24602);
and UO_1935 (O_1935,N_24375,N_24879);
and UO_1936 (O_1936,N_24409,N_24694);
and UO_1937 (O_1937,N_24985,N_24527);
or UO_1938 (O_1938,N_24905,N_24535);
or UO_1939 (O_1939,N_24678,N_24868);
and UO_1940 (O_1940,N_24938,N_24575);
xor UO_1941 (O_1941,N_24452,N_24484);
nor UO_1942 (O_1942,N_24532,N_24734);
xnor UO_1943 (O_1943,N_24543,N_24441);
nand UO_1944 (O_1944,N_24514,N_24641);
xor UO_1945 (O_1945,N_24703,N_24683);
nor UO_1946 (O_1946,N_24538,N_24752);
or UO_1947 (O_1947,N_24907,N_24820);
nand UO_1948 (O_1948,N_24977,N_24497);
xnor UO_1949 (O_1949,N_24596,N_24409);
nand UO_1950 (O_1950,N_24713,N_24967);
xor UO_1951 (O_1951,N_24508,N_24839);
nand UO_1952 (O_1952,N_24989,N_24567);
and UO_1953 (O_1953,N_24617,N_24592);
nand UO_1954 (O_1954,N_24884,N_24828);
or UO_1955 (O_1955,N_24858,N_24464);
xnor UO_1956 (O_1956,N_24896,N_24691);
nand UO_1957 (O_1957,N_24430,N_24585);
or UO_1958 (O_1958,N_24825,N_24749);
nor UO_1959 (O_1959,N_24874,N_24909);
nand UO_1960 (O_1960,N_24636,N_24776);
or UO_1961 (O_1961,N_24440,N_24989);
xnor UO_1962 (O_1962,N_24957,N_24413);
nand UO_1963 (O_1963,N_24829,N_24707);
xor UO_1964 (O_1964,N_24711,N_24598);
and UO_1965 (O_1965,N_24623,N_24729);
and UO_1966 (O_1966,N_24539,N_24692);
xnor UO_1967 (O_1967,N_24590,N_24846);
or UO_1968 (O_1968,N_24640,N_24550);
or UO_1969 (O_1969,N_24953,N_24940);
xnor UO_1970 (O_1970,N_24565,N_24555);
or UO_1971 (O_1971,N_24745,N_24791);
xor UO_1972 (O_1972,N_24887,N_24718);
and UO_1973 (O_1973,N_24949,N_24854);
nand UO_1974 (O_1974,N_24687,N_24384);
and UO_1975 (O_1975,N_24471,N_24639);
and UO_1976 (O_1976,N_24514,N_24733);
xnor UO_1977 (O_1977,N_24530,N_24445);
nand UO_1978 (O_1978,N_24517,N_24735);
or UO_1979 (O_1979,N_24573,N_24860);
nand UO_1980 (O_1980,N_24494,N_24958);
or UO_1981 (O_1981,N_24379,N_24826);
nand UO_1982 (O_1982,N_24457,N_24554);
xnor UO_1983 (O_1983,N_24526,N_24750);
or UO_1984 (O_1984,N_24911,N_24975);
and UO_1985 (O_1985,N_24573,N_24985);
nand UO_1986 (O_1986,N_24402,N_24857);
or UO_1987 (O_1987,N_24617,N_24953);
nor UO_1988 (O_1988,N_24884,N_24644);
nor UO_1989 (O_1989,N_24799,N_24911);
and UO_1990 (O_1990,N_24553,N_24576);
or UO_1991 (O_1991,N_24480,N_24911);
nor UO_1992 (O_1992,N_24463,N_24590);
and UO_1993 (O_1993,N_24564,N_24420);
or UO_1994 (O_1994,N_24440,N_24534);
xor UO_1995 (O_1995,N_24665,N_24383);
and UO_1996 (O_1996,N_24810,N_24532);
nor UO_1997 (O_1997,N_24647,N_24659);
or UO_1998 (O_1998,N_24748,N_24763);
and UO_1999 (O_1999,N_24993,N_24572);
and UO_2000 (O_2000,N_24450,N_24965);
or UO_2001 (O_2001,N_24663,N_24594);
xnor UO_2002 (O_2002,N_24378,N_24674);
and UO_2003 (O_2003,N_24573,N_24729);
xnor UO_2004 (O_2004,N_24958,N_24784);
xor UO_2005 (O_2005,N_24723,N_24909);
or UO_2006 (O_2006,N_24708,N_24723);
and UO_2007 (O_2007,N_24933,N_24811);
or UO_2008 (O_2008,N_24783,N_24494);
nor UO_2009 (O_2009,N_24651,N_24473);
nor UO_2010 (O_2010,N_24791,N_24695);
xnor UO_2011 (O_2011,N_24523,N_24730);
and UO_2012 (O_2012,N_24557,N_24385);
nand UO_2013 (O_2013,N_24743,N_24692);
and UO_2014 (O_2014,N_24709,N_24690);
xnor UO_2015 (O_2015,N_24958,N_24377);
nor UO_2016 (O_2016,N_24489,N_24407);
nor UO_2017 (O_2017,N_24967,N_24409);
and UO_2018 (O_2018,N_24767,N_24710);
nor UO_2019 (O_2019,N_24437,N_24566);
nor UO_2020 (O_2020,N_24393,N_24854);
xor UO_2021 (O_2021,N_24793,N_24390);
nand UO_2022 (O_2022,N_24530,N_24511);
nand UO_2023 (O_2023,N_24962,N_24662);
xor UO_2024 (O_2024,N_24913,N_24950);
nand UO_2025 (O_2025,N_24896,N_24412);
or UO_2026 (O_2026,N_24878,N_24711);
nand UO_2027 (O_2027,N_24504,N_24431);
and UO_2028 (O_2028,N_24672,N_24993);
nor UO_2029 (O_2029,N_24777,N_24807);
or UO_2030 (O_2030,N_24922,N_24386);
nor UO_2031 (O_2031,N_24745,N_24669);
xor UO_2032 (O_2032,N_24641,N_24380);
or UO_2033 (O_2033,N_24926,N_24777);
nand UO_2034 (O_2034,N_24553,N_24731);
and UO_2035 (O_2035,N_24809,N_24851);
nand UO_2036 (O_2036,N_24432,N_24717);
and UO_2037 (O_2037,N_24708,N_24731);
or UO_2038 (O_2038,N_24416,N_24619);
nand UO_2039 (O_2039,N_24485,N_24546);
nor UO_2040 (O_2040,N_24875,N_24412);
nand UO_2041 (O_2041,N_24619,N_24758);
nand UO_2042 (O_2042,N_24722,N_24634);
and UO_2043 (O_2043,N_24999,N_24952);
xnor UO_2044 (O_2044,N_24784,N_24699);
xor UO_2045 (O_2045,N_24946,N_24467);
and UO_2046 (O_2046,N_24719,N_24804);
xnor UO_2047 (O_2047,N_24592,N_24385);
xor UO_2048 (O_2048,N_24980,N_24533);
and UO_2049 (O_2049,N_24505,N_24845);
nor UO_2050 (O_2050,N_24675,N_24949);
nand UO_2051 (O_2051,N_24486,N_24926);
nor UO_2052 (O_2052,N_24745,N_24458);
or UO_2053 (O_2053,N_24602,N_24968);
nor UO_2054 (O_2054,N_24632,N_24565);
nand UO_2055 (O_2055,N_24578,N_24961);
nand UO_2056 (O_2056,N_24682,N_24683);
xor UO_2057 (O_2057,N_24848,N_24745);
and UO_2058 (O_2058,N_24870,N_24698);
or UO_2059 (O_2059,N_24683,N_24860);
xor UO_2060 (O_2060,N_24881,N_24875);
nand UO_2061 (O_2061,N_24672,N_24763);
or UO_2062 (O_2062,N_24782,N_24597);
and UO_2063 (O_2063,N_24820,N_24609);
and UO_2064 (O_2064,N_24377,N_24749);
or UO_2065 (O_2065,N_24789,N_24862);
or UO_2066 (O_2066,N_24455,N_24507);
nor UO_2067 (O_2067,N_24503,N_24806);
or UO_2068 (O_2068,N_24502,N_24579);
xor UO_2069 (O_2069,N_24747,N_24804);
nand UO_2070 (O_2070,N_24398,N_24410);
nor UO_2071 (O_2071,N_24967,N_24438);
or UO_2072 (O_2072,N_24591,N_24555);
xor UO_2073 (O_2073,N_24972,N_24829);
and UO_2074 (O_2074,N_24530,N_24964);
nor UO_2075 (O_2075,N_24799,N_24720);
and UO_2076 (O_2076,N_24756,N_24751);
nor UO_2077 (O_2077,N_24578,N_24935);
xor UO_2078 (O_2078,N_24967,N_24628);
xor UO_2079 (O_2079,N_24665,N_24478);
xnor UO_2080 (O_2080,N_24841,N_24576);
nand UO_2081 (O_2081,N_24385,N_24463);
or UO_2082 (O_2082,N_24674,N_24999);
xor UO_2083 (O_2083,N_24614,N_24389);
xnor UO_2084 (O_2084,N_24435,N_24878);
nor UO_2085 (O_2085,N_24961,N_24499);
or UO_2086 (O_2086,N_24641,N_24617);
nand UO_2087 (O_2087,N_24405,N_24811);
and UO_2088 (O_2088,N_24894,N_24567);
xor UO_2089 (O_2089,N_24536,N_24934);
nand UO_2090 (O_2090,N_24601,N_24431);
nor UO_2091 (O_2091,N_24925,N_24585);
xnor UO_2092 (O_2092,N_24999,N_24407);
and UO_2093 (O_2093,N_24572,N_24790);
nor UO_2094 (O_2094,N_24710,N_24848);
or UO_2095 (O_2095,N_24485,N_24436);
or UO_2096 (O_2096,N_24699,N_24477);
and UO_2097 (O_2097,N_24850,N_24397);
and UO_2098 (O_2098,N_24458,N_24461);
nand UO_2099 (O_2099,N_24687,N_24715);
nor UO_2100 (O_2100,N_24952,N_24376);
nand UO_2101 (O_2101,N_24501,N_24723);
or UO_2102 (O_2102,N_24638,N_24879);
nor UO_2103 (O_2103,N_24837,N_24649);
xor UO_2104 (O_2104,N_24734,N_24530);
and UO_2105 (O_2105,N_24782,N_24994);
or UO_2106 (O_2106,N_24376,N_24854);
nand UO_2107 (O_2107,N_24659,N_24482);
nand UO_2108 (O_2108,N_24701,N_24663);
nand UO_2109 (O_2109,N_24674,N_24825);
and UO_2110 (O_2110,N_24874,N_24483);
nand UO_2111 (O_2111,N_24996,N_24496);
nand UO_2112 (O_2112,N_24788,N_24600);
or UO_2113 (O_2113,N_24390,N_24832);
and UO_2114 (O_2114,N_24574,N_24630);
nand UO_2115 (O_2115,N_24838,N_24745);
xnor UO_2116 (O_2116,N_24650,N_24812);
or UO_2117 (O_2117,N_24996,N_24839);
or UO_2118 (O_2118,N_24970,N_24700);
xor UO_2119 (O_2119,N_24850,N_24759);
xnor UO_2120 (O_2120,N_24704,N_24686);
nand UO_2121 (O_2121,N_24705,N_24384);
xor UO_2122 (O_2122,N_24507,N_24727);
or UO_2123 (O_2123,N_24824,N_24544);
nor UO_2124 (O_2124,N_24492,N_24883);
nor UO_2125 (O_2125,N_24774,N_24636);
nor UO_2126 (O_2126,N_24998,N_24461);
and UO_2127 (O_2127,N_24636,N_24689);
nand UO_2128 (O_2128,N_24736,N_24583);
xnor UO_2129 (O_2129,N_24696,N_24495);
nand UO_2130 (O_2130,N_24944,N_24952);
and UO_2131 (O_2131,N_24882,N_24548);
nor UO_2132 (O_2132,N_24563,N_24865);
and UO_2133 (O_2133,N_24687,N_24416);
nor UO_2134 (O_2134,N_24515,N_24551);
xnor UO_2135 (O_2135,N_24384,N_24728);
or UO_2136 (O_2136,N_24727,N_24583);
nor UO_2137 (O_2137,N_24617,N_24398);
or UO_2138 (O_2138,N_24888,N_24853);
nor UO_2139 (O_2139,N_24629,N_24414);
or UO_2140 (O_2140,N_24653,N_24830);
or UO_2141 (O_2141,N_24710,N_24403);
nor UO_2142 (O_2142,N_24667,N_24937);
and UO_2143 (O_2143,N_24426,N_24512);
or UO_2144 (O_2144,N_24462,N_24996);
nand UO_2145 (O_2145,N_24666,N_24728);
or UO_2146 (O_2146,N_24617,N_24440);
nor UO_2147 (O_2147,N_24775,N_24417);
and UO_2148 (O_2148,N_24836,N_24925);
nand UO_2149 (O_2149,N_24482,N_24506);
and UO_2150 (O_2150,N_24875,N_24857);
nor UO_2151 (O_2151,N_24449,N_24409);
nand UO_2152 (O_2152,N_24821,N_24444);
nor UO_2153 (O_2153,N_24918,N_24609);
and UO_2154 (O_2154,N_24848,N_24407);
nand UO_2155 (O_2155,N_24995,N_24898);
xor UO_2156 (O_2156,N_24708,N_24918);
or UO_2157 (O_2157,N_24939,N_24965);
or UO_2158 (O_2158,N_24667,N_24996);
or UO_2159 (O_2159,N_24756,N_24606);
nor UO_2160 (O_2160,N_24632,N_24935);
xor UO_2161 (O_2161,N_24705,N_24603);
nor UO_2162 (O_2162,N_24636,N_24978);
or UO_2163 (O_2163,N_24566,N_24433);
nand UO_2164 (O_2164,N_24897,N_24529);
xor UO_2165 (O_2165,N_24956,N_24505);
or UO_2166 (O_2166,N_24614,N_24524);
or UO_2167 (O_2167,N_24480,N_24757);
or UO_2168 (O_2168,N_24449,N_24428);
nand UO_2169 (O_2169,N_24893,N_24981);
or UO_2170 (O_2170,N_24483,N_24622);
and UO_2171 (O_2171,N_24785,N_24798);
nand UO_2172 (O_2172,N_24815,N_24776);
or UO_2173 (O_2173,N_24610,N_24701);
xor UO_2174 (O_2174,N_24746,N_24700);
and UO_2175 (O_2175,N_24659,N_24906);
nor UO_2176 (O_2176,N_24922,N_24503);
nor UO_2177 (O_2177,N_24892,N_24801);
or UO_2178 (O_2178,N_24854,N_24551);
nand UO_2179 (O_2179,N_24706,N_24419);
and UO_2180 (O_2180,N_24781,N_24953);
xnor UO_2181 (O_2181,N_24915,N_24692);
nor UO_2182 (O_2182,N_24599,N_24692);
nand UO_2183 (O_2183,N_24582,N_24762);
nor UO_2184 (O_2184,N_24837,N_24599);
and UO_2185 (O_2185,N_24909,N_24694);
and UO_2186 (O_2186,N_24785,N_24601);
xnor UO_2187 (O_2187,N_24891,N_24500);
xnor UO_2188 (O_2188,N_24497,N_24767);
nand UO_2189 (O_2189,N_24827,N_24857);
nand UO_2190 (O_2190,N_24380,N_24547);
xor UO_2191 (O_2191,N_24867,N_24470);
and UO_2192 (O_2192,N_24417,N_24941);
xor UO_2193 (O_2193,N_24549,N_24935);
nand UO_2194 (O_2194,N_24466,N_24839);
nor UO_2195 (O_2195,N_24639,N_24706);
nor UO_2196 (O_2196,N_24994,N_24441);
nand UO_2197 (O_2197,N_24781,N_24420);
and UO_2198 (O_2198,N_24627,N_24636);
nand UO_2199 (O_2199,N_24978,N_24740);
xnor UO_2200 (O_2200,N_24923,N_24662);
nor UO_2201 (O_2201,N_24674,N_24717);
and UO_2202 (O_2202,N_24457,N_24855);
or UO_2203 (O_2203,N_24812,N_24500);
nor UO_2204 (O_2204,N_24724,N_24452);
or UO_2205 (O_2205,N_24887,N_24550);
and UO_2206 (O_2206,N_24727,N_24967);
or UO_2207 (O_2207,N_24626,N_24596);
or UO_2208 (O_2208,N_24567,N_24776);
xnor UO_2209 (O_2209,N_24870,N_24526);
or UO_2210 (O_2210,N_24424,N_24739);
nand UO_2211 (O_2211,N_24891,N_24957);
nor UO_2212 (O_2212,N_24540,N_24446);
xor UO_2213 (O_2213,N_24682,N_24939);
xnor UO_2214 (O_2214,N_24718,N_24429);
or UO_2215 (O_2215,N_24453,N_24417);
or UO_2216 (O_2216,N_24984,N_24784);
or UO_2217 (O_2217,N_24689,N_24714);
and UO_2218 (O_2218,N_24845,N_24416);
or UO_2219 (O_2219,N_24549,N_24577);
nand UO_2220 (O_2220,N_24493,N_24741);
xor UO_2221 (O_2221,N_24406,N_24458);
nor UO_2222 (O_2222,N_24744,N_24544);
and UO_2223 (O_2223,N_24739,N_24626);
and UO_2224 (O_2224,N_24659,N_24547);
nand UO_2225 (O_2225,N_24711,N_24869);
xor UO_2226 (O_2226,N_24927,N_24665);
and UO_2227 (O_2227,N_24839,N_24713);
and UO_2228 (O_2228,N_24939,N_24539);
nand UO_2229 (O_2229,N_24538,N_24763);
and UO_2230 (O_2230,N_24508,N_24494);
nor UO_2231 (O_2231,N_24994,N_24612);
and UO_2232 (O_2232,N_24592,N_24650);
nor UO_2233 (O_2233,N_24383,N_24990);
nor UO_2234 (O_2234,N_24831,N_24750);
and UO_2235 (O_2235,N_24532,N_24590);
or UO_2236 (O_2236,N_24977,N_24645);
nor UO_2237 (O_2237,N_24709,N_24405);
and UO_2238 (O_2238,N_24949,N_24543);
xor UO_2239 (O_2239,N_24977,N_24458);
or UO_2240 (O_2240,N_24823,N_24406);
and UO_2241 (O_2241,N_24701,N_24746);
and UO_2242 (O_2242,N_24465,N_24550);
xnor UO_2243 (O_2243,N_24489,N_24749);
and UO_2244 (O_2244,N_24695,N_24630);
nor UO_2245 (O_2245,N_24899,N_24860);
or UO_2246 (O_2246,N_24699,N_24668);
xor UO_2247 (O_2247,N_24632,N_24795);
nand UO_2248 (O_2248,N_24633,N_24490);
nand UO_2249 (O_2249,N_24649,N_24417);
nor UO_2250 (O_2250,N_24983,N_24949);
nor UO_2251 (O_2251,N_24875,N_24727);
xor UO_2252 (O_2252,N_24499,N_24706);
nor UO_2253 (O_2253,N_24406,N_24976);
xor UO_2254 (O_2254,N_24384,N_24866);
xor UO_2255 (O_2255,N_24461,N_24489);
and UO_2256 (O_2256,N_24566,N_24774);
nor UO_2257 (O_2257,N_24750,N_24911);
or UO_2258 (O_2258,N_24770,N_24402);
or UO_2259 (O_2259,N_24578,N_24375);
nor UO_2260 (O_2260,N_24465,N_24778);
xor UO_2261 (O_2261,N_24420,N_24848);
xnor UO_2262 (O_2262,N_24659,N_24442);
and UO_2263 (O_2263,N_24642,N_24883);
or UO_2264 (O_2264,N_24969,N_24428);
nand UO_2265 (O_2265,N_24717,N_24556);
nor UO_2266 (O_2266,N_24911,N_24457);
xor UO_2267 (O_2267,N_24443,N_24556);
and UO_2268 (O_2268,N_24813,N_24524);
xor UO_2269 (O_2269,N_24709,N_24916);
nand UO_2270 (O_2270,N_24816,N_24867);
nand UO_2271 (O_2271,N_24865,N_24561);
or UO_2272 (O_2272,N_24603,N_24449);
and UO_2273 (O_2273,N_24565,N_24462);
and UO_2274 (O_2274,N_24788,N_24693);
and UO_2275 (O_2275,N_24806,N_24885);
nand UO_2276 (O_2276,N_24683,N_24675);
nand UO_2277 (O_2277,N_24632,N_24476);
nor UO_2278 (O_2278,N_24581,N_24939);
nor UO_2279 (O_2279,N_24822,N_24799);
xor UO_2280 (O_2280,N_24989,N_24603);
nand UO_2281 (O_2281,N_24635,N_24437);
nand UO_2282 (O_2282,N_24847,N_24680);
and UO_2283 (O_2283,N_24630,N_24572);
nand UO_2284 (O_2284,N_24497,N_24598);
xnor UO_2285 (O_2285,N_24788,N_24496);
nor UO_2286 (O_2286,N_24981,N_24719);
nor UO_2287 (O_2287,N_24395,N_24611);
nand UO_2288 (O_2288,N_24574,N_24972);
xor UO_2289 (O_2289,N_24884,N_24713);
nand UO_2290 (O_2290,N_24953,N_24810);
nor UO_2291 (O_2291,N_24889,N_24489);
nor UO_2292 (O_2292,N_24394,N_24432);
nand UO_2293 (O_2293,N_24824,N_24474);
and UO_2294 (O_2294,N_24512,N_24683);
and UO_2295 (O_2295,N_24815,N_24585);
or UO_2296 (O_2296,N_24502,N_24852);
nand UO_2297 (O_2297,N_24762,N_24844);
and UO_2298 (O_2298,N_24625,N_24518);
xnor UO_2299 (O_2299,N_24618,N_24613);
xnor UO_2300 (O_2300,N_24879,N_24966);
nor UO_2301 (O_2301,N_24996,N_24733);
and UO_2302 (O_2302,N_24392,N_24764);
nor UO_2303 (O_2303,N_24916,N_24466);
and UO_2304 (O_2304,N_24472,N_24850);
and UO_2305 (O_2305,N_24484,N_24847);
nor UO_2306 (O_2306,N_24673,N_24741);
xnor UO_2307 (O_2307,N_24440,N_24537);
nor UO_2308 (O_2308,N_24918,N_24927);
xnor UO_2309 (O_2309,N_24531,N_24406);
nor UO_2310 (O_2310,N_24533,N_24955);
nand UO_2311 (O_2311,N_24412,N_24619);
nor UO_2312 (O_2312,N_24443,N_24929);
or UO_2313 (O_2313,N_24734,N_24411);
nor UO_2314 (O_2314,N_24520,N_24571);
xor UO_2315 (O_2315,N_24977,N_24572);
xnor UO_2316 (O_2316,N_24638,N_24904);
or UO_2317 (O_2317,N_24501,N_24910);
nand UO_2318 (O_2318,N_24846,N_24463);
and UO_2319 (O_2319,N_24906,N_24542);
and UO_2320 (O_2320,N_24680,N_24556);
or UO_2321 (O_2321,N_24832,N_24771);
nand UO_2322 (O_2322,N_24434,N_24792);
nand UO_2323 (O_2323,N_24525,N_24730);
or UO_2324 (O_2324,N_24722,N_24583);
and UO_2325 (O_2325,N_24405,N_24794);
xnor UO_2326 (O_2326,N_24975,N_24908);
and UO_2327 (O_2327,N_24563,N_24380);
and UO_2328 (O_2328,N_24879,N_24764);
and UO_2329 (O_2329,N_24902,N_24673);
xor UO_2330 (O_2330,N_24833,N_24778);
nand UO_2331 (O_2331,N_24441,N_24503);
xor UO_2332 (O_2332,N_24613,N_24388);
xor UO_2333 (O_2333,N_24733,N_24811);
nor UO_2334 (O_2334,N_24856,N_24981);
xnor UO_2335 (O_2335,N_24651,N_24691);
xor UO_2336 (O_2336,N_24645,N_24526);
nand UO_2337 (O_2337,N_24485,N_24869);
or UO_2338 (O_2338,N_24544,N_24499);
xor UO_2339 (O_2339,N_24523,N_24958);
nor UO_2340 (O_2340,N_24985,N_24438);
or UO_2341 (O_2341,N_24577,N_24499);
nor UO_2342 (O_2342,N_24625,N_24820);
nor UO_2343 (O_2343,N_24999,N_24990);
and UO_2344 (O_2344,N_24586,N_24418);
xor UO_2345 (O_2345,N_24532,N_24568);
nor UO_2346 (O_2346,N_24792,N_24778);
or UO_2347 (O_2347,N_24873,N_24956);
nand UO_2348 (O_2348,N_24920,N_24465);
and UO_2349 (O_2349,N_24533,N_24744);
and UO_2350 (O_2350,N_24393,N_24511);
nand UO_2351 (O_2351,N_24855,N_24836);
nor UO_2352 (O_2352,N_24484,N_24561);
nand UO_2353 (O_2353,N_24825,N_24559);
xnor UO_2354 (O_2354,N_24960,N_24927);
and UO_2355 (O_2355,N_24381,N_24623);
or UO_2356 (O_2356,N_24704,N_24540);
nor UO_2357 (O_2357,N_24865,N_24490);
nand UO_2358 (O_2358,N_24955,N_24863);
xor UO_2359 (O_2359,N_24584,N_24823);
or UO_2360 (O_2360,N_24702,N_24997);
nand UO_2361 (O_2361,N_24727,N_24529);
xnor UO_2362 (O_2362,N_24601,N_24477);
xor UO_2363 (O_2363,N_24707,N_24541);
nor UO_2364 (O_2364,N_24560,N_24861);
or UO_2365 (O_2365,N_24506,N_24699);
nor UO_2366 (O_2366,N_24884,N_24627);
nand UO_2367 (O_2367,N_24794,N_24880);
nand UO_2368 (O_2368,N_24793,N_24849);
or UO_2369 (O_2369,N_24731,N_24675);
xnor UO_2370 (O_2370,N_24621,N_24498);
or UO_2371 (O_2371,N_24593,N_24462);
nand UO_2372 (O_2372,N_24792,N_24953);
nor UO_2373 (O_2373,N_24716,N_24903);
and UO_2374 (O_2374,N_24544,N_24822);
xor UO_2375 (O_2375,N_24560,N_24724);
xor UO_2376 (O_2376,N_24968,N_24551);
and UO_2377 (O_2377,N_24557,N_24800);
nor UO_2378 (O_2378,N_24670,N_24788);
nand UO_2379 (O_2379,N_24776,N_24478);
xor UO_2380 (O_2380,N_24974,N_24521);
xor UO_2381 (O_2381,N_24995,N_24386);
nor UO_2382 (O_2382,N_24797,N_24385);
nor UO_2383 (O_2383,N_24852,N_24725);
xnor UO_2384 (O_2384,N_24459,N_24389);
nand UO_2385 (O_2385,N_24700,N_24870);
nor UO_2386 (O_2386,N_24644,N_24813);
and UO_2387 (O_2387,N_24943,N_24635);
nor UO_2388 (O_2388,N_24998,N_24628);
and UO_2389 (O_2389,N_24692,N_24497);
nor UO_2390 (O_2390,N_24846,N_24950);
nand UO_2391 (O_2391,N_24713,N_24385);
nand UO_2392 (O_2392,N_24568,N_24395);
nand UO_2393 (O_2393,N_24781,N_24399);
nor UO_2394 (O_2394,N_24546,N_24790);
xor UO_2395 (O_2395,N_24967,N_24912);
or UO_2396 (O_2396,N_24778,N_24954);
and UO_2397 (O_2397,N_24575,N_24736);
and UO_2398 (O_2398,N_24881,N_24396);
nand UO_2399 (O_2399,N_24444,N_24839);
nand UO_2400 (O_2400,N_24804,N_24409);
or UO_2401 (O_2401,N_24886,N_24642);
nand UO_2402 (O_2402,N_24735,N_24942);
and UO_2403 (O_2403,N_24825,N_24594);
nand UO_2404 (O_2404,N_24563,N_24581);
xnor UO_2405 (O_2405,N_24785,N_24562);
nor UO_2406 (O_2406,N_24468,N_24413);
nor UO_2407 (O_2407,N_24433,N_24722);
nand UO_2408 (O_2408,N_24460,N_24751);
or UO_2409 (O_2409,N_24642,N_24980);
nand UO_2410 (O_2410,N_24947,N_24744);
or UO_2411 (O_2411,N_24883,N_24776);
nor UO_2412 (O_2412,N_24468,N_24720);
xnor UO_2413 (O_2413,N_24721,N_24677);
xor UO_2414 (O_2414,N_24598,N_24758);
and UO_2415 (O_2415,N_24590,N_24682);
xor UO_2416 (O_2416,N_24526,N_24688);
and UO_2417 (O_2417,N_24624,N_24607);
or UO_2418 (O_2418,N_24929,N_24873);
or UO_2419 (O_2419,N_24764,N_24836);
or UO_2420 (O_2420,N_24531,N_24481);
nand UO_2421 (O_2421,N_24741,N_24565);
nor UO_2422 (O_2422,N_24949,N_24836);
xnor UO_2423 (O_2423,N_24428,N_24691);
nand UO_2424 (O_2424,N_24386,N_24849);
and UO_2425 (O_2425,N_24967,N_24651);
nand UO_2426 (O_2426,N_24408,N_24455);
and UO_2427 (O_2427,N_24677,N_24651);
nor UO_2428 (O_2428,N_24442,N_24573);
nand UO_2429 (O_2429,N_24649,N_24898);
nor UO_2430 (O_2430,N_24584,N_24434);
or UO_2431 (O_2431,N_24930,N_24793);
nand UO_2432 (O_2432,N_24855,N_24378);
nand UO_2433 (O_2433,N_24604,N_24795);
nor UO_2434 (O_2434,N_24570,N_24613);
nor UO_2435 (O_2435,N_24916,N_24721);
and UO_2436 (O_2436,N_24753,N_24839);
and UO_2437 (O_2437,N_24800,N_24556);
nor UO_2438 (O_2438,N_24876,N_24726);
or UO_2439 (O_2439,N_24676,N_24858);
and UO_2440 (O_2440,N_24515,N_24950);
and UO_2441 (O_2441,N_24486,N_24504);
xnor UO_2442 (O_2442,N_24544,N_24400);
or UO_2443 (O_2443,N_24724,N_24377);
or UO_2444 (O_2444,N_24826,N_24378);
and UO_2445 (O_2445,N_24711,N_24944);
xnor UO_2446 (O_2446,N_24628,N_24491);
or UO_2447 (O_2447,N_24886,N_24912);
nand UO_2448 (O_2448,N_24435,N_24534);
or UO_2449 (O_2449,N_24590,N_24937);
nand UO_2450 (O_2450,N_24886,N_24920);
xnor UO_2451 (O_2451,N_24794,N_24521);
and UO_2452 (O_2452,N_24687,N_24479);
and UO_2453 (O_2453,N_24469,N_24947);
or UO_2454 (O_2454,N_24986,N_24828);
nor UO_2455 (O_2455,N_24934,N_24740);
nand UO_2456 (O_2456,N_24455,N_24494);
xnor UO_2457 (O_2457,N_24440,N_24978);
nor UO_2458 (O_2458,N_24475,N_24646);
nand UO_2459 (O_2459,N_24803,N_24980);
and UO_2460 (O_2460,N_24733,N_24624);
and UO_2461 (O_2461,N_24451,N_24505);
nand UO_2462 (O_2462,N_24389,N_24796);
and UO_2463 (O_2463,N_24478,N_24991);
nand UO_2464 (O_2464,N_24760,N_24386);
nand UO_2465 (O_2465,N_24566,N_24695);
xor UO_2466 (O_2466,N_24511,N_24960);
xor UO_2467 (O_2467,N_24844,N_24847);
nor UO_2468 (O_2468,N_24809,N_24455);
nor UO_2469 (O_2469,N_24797,N_24876);
and UO_2470 (O_2470,N_24515,N_24999);
and UO_2471 (O_2471,N_24909,N_24675);
nand UO_2472 (O_2472,N_24998,N_24570);
and UO_2473 (O_2473,N_24462,N_24801);
or UO_2474 (O_2474,N_24435,N_24863);
or UO_2475 (O_2475,N_24670,N_24667);
nor UO_2476 (O_2476,N_24710,N_24690);
and UO_2477 (O_2477,N_24613,N_24533);
or UO_2478 (O_2478,N_24467,N_24532);
nor UO_2479 (O_2479,N_24623,N_24587);
or UO_2480 (O_2480,N_24791,N_24921);
or UO_2481 (O_2481,N_24945,N_24743);
nand UO_2482 (O_2482,N_24482,N_24833);
nand UO_2483 (O_2483,N_24387,N_24784);
and UO_2484 (O_2484,N_24823,N_24623);
nand UO_2485 (O_2485,N_24539,N_24866);
or UO_2486 (O_2486,N_24985,N_24585);
or UO_2487 (O_2487,N_24846,N_24607);
or UO_2488 (O_2488,N_24905,N_24446);
xnor UO_2489 (O_2489,N_24773,N_24499);
nor UO_2490 (O_2490,N_24955,N_24606);
nand UO_2491 (O_2491,N_24497,N_24614);
xor UO_2492 (O_2492,N_24552,N_24660);
nor UO_2493 (O_2493,N_24747,N_24531);
xnor UO_2494 (O_2494,N_24972,N_24916);
or UO_2495 (O_2495,N_24401,N_24724);
or UO_2496 (O_2496,N_24738,N_24840);
or UO_2497 (O_2497,N_24860,N_24498);
or UO_2498 (O_2498,N_24767,N_24587);
nand UO_2499 (O_2499,N_24641,N_24596);
xnor UO_2500 (O_2500,N_24477,N_24440);
xnor UO_2501 (O_2501,N_24438,N_24586);
or UO_2502 (O_2502,N_24649,N_24586);
xnor UO_2503 (O_2503,N_24405,N_24485);
or UO_2504 (O_2504,N_24841,N_24874);
and UO_2505 (O_2505,N_24825,N_24879);
xor UO_2506 (O_2506,N_24896,N_24444);
nor UO_2507 (O_2507,N_24476,N_24582);
and UO_2508 (O_2508,N_24378,N_24722);
xor UO_2509 (O_2509,N_24879,N_24865);
nand UO_2510 (O_2510,N_24730,N_24689);
nand UO_2511 (O_2511,N_24463,N_24899);
and UO_2512 (O_2512,N_24600,N_24499);
xnor UO_2513 (O_2513,N_24532,N_24426);
or UO_2514 (O_2514,N_24953,N_24524);
nand UO_2515 (O_2515,N_24396,N_24501);
nand UO_2516 (O_2516,N_24498,N_24849);
nand UO_2517 (O_2517,N_24584,N_24928);
xnor UO_2518 (O_2518,N_24528,N_24809);
nand UO_2519 (O_2519,N_24791,N_24685);
or UO_2520 (O_2520,N_24632,N_24463);
and UO_2521 (O_2521,N_24663,N_24489);
nand UO_2522 (O_2522,N_24765,N_24825);
nand UO_2523 (O_2523,N_24533,N_24482);
nor UO_2524 (O_2524,N_24511,N_24799);
and UO_2525 (O_2525,N_24580,N_24566);
nor UO_2526 (O_2526,N_24487,N_24803);
xor UO_2527 (O_2527,N_24443,N_24585);
nor UO_2528 (O_2528,N_24438,N_24461);
xor UO_2529 (O_2529,N_24999,N_24756);
nand UO_2530 (O_2530,N_24397,N_24792);
and UO_2531 (O_2531,N_24410,N_24400);
nand UO_2532 (O_2532,N_24931,N_24715);
nand UO_2533 (O_2533,N_24409,N_24791);
nand UO_2534 (O_2534,N_24695,N_24610);
or UO_2535 (O_2535,N_24430,N_24482);
nand UO_2536 (O_2536,N_24725,N_24733);
nand UO_2537 (O_2537,N_24973,N_24547);
nor UO_2538 (O_2538,N_24988,N_24723);
or UO_2539 (O_2539,N_24910,N_24953);
nand UO_2540 (O_2540,N_24832,N_24564);
xor UO_2541 (O_2541,N_24840,N_24806);
nor UO_2542 (O_2542,N_24503,N_24632);
and UO_2543 (O_2543,N_24428,N_24614);
nand UO_2544 (O_2544,N_24675,N_24628);
or UO_2545 (O_2545,N_24436,N_24650);
xnor UO_2546 (O_2546,N_24708,N_24796);
and UO_2547 (O_2547,N_24566,N_24606);
nor UO_2548 (O_2548,N_24643,N_24563);
or UO_2549 (O_2549,N_24855,N_24938);
nand UO_2550 (O_2550,N_24835,N_24790);
nor UO_2551 (O_2551,N_24526,N_24720);
nor UO_2552 (O_2552,N_24528,N_24959);
xor UO_2553 (O_2553,N_24951,N_24613);
nor UO_2554 (O_2554,N_24377,N_24710);
or UO_2555 (O_2555,N_24826,N_24436);
nand UO_2556 (O_2556,N_24861,N_24917);
nor UO_2557 (O_2557,N_24757,N_24484);
and UO_2558 (O_2558,N_24949,N_24952);
or UO_2559 (O_2559,N_24679,N_24808);
xor UO_2560 (O_2560,N_24790,N_24702);
or UO_2561 (O_2561,N_24589,N_24826);
and UO_2562 (O_2562,N_24841,N_24963);
or UO_2563 (O_2563,N_24721,N_24558);
or UO_2564 (O_2564,N_24824,N_24462);
xnor UO_2565 (O_2565,N_24556,N_24612);
or UO_2566 (O_2566,N_24653,N_24475);
or UO_2567 (O_2567,N_24832,N_24680);
nand UO_2568 (O_2568,N_24630,N_24773);
nor UO_2569 (O_2569,N_24719,N_24811);
or UO_2570 (O_2570,N_24633,N_24394);
or UO_2571 (O_2571,N_24511,N_24622);
and UO_2572 (O_2572,N_24392,N_24460);
nor UO_2573 (O_2573,N_24560,N_24476);
nor UO_2574 (O_2574,N_24513,N_24727);
xnor UO_2575 (O_2575,N_24685,N_24561);
nor UO_2576 (O_2576,N_24941,N_24749);
nand UO_2577 (O_2577,N_24618,N_24784);
nand UO_2578 (O_2578,N_24720,N_24690);
nor UO_2579 (O_2579,N_24424,N_24692);
or UO_2580 (O_2580,N_24401,N_24929);
xnor UO_2581 (O_2581,N_24789,N_24378);
xor UO_2582 (O_2582,N_24775,N_24967);
nor UO_2583 (O_2583,N_24491,N_24669);
nor UO_2584 (O_2584,N_24478,N_24979);
or UO_2585 (O_2585,N_24586,N_24489);
xor UO_2586 (O_2586,N_24866,N_24626);
or UO_2587 (O_2587,N_24553,N_24757);
and UO_2588 (O_2588,N_24913,N_24659);
and UO_2589 (O_2589,N_24490,N_24986);
nor UO_2590 (O_2590,N_24463,N_24824);
xor UO_2591 (O_2591,N_24621,N_24714);
and UO_2592 (O_2592,N_24933,N_24600);
or UO_2593 (O_2593,N_24971,N_24885);
nand UO_2594 (O_2594,N_24594,N_24413);
or UO_2595 (O_2595,N_24663,N_24889);
xor UO_2596 (O_2596,N_24629,N_24381);
or UO_2597 (O_2597,N_24733,N_24689);
nand UO_2598 (O_2598,N_24903,N_24482);
and UO_2599 (O_2599,N_24864,N_24415);
nor UO_2600 (O_2600,N_24817,N_24637);
or UO_2601 (O_2601,N_24922,N_24889);
nor UO_2602 (O_2602,N_24410,N_24600);
nand UO_2603 (O_2603,N_24843,N_24379);
and UO_2604 (O_2604,N_24471,N_24732);
nand UO_2605 (O_2605,N_24676,N_24797);
and UO_2606 (O_2606,N_24875,N_24506);
nand UO_2607 (O_2607,N_24456,N_24831);
and UO_2608 (O_2608,N_24449,N_24920);
nand UO_2609 (O_2609,N_24762,N_24521);
xnor UO_2610 (O_2610,N_24855,N_24716);
or UO_2611 (O_2611,N_24795,N_24953);
nand UO_2612 (O_2612,N_24737,N_24525);
or UO_2613 (O_2613,N_24872,N_24783);
and UO_2614 (O_2614,N_24613,N_24683);
xor UO_2615 (O_2615,N_24583,N_24628);
nor UO_2616 (O_2616,N_24638,N_24956);
and UO_2617 (O_2617,N_24778,N_24549);
nand UO_2618 (O_2618,N_24695,N_24739);
nand UO_2619 (O_2619,N_24807,N_24929);
nor UO_2620 (O_2620,N_24783,N_24782);
and UO_2621 (O_2621,N_24411,N_24435);
xnor UO_2622 (O_2622,N_24480,N_24440);
nor UO_2623 (O_2623,N_24604,N_24639);
xor UO_2624 (O_2624,N_24784,N_24463);
and UO_2625 (O_2625,N_24411,N_24547);
and UO_2626 (O_2626,N_24764,N_24460);
xnor UO_2627 (O_2627,N_24820,N_24919);
xnor UO_2628 (O_2628,N_24937,N_24865);
nor UO_2629 (O_2629,N_24505,N_24438);
and UO_2630 (O_2630,N_24754,N_24843);
xor UO_2631 (O_2631,N_24818,N_24883);
and UO_2632 (O_2632,N_24950,N_24562);
nor UO_2633 (O_2633,N_24466,N_24579);
and UO_2634 (O_2634,N_24400,N_24457);
xnor UO_2635 (O_2635,N_24867,N_24864);
nor UO_2636 (O_2636,N_24454,N_24824);
and UO_2637 (O_2637,N_24884,N_24832);
xnor UO_2638 (O_2638,N_24512,N_24771);
nand UO_2639 (O_2639,N_24833,N_24822);
xor UO_2640 (O_2640,N_24799,N_24453);
xnor UO_2641 (O_2641,N_24920,N_24833);
nor UO_2642 (O_2642,N_24701,N_24401);
xnor UO_2643 (O_2643,N_24537,N_24408);
xnor UO_2644 (O_2644,N_24518,N_24773);
nand UO_2645 (O_2645,N_24961,N_24761);
xor UO_2646 (O_2646,N_24678,N_24978);
nand UO_2647 (O_2647,N_24909,N_24733);
nand UO_2648 (O_2648,N_24428,N_24862);
and UO_2649 (O_2649,N_24504,N_24578);
or UO_2650 (O_2650,N_24640,N_24494);
nor UO_2651 (O_2651,N_24790,N_24628);
and UO_2652 (O_2652,N_24961,N_24598);
nor UO_2653 (O_2653,N_24695,N_24678);
or UO_2654 (O_2654,N_24620,N_24402);
xor UO_2655 (O_2655,N_24443,N_24888);
nor UO_2656 (O_2656,N_24600,N_24541);
nor UO_2657 (O_2657,N_24587,N_24737);
xnor UO_2658 (O_2658,N_24642,N_24576);
nand UO_2659 (O_2659,N_24922,N_24864);
and UO_2660 (O_2660,N_24983,N_24815);
and UO_2661 (O_2661,N_24937,N_24398);
nand UO_2662 (O_2662,N_24905,N_24721);
xnor UO_2663 (O_2663,N_24963,N_24391);
nor UO_2664 (O_2664,N_24393,N_24852);
xnor UO_2665 (O_2665,N_24815,N_24817);
xor UO_2666 (O_2666,N_24635,N_24450);
nor UO_2667 (O_2667,N_24553,N_24643);
nor UO_2668 (O_2668,N_24376,N_24761);
nand UO_2669 (O_2669,N_24843,N_24988);
nor UO_2670 (O_2670,N_24468,N_24402);
or UO_2671 (O_2671,N_24765,N_24882);
or UO_2672 (O_2672,N_24582,N_24483);
and UO_2673 (O_2673,N_24512,N_24902);
or UO_2674 (O_2674,N_24943,N_24697);
xor UO_2675 (O_2675,N_24713,N_24736);
nand UO_2676 (O_2676,N_24946,N_24792);
nand UO_2677 (O_2677,N_24671,N_24531);
nor UO_2678 (O_2678,N_24887,N_24782);
and UO_2679 (O_2679,N_24505,N_24405);
xnor UO_2680 (O_2680,N_24544,N_24437);
nor UO_2681 (O_2681,N_24922,N_24628);
nor UO_2682 (O_2682,N_24863,N_24706);
nor UO_2683 (O_2683,N_24524,N_24423);
nor UO_2684 (O_2684,N_24733,N_24968);
nor UO_2685 (O_2685,N_24494,N_24807);
and UO_2686 (O_2686,N_24675,N_24673);
and UO_2687 (O_2687,N_24421,N_24724);
nor UO_2688 (O_2688,N_24383,N_24474);
nand UO_2689 (O_2689,N_24506,N_24740);
and UO_2690 (O_2690,N_24825,N_24652);
nor UO_2691 (O_2691,N_24492,N_24451);
nand UO_2692 (O_2692,N_24597,N_24466);
nor UO_2693 (O_2693,N_24442,N_24699);
or UO_2694 (O_2694,N_24473,N_24808);
or UO_2695 (O_2695,N_24649,N_24816);
nor UO_2696 (O_2696,N_24543,N_24468);
and UO_2697 (O_2697,N_24995,N_24801);
xnor UO_2698 (O_2698,N_24479,N_24594);
nand UO_2699 (O_2699,N_24641,N_24963);
nor UO_2700 (O_2700,N_24503,N_24822);
nor UO_2701 (O_2701,N_24756,N_24569);
or UO_2702 (O_2702,N_24417,N_24600);
xnor UO_2703 (O_2703,N_24724,N_24568);
or UO_2704 (O_2704,N_24518,N_24734);
nand UO_2705 (O_2705,N_24604,N_24403);
and UO_2706 (O_2706,N_24627,N_24432);
xor UO_2707 (O_2707,N_24881,N_24666);
nor UO_2708 (O_2708,N_24673,N_24653);
nand UO_2709 (O_2709,N_24566,N_24852);
nor UO_2710 (O_2710,N_24567,N_24866);
nor UO_2711 (O_2711,N_24744,N_24577);
xor UO_2712 (O_2712,N_24762,N_24984);
nor UO_2713 (O_2713,N_24635,N_24799);
or UO_2714 (O_2714,N_24633,N_24934);
and UO_2715 (O_2715,N_24481,N_24933);
xor UO_2716 (O_2716,N_24797,N_24605);
and UO_2717 (O_2717,N_24381,N_24497);
xnor UO_2718 (O_2718,N_24599,N_24775);
nand UO_2719 (O_2719,N_24474,N_24403);
or UO_2720 (O_2720,N_24431,N_24886);
nor UO_2721 (O_2721,N_24544,N_24953);
xnor UO_2722 (O_2722,N_24394,N_24590);
or UO_2723 (O_2723,N_24809,N_24955);
nand UO_2724 (O_2724,N_24732,N_24796);
nor UO_2725 (O_2725,N_24721,N_24794);
nor UO_2726 (O_2726,N_24847,N_24738);
or UO_2727 (O_2727,N_24541,N_24721);
or UO_2728 (O_2728,N_24909,N_24965);
xor UO_2729 (O_2729,N_24557,N_24497);
nor UO_2730 (O_2730,N_24679,N_24535);
or UO_2731 (O_2731,N_24830,N_24724);
xor UO_2732 (O_2732,N_24816,N_24730);
and UO_2733 (O_2733,N_24481,N_24967);
nor UO_2734 (O_2734,N_24791,N_24594);
xor UO_2735 (O_2735,N_24619,N_24422);
and UO_2736 (O_2736,N_24558,N_24968);
or UO_2737 (O_2737,N_24842,N_24996);
xnor UO_2738 (O_2738,N_24833,N_24472);
and UO_2739 (O_2739,N_24467,N_24651);
and UO_2740 (O_2740,N_24485,N_24880);
or UO_2741 (O_2741,N_24972,N_24462);
xor UO_2742 (O_2742,N_24951,N_24690);
nor UO_2743 (O_2743,N_24952,N_24640);
xor UO_2744 (O_2744,N_24664,N_24861);
xor UO_2745 (O_2745,N_24818,N_24505);
and UO_2746 (O_2746,N_24417,N_24572);
xor UO_2747 (O_2747,N_24449,N_24827);
or UO_2748 (O_2748,N_24816,N_24453);
nor UO_2749 (O_2749,N_24537,N_24889);
or UO_2750 (O_2750,N_24863,N_24837);
nand UO_2751 (O_2751,N_24796,N_24698);
nor UO_2752 (O_2752,N_24688,N_24901);
xor UO_2753 (O_2753,N_24531,N_24758);
nor UO_2754 (O_2754,N_24866,N_24521);
nor UO_2755 (O_2755,N_24674,N_24713);
nor UO_2756 (O_2756,N_24716,N_24383);
nand UO_2757 (O_2757,N_24634,N_24830);
nand UO_2758 (O_2758,N_24908,N_24590);
xor UO_2759 (O_2759,N_24703,N_24517);
or UO_2760 (O_2760,N_24515,N_24459);
nor UO_2761 (O_2761,N_24591,N_24961);
nor UO_2762 (O_2762,N_24784,N_24445);
or UO_2763 (O_2763,N_24626,N_24476);
xor UO_2764 (O_2764,N_24479,N_24987);
and UO_2765 (O_2765,N_24748,N_24824);
nand UO_2766 (O_2766,N_24663,N_24463);
nor UO_2767 (O_2767,N_24623,N_24602);
xor UO_2768 (O_2768,N_24841,N_24816);
and UO_2769 (O_2769,N_24710,N_24433);
and UO_2770 (O_2770,N_24695,N_24565);
xnor UO_2771 (O_2771,N_24686,N_24759);
nand UO_2772 (O_2772,N_24481,N_24390);
nand UO_2773 (O_2773,N_24584,N_24419);
or UO_2774 (O_2774,N_24585,N_24690);
xor UO_2775 (O_2775,N_24987,N_24911);
nand UO_2776 (O_2776,N_24769,N_24504);
nand UO_2777 (O_2777,N_24825,N_24679);
nor UO_2778 (O_2778,N_24487,N_24825);
or UO_2779 (O_2779,N_24890,N_24848);
xor UO_2780 (O_2780,N_24472,N_24797);
or UO_2781 (O_2781,N_24788,N_24874);
and UO_2782 (O_2782,N_24928,N_24889);
xnor UO_2783 (O_2783,N_24828,N_24816);
nor UO_2784 (O_2784,N_24524,N_24974);
nand UO_2785 (O_2785,N_24628,N_24830);
nor UO_2786 (O_2786,N_24963,N_24724);
xor UO_2787 (O_2787,N_24403,N_24410);
nand UO_2788 (O_2788,N_24919,N_24708);
nand UO_2789 (O_2789,N_24770,N_24529);
xor UO_2790 (O_2790,N_24580,N_24961);
xor UO_2791 (O_2791,N_24512,N_24850);
or UO_2792 (O_2792,N_24433,N_24528);
and UO_2793 (O_2793,N_24876,N_24714);
xor UO_2794 (O_2794,N_24979,N_24653);
xnor UO_2795 (O_2795,N_24871,N_24395);
xnor UO_2796 (O_2796,N_24704,N_24495);
or UO_2797 (O_2797,N_24936,N_24633);
nor UO_2798 (O_2798,N_24764,N_24498);
or UO_2799 (O_2799,N_24508,N_24460);
xnor UO_2800 (O_2800,N_24684,N_24525);
nor UO_2801 (O_2801,N_24438,N_24454);
nor UO_2802 (O_2802,N_24723,N_24900);
nor UO_2803 (O_2803,N_24641,N_24607);
nor UO_2804 (O_2804,N_24936,N_24995);
or UO_2805 (O_2805,N_24972,N_24554);
nor UO_2806 (O_2806,N_24866,N_24542);
and UO_2807 (O_2807,N_24956,N_24816);
and UO_2808 (O_2808,N_24473,N_24833);
or UO_2809 (O_2809,N_24919,N_24481);
or UO_2810 (O_2810,N_24488,N_24934);
xor UO_2811 (O_2811,N_24399,N_24839);
nor UO_2812 (O_2812,N_24658,N_24766);
xor UO_2813 (O_2813,N_24599,N_24423);
nor UO_2814 (O_2814,N_24425,N_24933);
nand UO_2815 (O_2815,N_24906,N_24665);
or UO_2816 (O_2816,N_24897,N_24378);
or UO_2817 (O_2817,N_24454,N_24822);
and UO_2818 (O_2818,N_24384,N_24948);
nor UO_2819 (O_2819,N_24810,N_24471);
xnor UO_2820 (O_2820,N_24385,N_24838);
nor UO_2821 (O_2821,N_24805,N_24686);
and UO_2822 (O_2822,N_24451,N_24631);
and UO_2823 (O_2823,N_24765,N_24994);
nor UO_2824 (O_2824,N_24568,N_24877);
nor UO_2825 (O_2825,N_24914,N_24901);
or UO_2826 (O_2826,N_24904,N_24403);
nand UO_2827 (O_2827,N_24840,N_24827);
nand UO_2828 (O_2828,N_24483,N_24615);
nor UO_2829 (O_2829,N_24920,N_24587);
or UO_2830 (O_2830,N_24501,N_24630);
or UO_2831 (O_2831,N_24997,N_24669);
xor UO_2832 (O_2832,N_24914,N_24579);
xnor UO_2833 (O_2833,N_24748,N_24974);
nand UO_2834 (O_2834,N_24441,N_24960);
nand UO_2835 (O_2835,N_24646,N_24659);
nand UO_2836 (O_2836,N_24765,N_24834);
nand UO_2837 (O_2837,N_24884,N_24898);
or UO_2838 (O_2838,N_24743,N_24656);
and UO_2839 (O_2839,N_24442,N_24915);
or UO_2840 (O_2840,N_24553,N_24613);
and UO_2841 (O_2841,N_24500,N_24603);
or UO_2842 (O_2842,N_24981,N_24887);
nor UO_2843 (O_2843,N_24993,N_24444);
or UO_2844 (O_2844,N_24679,N_24455);
nor UO_2845 (O_2845,N_24399,N_24732);
nor UO_2846 (O_2846,N_24541,N_24691);
nand UO_2847 (O_2847,N_24632,N_24908);
or UO_2848 (O_2848,N_24723,N_24510);
or UO_2849 (O_2849,N_24772,N_24802);
or UO_2850 (O_2850,N_24977,N_24888);
nor UO_2851 (O_2851,N_24473,N_24479);
nor UO_2852 (O_2852,N_24488,N_24654);
and UO_2853 (O_2853,N_24420,N_24847);
nand UO_2854 (O_2854,N_24925,N_24436);
nor UO_2855 (O_2855,N_24788,N_24376);
nor UO_2856 (O_2856,N_24430,N_24711);
xor UO_2857 (O_2857,N_24464,N_24969);
xor UO_2858 (O_2858,N_24593,N_24803);
and UO_2859 (O_2859,N_24456,N_24784);
nor UO_2860 (O_2860,N_24686,N_24849);
nor UO_2861 (O_2861,N_24470,N_24830);
nor UO_2862 (O_2862,N_24498,N_24689);
or UO_2863 (O_2863,N_24877,N_24905);
nor UO_2864 (O_2864,N_24767,N_24531);
or UO_2865 (O_2865,N_24836,N_24656);
nor UO_2866 (O_2866,N_24755,N_24945);
nor UO_2867 (O_2867,N_24583,N_24497);
nor UO_2868 (O_2868,N_24970,N_24753);
nor UO_2869 (O_2869,N_24907,N_24669);
xnor UO_2870 (O_2870,N_24706,N_24787);
or UO_2871 (O_2871,N_24779,N_24762);
or UO_2872 (O_2872,N_24532,N_24599);
nand UO_2873 (O_2873,N_24824,N_24805);
nand UO_2874 (O_2874,N_24707,N_24801);
nor UO_2875 (O_2875,N_24986,N_24539);
or UO_2876 (O_2876,N_24402,N_24790);
nor UO_2877 (O_2877,N_24430,N_24842);
and UO_2878 (O_2878,N_24651,N_24940);
or UO_2879 (O_2879,N_24926,N_24585);
xor UO_2880 (O_2880,N_24502,N_24644);
xnor UO_2881 (O_2881,N_24781,N_24538);
xor UO_2882 (O_2882,N_24533,N_24858);
nor UO_2883 (O_2883,N_24891,N_24423);
xnor UO_2884 (O_2884,N_24925,N_24413);
and UO_2885 (O_2885,N_24991,N_24573);
or UO_2886 (O_2886,N_24414,N_24920);
and UO_2887 (O_2887,N_24450,N_24878);
or UO_2888 (O_2888,N_24795,N_24778);
xor UO_2889 (O_2889,N_24988,N_24778);
nor UO_2890 (O_2890,N_24610,N_24853);
or UO_2891 (O_2891,N_24605,N_24518);
xor UO_2892 (O_2892,N_24950,N_24437);
xnor UO_2893 (O_2893,N_24893,N_24918);
and UO_2894 (O_2894,N_24932,N_24781);
or UO_2895 (O_2895,N_24703,N_24974);
or UO_2896 (O_2896,N_24442,N_24682);
and UO_2897 (O_2897,N_24871,N_24765);
xnor UO_2898 (O_2898,N_24860,N_24438);
xor UO_2899 (O_2899,N_24847,N_24395);
and UO_2900 (O_2900,N_24434,N_24464);
or UO_2901 (O_2901,N_24527,N_24763);
nand UO_2902 (O_2902,N_24787,N_24552);
xor UO_2903 (O_2903,N_24912,N_24732);
xor UO_2904 (O_2904,N_24758,N_24846);
and UO_2905 (O_2905,N_24672,N_24697);
nor UO_2906 (O_2906,N_24688,N_24927);
or UO_2907 (O_2907,N_24690,N_24640);
nor UO_2908 (O_2908,N_24986,N_24399);
and UO_2909 (O_2909,N_24660,N_24827);
or UO_2910 (O_2910,N_24478,N_24510);
and UO_2911 (O_2911,N_24870,N_24815);
and UO_2912 (O_2912,N_24506,N_24849);
xnor UO_2913 (O_2913,N_24924,N_24740);
and UO_2914 (O_2914,N_24733,N_24838);
nand UO_2915 (O_2915,N_24691,N_24887);
nor UO_2916 (O_2916,N_24856,N_24772);
and UO_2917 (O_2917,N_24989,N_24848);
nor UO_2918 (O_2918,N_24894,N_24468);
nand UO_2919 (O_2919,N_24453,N_24621);
nor UO_2920 (O_2920,N_24766,N_24552);
nand UO_2921 (O_2921,N_24697,N_24888);
or UO_2922 (O_2922,N_24549,N_24418);
or UO_2923 (O_2923,N_24576,N_24871);
or UO_2924 (O_2924,N_24762,N_24883);
nand UO_2925 (O_2925,N_24519,N_24577);
or UO_2926 (O_2926,N_24496,N_24474);
xor UO_2927 (O_2927,N_24529,N_24971);
nor UO_2928 (O_2928,N_24645,N_24885);
xnor UO_2929 (O_2929,N_24845,N_24907);
nor UO_2930 (O_2930,N_24515,N_24641);
xor UO_2931 (O_2931,N_24816,N_24698);
or UO_2932 (O_2932,N_24639,N_24698);
or UO_2933 (O_2933,N_24691,N_24399);
nor UO_2934 (O_2934,N_24958,N_24822);
or UO_2935 (O_2935,N_24639,N_24691);
nand UO_2936 (O_2936,N_24381,N_24957);
or UO_2937 (O_2937,N_24488,N_24815);
xor UO_2938 (O_2938,N_24434,N_24387);
and UO_2939 (O_2939,N_24394,N_24383);
xor UO_2940 (O_2940,N_24827,N_24887);
xor UO_2941 (O_2941,N_24863,N_24963);
nand UO_2942 (O_2942,N_24469,N_24786);
and UO_2943 (O_2943,N_24648,N_24681);
or UO_2944 (O_2944,N_24514,N_24656);
or UO_2945 (O_2945,N_24994,N_24520);
xor UO_2946 (O_2946,N_24536,N_24558);
or UO_2947 (O_2947,N_24451,N_24646);
nand UO_2948 (O_2948,N_24889,N_24672);
or UO_2949 (O_2949,N_24645,N_24469);
xnor UO_2950 (O_2950,N_24790,N_24910);
and UO_2951 (O_2951,N_24957,N_24509);
nor UO_2952 (O_2952,N_24698,N_24715);
or UO_2953 (O_2953,N_24499,N_24942);
or UO_2954 (O_2954,N_24937,N_24570);
nand UO_2955 (O_2955,N_24461,N_24602);
nand UO_2956 (O_2956,N_24951,N_24410);
nor UO_2957 (O_2957,N_24705,N_24554);
or UO_2958 (O_2958,N_24804,N_24479);
nor UO_2959 (O_2959,N_24687,N_24973);
or UO_2960 (O_2960,N_24498,N_24963);
xor UO_2961 (O_2961,N_24486,N_24873);
nor UO_2962 (O_2962,N_24928,N_24820);
or UO_2963 (O_2963,N_24500,N_24568);
xnor UO_2964 (O_2964,N_24833,N_24853);
nand UO_2965 (O_2965,N_24434,N_24948);
nor UO_2966 (O_2966,N_24789,N_24411);
or UO_2967 (O_2967,N_24523,N_24775);
nand UO_2968 (O_2968,N_24717,N_24709);
nand UO_2969 (O_2969,N_24771,N_24827);
nor UO_2970 (O_2970,N_24643,N_24677);
nand UO_2971 (O_2971,N_24625,N_24783);
nor UO_2972 (O_2972,N_24765,N_24881);
nor UO_2973 (O_2973,N_24714,N_24504);
nor UO_2974 (O_2974,N_24664,N_24407);
nand UO_2975 (O_2975,N_24604,N_24630);
and UO_2976 (O_2976,N_24509,N_24714);
xor UO_2977 (O_2977,N_24520,N_24410);
xnor UO_2978 (O_2978,N_24736,N_24968);
xor UO_2979 (O_2979,N_24978,N_24984);
nor UO_2980 (O_2980,N_24796,N_24866);
nand UO_2981 (O_2981,N_24415,N_24447);
xor UO_2982 (O_2982,N_24872,N_24428);
xor UO_2983 (O_2983,N_24735,N_24450);
nor UO_2984 (O_2984,N_24944,N_24612);
nor UO_2985 (O_2985,N_24662,N_24468);
and UO_2986 (O_2986,N_24879,N_24962);
and UO_2987 (O_2987,N_24690,N_24608);
nand UO_2988 (O_2988,N_24908,N_24576);
nand UO_2989 (O_2989,N_24670,N_24540);
nand UO_2990 (O_2990,N_24504,N_24723);
and UO_2991 (O_2991,N_24645,N_24623);
xor UO_2992 (O_2992,N_24621,N_24899);
xor UO_2993 (O_2993,N_24553,N_24527);
or UO_2994 (O_2994,N_24946,N_24999);
nor UO_2995 (O_2995,N_24403,N_24514);
nor UO_2996 (O_2996,N_24565,N_24707);
xnor UO_2997 (O_2997,N_24958,N_24925);
nand UO_2998 (O_2998,N_24662,N_24963);
or UO_2999 (O_2999,N_24420,N_24745);
endmodule