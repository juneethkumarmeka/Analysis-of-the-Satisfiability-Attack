module basic_500_3000_500_4_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_295,In_265);
and U1 (N_1,In_442,In_241);
nor U2 (N_2,In_110,In_269);
or U3 (N_3,In_1,In_456);
and U4 (N_4,In_106,In_229);
xnor U5 (N_5,In_323,In_400);
nand U6 (N_6,In_471,In_118);
or U7 (N_7,In_416,In_22);
nand U8 (N_8,In_155,In_148);
nand U9 (N_9,In_117,In_112);
nand U10 (N_10,In_313,In_324);
nor U11 (N_11,In_177,In_13);
and U12 (N_12,In_250,In_429);
nand U13 (N_13,In_386,In_368);
nor U14 (N_14,In_35,In_174);
nor U15 (N_15,In_122,In_40);
nor U16 (N_16,In_84,In_453);
nand U17 (N_17,In_365,In_343);
or U18 (N_18,In_337,In_163);
or U19 (N_19,In_485,In_496);
and U20 (N_20,In_403,In_32);
or U21 (N_21,In_16,In_289);
nand U22 (N_22,In_55,In_82);
xnor U23 (N_23,In_192,In_385);
or U24 (N_24,In_433,In_204);
nand U25 (N_25,In_53,In_396);
nand U26 (N_26,In_72,In_197);
xnor U27 (N_27,In_256,In_320);
nand U28 (N_28,In_212,In_46);
nor U29 (N_29,In_316,In_460);
xor U30 (N_30,In_44,In_478);
or U31 (N_31,In_57,In_394);
nand U32 (N_32,In_183,In_131);
nor U33 (N_33,In_397,In_448);
nand U34 (N_34,In_211,In_205);
or U35 (N_35,In_186,In_24);
nand U36 (N_36,In_62,In_327);
and U37 (N_37,In_65,In_435);
or U38 (N_38,In_291,In_227);
nor U39 (N_39,In_206,In_367);
and U40 (N_40,In_251,In_281);
nand U41 (N_41,In_98,In_428);
nor U42 (N_42,In_200,In_372);
and U43 (N_43,In_263,In_321);
or U44 (N_44,In_102,In_481);
nor U45 (N_45,In_271,In_482);
or U46 (N_46,In_120,In_355);
or U47 (N_47,In_52,In_173);
nor U48 (N_48,In_449,In_28);
nand U49 (N_49,In_363,In_258);
and U50 (N_50,In_59,In_463);
or U51 (N_51,In_38,In_391);
nand U52 (N_52,In_268,In_259);
and U53 (N_53,In_243,In_114);
or U54 (N_54,In_199,In_290);
nor U55 (N_55,In_116,In_127);
nor U56 (N_56,In_375,In_308);
nor U57 (N_57,In_349,In_447);
or U58 (N_58,In_401,In_137);
xnor U59 (N_59,In_325,In_66);
or U60 (N_60,In_472,In_408);
nand U61 (N_61,In_350,In_220);
xnor U62 (N_62,In_392,In_474);
or U63 (N_63,In_79,In_415);
nand U64 (N_64,In_270,In_411);
nand U65 (N_65,In_412,In_348);
and U66 (N_66,In_314,In_73);
nor U67 (N_67,In_339,In_261);
and U68 (N_68,In_253,In_432);
or U69 (N_69,In_461,In_154);
and U70 (N_70,In_37,In_125);
nand U71 (N_71,In_364,In_172);
or U72 (N_72,In_376,In_115);
nand U73 (N_73,In_425,In_446);
or U74 (N_74,In_484,In_92);
and U75 (N_75,In_285,In_280);
nand U76 (N_76,In_132,In_277);
nor U77 (N_77,In_360,In_91);
nor U78 (N_78,In_25,In_344);
nor U79 (N_79,In_146,In_342);
or U80 (N_80,In_382,In_31);
xor U81 (N_81,In_233,In_336);
nand U82 (N_82,In_3,In_123);
nand U83 (N_83,In_443,In_498);
nand U84 (N_84,In_185,In_202);
or U85 (N_85,In_189,In_218);
nand U86 (N_86,In_414,In_18);
nor U87 (N_87,In_440,In_108);
xor U88 (N_88,In_109,In_143);
nor U89 (N_89,In_30,In_333);
nand U90 (N_90,In_225,In_399);
nor U91 (N_91,In_99,In_36);
nand U92 (N_92,In_21,In_222);
nand U93 (N_93,In_119,In_499);
nand U94 (N_94,In_68,In_83);
nand U95 (N_95,In_398,In_352);
nor U96 (N_96,In_39,In_464);
and U97 (N_97,In_113,In_240);
nand U98 (N_98,In_335,In_100);
and U99 (N_99,In_10,In_315);
nor U100 (N_100,In_492,In_423);
nor U101 (N_101,In_244,In_356);
and U102 (N_102,In_495,In_95);
nor U103 (N_103,In_147,In_158);
and U104 (N_104,In_34,In_266);
or U105 (N_105,In_418,In_319);
nor U106 (N_106,In_296,In_353);
xor U107 (N_107,In_462,In_152);
nand U108 (N_108,In_341,In_175);
and U109 (N_109,In_145,In_41);
nor U110 (N_110,In_300,In_284);
or U111 (N_111,In_167,In_219);
xor U112 (N_112,In_383,In_331);
or U113 (N_113,In_63,In_420);
or U114 (N_114,In_469,In_402);
nand U115 (N_115,In_198,In_326);
nand U116 (N_116,In_215,In_139);
and U117 (N_117,In_23,In_171);
or U118 (N_118,In_209,In_178);
and U119 (N_119,In_20,In_43);
or U120 (N_120,In_441,In_351);
or U121 (N_121,In_362,In_239);
or U122 (N_122,In_480,In_287);
xor U123 (N_123,In_278,In_151);
nor U124 (N_124,In_2,In_165);
nand U125 (N_125,In_201,In_304);
nor U126 (N_126,In_404,In_149);
and U127 (N_127,In_479,In_427);
nor U128 (N_128,In_217,In_431);
xor U129 (N_129,In_288,In_150);
nor U130 (N_130,In_87,In_221);
or U131 (N_131,In_128,In_332);
or U132 (N_132,In_179,In_208);
and U133 (N_133,In_242,In_377);
or U134 (N_134,In_48,In_69);
or U135 (N_135,In_370,In_465);
or U136 (N_136,In_235,In_224);
and U137 (N_137,In_407,In_387);
and U138 (N_138,In_193,In_359);
nor U139 (N_139,In_14,In_54);
nor U140 (N_140,In_161,In_76);
and U141 (N_141,In_417,In_168);
nor U142 (N_142,In_329,In_490);
nor U143 (N_143,In_70,In_267);
xnor U144 (N_144,In_390,In_111);
nor U145 (N_145,In_11,In_466);
or U146 (N_146,In_101,In_283);
nand U147 (N_147,In_67,In_153);
or U148 (N_148,In_473,In_434);
nand U149 (N_149,In_5,In_389);
or U150 (N_150,In_236,In_15);
and U151 (N_151,In_6,In_384);
nor U152 (N_152,In_366,In_121);
or U153 (N_153,In_438,In_156);
nor U154 (N_154,In_80,In_157);
or U155 (N_155,In_190,In_4);
nor U156 (N_156,In_56,In_105);
nand U157 (N_157,In_477,In_223);
nand U158 (N_158,In_107,In_488);
nand U159 (N_159,In_475,In_421);
xnor U160 (N_160,In_140,In_406);
nand U161 (N_161,In_395,In_164);
nand U162 (N_162,In_104,In_302);
nor U163 (N_163,In_237,In_292);
nand U164 (N_164,In_180,In_493);
or U165 (N_165,In_60,In_388);
nor U166 (N_166,In_459,In_486);
xor U167 (N_167,In_97,In_470);
nor U168 (N_168,In_454,In_358);
and U169 (N_169,In_245,In_124);
xor U170 (N_170,In_293,In_306);
and U171 (N_171,In_338,In_182);
and U172 (N_172,In_188,In_135);
nand U173 (N_173,In_136,In_159);
or U174 (N_174,In_216,In_297);
nor U175 (N_175,In_468,In_71);
nand U176 (N_176,In_176,In_86);
and U177 (N_177,In_238,In_317);
nand U178 (N_178,In_340,In_228);
or U179 (N_179,In_45,In_90);
xnor U180 (N_180,In_181,In_103);
and U181 (N_181,In_357,In_361);
or U182 (N_182,In_298,In_94);
or U183 (N_183,In_187,In_138);
or U184 (N_184,In_378,In_89);
nor U185 (N_185,In_294,In_279);
and U186 (N_186,In_444,In_272);
xnor U187 (N_187,In_234,In_78);
and U188 (N_188,In_330,In_7);
or U189 (N_189,In_42,In_195);
nand U190 (N_190,In_214,In_276);
nand U191 (N_191,In_9,In_213);
and U192 (N_192,In_318,In_12);
xnor U193 (N_193,In_450,In_409);
xnor U194 (N_194,In_457,In_437);
nand U195 (N_195,In_51,In_303);
nand U196 (N_196,In_50,In_322);
or U197 (N_197,In_286,In_452);
nor U198 (N_198,In_422,In_191);
xor U199 (N_199,In_371,In_166);
and U200 (N_200,In_184,In_93);
nor U201 (N_201,In_489,In_369);
nand U202 (N_202,In_451,In_194);
nor U203 (N_203,In_196,In_130);
or U204 (N_204,In_81,In_307);
nor U205 (N_205,In_476,In_75);
and U206 (N_206,In_346,In_405);
nand U207 (N_207,In_64,In_410);
and U208 (N_208,In_203,In_483);
xnor U209 (N_209,In_129,In_230);
nor U210 (N_210,In_419,In_299);
nand U211 (N_211,In_273,In_497);
nand U212 (N_212,In_257,In_458);
or U213 (N_213,In_430,In_162);
and U214 (N_214,In_17,In_373);
nor U215 (N_215,In_262,In_381);
or U216 (N_216,In_126,In_74);
and U217 (N_217,In_282,In_160);
nor U218 (N_218,In_354,In_77);
and U219 (N_219,In_248,In_27);
nand U220 (N_220,In_246,In_426);
or U221 (N_221,In_424,In_134);
nor U222 (N_222,In_170,In_467);
nor U223 (N_223,In_231,In_255);
or U224 (N_224,In_309,In_455);
and U225 (N_225,In_380,In_247);
xnor U226 (N_226,In_88,In_494);
and U227 (N_227,In_144,In_436);
nor U228 (N_228,In_210,In_226);
and U229 (N_229,In_310,In_19);
nand U230 (N_230,In_49,In_96);
nor U231 (N_231,In_305,In_0);
and U232 (N_232,In_274,In_301);
nand U233 (N_233,In_33,In_347);
nor U234 (N_234,In_85,In_207);
nor U235 (N_235,In_8,In_413);
nand U236 (N_236,In_379,In_169);
or U237 (N_237,In_491,In_133);
or U238 (N_238,In_445,In_58);
and U239 (N_239,In_487,In_252);
and U240 (N_240,In_26,In_141);
or U241 (N_241,In_249,In_29);
nor U242 (N_242,In_275,In_334);
and U243 (N_243,In_311,In_312);
and U244 (N_244,In_232,In_328);
and U245 (N_245,In_254,In_47);
or U246 (N_246,In_260,In_61);
nor U247 (N_247,In_345,In_439);
nor U248 (N_248,In_264,In_374);
or U249 (N_249,In_393,In_142);
and U250 (N_250,In_452,In_259);
nand U251 (N_251,In_248,In_16);
nor U252 (N_252,In_368,In_151);
and U253 (N_253,In_28,In_38);
xor U254 (N_254,In_20,In_245);
and U255 (N_255,In_286,In_12);
nand U256 (N_256,In_278,In_122);
and U257 (N_257,In_226,In_291);
nor U258 (N_258,In_198,In_488);
and U259 (N_259,In_151,In_78);
and U260 (N_260,In_241,In_396);
nand U261 (N_261,In_463,In_465);
nor U262 (N_262,In_50,In_433);
nand U263 (N_263,In_51,In_214);
nor U264 (N_264,In_356,In_388);
nand U265 (N_265,In_492,In_311);
and U266 (N_266,In_474,In_405);
nand U267 (N_267,In_299,In_133);
or U268 (N_268,In_358,In_300);
nand U269 (N_269,In_331,In_370);
and U270 (N_270,In_263,In_48);
and U271 (N_271,In_342,In_268);
or U272 (N_272,In_332,In_226);
nor U273 (N_273,In_6,In_131);
nand U274 (N_274,In_490,In_339);
and U275 (N_275,In_271,In_150);
or U276 (N_276,In_362,In_241);
and U277 (N_277,In_27,In_11);
or U278 (N_278,In_155,In_30);
nand U279 (N_279,In_196,In_387);
or U280 (N_280,In_102,In_466);
xor U281 (N_281,In_418,In_182);
or U282 (N_282,In_393,In_52);
nor U283 (N_283,In_213,In_111);
and U284 (N_284,In_375,In_183);
xor U285 (N_285,In_400,In_268);
or U286 (N_286,In_339,In_228);
and U287 (N_287,In_313,In_101);
and U288 (N_288,In_43,In_154);
nand U289 (N_289,In_45,In_129);
nand U290 (N_290,In_365,In_59);
xnor U291 (N_291,In_20,In_251);
and U292 (N_292,In_264,In_68);
nor U293 (N_293,In_224,In_158);
nor U294 (N_294,In_77,In_353);
nand U295 (N_295,In_384,In_294);
or U296 (N_296,In_389,In_126);
nor U297 (N_297,In_398,In_286);
nand U298 (N_298,In_208,In_400);
nand U299 (N_299,In_410,In_92);
nand U300 (N_300,In_492,In_478);
nand U301 (N_301,In_48,In_343);
or U302 (N_302,In_107,In_322);
nand U303 (N_303,In_375,In_18);
or U304 (N_304,In_204,In_9);
or U305 (N_305,In_80,In_138);
and U306 (N_306,In_293,In_244);
nor U307 (N_307,In_154,In_65);
nand U308 (N_308,In_481,In_472);
nor U309 (N_309,In_162,In_447);
nand U310 (N_310,In_24,In_333);
nor U311 (N_311,In_222,In_173);
and U312 (N_312,In_337,In_495);
nor U313 (N_313,In_270,In_349);
nand U314 (N_314,In_373,In_422);
nor U315 (N_315,In_358,In_254);
and U316 (N_316,In_440,In_65);
or U317 (N_317,In_286,In_231);
and U318 (N_318,In_121,In_389);
nand U319 (N_319,In_171,In_435);
nand U320 (N_320,In_343,In_47);
and U321 (N_321,In_490,In_163);
or U322 (N_322,In_47,In_10);
and U323 (N_323,In_372,In_188);
and U324 (N_324,In_36,In_125);
nor U325 (N_325,In_44,In_372);
nor U326 (N_326,In_309,In_261);
or U327 (N_327,In_175,In_454);
and U328 (N_328,In_289,In_89);
nor U329 (N_329,In_229,In_148);
and U330 (N_330,In_152,In_253);
or U331 (N_331,In_281,In_289);
nor U332 (N_332,In_380,In_40);
nand U333 (N_333,In_476,In_352);
and U334 (N_334,In_244,In_93);
nand U335 (N_335,In_23,In_200);
nor U336 (N_336,In_264,In_115);
xor U337 (N_337,In_17,In_111);
and U338 (N_338,In_435,In_409);
or U339 (N_339,In_40,In_115);
nor U340 (N_340,In_94,In_35);
or U341 (N_341,In_102,In_228);
and U342 (N_342,In_370,In_438);
nor U343 (N_343,In_212,In_316);
and U344 (N_344,In_92,In_120);
or U345 (N_345,In_303,In_120);
or U346 (N_346,In_137,In_308);
and U347 (N_347,In_425,In_439);
and U348 (N_348,In_12,In_349);
nor U349 (N_349,In_406,In_334);
or U350 (N_350,In_234,In_404);
nand U351 (N_351,In_458,In_410);
nor U352 (N_352,In_140,In_366);
nand U353 (N_353,In_46,In_67);
and U354 (N_354,In_391,In_415);
nor U355 (N_355,In_297,In_449);
and U356 (N_356,In_471,In_136);
xnor U357 (N_357,In_128,In_215);
nor U358 (N_358,In_241,In_300);
nand U359 (N_359,In_270,In_379);
or U360 (N_360,In_319,In_455);
nand U361 (N_361,In_141,In_486);
and U362 (N_362,In_255,In_203);
nor U363 (N_363,In_439,In_304);
or U364 (N_364,In_114,In_239);
or U365 (N_365,In_127,In_279);
nand U366 (N_366,In_159,In_41);
nand U367 (N_367,In_454,In_339);
nor U368 (N_368,In_42,In_474);
or U369 (N_369,In_273,In_361);
nor U370 (N_370,In_81,In_347);
or U371 (N_371,In_370,In_340);
nor U372 (N_372,In_82,In_493);
nor U373 (N_373,In_268,In_82);
nand U374 (N_374,In_135,In_407);
and U375 (N_375,In_217,In_422);
nand U376 (N_376,In_398,In_154);
nor U377 (N_377,In_373,In_51);
or U378 (N_378,In_467,In_255);
and U379 (N_379,In_333,In_109);
nor U380 (N_380,In_410,In_492);
nand U381 (N_381,In_288,In_40);
nor U382 (N_382,In_482,In_189);
nand U383 (N_383,In_474,In_387);
nor U384 (N_384,In_414,In_163);
or U385 (N_385,In_395,In_305);
or U386 (N_386,In_411,In_419);
or U387 (N_387,In_92,In_442);
nor U388 (N_388,In_5,In_463);
nor U389 (N_389,In_479,In_211);
nor U390 (N_390,In_244,In_192);
and U391 (N_391,In_169,In_389);
or U392 (N_392,In_273,In_216);
nor U393 (N_393,In_375,In_498);
xor U394 (N_394,In_54,In_442);
nand U395 (N_395,In_81,In_351);
nand U396 (N_396,In_125,In_237);
nand U397 (N_397,In_438,In_376);
and U398 (N_398,In_443,In_313);
and U399 (N_399,In_471,In_175);
or U400 (N_400,In_169,In_446);
or U401 (N_401,In_376,In_198);
nor U402 (N_402,In_306,In_72);
and U403 (N_403,In_163,In_408);
nand U404 (N_404,In_403,In_35);
nand U405 (N_405,In_85,In_100);
nor U406 (N_406,In_195,In_295);
and U407 (N_407,In_348,In_63);
nand U408 (N_408,In_135,In_169);
nor U409 (N_409,In_292,In_65);
and U410 (N_410,In_465,In_291);
nand U411 (N_411,In_90,In_436);
and U412 (N_412,In_6,In_151);
and U413 (N_413,In_281,In_398);
nand U414 (N_414,In_332,In_458);
or U415 (N_415,In_87,In_180);
nor U416 (N_416,In_278,In_478);
nand U417 (N_417,In_423,In_161);
xor U418 (N_418,In_137,In_336);
nand U419 (N_419,In_339,In_88);
or U420 (N_420,In_175,In_141);
and U421 (N_421,In_305,In_444);
or U422 (N_422,In_223,In_306);
and U423 (N_423,In_214,In_474);
nor U424 (N_424,In_404,In_401);
nor U425 (N_425,In_271,In_276);
nor U426 (N_426,In_376,In_192);
nand U427 (N_427,In_339,In_470);
and U428 (N_428,In_460,In_318);
or U429 (N_429,In_442,In_345);
and U430 (N_430,In_480,In_421);
or U431 (N_431,In_326,In_191);
nor U432 (N_432,In_59,In_171);
nor U433 (N_433,In_296,In_254);
nor U434 (N_434,In_403,In_18);
and U435 (N_435,In_140,In_356);
or U436 (N_436,In_253,In_207);
nor U437 (N_437,In_136,In_493);
nor U438 (N_438,In_36,In_216);
nand U439 (N_439,In_287,In_443);
or U440 (N_440,In_110,In_361);
or U441 (N_441,In_465,In_494);
nor U442 (N_442,In_358,In_312);
and U443 (N_443,In_239,In_430);
nand U444 (N_444,In_166,In_72);
nand U445 (N_445,In_336,In_124);
xor U446 (N_446,In_158,In_486);
and U447 (N_447,In_39,In_340);
and U448 (N_448,In_343,In_76);
and U449 (N_449,In_426,In_70);
and U450 (N_450,In_4,In_431);
and U451 (N_451,In_94,In_181);
nor U452 (N_452,In_32,In_349);
or U453 (N_453,In_82,In_33);
and U454 (N_454,In_476,In_414);
nor U455 (N_455,In_99,In_483);
or U456 (N_456,In_82,In_334);
nand U457 (N_457,In_128,In_147);
nand U458 (N_458,In_54,In_450);
and U459 (N_459,In_161,In_380);
or U460 (N_460,In_297,In_141);
or U461 (N_461,In_447,In_419);
nand U462 (N_462,In_55,In_113);
and U463 (N_463,In_13,In_203);
nand U464 (N_464,In_488,In_136);
nor U465 (N_465,In_413,In_163);
nor U466 (N_466,In_237,In_300);
or U467 (N_467,In_315,In_185);
xnor U468 (N_468,In_488,In_382);
nor U469 (N_469,In_481,In_483);
nor U470 (N_470,In_188,In_464);
and U471 (N_471,In_23,In_477);
nand U472 (N_472,In_303,In_121);
or U473 (N_473,In_402,In_15);
nor U474 (N_474,In_115,In_200);
or U475 (N_475,In_423,In_299);
xnor U476 (N_476,In_189,In_67);
and U477 (N_477,In_22,In_429);
and U478 (N_478,In_169,In_482);
nand U479 (N_479,In_79,In_464);
nand U480 (N_480,In_133,In_68);
nor U481 (N_481,In_429,In_451);
nand U482 (N_482,In_393,In_19);
and U483 (N_483,In_361,In_41);
xor U484 (N_484,In_235,In_259);
or U485 (N_485,In_26,In_200);
nand U486 (N_486,In_142,In_451);
and U487 (N_487,In_355,In_275);
nand U488 (N_488,In_496,In_2);
nor U489 (N_489,In_457,In_68);
and U490 (N_490,In_209,In_258);
nor U491 (N_491,In_161,In_335);
or U492 (N_492,In_137,In_199);
or U493 (N_493,In_454,In_68);
nand U494 (N_494,In_259,In_401);
or U495 (N_495,In_76,In_225);
or U496 (N_496,In_442,In_384);
nor U497 (N_497,In_268,In_420);
nor U498 (N_498,In_349,In_328);
xor U499 (N_499,In_227,In_276);
and U500 (N_500,In_250,In_378);
nand U501 (N_501,In_257,In_227);
or U502 (N_502,In_14,In_260);
xnor U503 (N_503,In_489,In_251);
nand U504 (N_504,In_172,In_365);
and U505 (N_505,In_389,In_313);
xnor U506 (N_506,In_142,In_192);
nand U507 (N_507,In_139,In_263);
and U508 (N_508,In_16,In_303);
xor U509 (N_509,In_293,In_130);
nor U510 (N_510,In_362,In_351);
nand U511 (N_511,In_152,In_330);
nor U512 (N_512,In_448,In_439);
and U513 (N_513,In_333,In_40);
nor U514 (N_514,In_65,In_107);
and U515 (N_515,In_128,In_390);
and U516 (N_516,In_304,In_187);
nor U517 (N_517,In_435,In_32);
nor U518 (N_518,In_121,In_359);
xor U519 (N_519,In_473,In_13);
xor U520 (N_520,In_333,In_403);
or U521 (N_521,In_185,In_80);
and U522 (N_522,In_403,In_349);
and U523 (N_523,In_319,In_341);
nor U524 (N_524,In_400,In_467);
or U525 (N_525,In_39,In_320);
xnor U526 (N_526,In_169,In_10);
or U527 (N_527,In_282,In_4);
and U528 (N_528,In_328,In_179);
xor U529 (N_529,In_358,In_234);
and U530 (N_530,In_83,In_34);
nor U531 (N_531,In_409,In_426);
or U532 (N_532,In_234,In_499);
nand U533 (N_533,In_464,In_26);
or U534 (N_534,In_429,In_444);
xnor U535 (N_535,In_96,In_209);
nand U536 (N_536,In_487,In_1);
nor U537 (N_537,In_129,In_315);
or U538 (N_538,In_227,In_273);
nand U539 (N_539,In_409,In_344);
nand U540 (N_540,In_74,In_467);
and U541 (N_541,In_387,In_95);
nor U542 (N_542,In_353,In_429);
xnor U543 (N_543,In_27,In_466);
and U544 (N_544,In_215,In_76);
nor U545 (N_545,In_273,In_85);
nor U546 (N_546,In_164,In_192);
nor U547 (N_547,In_24,In_21);
or U548 (N_548,In_257,In_442);
or U549 (N_549,In_297,In_247);
nand U550 (N_550,In_381,In_465);
or U551 (N_551,In_360,In_492);
or U552 (N_552,In_198,In_71);
and U553 (N_553,In_144,In_239);
nand U554 (N_554,In_354,In_331);
nand U555 (N_555,In_428,In_363);
and U556 (N_556,In_34,In_163);
xor U557 (N_557,In_482,In_347);
nor U558 (N_558,In_453,In_403);
nor U559 (N_559,In_370,In_45);
or U560 (N_560,In_483,In_47);
or U561 (N_561,In_149,In_247);
xnor U562 (N_562,In_404,In_116);
or U563 (N_563,In_390,In_329);
or U564 (N_564,In_261,In_139);
and U565 (N_565,In_264,In_388);
nand U566 (N_566,In_64,In_482);
and U567 (N_567,In_106,In_37);
and U568 (N_568,In_54,In_82);
nor U569 (N_569,In_87,In_137);
or U570 (N_570,In_431,In_320);
or U571 (N_571,In_47,In_85);
or U572 (N_572,In_43,In_64);
xor U573 (N_573,In_340,In_433);
nand U574 (N_574,In_8,In_450);
nor U575 (N_575,In_430,In_357);
or U576 (N_576,In_450,In_402);
and U577 (N_577,In_454,In_469);
or U578 (N_578,In_190,In_204);
nand U579 (N_579,In_142,In_316);
or U580 (N_580,In_219,In_418);
and U581 (N_581,In_68,In_195);
nor U582 (N_582,In_472,In_412);
or U583 (N_583,In_78,In_380);
or U584 (N_584,In_159,In_185);
and U585 (N_585,In_466,In_228);
nor U586 (N_586,In_458,In_472);
nor U587 (N_587,In_459,In_410);
nand U588 (N_588,In_279,In_142);
or U589 (N_589,In_435,In_159);
and U590 (N_590,In_149,In_250);
nand U591 (N_591,In_231,In_244);
nand U592 (N_592,In_295,In_448);
or U593 (N_593,In_475,In_435);
nand U594 (N_594,In_52,In_216);
or U595 (N_595,In_87,In_158);
or U596 (N_596,In_155,In_199);
or U597 (N_597,In_70,In_480);
nand U598 (N_598,In_258,In_429);
nand U599 (N_599,In_147,In_305);
nand U600 (N_600,In_470,In_265);
xnor U601 (N_601,In_309,In_77);
and U602 (N_602,In_171,In_459);
or U603 (N_603,In_454,In_111);
or U604 (N_604,In_194,In_442);
and U605 (N_605,In_88,In_131);
nor U606 (N_606,In_402,In_388);
or U607 (N_607,In_366,In_63);
nor U608 (N_608,In_115,In_368);
or U609 (N_609,In_265,In_494);
nand U610 (N_610,In_346,In_62);
xnor U611 (N_611,In_37,In_474);
nand U612 (N_612,In_326,In_455);
or U613 (N_613,In_488,In_395);
nor U614 (N_614,In_164,In_490);
or U615 (N_615,In_134,In_429);
xnor U616 (N_616,In_186,In_106);
or U617 (N_617,In_274,In_179);
or U618 (N_618,In_374,In_494);
xor U619 (N_619,In_242,In_159);
nor U620 (N_620,In_403,In_12);
or U621 (N_621,In_204,In_129);
nand U622 (N_622,In_281,In_147);
nor U623 (N_623,In_457,In_387);
nor U624 (N_624,In_341,In_89);
and U625 (N_625,In_478,In_340);
and U626 (N_626,In_446,In_150);
nor U627 (N_627,In_392,In_454);
or U628 (N_628,In_435,In_252);
nand U629 (N_629,In_296,In_102);
or U630 (N_630,In_148,In_372);
nor U631 (N_631,In_276,In_272);
or U632 (N_632,In_477,In_397);
nand U633 (N_633,In_0,In_270);
and U634 (N_634,In_313,In_260);
and U635 (N_635,In_174,In_385);
and U636 (N_636,In_499,In_281);
and U637 (N_637,In_380,In_306);
nor U638 (N_638,In_345,In_71);
or U639 (N_639,In_336,In_202);
nand U640 (N_640,In_72,In_260);
and U641 (N_641,In_461,In_352);
or U642 (N_642,In_278,In_354);
xor U643 (N_643,In_2,In_179);
and U644 (N_644,In_446,In_87);
or U645 (N_645,In_204,In_471);
and U646 (N_646,In_276,In_449);
and U647 (N_647,In_487,In_459);
xor U648 (N_648,In_127,In_46);
or U649 (N_649,In_497,In_319);
and U650 (N_650,In_438,In_130);
nand U651 (N_651,In_350,In_47);
and U652 (N_652,In_183,In_173);
and U653 (N_653,In_326,In_425);
nor U654 (N_654,In_78,In_391);
or U655 (N_655,In_339,In_44);
and U656 (N_656,In_221,In_163);
or U657 (N_657,In_168,In_255);
and U658 (N_658,In_124,In_498);
nand U659 (N_659,In_488,In_11);
nand U660 (N_660,In_421,In_133);
or U661 (N_661,In_492,In_495);
or U662 (N_662,In_5,In_329);
or U663 (N_663,In_217,In_386);
and U664 (N_664,In_31,In_203);
nor U665 (N_665,In_345,In_99);
or U666 (N_666,In_240,In_404);
nor U667 (N_667,In_78,In_267);
and U668 (N_668,In_388,In_387);
nand U669 (N_669,In_15,In_267);
xnor U670 (N_670,In_330,In_472);
nand U671 (N_671,In_476,In_406);
nor U672 (N_672,In_397,In_229);
nand U673 (N_673,In_79,In_238);
nor U674 (N_674,In_271,In_448);
xor U675 (N_675,In_395,In_215);
and U676 (N_676,In_146,In_414);
nor U677 (N_677,In_133,In_387);
and U678 (N_678,In_288,In_82);
nand U679 (N_679,In_239,In_478);
nand U680 (N_680,In_134,In_76);
and U681 (N_681,In_366,In_426);
nor U682 (N_682,In_466,In_127);
or U683 (N_683,In_44,In_28);
or U684 (N_684,In_408,In_320);
and U685 (N_685,In_204,In_431);
nand U686 (N_686,In_488,In_273);
xor U687 (N_687,In_413,In_393);
nor U688 (N_688,In_97,In_352);
or U689 (N_689,In_73,In_15);
nand U690 (N_690,In_66,In_188);
or U691 (N_691,In_474,In_356);
nand U692 (N_692,In_248,In_190);
or U693 (N_693,In_89,In_39);
and U694 (N_694,In_185,In_314);
xnor U695 (N_695,In_211,In_152);
nand U696 (N_696,In_448,In_89);
and U697 (N_697,In_278,In_464);
nor U698 (N_698,In_318,In_59);
nor U699 (N_699,In_475,In_3);
or U700 (N_700,In_12,In_332);
nand U701 (N_701,In_350,In_443);
nor U702 (N_702,In_361,In_410);
or U703 (N_703,In_389,In_331);
or U704 (N_704,In_207,In_380);
xor U705 (N_705,In_342,In_6);
xnor U706 (N_706,In_478,In_402);
nand U707 (N_707,In_331,In_457);
xnor U708 (N_708,In_357,In_144);
nor U709 (N_709,In_25,In_149);
and U710 (N_710,In_231,In_107);
nand U711 (N_711,In_202,In_33);
or U712 (N_712,In_332,In_66);
and U713 (N_713,In_210,In_262);
nand U714 (N_714,In_205,In_314);
and U715 (N_715,In_165,In_322);
nor U716 (N_716,In_36,In_250);
and U717 (N_717,In_341,In_182);
or U718 (N_718,In_302,In_339);
and U719 (N_719,In_114,In_159);
and U720 (N_720,In_313,In_352);
or U721 (N_721,In_298,In_263);
nand U722 (N_722,In_45,In_337);
or U723 (N_723,In_137,In_396);
and U724 (N_724,In_315,In_174);
or U725 (N_725,In_229,In_470);
nand U726 (N_726,In_159,In_141);
nand U727 (N_727,In_358,In_302);
nor U728 (N_728,In_239,In_441);
nand U729 (N_729,In_353,In_213);
and U730 (N_730,In_96,In_103);
or U731 (N_731,In_269,In_29);
nand U732 (N_732,In_403,In_257);
nor U733 (N_733,In_72,In_32);
or U734 (N_734,In_149,In_39);
xor U735 (N_735,In_87,In_251);
and U736 (N_736,In_357,In_131);
nor U737 (N_737,In_213,In_361);
nor U738 (N_738,In_0,In_2);
nand U739 (N_739,In_210,In_296);
nor U740 (N_740,In_495,In_245);
nor U741 (N_741,In_451,In_418);
nand U742 (N_742,In_346,In_16);
nor U743 (N_743,In_224,In_206);
nand U744 (N_744,In_408,In_275);
nand U745 (N_745,In_381,In_233);
and U746 (N_746,In_406,In_48);
and U747 (N_747,In_488,In_200);
and U748 (N_748,In_400,In_438);
and U749 (N_749,In_359,In_394);
or U750 (N_750,N_372,N_345);
and U751 (N_751,N_282,N_559);
nand U752 (N_752,N_160,N_679);
nor U753 (N_753,N_291,N_68);
and U754 (N_754,N_591,N_536);
or U755 (N_755,N_504,N_281);
xor U756 (N_756,N_147,N_94);
and U757 (N_757,N_623,N_292);
or U758 (N_758,N_299,N_601);
nor U759 (N_759,N_143,N_245);
xor U760 (N_760,N_438,N_335);
and U761 (N_761,N_563,N_379);
xnor U762 (N_762,N_736,N_541);
nor U763 (N_763,N_343,N_476);
nand U764 (N_764,N_229,N_191);
xnor U765 (N_765,N_456,N_682);
nor U766 (N_766,N_22,N_201);
or U767 (N_767,N_547,N_450);
nand U768 (N_768,N_499,N_97);
nand U769 (N_769,N_164,N_522);
nand U770 (N_770,N_706,N_669);
and U771 (N_771,N_444,N_703);
xor U772 (N_772,N_324,N_637);
xor U773 (N_773,N_569,N_220);
xnor U774 (N_774,N_197,N_214);
nor U775 (N_775,N_663,N_749);
and U776 (N_776,N_446,N_85);
xnor U777 (N_777,N_743,N_154);
and U778 (N_778,N_384,N_180);
xnor U779 (N_779,N_689,N_416);
nor U780 (N_780,N_422,N_678);
xor U781 (N_781,N_611,N_517);
xor U782 (N_782,N_358,N_149);
or U783 (N_783,N_8,N_91);
nand U784 (N_784,N_640,N_203);
nand U785 (N_785,N_120,N_35);
nand U786 (N_786,N_118,N_621);
or U787 (N_787,N_538,N_55);
xnor U788 (N_788,N_239,N_276);
nor U789 (N_789,N_205,N_532);
or U790 (N_790,N_179,N_674);
nor U791 (N_791,N_685,N_662);
and U792 (N_792,N_186,N_320);
or U793 (N_793,N_238,N_609);
nand U794 (N_794,N_465,N_13);
or U795 (N_795,N_138,N_426);
nor U796 (N_796,N_348,N_71);
or U797 (N_797,N_268,N_526);
and U798 (N_798,N_698,N_417);
nor U799 (N_799,N_382,N_624);
nor U800 (N_800,N_461,N_215);
xnor U801 (N_801,N_463,N_395);
or U802 (N_802,N_441,N_437);
nand U803 (N_803,N_159,N_712);
xor U804 (N_804,N_53,N_349);
or U805 (N_805,N_369,N_37);
nand U806 (N_806,N_58,N_651);
nand U807 (N_807,N_11,N_162);
nand U808 (N_808,N_515,N_259);
nand U809 (N_809,N_21,N_386);
and U810 (N_810,N_315,N_351);
or U811 (N_811,N_397,N_312);
xnor U812 (N_812,N_723,N_553);
and U813 (N_813,N_537,N_305);
and U814 (N_814,N_66,N_231);
nand U815 (N_815,N_347,N_46);
nor U816 (N_816,N_332,N_666);
nor U817 (N_817,N_468,N_146);
nand U818 (N_818,N_552,N_31);
and U819 (N_819,N_254,N_496);
nor U820 (N_820,N_294,N_524);
or U821 (N_821,N_337,N_396);
and U822 (N_822,N_746,N_664);
nand U823 (N_823,N_472,N_142);
nor U824 (N_824,N_236,N_131);
nor U825 (N_825,N_168,N_331);
xor U826 (N_826,N_399,N_424);
nor U827 (N_827,N_153,N_633);
or U828 (N_828,N_87,N_565);
nor U829 (N_829,N_602,N_230);
nor U830 (N_830,N_627,N_622);
nand U831 (N_831,N_346,N_708);
xor U832 (N_832,N_341,N_188);
nor U833 (N_833,N_725,N_728);
nor U834 (N_834,N_408,N_334);
or U835 (N_835,N_412,N_248);
xor U836 (N_836,N_199,N_356);
nand U837 (N_837,N_634,N_503);
and U838 (N_838,N_523,N_567);
nand U839 (N_839,N_19,N_413);
xor U840 (N_840,N_585,N_575);
and U841 (N_841,N_604,N_603);
or U842 (N_842,N_516,N_308);
nand U843 (N_843,N_256,N_491);
nor U844 (N_844,N_167,N_150);
nand U845 (N_845,N_302,N_610);
nand U846 (N_846,N_126,N_288);
nand U847 (N_847,N_218,N_459);
nand U848 (N_848,N_177,N_277);
or U849 (N_849,N_323,N_650);
nand U850 (N_850,N_132,N_139);
and U851 (N_851,N_605,N_580);
and U852 (N_852,N_740,N_724);
and U853 (N_853,N_551,N_30);
and U854 (N_854,N_270,N_727);
and U855 (N_855,N_612,N_630);
or U856 (N_856,N_701,N_592);
and U857 (N_857,N_649,N_200);
nor U858 (N_858,N_262,N_594);
and U859 (N_859,N_434,N_333);
xor U860 (N_860,N_415,N_208);
xnor U861 (N_861,N_129,N_449);
and U862 (N_862,N_726,N_653);
or U863 (N_863,N_187,N_88);
nand U864 (N_864,N_487,N_303);
and U865 (N_865,N_253,N_161);
nor U866 (N_866,N_16,N_629);
or U867 (N_867,N_325,N_738);
or U868 (N_868,N_598,N_638);
nand U869 (N_869,N_405,N_475);
or U870 (N_870,N_695,N_620);
or U871 (N_871,N_363,N_675);
nor U872 (N_872,N_579,N_520);
and U873 (N_873,N_364,N_133);
or U874 (N_874,N_57,N_272);
and U875 (N_875,N_170,N_462);
and U876 (N_876,N_251,N_387);
nor U877 (N_877,N_709,N_125);
nand U878 (N_878,N_490,N_572);
or U879 (N_879,N_466,N_165);
nor U880 (N_880,N_338,N_488);
or U881 (N_881,N_89,N_617);
nor U882 (N_882,N_717,N_586);
nor U883 (N_883,N_103,N_321);
xnor U884 (N_884,N_116,N_373);
and U885 (N_885,N_518,N_558);
nor U886 (N_886,N_696,N_216);
nand U887 (N_887,N_710,N_110);
nand U888 (N_888,N_148,N_583);
xnor U889 (N_889,N_112,N_119);
and U890 (N_890,N_92,N_407);
nor U891 (N_891,N_28,N_95);
xnor U892 (N_892,N_79,N_183);
and U893 (N_893,N_359,N_352);
and U894 (N_894,N_677,N_655);
and U895 (N_895,N_535,N_86);
nand U896 (N_896,N_484,N_430);
and U897 (N_897,N_309,N_137);
and U898 (N_898,N_322,N_70);
nand U899 (N_899,N_425,N_375);
or U900 (N_900,N_293,N_178);
and U901 (N_901,N_543,N_61);
nand U902 (N_902,N_562,N_127);
and U903 (N_903,N_534,N_684);
nand U904 (N_904,N_301,N_265);
and U905 (N_905,N_401,N_494);
or U906 (N_906,N_285,N_106);
and U907 (N_907,N_217,N_385);
or U908 (N_908,N_173,N_414);
or U909 (N_909,N_40,N_722);
nand U910 (N_910,N_298,N_295);
xnor U911 (N_911,N_700,N_402);
nand U912 (N_912,N_371,N_625);
nand U913 (N_913,N_33,N_419);
and U914 (N_914,N_39,N_495);
or U915 (N_915,N_246,N_613);
nor U916 (N_916,N_578,N_681);
or U917 (N_917,N_658,N_470);
nand U918 (N_918,N_307,N_63);
nand U919 (N_919,N_628,N_76);
nor U920 (N_920,N_519,N_531);
nor U921 (N_921,N_367,N_140);
and U922 (N_922,N_721,N_589);
and U923 (N_923,N_631,N_411);
nand U924 (N_924,N_243,N_157);
xor U925 (N_925,N_427,N_501);
or U926 (N_926,N_394,N_6);
nand U927 (N_927,N_680,N_152);
nand U928 (N_928,N_652,N_227);
nand U929 (N_929,N_497,N_554);
nor U930 (N_930,N_458,N_192);
or U931 (N_931,N_4,N_27);
nand U932 (N_932,N_745,N_720);
or U933 (N_933,N_711,N_557);
nor U934 (N_934,N_156,N_212);
and U935 (N_935,N_93,N_193);
and U936 (N_936,N_24,N_317);
nor U937 (N_937,N_287,N_467);
nor U938 (N_938,N_65,N_692);
nand U939 (N_939,N_544,N_690);
or U940 (N_940,N_353,N_659);
xnor U941 (N_941,N_584,N_699);
or U942 (N_942,N_365,N_460);
nor U943 (N_943,N_90,N_269);
and U944 (N_944,N_433,N_280);
xor U945 (N_945,N_566,N_48);
and U946 (N_946,N_533,N_542);
nor U947 (N_947,N_626,N_111);
or U948 (N_948,N_17,N_388);
and U949 (N_949,N_513,N_702);
or U950 (N_950,N_300,N_52);
nor U951 (N_951,N_508,N_432);
nor U952 (N_952,N_81,N_454);
and U953 (N_953,N_582,N_151);
or U954 (N_954,N_284,N_226);
nand U955 (N_955,N_41,N_117);
or U956 (N_956,N_296,N_383);
or U957 (N_957,N_32,N_12);
nor U958 (N_958,N_600,N_716);
and U959 (N_959,N_109,N_392);
and U960 (N_960,N_730,N_361);
or U961 (N_961,N_175,N_464);
or U962 (N_962,N_474,N_3);
nand U963 (N_963,N_639,N_431);
or U964 (N_964,N_206,N_577);
nor U965 (N_965,N_599,N_310);
xnor U966 (N_966,N_510,N_368);
or U967 (N_967,N_420,N_344);
or U968 (N_968,N_527,N_330);
and U969 (N_969,N_75,N_732);
and U970 (N_970,N_47,N_648);
and U971 (N_971,N_505,N_492);
and U972 (N_972,N_707,N_608);
and U973 (N_973,N_289,N_455);
and U974 (N_974,N_69,N_249);
nand U975 (N_975,N_443,N_99);
or U976 (N_976,N_687,N_279);
and U977 (N_977,N_130,N_548);
and U978 (N_978,N_645,N_469);
nor U979 (N_979,N_228,N_739);
or U980 (N_980,N_1,N_744);
and U981 (N_981,N_336,N_123);
nand U982 (N_982,N_485,N_18);
and U983 (N_983,N_378,N_439);
nor U984 (N_984,N_447,N_737);
xnor U985 (N_985,N_20,N_171);
nand U986 (N_986,N_340,N_619);
xor U987 (N_987,N_374,N_264);
or U988 (N_988,N_257,N_158);
nor U989 (N_989,N_670,N_440);
nand U990 (N_990,N_528,N_74);
or U991 (N_991,N_82,N_656);
or U992 (N_992,N_121,N_15);
nor U993 (N_993,N_290,N_241);
nor U994 (N_994,N_237,N_10);
nor U995 (N_995,N_530,N_135);
nor U996 (N_996,N_77,N_23);
nand U997 (N_997,N_478,N_51);
or U998 (N_998,N_261,N_445);
nor U999 (N_999,N_671,N_661);
xor U1000 (N_1000,N_145,N_45);
nand U1001 (N_1001,N_442,N_376);
nor U1002 (N_1002,N_451,N_113);
nand U1003 (N_1003,N_73,N_128);
nand U1004 (N_1004,N_357,N_509);
and U1005 (N_1005,N_715,N_350);
and U1006 (N_1006,N_360,N_83);
nor U1007 (N_1007,N_404,N_25);
nand U1008 (N_1008,N_693,N_204);
and U1009 (N_1009,N_222,N_550);
xnor U1010 (N_1010,N_172,N_252);
and U1011 (N_1011,N_98,N_641);
and U1012 (N_1012,N_174,N_570);
nand U1013 (N_1013,N_316,N_306);
nand U1014 (N_1014,N_44,N_688);
and U1015 (N_1015,N_719,N_748);
or U1016 (N_1016,N_713,N_0);
nand U1017 (N_1017,N_266,N_409);
nand U1018 (N_1018,N_105,N_221);
nor U1019 (N_1019,N_247,N_114);
nor U1020 (N_1020,N_525,N_54);
nor U1021 (N_1021,N_514,N_64);
and U1022 (N_1022,N_209,N_480);
or U1023 (N_1023,N_673,N_355);
or U1024 (N_1024,N_234,N_235);
nor U1025 (N_1025,N_122,N_546);
and U1026 (N_1026,N_481,N_225);
nand U1027 (N_1027,N_632,N_636);
nand U1028 (N_1028,N_311,N_194);
nor U1029 (N_1029,N_473,N_189);
nor U1030 (N_1030,N_741,N_498);
nand U1031 (N_1031,N_418,N_581);
xor U1032 (N_1032,N_274,N_42);
or U1033 (N_1033,N_576,N_381);
or U1034 (N_1034,N_185,N_448);
or U1035 (N_1035,N_568,N_328);
nand U1036 (N_1036,N_176,N_729);
and U1037 (N_1037,N_36,N_667);
nand U1038 (N_1038,N_271,N_452);
and U1039 (N_1039,N_400,N_618);
or U1040 (N_1040,N_587,N_607);
xor U1041 (N_1041,N_735,N_506);
or U1042 (N_1042,N_102,N_233);
xnor U1043 (N_1043,N_483,N_104);
or U1044 (N_1044,N_124,N_72);
nand U1045 (N_1045,N_2,N_223);
or U1046 (N_1046,N_297,N_595);
nand U1047 (N_1047,N_339,N_486);
nor U1048 (N_1048,N_511,N_314);
nor U1049 (N_1049,N_60,N_326);
and U1050 (N_1050,N_29,N_614);
nand U1051 (N_1051,N_67,N_198);
xor U1052 (N_1052,N_275,N_14);
nand U1053 (N_1053,N_232,N_144);
or U1054 (N_1054,N_255,N_676);
or U1055 (N_1055,N_616,N_471);
nand U1056 (N_1056,N_390,N_267);
nor U1057 (N_1057,N_107,N_342);
nand U1058 (N_1058,N_564,N_166);
nand U1059 (N_1059,N_304,N_529);
or U1060 (N_1060,N_590,N_100);
or U1061 (N_1061,N_377,N_313);
nand U1062 (N_1062,N_49,N_654);
nand U1063 (N_1063,N_457,N_588);
or U1064 (N_1064,N_59,N_683);
nand U1065 (N_1065,N_697,N_318);
or U1066 (N_1066,N_26,N_512);
nand U1067 (N_1067,N_115,N_380);
and U1068 (N_1068,N_286,N_555);
xnor U1069 (N_1069,N_660,N_169);
and U1070 (N_1070,N_665,N_9);
nor U1071 (N_1071,N_5,N_398);
or U1072 (N_1072,N_181,N_34);
and U1073 (N_1073,N_571,N_502);
xor U1074 (N_1074,N_410,N_327);
nand U1075 (N_1075,N_244,N_573);
or U1076 (N_1076,N_597,N_435);
nor U1077 (N_1077,N_521,N_545);
and U1078 (N_1078,N_136,N_428);
nand U1079 (N_1079,N_539,N_556);
xor U1080 (N_1080,N_163,N_733);
and U1081 (N_1081,N_38,N_134);
xor U1082 (N_1082,N_731,N_50);
nor U1083 (N_1083,N_207,N_182);
nand U1084 (N_1084,N_250,N_672);
nand U1085 (N_1085,N_354,N_647);
nor U1086 (N_1086,N_489,N_643);
or U1087 (N_1087,N_705,N_714);
and U1088 (N_1088,N_370,N_319);
or U1089 (N_1089,N_196,N_273);
nor U1090 (N_1090,N_393,N_644);
or U1091 (N_1091,N_202,N_747);
nand U1092 (N_1092,N_421,N_615);
and U1093 (N_1093,N_560,N_362);
or U1094 (N_1094,N_694,N_260);
and U1095 (N_1095,N_211,N_283);
and U1096 (N_1096,N_278,N_213);
xor U1097 (N_1097,N_155,N_657);
nand U1098 (N_1098,N_7,N_391);
nand U1099 (N_1099,N_686,N_561);
nor U1100 (N_1100,N_704,N_596);
nor U1101 (N_1101,N_646,N_718);
nor U1102 (N_1102,N_258,N_78);
and U1103 (N_1103,N_479,N_43);
and U1104 (N_1104,N_540,N_195);
and U1105 (N_1105,N_242,N_635);
or U1106 (N_1106,N_190,N_423);
nand U1107 (N_1107,N_574,N_101);
nor U1108 (N_1108,N_366,N_184);
and U1109 (N_1109,N_219,N_406);
nand U1110 (N_1110,N_507,N_96);
or U1111 (N_1111,N_436,N_642);
nor U1112 (N_1112,N_549,N_734);
nand U1113 (N_1113,N_482,N_141);
or U1114 (N_1114,N_389,N_453);
nand U1115 (N_1115,N_477,N_500);
and U1116 (N_1116,N_240,N_606);
nor U1117 (N_1117,N_593,N_742);
nor U1118 (N_1118,N_429,N_493);
and U1119 (N_1119,N_84,N_329);
nor U1120 (N_1120,N_56,N_80);
or U1121 (N_1121,N_691,N_263);
and U1122 (N_1122,N_224,N_62);
and U1123 (N_1123,N_668,N_108);
nor U1124 (N_1124,N_403,N_210);
and U1125 (N_1125,N_193,N_216);
and U1126 (N_1126,N_309,N_131);
nor U1127 (N_1127,N_15,N_629);
and U1128 (N_1128,N_166,N_232);
xor U1129 (N_1129,N_242,N_109);
and U1130 (N_1130,N_329,N_356);
nand U1131 (N_1131,N_579,N_70);
and U1132 (N_1132,N_555,N_637);
xor U1133 (N_1133,N_550,N_425);
and U1134 (N_1134,N_108,N_43);
nor U1135 (N_1135,N_178,N_636);
or U1136 (N_1136,N_146,N_280);
and U1137 (N_1137,N_366,N_247);
nor U1138 (N_1138,N_10,N_724);
and U1139 (N_1139,N_609,N_471);
and U1140 (N_1140,N_282,N_60);
or U1141 (N_1141,N_455,N_290);
and U1142 (N_1142,N_176,N_520);
or U1143 (N_1143,N_350,N_247);
nand U1144 (N_1144,N_358,N_167);
or U1145 (N_1145,N_93,N_735);
nand U1146 (N_1146,N_334,N_311);
nor U1147 (N_1147,N_741,N_364);
nand U1148 (N_1148,N_229,N_238);
nand U1149 (N_1149,N_697,N_28);
nor U1150 (N_1150,N_24,N_196);
nor U1151 (N_1151,N_554,N_331);
or U1152 (N_1152,N_563,N_105);
or U1153 (N_1153,N_303,N_374);
nand U1154 (N_1154,N_110,N_508);
and U1155 (N_1155,N_516,N_658);
xor U1156 (N_1156,N_475,N_735);
or U1157 (N_1157,N_252,N_46);
or U1158 (N_1158,N_550,N_593);
or U1159 (N_1159,N_569,N_104);
or U1160 (N_1160,N_687,N_641);
nor U1161 (N_1161,N_629,N_17);
nand U1162 (N_1162,N_356,N_670);
nor U1163 (N_1163,N_58,N_36);
xor U1164 (N_1164,N_183,N_43);
xor U1165 (N_1165,N_27,N_133);
xor U1166 (N_1166,N_70,N_445);
nor U1167 (N_1167,N_55,N_328);
nor U1168 (N_1168,N_258,N_384);
nand U1169 (N_1169,N_604,N_521);
xor U1170 (N_1170,N_32,N_2);
nor U1171 (N_1171,N_167,N_713);
nor U1172 (N_1172,N_237,N_174);
or U1173 (N_1173,N_227,N_119);
nand U1174 (N_1174,N_466,N_314);
nor U1175 (N_1175,N_217,N_41);
and U1176 (N_1176,N_436,N_118);
nand U1177 (N_1177,N_737,N_130);
and U1178 (N_1178,N_721,N_702);
nor U1179 (N_1179,N_250,N_26);
nor U1180 (N_1180,N_581,N_669);
nand U1181 (N_1181,N_711,N_597);
nand U1182 (N_1182,N_648,N_375);
nand U1183 (N_1183,N_546,N_291);
nand U1184 (N_1184,N_728,N_454);
and U1185 (N_1185,N_61,N_588);
and U1186 (N_1186,N_39,N_378);
nand U1187 (N_1187,N_714,N_492);
nand U1188 (N_1188,N_728,N_216);
or U1189 (N_1189,N_442,N_706);
nor U1190 (N_1190,N_521,N_231);
and U1191 (N_1191,N_159,N_693);
nor U1192 (N_1192,N_600,N_370);
or U1193 (N_1193,N_563,N_367);
nor U1194 (N_1194,N_748,N_492);
or U1195 (N_1195,N_493,N_156);
xnor U1196 (N_1196,N_551,N_0);
or U1197 (N_1197,N_574,N_98);
and U1198 (N_1198,N_481,N_336);
nor U1199 (N_1199,N_535,N_49);
and U1200 (N_1200,N_243,N_486);
or U1201 (N_1201,N_670,N_215);
or U1202 (N_1202,N_277,N_50);
nand U1203 (N_1203,N_745,N_349);
or U1204 (N_1204,N_509,N_668);
and U1205 (N_1205,N_705,N_593);
nand U1206 (N_1206,N_582,N_572);
and U1207 (N_1207,N_424,N_82);
nor U1208 (N_1208,N_559,N_488);
and U1209 (N_1209,N_160,N_617);
or U1210 (N_1210,N_499,N_130);
nand U1211 (N_1211,N_312,N_76);
and U1212 (N_1212,N_535,N_212);
nand U1213 (N_1213,N_494,N_261);
and U1214 (N_1214,N_238,N_648);
or U1215 (N_1215,N_349,N_2);
nand U1216 (N_1216,N_745,N_126);
nor U1217 (N_1217,N_678,N_582);
and U1218 (N_1218,N_132,N_681);
and U1219 (N_1219,N_535,N_33);
or U1220 (N_1220,N_721,N_348);
or U1221 (N_1221,N_743,N_118);
and U1222 (N_1222,N_683,N_108);
xnor U1223 (N_1223,N_645,N_532);
xnor U1224 (N_1224,N_58,N_153);
nand U1225 (N_1225,N_376,N_368);
xor U1226 (N_1226,N_46,N_101);
and U1227 (N_1227,N_638,N_571);
xor U1228 (N_1228,N_346,N_729);
xor U1229 (N_1229,N_502,N_261);
or U1230 (N_1230,N_512,N_668);
xnor U1231 (N_1231,N_450,N_164);
and U1232 (N_1232,N_418,N_709);
nand U1233 (N_1233,N_554,N_404);
or U1234 (N_1234,N_401,N_588);
nor U1235 (N_1235,N_479,N_205);
xnor U1236 (N_1236,N_339,N_364);
or U1237 (N_1237,N_513,N_442);
and U1238 (N_1238,N_171,N_361);
nor U1239 (N_1239,N_140,N_321);
and U1240 (N_1240,N_96,N_685);
xor U1241 (N_1241,N_53,N_649);
and U1242 (N_1242,N_703,N_302);
nand U1243 (N_1243,N_591,N_621);
nand U1244 (N_1244,N_25,N_335);
nor U1245 (N_1245,N_98,N_112);
nor U1246 (N_1246,N_340,N_384);
nor U1247 (N_1247,N_60,N_500);
and U1248 (N_1248,N_350,N_228);
and U1249 (N_1249,N_569,N_425);
nor U1250 (N_1250,N_624,N_611);
nand U1251 (N_1251,N_162,N_365);
or U1252 (N_1252,N_305,N_11);
or U1253 (N_1253,N_85,N_408);
and U1254 (N_1254,N_260,N_296);
or U1255 (N_1255,N_389,N_495);
nand U1256 (N_1256,N_165,N_188);
nand U1257 (N_1257,N_629,N_375);
nor U1258 (N_1258,N_715,N_696);
nor U1259 (N_1259,N_327,N_642);
nor U1260 (N_1260,N_168,N_697);
xor U1261 (N_1261,N_241,N_331);
xnor U1262 (N_1262,N_296,N_322);
and U1263 (N_1263,N_357,N_354);
xor U1264 (N_1264,N_710,N_74);
nor U1265 (N_1265,N_736,N_141);
and U1266 (N_1266,N_301,N_550);
or U1267 (N_1267,N_533,N_213);
nor U1268 (N_1268,N_583,N_47);
xnor U1269 (N_1269,N_724,N_163);
nor U1270 (N_1270,N_357,N_417);
or U1271 (N_1271,N_390,N_326);
and U1272 (N_1272,N_485,N_227);
or U1273 (N_1273,N_318,N_547);
nor U1274 (N_1274,N_7,N_387);
and U1275 (N_1275,N_697,N_372);
nand U1276 (N_1276,N_373,N_700);
nand U1277 (N_1277,N_476,N_369);
nor U1278 (N_1278,N_129,N_380);
nor U1279 (N_1279,N_296,N_215);
nor U1280 (N_1280,N_710,N_215);
or U1281 (N_1281,N_209,N_706);
nor U1282 (N_1282,N_282,N_592);
and U1283 (N_1283,N_639,N_728);
nand U1284 (N_1284,N_685,N_629);
and U1285 (N_1285,N_615,N_157);
or U1286 (N_1286,N_453,N_87);
and U1287 (N_1287,N_111,N_579);
or U1288 (N_1288,N_544,N_267);
or U1289 (N_1289,N_614,N_81);
or U1290 (N_1290,N_336,N_343);
nand U1291 (N_1291,N_403,N_718);
nand U1292 (N_1292,N_129,N_340);
or U1293 (N_1293,N_400,N_628);
xor U1294 (N_1294,N_212,N_610);
nand U1295 (N_1295,N_56,N_158);
or U1296 (N_1296,N_731,N_524);
and U1297 (N_1297,N_164,N_188);
nand U1298 (N_1298,N_77,N_161);
nand U1299 (N_1299,N_256,N_748);
nor U1300 (N_1300,N_524,N_170);
or U1301 (N_1301,N_191,N_388);
and U1302 (N_1302,N_599,N_366);
or U1303 (N_1303,N_144,N_112);
and U1304 (N_1304,N_614,N_171);
and U1305 (N_1305,N_57,N_223);
and U1306 (N_1306,N_331,N_567);
or U1307 (N_1307,N_669,N_464);
nand U1308 (N_1308,N_126,N_427);
or U1309 (N_1309,N_446,N_501);
or U1310 (N_1310,N_1,N_380);
nand U1311 (N_1311,N_681,N_540);
and U1312 (N_1312,N_306,N_664);
or U1313 (N_1313,N_540,N_328);
or U1314 (N_1314,N_438,N_262);
or U1315 (N_1315,N_663,N_72);
nand U1316 (N_1316,N_650,N_699);
and U1317 (N_1317,N_21,N_354);
and U1318 (N_1318,N_348,N_258);
and U1319 (N_1319,N_687,N_177);
and U1320 (N_1320,N_172,N_218);
nor U1321 (N_1321,N_213,N_415);
or U1322 (N_1322,N_79,N_1);
nand U1323 (N_1323,N_499,N_319);
and U1324 (N_1324,N_650,N_127);
or U1325 (N_1325,N_393,N_195);
xnor U1326 (N_1326,N_29,N_429);
nand U1327 (N_1327,N_236,N_667);
nand U1328 (N_1328,N_216,N_326);
nor U1329 (N_1329,N_386,N_116);
xor U1330 (N_1330,N_4,N_201);
or U1331 (N_1331,N_358,N_440);
nor U1332 (N_1332,N_74,N_296);
nand U1333 (N_1333,N_40,N_63);
nand U1334 (N_1334,N_119,N_534);
nand U1335 (N_1335,N_689,N_59);
and U1336 (N_1336,N_501,N_9);
or U1337 (N_1337,N_354,N_535);
nor U1338 (N_1338,N_116,N_94);
or U1339 (N_1339,N_493,N_665);
nor U1340 (N_1340,N_183,N_665);
xor U1341 (N_1341,N_474,N_476);
or U1342 (N_1342,N_286,N_153);
xnor U1343 (N_1343,N_561,N_40);
or U1344 (N_1344,N_146,N_60);
nand U1345 (N_1345,N_542,N_102);
xnor U1346 (N_1346,N_82,N_563);
and U1347 (N_1347,N_260,N_519);
xnor U1348 (N_1348,N_216,N_238);
nand U1349 (N_1349,N_329,N_164);
nand U1350 (N_1350,N_650,N_101);
xnor U1351 (N_1351,N_604,N_172);
nand U1352 (N_1352,N_551,N_227);
and U1353 (N_1353,N_597,N_710);
or U1354 (N_1354,N_237,N_134);
nand U1355 (N_1355,N_368,N_1);
nand U1356 (N_1356,N_438,N_603);
xnor U1357 (N_1357,N_453,N_124);
and U1358 (N_1358,N_670,N_428);
or U1359 (N_1359,N_556,N_495);
or U1360 (N_1360,N_702,N_596);
nand U1361 (N_1361,N_312,N_420);
or U1362 (N_1362,N_723,N_291);
nand U1363 (N_1363,N_25,N_138);
or U1364 (N_1364,N_380,N_544);
nor U1365 (N_1365,N_449,N_292);
nand U1366 (N_1366,N_118,N_378);
nand U1367 (N_1367,N_60,N_144);
nor U1368 (N_1368,N_705,N_451);
or U1369 (N_1369,N_182,N_484);
nor U1370 (N_1370,N_296,N_731);
or U1371 (N_1371,N_132,N_55);
nor U1372 (N_1372,N_213,N_409);
nand U1373 (N_1373,N_227,N_639);
nor U1374 (N_1374,N_465,N_267);
nand U1375 (N_1375,N_248,N_111);
or U1376 (N_1376,N_729,N_630);
xor U1377 (N_1377,N_734,N_53);
and U1378 (N_1378,N_183,N_722);
nor U1379 (N_1379,N_606,N_174);
nand U1380 (N_1380,N_681,N_724);
and U1381 (N_1381,N_712,N_141);
and U1382 (N_1382,N_53,N_748);
nor U1383 (N_1383,N_471,N_682);
and U1384 (N_1384,N_1,N_698);
or U1385 (N_1385,N_359,N_121);
or U1386 (N_1386,N_303,N_653);
and U1387 (N_1387,N_232,N_732);
nand U1388 (N_1388,N_483,N_677);
or U1389 (N_1389,N_690,N_659);
nor U1390 (N_1390,N_16,N_516);
xnor U1391 (N_1391,N_533,N_167);
or U1392 (N_1392,N_384,N_609);
nand U1393 (N_1393,N_394,N_382);
nand U1394 (N_1394,N_85,N_545);
nor U1395 (N_1395,N_142,N_0);
and U1396 (N_1396,N_443,N_199);
and U1397 (N_1397,N_219,N_582);
and U1398 (N_1398,N_114,N_514);
or U1399 (N_1399,N_414,N_418);
or U1400 (N_1400,N_537,N_748);
and U1401 (N_1401,N_532,N_142);
or U1402 (N_1402,N_519,N_597);
and U1403 (N_1403,N_462,N_409);
nor U1404 (N_1404,N_597,N_286);
or U1405 (N_1405,N_664,N_451);
nand U1406 (N_1406,N_85,N_470);
or U1407 (N_1407,N_676,N_524);
or U1408 (N_1408,N_181,N_386);
and U1409 (N_1409,N_540,N_415);
and U1410 (N_1410,N_148,N_455);
nor U1411 (N_1411,N_241,N_127);
xor U1412 (N_1412,N_636,N_461);
xnor U1413 (N_1413,N_525,N_468);
or U1414 (N_1414,N_372,N_584);
nor U1415 (N_1415,N_562,N_688);
nor U1416 (N_1416,N_181,N_308);
nor U1417 (N_1417,N_160,N_158);
or U1418 (N_1418,N_423,N_309);
and U1419 (N_1419,N_563,N_201);
nand U1420 (N_1420,N_532,N_162);
and U1421 (N_1421,N_298,N_740);
nand U1422 (N_1422,N_417,N_38);
nor U1423 (N_1423,N_160,N_406);
nor U1424 (N_1424,N_624,N_263);
and U1425 (N_1425,N_0,N_402);
nand U1426 (N_1426,N_601,N_392);
or U1427 (N_1427,N_203,N_749);
nand U1428 (N_1428,N_9,N_354);
nor U1429 (N_1429,N_162,N_553);
nand U1430 (N_1430,N_162,N_74);
and U1431 (N_1431,N_44,N_504);
xor U1432 (N_1432,N_739,N_746);
nand U1433 (N_1433,N_226,N_346);
or U1434 (N_1434,N_164,N_562);
or U1435 (N_1435,N_85,N_307);
and U1436 (N_1436,N_673,N_557);
nor U1437 (N_1437,N_387,N_477);
nor U1438 (N_1438,N_355,N_230);
and U1439 (N_1439,N_107,N_563);
and U1440 (N_1440,N_368,N_742);
and U1441 (N_1441,N_398,N_315);
nor U1442 (N_1442,N_336,N_565);
nor U1443 (N_1443,N_443,N_77);
and U1444 (N_1444,N_172,N_216);
or U1445 (N_1445,N_386,N_387);
nand U1446 (N_1446,N_652,N_270);
nor U1447 (N_1447,N_463,N_488);
or U1448 (N_1448,N_643,N_398);
and U1449 (N_1449,N_448,N_194);
and U1450 (N_1450,N_635,N_741);
nand U1451 (N_1451,N_466,N_664);
nor U1452 (N_1452,N_601,N_737);
nand U1453 (N_1453,N_708,N_402);
nor U1454 (N_1454,N_653,N_602);
nor U1455 (N_1455,N_325,N_374);
nor U1456 (N_1456,N_125,N_213);
or U1457 (N_1457,N_184,N_109);
or U1458 (N_1458,N_521,N_643);
and U1459 (N_1459,N_90,N_518);
and U1460 (N_1460,N_348,N_645);
and U1461 (N_1461,N_628,N_101);
or U1462 (N_1462,N_392,N_396);
nor U1463 (N_1463,N_411,N_562);
nand U1464 (N_1464,N_441,N_44);
nor U1465 (N_1465,N_395,N_423);
and U1466 (N_1466,N_638,N_652);
or U1467 (N_1467,N_214,N_486);
or U1468 (N_1468,N_485,N_347);
xnor U1469 (N_1469,N_668,N_476);
nand U1470 (N_1470,N_727,N_484);
and U1471 (N_1471,N_661,N_378);
xor U1472 (N_1472,N_633,N_575);
and U1473 (N_1473,N_183,N_361);
and U1474 (N_1474,N_225,N_153);
xor U1475 (N_1475,N_726,N_393);
or U1476 (N_1476,N_740,N_468);
and U1477 (N_1477,N_358,N_549);
or U1478 (N_1478,N_563,N_561);
nor U1479 (N_1479,N_109,N_231);
nor U1480 (N_1480,N_501,N_555);
and U1481 (N_1481,N_484,N_130);
and U1482 (N_1482,N_516,N_407);
and U1483 (N_1483,N_356,N_365);
and U1484 (N_1484,N_739,N_640);
nand U1485 (N_1485,N_135,N_520);
nand U1486 (N_1486,N_642,N_342);
nor U1487 (N_1487,N_151,N_589);
or U1488 (N_1488,N_77,N_10);
nand U1489 (N_1489,N_337,N_714);
nor U1490 (N_1490,N_570,N_697);
or U1491 (N_1491,N_76,N_43);
nor U1492 (N_1492,N_599,N_305);
xnor U1493 (N_1493,N_185,N_179);
and U1494 (N_1494,N_667,N_233);
nand U1495 (N_1495,N_39,N_629);
and U1496 (N_1496,N_740,N_693);
xnor U1497 (N_1497,N_293,N_749);
and U1498 (N_1498,N_523,N_130);
nor U1499 (N_1499,N_464,N_454);
or U1500 (N_1500,N_1417,N_1263);
and U1501 (N_1501,N_1177,N_766);
or U1502 (N_1502,N_1434,N_1428);
or U1503 (N_1503,N_1068,N_1002);
and U1504 (N_1504,N_941,N_1387);
nand U1505 (N_1505,N_1363,N_1091);
xor U1506 (N_1506,N_925,N_1338);
or U1507 (N_1507,N_966,N_785);
or U1508 (N_1508,N_1406,N_1132);
xor U1509 (N_1509,N_1321,N_1028);
nand U1510 (N_1510,N_1415,N_1009);
and U1511 (N_1511,N_1166,N_900);
nor U1512 (N_1512,N_827,N_770);
nor U1513 (N_1513,N_1025,N_1171);
or U1514 (N_1514,N_1113,N_876);
nand U1515 (N_1515,N_937,N_1441);
nor U1516 (N_1516,N_1401,N_1228);
and U1517 (N_1517,N_798,N_1144);
and U1518 (N_1518,N_1007,N_1054);
and U1519 (N_1519,N_1035,N_982);
and U1520 (N_1520,N_1433,N_793);
and U1521 (N_1521,N_1315,N_1150);
xor U1522 (N_1522,N_1271,N_1360);
nor U1523 (N_1523,N_1126,N_858);
xor U1524 (N_1524,N_1280,N_1129);
nor U1525 (N_1525,N_1257,N_902);
nand U1526 (N_1526,N_915,N_1033);
nand U1527 (N_1527,N_1104,N_1034);
xor U1528 (N_1528,N_799,N_1067);
or U1529 (N_1529,N_1096,N_1460);
nand U1530 (N_1530,N_1203,N_1403);
xor U1531 (N_1531,N_1413,N_1030);
nor U1532 (N_1532,N_1109,N_1165);
nor U1533 (N_1533,N_857,N_1374);
nand U1534 (N_1534,N_1044,N_859);
and U1535 (N_1535,N_1397,N_1452);
and U1536 (N_1536,N_1299,N_1013);
or U1537 (N_1537,N_1318,N_1247);
xor U1538 (N_1538,N_1341,N_1032);
nor U1539 (N_1539,N_1146,N_1252);
or U1540 (N_1540,N_1266,N_1337);
nor U1541 (N_1541,N_974,N_1075);
xnor U1542 (N_1542,N_1355,N_1422);
or U1543 (N_1543,N_947,N_936);
nand U1544 (N_1544,N_842,N_1041);
xor U1545 (N_1545,N_954,N_1380);
nand U1546 (N_1546,N_803,N_1285);
nand U1547 (N_1547,N_1463,N_1158);
or U1548 (N_1548,N_1453,N_1147);
or U1549 (N_1549,N_852,N_767);
or U1550 (N_1550,N_1099,N_867);
nand U1551 (N_1551,N_1004,N_1234);
or U1552 (N_1552,N_1213,N_774);
xor U1553 (N_1553,N_1462,N_1216);
nor U1554 (N_1554,N_924,N_1064);
nand U1555 (N_1555,N_1172,N_828);
or U1556 (N_1556,N_1130,N_1182);
and U1557 (N_1557,N_1449,N_1327);
or U1558 (N_1558,N_875,N_1442);
and U1559 (N_1559,N_1492,N_1268);
or U1560 (N_1560,N_1367,N_926);
nor U1561 (N_1561,N_805,N_1260);
nor U1562 (N_1562,N_841,N_984);
or U1563 (N_1563,N_1308,N_1201);
and U1564 (N_1564,N_1014,N_1479);
nand U1565 (N_1565,N_1480,N_1174);
and U1566 (N_1566,N_895,N_979);
nand U1567 (N_1567,N_1074,N_1061);
or U1568 (N_1568,N_1488,N_939);
xnor U1569 (N_1569,N_1491,N_801);
and U1570 (N_1570,N_1306,N_1135);
or U1571 (N_1571,N_958,N_878);
nor U1572 (N_1572,N_820,N_1421);
or U1573 (N_1573,N_1191,N_929);
nand U1574 (N_1574,N_1153,N_964);
or U1575 (N_1575,N_1371,N_1319);
and U1576 (N_1576,N_919,N_1092);
and U1577 (N_1577,N_991,N_1118);
and U1578 (N_1578,N_946,N_1197);
or U1579 (N_1579,N_1478,N_986);
nand U1580 (N_1580,N_1258,N_1499);
nor U1581 (N_1581,N_957,N_1365);
xor U1582 (N_1582,N_1362,N_1080);
or U1583 (N_1583,N_795,N_1088);
xnor U1584 (N_1584,N_1218,N_1282);
or U1585 (N_1585,N_866,N_1465);
nand U1586 (N_1586,N_775,N_791);
nor U1587 (N_1587,N_920,N_1168);
or U1588 (N_1588,N_1178,N_1382);
and U1589 (N_1589,N_1346,N_1141);
nor U1590 (N_1590,N_967,N_1008);
nand U1591 (N_1591,N_824,N_1354);
nor U1592 (N_1592,N_1196,N_877);
xnor U1593 (N_1593,N_1049,N_1432);
nand U1594 (N_1594,N_1272,N_1329);
or U1595 (N_1595,N_917,N_1388);
nand U1596 (N_1596,N_989,N_1485);
or U1597 (N_1597,N_837,N_787);
xor U1598 (N_1598,N_970,N_1063);
or U1599 (N_1599,N_1461,N_757);
nand U1600 (N_1600,N_848,N_840);
nor U1601 (N_1601,N_1426,N_765);
or U1602 (N_1602,N_1418,N_1475);
nor U1603 (N_1603,N_1438,N_845);
and U1604 (N_1604,N_1286,N_1134);
nor U1605 (N_1605,N_794,N_1469);
nor U1606 (N_1606,N_754,N_1200);
or U1607 (N_1607,N_948,N_999);
nor U1608 (N_1608,N_1467,N_861);
or U1609 (N_1609,N_1006,N_1078);
and U1610 (N_1610,N_1098,N_1240);
nor U1611 (N_1611,N_886,N_913);
or U1612 (N_1612,N_755,N_882);
xor U1613 (N_1613,N_1393,N_871);
nor U1614 (N_1614,N_809,N_1287);
nand U1615 (N_1615,N_1473,N_904);
nor U1616 (N_1616,N_1161,N_911);
nand U1617 (N_1617,N_1160,N_797);
or U1618 (N_1618,N_1190,N_1214);
and U1619 (N_1619,N_1303,N_1112);
nand U1620 (N_1620,N_1253,N_1167);
xor U1621 (N_1621,N_1262,N_872);
xor U1622 (N_1622,N_1137,N_975);
nor U1623 (N_1623,N_1339,N_1019);
xnor U1624 (N_1624,N_1395,N_1310);
nor U1625 (N_1625,N_980,N_1423);
and U1626 (N_1626,N_1486,N_952);
nor U1627 (N_1627,N_776,N_1375);
or U1628 (N_1628,N_1390,N_1373);
nand U1629 (N_1629,N_1281,N_1372);
nand U1630 (N_1630,N_1100,N_1052);
and U1631 (N_1631,N_1073,N_1192);
and U1632 (N_1632,N_1470,N_822);
and U1633 (N_1633,N_849,N_819);
nor U1634 (N_1634,N_1490,N_1187);
nor U1635 (N_1635,N_909,N_1036);
nand U1636 (N_1636,N_1425,N_1094);
xor U1637 (N_1637,N_1246,N_1439);
nand U1638 (N_1638,N_1116,N_914);
and U1639 (N_1639,N_1457,N_1392);
nor U1640 (N_1640,N_853,N_1450);
nor U1641 (N_1641,N_905,N_1121);
nand U1642 (N_1642,N_821,N_1489);
nor U1643 (N_1643,N_1199,N_1267);
xnor U1644 (N_1644,N_833,N_1076);
or U1645 (N_1645,N_1223,N_916);
nor U1646 (N_1646,N_1236,N_945);
or U1647 (N_1647,N_784,N_823);
and U1648 (N_1648,N_1224,N_1335);
xor U1649 (N_1649,N_816,N_1202);
and U1650 (N_1650,N_1176,N_781);
nor U1651 (N_1651,N_1229,N_1378);
and U1652 (N_1652,N_771,N_1250);
or U1653 (N_1653,N_890,N_1291);
nand U1654 (N_1654,N_1226,N_1336);
or U1655 (N_1655,N_1105,N_1069);
nand U1656 (N_1656,N_865,N_1404);
or U1657 (N_1657,N_1027,N_1039);
and U1658 (N_1658,N_1412,N_1241);
or U1659 (N_1659,N_1356,N_1468);
and U1660 (N_1660,N_1328,N_1204);
nor U1661 (N_1661,N_977,N_1139);
and U1662 (N_1662,N_978,N_1464);
or U1663 (N_1663,N_1095,N_1057);
or U1664 (N_1664,N_864,N_1017);
nor U1665 (N_1665,N_1265,N_1189);
nand U1666 (N_1666,N_1237,N_1437);
or U1667 (N_1667,N_800,N_1123);
or U1668 (N_1668,N_854,N_1142);
nand U1669 (N_1669,N_1003,N_1293);
or U1670 (N_1670,N_855,N_1345);
and U1671 (N_1671,N_1084,N_1115);
nor U1672 (N_1672,N_1060,N_1483);
or U1673 (N_1673,N_1083,N_894);
nor U1674 (N_1674,N_1256,N_1093);
nor U1675 (N_1675,N_1410,N_935);
nor U1676 (N_1676,N_1042,N_1451);
nor U1677 (N_1677,N_1435,N_1366);
and U1678 (N_1678,N_1305,N_1159);
nor U1679 (N_1679,N_1323,N_1498);
or U1680 (N_1680,N_1193,N_1255);
nand U1681 (N_1681,N_899,N_1347);
or U1682 (N_1682,N_1184,N_1037);
nand U1683 (N_1683,N_1209,N_1185);
nand U1684 (N_1684,N_1125,N_1409);
nor U1685 (N_1685,N_812,N_1011);
and U1686 (N_1686,N_1179,N_1408);
nand U1687 (N_1687,N_1152,N_750);
or U1688 (N_1688,N_1385,N_1055);
or U1689 (N_1689,N_778,N_1429);
and U1690 (N_1690,N_1359,N_1314);
nor U1691 (N_1691,N_1149,N_1304);
or U1692 (N_1692,N_1108,N_1322);
nand U1693 (N_1693,N_953,N_1277);
and U1694 (N_1694,N_887,N_1454);
nand U1695 (N_1695,N_1377,N_889);
nand U1696 (N_1696,N_1298,N_1261);
nor U1697 (N_1697,N_1148,N_1117);
and U1698 (N_1698,N_918,N_1173);
nor U1699 (N_1699,N_1379,N_1238);
nand U1700 (N_1700,N_1156,N_1021);
or U1701 (N_1701,N_912,N_1264);
or U1702 (N_1702,N_1133,N_987);
nor U1703 (N_1703,N_1046,N_1053);
or U1704 (N_1704,N_1233,N_1106);
xnor U1705 (N_1705,N_1138,N_783);
nand U1706 (N_1706,N_1368,N_1309);
nor U1707 (N_1707,N_1414,N_1169);
nand U1708 (N_1708,N_1496,N_1495);
nand U1709 (N_1709,N_811,N_1022);
nor U1710 (N_1710,N_773,N_1482);
nand U1711 (N_1711,N_1350,N_944);
nand U1712 (N_1712,N_1361,N_1402);
xor U1713 (N_1713,N_761,N_1140);
and U1714 (N_1714,N_1391,N_1056);
nor U1715 (N_1715,N_1000,N_908);
nor U1716 (N_1716,N_808,N_1005);
and U1717 (N_1717,N_831,N_1396);
and U1718 (N_1718,N_1254,N_1151);
or U1719 (N_1719,N_931,N_1381);
or U1720 (N_1720,N_1155,N_1352);
and U1721 (N_1721,N_1211,N_832);
nand U1722 (N_1722,N_1358,N_1188);
and U1723 (N_1723,N_1194,N_1444);
nor U1724 (N_1724,N_1407,N_1364);
nand U1725 (N_1725,N_1227,N_1273);
and U1726 (N_1726,N_1085,N_1270);
or U1727 (N_1727,N_1440,N_1170);
or U1728 (N_1728,N_792,N_896);
nand U1729 (N_1729,N_1207,N_1436);
and U1730 (N_1730,N_921,N_813);
or U1731 (N_1731,N_796,N_884);
nand U1732 (N_1732,N_1048,N_928);
nand U1733 (N_1733,N_1087,N_1332);
or U1734 (N_1734,N_1487,N_863);
nand U1735 (N_1735,N_1029,N_780);
nand U1736 (N_1736,N_1420,N_1269);
nand U1737 (N_1737,N_1333,N_880);
or U1738 (N_1738,N_934,N_1210);
nor U1739 (N_1739,N_1110,N_1430);
nand U1740 (N_1740,N_1231,N_764);
nand U1741 (N_1741,N_1276,N_992);
or U1742 (N_1742,N_873,N_1043);
nand U1743 (N_1743,N_752,N_1220);
or U1744 (N_1744,N_817,N_1343);
nand U1745 (N_1745,N_963,N_1376);
nand U1746 (N_1746,N_951,N_1275);
or U1747 (N_1747,N_1472,N_769);
and U1748 (N_1748,N_930,N_1079);
and U1749 (N_1749,N_1120,N_1058);
nand U1750 (N_1750,N_1143,N_1212);
nor U1751 (N_1751,N_1071,N_1302);
and U1752 (N_1752,N_1424,N_1419);
nand U1753 (N_1753,N_1111,N_1278);
or U1754 (N_1754,N_1244,N_1045);
and U1755 (N_1755,N_1090,N_1259);
nor U1756 (N_1756,N_844,N_856);
xnor U1757 (N_1757,N_753,N_1128);
nand U1758 (N_1758,N_806,N_779);
and U1759 (N_1759,N_1225,N_976);
and U1760 (N_1760,N_968,N_1398);
nand U1761 (N_1761,N_1394,N_906);
nand U1762 (N_1762,N_1274,N_1162);
nand U1763 (N_1763,N_758,N_961);
xor U1764 (N_1764,N_910,N_763);
or U1765 (N_1765,N_846,N_893);
nor U1766 (N_1766,N_1018,N_1294);
and U1767 (N_1767,N_1221,N_1232);
nand U1768 (N_1768,N_1186,N_1222);
nand U1769 (N_1769,N_1493,N_997);
and U1770 (N_1770,N_1427,N_1015);
and U1771 (N_1771,N_836,N_843);
nand U1772 (N_1772,N_815,N_985);
nor U1773 (N_1773,N_1324,N_891);
nand U1774 (N_1774,N_1353,N_789);
nand U1775 (N_1775,N_790,N_1136);
and U1776 (N_1776,N_777,N_1001);
xnor U1777 (N_1777,N_1330,N_826);
nor U1778 (N_1778,N_1459,N_1348);
or U1779 (N_1779,N_1290,N_1038);
or U1780 (N_1780,N_1307,N_1320);
xor U1781 (N_1781,N_1215,N_938);
xor U1782 (N_1782,N_1101,N_1131);
xor U1783 (N_1783,N_751,N_972);
nor U1784 (N_1784,N_1066,N_956);
or U1785 (N_1785,N_907,N_942);
or U1786 (N_1786,N_1047,N_1217);
or U1787 (N_1787,N_1349,N_932);
nand U1788 (N_1788,N_1062,N_1476);
nand U1789 (N_1789,N_1040,N_903);
nor U1790 (N_1790,N_1114,N_1284);
or U1791 (N_1791,N_1230,N_1208);
and U1792 (N_1792,N_1249,N_1154);
nand U1793 (N_1793,N_847,N_1431);
nand U1794 (N_1794,N_1411,N_1344);
or U1795 (N_1795,N_1494,N_1219);
nand U1796 (N_1796,N_1288,N_1458);
nor U1797 (N_1797,N_1103,N_1124);
nand U1798 (N_1798,N_1386,N_788);
nor U1799 (N_1799,N_1289,N_1446);
or U1800 (N_1800,N_969,N_1455);
and U1801 (N_1801,N_762,N_1195);
or U1802 (N_1802,N_1181,N_1072);
nand U1803 (N_1803,N_804,N_1239);
nand U1804 (N_1804,N_888,N_756);
xnor U1805 (N_1805,N_885,N_830);
or U1806 (N_1806,N_1023,N_1312);
nand U1807 (N_1807,N_981,N_818);
nand U1808 (N_1808,N_1340,N_1484);
or U1809 (N_1809,N_810,N_1107);
and U1810 (N_1810,N_1456,N_950);
xnor U1811 (N_1811,N_1466,N_1383);
nand U1812 (N_1812,N_850,N_1016);
or U1813 (N_1813,N_1326,N_1164);
nor U1814 (N_1814,N_851,N_1331);
and U1815 (N_1815,N_760,N_1157);
nand U1816 (N_1816,N_1295,N_1175);
and U1817 (N_1817,N_782,N_1082);
or U1818 (N_1818,N_993,N_1122);
nand U1819 (N_1819,N_802,N_898);
nor U1820 (N_1820,N_996,N_1400);
nand U1821 (N_1821,N_1102,N_1198);
and U1822 (N_1822,N_960,N_1051);
and U1823 (N_1823,N_1012,N_998);
and U1824 (N_1824,N_1292,N_868);
and U1825 (N_1825,N_1031,N_814);
xor U1826 (N_1826,N_1448,N_1279);
and U1827 (N_1827,N_1357,N_1010);
nor U1828 (N_1828,N_881,N_1086);
nand U1829 (N_1829,N_959,N_1065);
nand U1830 (N_1830,N_1180,N_1251);
and U1831 (N_1831,N_834,N_1059);
nor U1832 (N_1832,N_1325,N_1183);
or U1833 (N_1833,N_1389,N_1351);
nor U1834 (N_1834,N_1311,N_1077);
and U1835 (N_1835,N_1334,N_943);
nand U1836 (N_1836,N_923,N_1081);
and U1837 (N_1837,N_1097,N_965);
nor U1838 (N_1838,N_988,N_1481);
or U1839 (N_1839,N_995,N_973);
nor U1840 (N_1840,N_874,N_1050);
or U1841 (N_1841,N_839,N_825);
and U1842 (N_1842,N_1205,N_990);
nand U1843 (N_1843,N_1248,N_1317);
nand U1844 (N_1844,N_772,N_1163);
nor U1845 (N_1845,N_1342,N_1283);
nand U1846 (N_1846,N_1127,N_1384);
nor U1847 (N_1847,N_1296,N_1026);
nand U1848 (N_1848,N_1316,N_1497);
nand U1849 (N_1849,N_870,N_1206);
xor U1850 (N_1850,N_1145,N_1370);
nand U1851 (N_1851,N_883,N_1447);
and U1852 (N_1852,N_862,N_1477);
or U1853 (N_1853,N_835,N_1471);
and U1854 (N_1854,N_1399,N_962);
nand U1855 (N_1855,N_1243,N_927);
or U1856 (N_1856,N_1235,N_949);
or U1857 (N_1857,N_1416,N_1445);
nand U1858 (N_1858,N_971,N_879);
nand U1859 (N_1859,N_1119,N_1020);
nand U1860 (N_1860,N_933,N_1369);
nand U1861 (N_1861,N_1297,N_940);
nand U1862 (N_1862,N_1301,N_1313);
nor U1863 (N_1863,N_1474,N_1024);
nor U1864 (N_1864,N_786,N_869);
and U1865 (N_1865,N_838,N_901);
or U1866 (N_1866,N_759,N_829);
and U1867 (N_1867,N_1242,N_897);
nor U1868 (N_1868,N_892,N_1070);
xnor U1869 (N_1869,N_768,N_983);
nor U1870 (N_1870,N_1443,N_994);
nor U1871 (N_1871,N_807,N_1300);
or U1872 (N_1872,N_922,N_1405);
or U1873 (N_1873,N_1089,N_955);
nand U1874 (N_1874,N_860,N_1245);
xnor U1875 (N_1875,N_1185,N_1384);
xor U1876 (N_1876,N_958,N_1336);
or U1877 (N_1877,N_1262,N_1136);
nor U1878 (N_1878,N_1388,N_1436);
nand U1879 (N_1879,N_1343,N_913);
or U1880 (N_1880,N_942,N_1197);
or U1881 (N_1881,N_1454,N_1083);
or U1882 (N_1882,N_943,N_1309);
nor U1883 (N_1883,N_1301,N_1297);
and U1884 (N_1884,N_1460,N_1187);
and U1885 (N_1885,N_1064,N_1422);
nand U1886 (N_1886,N_1277,N_1027);
nand U1887 (N_1887,N_963,N_966);
nor U1888 (N_1888,N_1192,N_1375);
nand U1889 (N_1889,N_1139,N_963);
or U1890 (N_1890,N_765,N_1226);
nor U1891 (N_1891,N_890,N_1484);
or U1892 (N_1892,N_1272,N_1282);
nor U1893 (N_1893,N_874,N_1309);
nor U1894 (N_1894,N_965,N_969);
or U1895 (N_1895,N_896,N_1476);
nand U1896 (N_1896,N_962,N_903);
nand U1897 (N_1897,N_861,N_1212);
and U1898 (N_1898,N_1110,N_999);
nor U1899 (N_1899,N_1386,N_1274);
and U1900 (N_1900,N_1182,N_830);
and U1901 (N_1901,N_1310,N_857);
nor U1902 (N_1902,N_785,N_1065);
nor U1903 (N_1903,N_1113,N_1394);
nand U1904 (N_1904,N_1168,N_1029);
nand U1905 (N_1905,N_908,N_1045);
nand U1906 (N_1906,N_1461,N_1255);
xor U1907 (N_1907,N_1283,N_1349);
and U1908 (N_1908,N_1320,N_843);
or U1909 (N_1909,N_1470,N_1306);
nand U1910 (N_1910,N_889,N_1191);
or U1911 (N_1911,N_1170,N_1430);
nand U1912 (N_1912,N_1177,N_867);
nor U1913 (N_1913,N_937,N_795);
xor U1914 (N_1914,N_1042,N_1192);
nand U1915 (N_1915,N_886,N_1097);
xnor U1916 (N_1916,N_1208,N_1369);
or U1917 (N_1917,N_1002,N_1076);
or U1918 (N_1918,N_884,N_1245);
nand U1919 (N_1919,N_1153,N_873);
or U1920 (N_1920,N_750,N_1444);
nor U1921 (N_1921,N_1107,N_948);
or U1922 (N_1922,N_901,N_1108);
and U1923 (N_1923,N_990,N_1301);
nand U1924 (N_1924,N_1494,N_841);
nand U1925 (N_1925,N_766,N_1482);
and U1926 (N_1926,N_1115,N_810);
xnor U1927 (N_1927,N_1331,N_1050);
or U1928 (N_1928,N_1308,N_791);
and U1929 (N_1929,N_757,N_923);
nor U1930 (N_1930,N_1329,N_974);
or U1931 (N_1931,N_1395,N_1032);
nand U1932 (N_1932,N_867,N_1152);
nand U1933 (N_1933,N_890,N_831);
nor U1934 (N_1934,N_1482,N_1486);
or U1935 (N_1935,N_1158,N_1109);
and U1936 (N_1936,N_1129,N_1063);
nor U1937 (N_1937,N_837,N_1077);
nand U1938 (N_1938,N_1018,N_1397);
nor U1939 (N_1939,N_1455,N_1203);
and U1940 (N_1940,N_966,N_1208);
and U1941 (N_1941,N_1344,N_1379);
nor U1942 (N_1942,N_1042,N_870);
or U1943 (N_1943,N_820,N_894);
xnor U1944 (N_1944,N_1017,N_998);
nand U1945 (N_1945,N_899,N_1339);
nand U1946 (N_1946,N_843,N_827);
nor U1947 (N_1947,N_1399,N_1280);
nor U1948 (N_1948,N_1141,N_1398);
nand U1949 (N_1949,N_1422,N_771);
xnor U1950 (N_1950,N_1450,N_1240);
nand U1951 (N_1951,N_1185,N_1009);
nand U1952 (N_1952,N_1328,N_954);
nand U1953 (N_1953,N_1307,N_1434);
nor U1954 (N_1954,N_1264,N_1325);
xnor U1955 (N_1955,N_1277,N_1050);
xor U1956 (N_1956,N_1271,N_1347);
nor U1957 (N_1957,N_1043,N_968);
or U1958 (N_1958,N_1382,N_1319);
nand U1959 (N_1959,N_900,N_1126);
nor U1960 (N_1960,N_1316,N_1077);
or U1961 (N_1961,N_1032,N_1053);
nor U1962 (N_1962,N_1129,N_1437);
nand U1963 (N_1963,N_1336,N_850);
nor U1964 (N_1964,N_1467,N_986);
and U1965 (N_1965,N_883,N_1244);
and U1966 (N_1966,N_1018,N_1259);
and U1967 (N_1967,N_950,N_767);
and U1968 (N_1968,N_1144,N_1238);
and U1969 (N_1969,N_1195,N_1461);
or U1970 (N_1970,N_1281,N_1104);
xor U1971 (N_1971,N_795,N_1449);
or U1972 (N_1972,N_989,N_793);
xnor U1973 (N_1973,N_1435,N_764);
nand U1974 (N_1974,N_1119,N_1305);
nand U1975 (N_1975,N_760,N_879);
and U1976 (N_1976,N_879,N_1019);
nor U1977 (N_1977,N_755,N_1404);
nand U1978 (N_1978,N_773,N_976);
nor U1979 (N_1979,N_943,N_1296);
or U1980 (N_1980,N_1038,N_1338);
and U1981 (N_1981,N_869,N_1110);
xor U1982 (N_1982,N_1023,N_1137);
or U1983 (N_1983,N_963,N_1282);
xnor U1984 (N_1984,N_908,N_1172);
nor U1985 (N_1985,N_1374,N_975);
or U1986 (N_1986,N_1186,N_1130);
nor U1987 (N_1987,N_1414,N_1489);
nand U1988 (N_1988,N_1178,N_1454);
or U1989 (N_1989,N_1207,N_975);
nand U1990 (N_1990,N_1498,N_1049);
nand U1991 (N_1991,N_1070,N_896);
or U1992 (N_1992,N_888,N_1113);
nor U1993 (N_1993,N_763,N_1011);
nand U1994 (N_1994,N_1429,N_755);
and U1995 (N_1995,N_971,N_951);
and U1996 (N_1996,N_1109,N_1164);
or U1997 (N_1997,N_1413,N_929);
and U1998 (N_1998,N_992,N_997);
or U1999 (N_1999,N_906,N_1269);
nor U2000 (N_2000,N_895,N_954);
nand U2001 (N_2001,N_935,N_1499);
and U2002 (N_2002,N_1039,N_1120);
nor U2003 (N_2003,N_1377,N_1453);
nand U2004 (N_2004,N_1414,N_788);
or U2005 (N_2005,N_880,N_802);
nor U2006 (N_2006,N_989,N_1369);
nand U2007 (N_2007,N_1497,N_987);
and U2008 (N_2008,N_1391,N_1244);
or U2009 (N_2009,N_1450,N_1078);
nor U2010 (N_2010,N_1042,N_945);
nor U2011 (N_2011,N_822,N_1012);
or U2012 (N_2012,N_1364,N_934);
nand U2013 (N_2013,N_1324,N_760);
xor U2014 (N_2014,N_1355,N_927);
and U2015 (N_2015,N_946,N_852);
nand U2016 (N_2016,N_1049,N_1075);
nor U2017 (N_2017,N_1397,N_934);
nor U2018 (N_2018,N_1210,N_986);
or U2019 (N_2019,N_1400,N_1141);
nand U2020 (N_2020,N_845,N_905);
nand U2021 (N_2021,N_1167,N_1375);
and U2022 (N_2022,N_1409,N_1294);
or U2023 (N_2023,N_1222,N_1178);
and U2024 (N_2024,N_985,N_872);
or U2025 (N_2025,N_1356,N_810);
nor U2026 (N_2026,N_1304,N_1083);
nor U2027 (N_2027,N_1181,N_1363);
xnor U2028 (N_2028,N_1066,N_1286);
nor U2029 (N_2029,N_1158,N_1297);
nand U2030 (N_2030,N_1152,N_843);
and U2031 (N_2031,N_1440,N_876);
and U2032 (N_2032,N_861,N_1219);
nand U2033 (N_2033,N_1358,N_777);
nand U2034 (N_2034,N_1488,N_750);
and U2035 (N_2035,N_1231,N_1001);
nand U2036 (N_2036,N_1366,N_1379);
nor U2037 (N_2037,N_1185,N_783);
and U2038 (N_2038,N_934,N_1107);
or U2039 (N_2039,N_954,N_1041);
nor U2040 (N_2040,N_1392,N_905);
and U2041 (N_2041,N_933,N_1069);
nor U2042 (N_2042,N_1335,N_1228);
nand U2043 (N_2043,N_839,N_930);
nor U2044 (N_2044,N_1215,N_1029);
nand U2045 (N_2045,N_1434,N_1464);
nor U2046 (N_2046,N_1199,N_1486);
nand U2047 (N_2047,N_847,N_1033);
nor U2048 (N_2048,N_1299,N_1447);
and U2049 (N_2049,N_891,N_1430);
xnor U2050 (N_2050,N_1292,N_1394);
nor U2051 (N_2051,N_798,N_1254);
and U2052 (N_2052,N_922,N_1275);
and U2053 (N_2053,N_1214,N_1113);
and U2054 (N_2054,N_1183,N_1333);
nand U2055 (N_2055,N_1148,N_1069);
nor U2056 (N_2056,N_1435,N_1414);
and U2057 (N_2057,N_1012,N_1254);
nand U2058 (N_2058,N_1494,N_1184);
nand U2059 (N_2059,N_765,N_1343);
nand U2060 (N_2060,N_1095,N_1206);
nor U2061 (N_2061,N_1095,N_995);
or U2062 (N_2062,N_956,N_1159);
and U2063 (N_2063,N_1411,N_1498);
and U2064 (N_2064,N_1143,N_951);
or U2065 (N_2065,N_1380,N_766);
nand U2066 (N_2066,N_1239,N_1366);
nor U2067 (N_2067,N_1122,N_1223);
and U2068 (N_2068,N_917,N_1077);
or U2069 (N_2069,N_986,N_1154);
and U2070 (N_2070,N_1399,N_769);
nand U2071 (N_2071,N_1281,N_1492);
nand U2072 (N_2072,N_927,N_757);
nand U2073 (N_2073,N_845,N_1391);
and U2074 (N_2074,N_1305,N_1059);
nor U2075 (N_2075,N_1466,N_1385);
nor U2076 (N_2076,N_944,N_1387);
nor U2077 (N_2077,N_1088,N_826);
or U2078 (N_2078,N_996,N_1330);
or U2079 (N_2079,N_1310,N_1248);
nor U2080 (N_2080,N_1459,N_783);
nor U2081 (N_2081,N_1150,N_760);
or U2082 (N_2082,N_1440,N_1171);
nor U2083 (N_2083,N_1233,N_769);
and U2084 (N_2084,N_1370,N_1204);
and U2085 (N_2085,N_1215,N_759);
nand U2086 (N_2086,N_1171,N_1485);
nor U2087 (N_2087,N_1168,N_985);
nand U2088 (N_2088,N_779,N_1228);
xnor U2089 (N_2089,N_1446,N_1194);
or U2090 (N_2090,N_1054,N_1326);
or U2091 (N_2091,N_1234,N_1351);
or U2092 (N_2092,N_1257,N_888);
or U2093 (N_2093,N_1459,N_1132);
xor U2094 (N_2094,N_878,N_1224);
or U2095 (N_2095,N_1154,N_800);
and U2096 (N_2096,N_1327,N_1470);
nand U2097 (N_2097,N_1316,N_859);
and U2098 (N_2098,N_1388,N_1350);
nor U2099 (N_2099,N_821,N_1373);
and U2100 (N_2100,N_896,N_890);
or U2101 (N_2101,N_973,N_904);
nor U2102 (N_2102,N_1431,N_842);
nor U2103 (N_2103,N_961,N_1084);
xnor U2104 (N_2104,N_1052,N_1248);
nand U2105 (N_2105,N_931,N_960);
nand U2106 (N_2106,N_1184,N_934);
nand U2107 (N_2107,N_1469,N_934);
nor U2108 (N_2108,N_878,N_879);
or U2109 (N_2109,N_870,N_1110);
nand U2110 (N_2110,N_1245,N_865);
nor U2111 (N_2111,N_787,N_1103);
or U2112 (N_2112,N_1196,N_935);
or U2113 (N_2113,N_1178,N_1485);
nor U2114 (N_2114,N_809,N_1279);
or U2115 (N_2115,N_1196,N_793);
nand U2116 (N_2116,N_1097,N_1353);
nand U2117 (N_2117,N_1416,N_768);
or U2118 (N_2118,N_861,N_1090);
and U2119 (N_2119,N_874,N_781);
or U2120 (N_2120,N_970,N_1281);
nand U2121 (N_2121,N_961,N_1432);
or U2122 (N_2122,N_1438,N_1061);
nand U2123 (N_2123,N_750,N_1489);
nor U2124 (N_2124,N_1249,N_1402);
and U2125 (N_2125,N_1320,N_781);
nand U2126 (N_2126,N_1004,N_1022);
nor U2127 (N_2127,N_1488,N_1407);
xnor U2128 (N_2128,N_954,N_1255);
and U2129 (N_2129,N_1330,N_1190);
xnor U2130 (N_2130,N_920,N_1368);
nand U2131 (N_2131,N_1068,N_951);
and U2132 (N_2132,N_1145,N_1412);
nor U2133 (N_2133,N_1357,N_831);
xnor U2134 (N_2134,N_1346,N_999);
xnor U2135 (N_2135,N_1456,N_818);
nand U2136 (N_2136,N_1213,N_1154);
nor U2137 (N_2137,N_1241,N_1121);
and U2138 (N_2138,N_880,N_1390);
nor U2139 (N_2139,N_1235,N_1474);
xnor U2140 (N_2140,N_767,N_989);
nor U2141 (N_2141,N_1222,N_986);
nor U2142 (N_2142,N_884,N_1168);
or U2143 (N_2143,N_1196,N_1131);
nand U2144 (N_2144,N_896,N_1422);
and U2145 (N_2145,N_1488,N_996);
xnor U2146 (N_2146,N_1074,N_826);
or U2147 (N_2147,N_1448,N_779);
and U2148 (N_2148,N_996,N_1375);
nand U2149 (N_2149,N_1277,N_1372);
or U2150 (N_2150,N_1481,N_1032);
and U2151 (N_2151,N_1294,N_1014);
and U2152 (N_2152,N_835,N_850);
nand U2153 (N_2153,N_854,N_991);
and U2154 (N_2154,N_993,N_841);
or U2155 (N_2155,N_1201,N_1321);
or U2156 (N_2156,N_1039,N_1333);
and U2157 (N_2157,N_1065,N_1422);
xnor U2158 (N_2158,N_1154,N_755);
nand U2159 (N_2159,N_965,N_1297);
nand U2160 (N_2160,N_1212,N_812);
nand U2161 (N_2161,N_1162,N_970);
nand U2162 (N_2162,N_1382,N_776);
xnor U2163 (N_2163,N_973,N_1219);
or U2164 (N_2164,N_1343,N_941);
xor U2165 (N_2165,N_1190,N_859);
and U2166 (N_2166,N_1094,N_1153);
xnor U2167 (N_2167,N_1452,N_1381);
nor U2168 (N_2168,N_769,N_883);
xnor U2169 (N_2169,N_1317,N_1442);
and U2170 (N_2170,N_792,N_1445);
xor U2171 (N_2171,N_1189,N_909);
xnor U2172 (N_2172,N_780,N_1039);
and U2173 (N_2173,N_1135,N_1064);
or U2174 (N_2174,N_790,N_1238);
nor U2175 (N_2175,N_1263,N_1393);
nand U2176 (N_2176,N_750,N_867);
or U2177 (N_2177,N_813,N_894);
nand U2178 (N_2178,N_1375,N_890);
and U2179 (N_2179,N_1296,N_898);
and U2180 (N_2180,N_865,N_1004);
xnor U2181 (N_2181,N_1163,N_1276);
nor U2182 (N_2182,N_864,N_1369);
nor U2183 (N_2183,N_1317,N_1374);
and U2184 (N_2184,N_1220,N_1396);
nor U2185 (N_2185,N_1094,N_1267);
or U2186 (N_2186,N_885,N_1341);
xnor U2187 (N_2187,N_1183,N_1305);
or U2188 (N_2188,N_971,N_1372);
or U2189 (N_2189,N_893,N_1394);
and U2190 (N_2190,N_1313,N_1334);
nor U2191 (N_2191,N_1333,N_1131);
nor U2192 (N_2192,N_1013,N_1388);
and U2193 (N_2193,N_1290,N_977);
xnor U2194 (N_2194,N_1126,N_1218);
nand U2195 (N_2195,N_878,N_843);
nor U2196 (N_2196,N_1077,N_1480);
nand U2197 (N_2197,N_1105,N_1238);
or U2198 (N_2198,N_1077,N_1121);
and U2199 (N_2199,N_1042,N_886);
nand U2200 (N_2200,N_1093,N_770);
nor U2201 (N_2201,N_1455,N_1208);
and U2202 (N_2202,N_1111,N_1113);
nand U2203 (N_2203,N_899,N_1350);
xnor U2204 (N_2204,N_1315,N_1367);
nand U2205 (N_2205,N_1052,N_887);
or U2206 (N_2206,N_1378,N_1171);
and U2207 (N_2207,N_1327,N_1411);
and U2208 (N_2208,N_1354,N_1045);
nand U2209 (N_2209,N_828,N_1449);
or U2210 (N_2210,N_1174,N_1310);
nand U2211 (N_2211,N_829,N_1439);
or U2212 (N_2212,N_767,N_1282);
nand U2213 (N_2213,N_1455,N_870);
nand U2214 (N_2214,N_1182,N_775);
nor U2215 (N_2215,N_775,N_895);
nor U2216 (N_2216,N_1162,N_1251);
nor U2217 (N_2217,N_1176,N_1204);
and U2218 (N_2218,N_938,N_1393);
nor U2219 (N_2219,N_1354,N_1460);
nand U2220 (N_2220,N_964,N_1458);
nand U2221 (N_2221,N_1135,N_1152);
and U2222 (N_2222,N_1367,N_834);
nor U2223 (N_2223,N_1218,N_1136);
nor U2224 (N_2224,N_1175,N_1105);
xnor U2225 (N_2225,N_1271,N_790);
nor U2226 (N_2226,N_906,N_808);
and U2227 (N_2227,N_1407,N_768);
or U2228 (N_2228,N_1461,N_916);
and U2229 (N_2229,N_872,N_1498);
nor U2230 (N_2230,N_1352,N_806);
nor U2231 (N_2231,N_1137,N_1193);
or U2232 (N_2232,N_1292,N_1090);
and U2233 (N_2233,N_789,N_1280);
nand U2234 (N_2234,N_890,N_1419);
nand U2235 (N_2235,N_1316,N_771);
nand U2236 (N_2236,N_1135,N_807);
or U2237 (N_2237,N_1417,N_1323);
xnor U2238 (N_2238,N_1418,N_817);
nor U2239 (N_2239,N_1182,N_957);
or U2240 (N_2240,N_1420,N_1186);
and U2241 (N_2241,N_1303,N_918);
and U2242 (N_2242,N_1495,N_1064);
xor U2243 (N_2243,N_1218,N_827);
nand U2244 (N_2244,N_922,N_1326);
or U2245 (N_2245,N_932,N_927);
nand U2246 (N_2246,N_1479,N_979);
nor U2247 (N_2247,N_1252,N_1365);
xnor U2248 (N_2248,N_1163,N_1395);
and U2249 (N_2249,N_963,N_999);
and U2250 (N_2250,N_2183,N_1812);
or U2251 (N_2251,N_2096,N_2139);
nor U2252 (N_2252,N_1710,N_1790);
and U2253 (N_2253,N_1838,N_2202);
and U2254 (N_2254,N_1846,N_1713);
nor U2255 (N_2255,N_1945,N_2094);
nand U2256 (N_2256,N_1515,N_1941);
and U2257 (N_2257,N_1773,N_1841);
and U2258 (N_2258,N_1850,N_1525);
and U2259 (N_2259,N_1662,N_2204);
nor U2260 (N_2260,N_2165,N_1611);
or U2261 (N_2261,N_1882,N_2176);
nor U2262 (N_2262,N_2113,N_2198);
or U2263 (N_2263,N_2076,N_1533);
nor U2264 (N_2264,N_2177,N_1683);
and U2265 (N_2265,N_2024,N_1982);
and U2266 (N_2266,N_1736,N_1535);
nor U2267 (N_2267,N_2144,N_2081);
or U2268 (N_2268,N_1897,N_1800);
nand U2269 (N_2269,N_1952,N_1877);
or U2270 (N_2270,N_1682,N_1810);
and U2271 (N_2271,N_1906,N_2121);
or U2272 (N_2272,N_1577,N_2194);
or U2273 (N_2273,N_2103,N_1762);
nand U2274 (N_2274,N_1648,N_1777);
and U2275 (N_2275,N_2141,N_2133);
nor U2276 (N_2276,N_2209,N_1604);
or U2277 (N_2277,N_1962,N_2243);
xnor U2278 (N_2278,N_2112,N_1609);
nor U2279 (N_2279,N_1717,N_2119);
nand U2280 (N_2280,N_2179,N_2151);
or U2281 (N_2281,N_1749,N_1509);
nor U2282 (N_2282,N_1538,N_2167);
and U2283 (N_2283,N_1776,N_2124);
and U2284 (N_2284,N_2062,N_1778);
nand U2285 (N_2285,N_1964,N_1892);
or U2286 (N_2286,N_1645,N_2145);
nor U2287 (N_2287,N_1861,N_1744);
and U2288 (N_2288,N_1903,N_2162);
xnor U2289 (N_2289,N_1669,N_2182);
nor U2290 (N_2290,N_1907,N_1524);
and U2291 (N_2291,N_1751,N_1862);
nor U2292 (N_2292,N_2193,N_1786);
nand U2293 (N_2293,N_1613,N_2027);
xor U2294 (N_2294,N_1804,N_1832);
nand U2295 (N_2295,N_2012,N_1792);
nand U2296 (N_2296,N_1559,N_2017);
nor U2297 (N_2297,N_1876,N_2042);
nand U2298 (N_2298,N_1798,N_2231);
and U2299 (N_2299,N_1597,N_1935);
or U2300 (N_2300,N_2000,N_1652);
or U2301 (N_2301,N_2093,N_1901);
nor U2302 (N_2302,N_2152,N_1995);
nor U2303 (N_2303,N_2217,N_1988);
xnor U2304 (N_2304,N_2157,N_1508);
nand U2305 (N_2305,N_1573,N_1771);
nor U2306 (N_2306,N_2004,N_2160);
and U2307 (N_2307,N_2210,N_1830);
or U2308 (N_2308,N_2180,N_1546);
nor U2309 (N_2309,N_1851,N_1829);
nand U2310 (N_2310,N_1701,N_2115);
xnor U2311 (N_2311,N_1925,N_1621);
and U2312 (N_2312,N_2080,N_1722);
and U2313 (N_2313,N_2129,N_2086);
and U2314 (N_2314,N_1822,N_1872);
nand U2315 (N_2315,N_1680,N_1864);
nor U2316 (N_2316,N_1818,N_1808);
nor U2317 (N_2317,N_2154,N_1527);
nand U2318 (N_2318,N_1689,N_1765);
or U2319 (N_2319,N_1551,N_1900);
xnor U2320 (N_2320,N_1581,N_1658);
xnor U2321 (N_2321,N_1780,N_2127);
or U2322 (N_2322,N_2207,N_1998);
nand U2323 (N_2323,N_1735,N_2238);
xnor U2324 (N_2324,N_1705,N_2072);
xor U2325 (N_2325,N_1550,N_2242);
nand U2326 (N_2326,N_2116,N_2146);
nor U2327 (N_2327,N_1819,N_1575);
nand U2328 (N_2328,N_1750,N_1927);
nor U2329 (N_2329,N_1625,N_1895);
nor U2330 (N_2330,N_1547,N_2232);
nand U2331 (N_2331,N_1562,N_2101);
xnor U2332 (N_2332,N_2130,N_1899);
or U2333 (N_2333,N_1920,N_1879);
nand U2334 (N_2334,N_1950,N_1653);
or U2335 (N_2335,N_1685,N_1728);
and U2336 (N_2336,N_1628,N_1972);
xnor U2337 (N_2337,N_1840,N_1878);
or U2338 (N_2338,N_2082,N_1983);
nand U2339 (N_2339,N_1811,N_1794);
or U2340 (N_2340,N_1724,N_1757);
nand U2341 (N_2341,N_2097,N_2098);
nand U2342 (N_2342,N_1937,N_2197);
and U2343 (N_2343,N_1960,N_1943);
xnor U2344 (N_2344,N_1855,N_2018);
nor U2345 (N_2345,N_2228,N_1865);
or U2346 (N_2346,N_1591,N_1867);
nand U2347 (N_2347,N_2033,N_1536);
nand U2348 (N_2348,N_1820,N_1809);
nor U2349 (N_2349,N_1843,N_2218);
or U2350 (N_2350,N_1993,N_1636);
and U2351 (N_2351,N_1886,N_1593);
nand U2352 (N_2352,N_1957,N_1631);
or U2353 (N_2353,N_1542,N_1874);
nand U2354 (N_2354,N_2047,N_1714);
nor U2355 (N_2355,N_1959,N_1672);
nand U2356 (N_2356,N_1918,N_1720);
and U2357 (N_2357,N_2002,N_1707);
and U2358 (N_2358,N_2178,N_1990);
and U2359 (N_2359,N_1534,N_1549);
and U2360 (N_2360,N_1803,N_1640);
or U2361 (N_2361,N_2205,N_1727);
and U2362 (N_2362,N_2057,N_2009);
nand U2363 (N_2363,N_2169,N_1913);
and U2364 (N_2364,N_1940,N_1583);
or U2365 (N_2365,N_1999,N_1603);
nor U2366 (N_2366,N_2142,N_1815);
xnor U2367 (N_2367,N_1712,N_2037);
nand U2368 (N_2368,N_1719,N_1635);
and U2369 (N_2369,N_1791,N_2244);
nand U2370 (N_2370,N_1684,N_1737);
and U2371 (N_2371,N_1526,N_1734);
nor U2372 (N_2372,N_2028,N_2034);
and U2373 (N_2373,N_1799,N_1620);
nand U2374 (N_2374,N_1555,N_2046);
nand U2375 (N_2375,N_2029,N_1976);
or U2376 (N_2376,N_1514,N_1761);
nand U2377 (N_2377,N_1503,N_1989);
or U2378 (N_2378,N_1958,N_1805);
or U2379 (N_2379,N_1698,N_1934);
nor U2380 (N_2380,N_1585,N_1632);
xnor U2381 (N_2381,N_2088,N_2156);
nor U2382 (N_2382,N_1571,N_1731);
or U2383 (N_2383,N_1847,N_1980);
and U2384 (N_2384,N_2114,N_1711);
or U2385 (N_2385,N_1733,N_1606);
and U2386 (N_2386,N_1963,N_1833);
nor U2387 (N_2387,N_2233,N_1917);
nor U2388 (N_2388,N_1730,N_2161);
nor U2389 (N_2389,N_2105,N_1574);
xor U2390 (N_2390,N_1806,N_1755);
nor U2391 (N_2391,N_1661,N_2234);
and U2392 (N_2392,N_1823,N_1979);
nand U2393 (N_2393,N_1890,N_1852);
nor U2394 (N_2394,N_1985,N_2149);
nor U2395 (N_2395,N_1693,N_1646);
nor U2396 (N_2396,N_1802,N_2071);
or U2397 (N_2397,N_1857,N_1789);
or U2398 (N_2398,N_1660,N_1931);
nor U2399 (N_2399,N_2206,N_2230);
nand U2400 (N_2400,N_1715,N_2065);
and U2401 (N_2401,N_2039,N_1814);
or U2402 (N_2402,N_2173,N_1747);
or U2403 (N_2403,N_1914,N_1760);
or U2404 (N_2404,N_1974,N_2188);
nor U2405 (N_2405,N_2064,N_1997);
and U2406 (N_2406,N_2239,N_1987);
nand U2407 (N_2407,N_1991,N_1563);
nor U2408 (N_2408,N_2181,N_1570);
or U2409 (N_2409,N_1994,N_1739);
nand U2410 (N_2410,N_1670,N_1586);
nor U2411 (N_2411,N_1970,N_2148);
or U2412 (N_2412,N_1610,N_1567);
or U2413 (N_2413,N_1947,N_2184);
nand U2414 (N_2414,N_1647,N_1986);
or U2415 (N_2415,N_1908,N_1665);
and U2416 (N_2416,N_1881,N_2211);
or U2417 (N_2417,N_2050,N_1898);
and U2418 (N_2418,N_2052,N_1537);
and U2419 (N_2419,N_2219,N_2010);
or U2420 (N_2420,N_1854,N_2038);
or U2421 (N_2421,N_2158,N_1825);
or U2422 (N_2422,N_1568,N_2109);
and U2423 (N_2423,N_1654,N_1596);
xor U2424 (N_2424,N_2077,N_2137);
and U2425 (N_2425,N_1837,N_1759);
nor U2426 (N_2426,N_2245,N_2008);
nor U2427 (N_2427,N_2168,N_1687);
nand U2428 (N_2428,N_2227,N_1602);
and U2429 (N_2429,N_2091,N_1594);
nor U2430 (N_2430,N_1826,N_2053);
xor U2431 (N_2431,N_2135,N_1894);
nand U2432 (N_2432,N_1929,N_1772);
and U2433 (N_2433,N_1844,N_1502);
nand U2434 (N_2434,N_1651,N_2222);
and U2435 (N_2435,N_1605,N_2019);
nor U2436 (N_2436,N_1520,N_1726);
or U2437 (N_2437,N_2099,N_2164);
nor U2438 (N_2438,N_1746,N_1531);
nor U2439 (N_2439,N_1633,N_2068);
nand U2440 (N_2440,N_1691,N_1748);
and U2441 (N_2441,N_2069,N_1540);
nand U2442 (N_2442,N_1949,N_2166);
nor U2443 (N_2443,N_1572,N_1853);
nor U2444 (N_2444,N_2214,N_1930);
or U2445 (N_2445,N_1909,N_1787);
nand U2446 (N_2446,N_2163,N_1578);
and U2447 (N_2447,N_1919,N_2030);
or U2448 (N_2448,N_1885,N_1557);
nor U2449 (N_2449,N_1599,N_1637);
nand U2450 (N_2450,N_2138,N_1911);
and U2451 (N_2451,N_1518,N_1500);
or U2452 (N_2452,N_1675,N_1768);
and U2453 (N_2453,N_1639,N_1875);
nor U2454 (N_2454,N_1592,N_1860);
xor U2455 (N_2455,N_2044,N_1942);
or U2456 (N_2456,N_1828,N_1560);
nor U2457 (N_2457,N_1643,N_2174);
xnor U2458 (N_2458,N_1912,N_1706);
nand U2459 (N_2459,N_2003,N_2125);
nand U2460 (N_2460,N_2036,N_1741);
and U2461 (N_2461,N_2226,N_2235);
nand U2462 (N_2462,N_2147,N_1624);
nor U2463 (N_2463,N_1782,N_1924);
nand U2464 (N_2464,N_1729,N_1576);
nand U2465 (N_2465,N_1650,N_1992);
nand U2466 (N_2466,N_2200,N_2035);
or U2467 (N_2467,N_1922,N_1558);
nand U2468 (N_2468,N_2060,N_1785);
nand U2469 (N_2469,N_1601,N_2189);
or U2470 (N_2470,N_1686,N_2224);
or U2471 (N_2471,N_1887,N_2134);
or U2472 (N_2472,N_2132,N_1552);
and U2473 (N_2473,N_1888,N_1529);
or U2474 (N_2474,N_1968,N_1905);
or U2475 (N_2475,N_1775,N_1793);
nand U2476 (N_2476,N_2007,N_1936);
nand U2477 (N_2477,N_1981,N_2199);
nor U2478 (N_2478,N_2192,N_1543);
nand U2479 (N_2479,N_2058,N_2171);
and U2480 (N_2480,N_1622,N_1590);
nand U2481 (N_2481,N_1965,N_1921);
nor U2482 (N_2482,N_2067,N_1692);
and U2483 (N_2483,N_1781,N_1655);
or U2484 (N_2484,N_2056,N_2212);
nor U2485 (N_2485,N_1673,N_1566);
nor U2486 (N_2486,N_1516,N_1598);
and U2487 (N_2487,N_1893,N_1511);
and U2488 (N_2488,N_1745,N_2020);
nand U2489 (N_2489,N_1946,N_1764);
nand U2490 (N_2490,N_1767,N_1580);
nand U2491 (N_2491,N_1700,N_2063);
or U2492 (N_2492,N_1545,N_1953);
xor U2493 (N_2493,N_1589,N_2128);
and U2494 (N_2494,N_1753,N_2203);
and U2495 (N_2495,N_1505,N_1817);
nand U2496 (N_2496,N_2061,N_1716);
nand U2497 (N_2497,N_2078,N_1626);
and U2498 (N_2498,N_2104,N_1770);
or U2499 (N_2499,N_2040,N_1629);
nand U2500 (N_2500,N_2237,N_2048);
and U2501 (N_2501,N_1896,N_1696);
and U2502 (N_2502,N_1721,N_1649);
or U2503 (N_2503,N_1816,N_1584);
or U2504 (N_2504,N_2123,N_1630);
nor U2505 (N_2505,N_1679,N_1834);
nand U2506 (N_2506,N_1856,N_2175);
or U2507 (N_2507,N_1513,N_2074);
nor U2508 (N_2508,N_2085,N_1544);
nand U2509 (N_2509,N_1708,N_1723);
nor U2510 (N_2510,N_1532,N_2015);
nand U2511 (N_2511,N_2221,N_1969);
nand U2512 (N_2512,N_2051,N_1866);
or U2513 (N_2513,N_1948,N_1541);
or U2514 (N_2514,N_1699,N_2170);
nand U2515 (N_2515,N_2013,N_1756);
and U2516 (N_2516,N_1961,N_2005);
or U2517 (N_2517,N_2021,N_1659);
or U2518 (N_2518,N_1663,N_1868);
xnor U2519 (N_2519,N_2026,N_2001);
nor U2520 (N_2520,N_1530,N_1564);
and U2521 (N_2521,N_1612,N_2014);
or U2522 (N_2522,N_1774,N_2117);
nor U2523 (N_2523,N_1678,N_2022);
and U2524 (N_2524,N_1709,N_1587);
nor U2525 (N_2525,N_1902,N_1556);
or U2526 (N_2526,N_1758,N_1666);
nand U2527 (N_2527,N_1928,N_1795);
nand U2528 (N_2528,N_1501,N_1973);
and U2529 (N_2529,N_1638,N_2100);
or U2530 (N_2530,N_2223,N_1763);
and U2531 (N_2531,N_1506,N_2190);
nand U2532 (N_2532,N_1971,N_1623);
and U2533 (N_2533,N_1944,N_1939);
nand U2534 (N_2534,N_1694,N_1967);
or U2535 (N_2535,N_2201,N_1932);
and U2536 (N_2536,N_2089,N_1891);
nor U2537 (N_2537,N_1579,N_2059);
nand U2538 (N_2538,N_1954,N_2102);
nor U2539 (N_2539,N_1788,N_1703);
nand U2540 (N_2540,N_2011,N_1996);
and U2541 (N_2541,N_1779,N_2220);
nor U2542 (N_2542,N_1674,N_1858);
and U2543 (N_2543,N_2084,N_2111);
or U2544 (N_2544,N_1845,N_1743);
nor U2545 (N_2545,N_2087,N_1923);
nand U2546 (N_2546,N_2066,N_1807);
or U2547 (N_2547,N_2216,N_1539);
and U2548 (N_2548,N_1582,N_2045);
and U2549 (N_2549,N_1978,N_2196);
nor U2550 (N_2550,N_1884,N_1554);
nand U2551 (N_2551,N_1836,N_1504);
nor U2552 (N_2552,N_2229,N_2195);
nor U2553 (N_2553,N_2246,N_2023);
and U2554 (N_2554,N_1608,N_1522);
nand U2555 (N_2555,N_1619,N_1938);
or U2556 (N_2556,N_1955,N_1695);
nor U2557 (N_2557,N_1681,N_1588);
and U2558 (N_2558,N_2172,N_2247);
nand U2559 (N_2559,N_2075,N_1889);
or U2560 (N_2560,N_1740,N_1702);
or U2561 (N_2561,N_1671,N_2131);
and U2562 (N_2562,N_1616,N_1676);
nand U2563 (N_2563,N_2070,N_2090);
or U2564 (N_2564,N_1752,N_1668);
and U2565 (N_2565,N_2153,N_2140);
nor U2566 (N_2566,N_2110,N_1519);
nand U2567 (N_2567,N_1827,N_1521);
and U2568 (N_2568,N_2191,N_1839);
and U2569 (N_2569,N_1641,N_1951);
and U2570 (N_2570,N_1870,N_1553);
nand U2571 (N_2571,N_1975,N_1849);
or U2572 (N_2572,N_1797,N_1796);
and U2573 (N_2573,N_2236,N_1732);
xnor U2574 (N_2574,N_1742,N_2049);
nor U2575 (N_2575,N_1933,N_1565);
or U2576 (N_2576,N_2159,N_1915);
nand U2577 (N_2577,N_1926,N_2187);
xnor U2578 (N_2578,N_1966,N_1904);
xnor U2579 (N_2579,N_1801,N_1821);
nand U2580 (N_2580,N_1642,N_1615);
and U2581 (N_2581,N_1614,N_2150);
or U2582 (N_2582,N_2092,N_2006);
or U2583 (N_2583,N_1627,N_2136);
nor U2584 (N_2584,N_2213,N_1657);
and U2585 (N_2585,N_1569,N_2185);
nand U2586 (N_2586,N_1600,N_1507);
or U2587 (N_2587,N_1977,N_2031);
and U2588 (N_2588,N_2143,N_2083);
xor U2589 (N_2589,N_1688,N_2126);
nor U2590 (N_2590,N_1718,N_1548);
and U2591 (N_2591,N_2240,N_1848);
or U2592 (N_2592,N_1725,N_2032);
nand U2593 (N_2593,N_1956,N_1607);
xnor U2594 (N_2594,N_2054,N_1677);
nor U2595 (N_2595,N_2155,N_1813);
or U2596 (N_2596,N_2055,N_2241);
and U2597 (N_2597,N_1835,N_1634);
nand U2598 (N_2598,N_1618,N_1824);
nor U2599 (N_2599,N_1754,N_1644);
and U2600 (N_2600,N_1738,N_1704);
and U2601 (N_2601,N_1595,N_1783);
xnor U2602 (N_2602,N_2120,N_1517);
nand U2603 (N_2603,N_2208,N_1656);
nor U2604 (N_2604,N_1869,N_2079);
nand U2605 (N_2605,N_1871,N_2118);
or U2606 (N_2606,N_1831,N_1523);
or U2607 (N_2607,N_2107,N_1690);
xor U2608 (N_2608,N_2122,N_1697);
nand U2609 (N_2609,N_1617,N_1910);
and U2610 (N_2610,N_1510,N_1561);
or U2611 (N_2611,N_2248,N_2041);
and U2612 (N_2612,N_1528,N_2215);
or U2613 (N_2613,N_2108,N_2095);
and U2614 (N_2614,N_1880,N_1766);
nand U2615 (N_2615,N_2186,N_2225);
and U2616 (N_2616,N_1512,N_1842);
nand U2617 (N_2617,N_1873,N_2073);
or U2618 (N_2618,N_1664,N_2249);
nand U2619 (N_2619,N_1863,N_1784);
or U2620 (N_2620,N_1859,N_1883);
or U2621 (N_2621,N_2025,N_1916);
nand U2622 (N_2622,N_1984,N_2106);
or U2623 (N_2623,N_2016,N_1769);
and U2624 (N_2624,N_2043,N_1667);
or U2625 (N_2625,N_2212,N_2134);
nor U2626 (N_2626,N_1633,N_1884);
nor U2627 (N_2627,N_1722,N_1883);
and U2628 (N_2628,N_1744,N_2161);
nand U2629 (N_2629,N_1738,N_1791);
nand U2630 (N_2630,N_1730,N_2173);
nor U2631 (N_2631,N_1695,N_1504);
nand U2632 (N_2632,N_1833,N_2211);
and U2633 (N_2633,N_2022,N_1863);
nor U2634 (N_2634,N_1902,N_1751);
nor U2635 (N_2635,N_1563,N_2245);
or U2636 (N_2636,N_1981,N_2220);
nand U2637 (N_2637,N_1880,N_1715);
or U2638 (N_2638,N_2079,N_1912);
xnor U2639 (N_2639,N_1607,N_1664);
and U2640 (N_2640,N_2019,N_2066);
xnor U2641 (N_2641,N_2033,N_2134);
nand U2642 (N_2642,N_2110,N_2236);
or U2643 (N_2643,N_2230,N_1907);
or U2644 (N_2644,N_2237,N_1697);
or U2645 (N_2645,N_1736,N_1979);
nor U2646 (N_2646,N_2146,N_2088);
and U2647 (N_2647,N_2066,N_1679);
nand U2648 (N_2648,N_2039,N_1922);
nand U2649 (N_2649,N_2012,N_2083);
or U2650 (N_2650,N_1541,N_1902);
nand U2651 (N_2651,N_2212,N_1820);
nor U2652 (N_2652,N_2023,N_1871);
and U2653 (N_2653,N_1715,N_2173);
and U2654 (N_2654,N_2147,N_1692);
and U2655 (N_2655,N_1573,N_1518);
nand U2656 (N_2656,N_1838,N_2128);
nand U2657 (N_2657,N_1759,N_1739);
nor U2658 (N_2658,N_1560,N_1758);
and U2659 (N_2659,N_1501,N_1627);
nand U2660 (N_2660,N_1719,N_1935);
nor U2661 (N_2661,N_2151,N_2145);
and U2662 (N_2662,N_2065,N_1784);
or U2663 (N_2663,N_1580,N_2235);
nor U2664 (N_2664,N_1751,N_1910);
xor U2665 (N_2665,N_1961,N_1836);
and U2666 (N_2666,N_1856,N_1793);
and U2667 (N_2667,N_1819,N_1666);
or U2668 (N_2668,N_2247,N_2214);
xor U2669 (N_2669,N_1651,N_1562);
nor U2670 (N_2670,N_1742,N_1876);
nand U2671 (N_2671,N_1913,N_2205);
or U2672 (N_2672,N_1920,N_1925);
nor U2673 (N_2673,N_1782,N_1779);
xnor U2674 (N_2674,N_1503,N_1926);
and U2675 (N_2675,N_2170,N_1627);
nor U2676 (N_2676,N_1913,N_1516);
and U2677 (N_2677,N_2050,N_1824);
nor U2678 (N_2678,N_2033,N_1880);
xor U2679 (N_2679,N_1797,N_1506);
nand U2680 (N_2680,N_1511,N_1838);
nor U2681 (N_2681,N_2004,N_1764);
and U2682 (N_2682,N_2151,N_1974);
xor U2683 (N_2683,N_2065,N_1565);
nand U2684 (N_2684,N_1533,N_1819);
nor U2685 (N_2685,N_1914,N_1849);
nand U2686 (N_2686,N_1698,N_1837);
or U2687 (N_2687,N_1795,N_1513);
nor U2688 (N_2688,N_1503,N_1819);
nand U2689 (N_2689,N_1602,N_2083);
or U2690 (N_2690,N_1678,N_1889);
and U2691 (N_2691,N_1541,N_1821);
nand U2692 (N_2692,N_1726,N_2057);
and U2693 (N_2693,N_2027,N_1581);
nand U2694 (N_2694,N_1773,N_2226);
nor U2695 (N_2695,N_1860,N_2043);
xor U2696 (N_2696,N_1577,N_2216);
xor U2697 (N_2697,N_1874,N_1601);
nor U2698 (N_2698,N_1602,N_1741);
or U2699 (N_2699,N_1500,N_1829);
xor U2700 (N_2700,N_1506,N_2125);
or U2701 (N_2701,N_2170,N_1768);
nand U2702 (N_2702,N_1988,N_2156);
nand U2703 (N_2703,N_1672,N_1848);
and U2704 (N_2704,N_1610,N_1750);
and U2705 (N_2705,N_1797,N_1718);
nor U2706 (N_2706,N_2142,N_2168);
xnor U2707 (N_2707,N_1893,N_2103);
or U2708 (N_2708,N_2134,N_1826);
or U2709 (N_2709,N_2145,N_1802);
or U2710 (N_2710,N_1614,N_1770);
nand U2711 (N_2711,N_1565,N_2066);
and U2712 (N_2712,N_1624,N_1869);
or U2713 (N_2713,N_1779,N_1614);
or U2714 (N_2714,N_1871,N_2224);
nand U2715 (N_2715,N_1719,N_1796);
or U2716 (N_2716,N_1617,N_2048);
and U2717 (N_2717,N_1725,N_1516);
nand U2718 (N_2718,N_1611,N_1880);
or U2719 (N_2719,N_1952,N_2126);
and U2720 (N_2720,N_2096,N_1873);
or U2721 (N_2721,N_2193,N_1947);
nand U2722 (N_2722,N_1709,N_1796);
and U2723 (N_2723,N_2003,N_1740);
or U2724 (N_2724,N_2117,N_1907);
and U2725 (N_2725,N_2027,N_2037);
nand U2726 (N_2726,N_1634,N_2230);
and U2727 (N_2727,N_2249,N_1717);
nand U2728 (N_2728,N_2026,N_1815);
or U2729 (N_2729,N_1534,N_1887);
or U2730 (N_2730,N_1819,N_2014);
xor U2731 (N_2731,N_2113,N_2140);
xnor U2732 (N_2732,N_1605,N_2231);
or U2733 (N_2733,N_1983,N_1585);
nand U2734 (N_2734,N_2217,N_2238);
and U2735 (N_2735,N_1562,N_1686);
nand U2736 (N_2736,N_1646,N_1556);
xor U2737 (N_2737,N_1570,N_1501);
nor U2738 (N_2738,N_2230,N_1520);
nor U2739 (N_2739,N_2030,N_1933);
nand U2740 (N_2740,N_1968,N_1561);
nor U2741 (N_2741,N_1930,N_2161);
nand U2742 (N_2742,N_1543,N_2014);
nand U2743 (N_2743,N_2139,N_2078);
nor U2744 (N_2744,N_1503,N_2249);
and U2745 (N_2745,N_1618,N_1978);
and U2746 (N_2746,N_2244,N_1743);
and U2747 (N_2747,N_1790,N_1733);
or U2748 (N_2748,N_2137,N_1763);
nor U2749 (N_2749,N_1706,N_1796);
nor U2750 (N_2750,N_1688,N_2212);
nor U2751 (N_2751,N_2220,N_1940);
and U2752 (N_2752,N_2162,N_1869);
nand U2753 (N_2753,N_1781,N_1615);
nor U2754 (N_2754,N_1775,N_2065);
and U2755 (N_2755,N_2207,N_2153);
nand U2756 (N_2756,N_1827,N_2186);
and U2757 (N_2757,N_1918,N_2177);
or U2758 (N_2758,N_2061,N_1830);
and U2759 (N_2759,N_1648,N_1763);
or U2760 (N_2760,N_1514,N_2211);
nor U2761 (N_2761,N_1639,N_2204);
nand U2762 (N_2762,N_2163,N_1788);
xnor U2763 (N_2763,N_1633,N_2142);
xor U2764 (N_2764,N_1947,N_1733);
and U2765 (N_2765,N_1506,N_2057);
nor U2766 (N_2766,N_2209,N_2223);
or U2767 (N_2767,N_2159,N_1856);
or U2768 (N_2768,N_1730,N_2172);
and U2769 (N_2769,N_2035,N_2197);
nand U2770 (N_2770,N_1681,N_1695);
and U2771 (N_2771,N_2075,N_1781);
or U2772 (N_2772,N_1684,N_2128);
or U2773 (N_2773,N_2051,N_1746);
and U2774 (N_2774,N_1794,N_2136);
nor U2775 (N_2775,N_1924,N_1777);
xnor U2776 (N_2776,N_1548,N_1996);
nand U2777 (N_2777,N_2170,N_2205);
and U2778 (N_2778,N_1952,N_1939);
nor U2779 (N_2779,N_2093,N_1559);
or U2780 (N_2780,N_2207,N_2162);
and U2781 (N_2781,N_1996,N_2025);
or U2782 (N_2782,N_1733,N_1513);
and U2783 (N_2783,N_1706,N_1772);
or U2784 (N_2784,N_1897,N_1716);
nand U2785 (N_2785,N_2090,N_2055);
nor U2786 (N_2786,N_1588,N_1613);
and U2787 (N_2787,N_1963,N_1853);
nand U2788 (N_2788,N_1733,N_1927);
xor U2789 (N_2789,N_1959,N_1609);
nand U2790 (N_2790,N_1793,N_2217);
nand U2791 (N_2791,N_1859,N_1595);
nand U2792 (N_2792,N_1945,N_1746);
or U2793 (N_2793,N_2169,N_2246);
nand U2794 (N_2794,N_1965,N_2004);
or U2795 (N_2795,N_2233,N_1690);
nor U2796 (N_2796,N_2134,N_1586);
and U2797 (N_2797,N_1879,N_2204);
nor U2798 (N_2798,N_2203,N_1965);
or U2799 (N_2799,N_1972,N_1646);
or U2800 (N_2800,N_1891,N_2128);
and U2801 (N_2801,N_1862,N_1948);
nand U2802 (N_2802,N_2229,N_1579);
and U2803 (N_2803,N_2096,N_1858);
nand U2804 (N_2804,N_2133,N_1707);
or U2805 (N_2805,N_1865,N_1788);
nor U2806 (N_2806,N_1870,N_1829);
xnor U2807 (N_2807,N_1628,N_1597);
and U2808 (N_2808,N_1589,N_1577);
and U2809 (N_2809,N_1871,N_1883);
or U2810 (N_2810,N_2179,N_1831);
or U2811 (N_2811,N_1591,N_1953);
or U2812 (N_2812,N_2044,N_1684);
or U2813 (N_2813,N_1617,N_1836);
and U2814 (N_2814,N_1943,N_1820);
nand U2815 (N_2815,N_1639,N_1750);
nor U2816 (N_2816,N_1859,N_2092);
nor U2817 (N_2817,N_1793,N_1882);
xnor U2818 (N_2818,N_2072,N_1555);
nor U2819 (N_2819,N_1918,N_1979);
or U2820 (N_2820,N_1757,N_1798);
or U2821 (N_2821,N_2103,N_1914);
and U2822 (N_2822,N_1814,N_2063);
nand U2823 (N_2823,N_1895,N_1622);
and U2824 (N_2824,N_1914,N_1866);
nor U2825 (N_2825,N_1892,N_2058);
nor U2826 (N_2826,N_1849,N_2169);
nor U2827 (N_2827,N_1576,N_1996);
nor U2828 (N_2828,N_2122,N_1857);
nand U2829 (N_2829,N_2171,N_1724);
and U2830 (N_2830,N_2234,N_2133);
nor U2831 (N_2831,N_2117,N_1892);
or U2832 (N_2832,N_1930,N_1866);
or U2833 (N_2833,N_2130,N_2045);
and U2834 (N_2834,N_2224,N_1665);
and U2835 (N_2835,N_1862,N_1796);
nand U2836 (N_2836,N_1943,N_2085);
or U2837 (N_2837,N_2136,N_1680);
nor U2838 (N_2838,N_2061,N_1874);
nor U2839 (N_2839,N_1577,N_1595);
or U2840 (N_2840,N_1991,N_1578);
and U2841 (N_2841,N_1976,N_2120);
nor U2842 (N_2842,N_1754,N_2243);
and U2843 (N_2843,N_2211,N_1953);
or U2844 (N_2844,N_1998,N_1931);
or U2845 (N_2845,N_2021,N_1611);
nor U2846 (N_2846,N_1618,N_1523);
and U2847 (N_2847,N_1825,N_1642);
xor U2848 (N_2848,N_1972,N_2000);
and U2849 (N_2849,N_2070,N_1792);
or U2850 (N_2850,N_2109,N_1663);
nand U2851 (N_2851,N_1973,N_2196);
nand U2852 (N_2852,N_1826,N_1663);
nand U2853 (N_2853,N_1576,N_1946);
nand U2854 (N_2854,N_1845,N_2032);
nand U2855 (N_2855,N_2197,N_1665);
and U2856 (N_2856,N_1549,N_1716);
and U2857 (N_2857,N_2152,N_1586);
and U2858 (N_2858,N_1978,N_1716);
nor U2859 (N_2859,N_1605,N_1767);
and U2860 (N_2860,N_2116,N_1835);
nor U2861 (N_2861,N_1735,N_1923);
and U2862 (N_2862,N_1564,N_1933);
nand U2863 (N_2863,N_1730,N_2030);
nand U2864 (N_2864,N_1835,N_1693);
nand U2865 (N_2865,N_1937,N_1670);
and U2866 (N_2866,N_2094,N_1646);
and U2867 (N_2867,N_1584,N_2187);
nand U2868 (N_2868,N_1738,N_1732);
nor U2869 (N_2869,N_1672,N_1996);
and U2870 (N_2870,N_2080,N_1836);
nor U2871 (N_2871,N_1820,N_1545);
nand U2872 (N_2872,N_2133,N_1799);
xor U2873 (N_2873,N_1595,N_1811);
or U2874 (N_2874,N_2223,N_1637);
nor U2875 (N_2875,N_1675,N_1574);
or U2876 (N_2876,N_1644,N_1706);
nor U2877 (N_2877,N_1932,N_1589);
and U2878 (N_2878,N_1787,N_2120);
and U2879 (N_2879,N_1681,N_1766);
nand U2880 (N_2880,N_2112,N_2131);
or U2881 (N_2881,N_2207,N_1901);
or U2882 (N_2882,N_1762,N_1700);
xor U2883 (N_2883,N_2087,N_2120);
nand U2884 (N_2884,N_2021,N_2083);
nand U2885 (N_2885,N_1616,N_1710);
xnor U2886 (N_2886,N_1959,N_1694);
xnor U2887 (N_2887,N_2124,N_2147);
and U2888 (N_2888,N_1691,N_1500);
and U2889 (N_2889,N_2236,N_1503);
nor U2890 (N_2890,N_1804,N_2023);
nor U2891 (N_2891,N_1608,N_1856);
nor U2892 (N_2892,N_1688,N_1787);
nand U2893 (N_2893,N_1885,N_2143);
xor U2894 (N_2894,N_1969,N_1809);
nor U2895 (N_2895,N_1695,N_2056);
or U2896 (N_2896,N_1574,N_1725);
xnor U2897 (N_2897,N_2057,N_1909);
xor U2898 (N_2898,N_1941,N_1817);
nor U2899 (N_2899,N_2113,N_1777);
and U2900 (N_2900,N_2242,N_2190);
nor U2901 (N_2901,N_1621,N_1569);
or U2902 (N_2902,N_2015,N_1696);
nor U2903 (N_2903,N_1654,N_2120);
or U2904 (N_2904,N_1809,N_2192);
or U2905 (N_2905,N_2075,N_1872);
xnor U2906 (N_2906,N_1613,N_1751);
nand U2907 (N_2907,N_2062,N_1835);
and U2908 (N_2908,N_1963,N_1836);
nor U2909 (N_2909,N_2120,N_1642);
nand U2910 (N_2910,N_1577,N_1746);
nor U2911 (N_2911,N_1880,N_1705);
and U2912 (N_2912,N_2157,N_1551);
xnor U2913 (N_2913,N_1780,N_1880);
or U2914 (N_2914,N_2132,N_1881);
or U2915 (N_2915,N_1949,N_2147);
or U2916 (N_2916,N_2100,N_1672);
and U2917 (N_2917,N_1847,N_1915);
and U2918 (N_2918,N_1630,N_1814);
nor U2919 (N_2919,N_2181,N_2217);
and U2920 (N_2920,N_2180,N_1758);
nand U2921 (N_2921,N_2235,N_1672);
and U2922 (N_2922,N_1563,N_1546);
nand U2923 (N_2923,N_1624,N_1967);
nor U2924 (N_2924,N_1749,N_1642);
and U2925 (N_2925,N_1647,N_1890);
and U2926 (N_2926,N_2027,N_1598);
nand U2927 (N_2927,N_1684,N_1916);
xnor U2928 (N_2928,N_2033,N_1665);
or U2929 (N_2929,N_2238,N_1917);
or U2930 (N_2930,N_1518,N_1795);
xor U2931 (N_2931,N_2025,N_1928);
or U2932 (N_2932,N_2188,N_1547);
or U2933 (N_2933,N_1756,N_1590);
xnor U2934 (N_2934,N_2040,N_2242);
nand U2935 (N_2935,N_1559,N_1548);
and U2936 (N_2936,N_1798,N_1667);
nor U2937 (N_2937,N_1742,N_2222);
or U2938 (N_2938,N_1965,N_1786);
nand U2939 (N_2939,N_1782,N_2163);
or U2940 (N_2940,N_1655,N_1975);
nor U2941 (N_2941,N_2129,N_1505);
or U2942 (N_2942,N_1596,N_1738);
and U2943 (N_2943,N_1766,N_1780);
and U2944 (N_2944,N_1722,N_1789);
nand U2945 (N_2945,N_1700,N_2174);
or U2946 (N_2946,N_2105,N_1981);
and U2947 (N_2947,N_1554,N_1711);
nand U2948 (N_2948,N_1696,N_1644);
nor U2949 (N_2949,N_1654,N_1591);
xor U2950 (N_2950,N_1526,N_1621);
nor U2951 (N_2951,N_1521,N_2109);
and U2952 (N_2952,N_2009,N_1656);
nor U2953 (N_2953,N_1669,N_2003);
and U2954 (N_2954,N_2073,N_1594);
nor U2955 (N_2955,N_1550,N_1820);
nand U2956 (N_2956,N_1859,N_1974);
nand U2957 (N_2957,N_2163,N_1741);
or U2958 (N_2958,N_2187,N_2034);
or U2959 (N_2959,N_1599,N_1533);
and U2960 (N_2960,N_2232,N_1966);
or U2961 (N_2961,N_1694,N_2141);
xnor U2962 (N_2962,N_1565,N_1576);
nor U2963 (N_2963,N_1885,N_1964);
or U2964 (N_2964,N_1946,N_2135);
and U2965 (N_2965,N_2138,N_1897);
or U2966 (N_2966,N_2196,N_1703);
nor U2967 (N_2967,N_1851,N_1538);
nor U2968 (N_2968,N_1928,N_2119);
and U2969 (N_2969,N_1667,N_1633);
or U2970 (N_2970,N_1520,N_1626);
nor U2971 (N_2971,N_1582,N_2227);
or U2972 (N_2972,N_1694,N_2219);
xnor U2973 (N_2973,N_2145,N_1589);
xor U2974 (N_2974,N_1771,N_1805);
and U2975 (N_2975,N_2059,N_2073);
nor U2976 (N_2976,N_1984,N_2104);
nand U2977 (N_2977,N_2107,N_2243);
nand U2978 (N_2978,N_2201,N_2233);
and U2979 (N_2979,N_2109,N_1743);
nand U2980 (N_2980,N_1855,N_1757);
and U2981 (N_2981,N_2073,N_2149);
nand U2982 (N_2982,N_1980,N_1743);
and U2983 (N_2983,N_1559,N_1840);
or U2984 (N_2984,N_1798,N_1696);
and U2985 (N_2985,N_2070,N_2071);
nor U2986 (N_2986,N_1522,N_2114);
and U2987 (N_2987,N_2129,N_2056);
and U2988 (N_2988,N_1608,N_1822);
nand U2989 (N_2989,N_1717,N_1920);
nand U2990 (N_2990,N_2240,N_1599);
nor U2991 (N_2991,N_2243,N_1640);
nand U2992 (N_2992,N_2198,N_1721);
or U2993 (N_2993,N_1585,N_2186);
or U2994 (N_2994,N_2090,N_2249);
nand U2995 (N_2995,N_1874,N_2043);
nand U2996 (N_2996,N_2011,N_1858);
xor U2997 (N_2997,N_1871,N_1829);
and U2998 (N_2998,N_1519,N_1684);
xnor U2999 (N_2999,N_1971,N_1917);
nand UO_0 (O_0,N_2920,N_2679);
or UO_1 (O_1,N_2922,N_2762);
and UO_2 (O_2,N_2828,N_2687);
or UO_3 (O_3,N_2819,N_2694);
or UO_4 (O_4,N_2529,N_2989);
or UO_5 (O_5,N_2788,N_2881);
or UO_6 (O_6,N_2923,N_2314);
xor UO_7 (O_7,N_2611,N_2477);
nand UO_8 (O_8,N_2421,N_2478);
nor UO_9 (O_9,N_2897,N_2970);
nand UO_10 (O_10,N_2791,N_2531);
nand UO_11 (O_11,N_2825,N_2340);
xor UO_12 (O_12,N_2524,N_2842);
and UO_13 (O_13,N_2290,N_2304);
and UO_14 (O_14,N_2625,N_2769);
nor UO_15 (O_15,N_2583,N_2732);
and UO_16 (O_16,N_2849,N_2676);
and UO_17 (O_17,N_2398,N_2467);
nand UO_18 (O_18,N_2746,N_2269);
or UO_19 (O_19,N_2725,N_2628);
and UO_20 (O_20,N_2613,N_2723);
nor UO_21 (O_21,N_2609,N_2466);
or UO_22 (O_22,N_2593,N_2312);
nand UO_23 (O_23,N_2615,N_2858);
or UO_24 (O_24,N_2502,N_2517);
nand UO_25 (O_25,N_2281,N_2957);
or UO_26 (O_26,N_2992,N_2298);
or UO_27 (O_27,N_2480,N_2802);
nand UO_28 (O_28,N_2864,N_2280);
nor UO_29 (O_29,N_2322,N_2665);
nor UO_30 (O_30,N_2379,N_2815);
nor UO_31 (O_31,N_2258,N_2488);
nor UO_32 (O_32,N_2342,N_2595);
nor UO_33 (O_33,N_2397,N_2677);
nor UO_34 (O_34,N_2741,N_2614);
or UO_35 (O_35,N_2737,N_2689);
nor UO_36 (O_36,N_2945,N_2977);
and UO_37 (O_37,N_2823,N_2297);
or UO_38 (O_38,N_2981,N_2994);
and UO_39 (O_39,N_2630,N_2956);
nor UO_40 (O_40,N_2429,N_2303);
xnor UO_41 (O_41,N_2939,N_2797);
nand UO_42 (O_42,N_2460,N_2526);
or UO_43 (O_43,N_2446,N_2926);
xnor UO_44 (O_44,N_2890,N_2867);
or UO_45 (O_45,N_2377,N_2557);
or UO_46 (O_46,N_2693,N_2866);
and UO_47 (O_47,N_2899,N_2461);
or UO_48 (O_48,N_2913,N_2711);
xnor UO_49 (O_49,N_2728,N_2577);
xnor UO_50 (O_50,N_2410,N_2789);
or UO_51 (O_51,N_2395,N_2950);
xnor UO_52 (O_52,N_2877,N_2492);
and UO_53 (O_53,N_2850,N_2841);
nand UO_54 (O_54,N_2617,N_2982);
and UO_55 (O_55,N_2779,N_2387);
or UO_56 (O_56,N_2715,N_2562);
nor UO_57 (O_57,N_2589,N_2515);
or UO_58 (O_58,N_2808,N_2293);
nor UO_59 (O_59,N_2958,N_2855);
nand UO_60 (O_60,N_2766,N_2471);
nand UO_61 (O_61,N_2836,N_2424);
nand UO_62 (O_62,N_2869,N_2306);
and UO_63 (O_63,N_2636,N_2390);
nand UO_64 (O_64,N_2868,N_2282);
and UO_65 (O_65,N_2938,N_2464);
or UO_66 (O_66,N_2667,N_2697);
nor UO_67 (O_67,N_2454,N_2742);
or UO_68 (O_68,N_2533,N_2400);
and UO_69 (O_69,N_2432,N_2498);
nand UO_70 (O_70,N_2317,N_2835);
nand UO_71 (O_71,N_2627,N_2642);
and UO_72 (O_72,N_2556,N_2635);
and UO_73 (O_73,N_2680,N_2599);
nand UO_74 (O_74,N_2942,N_2428);
nand UO_75 (O_75,N_2907,N_2946);
and UO_76 (O_76,N_2817,N_2829);
nor UO_77 (O_77,N_2623,N_2986);
or UO_78 (O_78,N_2404,N_2278);
and UO_79 (O_79,N_2575,N_2504);
or UO_80 (O_80,N_2494,N_2873);
nor UO_81 (O_81,N_2479,N_2933);
and UO_82 (O_82,N_2417,N_2536);
or UO_83 (O_83,N_2339,N_2323);
or UO_84 (O_84,N_2754,N_2500);
or UO_85 (O_85,N_2853,N_2931);
and UO_86 (O_86,N_2389,N_2704);
or UO_87 (O_87,N_2888,N_2580);
and UO_88 (O_88,N_2261,N_2618);
and UO_89 (O_89,N_2541,N_2772);
or UO_90 (O_90,N_2889,N_2846);
nand UO_91 (O_91,N_2394,N_2987);
and UO_92 (O_92,N_2646,N_2528);
and UO_93 (O_93,N_2874,N_2978);
and UO_94 (O_94,N_2594,N_2326);
nand UO_95 (O_95,N_2671,N_2784);
nand UO_96 (O_96,N_2554,N_2796);
or UO_97 (O_97,N_2684,N_2639);
and UO_98 (O_98,N_2449,N_2940);
nor UO_99 (O_99,N_2718,N_2380);
nand UO_100 (O_100,N_2329,N_2925);
xor UO_101 (O_101,N_2979,N_2906);
nand UO_102 (O_102,N_2356,N_2993);
nand UO_103 (O_103,N_2706,N_2672);
nand UO_104 (O_104,N_2837,N_2810);
nor UO_105 (O_105,N_2337,N_2727);
or UO_106 (O_106,N_2807,N_2696);
and UO_107 (O_107,N_2674,N_2255);
xnor UO_108 (O_108,N_2457,N_2830);
or UO_109 (O_109,N_2903,N_2820);
or UO_110 (O_110,N_2512,N_2943);
nand UO_111 (O_111,N_2730,N_2681);
or UO_112 (O_112,N_2288,N_2844);
xnor UO_113 (O_113,N_2341,N_2425);
nand UO_114 (O_114,N_2909,N_2682);
or UO_115 (O_115,N_2451,N_2717);
nor UO_116 (O_116,N_2590,N_2756);
and UO_117 (O_117,N_2947,N_2904);
xnor UO_118 (O_118,N_2537,N_2546);
nor UO_119 (O_119,N_2521,N_2900);
nor UO_120 (O_120,N_2362,N_2259);
xnor UO_121 (O_121,N_2438,N_2721);
or UO_122 (O_122,N_2710,N_2882);
nand UO_123 (O_123,N_2731,N_2893);
or UO_124 (O_124,N_2865,N_2364);
or UO_125 (O_125,N_2770,N_2499);
xnor UO_126 (O_126,N_2649,N_2840);
nand UO_127 (O_127,N_2405,N_2313);
nor UO_128 (O_128,N_2690,N_2937);
and UO_129 (O_129,N_2481,N_2491);
nor UO_130 (O_130,N_2700,N_2980);
or UO_131 (O_131,N_2824,N_2547);
nor UO_132 (O_132,N_2738,N_2474);
and UO_133 (O_133,N_2476,N_2863);
and UO_134 (O_134,N_2596,N_2365);
nand UO_135 (O_135,N_2431,N_2932);
or UO_136 (O_136,N_2875,N_2834);
nand UO_137 (O_137,N_2445,N_2332);
xor UO_138 (O_138,N_2487,N_2964);
nor UO_139 (O_139,N_2921,N_2252);
or UO_140 (O_140,N_2386,N_2503);
and UO_141 (O_141,N_2335,N_2525);
or UO_142 (O_142,N_2299,N_2654);
nor UO_143 (O_143,N_2582,N_2702);
and UO_144 (O_144,N_2442,N_2780);
nor UO_145 (O_145,N_2607,N_2415);
xor UO_146 (O_146,N_2871,N_2826);
nor UO_147 (O_147,N_2734,N_2917);
and UO_148 (O_148,N_2886,N_2523);
nand UO_149 (O_149,N_2407,N_2578);
xnor UO_150 (O_150,N_2744,N_2751);
nand UO_151 (O_151,N_2565,N_2894);
or UO_152 (O_152,N_2378,N_2602);
and UO_153 (O_153,N_2287,N_2847);
and UO_154 (O_154,N_2396,N_2475);
and UO_155 (O_155,N_2719,N_2345);
nand UO_156 (O_156,N_2321,N_2934);
nor UO_157 (O_157,N_2972,N_2427);
or UO_158 (O_158,N_2600,N_2967);
nand UO_159 (O_159,N_2912,N_2505);
and UO_160 (O_160,N_2453,N_2966);
xor UO_161 (O_161,N_2643,N_2857);
or UO_162 (O_162,N_2308,N_2413);
or UO_163 (O_163,N_2485,N_2567);
and UO_164 (O_164,N_2902,N_2859);
or UO_165 (O_165,N_2519,N_2709);
and UO_166 (O_166,N_2291,N_2539);
nand UO_167 (O_167,N_2419,N_2349);
nor UO_168 (O_168,N_2898,N_2358);
nor UO_169 (O_169,N_2579,N_2535);
nand UO_170 (O_170,N_2765,N_2722);
and UO_171 (O_171,N_2253,N_2587);
xnor UO_172 (O_172,N_2891,N_2975);
nand UO_173 (O_173,N_2801,N_2763);
xor UO_174 (O_174,N_2436,N_2566);
and UO_175 (O_175,N_2352,N_2591);
nand UO_176 (O_176,N_2574,N_2666);
nand UO_177 (O_177,N_2959,N_2838);
xor UO_178 (O_178,N_2716,N_2344);
nor UO_179 (O_179,N_2509,N_2520);
nand UO_180 (O_180,N_2692,N_2930);
nor UO_181 (O_181,N_2990,N_2759);
and UO_182 (O_182,N_2729,N_2648);
nor UO_183 (O_183,N_2373,N_2402);
nand UO_184 (O_184,N_2929,N_2270);
or UO_185 (O_185,N_2799,N_2265);
nor UO_186 (O_186,N_2792,N_2441);
xor UO_187 (O_187,N_2532,N_2678);
and UO_188 (O_188,N_2581,N_2250);
nor UO_189 (O_189,N_2918,N_2862);
or UO_190 (O_190,N_2610,N_2560);
and UO_191 (O_191,N_2507,N_2330);
nand UO_192 (O_192,N_2805,N_2758);
xnor UO_193 (O_193,N_2576,N_2668);
nor UO_194 (O_194,N_2622,N_2385);
nand UO_195 (O_195,N_2391,N_2334);
nand UO_196 (O_196,N_2786,N_2750);
or UO_197 (O_197,N_2658,N_2310);
nor UO_198 (O_198,N_2971,N_2673);
nand UO_199 (O_199,N_2634,N_2775);
nand UO_200 (O_200,N_2496,N_2916);
nor UO_201 (O_201,N_2739,N_2604);
or UO_202 (O_202,N_2274,N_2256);
nand UO_203 (O_203,N_2354,N_2953);
or UO_204 (O_204,N_2851,N_2490);
and UO_205 (O_205,N_2724,N_2559);
nand UO_206 (O_206,N_2418,N_2254);
or UO_207 (O_207,N_2495,N_2586);
nor UO_208 (O_208,N_2936,N_2448);
nand UO_209 (O_209,N_2887,N_2659);
and UO_210 (O_210,N_2663,N_2695);
or UO_211 (O_211,N_2661,N_2435);
nor UO_212 (O_212,N_2497,N_2621);
nand UO_213 (O_213,N_2908,N_2414);
xnor UO_214 (O_214,N_2462,N_2371);
and UO_215 (O_215,N_2292,N_2773);
nor UO_216 (O_216,N_2878,N_2279);
and UO_217 (O_217,N_2713,N_2571);
nand UO_218 (O_218,N_2633,N_2827);
xnor UO_219 (O_219,N_2263,N_2753);
nor UO_220 (O_220,N_2800,N_2375);
or UO_221 (O_221,N_2264,N_2703);
nor UO_222 (O_222,N_2434,N_2319);
xor UO_223 (O_223,N_2736,N_2455);
nand UO_224 (O_224,N_2311,N_2359);
nand UO_225 (O_225,N_2914,N_2315);
and UO_226 (O_226,N_2876,N_2708);
nand UO_227 (O_227,N_2748,N_2508);
and UO_228 (O_228,N_2289,N_2584);
or UO_229 (O_229,N_2821,N_2403);
nor UO_230 (O_230,N_2656,N_2774);
and UO_231 (O_231,N_2804,N_2300);
nor UO_232 (O_232,N_2440,N_2657);
or UO_233 (O_233,N_2423,N_2670);
or UO_234 (O_234,N_2752,N_2782);
or UO_235 (O_235,N_2486,N_2941);
nand UO_236 (O_236,N_2733,N_2472);
or UO_237 (O_237,N_2861,N_2412);
xor UO_238 (O_238,N_2527,N_2569);
and UO_239 (O_239,N_2483,N_2901);
nand UO_240 (O_240,N_2470,N_2585);
or UO_241 (O_241,N_2608,N_2601);
and UO_242 (O_242,N_2845,N_2372);
or UO_243 (O_243,N_2411,N_2384);
or UO_244 (O_244,N_2776,N_2641);
nor UO_245 (O_245,N_2856,N_2948);
or UO_246 (O_246,N_2885,N_2691);
nor UO_247 (O_247,N_2701,N_2388);
or UO_248 (O_248,N_2745,N_2551);
nand UO_249 (O_249,N_2338,N_2698);
nand UO_250 (O_250,N_2976,N_2284);
nor UO_251 (O_251,N_2785,N_2333);
nand UO_252 (O_252,N_2570,N_2652);
nor UO_253 (O_253,N_2433,N_2675);
and UO_254 (O_254,N_2381,N_2927);
nand UO_255 (O_255,N_2619,N_2416);
nand UO_256 (O_256,N_2951,N_2268);
and UO_257 (O_257,N_2283,N_2647);
nand UO_258 (O_258,N_2473,N_2767);
nor UO_259 (O_259,N_2518,N_2818);
or UO_260 (O_260,N_2852,N_2355);
nand UO_261 (O_261,N_2795,N_2812);
and UO_262 (O_262,N_2357,N_2257);
and UO_263 (O_263,N_2757,N_2624);
and UO_264 (O_264,N_2777,N_2809);
and UO_265 (O_265,N_2296,N_2392);
nor UO_266 (O_266,N_2870,N_2353);
or UO_267 (O_267,N_2811,N_2638);
nand UO_268 (O_268,N_2458,N_2463);
nand UO_269 (O_269,N_2251,N_2530);
or UO_270 (O_270,N_2318,N_2720);
or UO_271 (O_271,N_2879,N_2437);
xor UO_272 (O_272,N_2960,N_2267);
or UO_273 (O_273,N_2640,N_2984);
nor UO_274 (O_274,N_2563,N_2749);
and UO_275 (O_275,N_2266,N_2983);
or UO_276 (O_276,N_2998,N_2309);
and UO_277 (O_277,N_2631,N_2272);
or UO_278 (O_278,N_2285,N_2988);
nand UO_279 (O_279,N_2793,N_2409);
nor UO_280 (O_280,N_2360,N_2771);
and UO_281 (O_281,N_2714,N_2644);
nand UO_282 (O_282,N_2803,N_2555);
nor UO_283 (O_283,N_2949,N_2952);
or UO_284 (O_284,N_2707,N_2383);
nor UO_285 (O_285,N_2393,N_2798);
xor UO_286 (O_286,N_2598,N_2343);
xor UO_287 (O_287,N_2944,N_2895);
xor UO_288 (O_288,N_2832,N_2295);
nor UO_289 (O_289,N_2626,N_2833);
nor UO_290 (O_290,N_2962,N_2974);
nand UO_291 (O_291,N_2511,N_2406);
nor UO_292 (O_292,N_2860,N_2735);
or UO_293 (O_293,N_2561,N_2327);
and UO_294 (O_294,N_2726,N_2336);
and UO_295 (O_295,N_2740,N_2655);
and UO_296 (O_296,N_2420,N_2513);
nor UO_297 (O_297,N_2376,N_2346);
and UO_298 (O_298,N_2260,N_2848);
or UO_299 (O_299,N_2361,N_2493);
and UO_300 (O_300,N_2506,N_2294);
nand UO_301 (O_301,N_2629,N_2331);
nor UO_302 (O_302,N_2664,N_2854);
nand UO_303 (O_303,N_2540,N_2347);
or UO_304 (O_304,N_2761,N_2790);
xor UO_305 (O_305,N_2307,N_2568);
nor UO_306 (O_306,N_2305,N_2538);
and UO_307 (O_307,N_2603,N_2549);
nand UO_308 (O_308,N_2426,N_2928);
nand UO_309 (O_309,N_2370,N_2348);
nor UO_310 (O_310,N_2778,N_2822);
and UO_311 (O_311,N_2351,N_2382);
and UO_312 (O_312,N_2262,N_2366);
and UO_313 (O_313,N_2915,N_2456);
nand UO_314 (O_314,N_2880,N_2367);
xor UO_315 (O_315,N_2831,N_2685);
and UO_316 (O_316,N_2363,N_2872);
nor UO_317 (O_317,N_2616,N_2650);
nor UO_318 (O_318,N_2401,N_2408);
or UO_319 (O_319,N_2787,N_2764);
nand UO_320 (O_320,N_2516,N_2459);
or UO_321 (O_321,N_2910,N_2896);
xor UO_322 (O_322,N_2997,N_2452);
and UO_323 (O_323,N_2969,N_2606);
xnor UO_324 (O_324,N_2919,N_2422);
or UO_325 (O_325,N_2374,N_2905);
and UO_326 (O_326,N_2605,N_2522);
nor UO_327 (O_327,N_2892,N_2443);
and UO_328 (O_328,N_2686,N_2705);
and UO_329 (O_329,N_2325,N_2883);
and UO_330 (O_330,N_2924,N_2839);
or UO_331 (O_331,N_2683,N_2688);
nor UO_332 (O_332,N_2301,N_2843);
nor UO_333 (O_333,N_2302,N_2545);
and UO_334 (O_334,N_2469,N_2743);
and UO_335 (O_335,N_2286,N_2813);
nand UO_336 (O_336,N_2632,N_2465);
nand UO_337 (O_337,N_2548,N_2399);
or UO_338 (O_338,N_2999,N_2955);
nor UO_339 (O_339,N_2328,N_2514);
nand UO_340 (O_340,N_2996,N_2447);
and UO_341 (O_341,N_2482,N_2275);
nand UO_342 (O_342,N_2573,N_2592);
nand UO_343 (O_343,N_2669,N_2814);
nor UO_344 (O_344,N_2645,N_2369);
nor UO_345 (O_345,N_2651,N_2510);
and UO_346 (O_346,N_2324,N_2542);
nor UO_347 (O_347,N_2350,N_2965);
nand UO_348 (O_348,N_2662,N_2783);
nand UO_349 (O_349,N_2501,N_2712);
or UO_350 (O_350,N_2755,N_2768);
nor UO_351 (O_351,N_2781,N_2273);
nor UO_352 (O_352,N_2572,N_2430);
nand UO_353 (O_353,N_2884,N_2816);
or UO_354 (O_354,N_2991,N_2954);
or UO_355 (O_355,N_2973,N_2484);
xor UO_356 (O_356,N_2550,N_2489);
and UO_357 (O_357,N_2316,N_2653);
or UO_358 (O_358,N_2534,N_2368);
and UO_359 (O_359,N_2450,N_2637);
nand UO_360 (O_360,N_2544,N_2620);
nor UO_361 (O_361,N_2935,N_2271);
and UO_362 (O_362,N_2564,N_2699);
and UO_363 (O_363,N_2961,N_2320);
nand UO_364 (O_364,N_2660,N_2588);
nor UO_365 (O_365,N_2963,N_2985);
nand UO_366 (O_366,N_2552,N_2612);
and UO_367 (O_367,N_2468,N_2553);
nand UO_368 (O_368,N_2543,N_2806);
nor UO_369 (O_369,N_2968,N_2276);
and UO_370 (O_370,N_2995,N_2558);
xnor UO_371 (O_371,N_2444,N_2277);
nor UO_372 (O_372,N_2760,N_2794);
nor UO_373 (O_373,N_2911,N_2747);
nor UO_374 (O_374,N_2597,N_2439);
and UO_375 (O_375,N_2438,N_2707);
nand UO_376 (O_376,N_2899,N_2253);
nor UO_377 (O_377,N_2437,N_2927);
or UO_378 (O_378,N_2782,N_2680);
and UO_379 (O_379,N_2535,N_2952);
nand UO_380 (O_380,N_2503,N_2276);
nor UO_381 (O_381,N_2960,N_2840);
nor UO_382 (O_382,N_2414,N_2404);
nor UO_383 (O_383,N_2405,N_2967);
nand UO_384 (O_384,N_2260,N_2568);
nand UO_385 (O_385,N_2302,N_2539);
and UO_386 (O_386,N_2258,N_2460);
nand UO_387 (O_387,N_2805,N_2380);
nand UO_388 (O_388,N_2985,N_2704);
nand UO_389 (O_389,N_2912,N_2847);
or UO_390 (O_390,N_2546,N_2421);
nor UO_391 (O_391,N_2612,N_2657);
nand UO_392 (O_392,N_2471,N_2684);
and UO_393 (O_393,N_2476,N_2302);
and UO_394 (O_394,N_2353,N_2474);
and UO_395 (O_395,N_2487,N_2565);
and UO_396 (O_396,N_2458,N_2436);
or UO_397 (O_397,N_2297,N_2332);
nor UO_398 (O_398,N_2625,N_2862);
nand UO_399 (O_399,N_2679,N_2859);
or UO_400 (O_400,N_2281,N_2463);
nor UO_401 (O_401,N_2941,N_2993);
or UO_402 (O_402,N_2692,N_2753);
or UO_403 (O_403,N_2725,N_2825);
or UO_404 (O_404,N_2917,N_2939);
or UO_405 (O_405,N_2542,N_2377);
nor UO_406 (O_406,N_2448,N_2999);
nor UO_407 (O_407,N_2658,N_2486);
nand UO_408 (O_408,N_2539,N_2840);
or UO_409 (O_409,N_2843,N_2298);
and UO_410 (O_410,N_2827,N_2587);
xnor UO_411 (O_411,N_2621,N_2946);
nor UO_412 (O_412,N_2430,N_2271);
or UO_413 (O_413,N_2865,N_2313);
nor UO_414 (O_414,N_2276,N_2408);
and UO_415 (O_415,N_2319,N_2779);
or UO_416 (O_416,N_2468,N_2313);
nor UO_417 (O_417,N_2314,N_2915);
nand UO_418 (O_418,N_2905,N_2681);
nand UO_419 (O_419,N_2391,N_2921);
and UO_420 (O_420,N_2894,N_2793);
and UO_421 (O_421,N_2739,N_2341);
nor UO_422 (O_422,N_2493,N_2266);
and UO_423 (O_423,N_2616,N_2983);
nand UO_424 (O_424,N_2496,N_2984);
or UO_425 (O_425,N_2360,N_2414);
nand UO_426 (O_426,N_2400,N_2728);
nor UO_427 (O_427,N_2735,N_2802);
xnor UO_428 (O_428,N_2637,N_2872);
nand UO_429 (O_429,N_2602,N_2281);
and UO_430 (O_430,N_2688,N_2725);
nand UO_431 (O_431,N_2333,N_2530);
nor UO_432 (O_432,N_2553,N_2490);
or UO_433 (O_433,N_2542,N_2434);
or UO_434 (O_434,N_2531,N_2869);
or UO_435 (O_435,N_2321,N_2431);
and UO_436 (O_436,N_2550,N_2314);
and UO_437 (O_437,N_2910,N_2974);
or UO_438 (O_438,N_2624,N_2789);
and UO_439 (O_439,N_2267,N_2619);
nor UO_440 (O_440,N_2695,N_2484);
nor UO_441 (O_441,N_2775,N_2337);
or UO_442 (O_442,N_2760,N_2622);
or UO_443 (O_443,N_2766,N_2666);
nor UO_444 (O_444,N_2949,N_2872);
xnor UO_445 (O_445,N_2283,N_2534);
nor UO_446 (O_446,N_2601,N_2907);
nand UO_447 (O_447,N_2606,N_2531);
nand UO_448 (O_448,N_2288,N_2675);
and UO_449 (O_449,N_2727,N_2926);
xnor UO_450 (O_450,N_2942,N_2449);
nor UO_451 (O_451,N_2840,N_2694);
and UO_452 (O_452,N_2334,N_2536);
nand UO_453 (O_453,N_2300,N_2463);
xnor UO_454 (O_454,N_2404,N_2321);
xnor UO_455 (O_455,N_2281,N_2405);
or UO_456 (O_456,N_2622,N_2604);
nor UO_457 (O_457,N_2520,N_2414);
nor UO_458 (O_458,N_2750,N_2961);
nor UO_459 (O_459,N_2616,N_2662);
or UO_460 (O_460,N_2803,N_2374);
nand UO_461 (O_461,N_2391,N_2493);
and UO_462 (O_462,N_2866,N_2854);
nor UO_463 (O_463,N_2684,N_2870);
nor UO_464 (O_464,N_2417,N_2385);
nand UO_465 (O_465,N_2442,N_2282);
or UO_466 (O_466,N_2528,N_2966);
nand UO_467 (O_467,N_2684,N_2875);
nand UO_468 (O_468,N_2926,N_2277);
nand UO_469 (O_469,N_2721,N_2770);
or UO_470 (O_470,N_2802,N_2443);
nand UO_471 (O_471,N_2810,N_2429);
nand UO_472 (O_472,N_2445,N_2378);
xnor UO_473 (O_473,N_2673,N_2833);
and UO_474 (O_474,N_2255,N_2930);
and UO_475 (O_475,N_2910,N_2726);
or UO_476 (O_476,N_2504,N_2444);
nand UO_477 (O_477,N_2772,N_2444);
nand UO_478 (O_478,N_2715,N_2681);
nor UO_479 (O_479,N_2625,N_2258);
nor UO_480 (O_480,N_2981,N_2308);
nand UO_481 (O_481,N_2862,N_2676);
nand UO_482 (O_482,N_2301,N_2874);
nor UO_483 (O_483,N_2961,N_2870);
nand UO_484 (O_484,N_2509,N_2326);
xor UO_485 (O_485,N_2809,N_2988);
nand UO_486 (O_486,N_2496,N_2670);
xnor UO_487 (O_487,N_2882,N_2842);
xnor UO_488 (O_488,N_2893,N_2773);
or UO_489 (O_489,N_2694,N_2946);
xor UO_490 (O_490,N_2742,N_2942);
or UO_491 (O_491,N_2338,N_2604);
nor UO_492 (O_492,N_2739,N_2299);
or UO_493 (O_493,N_2505,N_2758);
xor UO_494 (O_494,N_2277,N_2487);
and UO_495 (O_495,N_2672,N_2519);
xor UO_496 (O_496,N_2387,N_2990);
or UO_497 (O_497,N_2365,N_2516);
nor UO_498 (O_498,N_2804,N_2486);
or UO_499 (O_499,N_2298,N_2741);
endmodule