module basic_500_3000_500_15_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_33,In_402);
or U1 (N_1,In_309,In_4);
or U2 (N_2,In_274,In_186);
or U3 (N_3,In_269,In_146);
nand U4 (N_4,In_130,In_190);
nand U5 (N_5,In_387,In_127);
nor U6 (N_6,In_247,In_404);
or U7 (N_7,In_494,In_430);
nand U8 (N_8,In_306,In_480);
or U9 (N_9,In_245,In_40);
nor U10 (N_10,In_117,In_482);
and U11 (N_11,In_357,In_272);
and U12 (N_12,In_23,In_453);
nand U13 (N_13,In_188,In_162);
nand U14 (N_14,In_267,In_458);
and U15 (N_15,In_429,In_213);
nand U16 (N_16,In_3,In_340);
or U17 (N_17,In_37,In_449);
nor U18 (N_18,In_165,In_184);
nor U19 (N_19,In_488,In_388);
nor U20 (N_20,In_136,In_181);
nand U21 (N_21,In_313,In_195);
or U22 (N_22,In_305,In_81);
nand U23 (N_23,In_60,In_422);
and U24 (N_24,In_364,In_177);
nor U25 (N_25,In_377,In_375);
nand U26 (N_26,In_444,In_191);
or U27 (N_27,In_134,In_5);
nand U28 (N_28,In_440,In_34);
nor U29 (N_29,In_211,In_210);
nand U30 (N_30,In_443,In_289);
and U31 (N_31,In_253,In_233);
and U32 (N_32,In_303,In_329);
and U33 (N_33,In_132,In_87);
and U34 (N_34,In_137,In_408);
or U35 (N_35,In_380,In_112);
and U36 (N_36,In_13,In_467);
and U37 (N_37,In_456,In_27);
and U38 (N_38,In_341,In_105);
nor U39 (N_39,In_261,In_38);
or U40 (N_40,In_486,In_337);
and U41 (N_41,In_325,In_176);
nand U42 (N_42,In_266,In_32);
and U43 (N_43,In_241,In_320);
and U44 (N_44,In_56,In_386);
nor U45 (N_45,In_118,In_356);
nor U46 (N_46,In_62,In_291);
and U47 (N_47,In_483,In_161);
or U48 (N_48,In_248,In_205);
or U49 (N_49,In_209,In_415);
and U50 (N_50,In_164,In_90);
nor U51 (N_51,In_316,In_295);
and U52 (N_52,In_0,In_61);
and U53 (N_53,In_376,In_399);
or U54 (N_54,In_113,In_296);
or U55 (N_55,In_128,In_59);
or U56 (N_56,In_499,In_319);
or U57 (N_57,In_333,In_401);
nor U58 (N_58,In_99,In_91);
nor U59 (N_59,In_436,In_416);
xor U60 (N_60,In_263,In_351);
nand U61 (N_61,In_414,In_411);
or U62 (N_62,In_63,In_133);
nor U63 (N_63,In_44,In_469);
nand U64 (N_64,In_300,In_265);
nand U65 (N_65,In_72,In_439);
nand U66 (N_66,In_17,In_317);
or U67 (N_67,In_79,In_204);
or U68 (N_68,In_203,In_77);
nor U69 (N_69,In_64,In_400);
or U70 (N_70,In_489,In_160);
nand U71 (N_71,In_173,In_276);
nor U72 (N_72,In_35,In_143);
and U73 (N_73,In_497,In_487);
nand U74 (N_74,In_428,In_171);
and U75 (N_75,In_334,In_144);
or U76 (N_76,In_158,In_452);
and U77 (N_77,In_168,In_448);
nor U78 (N_78,In_145,In_104);
and U79 (N_79,In_18,In_239);
nand U80 (N_80,In_121,In_30);
or U81 (N_81,In_55,In_286);
xor U82 (N_82,In_397,In_338);
or U83 (N_83,In_16,In_366);
nand U84 (N_84,In_242,In_374);
nand U85 (N_85,In_151,In_373);
or U86 (N_86,In_222,In_421);
nor U87 (N_87,In_78,In_354);
or U88 (N_88,In_407,In_106);
nand U89 (N_89,In_259,In_28);
xnor U90 (N_90,In_229,In_119);
or U91 (N_91,In_218,In_221);
nand U92 (N_92,In_466,In_350);
nor U93 (N_93,In_352,In_326);
and U94 (N_94,In_116,In_93);
nor U95 (N_95,In_82,In_175);
xnor U96 (N_96,In_315,In_437);
or U97 (N_97,In_148,In_19);
and U98 (N_98,In_199,In_277);
and U99 (N_99,In_123,In_293);
nor U100 (N_100,In_264,In_92);
or U101 (N_101,In_447,In_43);
nor U102 (N_102,In_464,In_189);
and U103 (N_103,In_200,In_463);
and U104 (N_104,In_257,In_361);
nor U105 (N_105,In_53,In_365);
nand U106 (N_106,In_141,In_348);
nor U107 (N_107,In_470,In_67);
nor U108 (N_108,In_445,In_73);
or U109 (N_109,In_153,In_122);
and U110 (N_110,In_288,In_282);
and U111 (N_111,In_258,In_39);
or U112 (N_112,In_196,In_394);
nand U113 (N_113,In_260,In_403);
and U114 (N_114,In_159,In_379);
nor U115 (N_115,In_202,In_327);
nor U116 (N_116,In_187,In_308);
nor U117 (N_117,In_432,In_100);
and U118 (N_118,In_324,In_51);
or U119 (N_119,In_1,In_438);
and U120 (N_120,In_298,In_231);
nor U121 (N_121,In_474,In_66);
and U122 (N_122,In_271,In_115);
nor U123 (N_123,In_26,In_485);
nand U124 (N_124,In_70,In_412);
nor U125 (N_125,In_235,In_435);
or U126 (N_126,In_462,In_36);
or U127 (N_127,In_232,In_311);
or U128 (N_128,In_249,In_150);
or U129 (N_129,In_75,In_353);
or U130 (N_130,In_262,In_157);
or U131 (N_131,In_299,In_498);
nand U132 (N_132,In_102,In_212);
nand U133 (N_133,In_423,In_419);
nor U134 (N_134,In_152,In_120);
and U135 (N_135,In_155,In_111);
and U136 (N_136,In_230,In_285);
nor U137 (N_137,In_331,In_29);
and U138 (N_138,In_83,In_193);
and U139 (N_139,In_243,In_455);
nor U140 (N_140,In_109,In_101);
nor U141 (N_141,In_124,In_108);
nand U142 (N_142,In_367,In_427);
nor U143 (N_143,In_347,In_336);
and U144 (N_144,In_339,In_281);
nand U145 (N_145,In_89,In_278);
nand U146 (N_146,In_172,In_254);
and U147 (N_147,In_344,In_98);
nor U148 (N_148,In_360,In_154);
or U149 (N_149,In_135,In_208);
nand U150 (N_150,In_174,In_96);
nor U151 (N_151,In_9,In_476);
and U152 (N_152,In_228,In_46);
nand U153 (N_153,In_216,In_410);
nand U154 (N_154,In_383,In_302);
nand U155 (N_155,In_398,In_314);
nand U156 (N_156,In_323,In_479);
and U157 (N_157,In_409,In_446);
nor U158 (N_158,In_76,In_318);
nor U159 (N_159,In_25,In_215);
or U160 (N_160,In_49,In_426);
or U161 (N_161,In_94,In_224);
or U162 (N_162,In_2,In_275);
and U163 (N_163,In_393,In_406);
nor U164 (N_164,In_8,In_280);
nor U165 (N_165,In_41,In_273);
nor U166 (N_166,In_246,In_45);
nor U167 (N_167,In_206,In_481);
nor U168 (N_168,In_392,In_475);
or U169 (N_169,In_10,In_292);
and U170 (N_170,In_378,In_142);
nand U171 (N_171,In_110,In_396);
or U172 (N_172,In_363,In_54);
nor U173 (N_173,In_420,In_166);
nand U174 (N_174,In_330,In_107);
and U175 (N_175,In_147,In_129);
or U176 (N_176,In_178,In_425);
nand U177 (N_177,In_310,In_194);
or U178 (N_178,In_368,In_207);
nand U179 (N_179,In_95,In_461);
and U180 (N_180,In_183,In_179);
and U181 (N_181,In_7,In_391);
nand U182 (N_182,In_149,In_381);
nand U183 (N_183,In_14,In_450);
and U184 (N_184,In_477,In_328);
nor U185 (N_185,In_395,In_74);
and U186 (N_186,In_244,In_355);
nor U187 (N_187,In_270,In_294);
and U188 (N_188,In_442,In_413);
or U189 (N_189,In_284,In_50);
nor U190 (N_190,In_287,In_389);
or U191 (N_191,In_493,In_201);
and U192 (N_192,In_371,In_131);
nand U193 (N_193,In_217,In_86);
nor U194 (N_194,In_214,In_80);
nand U195 (N_195,In_362,In_346);
and U196 (N_196,In_192,In_496);
and U197 (N_197,In_424,In_332);
or U198 (N_198,In_441,In_12);
or U199 (N_199,In_84,In_491);
or U200 (N_200,N_114,N_82);
nor U201 (N_201,N_182,N_0);
nand U202 (N_202,N_27,In_321);
nor U203 (N_203,N_190,N_163);
or U204 (N_204,N_79,N_140);
or U205 (N_205,N_96,N_172);
and U206 (N_206,N_127,In_240);
nor U207 (N_207,N_72,N_105);
or U208 (N_208,In_57,N_141);
and U209 (N_209,In_342,N_138);
and U210 (N_210,In_69,N_76);
nand U211 (N_211,In_85,In_471);
nand U212 (N_212,N_40,N_158);
and U213 (N_213,In_301,N_18);
nor U214 (N_214,N_122,In_20);
nor U215 (N_215,N_25,N_148);
nand U216 (N_216,In_114,N_34);
and U217 (N_217,N_58,N_30);
or U218 (N_218,N_102,In_472);
and U219 (N_219,N_171,N_74);
or U220 (N_220,N_28,N_100);
nor U221 (N_221,In_473,N_130);
nor U222 (N_222,N_156,N_170);
nor U223 (N_223,N_198,N_63);
nor U224 (N_224,N_62,N_87);
nor U225 (N_225,N_35,N_136);
nor U226 (N_226,N_19,In_478);
nand U227 (N_227,N_174,N_64);
nor U228 (N_228,N_161,N_121);
and U229 (N_229,N_70,In_167);
or U230 (N_230,In_198,In_307);
nand U231 (N_231,N_36,N_15);
nor U232 (N_232,N_152,In_484);
or U233 (N_233,In_227,In_417);
and U234 (N_234,In_434,In_22);
nor U235 (N_235,N_92,N_51);
or U236 (N_236,N_123,N_7);
nor U237 (N_237,N_57,In_459);
and U238 (N_238,N_53,N_146);
or U239 (N_239,In_359,In_88);
or U240 (N_240,N_160,N_12);
nand U241 (N_241,N_81,In_290);
and U242 (N_242,N_93,In_180);
nand U243 (N_243,N_192,N_185);
and U244 (N_244,In_65,In_6);
nand U245 (N_245,N_133,In_418);
and U246 (N_246,N_38,N_147);
nand U247 (N_247,N_150,N_67);
and U248 (N_248,In_335,N_103);
or U249 (N_249,N_115,N_31);
nand U250 (N_250,N_16,N_24);
nand U251 (N_251,In_238,In_297);
nor U252 (N_252,N_86,In_322);
nor U253 (N_253,N_120,N_107);
and U254 (N_254,In_495,In_169);
nor U255 (N_255,N_144,In_103);
nand U256 (N_256,N_61,In_268);
nand U257 (N_257,N_189,N_110);
nor U258 (N_258,N_112,N_71);
nand U259 (N_259,In_304,N_142);
or U260 (N_260,N_99,N_149);
and U261 (N_261,In_197,In_465);
and U262 (N_262,N_173,In_138);
and U263 (N_263,N_33,In_225);
and U264 (N_264,N_54,In_384);
and U265 (N_265,N_193,In_219);
nand U266 (N_266,In_256,N_199);
or U267 (N_267,In_385,N_42);
or U268 (N_268,N_143,N_108);
nor U269 (N_269,N_68,In_15);
and U270 (N_270,In_370,N_84);
nor U271 (N_271,In_21,In_454);
and U272 (N_272,N_89,N_128);
nor U273 (N_273,N_66,N_29);
nand U274 (N_274,N_157,N_41);
and U275 (N_275,In_48,N_47);
nand U276 (N_276,N_134,N_164);
or U277 (N_277,In_126,In_236);
and U278 (N_278,In_139,In_58);
nand U279 (N_279,N_162,N_118);
nand U280 (N_280,N_20,N_90);
nand U281 (N_281,N_52,N_117);
nand U282 (N_282,In_283,In_226);
or U283 (N_283,In_182,N_124);
nor U284 (N_284,N_83,N_111);
nand U285 (N_285,In_252,N_91);
and U286 (N_286,In_345,In_97);
or U287 (N_287,In_312,N_94);
nand U288 (N_288,In_382,In_237);
nor U289 (N_289,In_251,N_197);
nor U290 (N_290,N_26,N_153);
and U291 (N_291,N_126,N_80);
or U292 (N_292,In_457,In_156);
and U293 (N_293,In_451,N_177);
nand U294 (N_294,N_50,In_358);
nor U295 (N_295,In_433,N_46);
or U296 (N_296,In_490,N_8);
nor U297 (N_297,N_44,N_10);
or U298 (N_298,N_159,In_349);
or U299 (N_299,N_59,In_492);
and U300 (N_300,N_180,In_372);
or U301 (N_301,N_151,N_166);
nor U302 (N_302,N_49,In_71);
nor U303 (N_303,N_78,N_85);
and U304 (N_304,N_154,N_179);
and U305 (N_305,N_181,N_125);
or U306 (N_306,N_104,N_145);
nor U307 (N_307,N_169,N_113);
and U308 (N_308,N_95,N_56);
or U309 (N_309,In_234,N_119);
or U310 (N_310,N_186,N_4);
nand U311 (N_311,N_69,N_5);
or U312 (N_312,N_183,In_11);
nand U313 (N_313,N_88,In_250);
nand U314 (N_314,N_109,N_101);
nor U315 (N_315,N_195,N_116);
nor U316 (N_316,In_68,N_9);
or U317 (N_317,N_187,N_98);
or U318 (N_318,In_52,In_163);
or U319 (N_319,N_22,In_460);
nor U320 (N_320,In_42,In_170);
and U321 (N_321,N_97,N_178);
nand U322 (N_322,N_106,N_132);
nand U323 (N_323,N_137,N_21);
and U324 (N_324,N_194,In_255);
nand U325 (N_325,In_343,N_191);
and U326 (N_326,In_31,N_165);
and U327 (N_327,N_155,In_140);
and U328 (N_328,N_23,N_167);
or U329 (N_329,In_220,N_39);
or U330 (N_330,N_32,N_3);
nand U331 (N_331,In_47,N_77);
or U332 (N_332,N_135,N_176);
or U333 (N_333,N_139,In_24);
nand U334 (N_334,N_43,N_60);
nand U335 (N_335,N_168,N_188);
nor U336 (N_336,N_131,In_223);
or U337 (N_337,N_175,N_73);
nand U338 (N_338,N_37,In_185);
or U339 (N_339,N_196,N_14);
nor U340 (N_340,In_390,N_184);
nor U341 (N_341,In_279,In_405);
or U342 (N_342,N_11,N_75);
nand U343 (N_343,N_2,N_17);
nor U344 (N_344,N_6,N_48);
nand U345 (N_345,N_129,In_369);
or U346 (N_346,N_65,In_468);
nand U347 (N_347,N_45,In_125);
nor U348 (N_348,N_1,N_13);
nor U349 (N_349,N_55,In_431);
nand U350 (N_350,In_418,In_68);
or U351 (N_351,N_98,N_194);
or U352 (N_352,In_21,N_7);
nor U353 (N_353,N_116,In_22);
or U354 (N_354,N_199,N_158);
and U355 (N_355,N_80,N_21);
or U356 (N_356,In_225,In_237);
or U357 (N_357,N_156,N_172);
nor U358 (N_358,N_158,N_91);
nor U359 (N_359,N_3,N_165);
nor U360 (N_360,N_43,N_145);
or U361 (N_361,N_168,In_225);
and U362 (N_362,N_60,N_100);
nand U363 (N_363,In_22,N_16);
and U364 (N_364,N_199,In_227);
or U365 (N_365,N_185,N_4);
nand U366 (N_366,In_335,In_182);
or U367 (N_367,N_125,N_196);
nor U368 (N_368,N_124,In_219);
and U369 (N_369,N_154,N_10);
nand U370 (N_370,In_322,N_45);
and U371 (N_371,N_76,N_177);
and U372 (N_372,N_5,N_81);
nand U373 (N_373,N_24,In_478);
nand U374 (N_374,In_335,In_484);
nor U375 (N_375,In_492,N_80);
nor U376 (N_376,In_473,N_166);
or U377 (N_377,N_13,In_138);
nor U378 (N_378,N_171,In_390);
nand U379 (N_379,N_6,N_144);
and U380 (N_380,N_115,N_37);
and U381 (N_381,N_140,N_12);
and U382 (N_382,In_234,In_126);
nor U383 (N_383,In_451,N_162);
and U384 (N_384,In_372,N_126);
nor U385 (N_385,In_88,N_44);
and U386 (N_386,N_36,N_158);
and U387 (N_387,N_159,In_22);
and U388 (N_388,In_434,In_322);
nor U389 (N_389,N_134,N_16);
and U390 (N_390,N_191,In_301);
and U391 (N_391,N_198,N_188);
or U392 (N_392,N_110,In_457);
and U393 (N_393,N_25,N_32);
nand U394 (N_394,In_223,In_343);
and U395 (N_395,N_15,N_143);
and U396 (N_396,N_148,N_1);
nor U397 (N_397,In_57,N_74);
nand U398 (N_398,In_103,N_165);
nand U399 (N_399,In_220,N_45);
and U400 (N_400,N_354,N_261);
nand U401 (N_401,N_392,N_312);
or U402 (N_402,N_340,N_317);
nor U403 (N_403,N_241,N_376);
and U404 (N_404,N_362,N_379);
and U405 (N_405,N_239,N_283);
nand U406 (N_406,N_243,N_217);
or U407 (N_407,N_389,N_366);
or U408 (N_408,N_298,N_396);
nor U409 (N_409,N_204,N_201);
nor U410 (N_410,N_287,N_351);
or U411 (N_411,N_321,N_349);
nor U412 (N_412,N_288,N_314);
xnor U413 (N_413,N_277,N_368);
and U414 (N_414,N_297,N_350);
nor U415 (N_415,N_306,N_384);
or U416 (N_416,N_330,N_395);
nand U417 (N_417,N_352,N_335);
nand U418 (N_418,N_381,N_248);
and U419 (N_419,N_347,N_226);
or U420 (N_420,N_294,N_268);
and U421 (N_421,N_371,N_210);
nor U422 (N_422,N_383,N_219);
and U423 (N_423,N_291,N_266);
or U424 (N_424,N_229,N_355);
or U425 (N_425,N_380,N_397);
nand U426 (N_426,N_394,N_387);
nand U427 (N_427,N_228,N_273);
or U428 (N_428,N_256,N_225);
or U429 (N_429,N_233,N_245);
or U430 (N_430,N_393,N_215);
nor U431 (N_431,N_275,N_367);
nor U432 (N_432,N_203,N_338);
or U433 (N_433,N_222,N_202);
and U434 (N_434,N_258,N_382);
nor U435 (N_435,N_333,N_348);
nor U436 (N_436,N_274,N_254);
nand U437 (N_437,N_308,N_237);
nor U438 (N_438,N_208,N_206);
nor U439 (N_439,N_255,N_227);
and U440 (N_440,N_220,N_358);
nor U441 (N_441,N_279,N_249);
nand U442 (N_442,N_316,N_374);
or U443 (N_443,N_301,N_238);
or U444 (N_444,N_205,N_234);
nand U445 (N_445,N_260,N_286);
nand U446 (N_446,N_398,N_271);
nor U447 (N_447,N_325,N_339);
nor U448 (N_448,N_334,N_327);
nor U449 (N_449,N_280,N_307);
or U450 (N_450,N_251,N_257);
or U451 (N_451,N_328,N_244);
or U452 (N_452,N_372,N_343);
and U453 (N_453,N_259,N_337);
nand U454 (N_454,N_363,N_231);
nand U455 (N_455,N_270,N_386);
nor U456 (N_456,N_216,N_311);
nand U457 (N_457,N_322,N_281);
or U458 (N_458,N_224,N_329);
nand U459 (N_459,N_253,N_299);
or U460 (N_460,N_292,N_353);
or U461 (N_461,N_212,N_315);
nand U462 (N_462,N_214,N_385);
nor U463 (N_463,N_323,N_356);
and U464 (N_464,N_341,N_344);
or U465 (N_465,N_310,N_319);
nand U466 (N_466,N_296,N_326);
or U467 (N_467,N_346,N_272);
nor U468 (N_468,N_282,N_242);
and U469 (N_469,N_264,N_345);
nand U470 (N_470,N_309,N_300);
nor U471 (N_471,N_269,N_276);
nor U472 (N_472,N_364,N_377);
nand U473 (N_473,N_207,N_378);
and U474 (N_474,N_365,N_289);
or U475 (N_475,N_324,N_359);
and U476 (N_476,N_318,N_373);
and U477 (N_477,N_252,N_246);
nor U478 (N_478,N_235,N_360);
nand U479 (N_479,N_313,N_361);
or U480 (N_480,N_290,N_211);
nor U481 (N_481,N_375,N_200);
nor U482 (N_482,N_305,N_342);
nand U483 (N_483,N_278,N_230);
or U484 (N_484,N_370,N_262);
nand U485 (N_485,N_357,N_331);
or U486 (N_486,N_263,N_369);
nor U487 (N_487,N_223,N_232);
nor U488 (N_488,N_320,N_303);
nor U489 (N_489,N_236,N_285);
or U490 (N_490,N_221,N_388);
nor U491 (N_491,N_399,N_332);
nand U492 (N_492,N_293,N_218);
and U493 (N_493,N_390,N_304);
and U494 (N_494,N_267,N_265);
or U495 (N_495,N_284,N_209);
nand U496 (N_496,N_336,N_302);
nand U497 (N_497,N_295,N_250);
nor U498 (N_498,N_247,N_213);
nor U499 (N_499,N_391,N_240);
nor U500 (N_500,N_358,N_233);
or U501 (N_501,N_365,N_268);
or U502 (N_502,N_345,N_386);
or U503 (N_503,N_395,N_224);
and U504 (N_504,N_256,N_383);
nand U505 (N_505,N_385,N_210);
and U506 (N_506,N_221,N_365);
nand U507 (N_507,N_363,N_324);
nand U508 (N_508,N_239,N_276);
or U509 (N_509,N_361,N_201);
nor U510 (N_510,N_206,N_353);
and U511 (N_511,N_215,N_326);
nor U512 (N_512,N_223,N_247);
or U513 (N_513,N_388,N_206);
nand U514 (N_514,N_378,N_310);
nor U515 (N_515,N_221,N_355);
or U516 (N_516,N_287,N_355);
and U517 (N_517,N_260,N_358);
and U518 (N_518,N_215,N_253);
nand U519 (N_519,N_335,N_342);
or U520 (N_520,N_340,N_378);
nand U521 (N_521,N_288,N_225);
or U522 (N_522,N_243,N_360);
nor U523 (N_523,N_206,N_216);
or U524 (N_524,N_337,N_308);
nand U525 (N_525,N_352,N_319);
or U526 (N_526,N_284,N_307);
and U527 (N_527,N_390,N_225);
or U528 (N_528,N_330,N_398);
and U529 (N_529,N_381,N_359);
and U530 (N_530,N_319,N_234);
and U531 (N_531,N_341,N_380);
and U532 (N_532,N_278,N_263);
nand U533 (N_533,N_283,N_278);
and U534 (N_534,N_215,N_360);
or U535 (N_535,N_207,N_297);
nor U536 (N_536,N_257,N_265);
or U537 (N_537,N_362,N_279);
nor U538 (N_538,N_325,N_283);
or U539 (N_539,N_318,N_288);
nand U540 (N_540,N_365,N_258);
and U541 (N_541,N_217,N_384);
or U542 (N_542,N_305,N_313);
nand U543 (N_543,N_266,N_394);
nand U544 (N_544,N_253,N_324);
nor U545 (N_545,N_379,N_230);
and U546 (N_546,N_262,N_380);
nor U547 (N_547,N_233,N_266);
nand U548 (N_548,N_290,N_233);
nand U549 (N_549,N_305,N_238);
nand U550 (N_550,N_354,N_376);
and U551 (N_551,N_254,N_374);
nand U552 (N_552,N_319,N_357);
nand U553 (N_553,N_260,N_294);
or U554 (N_554,N_201,N_329);
or U555 (N_555,N_370,N_251);
nand U556 (N_556,N_338,N_363);
nand U557 (N_557,N_332,N_263);
xnor U558 (N_558,N_317,N_344);
nand U559 (N_559,N_359,N_269);
and U560 (N_560,N_315,N_259);
or U561 (N_561,N_387,N_324);
or U562 (N_562,N_293,N_349);
nor U563 (N_563,N_308,N_239);
nand U564 (N_564,N_312,N_357);
nand U565 (N_565,N_210,N_292);
or U566 (N_566,N_265,N_307);
nand U567 (N_567,N_327,N_388);
and U568 (N_568,N_244,N_214);
and U569 (N_569,N_258,N_268);
and U570 (N_570,N_307,N_305);
nor U571 (N_571,N_320,N_307);
and U572 (N_572,N_266,N_389);
nand U573 (N_573,N_358,N_362);
nand U574 (N_574,N_278,N_398);
nor U575 (N_575,N_279,N_248);
nand U576 (N_576,N_364,N_209);
nand U577 (N_577,N_319,N_251);
or U578 (N_578,N_213,N_235);
or U579 (N_579,N_281,N_328);
or U580 (N_580,N_320,N_272);
nor U581 (N_581,N_287,N_247);
nand U582 (N_582,N_266,N_293);
or U583 (N_583,N_231,N_339);
nand U584 (N_584,N_289,N_336);
nor U585 (N_585,N_235,N_273);
nor U586 (N_586,N_337,N_231);
and U587 (N_587,N_388,N_376);
nor U588 (N_588,N_331,N_347);
and U589 (N_589,N_303,N_322);
or U590 (N_590,N_361,N_303);
nand U591 (N_591,N_312,N_280);
nor U592 (N_592,N_250,N_327);
and U593 (N_593,N_379,N_200);
nand U594 (N_594,N_228,N_246);
nand U595 (N_595,N_382,N_299);
and U596 (N_596,N_212,N_273);
or U597 (N_597,N_275,N_203);
nand U598 (N_598,N_236,N_390);
nand U599 (N_599,N_389,N_392);
nand U600 (N_600,N_595,N_587);
and U601 (N_601,N_426,N_440);
nor U602 (N_602,N_554,N_438);
and U603 (N_603,N_461,N_588);
nand U604 (N_604,N_533,N_403);
or U605 (N_605,N_464,N_580);
or U606 (N_606,N_418,N_512);
and U607 (N_607,N_527,N_474);
and U608 (N_608,N_547,N_549);
or U609 (N_609,N_433,N_445);
nand U610 (N_610,N_525,N_489);
and U611 (N_611,N_422,N_538);
or U612 (N_612,N_496,N_468);
nor U613 (N_613,N_408,N_480);
or U614 (N_614,N_524,N_495);
or U615 (N_615,N_473,N_485);
and U616 (N_616,N_592,N_486);
or U617 (N_617,N_471,N_419);
nor U618 (N_618,N_570,N_405);
nor U619 (N_619,N_511,N_487);
nor U620 (N_620,N_400,N_558);
or U621 (N_621,N_566,N_425);
or U622 (N_622,N_413,N_574);
nand U623 (N_623,N_492,N_494);
and U624 (N_624,N_517,N_559);
and U625 (N_625,N_594,N_424);
or U626 (N_626,N_569,N_583);
or U627 (N_627,N_539,N_585);
nand U628 (N_628,N_515,N_548);
nand U629 (N_629,N_540,N_450);
nand U630 (N_630,N_555,N_545);
and U631 (N_631,N_514,N_455);
and U632 (N_632,N_441,N_541);
nor U633 (N_633,N_502,N_597);
nand U634 (N_634,N_535,N_534);
nor U635 (N_635,N_478,N_449);
or U636 (N_636,N_465,N_409);
and U637 (N_637,N_453,N_467);
or U638 (N_638,N_551,N_475);
and U639 (N_639,N_443,N_488);
nor U640 (N_640,N_499,N_469);
nand U641 (N_641,N_546,N_463);
or U642 (N_642,N_452,N_421);
nor U643 (N_643,N_528,N_578);
or U644 (N_644,N_522,N_513);
or U645 (N_645,N_564,N_508);
nor U646 (N_646,N_526,N_412);
and U647 (N_647,N_589,N_544);
nor U648 (N_648,N_430,N_503);
nand U649 (N_649,N_586,N_573);
nand U650 (N_650,N_420,N_504);
and U651 (N_651,N_531,N_431);
and U652 (N_652,N_576,N_428);
nand U653 (N_653,N_556,N_596);
nand U654 (N_654,N_568,N_567);
and U655 (N_655,N_537,N_429);
nor U656 (N_656,N_542,N_577);
or U657 (N_657,N_582,N_435);
and U658 (N_658,N_500,N_584);
or U659 (N_659,N_560,N_451);
and U660 (N_660,N_493,N_519);
or U661 (N_661,N_507,N_529);
nand U662 (N_662,N_593,N_470);
nand U663 (N_663,N_575,N_476);
or U664 (N_664,N_510,N_509);
and U665 (N_665,N_446,N_423);
or U666 (N_666,N_447,N_466);
nor U667 (N_667,N_472,N_553);
or U668 (N_668,N_557,N_457);
and U669 (N_669,N_483,N_523);
nand U670 (N_670,N_484,N_490);
or U671 (N_671,N_414,N_590);
nor U672 (N_672,N_477,N_456);
or U673 (N_673,N_598,N_562);
nand U674 (N_674,N_444,N_550);
or U675 (N_675,N_454,N_459);
or U676 (N_676,N_439,N_520);
or U677 (N_677,N_427,N_572);
and U678 (N_678,N_571,N_481);
and U679 (N_679,N_565,N_406);
or U680 (N_680,N_591,N_462);
and U681 (N_681,N_536,N_432);
and U682 (N_682,N_402,N_482);
nand U683 (N_683,N_479,N_552);
nor U684 (N_684,N_407,N_505);
or U685 (N_685,N_543,N_448);
nor U686 (N_686,N_491,N_410);
and U687 (N_687,N_521,N_501);
and U688 (N_688,N_434,N_506);
nand U689 (N_689,N_460,N_404);
nand U690 (N_690,N_401,N_561);
and U691 (N_691,N_579,N_498);
and U692 (N_692,N_581,N_516);
and U693 (N_693,N_415,N_436);
nor U694 (N_694,N_497,N_518);
nor U695 (N_695,N_416,N_530);
or U696 (N_696,N_599,N_437);
and U697 (N_697,N_532,N_417);
nand U698 (N_698,N_411,N_563);
nand U699 (N_699,N_442,N_458);
nand U700 (N_700,N_470,N_468);
or U701 (N_701,N_458,N_496);
or U702 (N_702,N_584,N_444);
nor U703 (N_703,N_484,N_472);
nor U704 (N_704,N_422,N_436);
nand U705 (N_705,N_513,N_414);
and U706 (N_706,N_416,N_506);
or U707 (N_707,N_424,N_484);
nand U708 (N_708,N_496,N_508);
nor U709 (N_709,N_477,N_561);
and U710 (N_710,N_475,N_453);
nor U711 (N_711,N_419,N_574);
nand U712 (N_712,N_484,N_563);
nand U713 (N_713,N_487,N_406);
or U714 (N_714,N_427,N_589);
or U715 (N_715,N_552,N_543);
xnor U716 (N_716,N_453,N_473);
and U717 (N_717,N_582,N_440);
nor U718 (N_718,N_574,N_464);
and U719 (N_719,N_460,N_546);
nor U720 (N_720,N_547,N_427);
nor U721 (N_721,N_449,N_433);
and U722 (N_722,N_469,N_439);
nand U723 (N_723,N_535,N_443);
nand U724 (N_724,N_407,N_499);
nor U725 (N_725,N_476,N_418);
or U726 (N_726,N_504,N_425);
nor U727 (N_727,N_540,N_484);
nor U728 (N_728,N_451,N_599);
nor U729 (N_729,N_467,N_552);
nand U730 (N_730,N_596,N_549);
nor U731 (N_731,N_583,N_571);
nand U732 (N_732,N_598,N_469);
and U733 (N_733,N_418,N_452);
nor U734 (N_734,N_529,N_438);
and U735 (N_735,N_533,N_413);
nor U736 (N_736,N_439,N_456);
or U737 (N_737,N_429,N_487);
xor U738 (N_738,N_581,N_597);
and U739 (N_739,N_442,N_499);
or U740 (N_740,N_435,N_474);
nor U741 (N_741,N_500,N_484);
or U742 (N_742,N_448,N_531);
nor U743 (N_743,N_568,N_548);
nor U744 (N_744,N_524,N_563);
nor U745 (N_745,N_443,N_415);
and U746 (N_746,N_416,N_594);
nand U747 (N_747,N_500,N_589);
or U748 (N_748,N_458,N_472);
nand U749 (N_749,N_550,N_508);
nand U750 (N_750,N_451,N_555);
and U751 (N_751,N_453,N_492);
or U752 (N_752,N_446,N_565);
nand U753 (N_753,N_502,N_551);
nor U754 (N_754,N_567,N_478);
nand U755 (N_755,N_500,N_474);
nor U756 (N_756,N_491,N_457);
and U757 (N_757,N_523,N_537);
and U758 (N_758,N_536,N_443);
nor U759 (N_759,N_417,N_508);
nand U760 (N_760,N_598,N_410);
and U761 (N_761,N_480,N_487);
nor U762 (N_762,N_472,N_591);
and U763 (N_763,N_579,N_418);
and U764 (N_764,N_584,N_413);
nand U765 (N_765,N_449,N_553);
or U766 (N_766,N_512,N_415);
nand U767 (N_767,N_443,N_438);
and U768 (N_768,N_515,N_445);
and U769 (N_769,N_542,N_496);
and U770 (N_770,N_435,N_421);
nand U771 (N_771,N_517,N_501);
nor U772 (N_772,N_534,N_569);
nor U773 (N_773,N_599,N_473);
or U774 (N_774,N_548,N_428);
and U775 (N_775,N_558,N_591);
nor U776 (N_776,N_515,N_437);
nand U777 (N_777,N_428,N_443);
nor U778 (N_778,N_417,N_543);
and U779 (N_779,N_424,N_431);
nand U780 (N_780,N_498,N_559);
nand U781 (N_781,N_485,N_466);
nand U782 (N_782,N_422,N_516);
nand U783 (N_783,N_416,N_575);
or U784 (N_784,N_503,N_448);
nand U785 (N_785,N_516,N_523);
and U786 (N_786,N_533,N_534);
nor U787 (N_787,N_500,N_519);
or U788 (N_788,N_586,N_439);
nand U789 (N_789,N_419,N_535);
or U790 (N_790,N_442,N_429);
nand U791 (N_791,N_575,N_466);
nor U792 (N_792,N_411,N_495);
nor U793 (N_793,N_598,N_590);
and U794 (N_794,N_501,N_575);
or U795 (N_795,N_460,N_532);
nand U796 (N_796,N_578,N_588);
nand U797 (N_797,N_410,N_432);
nor U798 (N_798,N_509,N_430);
nor U799 (N_799,N_450,N_582);
nor U800 (N_800,N_600,N_708);
or U801 (N_801,N_639,N_724);
or U802 (N_802,N_674,N_725);
nor U803 (N_803,N_676,N_787);
nor U804 (N_804,N_665,N_617);
nor U805 (N_805,N_785,N_700);
nor U806 (N_806,N_680,N_623);
and U807 (N_807,N_721,N_633);
nor U808 (N_808,N_796,N_627);
nand U809 (N_809,N_630,N_686);
nor U810 (N_810,N_652,N_682);
nor U811 (N_811,N_656,N_745);
nand U812 (N_812,N_766,N_770);
and U813 (N_813,N_655,N_612);
or U814 (N_814,N_769,N_677);
or U815 (N_815,N_668,N_752);
nor U816 (N_816,N_698,N_768);
or U817 (N_817,N_691,N_651);
and U818 (N_818,N_797,N_703);
nor U819 (N_819,N_730,N_722);
nand U820 (N_820,N_783,N_748);
nor U821 (N_821,N_688,N_736);
or U822 (N_822,N_731,N_789);
nor U823 (N_823,N_728,N_664);
nand U824 (N_824,N_739,N_660);
and U825 (N_825,N_695,N_793);
nand U826 (N_826,N_788,N_616);
or U827 (N_827,N_758,N_608);
nor U828 (N_828,N_798,N_646);
and U829 (N_829,N_777,N_625);
and U830 (N_830,N_718,N_693);
or U831 (N_831,N_707,N_753);
nand U832 (N_832,N_605,N_714);
or U833 (N_833,N_778,N_772);
or U834 (N_834,N_776,N_712);
nand U835 (N_835,N_618,N_624);
nor U836 (N_836,N_663,N_621);
and U837 (N_837,N_644,N_791);
or U838 (N_838,N_678,N_715);
or U839 (N_839,N_751,N_734);
or U840 (N_840,N_645,N_641);
or U841 (N_841,N_657,N_779);
or U842 (N_842,N_604,N_642);
nand U843 (N_843,N_611,N_799);
or U844 (N_844,N_732,N_620);
nand U845 (N_845,N_759,N_729);
nand U846 (N_846,N_781,N_749);
or U847 (N_847,N_774,N_726);
and U848 (N_848,N_670,N_701);
nand U849 (N_849,N_790,N_784);
or U850 (N_850,N_672,N_705);
nor U851 (N_851,N_634,N_635);
and U852 (N_852,N_761,N_754);
nand U853 (N_853,N_649,N_683);
nor U854 (N_854,N_738,N_632);
nand U855 (N_855,N_636,N_637);
and U856 (N_856,N_773,N_607);
and U857 (N_857,N_654,N_786);
nand U858 (N_858,N_610,N_606);
and U859 (N_859,N_720,N_692);
or U860 (N_860,N_792,N_702);
nor U861 (N_861,N_647,N_767);
nand U862 (N_862,N_628,N_603);
nand U863 (N_863,N_640,N_723);
or U864 (N_864,N_794,N_669);
and U865 (N_865,N_763,N_667);
and U866 (N_866,N_764,N_694);
nand U867 (N_867,N_711,N_775);
or U868 (N_868,N_706,N_744);
and U869 (N_869,N_709,N_648);
nor U870 (N_870,N_661,N_771);
or U871 (N_871,N_681,N_653);
nor U872 (N_872,N_643,N_622);
nand U873 (N_873,N_765,N_629);
nand U874 (N_874,N_684,N_743);
nand U875 (N_875,N_710,N_601);
or U876 (N_876,N_719,N_666);
or U877 (N_877,N_689,N_737);
nor U878 (N_878,N_740,N_658);
nand U879 (N_879,N_755,N_673);
and U880 (N_880,N_638,N_679);
or U881 (N_881,N_757,N_742);
and U882 (N_882,N_609,N_671);
nor U883 (N_883,N_690,N_615);
nand U884 (N_884,N_756,N_733);
nand U885 (N_885,N_613,N_696);
or U886 (N_886,N_735,N_762);
and U887 (N_887,N_631,N_675);
nand U888 (N_888,N_747,N_697);
or U889 (N_889,N_659,N_662);
or U890 (N_890,N_782,N_704);
nand U891 (N_891,N_746,N_626);
nand U892 (N_892,N_619,N_699);
and U893 (N_893,N_760,N_780);
or U894 (N_894,N_685,N_717);
nor U895 (N_895,N_741,N_687);
and U896 (N_896,N_650,N_713);
or U897 (N_897,N_716,N_602);
nor U898 (N_898,N_750,N_727);
and U899 (N_899,N_614,N_795);
and U900 (N_900,N_610,N_615);
nor U901 (N_901,N_608,N_732);
or U902 (N_902,N_758,N_621);
nand U903 (N_903,N_768,N_765);
and U904 (N_904,N_691,N_769);
nand U905 (N_905,N_670,N_627);
nor U906 (N_906,N_742,N_744);
nor U907 (N_907,N_606,N_796);
nand U908 (N_908,N_787,N_656);
and U909 (N_909,N_652,N_648);
and U910 (N_910,N_702,N_710);
or U911 (N_911,N_717,N_733);
or U912 (N_912,N_649,N_635);
xnor U913 (N_913,N_687,N_779);
or U914 (N_914,N_760,N_662);
or U915 (N_915,N_749,N_667);
and U916 (N_916,N_753,N_651);
or U917 (N_917,N_781,N_601);
and U918 (N_918,N_632,N_702);
or U919 (N_919,N_666,N_717);
and U920 (N_920,N_683,N_685);
and U921 (N_921,N_708,N_712);
or U922 (N_922,N_711,N_700);
and U923 (N_923,N_729,N_661);
and U924 (N_924,N_718,N_795);
or U925 (N_925,N_742,N_740);
nand U926 (N_926,N_787,N_689);
or U927 (N_927,N_670,N_631);
and U928 (N_928,N_690,N_731);
or U929 (N_929,N_687,N_773);
nand U930 (N_930,N_744,N_788);
nor U931 (N_931,N_779,N_682);
or U932 (N_932,N_676,N_733);
nand U933 (N_933,N_750,N_605);
and U934 (N_934,N_765,N_659);
and U935 (N_935,N_792,N_784);
nand U936 (N_936,N_768,N_774);
nand U937 (N_937,N_767,N_611);
nand U938 (N_938,N_738,N_619);
nor U939 (N_939,N_675,N_727);
or U940 (N_940,N_621,N_778);
or U941 (N_941,N_771,N_769);
nor U942 (N_942,N_630,N_792);
or U943 (N_943,N_617,N_627);
nor U944 (N_944,N_781,N_670);
or U945 (N_945,N_715,N_674);
and U946 (N_946,N_722,N_657);
and U947 (N_947,N_621,N_666);
nor U948 (N_948,N_722,N_680);
nor U949 (N_949,N_640,N_637);
and U950 (N_950,N_745,N_699);
or U951 (N_951,N_684,N_782);
or U952 (N_952,N_715,N_764);
or U953 (N_953,N_727,N_797);
and U954 (N_954,N_652,N_746);
nand U955 (N_955,N_611,N_760);
and U956 (N_956,N_755,N_628);
and U957 (N_957,N_685,N_734);
nor U958 (N_958,N_731,N_729);
nand U959 (N_959,N_659,N_683);
and U960 (N_960,N_676,N_604);
nor U961 (N_961,N_781,N_712);
nand U962 (N_962,N_768,N_661);
or U963 (N_963,N_788,N_650);
or U964 (N_964,N_789,N_683);
and U965 (N_965,N_759,N_746);
nand U966 (N_966,N_755,N_624);
nor U967 (N_967,N_772,N_672);
nand U968 (N_968,N_627,N_740);
nor U969 (N_969,N_658,N_619);
nand U970 (N_970,N_773,N_602);
or U971 (N_971,N_637,N_600);
and U972 (N_972,N_637,N_743);
or U973 (N_973,N_784,N_677);
nand U974 (N_974,N_733,N_791);
nor U975 (N_975,N_616,N_754);
nand U976 (N_976,N_767,N_762);
nor U977 (N_977,N_757,N_655);
nor U978 (N_978,N_773,N_666);
and U979 (N_979,N_744,N_661);
and U980 (N_980,N_760,N_661);
nand U981 (N_981,N_645,N_729);
and U982 (N_982,N_650,N_652);
xor U983 (N_983,N_756,N_662);
or U984 (N_984,N_772,N_676);
and U985 (N_985,N_755,N_700);
nand U986 (N_986,N_671,N_668);
nand U987 (N_987,N_719,N_655);
and U988 (N_988,N_751,N_728);
or U989 (N_989,N_771,N_699);
or U990 (N_990,N_758,N_740);
and U991 (N_991,N_768,N_684);
xnor U992 (N_992,N_665,N_754);
and U993 (N_993,N_752,N_623);
or U994 (N_994,N_769,N_614);
nor U995 (N_995,N_794,N_646);
nand U996 (N_996,N_680,N_679);
nor U997 (N_997,N_681,N_734);
nand U998 (N_998,N_798,N_661);
nand U999 (N_999,N_738,N_728);
nor U1000 (N_1000,N_812,N_945);
nand U1001 (N_1001,N_914,N_826);
or U1002 (N_1002,N_920,N_807);
and U1003 (N_1003,N_853,N_922);
nor U1004 (N_1004,N_904,N_973);
nor U1005 (N_1005,N_854,N_856);
nor U1006 (N_1006,N_907,N_846);
and U1007 (N_1007,N_992,N_848);
or U1008 (N_1008,N_836,N_892);
nor U1009 (N_1009,N_840,N_911);
and U1010 (N_1010,N_942,N_936);
nand U1011 (N_1011,N_841,N_921);
or U1012 (N_1012,N_970,N_981);
nand U1013 (N_1013,N_838,N_993);
and U1014 (N_1014,N_972,N_974);
or U1015 (N_1015,N_969,N_900);
or U1016 (N_1016,N_937,N_824);
nand U1017 (N_1017,N_961,N_873);
nand U1018 (N_1018,N_849,N_845);
nor U1019 (N_1019,N_834,N_822);
and U1020 (N_1020,N_967,N_863);
nand U1021 (N_1021,N_929,N_978);
and U1022 (N_1022,N_996,N_805);
and U1023 (N_1023,N_964,N_913);
and U1024 (N_1024,N_924,N_948);
or U1025 (N_1025,N_966,N_851);
nor U1026 (N_1026,N_938,N_896);
nor U1027 (N_1027,N_864,N_808);
nand U1028 (N_1028,N_815,N_935);
and U1029 (N_1029,N_891,N_949);
nand U1030 (N_1030,N_820,N_857);
and U1031 (N_1031,N_843,N_988);
and U1032 (N_1032,N_987,N_979);
nor U1033 (N_1033,N_901,N_902);
and U1034 (N_1034,N_852,N_888);
and U1035 (N_1035,N_931,N_917);
nand U1036 (N_1036,N_977,N_905);
nand U1037 (N_1037,N_816,N_821);
or U1038 (N_1038,N_871,N_819);
and U1039 (N_1039,N_866,N_958);
or U1040 (N_1040,N_882,N_919);
or U1041 (N_1041,N_889,N_875);
nor U1042 (N_1042,N_918,N_802);
nand U1043 (N_1043,N_941,N_886);
nor U1044 (N_1044,N_818,N_939);
and U1045 (N_1045,N_984,N_906);
nor U1046 (N_1046,N_809,N_810);
nand U1047 (N_1047,N_860,N_926);
nor U1048 (N_1048,N_950,N_874);
nand U1049 (N_1049,N_932,N_858);
nand U1050 (N_1050,N_833,N_835);
and U1051 (N_1051,N_957,N_825);
nand U1052 (N_1052,N_837,N_930);
or U1053 (N_1053,N_829,N_983);
nor U1054 (N_1054,N_803,N_868);
nor U1055 (N_1055,N_839,N_850);
or U1056 (N_1056,N_859,N_847);
nor U1057 (N_1057,N_903,N_940);
and U1058 (N_1058,N_883,N_842);
or U1059 (N_1059,N_817,N_963);
and U1060 (N_1060,N_879,N_946);
and U1061 (N_1061,N_965,N_885);
or U1062 (N_1062,N_971,N_823);
or U1063 (N_1063,N_916,N_912);
and U1064 (N_1064,N_999,N_985);
and U1065 (N_1065,N_954,N_890);
or U1066 (N_1066,N_934,N_830);
nand U1067 (N_1067,N_894,N_951);
and U1068 (N_1068,N_976,N_801);
nand U1069 (N_1069,N_980,N_908);
nand U1070 (N_1070,N_869,N_952);
and U1071 (N_1071,N_881,N_811);
nand U1072 (N_1072,N_944,N_925);
nor U1073 (N_1073,N_832,N_933);
nand U1074 (N_1074,N_870,N_813);
or U1075 (N_1075,N_800,N_806);
or U1076 (N_1076,N_880,N_887);
nor U1077 (N_1077,N_997,N_990);
nand U1078 (N_1078,N_982,N_991);
xor U1079 (N_1079,N_960,N_898);
and U1080 (N_1080,N_855,N_895);
or U1081 (N_1081,N_928,N_814);
nand U1082 (N_1082,N_877,N_959);
and U1083 (N_1083,N_923,N_956);
or U1084 (N_1084,N_998,N_947);
nand U1085 (N_1085,N_862,N_968);
and U1086 (N_1086,N_893,N_995);
nand U1087 (N_1087,N_804,N_989);
nor U1088 (N_1088,N_899,N_927);
nand U1089 (N_1089,N_962,N_915);
and U1090 (N_1090,N_876,N_953);
and U1091 (N_1091,N_867,N_943);
nand U1092 (N_1092,N_828,N_878);
nand U1093 (N_1093,N_910,N_986);
and U1094 (N_1094,N_844,N_955);
or U1095 (N_1095,N_884,N_831);
nor U1096 (N_1096,N_897,N_865);
nand U1097 (N_1097,N_827,N_861);
and U1098 (N_1098,N_872,N_909);
nand U1099 (N_1099,N_975,N_994);
or U1100 (N_1100,N_928,N_828);
nand U1101 (N_1101,N_966,N_985);
nor U1102 (N_1102,N_897,N_965);
nor U1103 (N_1103,N_827,N_868);
and U1104 (N_1104,N_948,N_986);
or U1105 (N_1105,N_889,N_976);
nand U1106 (N_1106,N_964,N_815);
nand U1107 (N_1107,N_927,N_895);
nor U1108 (N_1108,N_860,N_910);
and U1109 (N_1109,N_898,N_893);
nand U1110 (N_1110,N_896,N_976);
or U1111 (N_1111,N_938,N_875);
nor U1112 (N_1112,N_851,N_932);
nand U1113 (N_1113,N_924,N_828);
nand U1114 (N_1114,N_921,N_933);
or U1115 (N_1115,N_894,N_943);
and U1116 (N_1116,N_868,N_883);
nor U1117 (N_1117,N_947,N_844);
nor U1118 (N_1118,N_896,N_855);
and U1119 (N_1119,N_988,N_927);
or U1120 (N_1120,N_824,N_962);
or U1121 (N_1121,N_852,N_808);
nand U1122 (N_1122,N_831,N_932);
and U1123 (N_1123,N_848,N_816);
nand U1124 (N_1124,N_867,N_958);
nor U1125 (N_1125,N_998,N_892);
nor U1126 (N_1126,N_946,N_831);
and U1127 (N_1127,N_810,N_936);
and U1128 (N_1128,N_918,N_832);
nor U1129 (N_1129,N_878,N_886);
or U1130 (N_1130,N_959,N_816);
nor U1131 (N_1131,N_857,N_931);
or U1132 (N_1132,N_825,N_966);
and U1133 (N_1133,N_861,N_851);
nand U1134 (N_1134,N_934,N_840);
and U1135 (N_1135,N_894,N_938);
or U1136 (N_1136,N_930,N_886);
and U1137 (N_1137,N_889,N_885);
and U1138 (N_1138,N_850,N_831);
and U1139 (N_1139,N_809,N_878);
or U1140 (N_1140,N_839,N_862);
or U1141 (N_1141,N_921,N_848);
nand U1142 (N_1142,N_870,N_835);
or U1143 (N_1143,N_905,N_934);
or U1144 (N_1144,N_861,N_935);
nor U1145 (N_1145,N_877,N_860);
nand U1146 (N_1146,N_845,N_931);
and U1147 (N_1147,N_840,N_982);
or U1148 (N_1148,N_877,N_876);
nand U1149 (N_1149,N_861,N_811);
or U1150 (N_1150,N_833,N_874);
nor U1151 (N_1151,N_883,N_933);
and U1152 (N_1152,N_926,N_875);
nor U1153 (N_1153,N_801,N_926);
or U1154 (N_1154,N_890,N_999);
or U1155 (N_1155,N_973,N_883);
nand U1156 (N_1156,N_987,N_941);
nor U1157 (N_1157,N_991,N_955);
and U1158 (N_1158,N_813,N_881);
nor U1159 (N_1159,N_855,N_812);
nor U1160 (N_1160,N_919,N_812);
nor U1161 (N_1161,N_913,N_872);
and U1162 (N_1162,N_995,N_819);
nor U1163 (N_1163,N_834,N_877);
nor U1164 (N_1164,N_825,N_805);
or U1165 (N_1165,N_840,N_959);
nand U1166 (N_1166,N_988,N_806);
nor U1167 (N_1167,N_970,N_829);
nor U1168 (N_1168,N_815,N_859);
or U1169 (N_1169,N_823,N_912);
nand U1170 (N_1170,N_931,N_854);
nand U1171 (N_1171,N_837,N_968);
or U1172 (N_1172,N_934,N_976);
nor U1173 (N_1173,N_893,N_828);
and U1174 (N_1174,N_853,N_878);
nor U1175 (N_1175,N_803,N_958);
or U1176 (N_1176,N_825,N_969);
nand U1177 (N_1177,N_851,N_844);
and U1178 (N_1178,N_800,N_915);
and U1179 (N_1179,N_871,N_888);
and U1180 (N_1180,N_967,N_919);
nor U1181 (N_1181,N_985,N_884);
or U1182 (N_1182,N_821,N_909);
nor U1183 (N_1183,N_950,N_961);
or U1184 (N_1184,N_801,N_960);
nor U1185 (N_1185,N_860,N_944);
nand U1186 (N_1186,N_897,N_907);
nor U1187 (N_1187,N_876,N_803);
nor U1188 (N_1188,N_833,N_923);
and U1189 (N_1189,N_932,N_853);
and U1190 (N_1190,N_811,N_952);
or U1191 (N_1191,N_856,N_833);
nor U1192 (N_1192,N_913,N_934);
xnor U1193 (N_1193,N_964,N_993);
or U1194 (N_1194,N_898,N_875);
nor U1195 (N_1195,N_938,N_987);
or U1196 (N_1196,N_975,N_838);
and U1197 (N_1197,N_924,N_832);
nand U1198 (N_1198,N_986,N_972);
and U1199 (N_1199,N_914,N_969);
or U1200 (N_1200,N_1172,N_1169);
or U1201 (N_1201,N_1117,N_1018);
nand U1202 (N_1202,N_1083,N_1016);
nor U1203 (N_1203,N_1140,N_1154);
nor U1204 (N_1204,N_1006,N_1070);
nand U1205 (N_1205,N_1021,N_1015);
or U1206 (N_1206,N_1056,N_1012);
nor U1207 (N_1207,N_1050,N_1030);
or U1208 (N_1208,N_1065,N_1183);
and U1209 (N_1209,N_1168,N_1158);
nand U1210 (N_1210,N_1123,N_1141);
nor U1211 (N_1211,N_1062,N_1106);
or U1212 (N_1212,N_1101,N_1185);
and U1213 (N_1213,N_1026,N_1167);
nor U1214 (N_1214,N_1010,N_1053);
or U1215 (N_1215,N_1043,N_1113);
and U1216 (N_1216,N_1142,N_1092);
nand U1217 (N_1217,N_1130,N_1115);
xor U1218 (N_1218,N_1046,N_1198);
xor U1219 (N_1219,N_1136,N_1013);
nor U1220 (N_1220,N_1004,N_1137);
or U1221 (N_1221,N_1180,N_1052);
nor U1222 (N_1222,N_1163,N_1190);
and U1223 (N_1223,N_1191,N_1093);
and U1224 (N_1224,N_1014,N_1039);
nor U1225 (N_1225,N_1189,N_1036);
or U1226 (N_1226,N_1160,N_1054);
and U1227 (N_1227,N_1104,N_1145);
and U1228 (N_1228,N_1034,N_1085);
nor U1229 (N_1229,N_1146,N_1131);
nor U1230 (N_1230,N_1061,N_1152);
or U1231 (N_1231,N_1143,N_1103);
xor U1232 (N_1232,N_1059,N_1111);
and U1233 (N_1233,N_1023,N_1066);
nand U1234 (N_1234,N_1008,N_1020);
or U1235 (N_1235,N_1124,N_1120);
or U1236 (N_1236,N_1017,N_1155);
nor U1237 (N_1237,N_1157,N_1077);
or U1238 (N_1238,N_1098,N_1024);
and U1239 (N_1239,N_1195,N_1074);
nand U1240 (N_1240,N_1082,N_1097);
nor U1241 (N_1241,N_1048,N_1071);
nor U1242 (N_1242,N_1086,N_1164);
nor U1243 (N_1243,N_1162,N_1011);
nor U1244 (N_1244,N_1139,N_1044);
nor U1245 (N_1245,N_1028,N_1109);
nor U1246 (N_1246,N_1073,N_1153);
nand U1247 (N_1247,N_1094,N_1116);
nand U1248 (N_1248,N_1081,N_1005);
nor U1249 (N_1249,N_1007,N_1122);
nand U1250 (N_1250,N_1177,N_1110);
nand U1251 (N_1251,N_1051,N_1089);
or U1252 (N_1252,N_1064,N_1058);
nor U1253 (N_1253,N_1133,N_1174);
nand U1254 (N_1254,N_1057,N_1184);
nand U1255 (N_1255,N_1068,N_1002);
nand U1256 (N_1256,N_1194,N_1105);
nor U1257 (N_1257,N_1129,N_1090);
nor U1258 (N_1258,N_1151,N_1192);
and U1259 (N_1259,N_1009,N_1118);
xnor U1260 (N_1260,N_1076,N_1038);
or U1261 (N_1261,N_1134,N_1128);
and U1262 (N_1262,N_1171,N_1173);
nand U1263 (N_1263,N_1080,N_1127);
nand U1264 (N_1264,N_1022,N_1186);
and U1265 (N_1265,N_1144,N_1108);
or U1266 (N_1266,N_1045,N_1135);
and U1267 (N_1267,N_1121,N_1000);
nor U1268 (N_1268,N_1170,N_1096);
or U1269 (N_1269,N_1035,N_1156);
or U1270 (N_1270,N_1119,N_1138);
nand U1271 (N_1271,N_1060,N_1072);
or U1272 (N_1272,N_1079,N_1025);
and U1273 (N_1273,N_1084,N_1161);
nor U1274 (N_1274,N_1037,N_1047);
or U1275 (N_1275,N_1078,N_1033);
or U1276 (N_1276,N_1067,N_1100);
nor U1277 (N_1277,N_1003,N_1087);
and U1278 (N_1278,N_1032,N_1040);
or U1279 (N_1279,N_1147,N_1027);
nor U1280 (N_1280,N_1112,N_1150);
and U1281 (N_1281,N_1001,N_1179);
or U1282 (N_1282,N_1091,N_1187);
and U1283 (N_1283,N_1099,N_1029);
and U1284 (N_1284,N_1075,N_1199);
nor U1285 (N_1285,N_1125,N_1197);
nor U1286 (N_1286,N_1132,N_1149);
or U1287 (N_1287,N_1196,N_1175);
or U1288 (N_1288,N_1182,N_1114);
nor U1289 (N_1289,N_1188,N_1166);
or U1290 (N_1290,N_1095,N_1148);
nor U1291 (N_1291,N_1193,N_1178);
and U1292 (N_1292,N_1165,N_1107);
nor U1293 (N_1293,N_1176,N_1041);
nor U1294 (N_1294,N_1031,N_1102);
or U1295 (N_1295,N_1069,N_1049);
or U1296 (N_1296,N_1063,N_1159);
and U1297 (N_1297,N_1042,N_1019);
or U1298 (N_1298,N_1055,N_1088);
or U1299 (N_1299,N_1181,N_1126);
or U1300 (N_1300,N_1183,N_1177);
or U1301 (N_1301,N_1066,N_1080);
nor U1302 (N_1302,N_1079,N_1006);
and U1303 (N_1303,N_1101,N_1191);
nand U1304 (N_1304,N_1003,N_1152);
and U1305 (N_1305,N_1166,N_1092);
nand U1306 (N_1306,N_1137,N_1071);
and U1307 (N_1307,N_1195,N_1120);
nand U1308 (N_1308,N_1150,N_1078);
nor U1309 (N_1309,N_1177,N_1099);
nor U1310 (N_1310,N_1025,N_1068);
nand U1311 (N_1311,N_1080,N_1028);
nand U1312 (N_1312,N_1021,N_1035);
nor U1313 (N_1313,N_1015,N_1177);
or U1314 (N_1314,N_1140,N_1046);
nor U1315 (N_1315,N_1001,N_1155);
and U1316 (N_1316,N_1000,N_1099);
or U1317 (N_1317,N_1015,N_1019);
or U1318 (N_1318,N_1170,N_1079);
nand U1319 (N_1319,N_1171,N_1184);
nor U1320 (N_1320,N_1096,N_1032);
and U1321 (N_1321,N_1038,N_1035);
nand U1322 (N_1322,N_1166,N_1140);
nand U1323 (N_1323,N_1145,N_1063);
and U1324 (N_1324,N_1147,N_1156);
nor U1325 (N_1325,N_1038,N_1159);
nor U1326 (N_1326,N_1189,N_1065);
nand U1327 (N_1327,N_1139,N_1126);
and U1328 (N_1328,N_1172,N_1147);
and U1329 (N_1329,N_1062,N_1155);
or U1330 (N_1330,N_1149,N_1172);
nor U1331 (N_1331,N_1165,N_1082);
or U1332 (N_1332,N_1188,N_1064);
and U1333 (N_1333,N_1171,N_1049);
or U1334 (N_1334,N_1108,N_1139);
nand U1335 (N_1335,N_1137,N_1107);
and U1336 (N_1336,N_1199,N_1027);
and U1337 (N_1337,N_1191,N_1183);
and U1338 (N_1338,N_1063,N_1189);
nand U1339 (N_1339,N_1148,N_1181);
and U1340 (N_1340,N_1100,N_1156);
and U1341 (N_1341,N_1144,N_1046);
nand U1342 (N_1342,N_1127,N_1067);
or U1343 (N_1343,N_1029,N_1144);
and U1344 (N_1344,N_1084,N_1103);
or U1345 (N_1345,N_1104,N_1093);
and U1346 (N_1346,N_1130,N_1128);
or U1347 (N_1347,N_1127,N_1013);
nor U1348 (N_1348,N_1164,N_1111);
nand U1349 (N_1349,N_1172,N_1151);
and U1350 (N_1350,N_1089,N_1144);
or U1351 (N_1351,N_1071,N_1067);
or U1352 (N_1352,N_1181,N_1041);
nand U1353 (N_1353,N_1039,N_1172);
nor U1354 (N_1354,N_1103,N_1128);
nand U1355 (N_1355,N_1058,N_1091);
or U1356 (N_1356,N_1158,N_1025);
nand U1357 (N_1357,N_1123,N_1081);
or U1358 (N_1358,N_1175,N_1017);
and U1359 (N_1359,N_1027,N_1035);
or U1360 (N_1360,N_1061,N_1176);
nand U1361 (N_1361,N_1101,N_1134);
and U1362 (N_1362,N_1035,N_1130);
nand U1363 (N_1363,N_1147,N_1040);
nor U1364 (N_1364,N_1011,N_1021);
or U1365 (N_1365,N_1146,N_1172);
nand U1366 (N_1366,N_1130,N_1123);
nand U1367 (N_1367,N_1056,N_1083);
nand U1368 (N_1368,N_1140,N_1090);
nand U1369 (N_1369,N_1117,N_1027);
nand U1370 (N_1370,N_1081,N_1030);
and U1371 (N_1371,N_1042,N_1109);
or U1372 (N_1372,N_1066,N_1182);
and U1373 (N_1373,N_1001,N_1028);
and U1374 (N_1374,N_1157,N_1090);
and U1375 (N_1375,N_1029,N_1091);
nand U1376 (N_1376,N_1042,N_1013);
and U1377 (N_1377,N_1002,N_1171);
and U1378 (N_1378,N_1091,N_1031);
or U1379 (N_1379,N_1121,N_1161);
nand U1380 (N_1380,N_1037,N_1145);
or U1381 (N_1381,N_1168,N_1113);
and U1382 (N_1382,N_1145,N_1073);
or U1383 (N_1383,N_1130,N_1114);
nor U1384 (N_1384,N_1051,N_1136);
xor U1385 (N_1385,N_1070,N_1152);
nor U1386 (N_1386,N_1001,N_1092);
nand U1387 (N_1387,N_1113,N_1122);
and U1388 (N_1388,N_1014,N_1037);
xnor U1389 (N_1389,N_1164,N_1014);
nor U1390 (N_1390,N_1065,N_1136);
nand U1391 (N_1391,N_1031,N_1063);
nor U1392 (N_1392,N_1094,N_1125);
nand U1393 (N_1393,N_1011,N_1136);
or U1394 (N_1394,N_1086,N_1027);
and U1395 (N_1395,N_1199,N_1060);
or U1396 (N_1396,N_1040,N_1053);
nand U1397 (N_1397,N_1139,N_1019);
or U1398 (N_1398,N_1135,N_1043);
nor U1399 (N_1399,N_1070,N_1047);
and U1400 (N_1400,N_1387,N_1230);
and U1401 (N_1401,N_1225,N_1228);
nor U1402 (N_1402,N_1216,N_1292);
and U1403 (N_1403,N_1311,N_1386);
or U1404 (N_1404,N_1284,N_1276);
or U1405 (N_1405,N_1394,N_1278);
or U1406 (N_1406,N_1294,N_1347);
nor U1407 (N_1407,N_1378,N_1302);
nand U1408 (N_1408,N_1371,N_1330);
nand U1409 (N_1409,N_1391,N_1383);
nand U1410 (N_1410,N_1261,N_1293);
or U1411 (N_1411,N_1325,N_1344);
or U1412 (N_1412,N_1301,N_1247);
nand U1413 (N_1413,N_1314,N_1291);
nand U1414 (N_1414,N_1323,N_1359);
and U1415 (N_1415,N_1237,N_1223);
nand U1416 (N_1416,N_1262,N_1218);
or U1417 (N_1417,N_1370,N_1274);
nor U1418 (N_1418,N_1339,N_1307);
nor U1419 (N_1419,N_1285,N_1235);
nand U1420 (N_1420,N_1376,N_1310);
nand U1421 (N_1421,N_1268,N_1354);
nand U1422 (N_1422,N_1340,N_1254);
nand U1423 (N_1423,N_1288,N_1306);
or U1424 (N_1424,N_1249,N_1279);
nor U1425 (N_1425,N_1229,N_1267);
nand U1426 (N_1426,N_1318,N_1243);
nand U1427 (N_1427,N_1342,N_1263);
and U1428 (N_1428,N_1208,N_1260);
nand U1429 (N_1429,N_1255,N_1374);
or U1430 (N_1430,N_1227,N_1313);
and U1431 (N_1431,N_1205,N_1281);
and U1432 (N_1432,N_1283,N_1331);
nand U1433 (N_1433,N_1369,N_1206);
nand U1434 (N_1434,N_1303,N_1353);
and U1435 (N_1435,N_1280,N_1209);
or U1436 (N_1436,N_1326,N_1214);
nand U1437 (N_1437,N_1327,N_1346);
or U1438 (N_1438,N_1385,N_1265);
and U1439 (N_1439,N_1329,N_1357);
nand U1440 (N_1440,N_1343,N_1337);
nor U1441 (N_1441,N_1304,N_1211);
or U1442 (N_1442,N_1350,N_1202);
nand U1443 (N_1443,N_1392,N_1246);
nor U1444 (N_1444,N_1287,N_1221);
and U1445 (N_1445,N_1201,N_1351);
and U1446 (N_1446,N_1258,N_1236);
nand U1447 (N_1447,N_1298,N_1286);
nand U1448 (N_1448,N_1319,N_1389);
and U1449 (N_1449,N_1253,N_1240);
nor U1450 (N_1450,N_1360,N_1365);
or U1451 (N_1451,N_1200,N_1309);
nand U1452 (N_1452,N_1396,N_1308);
and U1453 (N_1453,N_1297,N_1317);
and U1454 (N_1454,N_1231,N_1372);
or U1455 (N_1455,N_1244,N_1256);
and U1456 (N_1456,N_1375,N_1275);
nand U1457 (N_1457,N_1393,N_1204);
nand U1458 (N_1458,N_1397,N_1271);
or U1459 (N_1459,N_1232,N_1356);
nor U1460 (N_1460,N_1245,N_1358);
nand U1461 (N_1461,N_1373,N_1224);
nor U1462 (N_1462,N_1315,N_1251);
nand U1463 (N_1463,N_1273,N_1366);
or U1464 (N_1464,N_1238,N_1215);
or U1465 (N_1465,N_1295,N_1277);
nor U1466 (N_1466,N_1381,N_1361);
nand U1467 (N_1467,N_1334,N_1270);
and U1468 (N_1468,N_1322,N_1355);
xnor U1469 (N_1469,N_1364,N_1226);
and U1470 (N_1470,N_1395,N_1399);
or U1471 (N_1471,N_1217,N_1349);
nor U1472 (N_1472,N_1252,N_1382);
or U1473 (N_1473,N_1335,N_1296);
or U1474 (N_1474,N_1212,N_1380);
nand U1475 (N_1475,N_1272,N_1220);
nand U1476 (N_1476,N_1269,N_1352);
or U1477 (N_1477,N_1248,N_1362);
nor U1478 (N_1478,N_1320,N_1289);
or U1479 (N_1479,N_1321,N_1324);
and U1480 (N_1480,N_1259,N_1241);
and U1481 (N_1481,N_1300,N_1312);
nor U1482 (N_1482,N_1379,N_1377);
and U1483 (N_1483,N_1338,N_1333);
or U1484 (N_1484,N_1282,N_1328);
or U1485 (N_1485,N_1368,N_1316);
nor U1486 (N_1486,N_1266,N_1336);
nor U1487 (N_1487,N_1348,N_1207);
nor U1488 (N_1488,N_1290,N_1332);
xnor U1489 (N_1489,N_1222,N_1388);
nand U1490 (N_1490,N_1345,N_1363);
nor U1491 (N_1491,N_1257,N_1398);
nand U1492 (N_1492,N_1203,N_1239);
and U1493 (N_1493,N_1367,N_1390);
nor U1494 (N_1494,N_1250,N_1341);
nor U1495 (N_1495,N_1264,N_1384);
or U1496 (N_1496,N_1305,N_1233);
nor U1497 (N_1497,N_1234,N_1299);
nor U1498 (N_1498,N_1242,N_1210);
nor U1499 (N_1499,N_1219,N_1213);
xor U1500 (N_1500,N_1248,N_1324);
nor U1501 (N_1501,N_1219,N_1315);
nand U1502 (N_1502,N_1285,N_1323);
or U1503 (N_1503,N_1276,N_1363);
or U1504 (N_1504,N_1305,N_1227);
nand U1505 (N_1505,N_1202,N_1354);
nor U1506 (N_1506,N_1393,N_1232);
nor U1507 (N_1507,N_1387,N_1323);
or U1508 (N_1508,N_1231,N_1353);
nand U1509 (N_1509,N_1338,N_1200);
nand U1510 (N_1510,N_1305,N_1377);
nor U1511 (N_1511,N_1251,N_1246);
nand U1512 (N_1512,N_1261,N_1203);
or U1513 (N_1513,N_1234,N_1344);
nand U1514 (N_1514,N_1323,N_1311);
nor U1515 (N_1515,N_1233,N_1387);
or U1516 (N_1516,N_1362,N_1236);
nor U1517 (N_1517,N_1255,N_1348);
and U1518 (N_1518,N_1307,N_1358);
nand U1519 (N_1519,N_1250,N_1303);
and U1520 (N_1520,N_1392,N_1351);
nand U1521 (N_1521,N_1235,N_1357);
nor U1522 (N_1522,N_1350,N_1317);
nand U1523 (N_1523,N_1327,N_1296);
nor U1524 (N_1524,N_1335,N_1311);
nor U1525 (N_1525,N_1301,N_1271);
nor U1526 (N_1526,N_1302,N_1393);
nor U1527 (N_1527,N_1345,N_1326);
nor U1528 (N_1528,N_1349,N_1321);
nor U1529 (N_1529,N_1259,N_1213);
or U1530 (N_1530,N_1224,N_1201);
nand U1531 (N_1531,N_1303,N_1228);
nand U1532 (N_1532,N_1270,N_1367);
or U1533 (N_1533,N_1326,N_1328);
nand U1534 (N_1534,N_1221,N_1397);
xnor U1535 (N_1535,N_1276,N_1360);
and U1536 (N_1536,N_1362,N_1267);
nand U1537 (N_1537,N_1297,N_1378);
nor U1538 (N_1538,N_1332,N_1386);
and U1539 (N_1539,N_1308,N_1289);
or U1540 (N_1540,N_1301,N_1394);
nand U1541 (N_1541,N_1245,N_1299);
and U1542 (N_1542,N_1249,N_1285);
or U1543 (N_1543,N_1335,N_1308);
and U1544 (N_1544,N_1307,N_1361);
nor U1545 (N_1545,N_1284,N_1399);
nand U1546 (N_1546,N_1337,N_1380);
nor U1547 (N_1547,N_1250,N_1297);
nand U1548 (N_1548,N_1233,N_1237);
or U1549 (N_1549,N_1259,N_1243);
and U1550 (N_1550,N_1364,N_1385);
nand U1551 (N_1551,N_1341,N_1324);
nor U1552 (N_1552,N_1309,N_1241);
or U1553 (N_1553,N_1250,N_1316);
nor U1554 (N_1554,N_1292,N_1339);
nand U1555 (N_1555,N_1301,N_1294);
or U1556 (N_1556,N_1259,N_1262);
nand U1557 (N_1557,N_1283,N_1221);
nand U1558 (N_1558,N_1209,N_1204);
and U1559 (N_1559,N_1284,N_1340);
nor U1560 (N_1560,N_1241,N_1390);
and U1561 (N_1561,N_1382,N_1280);
or U1562 (N_1562,N_1373,N_1318);
nand U1563 (N_1563,N_1331,N_1261);
nor U1564 (N_1564,N_1202,N_1324);
or U1565 (N_1565,N_1229,N_1242);
nand U1566 (N_1566,N_1243,N_1274);
or U1567 (N_1567,N_1313,N_1259);
and U1568 (N_1568,N_1346,N_1228);
nor U1569 (N_1569,N_1239,N_1341);
nor U1570 (N_1570,N_1253,N_1250);
nand U1571 (N_1571,N_1330,N_1366);
or U1572 (N_1572,N_1315,N_1227);
nor U1573 (N_1573,N_1347,N_1240);
nand U1574 (N_1574,N_1241,N_1271);
nand U1575 (N_1575,N_1357,N_1342);
nor U1576 (N_1576,N_1320,N_1264);
nand U1577 (N_1577,N_1214,N_1240);
or U1578 (N_1578,N_1278,N_1373);
and U1579 (N_1579,N_1234,N_1218);
or U1580 (N_1580,N_1302,N_1221);
or U1581 (N_1581,N_1283,N_1238);
and U1582 (N_1582,N_1355,N_1257);
nand U1583 (N_1583,N_1303,N_1246);
and U1584 (N_1584,N_1398,N_1393);
and U1585 (N_1585,N_1267,N_1273);
and U1586 (N_1586,N_1262,N_1219);
and U1587 (N_1587,N_1322,N_1209);
nor U1588 (N_1588,N_1288,N_1356);
nand U1589 (N_1589,N_1361,N_1335);
or U1590 (N_1590,N_1365,N_1395);
and U1591 (N_1591,N_1307,N_1372);
and U1592 (N_1592,N_1341,N_1251);
and U1593 (N_1593,N_1245,N_1219);
and U1594 (N_1594,N_1352,N_1278);
nor U1595 (N_1595,N_1233,N_1306);
nor U1596 (N_1596,N_1280,N_1291);
nand U1597 (N_1597,N_1309,N_1268);
or U1598 (N_1598,N_1399,N_1249);
and U1599 (N_1599,N_1225,N_1284);
nor U1600 (N_1600,N_1406,N_1560);
and U1601 (N_1601,N_1517,N_1515);
nand U1602 (N_1602,N_1443,N_1558);
nor U1603 (N_1603,N_1401,N_1564);
nor U1604 (N_1604,N_1538,N_1599);
or U1605 (N_1605,N_1415,N_1403);
or U1606 (N_1606,N_1500,N_1594);
nand U1607 (N_1607,N_1405,N_1510);
or U1608 (N_1608,N_1530,N_1485);
or U1609 (N_1609,N_1489,N_1459);
nand U1610 (N_1610,N_1471,N_1573);
or U1611 (N_1611,N_1547,N_1446);
nand U1612 (N_1612,N_1408,N_1523);
and U1613 (N_1613,N_1435,N_1456);
and U1614 (N_1614,N_1482,N_1429);
and U1615 (N_1615,N_1535,N_1585);
nand U1616 (N_1616,N_1514,N_1484);
nand U1617 (N_1617,N_1404,N_1513);
and U1618 (N_1618,N_1498,N_1568);
nand U1619 (N_1619,N_1424,N_1508);
xnor U1620 (N_1620,N_1587,N_1527);
nor U1621 (N_1621,N_1522,N_1409);
nand U1622 (N_1622,N_1411,N_1524);
and U1623 (N_1623,N_1569,N_1575);
nand U1624 (N_1624,N_1468,N_1539);
nor U1625 (N_1625,N_1525,N_1554);
and U1626 (N_1626,N_1467,N_1534);
nand U1627 (N_1627,N_1453,N_1462);
nor U1628 (N_1628,N_1502,N_1416);
nand U1629 (N_1629,N_1487,N_1407);
nor U1630 (N_1630,N_1496,N_1447);
nand U1631 (N_1631,N_1437,N_1563);
or U1632 (N_1632,N_1492,N_1476);
and U1633 (N_1633,N_1532,N_1555);
nand U1634 (N_1634,N_1440,N_1444);
xnor U1635 (N_1635,N_1590,N_1592);
and U1636 (N_1636,N_1549,N_1457);
or U1637 (N_1637,N_1458,N_1509);
nand U1638 (N_1638,N_1507,N_1475);
nand U1639 (N_1639,N_1448,N_1561);
and U1640 (N_1640,N_1412,N_1543);
and U1641 (N_1641,N_1491,N_1520);
or U1642 (N_1642,N_1551,N_1578);
nand U1643 (N_1643,N_1544,N_1503);
nor U1644 (N_1644,N_1478,N_1497);
nor U1645 (N_1645,N_1533,N_1531);
and U1646 (N_1646,N_1537,N_1418);
or U1647 (N_1647,N_1425,N_1574);
or U1648 (N_1648,N_1432,N_1516);
or U1649 (N_1649,N_1477,N_1505);
nor U1650 (N_1650,N_1460,N_1450);
nand U1651 (N_1651,N_1583,N_1434);
nor U1652 (N_1652,N_1494,N_1566);
and U1653 (N_1653,N_1422,N_1421);
and U1654 (N_1654,N_1546,N_1529);
and U1655 (N_1655,N_1466,N_1596);
or U1656 (N_1656,N_1490,N_1427);
or U1657 (N_1657,N_1483,N_1428);
nand U1658 (N_1658,N_1519,N_1548);
and U1659 (N_1659,N_1451,N_1545);
nor U1660 (N_1660,N_1526,N_1439);
and U1661 (N_1661,N_1442,N_1598);
and U1662 (N_1662,N_1511,N_1413);
nor U1663 (N_1663,N_1480,N_1586);
or U1664 (N_1664,N_1576,N_1463);
nand U1665 (N_1665,N_1430,N_1572);
nand U1666 (N_1666,N_1506,N_1495);
and U1667 (N_1667,N_1402,N_1419);
or U1668 (N_1668,N_1474,N_1571);
or U1669 (N_1669,N_1562,N_1454);
nand U1670 (N_1670,N_1552,N_1465);
and U1671 (N_1671,N_1595,N_1559);
or U1672 (N_1672,N_1581,N_1540);
nor U1673 (N_1673,N_1486,N_1436);
nand U1674 (N_1674,N_1504,N_1433);
or U1675 (N_1675,N_1423,N_1501);
nor U1676 (N_1676,N_1536,N_1582);
nor U1677 (N_1677,N_1445,N_1550);
or U1678 (N_1678,N_1449,N_1567);
and U1679 (N_1679,N_1410,N_1493);
nand U1680 (N_1680,N_1469,N_1441);
nor U1681 (N_1681,N_1461,N_1473);
or U1682 (N_1682,N_1499,N_1464);
nor U1683 (N_1683,N_1417,N_1481);
nand U1684 (N_1684,N_1579,N_1521);
and U1685 (N_1685,N_1472,N_1479);
and U1686 (N_1686,N_1488,N_1470);
nor U1687 (N_1687,N_1584,N_1420);
xnor U1688 (N_1688,N_1553,N_1400);
nand U1689 (N_1689,N_1577,N_1414);
and U1690 (N_1690,N_1426,N_1431);
nand U1691 (N_1691,N_1557,N_1542);
nand U1692 (N_1692,N_1588,N_1518);
and U1693 (N_1693,N_1528,N_1597);
nand U1694 (N_1694,N_1455,N_1438);
nand U1695 (N_1695,N_1570,N_1556);
or U1696 (N_1696,N_1593,N_1512);
or U1697 (N_1697,N_1589,N_1452);
and U1698 (N_1698,N_1580,N_1541);
and U1699 (N_1699,N_1565,N_1591);
nor U1700 (N_1700,N_1400,N_1466);
and U1701 (N_1701,N_1537,N_1476);
or U1702 (N_1702,N_1419,N_1439);
and U1703 (N_1703,N_1433,N_1512);
xor U1704 (N_1704,N_1435,N_1589);
or U1705 (N_1705,N_1444,N_1581);
and U1706 (N_1706,N_1593,N_1529);
or U1707 (N_1707,N_1534,N_1479);
nand U1708 (N_1708,N_1463,N_1471);
or U1709 (N_1709,N_1563,N_1438);
or U1710 (N_1710,N_1551,N_1461);
or U1711 (N_1711,N_1489,N_1583);
xor U1712 (N_1712,N_1560,N_1512);
and U1713 (N_1713,N_1429,N_1582);
nor U1714 (N_1714,N_1470,N_1409);
or U1715 (N_1715,N_1447,N_1554);
nand U1716 (N_1716,N_1513,N_1495);
and U1717 (N_1717,N_1527,N_1429);
or U1718 (N_1718,N_1477,N_1492);
nand U1719 (N_1719,N_1534,N_1461);
and U1720 (N_1720,N_1535,N_1545);
or U1721 (N_1721,N_1565,N_1472);
and U1722 (N_1722,N_1437,N_1444);
or U1723 (N_1723,N_1572,N_1438);
and U1724 (N_1724,N_1498,N_1464);
nand U1725 (N_1725,N_1513,N_1430);
and U1726 (N_1726,N_1524,N_1589);
or U1727 (N_1727,N_1407,N_1570);
nand U1728 (N_1728,N_1447,N_1597);
and U1729 (N_1729,N_1505,N_1456);
nand U1730 (N_1730,N_1515,N_1533);
and U1731 (N_1731,N_1552,N_1560);
nor U1732 (N_1732,N_1498,N_1574);
nand U1733 (N_1733,N_1411,N_1547);
nor U1734 (N_1734,N_1530,N_1452);
nand U1735 (N_1735,N_1544,N_1577);
nand U1736 (N_1736,N_1554,N_1541);
nor U1737 (N_1737,N_1495,N_1470);
nor U1738 (N_1738,N_1419,N_1503);
nor U1739 (N_1739,N_1487,N_1459);
and U1740 (N_1740,N_1580,N_1577);
nor U1741 (N_1741,N_1581,N_1446);
nor U1742 (N_1742,N_1543,N_1513);
nor U1743 (N_1743,N_1517,N_1586);
and U1744 (N_1744,N_1456,N_1565);
or U1745 (N_1745,N_1410,N_1432);
and U1746 (N_1746,N_1467,N_1524);
or U1747 (N_1747,N_1490,N_1428);
and U1748 (N_1748,N_1463,N_1580);
nand U1749 (N_1749,N_1533,N_1558);
nand U1750 (N_1750,N_1468,N_1487);
nand U1751 (N_1751,N_1484,N_1526);
nand U1752 (N_1752,N_1558,N_1524);
and U1753 (N_1753,N_1425,N_1441);
nand U1754 (N_1754,N_1516,N_1515);
nand U1755 (N_1755,N_1590,N_1419);
or U1756 (N_1756,N_1571,N_1432);
nor U1757 (N_1757,N_1473,N_1535);
nand U1758 (N_1758,N_1579,N_1520);
or U1759 (N_1759,N_1455,N_1533);
nor U1760 (N_1760,N_1538,N_1591);
or U1761 (N_1761,N_1500,N_1410);
or U1762 (N_1762,N_1505,N_1541);
nand U1763 (N_1763,N_1481,N_1441);
and U1764 (N_1764,N_1504,N_1476);
nand U1765 (N_1765,N_1583,N_1568);
nor U1766 (N_1766,N_1448,N_1447);
nand U1767 (N_1767,N_1449,N_1495);
nand U1768 (N_1768,N_1495,N_1494);
or U1769 (N_1769,N_1573,N_1444);
or U1770 (N_1770,N_1533,N_1513);
nand U1771 (N_1771,N_1572,N_1476);
or U1772 (N_1772,N_1554,N_1483);
nand U1773 (N_1773,N_1507,N_1567);
nand U1774 (N_1774,N_1519,N_1430);
nor U1775 (N_1775,N_1485,N_1537);
nor U1776 (N_1776,N_1478,N_1582);
and U1777 (N_1777,N_1561,N_1466);
nor U1778 (N_1778,N_1449,N_1457);
or U1779 (N_1779,N_1475,N_1405);
xor U1780 (N_1780,N_1592,N_1435);
or U1781 (N_1781,N_1461,N_1518);
or U1782 (N_1782,N_1474,N_1427);
nand U1783 (N_1783,N_1478,N_1463);
or U1784 (N_1784,N_1571,N_1413);
nor U1785 (N_1785,N_1491,N_1557);
nor U1786 (N_1786,N_1453,N_1587);
and U1787 (N_1787,N_1531,N_1554);
nor U1788 (N_1788,N_1479,N_1579);
or U1789 (N_1789,N_1423,N_1573);
nand U1790 (N_1790,N_1410,N_1401);
and U1791 (N_1791,N_1519,N_1532);
and U1792 (N_1792,N_1591,N_1467);
nor U1793 (N_1793,N_1423,N_1424);
nand U1794 (N_1794,N_1461,N_1530);
and U1795 (N_1795,N_1544,N_1564);
or U1796 (N_1796,N_1476,N_1553);
nand U1797 (N_1797,N_1501,N_1475);
and U1798 (N_1798,N_1459,N_1562);
and U1799 (N_1799,N_1491,N_1509);
nand U1800 (N_1800,N_1736,N_1671);
nand U1801 (N_1801,N_1641,N_1730);
nor U1802 (N_1802,N_1630,N_1746);
and U1803 (N_1803,N_1643,N_1667);
or U1804 (N_1804,N_1642,N_1732);
or U1805 (N_1805,N_1632,N_1607);
nor U1806 (N_1806,N_1769,N_1647);
or U1807 (N_1807,N_1770,N_1706);
nor U1808 (N_1808,N_1619,N_1654);
or U1809 (N_1809,N_1628,N_1659);
or U1810 (N_1810,N_1629,N_1681);
and U1811 (N_1811,N_1758,N_1756);
nor U1812 (N_1812,N_1783,N_1785);
nor U1813 (N_1813,N_1744,N_1743);
and U1814 (N_1814,N_1793,N_1613);
and U1815 (N_1815,N_1658,N_1677);
or U1816 (N_1816,N_1765,N_1788);
nor U1817 (N_1817,N_1738,N_1694);
nor U1818 (N_1818,N_1734,N_1676);
and U1819 (N_1819,N_1776,N_1764);
nor U1820 (N_1820,N_1726,N_1768);
and U1821 (N_1821,N_1648,N_1655);
nor U1822 (N_1822,N_1686,N_1645);
nand U1823 (N_1823,N_1622,N_1751);
nand U1824 (N_1824,N_1737,N_1650);
nor U1825 (N_1825,N_1623,N_1749);
nor U1826 (N_1826,N_1710,N_1675);
nor U1827 (N_1827,N_1774,N_1733);
nor U1828 (N_1828,N_1773,N_1798);
nor U1829 (N_1829,N_1618,N_1684);
nor U1830 (N_1830,N_1636,N_1704);
nor U1831 (N_1831,N_1712,N_1673);
or U1832 (N_1832,N_1724,N_1797);
and U1833 (N_1833,N_1719,N_1617);
or U1834 (N_1834,N_1646,N_1766);
or U1835 (N_1835,N_1729,N_1669);
or U1836 (N_1836,N_1674,N_1721);
nand U1837 (N_1837,N_1735,N_1755);
nor U1838 (N_1838,N_1626,N_1631);
or U1839 (N_1839,N_1668,N_1621);
nand U1840 (N_1840,N_1602,N_1692);
nand U1841 (N_1841,N_1731,N_1711);
or U1842 (N_1842,N_1705,N_1615);
nand U1843 (N_1843,N_1723,N_1759);
nor U1844 (N_1844,N_1653,N_1604);
nand U1845 (N_1845,N_1662,N_1791);
and U1846 (N_1846,N_1624,N_1634);
nand U1847 (N_1847,N_1687,N_1666);
and U1848 (N_1848,N_1695,N_1767);
and U1849 (N_1849,N_1600,N_1644);
and U1850 (N_1850,N_1657,N_1635);
or U1851 (N_1851,N_1728,N_1780);
or U1852 (N_1852,N_1727,N_1638);
nor U1853 (N_1853,N_1703,N_1790);
nor U1854 (N_1854,N_1777,N_1656);
nor U1855 (N_1855,N_1649,N_1661);
nand U1856 (N_1856,N_1714,N_1665);
nand U1857 (N_1857,N_1725,N_1660);
or U1858 (N_1858,N_1796,N_1708);
or U1859 (N_1859,N_1688,N_1672);
and U1860 (N_1860,N_1750,N_1637);
or U1861 (N_1861,N_1606,N_1678);
or U1862 (N_1862,N_1612,N_1605);
nand U1863 (N_1863,N_1772,N_1745);
or U1864 (N_1864,N_1779,N_1761);
nand U1865 (N_1865,N_1640,N_1782);
nor U1866 (N_1866,N_1693,N_1789);
xnor U1867 (N_1867,N_1792,N_1718);
nor U1868 (N_1868,N_1757,N_1699);
or U1869 (N_1869,N_1609,N_1700);
or U1870 (N_1870,N_1799,N_1709);
and U1871 (N_1871,N_1753,N_1616);
nor U1872 (N_1872,N_1784,N_1625);
and U1873 (N_1873,N_1722,N_1760);
and U1874 (N_1874,N_1610,N_1762);
or U1875 (N_1875,N_1763,N_1794);
or U1876 (N_1876,N_1633,N_1787);
or U1877 (N_1877,N_1696,N_1781);
or U1878 (N_1878,N_1689,N_1752);
nand U1879 (N_1879,N_1664,N_1679);
or U1880 (N_1880,N_1739,N_1701);
and U1881 (N_1881,N_1747,N_1741);
or U1882 (N_1882,N_1717,N_1697);
nor U1883 (N_1883,N_1778,N_1652);
or U1884 (N_1884,N_1651,N_1748);
or U1885 (N_1885,N_1603,N_1713);
nand U1886 (N_1886,N_1707,N_1601);
or U1887 (N_1887,N_1754,N_1691);
nor U1888 (N_1888,N_1716,N_1683);
or U1889 (N_1889,N_1639,N_1786);
or U1890 (N_1890,N_1690,N_1627);
nor U1891 (N_1891,N_1742,N_1740);
or U1892 (N_1892,N_1771,N_1682);
nand U1893 (N_1893,N_1715,N_1670);
or U1894 (N_1894,N_1720,N_1611);
or U1895 (N_1895,N_1680,N_1620);
nand U1896 (N_1896,N_1698,N_1608);
nor U1897 (N_1897,N_1614,N_1702);
and U1898 (N_1898,N_1663,N_1775);
or U1899 (N_1899,N_1685,N_1795);
nor U1900 (N_1900,N_1766,N_1671);
and U1901 (N_1901,N_1703,N_1734);
xor U1902 (N_1902,N_1649,N_1610);
xor U1903 (N_1903,N_1666,N_1612);
nand U1904 (N_1904,N_1621,N_1798);
nor U1905 (N_1905,N_1751,N_1730);
nand U1906 (N_1906,N_1651,N_1738);
or U1907 (N_1907,N_1726,N_1610);
nand U1908 (N_1908,N_1677,N_1731);
nor U1909 (N_1909,N_1634,N_1601);
nor U1910 (N_1910,N_1776,N_1732);
or U1911 (N_1911,N_1680,N_1655);
xnor U1912 (N_1912,N_1641,N_1746);
nor U1913 (N_1913,N_1675,N_1677);
or U1914 (N_1914,N_1760,N_1724);
or U1915 (N_1915,N_1725,N_1639);
or U1916 (N_1916,N_1732,N_1604);
or U1917 (N_1917,N_1747,N_1661);
nor U1918 (N_1918,N_1739,N_1660);
and U1919 (N_1919,N_1797,N_1690);
nor U1920 (N_1920,N_1760,N_1731);
or U1921 (N_1921,N_1608,N_1627);
or U1922 (N_1922,N_1782,N_1772);
nand U1923 (N_1923,N_1723,N_1745);
or U1924 (N_1924,N_1729,N_1780);
or U1925 (N_1925,N_1719,N_1699);
nand U1926 (N_1926,N_1798,N_1702);
or U1927 (N_1927,N_1705,N_1782);
or U1928 (N_1928,N_1604,N_1674);
nor U1929 (N_1929,N_1717,N_1711);
nor U1930 (N_1930,N_1718,N_1697);
nand U1931 (N_1931,N_1694,N_1778);
nor U1932 (N_1932,N_1791,N_1734);
nor U1933 (N_1933,N_1674,N_1691);
nor U1934 (N_1934,N_1704,N_1771);
nor U1935 (N_1935,N_1739,N_1726);
or U1936 (N_1936,N_1693,N_1614);
or U1937 (N_1937,N_1779,N_1729);
and U1938 (N_1938,N_1614,N_1733);
nand U1939 (N_1939,N_1732,N_1609);
nor U1940 (N_1940,N_1630,N_1762);
nor U1941 (N_1941,N_1688,N_1741);
or U1942 (N_1942,N_1696,N_1713);
nand U1943 (N_1943,N_1622,N_1663);
nand U1944 (N_1944,N_1705,N_1703);
or U1945 (N_1945,N_1758,N_1766);
and U1946 (N_1946,N_1690,N_1695);
and U1947 (N_1947,N_1796,N_1749);
and U1948 (N_1948,N_1667,N_1602);
or U1949 (N_1949,N_1689,N_1710);
and U1950 (N_1950,N_1746,N_1718);
and U1951 (N_1951,N_1675,N_1668);
and U1952 (N_1952,N_1666,N_1794);
xor U1953 (N_1953,N_1757,N_1622);
and U1954 (N_1954,N_1729,N_1672);
nor U1955 (N_1955,N_1791,N_1745);
or U1956 (N_1956,N_1743,N_1778);
nor U1957 (N_1957,N_1627,N_1602);
or U1958 (N_1958,N_1721,N_1666);
and U1959 (N_1959,N_1652,N_1631);
nor U1960 (N_1960,N_1675,N_1690);
nor U1961 (N_1961,N_1747,N_1751);
or U1962 (N_1962,N_1745,N_1604);
or U1963 (N_1963,N_1757,N_1714);
nor U1964 (N_1964,N_1605,N_1604);
and U1965 (N_1965,N_1618,N_1763);
or U1966 (N_1966,N_1639,N_1770);
and U1967 (N_1967,N_1602,N_1660);
or U1968 (N_1968,N_1621,N_1715);
and U1969 (N_1969,N_1782,N_1729);
nand U1970 (N_1970,N_1743,N_1625);
and U1971 (N_1971,N_1741,N_1703);
and U1972 (N_1972,N_1634,N_1754);
and U1973 (N_1973,N_1715,N_1631);
nor U1974 (N_1974,N_1728,N_1710);
and U1975 (N_1975,N_1761,N_1660);
nor U1976 (N_1976,N_1716,N_1720);
nand U1977 (N_1977,N_1759,N_1666);
and U1978 (N_1978,N_1634,N_1623);
nand U1979 (N_1979,N_1635,N_1679);
and U1980 (N_1980,N_1606,N_1673);
nor U1981 (N_1981,N_1621,N_1712);
or U1982 (N_1982,N_1662,N_1722);
or U1983 (N_1983,N_1636,N_1728);
nor U1984 (N_1984,N_1794,N_1651);
or U1985 (N_1985,N_1666,N_1764);
nand U1986 (N_1986,N_1668,N_1760);
or U1987 (N_1987,N_1613,N_1733);
nand U1988 (N_1988,N_1709,N_1649);
or U1989 (N_1989,N_1650,N_1607);
nor U1990 (N_1990,N_1791,N_1660);
and U1991 (N_1991,N_1613,N_1654);
or U1992 (N_1992,N_1697,N_1726);
nor U1993 (N_1993,N_1773,N_1682);
nor U1994 (N_1994,N_1727,N_1752);
or U1995 (N_1995,N_1773,N_1615);
or U1996 (N_1996,N_1700,N_1715);
nor U1997 (N_1997,N_1630,N_1743);
nand U1998 (N_1998,N_1606,N_1717);
nand U1999 (N_1999,N_1734,N_1633);
nor U2000 (N_2000,N_1915,N_1823);
and U2001 (N_2001,N_1834,N_1814);
nand U2002 (N_2002,N_1907,N_1859);
nor U2003 (N_2003,N_1857,N_1992);
nand U2004 (N_2004,N_1961,N_1960);
or U2005 (N_2005,N_1901,N_1844);
and U2006 (N_2006,N_1995,N_1965);
or U2007 (N_2007,N_1886,N_1950);
or U2008 (N_2008,N_1988,N_1912);
or U2009 (N_2009,N_1941,N_1876);
nand U2010 (N_2010,N_1968,N_1926);
nand U2011 (N_2011,N_1999,N_1991);
nand U2012 (N_2012,N_1937,N_1863);
and U2013 (N_2013,N_1973,N_1980);
nor U2014 (N_2014,N_1986,N_1963);
or U2015 (N_2015,N_1864,N_1865);
and U2016 (N_2016,N_1852,N_1855);
and U2017 (N_2017,N_1874,N_1888);
nor U2018 (N_2018,N_1957,N_1841);
nor U2019 (N_2019,N_1867,N_1958);
nor U2020 (N_2020,N_1818,N_1933);
nor U2021 (N_2021,N_1889,N_1938);
and U2022 (N_2022,N_1908,N_1861);
nor U2023 (N_2023,N_1977,N_1948);
and U2024 (N_2024,N_1880,N_1824);
nor U2025 (N_2025,N_1930,N_1872);
nor U2026 (N_2026,N_1964,N_1913);
nand U2027 (N_2027,N_1928,N_1803);
or U2028 (N_2028,N_1800,N_1809);
or U2029 (N_2029,N_1842,N_1843);
xor U2030 (N_2030,N_1832,N_1891);
nor U2031 (N_2031,N_1984,N_1879);
nor U2032 (N_2032,N_1940,N_1827);
nand U2033 (N_2033,N_1982,N_1875);
and U2034 (N_2034,N_1946,N_1856);
nor U2035 (N_2035,N_1929,N_1810);
nand U2036 (N_2036,N_1944,N_1897);
nor U2037 (N_2037,N_1887,N_1830);
or U2038 (N_2038,N_1862,N_1975);
nor U2039 (N_2039,N_1945,N_1833);
nand U2040 (N_2040,N_1916,N_1839);
nor U2041 (N_2041,N_1909,N_1903);
nand U2042 (N_2042,N_1877,N_1836);
and U2043 (N_2043,N_1990,N_1936);
and U2044 (N_2044,N_1959,N_1802);
nor U2045 (N_2045,N_1881,N_1846);
and U2046 (N_2046,N_1893,N_1955);
nor U2047 (N_2047,N_1835,N_1983);
nor U2048 (N_2048,N_1837,N_1979);
and U2049 (N_2049,N_1898,N_1918);
nor U2050 (N_2050,N_1978,N_1858);
and U2051 (N_2051,N_1920,N_1817);
and U2052 (N_2052,N_1819,N_1974);
or U2053 (N_2053,N_1923,N_1813);
or U2054 (N_2054,N_1828,N_1801);
or U2055 (N_2055,N_1831,N_1847);
nand U2056 (N_2056,N_1812,N_1821);
and U2057 (N_2057,N_1849,N_1890);
and U2058 (N_2058,N_1943,N_1866);
nand U2059 (N_2059,N_1878,N_1970);
nand U2060 (N_2060,N_1829,N_1871);
and U2061 (N_2061,N_1935,N_1895);
nor U2062 (N_2062,N_1808,N_1868);
nor U2063 (N_2063,N_1870,N_1953);
or U2064 (N_2064,N_1805,N_1850);
nand U2065 (N_2065,N_1911,N_1922);
xor U2066 (N_2066,N_1994,N_1925);
or U2067 (N_2067,N_1996,N_1873);
or U2068 (N_2068,N_1972,N_1820);
or U2069 (N_2069,N_1917,N_1848);
and U2070 (N_2070,N_1838,N_1969);
nand U2071 (N_2071,N_1952,N_1899);
nand U2072 (N_2072,N_1906,N_1966);
nand U2073 (N_2073,N_1989,N_1804);
nor U2074 (N_2074,N_1845,N_1924);
and U2075 (N_2075,N_1900,N_1811);
or U2076 (N_2076,N_1851,N_1896);
and U2077 (N_2077,N_1942,N_1998);
nand U2078 (N_2078,N_1993,N_1905);
nor U2079 (N_2079,N_1919,N_1947);
and U2080 (N_2080,N_1854,N_1869);
nor U2081 (N_2081,N_1885,N_1949);
nand U2082 (N_2082,N_1939,N_1910);
or U2083 (N_2083,N_1822,N_1931);
and U2084 (N_2084,N_1997,N_1956);
and U2085 (N_2085,N_1894,N_1853);
nor U2086 (N_2086,N_1954,N_1902);
or U2087 (N_2087,N_1884,N_1807);
nand U2088 (N_2088,N_1904,N_1815);
nand U2089 (N_2089,N_1860,N_1971);
and U2090 (N_2090,N_1825,N_1921);
nor U2091 (N_2091,N_1962,N_1967);
nand U2092 (N_2092,N_1927,N_1987);
nor U2093 (N_2093,N_1826,N_1934);
or U2094 (N_2094,N_1892,N_1976);
or U2095 (N_2095,N_1882,N_1883);
nand U2096 (N_2096,N_1981,N_1816);
or U2097 (N_2097,N_1951,N_1806);
nor U2098 (N_2098,N_1840,N_1985);
nor U2099 (N_2099,N_1932,N_1914);
nand U2100 (N_2100,N_1911,N_1935);
or U2101 (N_2101,N_1905,N_1951);
or U2102 (N_2102,N_1987,N_1970);
nor U2103 (N_2103,N_1857,N_1924);
nand U2104 (N_2104,N_1999,N_1927);
nand U2105 (N_2105,N_1803,N_1957);
or U2106 (N_2106,N_1908,N_1957);
nor U2107 (N_2107,N_1876,N_1849);
nor U2108 (N_2108,N_1822,N_1937);
nand U2109 (N_2109,N_1857,N_1872);
nand U2110 (N_2110,N_1949,N_1957);
nor U2111 (N_2111,N_1862,N_1820);
and U2112 (N_2112,N_1885,N_1818);
nand U2113 (N_2113,N_1993,N_1939);
nand U2114 (N_2114,N_1807,N_1900);
nand U2115 (N_2115,N_1915,N_1979);
nor U2116 (N_2116,N_1810,N_1910);
or U2117 (N_2117,N_1849,N_1871);
nor U2118 (N_2118,N_1877,N_1938);
or U2119 (N_2119,N_1940,N_1917);
and U2120 (N_2120,N_1849,N_1979);
nand U2121 (N_2121,N_1993,N_1988);
nand U2122 (N_2122,N_1915,N_1853);
nand U2123 (N_2123,N_1842,N_1911);
or U2124 (N_2124,N_1898,N_1805);
nand U2125 (N_2125,N_1842,N_1954);
nand U2126 (N_2126,N_1902,N_1975);
and U2127 (N_2127,N_1881,N_1876);
and U2128 (N_2128,N_1825,N_1850);
nor U2129 (N_2129,N_1937,N_1952);
or U2130 (N_2130,N_1887,N_1829);
nor U2131 (N_2131,N_1914,N_1869);
nor U2132 (N_2132,N_1824,N_1975);
xor U2133 (N_2133,N_1857,N_1913);
nand U2134 (N_2134,N_1902,N_1822);
nand U2135 (N_2135,N_1881,N_1961);
and U2136 (N_2136,N_1942,N_1808);
nor U2137 (N_2137,N_1945,N_1987);
and U2138 (N_2138,N_1953,N_1864);
and U2139 (N_2139,N_1906,N_1920);
or U2140 (N_2140,N_1844,N_1874);
and U2141 (N_2141,N_1872,N_1938);
nand U2142 (N_2142,N_1927,N_1953);
nor U2143 (N_2143,N_1927,N_1941);
nand U2144 (N_2144,N_1848,N_1857);
and U2145 (N_2145,N_1899,N_1879);
nor U2146 (N_2146,N_1831,N_1992);
and U2147 (N_2147,N_1942,N_1959);
or U2148 (N_2148,N_1838,N_1951);
nor U2149 (N_2149,N_1955,N_1957);
nor U2150 (N_2150,N_1949,N_1895);
nand U2151 (N_2151,N_1873,N_1971);
or U2152 (N_2152,N_1925,N_1853);
and U2153 (N_2153,N_1840,N_1854);
and U2154 (N_2154,N_1983,N_1803);
nand U2155 (N_2155,N_1988,N_1914);
or U2156 (N_2156,N_1806,N_1854);
or U2157 (N_2157,N_1912,N_1984);
nand U2158 (N_2158,N_1874,N_1809);
and U2159 (N_2159,N_1962,N_1947);
and U2160 (N_2160,N_1945,N_1857);
and U2161 (N_2161,N_1986,N_1815);
nand U2162 (N_2162,N_1989,N_1964);
and U2163 (N_2163,N_1852,N_1934);
or U2164 (N_2164,N_1887,N_1880);
or U2165 (N_2165,N_1990,N_1857);
and U2166 (N_2166,N_1966,N_1900);
nand U2167 (N_2167,N_1898,N_1914);
or U2168 (N_2168,N_1904,N_1801);
or U2169 (N_2169,N_1937,N_1836);
or U2170 (N_2170,N_1816,N_1883);
and U2171 (N_2171,N_1808,N_1944);
and U2172 (N_2172,N_1837,N_1864);
and U2173 (N_2173,N_1924,N_1869);
and U2174 (N_2174,N_1862,N_1980);
and U2175 (N_2175,N_1907,N_1970);
nand U2176 (N_2176,N_1904,N_1912);
nand U2177 (N_2177,N_1904,N_1876);
or U2178 (N_2178,N_1895,N_1868);
or U2179 (N_2179,N_1952,N_1962);
and U2180 (N_2180,N_1909,N_1819);
or U2181 (N_2181,N_1825,N_1969);
or U2182 (N_2182,N_1834,N_1853);
nor U2183 (N_2183,N_1912,N_1920);
and U2184 (N_2184,N_1948,N_1826);
and U2185 (N_2185,N_1944,N_1896);
and U2186 (N_2186,N_1973,N_1844);
or U2187 (N_2187,N_1894,N_1863);
nor U2188 (N_2188,N_1859,N_1878);
nand U2189 (N_2189,N_1986,N_1906);
nand U2190 (N_2190,N_1903,N_1892);
and U2191 (N_2191,N_1844,N_1987);
or U2192 (N_2192,N_1893,N_1823);
or U2193 (N_2193,N_1847,N_1939);
or U2194 (N_2194,N_1804,N_1902);
and U2195 (N_2195,N_1880,N_1996);
nor U2196 (N_2196,N_1887,N_1909);
and U2197 (N_2197,N_1912,N_1978);
nor U2198 (N_2198,N_1855,N_1897);
nand U2199 (N_2199,N_1907,N_1815);
or U2200 (N_2200,N_2049,N_2150);
nor U2201 (N_2201,N_2035,N_2122);
nor U2202 (N_2202,N_2105,N_2017);
nand U2203 (N_2203,N_2086,N_2074);
nand U2204 (N_2204,N_2072,N_2084);
nand U2205 (N_2205,N_2158,N_2160);
nand U2206 (N_2206,N_2115,N_2162);
nor U2207 (N_2207,N_2143,N_2170);
and U2208 (N_2208,N_2075,N_2024);
nor U2209 (N_2209,N_2007,N_2040);
and U2210 (N_2210,N_2116,N_2023);
nor U2211 (N_2211,N_2113,N_2106);
or U2212 (N_2212,N_2124,N_2163);
or U2213 (N_2213,N_2192,N_2135);
nand U2214 (N_2214,N_2021,N_2019);
or U2215 (N_2215,N_2153,N_2175);
or U2216 (N_2216,N_2181,N_2148);
nand U2217 (N_2217,N_2125,N_2161);
and U2218 (N_2218,N_2048,N_2171);
and U2219 (N_2219,N_2144,N_2131);
and U2220 (N_2220,N_2002,N_2027);
or U2221 (N_2221,N_2031,N_2119);
or U2222 (N_2222,N_2093,N_2114);
nand U2223 (N_2223,N_2026,N_2195);
or U2224 (N_2224,N_2168,N_2110);
nand U2225 (N_2225,N_2070,N_2059);
and U2226 (N_2226,N_2184,N_2013);
nor U2227 (N_2227,N_2141,N_2029);
or U2228 (N_2228,N_2063,N_2069);
or U2229 (N_2229,N_2198,N_2130);
and U2230 (N_2230,N_2009,N_2111);
and U2231 (N_2231,N_2011,N_2095);
nor U2232 (N_2232,N_2134,N_2028);
nor U2233 (N_2233,N_2112,N_2041);
nand U2234 (N_2234,N_2052,N_2169);
nor U2235 (N_2235,N_2057,N_2078);
or U2236 (N_2236,N_2136,N_2145);
nand U2237 (N_2237,N_2046,N_2036);
and U2238 (N_2238,N_2118,N_2197);
and U2239 (N_2239,N_2058,N_2196);
and U2240 (N_2240,N_2194,N_2071);
nor U2241 (N_2241,N_2133,N_2199);
and U2242 (N_2242,N_2178,N_2172);
nand U2243 (N_2243,N_2188,N_2088);
and U2244 (N_2244,N_2102,N_2176);
and U2245 (N_2245,N_2025,N_2016);
nand U2246 (N_2246,N_2132,N_2065);
and U2247 (N_2247,N_2117,N_2109);
nor U2248 (N_2248,N_2053,N_2185);
nor U2249 (N_2249,N_2068,N_2047);
nand U2250 (N_2250,N_2008,N_2098);
nor U2251 (N_2251,N_2166,N_2087);
nor U2252 (N_2252,N_2120,N_2060);
nor U2253 (N_2253,N_2123,N_2000);
nor U2254 (N_2254,N_2155,N_2055);
and U2255 (N_2255,N_2152,N_2004);
nor U2256 (N_2256,N_2003,N_2129);
nor U2257 (N_2257,N_2146,N_2186);
or U2258 (N_2258,N_2030,N_2045);
nor U2259 (N_2259,N_2067,N_2103);
or U2260 (N_2260,N_2138,N_2179);
xor U2261 (N_2261,N_2061,N_2174);
xnor U2262 (N_2262,N_2050,N_2099);
nand U2263 (N_2263,N_2037,N_2080);
and U2264 (N_2264,N_2104,N_2092);
nor U2265 (N_2265,N_2164,N_2073);
and U2266 (N_2266,N_2020,N_2156);
xor U2267 (N_2267,N_2079,N_2051);
nand U2268 (N_2268,N_2066,N_2010);
nor U2269 (N_2269,N_2189,N_2139);
nand U2270 (N_2270,N_2137,N_2081);
nor U2271 (N_2271,N_2191,N_2147);
and U2272 (N_2272,N_2014,N_2151);
nor U2273 (N_2273,N_2167,N_2159);
or U2274 (N_2274,N_2018,N_2044);
nor U2275 (N_2275,N_2090,N_2190);
nand U2276 (N_2276,N_2082,N_2038);
and U2277 (N_2277,N_2062,N_2101);
and U2278 (N_2278,N_2085,N_2187);
nand U2279 (N_2279,N_2097,N_2173);
nand U2280 (N_2280,N_2182,N_2091);
nand U2281 (N_2281,N_2034,N_2165);
nand U2282 (N_2282,N_2022,N_2083);
or U2283 (N_2283,N_2127,N_2054);
nand U2284 (N_2284,N_2001,N_2126);
and U2285 (N_2285,N_2064,N_2154);
nand U2286 (N_2286,N_2128,N_2108);
and U2287 (N_2287,N_2077,N_2149);
nor U2288 (N_2288,N_2042,N_2177);
nor U2289 (N_2289,N_2180,N_2043);
and U2290 (N_2290,N_2094,N_2193);
nand U2291 (N_2291,N_2006,N_2032);
nor U2292 (N_2292,N_2096,N_2140);
xor U2293 (N_2293,N_2121,N_2076);
or U2294 (N_2294,N_2056,N_2012);
nand U2295 (N_2295,N_2005,N_2100);
nor U2296 (N_2296,N_2183,N_2157);
nor U2297 (N_2297,N_2015,N_2107);
and U2298 (N_2298,N_2033,N_2039);
and U2299 (N_2299,N_2142,N_2089);
or U2300 (N_2300,N_2124,N_2173);
nor U2301 (N_2301,N_2199,N_2113);
nand U2302 (N_2302,N_2180,N_2104);
nor U2303 (N_2303,N_2140,N_2138);
nor U2304 (N_2304,N_2007,N_2047);
and U2305 (N_2305,N_2148,N_2155);
nor U2306 (N_2306,N_2190,N_2068);
nand U2307 (N_2307,N_2186,N_2043);
or U2308 (N_2308,N_2096,N_2119);
nand U2309 (N_2309,N_2170,N_2184);
and U2310 (N_2310,N_2125,N_2153);
nand U2311 (N_2311,N_2032,N_2025);
or U2312 (N_2312,N_2107,N_2113);
nand U2313 (N_2313,N_2172,N_2005);
and U2314 (N_2314,N_2019,N_2095);
nor U2315 (N_2315,N_2056,N_2123);
nor U2316 (N_2316,N_2094,N_2183);
or U2317 (N_2317,N_2128,N_2129);
and U2318 (N_2318,N_2111,N_2168);
or U2319 (N_2319,N_2125,N_2058);
nand U2320 (N_2320,N_2186,N_2148);
and U2321 (N_2321,N_2091,N_2050);
nor U2322 (N_2322,N_2112,N_2176);
or U2323 (N_2323,N_2112,N_2188);
xor U2324 (N_2324,N_2142,N_2192);
nand U2325 (N_2325,N_2192,N_2170);
or U2326 (N_2326,N_2191,N_2164);
or U2327 (N_2327,N_2145,N_2079);
nand U2328 (N_2328,N_2104,N_2107);
nand U2329 (N_2329,N_2120,N_2140);
nand U2330 (N_2330,N_2173,N_2045);
nand U2331 (N_2331,N_2149,N_2159);
or U2332 (N_2332,N_2053,N_2052);
nand U2333 (N_2333,N_2081,N_2012);
and U2334 (N_2334,N_2047,N_2034);
nor U2335 (N_2335,N_2066,N_2113);
nor U2336 (N_2336,N_2069,N_2166);
nand U2337 (N_2337,N_2127,N_2175);
nor U2338 (N_2338,N_2135,N_2156);
or U2339 (N_2339,N_2197,N_2002);
and U2340 (N_2340,N_2134,N_2125);
or U2341 (N_2341,N_2007,N_2164);
and U2342 (N_2342,N_2042,N_2019);
or U2343 (N_2343,N_2080,N_2079);
and U2344 (N_2344,N_2124,N_2034);
and U2345 (N_2345,N_2004,N_2167);
xnor U2346 (N_2346,N_2108,N_2135);
or U2347 (N_2347,N_2057,N_2152);
nor U2348 (N_2348,N_2003,N_2106);
nor U2349 (N_2349,N_2118,N_2133);
or U2350 (N_2350,N_2001,N_2040);
nor U2351 (N_2351,N_2026,N_2093);
nand U2352 (N_2352,N_2104,N_2068);
nand U2353 (N_2353,N_2024,N_2014);
nor U2354 (N_2354,N_2159,N_2006);
or U2355 (N_2355,N_2142,N_2121);
and U2356 (N_2356,N_2040,N_2196);
nand U2357 (N_2357,N_2045,N_2163);
and U2358 (N_2358,N_2024,N_2015);
nand U2359 (N_2359,N_2179,N_2065);
and U2360 (N_2360,N_2159,N_2185);
nor U2361 (N_2361,N_2178,N_2159);
and U2362 (N_2362,N_2121,N_2100);
nand U2363 (N_2363,N_2116,N_2138);
or U2364 (N_2364,N_2160,N_2002);
and U2365 (N_2365,N_2001,N_2130);
and U2366 (N_2366,N_2183,N_2097);
and U2367 (N_2367,N_2011,N_2154);
xnor U2368 (N_2368,N_2144,N_2137);
nor U2369 (N_2369,N_2083,N_2072);
nand U2370 (N_2370,N_2141,N_2081);
nor U2371 (N_2371,N_2138,N_2174);
and U2372 (N_2372,N_2010,N_2003);
and U2373 (N_2373,N_2153,N_2161);
nand U2374 (N_2374,N_2003,N_2066);
nand U2375 (N_2375,N_2032,N_2136);
nand U2376 (N_2376,N_2080,N_2181);
or U2377 (N_2377,N_2187,N_2029);
and U2378 (N_2378,N_2090,N_2150);
and U2379 (N_2379,N_2181,N_2053);
or U2380 (N_2380,N_2078,N_2159);
nand U2381 (N_2381,N_2083,N_2104);
xor U2382 (N_2382,N_2177,N_2081);
or U2383 (N_2383,N_2067,N_2131);
nor U2384 (N_2384,N_2052,N_2050);
nand U2385 (N_2385,N_2020,N_2019);
or U2386 (N_2386,N_2022,N_2056);
or U2387 (N_2387,N_2032,N_2160);
nand U2388 (N_2388,N_2078,N_2175);
or U2389 (N_2389,N_2181,N_2059);
or U2390 (N_2390,N_2156,N_2136);
and U2391 (N_2391,N_2151,N_2109);
nor U2392 (N_2392,N_2000,N_2089);
or U2393 (N_2393,N_2062,N_2189);
and U2394 (N_2394,N_2178,N_2092);
nor U2395 (N_2395,N_2054,N_2078);
nand U2396 (N_2396,N_2017,N_2051);
nor U2397 (N_2397,N_2050,N_2141);
or U2398 (N_2398,N_2017,N_2080);
nor U2399 (N_2399,N_2016,N_2167);
and U2400 (N_2400,N_2367,N_2373);
or U2401 (N_2401,N_2392,N_2212);
nand U2402 (N_2402,N_2394,N_2331);
and U2403 (N_2403,N_2232,N_2345);
or U2404 (N_2404,N_2388,N_2281);
nand U2405 (N_2405,N_2280,N_2202);
and U2406 (N_2406,N_2380,N_2213);
and U2407 (N_2407,N_2353,N_2314);
or U2408 (N_2408,N_2270,N_2294);
or U2409 (N_2409,N_2205,N_2330);
nand U2410 (N_2410,N_2290,N_2275);
nand U2411 (N_2411,N_2297,N_2268);
or U2412 (N_2412,N_2333,N_2240);
nor U2413 (N_2413,N_2379,N_2256);
nor U2414 (N_2414,N_2376,N_2356);
and U2415 (N_2415,N_2340,N_2233);
and U2416 (N_2416,N_2234,N_2245);
nand U2417 (N_2417,N_2239,N_2271);
and U2418 (N_2418,N_2282,N_2378);
or U2419 (N_2419,N_2273,N_2386);
nor U2420 (N_2420,N_2387,N_2288);
and U2421 (N_2421,N_2313,N_2338);
or U2422 (N_2422,N_2358,N_2291);
nor U2423 (N_2423,N_2266,N_2203);
or U2424 (N_2424,N_2366,N_2200);
and U2425 (N_2425,N_2237,N_2311);
nand U2426 (N_2426,N_2385,N_2397);
or U2427 (N_2427,N_2354,N_2324);
nand U2428 (N_2428,N_2363,N_2320);
nand U2429 (N_2429,N_2253,N_2231);
nand U2430 (N_2430,N_2364,N_2230);
and U2431 (N_2431,N_2225,N_2326);
nand U2432 (N_2432,N_2257,N_2329);
nor U2433 (N_2433,N_2223,N_2342);
nand U2434 (N_2434,N_2299,N_2362);
or U2435 (N_2435,N_2260,N_2377);
or U2436 (N_2436,N_2344,N_2252);
nor U2437 (N_2437,N_2283,N_2279);
or U2438 (N_2438,N_2251,N_2308);
nor U2439 (N_2439,N_2250,N_2278);
or U2440 (N_2440,N_2389,N_2352);
nor U2441 (N_2441,N_2287,N_2360);
nand U2442 (N_2442,N_2296,N_2210);
nor U2443 (N_2443,N_2355,N_2334);
nand U2444 (N_2444,N_2372,N_2346);
and U2445 (N_2445,N_2226,N_2277);
and U2446 (N_2446,N_2236,N_2243);
nand U2447 (N_2447,N_2390,N_2359);
and U2448 (N_2448,N_2292,N_2289);
nand U2449 (N_2449,N_2321,N_2207);
nor U2450 (N_2450,N_2272,N_2327);
nand U2451 (N_2451,N_2258,N_2393);
and U2452 (N_2452,N_2317,N_2399);
nand U2453 (N_2453,N_2337,N_2254);
or U2454 (N_2454,N_2248,N_2235);
nor U2455 (N_2455,N_2336,N_2261);
and U2456 (N_2456,N_2365,N_2218);
or U2457 (N_2457,N_2323,N_2381);
nor U2458 (N_2458,N_2300,N_2383);
nand U2459 (N_2459,N_2263,N_2220);
nor U2460 (N_2460,N_2370,N_2395);
or U2461 (N_2461,N_2348,N_2343);
or U2462 (N_2462,N_2229,N_2304);
xnor U2463 (N_2463,N_2351,N_2265);
nor U2464 (N_2464,N_2332,N_2215);
and U2465 (N_2465,N_2214,N_2371);
or U2466 (N_2466,N_2309,N_2208);
and U2467 (N_2467,N_2295,N_2284);
and U2468 (N_2468,N_2302,N_2228);
nor U2469 (N_2469,N_2310,N_2347);
nor U2470 (N_2470,N_2255,N_2259);
nand U2471 (N_2471,N_2306,N_2357);
and U2472 (N_2472,N_2276,N_2211);
nand U2473 (N_2473,N_2374,N_2298);
nand U2474 (N_2474,N_2368,N_2242);
or U2475 (N_2475,N_2216,N_2398);
nor U2476 (N_2476,N_2328,N_2219);
and U2477 (N_2477,N_2335,N_2238);
nand U2478 (N_2478,N_2361,N_2382);
nor U2479 (N_2479,N_2303,N_2224);
nor U2480 (N_2480,N_2217,N_2209);
nor U2481 (N_2481,N_2339,N_2396);
nor U2482 (N_2482,N_2206,N_2307);
nand U2483 (N_2483,N_2264,N_2246);
and U2484 (N_2484,N_2262,N_2269);
nor U2485 (N_2485,N_2247,N_2305);
nor U2486 (N_2486,N_2267,N_2222);
nor U2487 (N_2487,N_2384,N_2318);
and U2488 (N_2488,N_2391,N_2274);
nand U2489 (N_2489,N_2221,N_2293);
and U2490 (N_2490,N_2301,N_2249);
nand U2491 (N_2491,N_2241,N_2350);
nor U2492 (N_2492,N_2325,N_2204);
nand U2493 (N_2493,N_2244,N_2369);
nand U2494 (N_2494,N_2341,N_2286);
nand U2495 (N_2495,N_2349,N_2227);
or U2496 (N_2496,N_2201,N_2316);
or U2497 (N_2497,N_2319,N_2285);
nor U2498 (N_2498,N_2375,N_2322);
nand U2499 (N_2499,N_2312,N_2315);
or U2500 (N_2500,N_2268,N_2231);
nor U2501 (N_2501,N_2281,N_2272);
nand U2502 (N_2502,N_2281,N_2271);
and U2503 (N_2503,N_2291,N_2351);
nor U2504 (N_2504,N_2393,N_2385);
nand U2505 (N_2505,N_2371,N_2250);
and U2506 (N_2506,N_2337,N_2209);
nand U2507 (N_2507,N_2385,N_2216);
nand U2508 (N_2508,N_2394,N_2235);
nor U2509 (N_2509,N_2390,N_2389);
or U2510 (N_2510,N_2293,N_2286);
and U2511 (N_2511,N_2275,N_2337);
nor U2512 (N_2512,N_2252,N_2357);
nand U2513 (N_2513,N_2367,N_2258);
or U2514 (N_2514,N_2268,N_2272);
or U2515 (N_2515,N_2319,N_2333);
and U2516 (N_2516,N_2290,N_2271);
and U2517 (N_2517,N_2317,N_2286);
xor U2518 (N_2518,N_2235,N_2347);
nand U2519 (N_2519,N_2292,N_2387);
nor U2520 (N_2520,N_2265,N_2336);
or U2521 (N_2521,N_2360,N_2215);
nand U2522 (N_2522,N_2310,N_2298);
nand U2523 (N_2523,N_2320,N_2278);
nor U2524 (N_2524,N_2367,N_2209);
nor U2525 (N_2525,N_2252,N_2251);
or U2526 (N_2526,N_2334,N_2240);
or U2527 (N_2527,N_2351,N_2334);
and U2528 (N_2528,N_2364,N_2334);
nand U2529 (N_2529,N_2248,N_2259);
nand U2530 (N_2530,N_2301,N_2290);
nor U2531 (N_2531,N_2214,N_2304);
or U2532 (N_2532,N_2303,N_2279);
nand U2533 (N_2533,N_2333,N_2231);
and U2534 (N_2534,N_2308,N_2399);
nand U2535 (N_2535,N_2309,N_2246);
and U2536 (N_2536,N_2295,N_2277);
or U2537 (N_2537,N_2243,N_2267);
and U2538 (N_2538,N_2222,N_2302);
nor U2539 (N_2539,N_2244,N_2260);
nand U2540 (N_2540,N_2303,N_2363);
and U2541 (N_2541,N_2359,N_2329);
or U2542 (N_2542,N_2294,N_2335);
or U2543 (N_2543,N_2306,N_2391);
nand U2544 (N_2544,N_2397,N_2263);
nor U2545 (N_2545,N_2262,N_2212);
nor U2546 (N_2546,N_2291,N_2359);
or U2547 (N_2547,N_2248,N_2329);
nor U2548 (N_2548,N_2315,N_2323);
nor U2549 (N_2549,N_2218,N_2374);
xnor U2550 (N_2550,N_2372,N_2289);
nand U2551 (N_2551,N_2319,N_2223);
and U2552 (N_2552,N_2357,N_2249);
nor U2553 (N_2553,N_2339,N_2228);
and U2554 (N_2554,N_2306,N_2292);
and U2555 (N_2555,N_2301,N_2257);
or U2556 (N_2556,N_2385,N_2205);
nor U2557 (N_2557,N_2313,N_2278);
or U2558 (N_2558,N_2330,N_2327);
or U2559 (N_2559,N_2363,N_2210);
and U2560 (N_2560,N_2229,N_2344);
and U2561 (N_2561,N_2260,N_2323);
or U2562 (N_2562,N_2218,N_2303);
and U2563 (N_2563,N_2295,N_2356);
nand U2564 (N_2564,N_2288,N_2265);
and U2565 (N_2565,N_2364,N_2211);
and U2566 (N_2566,N_2289,N_2349);
and U2567 (N_2567,N_2238,N_2250);
nor U2568 (N_2568,N_2239,N_2273);
nand U2569 (N_2569,N_2285,N_2257);
and U2570 (N_2570,N_2329,N_2279);
nand U2571 (N_2571,N_2236,N_2222);
and U2572 (N_2572,N_2286,N_2362);
and U2573 (N_2573,N_2252,N_2388);
and U2574 (N_2574,N_2237,N_2372);
nand U2575 (N_2575,N_2384,N_2220);
or U2576 (N_2576,N_2309,N_2304);
nor U2577 (N_2577,N_2286,N_2375);
and U2578 (N_2578,N_2340,N_2374);
and U2579 (N_2579,N_2376,N_2354);
or U2580 (N_2580,N_2307,N_2296);
or U2581 (N_2581,N_2334,N_2252);
nand U2582 (N_2582,N_2344,N_2203);
or U2583 (N_2583,N_2354,N_2234);
or U2584 (N_2584,N_2228,N_2354);
or U2585 (N_2585,N_2282,N_2331);
nor U2586 (N_2586,N_2256,N_2308);
and U2587 (N_2587,N_2357,N_2205);
nor U2588 (N_2588,N_2377,N_2330);
nor U2589 (N_2589,N_2297,N_2208);
nor U2590 (N_2590,N_2294,N_2297);
nand U2591 (N_2591,N_2281,N_2308);
and U2592 (N_2592,N_2267,N_2335);
or U2593 (N_2593,N_2227,N_2382);
nand U2594 (N_2594,N_2316,N_2252);
nand U2595 (N_2595,N_2311,N_2298);
nand U2596 (N_2596,N_2257,N_2231);
nor U2597 (N_2597,N_2230,N_2368);
nor U2598 (N_2598,N_2254,N_2386);
or U2599 (N_2599,N_2285,N_2396);
or U2600 (N_2600,N_2469,N_2429);
xnor U2601 (N_2601,N_2451,N_2485);
nor U2602 (N_2602,N_2500,N_2521);
or U2603 (N_2603,N_2417,N_2524);
and U2604 (N_2604,N_2413,N_2586);
and U2605 (N_2605,N_2437,N_2520);
nor U2606 (N_2606,N_2438,N_2553);
or U2607 (N_2607,N_2446,N_2545);
or U2608 (N_2608,N_2540,N_2426);
or U2609 (N_2609,N_2472,N_2573);
nand U2610 (N_2610,N_2489,N_2465);
nand U2611 (N_2611,N_2423,N_2562);
nor U2612 (N_2612,N_2499,N_2447);
nand U2613 (N_2613,N_2415,N_2444);
and U2614 (N_2614,N_2463,N_2408);
and U2615 (N_2615,N_2583,N_2512);
and U2616 (N_2616,N_2537,N_2559);
nor U2617 (N_2617,N_2421,N_2486);
nor U2618 (N_2618,N_2536,N_2414);
and U2619 (N_2619,N_2544,N_2502);
and U2620 (N_2620,N_2492,N_2542);
nand U2621 (N_2621,N_2580,N_2576);
nor U2622 (N_2622,N_2584,N_2440);
nand U2623 (N_2623,N_2550,N_2496);
nand U2624 (N_2624,N_2527,N_2443);
or U2625 (N_2625,N_2457,N_2511);
and U2626 (N_2626,N_2557,N_2407);
nor U2627 (N_2627,N_2481,N_2484);
or U2628 (N_2628,N_2452,N_2530);
and U2629 (N_2629,N_2420,N_2442);
nor U2630 (N_2630,N_2497,N_2478);
nor U2631 (N_2631,N_2522,N_2464);
nor U2632 (N_2632,N_2556,N_2582);
nand U2633 (N_2633,N_2532,N_2543);
nor U2634 (N_2634,N_2596,N_2593);
nand U2635 (N_2635,N_2514,N_2506);
and U2636 (N_2636,N_2552,N_2598);
nor U2637 (N_2637,N_2468,N_2475);
nand U2638 (N_2638,N_2498,N_2403);
nor U2639 (N_2639,N_2505,N_2479);
and U2640 (N_2640,N_2528,N_2401);
and U2641 (N_2641,N_2483,N_2435);
or U2642 (N_2642,N_2462,N_2534);
and U2643 (N_2643,N_2461,N_2538);
nor U2644 (N_2644,N_2519,N_2504);
and U2645 (N_2645,N_2513,N_2488);
nor U2646 (N_2646,N_2516,N_2501);
or U2647 (N_2647,N_2529,N_2594);
or U2648 (N_2648,N_2591,N_2546);
and U2649 (N_2649,N_2418,N_2585);
or U2650 (N_2650,N_2419,N_2471);
nor U2651 (N_2651,N_2526,N_2491);
or U2652 (N_2652,N_2445,N_2510);
nand U2653 (N_2653,N_2494,N_2436);
nand U2654 (N_2654,N_2427,N_2433);
nand U2655 (N_2655,N_2455,N_2507);
or U2656 (N_2656,N_2473,N_2493);
or U2657 (N_2657,N_2539,N_2579);
or U2658 (N_2658,N_2571,N_2480);
or U2659 (N_2659,N_2590,N_2595);
and U2660 (N_2660,N_2412,N_2450);
nor U2661 (N_2661,N_2525,N_2533);
and U2662 (N_2662,N_2565,N_2517);
or U2663 (N_2663,N_2569,N_2449);
nor U2664 (N_2664,N_2474,N_2567);
and U2665 (N_2665,N_2575,N_2509);
nor U2666 (N_2666,N_2578,N_2487);
nand U2667 (N_2667,N_2411,N_2570);
and U2668 (N_2668,N_2508,N_2477);
nor U2669 (N_2669,N_2568,N_2476);
nor U2670 (N_2670,N_2541,N_2482);
nor U2671 (N_2671,N_2431,N_2581);
or U2672 (N_2672,N_2410,N_2574);
and U2673 (N_2673,N_2566,N_2535);
and U2674 (N_2674,N_2561,N_2402);
or U2675 (N_2675,N_2422,N_2547);
nand U2676 (N_2676,N_2460,N_2441);
nor U2677 (N_2677,N_2467,N_2563);
and U2678 (N_2678,N_2577,N_2448);
or U2679 (N_2679,N_2503,N_2599);
nor U2680 (N_2680,N_2425,N_2515);
nand U2681 (N_2681,N_2406,N_2554);
nor U2682 (N_2682,N_2466,N_2587);
or U2683 (N_2683,N_2459,N_2430);
nand U2684 (N_2684,N_2405,N_2404);
nor U2685 (N_2685,N_2549,N_2572);
or U2686 (N_2686,N_2490,N_2597);
nor U2687 (N_2687,N_2434,N_2518);
nand U2688 (N_2688,N_2428,N_2439);
nor U2689 (N_2689,N_2453,N_2592);
or U2690 (N_2690,N_2454,N_2564);
nor U2691 (N_2691,N_2424,N_2432);
and U2692 (N_2692,N_2531,N_2560);
or U2693 (N_2693,N_2523,N_2470);
nor U2694 (N_2694,N_2400,N_2495);
and U2695 (N_2695,N_2548,N_2456);
nand U2696 (N_2696,N_2551,N_2416);
nor U2697 (N_2697,N_2589,N_2558);
or U2698 (N_2698,N_2458,N_2555);
nor U2699 (N_2699,N_2588,N_2409);
or U2700 (N_2700,N_2463,N_2574);
or U2701 (N_2701,N_2501,N_2519);
nor U2702 (N_2702,N_2406,N_2411);
and U2703 (N_2703,N_2514,N_2591);
nand U2704 (N_2704,N_2535,N_2522);
or U2705 (N_2705,N_2514,N_2442);
and U2706 (N_2706,N_2503,N_2440);
or U2707 (N_2707,N_2500,N_2446);
nand U2708 (N_2708,N_2537,N_2450);
or U2709 (N_2709,N_2551,N_2495);
or U2710 (N_2710,N_2489,N_2490);
and U2711 (N_2711,N_2582,N_2463);
nand U2712 (N_2712,N_2403,N_2597);
nor U2713 (N_2713,N_2511,N_2585);
or U2714 (N_2714,N_2588,N_2460);
nand U2715 (N_2715,N_2409,N_2519);
or U2716 (N_2716,N_2424,N_2527);
or U2717 (N_2717,N_2524,N_2567);
or U2718 (N_2718,N_2482,N_2585);
and U2719 (N_2719,N_2501,N_2512);
nand U2720 (N_2720,N_2486,N_2498);
and U2721 (N_2721,N_2460,N_2583);
and U2722 (N_2722,N_2544,N_2449);
or U2723 (N_2723,N_2586,N_2590);
and U2724 (N_2724,N_2513,N_2480);
xor U2725 (N_2725,N_2484,N_2460);
nor U2726 (N_2726,N_2407,N_2581);
and U2727 (N_2727,N_2510,N_2423);
and U2728 (N_2728,N_2484,N_2411);
or U2729 (N_2729,N_2583,N_2461);
or U2730 (N_2730,N_2462,N_2584);
and U2731 (N_2731,N_2465,N_2591);
nand U2732 (N_2732,N_2503,N_2566);
nand U2733 (N_2733,N_2464,N_2577);
or U2734 (N_2734,N_2572,N_2423);
nand U2735 (N_2735,N_2586,N_2529);
or U2736 (N_2736,N_2404,N_2485);
nand U2737 (N_2737,N_2502,N_2446);
nand U2738 (N_2738,N_2496,N_2445);
or U2739 (N_2739,N_2552,N_2411);
nor U2740 (N_2740,N_2501,N_2518);
nand U2741 (N_2741,N_2468,N_2585);
and U2742 (N_2742,N_2444,N_2477);
and U2743 (N_2743,N_2483,N_2589);
and U2744 (N_2744,N_2525,N_2425);
and U2745 (N_2745,N_2428,N_2408);
and U2746 (N_2746,N_2476,N_2531);
nor U2747 (N_2747,N_2539,N_2570);
nor U2748 (N_2748,N_2445,N_2448);
and U2749 (N_2749,N_2543,N_2558);
and U2750 (N_2750,N_2520,N_2534);
and U2751 (N_2751,N_2517,N_2567);
and U2752 (N_2752,N_2437,N_2550);
nor U2753 (N_2753,N_2402,N_2422);
and U2754 (N_2754,N_2575,N_2436);
nand U2755 (N_2755,N_2478,N_2470);
nor U2756 (N_2756,N_2417,N_2499);
nand U2757 (N_2757,N_2491,N_2593);
and U2758 (N_2758,N_2523,N_2438);
nand U2759 (N_2759,N_2549,N_2544);
nand U2760 (N_2760,N_2463,N_2430);
nor U2761 (N_2761,N_2408,N_2424);
or U2762 (N_2762,N_2567,N_2461);
or U2763 (N_2763,N_2476,N_2483);
xnor U2764 (N_2764,N_2518,N_2496);
and U2765 (N_2765,N_2401,N_2578);
or U2766 (N_2766,N_2523,N_2578);
nand U2767 (N_2767,N_2448,N_2543);
or U2768 (N_2768,N_2467,N_2535);
and U2769 (N_2769,N_2496,N_2521);
and U2770 (N_2770,N_2515,N_2502);
nand U2771 (N_2771,N_2479,N_2513);
nand U2772 (N_2772,N_2588,N_2563);
and U2773 (N_2773,N_2414,N_2530);
nand U2774 (N_2774,N_2590,N_2506);
and U2775 (N_2775,N_2505,N_2406);
and U2776 (N_2776,N_2597,N_2549);
nand U2777 (N_2777,N_2519,N_2470);
or U2778 (N_2778,N_2556,N_2456);
nand U2779 (N_2779,N_2444,N_2519);
and U2780 (N_2780,N_2573,N_2580);
nor U2781 (N_2781,N_2512,N_2510);
and U2782 (N_2782,N_2405,N_2586);
nor U2783 (N_2783,N_2527,N_2514);
nand U2784 (N_2784,N_2409,N_2500);
nand U2785 (N_2785,N_2447,N_2450);
and U2786 (N_2786,N_2470,N_2417);
nor U2787 (N_2787,N_2475,N_2455);
nand U2788 (N_2788,N_2572,N_2571);
nor U2789 (N_2789,N_2527,N_2432);
nand U2790 (N_2790,N_2581,N_2474);
nand U2791 (N_2791,N_2568,N_2578);
and U2792 (N_2792,N_2567,N_2433);
nor U2793 (N_2793,N_2416,N_2406);
or U2794 (N_2794,N_2458,N_2499);
nor U2795 (N_2795,N_2531,N_2504);
and U2796 (N_2796,N_2512,N_2533);
or U2797 (N_2797,N_2487,N_2488);
and U2798 (N_2798,N_2487,N_2410);
nor U2799 (N_2799,N_2492,N_2582);
nor U2800 (N_2800,N_2749,N_2739);
nor U2801 (N_2801,N_2682,N_2684);
and U2802 (N_2802,N_2723,N_2608);
and U2803 (N_2803,N_2626,N_2797);
nand U2804 (N_2804,N_2664,N_2706);
nand U2805 (N_2805,N_2656,N_2637);
nor U2806 (N_2806,N_2607,N_2777);
and U2807 (N_2807,N_2776,N_2655);
or U2808 (N_2808,N_2719,N_2686);
or U2809 (N_2809,N_2725,N_2649);
nor U2810 (N_2810,N_2622,N_2623);
nor U2811 (N_2811,N_2699,N_2653);
nand U2812 (N_2812,N_2730,N_2736);
or U2813 (N_2813,N_2732,N_2716);
or U2814 (N_2814,N_2687,N_2636);
and U2815 (N_2815,N_2761,N_2691);
and U2816 (N_2816,N_2671,N_2600);
and U2817 (N_2817,N_2644,N_2789);
nor U2818 (N_2818,N_2602,N_2657);
nand U2819 (N_2819,N_2717,N_2680);
nand U2820 (N_2820,N_2605,N_2782);
nor U2821 (N_2821,N_2737,N_2780);
nand U2822 (N_2822,N_2708,N_2721);
nand U2823 (N_2823,N_2648,N_2697);
nand U2824 (N_2824,N_2775,N_2750);
nand U2825 (N_2825,N_2707,N_2766);
nand U2826 (N_2826,N_2698,N_2669);
nand U2827 (N_2827,N_2640,N_2619);
or U2828 (N_2828,N_2615,N_2704);
nor U2829 (N_2829,N_2658,N_2666);
and U2830 (N_2830,N_2773,N_2613);
or U2831 (N_2831,N_2770,N_2692);
and U2832 (N_2832,N_2612,N_2790);
nor U2833 (N_2833,N_2784,N_2753);
nor U2834 (N_2834,N_2792,N_2695);
or U2835 (N_2835,N_2781,N_2620);
and U2836 (N_2836,N_2645,N_2774);
nand U2837 (N_2837,N_2769,N_2763);
nand U2838 (N_2838,N_2743,N_2689);
nand U2839 (N_2839,N_2688,N_2788);
nor U2840 (N_2840,N_2731,N_2651);
and U2841 (N_2841,N_2724,N_2635);
or U2842 (N_2842,N_2764,N_2670);
nor U2843 (N_2843,N_2673,N_2617);
nor U2844 (N_2844,N_2738,N_2614);
nor U2845 (N_2845,N_2601,N_2728);
and U2846 (N_2846,N_2744,N_2633);
nor U2847 (N_2847,N_2634,N_2727);
or U2848 (N_2848,N_2621,N_2778);
or U2849 (N_2849,N_2638,N_2618);
or U2850 (N_2850,N_2734,N_2709);
and U2851 (N_2851,N_2742,N_2604);
nand U2852 (N_2852,N_2747,N_2683);
or U2853 (N_2853,N_2767,N_2696);
nor U2854 (N_2854,N_2668,N_2759);
nor U2855 (N_2855,N_2660,N_2611);
or U2856 (N_2856,N_2745,N_2754);
or U2857 (N_2857,N_2641,N_2720);
nor U2858 (N_2858,N_2722,N_2765);
nand U2859 (N_2859,N_2799,N_2610);
and U2860 (N_2860,N_2755,N_2712);
nor U2861 (N_2861,N_2659,N_2625);
nand U2862 (N_2862,N_2693,N_2629);
or U2863 (N_2863,N_2667,N_2735);
nor U2864 (N_2864,N_2701,N_2795);
nor U2865 (N_2865,N_2787,N_2756);
nand U2866 (N_2866,N_2711,N_2685);
xor U2867 (N_2867,N_2751,N_2733);
nand U2868 (N_2868,N_2681,N_2715);
nand U2869 (N_2869,N_2654,N_2758);
nand U2870 (N_2870,N_2646,N_2741);
nor U2871 (N_2871,N_2603,N_2771);
and U2872 (N_2872,N_2740,N_2647);
nor U2873 (N_2873,N_2752,N_2627);
nor U2874 (N_2874,N_2616,N_2606);
nand U2875 (N_2875,N_2705,N_2665);
nor U2876 (N_2876,N_2710,N_2729);
nand U2877 (N_2877,N_2793,N_2772);
nand U2878 (N_2878,N_2630,N_2703);
and U2879 (N_2879,N_2677,N_2632);
nor U2880 (N_2880,N_2757,N_2713);
nor U2881 (N_2881,N_2639,N_2661);
nor U2882 (N_2882,N_2663,N_2726);
nor U2883 (N_2883,N_2624,N_2662);
nand U2884 (N_2884,N_2643,N_2702);
nor U2885 (N_2885,N_2794,N_2672);
and U2886 (N_2886,N_2714,N_2628);
and U2887 (N_2887,N_2762,N_2748);
and U2888 (N_2888,N_2798,N_2679);
and U2889 (N_2889,N_2690,N_2718);
nand U2890 (N_2890,N_2791,N_2694);
or U2891 (N_2891,N_2768,N_2760);
or U2892 (N_2892,N_2785,N_2650);
or U2893 (N_2893,N_2652,N_2676);
nand U2894 (N_2894,N_2609,N_2746);
nand U2895 (N_2895,N_2796,N_2678);
nand U2896 (N_2896,N_2783,N_2700);
nor U2897 (N_2897,N_2642,N_2631);
nand U2898 (N_2898,N_2786,N_2675);
and U2899 (N_2899,N_2674,N_2779);
nand U2900 (N_2900,N_2617,N_2697);
or U2901 (N_2901,N_2678,N_2746);
nand U2902 (N_2902,N_2679,N_2780);
nand U2903 (N_2903,N_2680,N_2736);
nand U2904 (N_2904,N_2788,N_2603);
or U2905 (N_2905,N_2711,N_2669);
or U2906 (N_2906,N_2792,N_2616);
nor U2907 (N_2907,N_2717,N_2601);
or U2908 (N_2908,N_2759,N_2697);
nand U2909 (N_2909,N_2797,N_2736);
and U2910 (N_2910,N_2740,N_2710);
nor U2911 (N_2911,N_2738,N_2632);
and U2912 (N_2912,N_2683,N_2708);
or U2913 (N_2913,N_2769,N_2771);
nor U2914 (N_2914,N_2729,N_2642);
and U2915 (N_2915,N_2792,N_2624);
and U2916 (N_2916,N_2630,N_2779);
nor U2917 (N_2917,N_2779,N_2750);
and U2918 (N_2918,N_2719,N_2784);
and U2919 (N_2919,N_2610,N_2795);
nand U2920 (N_2920,N_2639,N_2725);
or U2921 (N_2921,N_2665,N_2671);
and U2922 (N_2922,N_2759,N_2640);
nand U2923 (N_2923,N_2612,N_2784);
and U2924 (N_2924,N_2659,N_2669);
and U2925 (N_2925,N_2775,N_2688);
or U2926 (N_2926,N_2604,N_2635);
and U2927 (N_2927,N_2691,N_2789);
nor U2928 (N_2928,N_2791,N_2706);
and U2929 (N_2929,N_2714,N_2738);
nand U2930 (N_2930,N_2763,N_2691);
nand U2931 (N_2931,N_2735,N_2724);
and U2932 (N_2932,N_2680,N_2718);
nor U2933 (N_2933,N_2618,N_2782);
nor U2934 (N_2934,N_2653,N_2661);
or U2935 (N_2935,N_2757,N_2789);
nor U2936 (N_2936,N_2765,N_2697);
and U2937 (N_2937,N_2742,N_2792);
nor U2938 (N_2938,N_2671,N_2656);
and U2939 (N_2939,N_2651,N_2634);
nand U2940 (N_2940,N_2643,N_2731);
nand U2941 (N_2941,N_2762,N_2760);
or U2942 (N_2942,N_2665,N_2687);
nor U2943 (N_2943,N_2795,N_2616);
nand U2944 (N_2944,N_2788,N_2698);
nand U2945 (N_2945,N_2716,N_2775);
or U2946 (N_2946,N_2651,N_2709);
nand U2947 (N_2947,N_2705,N_2775);
nor U2948 (N_2948,N_2796,N_2759);
nand U2949 (N_2949,N_2721,N_2780);
and U2950 (N_2950,N_2721,N_2755);
nand U2951 (N_2951,N_2785,N_2774);
nor U2952 (N_2952,N_2688,N_2718);
nor U2953 (N_2953,N_2733,N_2643);
or U2954 (N_2954,N_2693,N_2758);
xor U2955 (N_2955,N_2798,N_2778);
nand U2956 (N_2956,N_2647,N_2632);
and U2957 (N_2957,N_2675,N_2614);
and U2958 (N_2958,N_2623,N_2633);
or U2959 (N_2959,N_2687,N_2612);
and U2960 (N_2960,N_2752,N_2786);
or U2961 (N_2961,N_2743,N_2605);
or U2962 (N_2962,N_2611,N_2678);
or U2963 (N_2963,N_2616,N_2736);
or U2964 (N_2964,N_2673,N_2611);
and U2965 (N_2965,N_2772,N_2728);
or U2966 (N_2966,N_2683,N_2626);
and U2967 (N_2967,N_2797,N_2727);
and U2968 (N_2968,N_2677,N_2667);
or U2969 (N_2969,N_2730,N_2609);
nand U2970 (N_2970,N_2782,N_2624);
nor U2971 (N_2971,N_2766,N_2748);
or U2972 (N_2972,N_2633,N_2610);
nand U2973 (N_2973,N_2747,N_2607);
nand U2974 (N_2974,N_2783,N_2635);
or U2975 (N_2975,N_2725,N_2728);
nor U2976 (N_2976,N_2765,N_2607);
nand U2977 (N_2977,N_2660,N_2629);
nand U2978 (N_2978,N_2609,N_2721);
or U2979 (N_2979,N_2690,N_2678);
or U2980 (N_2980,N_2688,N_2738);
and U2981 (N_2981,N_2724,N_2636);
nand U2982 (N_2982,N_2657,N_2754);
xnor U2983 (N_2983,N_2742,N_2632);
and U2984 (N_2984,N_2713,N_2614);
nand U2985 (N_2985,N_2655,N_2729);
nor U2986 (N_2986,N_2626,N_2632);
nor U2987 (N_2987,N_2684,N_2707);
nand U2988 (N_2988,N_2760,N_2657);
nand U2989 (N_2989,N_2707,N_2664);
nand U2990 (N_2990,N_2674,N_2786);
or U2991 (N_2991,N_2610,N_2647);
nand U2992 (N_2992,N_2648,N_2644);
or U2993 (N_2993,N_2657,N_2692);
or U2994 (N_2994,N_2638,N_2601);
nand U2995 (N_2995,N_2717,N_2768);
nand U2996 (N_2996,N_2699,N_2763);
or U2997 (N_2997,N_2612,N_2736);
nor U2998 (N_2998,N_2721,N_2762);
or U2999 (N_2999,N_2754,N_2759);
and UO_0 (O_0,N_2808,N_2905);
and UO_1 (O_1,N_2851,N_2814);
and UO_2 (O_2,N_2977,N_2994);
nor UO_3 (O_3,N_2967,N_2913);
or UO_4 (O_4,N_2912,N_2831);
and UO_5 (O_5,N_2926,N_2930);
nor UO_6 (O_6,N_2920,N_2988);
and UO_7 (O_7,N_2815,N_2868);
nor UO_8 (O_8,N_2844,N_2863);
nor UO_9 (O_9,N_2933,N_2874);
and UO_10 (O_10,N_2852,N_2878);
or UO_11 (O_11,N_2879,N_2915);
nor UO_12 (O_12,N_2949,N_2965);
and UO_13 (O_13,N_2973,N_2827);
nand UO_14 (O_14,N_2824,N_2989);
nor UO_15 (O_15,N_2999,N_2821);
and UO_16 (O_16,N_2845,N_2986);
or UO_17 (O_17,N_2961,N_2972);
nand UO_18 (O_18,N_2880,N_2962);
nand UO_19 (O_19,N_2974,N_2960);
or UO_20 (O_20,N_2979,N_2820);
xnor UO_21 (O_21,N_2904,N_2829);
or UO_22 (O_22,N_2876,N_2895);
or UO_23 (O_23,N_2853,N_2883);
nor UO_24 (O_24,N_2801,N_2936);
nand UO_25 (O_25,N_2881,N_2865);
nand UO_26 (O_26,N_2850,N_2871);
nand UO_27 (O_27,N_2980,N_2996);
nor UO_28 (O_28,N_2804,N_2935);
nor UO_29 (O_29,N_2993,N_2860);
nor UO_30 (O_30,N_2810,N_2957);
or UO_31 (O_31,N_2901,N_2998);
nor UO_32 (O_32,N_2898,N_2902);
nor UO_33 (O_33,N_2894,N_2893);
nand UO_34 (O_34,N_2909,N_2976);
nor UO_35 (O_35,N_2832,N_2864);
nor UO_36 (O_36,N_2854,N_2813);
nor UO_37 (O_37,N_2997,N_2855);
or UO_38 (O_38,N_2836,N_2978);
and UO_39 (O_39,N_2983,N_2927);
or UO_40 (O_40,N_2849,N_2959);
nor UO_41 (O_41,N_2981,N_2908);
and UO_42 (O_42,N_2846,N_2803);
or UO_43 (O_43,N_2966,N_2872);
nand UO_44 (O_44,N_2802,N_2985);
and UO_45 (O_45,N_2866,N_2809);
and UO_46 (O_46,N_2800,N_2877);
nand UO_47 (O_47,N_2955,N_2919);
nor UO_48 (O_48,N_2807,N_2910);
and UO_49 (O_49,N_2888,N_2918);
nor UO_50 (O_50,N_2870,N_2843);
nor UO_51 (O_51,N_2968,N_2856);
nand UO_52 (O_52,N_2928,N_2942);
or UO_53 (O_53,N_2964,N_2861);
and UO_54 (O_54,N_2984,N_2817);
nand UO_55 (O_55,N_2995,N_2811);
nor UO_56 (O_56,N_2833,N_2943);
and UO_57 (O_57,N_2929,N_2907);
or UO_58 (O_58,N_2982,N_2916);
and UO_59 (O_59,N_2958,N_2937);
nor UO_60 (O_60,N_2954,N_2873);
or UO_61 (O_61,N_2838,N_2835);
nor UO_62 (O_62,N_2859,N_2896);
and UO_63 (O_63,N_2931,N_2903);
nand UO_64 (O_64,N_2948,N_2897);
nor UO_65 (O_65,N_2946,N_2941);
nor UO_66 (O_66,N_2823,N_2875);
nor UO_67 (O_67,N_2805,N_2858);
and UO_68 (O_68,N_2882,N_2890);
or UO_69 (O_69,N_2924,N_2834);
or UO_70 (O_70,N_2963,N_2947);
nor UO_71 (O_71,N_2837,N_2885);
nor UO_72 (O_72,N_2822,N_2970);
nand UO_73 (O_73,N_2914,N_2940);
nor UO_74 (O_74,N_2825,N_2900);
or UO_75 (O_75,N_2828,N_2847);
or UO_76 (O_76,N_2889,N_2899);
nand UO_77 (O_77,N_2987,N_2840);
and UO_78 (O_78,N_2991,N_2939);
and UO_79 (O_79,N_2922,N_2969);
nand UO_80 (O_80,N_2975,N_2839);
nor UO_81 (O_81,N_2956,N_2819);
and UO_82 (O_82,N_2848,N_2812);
or UO_83 (O_83,N_2869,N_2971);
and UO_84 (O_84,N_2992,N_2892);
and UO_85 (O_85,N_2951,N_2826);
nand UO_86 (O_86,N_2816,N_2806);
nand UO_87 (O_87,N_2953,N_2944);
and UO_88 (O_88,N_2917,N_2932);
nand UO_89 (O_89,N_2842,N_2818);
nand UO_90 (O_90,N_2945,N_2934);
and UO_91 (O_91,N_2911,N_2990);
and UO_92 (O_92,N_2867,N_2921);
and UO_93 (O_93,N_2906,N_2841);
nor UO_94 (O_94,N_2862,N_2952);
or UO_95 (O_95,N_2884,N_2925);
and UO_96 (O_96,N_2891,N_2938);
and UO_97 (O_97,N_2886,N_2830);
nor UO_98 (O_98,N_2857,N_2950);
or UO_99 (O_99,N_2887,N_2923);
nand UO_100 (O_100,N_2953,N_2931);
nor UO_101 (O_101,N_2881,N_2845);
nor UO_102 (O_102,N_2949,N_2886);
and UO_103 (O_103,N_2813,N_2900);
nor UO_104 (O_104,N_2925,N_2990);
and UO_105 (O_105,N_2972,N_2807);
nor UO_106 (O_106,N_2894,N_2852);
nand UO_107 (O_107,N_2814,N_2885);
nand UO_108 (O_108,N_2989,N_2993);
nor UO_109 (O_109,N_2980,N_2849);
or UO_110 (O_110,N_2991,N_2883);
and UO_111 (O_111,N_2826,N_2891);
or UO_112 (O_112,N_2827,N_2901);
or UO_113 (O_113,N_2900,N_2800);
and UO_114 (O_114,N_2986,N_2979);
and UO_115 (O_115,N_2837,N_2886);
or UO_116 (O_116,N_2815,N_2844);
xor UO_117 (O_117,N_2894,N_2995);
or UO_118 (O_118,N_2930,N_2911);
and UO_119 (O_119,N_2855,N_2853);
or UO_120 (O_120,N_2940,N_2991);
nand UO_121 (O_121,N_2858,N_2997);
and UO_122 (O_122,N_2874,N_2870);
nor UO_123 (O_123,N_2832,N_2943);
or UO_124 (O_124,N_2996,N_2821);
and UO_125 (O_125,N_2934,N_2825);
nand UO_126 (O_126,N_2896,N_2805);
nand UO_127 (O_127,N_2887,N_2984);
or UO_128 (O_128,N_2829,N_2922);
nand UO_129 (O_129,N_2954,N_2959);
or UO_130 (O_130,N_2944,N_2971);
and UO_131 (O_131,N_2980,N_2884);
or UO_132 (O_132,N_2975,N_2876);
or UO_133 (O_133,N_2830,N_2838);
or UO_134 (O_134,N_2977,N_2904);
and UO_135 (O_135,N_2893,N_2907);
and UO_136 (O_136,N_2809,N_2849);
or UO_137 (O_137,N_2878,N_2904);
nand UO_138 (O_138,N_2895,N_2901);
and UO_139 (O_139,N_2884,N_2984);
nor UO_140 (O_140,N_2926,N_2830);
nand UO_141 (O_141,N_2937,N_2836);
nor UO_142 (O_142,N_2832,N_2835);
nor UO_143 (O_143,N_2936,N_2964);
nand UO_144 (O_144,N_2891,N_2852);
nor UO_145 (O_145,N_2926,N_2834);
nand UO_146 (O_146,N_2876,N_2918);
nor UO_147 (O_147,N_2803,N_2937);
nand UO_148 (O_148,N_2807,N_2854);
or UO_149 (O_149,N_2944,N_2957);
or UO_150 (O_150,N_2926,N_2873);
or UO_151 (O_151,N_2980,N_2871);
nand UO_152 (O_152,N_2995,N_2850);
xor UO_153 (O_153,N_2958,N_2947);
and UO_154 (O_154,N_2829,N_2944);
or UO_155 (O_155,N_2843,N_2939);
or UO_156 (O_156,N_2865,N_2880);
and UO_157 (O_157,N_2912,N_2903);
and UO_158 (O_158,N_2928,N_2829);
nand UO_159 (O_159,N_2881,N_2823);
and UO_160 (O_160,N_2971,N_2863);
or UO_161 (O_161,N_2879,N_2917);
and UO_162 (O_162,N_2979,N_2983);
nor UO_163 (O_163,N_2806,N_2804);
xnor UO_164 (O_164,N_2841,N_2920);
and UO_165 (O_165,N_2840,N_2866);
or UO_166 (O_166,N_2949,N_2879);
nor UO_167 (O_167,N_2858,N_2848);
nand UO_168 (O_168,N_2816,N_2992);
and UO_169 (O_169,N_2980,N_2813);
and UO_170 (O_170,N_2898,N_2823);
nor UO_171 (O_171,N_2823,N_2931);
and UO_172 (O_172,N_2876,N_2957);
and UO_173 (O_173,N_2968,N_2991);
nor UO_174 (O_174,N_2896,N_2837);
and UO_175 (O_175,N_2825,N_2929);
nor UO_176 (O_176,N_2949,N_2889);
and UO_177 (O_177,N_2985,N_2865);
nand UO_178 (O_178,N_2828,N_2852);
and UO_179 (O_179,N_2963,N_2852);
or UO_180 (O_180,N_2980,N_2976);
or UO_181 (O_181,N_2923,N_2800);
or UO_182 (O_182,N_2896,N_2845);
or UO_183 (O_183,N_2954,N_2864);
or UO_184 (O_184,N_2979,N_2877);
nand UO_185 (O_185,N_2953,N_2913);
and UO_186 (O_186,N_2837,N_2816);
nor UO_187 (O_187,N_2964,N_2925);
nor UO_188 (O_188,N_2804,N_2899);
or UO_189 (O_189,N_2849,N_2986);
and UO_190 (O_190,N_2981,N_2828);
or UO_191 (O_191,N_2802,N_2986);
nand UO_192 (O_192,N_2984,N_2804);
nor UO_193 (O_193,N_2829,N_2964);
nor UO_194 (O_194,N_2867,N_2923);
nor UO_195 (O_195,N_2891,N_2868);
nand UO_196 (O_196,N_2882,N_2936);
or UO_197 (O_197,N_2917,N_2908);
or UO_198 (O_198,N_2980,N_2915);
nand UO_199 (O_199,N_2904,N_2935);
and UO_200 (O_200,N_2978,N_2905);
and UO_201 (O_201,N_2862,N_2826);
or UO_202 (O_202,N_2829,N_2955);
or UO_203 (O_203,N_2880,N_2983);
nor UO_204 (O_204,N_2998,N_2896);
or UO_205 (O_205,N_2838,N_2854);
nand UO_206 (O_206,N_2964,N_2815);
or UO_207 (O_207,N_2989,N_2849);
or UO_208 (O_208,N_2969,N_2975);
and UO_209 (O_209,N_2860,N_2867);
or UO_210 (O_210,N_2875,N_2879);
nand UO_211 (O_211,N_2936,N_2982);
or UO_212 (O_212,N_2974,N_2804);
or UO_213 (O_213,N_2828,N_2999);
and UO_214 (O_214,N_2840,N_2844);
or UO_215 (O_215,N_2875,N_2800);
and UO_216 (O_216,N_2806,N_2867);
or UO_217 (O_217,N_2879,N_2931);
nor UO_218 (O_218,N_2927,N_2857);
nand UO_219 (O_219,N_2972,N_2999);
or UO_220 (O_220,N_2847,N_2881);
nand UO_221 (O_221,N_2898,N_2950);
and UO_222 (O_222,N_2928,N_2981);
nand UO_223 (O_223,N_2875,N_2935);
and UO_224 (O_224,N_2973,N_2943);
nor UO_225 (O_225,N_2806,N_2885);
nor UO_226 (O_226,N_2875,N_2822);
nand UO_227 (O_227,N_2979,N_2856);
nand UO_228 (O_228,N_2918,N_2966);
nand UO_229 (O_229,N_2865,N_2964);
or UO_230 (O_230,N_2972,N_2825);
or UO_231 (O_231,N_2857,N_2889);
and UO_232 (O_232,N_2943,N_2931);
or UO_233 (O_233,N_2936,N_2989);
and UO_234 (O_234,N_2971,N_2928);
nand UO_235 (O_235,N_2985,N_2903);
or UO_236 (O_236,N_2835,N_2840);
or UO_237 (O_237,N_2947,N_2849);
and UO_238 (O_238,N_2932,N_2827);
nor UO_239 (O_239,N_2979,N_2868);
nor UO_240 (O_240,N_2873,N_2916);
nor UO_241 (O_241,N_2872,N_2861);
nand UO_242 (O_242,N_2933,N_2879);
and UO_243 (O_243,N_2871,N_2975);
nand UO_244 (O_244,N_2853,N_2968);
or UO_245 (O_245,N_2825,N_2928);
nand UO_246 (O_246,N_2992,N_2991);
nor UO_247 (O_247,N_2988,N_2828);
and UO_248 (O_248,N_2923,N_2929);
or UO_249 (O_249,N_2906,N_2944);
nor UO_250 (O_250,N_2800,N_2861);
or UO_251 (O_251,N_2883,N_2913);
nand UO_252 (O_252,N_2923,N_2807);
nand UO_253 (O_253,N_2856,N_2978);
or UO_254 (O_254,N_2885,N_2907);
or UO_255 (O_255,N_2834,N_2802);
nand UO_256 (O_256,N_2879,N_2828);
or UO_257 (O_257,N_2986,N_2815);
xor UO_258 (O_258,N_2826,N_2972);
nor UO_259 (O_259,N_2912,N_2890);
or UO_260 (O_260,N_2888,N_2948);
or UO_261 (O_261,N_2996,N_2981);
nand UO_262 (O_262,N_2902,N_2831);
nand UO_263 (O_263,N_2916,N_2953);
nand UO_264 (O_264,N_2984,N_2823);
and UO_265 (O_265,N_2871,N_2954);
and UO_266 (O_266,N_2960,N_2838);
nor UO_267 (O_267,N_2968,N_2938);
nor UO_268 (O_268,N_2924,N_2858);
nand UO_269 (O_269,N_2975,N_2919);
nand UO_270 (O_270,N_2852,N_2809);
nand UO_271 (O_271,N_2984,N_2903);
nor UO_272 (O_272,N_2899,N_2949);
nor UO_273 (O_273,N_2935,N_2829);
or UO_274 (O_274,N_2951,N_2942);
nand UO_275 (O_275,N_2974,N_2854);
or UO_276 (O_276,N_2809,N_2915);
nor UO_277 (O_277,N_2898,N_2907);
nor UO_278 (O_278,N_2855,N_2980);
nand UO_279 (O_279,N_2922,N_2877);
nor UO_280 (O_280,N_2847,N_2867);
nor UO_281 (O_281,N_2921,N_2989);
nand UO_282 (O_282,N_2887,N_2895);
and UO_283 (O_283,N_2894,N_2816);
nor UO_284 (O_284,N_2969,N_2963);
or UO_285 (O_285,N_2986,N_2891);
and UO_286 (O_286,N_2856,N_2883);
nand UO_287 (O_287,N_2933,N_2892);
and UO_288 (O_288,N_2964,N_2923);
and UO_289 (O_289,N_2802,N_2987);
xor UO_290 (O_290,N_2940,N_2859);
xor UO_291 (O_291,N_2871,N_2804);
and UO_292 (O_292,N_2838,N_2915);
and UO_293 (O_293,N_2881,N_2935);
and UO_294 (O_294,N_2972,N_2833);
or UO_295 (O_295,N_2895,N_2836);
or UO_296 (O_296,N_2816,N_2927);
or UO_297 (O_297,N_2826,N_2901);
and UO_298 (O_298,N_2983,N_2913);
or UO_299 (O_299,N_2811,N_2955);
nor UO_300 (O_300,N_2934,N_2859);
nand UO_301 (O_301,N_2862,N_2944);
nor UO_302 (O_302,N_2963,N_2872);
nor UO_303 (O_303,N_2808,N_2838);
xor UO_304 (O_304,N_2943,N_2997);
xor UO_305 (O_305,N_2997,N_2814);
or UO_306 (O_306,N_2851,N_2857);
nor UO_307 (O_307,N_2930,N_2895);
nand UO_308 (O_308,N_2878,N_2818);
nand UO_309 (O_309,N_2847,N_2837);
and UO_310 (O_310,N_2990,N_2834);
nor UO_311 (O_311,N_2800,N_2899);
nand UO_312 (O_312,N_2971,N_2978);
nand UO_313 (O_313,N_2842,N_2954);
nor UO_314 (O_314,N_2829,N_2914);
and UO_315 (O_315,N_2843,N_2829);
nor UO_316 (O_316,N_2854,N_2852);
or UO_317 (O_317,N_2903,N_2983);
nor UO_318 (O_318,N_2922,N_2903);
or UO_319 (O_319,N_2904,N_2917);
nand UO_320 (O_320,N_2970,N_2847);
nand UO_321 (O_321,N_2860,N_2937);
nand UO_322 (O_322,N_2898,N_2975);
nand UO_323 (O_323,N_2819,N_2890);
nor UO_324 (O_324,N_2834,N_2910);
and UO_325 (O_325,N_2895,N_2890);
nor UO_326 (O_326,N_2858,N_2857);
nor UO_327 (O_327,N_2849,N_2914);
nor UO_328 (O_328,N_2895,N_2988);
nor UO_329 (O_329,N_2860,N_2966);
nor UO_330 (O_330,N_2819,N_2904);
nor UO_331 (O_331,N_2811,N_2932);
nand UO_332 (O_332,N_2836,N_2889);
or UO_333 (O_333,N_2839,N_2843);
or UO_334 (O_334,N_2991,N_2936);
and UO_335 (O_335,N_2947,N_2866);
nor UO_336 (O_336,N_2814,N_2812);
or UO_337 (O_337,N_2808,N_2971);
nand UO_338 (O_338,N_2903,N_2989);
and UO_339 (O_339,N_2952,N_2867);
nor UO_340 (O_340,N_2950,N_2933);
nor UO_341 (O_341,N_2894,N_2880);
or UO_342 (O_342,N_2966,N_2848);
or UO_343 (O_343,N_2819,N_2929);
nor UO_344 (O_344,N_2922,N_2952);
nor UO_345 (O_345,N_2880,N_2873);
nor UO_346 (O_346,N_2962,N_2930);
and UO_347 (O_347,N_2888,N_2983);
and UO_348 (O_348,N_2944,N_2895);
nor UO_349 (O_349,N_2971,N_2861);
nand UO_350 (O_350,N_2917,N_2871);
and UO_351 (O_351,N_2995,N_2910);
and UO_352 (O_352,N_2880,N_2847);
nor UO_353 (O_353,N_2927,N_2884);
nand UO_354 (O_354,N_2986,N_2865);
and UO_355 (O_355,N_2847,N_2815);
nor UO_356 (O_356,N_2823,N_2810);
nand UO_357 (O_357,N_2866,N_2894);
and UO_358 (O_358,N_2913,N_2985);
nor UO_359 (O_359,N_2978,N_2842);
nor UO_360 (O_360,N_2940,N_2994);
nor UO_361 (O_361,N_2900,N_2898);
or UO_362 (O_362,N_2848,N_2999);
nor UO_363 (O_363,N_2949,N_2874);
nand UO_364 (O_364,N_2851,N_2930);
and UO_365 (O_365,N_2915,N_2857);
and UO_366 (O_366,N_2976,N_2816);
nor UO_367 (O_367,N_2826,N_2946);
or UO_368 (O_368,N_2979,N_2872);
nor UO_369 (O_369,N_2965,N_2916);
nand UO_370 (O_370,N_2826,N_2809);
nand UO_371 (O_371,N_2980,N_2893);
xnor UO_372 (O_372,N_2990,N_2956);
and UO_373 (O_373,N_2835,N_2897);
or UO_374 (O_374,N_2883,N_2843);
or UO_375 (O_375,N_2963,N_2871);
nor UO_376 (O_376,N_2803,N_2901);
nor UO_377 (O_377,N_2855,N_2934);
nand UO_378 (O_378,N_2937,N_2955);
or UO_379 (O_379,N_2953,N_2992);
nand UO_380 (O_380,N_2899,N_2809);
or UO_381 (O_381,N_2928,N_2992);
and UO_382 (O_382,N_2940,N_2867);
and UO_383 (O_383,N_2990,N_2902);
xnor UO_384 (O_384,N_2981,N_2816);
or UO_385 (O_385,N_2936,N_2984);
nand UO_386 (O_386,N_2820,N_2899);
nor UO_387 (O_387,N_2905,N_2907);
nor UO_388 (O_388,N_2917,N_2996);
and UO_389 (O_389,N_2865,N_2949);
nor UO_390 (O_390,N_2994,N_2858);
nand UO_391 (O_391,N_2894,N_2862);
or UO_392 (O_392,N_2868,N_2841);
or UO_393 (O_393,N_2953,N_2833);
nand UO_394 (O_394,N_2829,N_2996);
and UO_395 (O_395,N_2879,N_2808);
nor UO_396 (O_396,N_2995,N_2975);
and UO_397 (O_397,N_2962,N_2903);
xor UO_398 (O_398,N_2859,N_2947);
or UO_399 (O_399,N_2823,N_2971);
nor UO_400 (O_400,N_2809,N_2964);
or UO_401 (O_401,N_2889,N_2877);
nand UO_402 (O_402,N_2965,N_2944);
xor UO_403 (O_403,N_2908,N_2817);
and UO_404 (O_404,N_2957,N_2835);
nor UO_405 (O_405,N_2962,N_2840);
nor UO_406 (O_406,N_2917,N_2863);
nand UO_407 (O_407,N_2984,N_2945);
or UO_408 (O_408,N_2852,N_2945);
or UO_409 (O_409,N_2823,N_2960);
nand UO_410 (O_410,N_2872,N_2923);
and UO_411 (O_411,N_2914,N_2873);
nand UO_412 (O_412,N_2878,N_2879);
nor UO_413 (O_413,N_2870,N_2908);
nand UO_414 (O_414,N_2965,N_2863);
nor UO_415 (O_415,N_2826,N_2817);
nor UO_416 (O_416,N_2893,N_2966);
nor UO_417 (O_417,N_2838,N_2911);
or UO_418 (O_418,N_2802,N_2977);
or UO_419 (O_419,N_2839,N_2848);
or UO_420 (O_420,N_2878,N_2918);
nor UO_421 (O_421,N_2879,N_2840);
and UO_422 (O_422,N_2877,N_2996);
nor UO_423 (O_423,N_2927,N_2863);
or UO_424 (O_424,N_2949,N_2853);
or UO_425 (O_425,N_2865,N_2898);
nand UO_426 (O_426,N_2932,N_2899);
nand UO_427 (O_427,N_2851,N_2945);
or UO_428 (O_428,N_2874,N_2914);
nand UO_429 (O_429,N_2873,N_2805);
nand UO_430 (O_430,N_2919,N_2986);
and UO_431 (O_431,N_2863,N_2872);
and UO_432 (O_432,N_2813,N_2921);
nor UO_433 (O_433,N_2868,N_2884);
xor UO_434 (O_434,N_2810,N_2885);
nor UO_435 (O_435,N_2986,N_2951);
or UO_436 (O_436,N_2827,N_2885);
nor UO_437 (O_437,N_2898,N_2960);
nand UO_438 (O_438,N_2982,N_2942);
and UO_439 (O_439,N_2943,N_2927);
and UO_440 (O_440,N_2937,N_2816);
and UO_441 (O_441,N_2981,N_2954);
or UO_442 (O_442,N_2995,N_2809);
and UO_443 (O_443,N_2962,N_2995);
or UO_444 (O_444,N_2871,N_2806);
nand UO_445 (O_445,N_2889,N_2825);
or UO_446 (O_446,N_2836,N_2998);
nand UO_447 (O_447,N_2977,N_2852);
and UO_448 (O_448,N_2984,N_2886);
or UO_449 (O_449,N_2924,N_2891);
nor UO_450 (O_450,N_2985,N_2984);
or UO_451 (O_451,N_2914,N_2977);
nand UO_452 (O_452,N_2826,N_2914);
nand UO_453 (O_453,N_2942,N_2989);
and UO_454 (O_454,N_2955,N_2872);
and UO_455 (O_455,N_2950,N_2801);
xnor UO_456 (O_456,N_2906,N_2879);
and UO_457 (O_457,N_2951,N_2975);
nor UO_458 (O_458,N_2906,N_2959);
and UO_459 (O_459,N_2984,N_2980);
nand UO_460 (O_460,N_2866,N_2887);
or UO_461 (O_461,N_2930,N_2858);
nor UO_462 (O_462,N_2870,N_2994);
and UO_463 (O_463,N_2969,N_2925);
nor UO_464 (O_464,N_2900,N_2816);
nand UO_465 (O_465,N_2949,N_2877);
nor UO_466 (O_466,N_2960,N_2808);
or UO_467 (O_467,N_2818,N_2997);
or UO_468 (O_468,N_2957,N_2967);
nand UO_469 (O_469,N_2884,N_2974);
nand UO_470 (O_470,N_2992,N_2861);
nand UO_471 (O_471,N_2966,N_2853);
nor UO_472 (O_472,N_2874,N_2905);
or UO_473 (O_473,N_2845,N_2908);
nand UO_474 (O_474,N_2964,N_2853);
or UO_475 (O_475,N_2852,N_2803);
nor UO_476 (O_476,N_2955,N_2901);
and UO_477 (O_477,N_2850,N_2825);
nor UO_478 (O_478,N_2833,N_2867);
nor UO_479 (O_479,N_2944,N_2922);
nor UO_480 (O_480,N_2962,N_2952);
nand UO_481 (O_481,N_2814,N_2910);
nor UO_482 (O_482,N_2992,N_2825);
nand UO_483 (O_483,N_2978,N_2923);
and UO_484 (O_484,N_2919,N_2855);
nor UO_485 (O_485,N_2866,N_2843);
and UO_486 (O_486,N_2952,N_2979);
and UO_487 (O_487,N_2828,N_2809);
nor UO_488 (O_488,N_2838,N_2906);
and UO_489 (O_489,N_2877,N_2909);
nor UO_490 (O_490,N_2840,N_2982);
and UO_491 (O_491,N_2897,N_2900);
and UO_492 (O_492,N_2811,N_2914);
nand UO_493 (O_493,N_2921,N_2885);
and UO_494 (O_494,N_2887,N_2810);
nor UO_495 (O_495,N_2987,N_2950);
and UO_496 (O_496,N_2971,N_2854);
nor UO_497 (O_497,N_2991,N_2872);
and UO_498 (O_498,N_2911,N_2801);
nor UO_499 (O_499,N_2840,N_2875);
endmodule