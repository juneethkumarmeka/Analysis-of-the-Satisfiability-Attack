module basic_1000_10000_1500_4_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_697,In_390);
nand U1 (N_1,In_475,In_889);
or U2 (N_2,In_853,In_454);
nor U3 (N_3,In_716,In_20);
nor U4 (N_4,In_494,In_649);
or U5 (N_5,In_94,In_804);
nand U6 (N_6,In_336,In_451);
nand U7 (N_7,In_112,In_995);
and U8 (N_8,In_898,In_386);
nand U9 (N_9,In_815,In_295);
nand U10 (N_10,In_514,In_849);
or U11 (N_11,In_724,In_512);
and U12 (N_12,In_675,In_587);
nand U13 (N_13,In_405,In_571);
nor U14 (N_14,In_49,In_518);
and U15 (N_15,In_755,In_281);
or U16 (N_16,In_642,In_600);
nor U17 (N_17,In_994,In_318);
or U18 (N_18,In_51,In_958);
or U19 (N_19,In_355,In_733);
or U20 (N_20,In_694,In_291);
or U21 (N_21,In_315,In_781);
nand U22 (N_22,In_420,In_885);
and U23 (N_23,In_776,In_822);
nor U24 (N_24,In_303,In_188);
and U25 (N_25,In_865,In_610);
nor U26 (N_26,In_184,In_113);
nand U27 (N_27,In_81,In_984);
and U28 (N_28,In_554,In_828);
and U29 (N_29,In_75,In_977);
or U30 (N_30,In_799,In_873);
or U31 (N_31,In_695,In_578);
nand U32 (N_32,In_952,In_147);
and U33 (N_33,In_786,In_686);
nand U34 (N_34,In_125,In_845);
nor U35 (N_35,In_167,In_68);
nand U36 (N_36,In_640,In_831);
and U37 (N_37,In_987,In_537);
nor U38 (N_38,In_955,In_961);
or U39 (N_39,In_651,In_878);
nand U40 (N_40,In_161,In_641);
nand U41 (N_41,In_489,In_748);
and U42 (N_42,In_637,In_462);
or U43 (N_43,In_389,In_121);
and U44 (N_44,In_586,In_784);
nand U45 (N_45,In_403,In_509);
nor U46 (N_46,In_198,In_399);
nor U47 (N_47,In_194,In_939);
nand U48 (N_48,In_813,In_193);
nor U49 (N_49,In_567,In_681);
nand U50 (N_50,In_553,In_42);
nand U51 (N_51,In_319,In_38);
nor U52 (N_52,In_169,In_983);
and U53 (N_53,In_674,In_759);
and U54 (N_54,In_360,In_338);
nor U55 (N_55,In_954,In_372);
or U56 (N_56,In_215,In_385);
nor U57 (N_57,In_887,In_304);
or U58 (N_58,In_912,In_682);
and U59 (N_59,In_497,In_325);
nand U60 (N_60,In_673,In_635);
nand U61 (N_61,In_902,In_397);
and U62 (N_62,In_840,In_923);
or U63 (N_63,In_52,In_988);
nor U64 (N_64,In_422,In_615);
nand U65 (N_65,In_79,In_36);
nor U66 (N_66,In_880,In_190);
nand U67 (N_67,In_572,In_827);
and U68 (N_68,In_82,In_23);
nor U69 (N_69,In_408,In_8);
nand U70 (N_70,In_86,In_608);
nor U71 (N_71,In_914,In_824);
and U72 (N_72,In_529,In_505);
nor U73 (N_73,In_848,In_138);
and U74 (N_74,In_585,In_140);
nand U75 (N_75,In_783,In_279);
nand U76 (N_76,In_78,In_407);
or U77 (N_77,In_219,In_974);
nor U78 (N_78,In_807,In_469);
and U79 (N_79,In_387,In_523);
or U80 (N_80,In_237,In_119);
or U81 (N_81,In_285,In_738);
nand U82 (N_82,In_91,In_750);
nand U83 (N_83,In_897,In_569);
nand U84 (N_84,In_270,In_671);
or U85 (N_85,In_267,In_177);
and U86 (N_86,In_660,In_966);
xor U87 (N_87,In_526,In_524);
or U88 (N_88,In_468,In_691);
or U89 (N_89,In_756,In_427);
or U90 (N_90,In_61,In_588);
or U91 (N_91,In_752,In_260);
or U92 (N_92,In_749,In_255);
nor U93 (N_93,In_111,In_525);
nand U94 (N_94,In_609,In_120);
or U95 (N_95,In_820,In_570);
nor U96 (N_96,In_143,In_678);
nor U97 (N_97,In_591,In_593);
nor U98 (N_98,In_409,In_13);
nand U99 (N_99,In_904,In_737);
and U100 (N_100,In_398,In_705);
or U101 (N_101,In_344,In_657);
nand U102 (N_102,In_234,In_973);
xnor U103 (N_103,In_688,In_178);
or U104 (N_104,In_266,In_991);
or U105 (N_105,In_577,In_362);
or U106 (N_106,In_661,In_174);
or U107 (N_107,In_544,In_400);
or U108 (N_108,In_683,In_861);
nor U109 (N_109,In_645,In_32);
or U110 (N_110,In_773,In_156);
or U111 (N_111,In_877,In_780);
nand U112 (N_112,In_11,In_937);
and U113 (N_113,In_88,In_47);
nor U114 (N_114,In_40,In_4);
nor U115 (N_115,In_208,In_223);
or U116 (N_116,In_248,In_351);
nand U117 (N_117,In_7,In_298);
nor U118 (N_118,In_731,In_864);
nor U119 (N_119,In_732,In_742);
nor U120 (N_120,In_986,In_720);
or U121 (N_121,In_154,In_703);
nand U122 (N_122,In_187,In_626);
nor U123 (N_123,In_765,In_150);
or U124 (N_124,In_825,In_37);
nand U125 (N_125,In_485,In_6);
nand U126 (N_126,In_690,In_216);
nor U127 (N_127,In_774,In_445);
nand U128 (N_128,In_448,In_630);
and U129 (N_129,In_806,In_361);
or U130 (N_130,In_998,In_348);
nand U131 (N_131,In_483,In_496);
and U132 (N_132,In_54,In_614);
and U133 (N_133,In_264,In_166);
nor U134 (N_134,In_596,In_326);
nor U135 (N_135,In_711,In_391);
or U136 (N_136,In_132,In_313);
nand U137 (N_137,In_796,In_200);
nand U138 (N_138,In_943,In_808);
or U139 (N_139,In_253,In_627);
or U140 (N_140,In_417,In_838);
nor U141 (N_141,In_35,In_57);
and U142 (N_142,In_706,In_792);
nand U143 (N_143,In_490,In_459);
and U144 (N_144,In_250,In_746);
and U145 (N_145,In_339,In_564);
or U146 (N_146,In_975,In_863);
or U147 (N_147,In_242,In_340);
or U148 (N_148,In_947,In_666);
nor U149 (N_149,In_527,In_624);
or U150 (N_150,In_379,In_546);
and U151 (N_151,In_548,In_352);
nand U152 (N_152,In_41,In_214);
or U153 (N_153,In_830,In_498);
nor U154 (N_154,In_979,In_927);
nand U155 (N_155,In_823,In_21);
and U156 (N_156,In_382,In_282);
nor U157 (N_157,In_718,In_740);
nand U158 (N_158,In_443,In_16);
nand U159 (N_159,In_413,In_918);
and U160 (N_160,In_894,In_693);
nor U161 (N_161,In_369,In_655);
or U162 (N_162,In_753,In_185);
and U163 (N_163,In_930,In_758);
nor U164 (N_164,In_932,In_10);
or U165 (N_165,In_231,In_402);
or U166 (N_166,In_180,In_327);
nor U167 (N_167,In_476,In_871);
nor U168 (N_168,In_990,In_109);
and U169 (N_169,In_946,In_106);
nor U170 (N_170,In_87,In_757);
and U171 (N_171,In_296,In_31);
or U172 (N_172,In_829,In_648);
and U173 (N_173,In_719,In_258);
nor U174 (N_174,In_633,In_371);
nor U175 (N_175,In_359,In_510);
nor U176 (N_176,In_891,In_333);
and U177 (N_177,In_1,In_832);
nand U178 (N_178,In_936,In_560);
nand U179 (N_179,In_760,In_522);
and U180 (N_180,In_713,In_816);
or U181 (N_181,In_658,In_805);
nand U182 (N_182,In_934,In_652);
and U183 (N_183,In_613,In_884);
nor U184 (N_184,In_317,In_71);
and U185 (N_185,In_584,In_687);
nor U186 (N_186,In_676,In_201);
and U187 (N_187,In_426,In_725);
nor U188 (N_188,In_739,In_115);
and U189 (N_189,In_2,In_501);
and U190 (N_190,In_364,In_328);
nor U191 (N_191,In_558,In_899);
and U192 (N_192,In_941,In_775);
or U193 (N_193,In_911,In_539);
and U194 (N_194,In_940,In_704);
xnor U195 (N_195,In_274,In_965);
and U196 (N_196,In_90,In_908);
nor U197 (N_197,In_346,In_769);
nor U198 (N_198,In_436,In_684);
xnor U199 (N_199,In_305,In_948);
nor U200 (N_200,In_680,In_888);
nand U201 (N_201,In_347,In_243);
nand U202 (N_202,In_25,In_528);
nand U203 (N_203,In_284,In_472);
nor U204 (N_204,In_971,In_331);
nand U205 (N_205,In_481,In_730);
nor U206 (N_206,In_559,In_550);
nor U207 (N_207,In_341,In_104);
and U208 (N_208,In_579,In_129);
nand U209 (N_209,In_394,In_920);
nor U210 (N_210,In_962,In_165);
nor U211 (N_211,In_314,In_826);
and U212 (N_212,In_404,In_24);
nand U213 (N_213,In_771,In_100);
nand U214 (N_214,In_181,In_310);
or U215 (N_215,In_375,In_43);
nand U216 (N_216,In_870,In_502);
nor U217 (N_217,In_557,In_477);
and U218 (N_218,In_556,In_337);
nor U219 (N_219,In_65,In_798);
nand U220 (N_220,In_513,In_460);
or U221 (N_221,In_874,In_197);
and U222 (N_222,In_886,In_667);
or U223 (N_223,In_97,In_745);
nor U224 (N_224,In_601,In_555);
and U225 (N_225,In_329,In_220);
or U226 (N_226,In_101,In_883);
nor U227 (N_227,In_967,In_280);
nor U228 (N_228,In_721,In_449);
nor U229 (N_229,In_72,In_142);
and U230 (N_230,In_392,In_493);
and U231 (N_231,In_441,In_935);
or U232 (N_232,In_159,In_532);
nor U233 (N_233,In_412,In_334);
and U234 (N_234,In_672,In_98);
nand U235 (N_235,In_252,In_698);
nor U236 (N_236,In_604,In_599);
or U237 (N_237,In_15,In_903);
and U238 (N_238,In_980,In_707);
nand U239 (N_239,In_70,In_989);
nand U240 (N_240,In_793,In_136);
and U241 (N_241,In_450,In_900);
nand U242 (N_242,In_452,In_530);
nor U243 (N_243,In_357,In_517);
and U244 (N_244,In_603,In_788);
nor U245 (N_245,In_393,In_162);
nor U246 (N_246,In_696,In_229);
nand U247 (N_247,In_638,In_964);
nand U248 (N_248,In_269,In_850);
nand U249 (N_249,In_235,In_743);
nor U250 (N_250,In_320,In_175);
nand U251 (N_251,In_191,In_416);
nor U252 (N_252,In_251,In_944);
nand U253 (N_253,In_881,In_879);
nand U254 (N_254,In_464,In_254);
nand U255 (N_255,In_263,In_479);
and U256 (N_256,In_286,In_616);
or U257 (N_257,In_240,In_33);
xnor U258 (N_258,In_425,In_520);
and U259 (N_259,In_636,In_581);
or U260 (N_260,In_551,In_434);
nand U261 (N_261,In_224,In_95);
nor U262 (N_262,In_116,In_985);
and U263 (N_263,In_860,In_423);
nor U264 (N_264,In_504,In_380);
nand U265 (N_265,In_699,In_541);
nand U266 (N_266,In_302,In_447);
or U267 (N_267,In_929,In_621);
nor U268 (N_268,In_906,In_656);
or U269 (N_269,In_204,In_992);
or U270 (N_270,In_857,In_257);
and U271 (N_271,In_418,In_741);
nand U272 (N_272,In_875,In_597);
nor U273 (N_273,In_470,In_373);
or U274 (N_274,In_69,In_276);
and U275 (N_275,In_854,In_486);
and U276 (N_276,In_83,In_942);
xor U277 (N_277,In_146,In_126);
nand U278 (N_278,In_933,In_192);
and U279 (N_279,In_618,In_632);
nand U280 (N_280,In_288,In_383);
nor U281 (N_281,In_785,In_366);
and U282 (N_282,In_213,In_976);
nand U283 (N_283,In_259,In_316);
or U284 (N_284,In_268,In_271);
or U285 (N_285,In_414,In_957);
or U286 (N_286,In_151,In_92);
nor U287 (N_287,In_602,In_620);
nor U288 (N_288,In_797,In_168);
and U289 (N_289,In_283,In_821);
nand U290 (N_290,In_931,In_332);
and U291 (N_291,In_152,In_814);
nor U292 (N_292,In_890,In_131);
nor U293 (N_293,In_945,In_679);
and U294 (N_294,In_155,In_350);
and U295 (N_295,In_128,In_163);
and U296 (N_296,In_852,In_217);
or U297 (N_297,In_12,In_924);
nor U298 (N_298,In_108,In_960);
xnor U299 (N_299,In_536,In_236);
and U300 (N_300,In_227,In_778);
nand U301 (N_301,In_293,In_103);
and U302 (N_302,In_503,In_729);
or U303 (N_303,In_130,In_107);
or U304 (N_304,In_777,In_818);
nand U305 (N_305,In_812,In_801);
nor U306 (N_306,In_791,In_670);
or U307 (N_307,In_96,In_195);
nand U308 (N_308,In_478,In_367);
nor U309 (N_309,In_199,In_471);
nand U310 (N_310,In_768,In_810);
nor U311 (N_311,In_354,In_702);
and U312 (N_312,In_547,In_148);
or U313 (N_313,In_135,In_46);
or U314 (N_314,In_907,In_744);
xnor U315 (N_315,In_376,In_997);
nand U316 (N_316,In_735,In_463);
and U317 (N_317,In_643,In_73);
or U318 (N_318,In_466,In_896);
and U319 (N_319,In_323,In_612);
or U320 (N_320,In_639,In_949);
and U321 (N_321,In_766,In_482);
nand U322 (N_322,In_467,In_461);
and U323 (N_323,In_747,In_842);
or U324 (N_324,In_358,In_145);
and U325 (N_325,In_421,In_917);
and U326 (N_326,In_45,In_619);
nor U327 (N_327,In_353,In_545);
or U328 (N_328,In_993,In_542);
nand U329 (N_329,In_800,In_186);
and U330 (N_330,In_654,In_708);
nor U331 (N_331,In_218,In_80);
and U332 (N_332,In_27,In_726);
nor U333 (N_333,In_210,In_349);
or U334 (N_334,In_230,In_605);
and U335 (N_335,In_432,In_611);
nand U336 (N_336,In_442,In_487);
nand U337 (N_337,In_160,In_710);
and U338 (N_338,In_289,In_370);
and U339 (N_339,In_916,In_458);
and U340 (N_340,In_446,In_249);
or U341 (N_341,In_790,In_244);
nor U342 (N_342,In_607,In_566);
and U343 (N_343,In_764,In_374);
nand U344 (N_344,In_701,In_309);
or U345 (N_345,In_76,In_311);
nand U346 (N_346,In_722,In_782);
and U347 (N_347,In_623,In_171);
and U348 (N_348,In_278,In_928);
and U349 (N_349,In_728,In_905);
or U350 (N_350,In_909,In_239);
nand U351 (N_351,In_659,In_583);
nor U352 (N_352,In_969,In_307);
nor U353 (N_353,In_589,In_238);
or U354 (N_354,In_919,In_368);
or U355 (N_355,In_196,In_892);
and U356 (N_356,In_953,In_202);
and U357 (N_357,In_225,In_308);
and U358 (N_358,In_134,In_411);
nor U359 (N_359,In_817,In_170);
nor U360 (N_360,In_406,In_959);
and U361 (N_361,In_67,In_183);
or U362 (N_362,In_149,In_3);
nand U363 (N_363,In_869,In_395);
nand U364 (N_364,In_396,In_484);
or U365 (N_365,In_843,In_495);
nor U366 (N_366,In_662,In_465);
or U367 (N_367,In_226,In_99);
and U368 (N_368,In_233,In_164);
nor U369 (N_369,In_14,In_455);
or U370 (N_370,In_439,In_500);
and U371 (N_371,In_692,In_819);
nand U372 (N_372,In_751,In_982);
nand U373 (N_373,In_58,In_895);
nor U374 (N_374,In_925,In_122);
nor U375 (N_375,In_543,In_491);
nand U376 (N_376,In_951,In_342);
or U377 (N_377,In_105,In_34);
or U378 (N_378,In_647,In_938);
nand U379 (N_379,In_55,In_963);
and U380 (N_380,In_290,In_287);
or U381 (N_381,In_39,In_794);
nor U382 (N_382,In_66,In_322);
and U383 (N_383,In_301,In_669);
or U384 (N_384,In_772,In_665);
and U385 (N_385,In_124,In_552);
nor U386 (N_386,In_855,In_634);
nand U387 (N_387,In_996,In_734);
and U388 (N_388,In_802,In_859);
nor U389 (N_389,In_646,In_30);
or U390 (N_390,In_141,In_48);
nand U391 (N_391,In_575,In_60);
or U392 (N_392,In_294,In_893);
nor U393 (N_393,In_915,In_273);
nand U394 (N_394,In_433,In_114);
and U395 (N_395,In_9,In_437);
and U396 (N_396,In_438,In_779);
xnor U397 (N_397,In_245,In_232);
nor U398 (N_398,In_457,In_22);
nor U399 (N_399,In_110,In_594);
or U400 (N_400,In_576,In_365);
nand U401 (N_401,In_26,In_410);
and U402 (N_402,In_118,In_221);
or U403 (N_403,In_754,In_787);
nor U404 (N_404,In_176,In_324);
nor U405 (N_405,In_189,In_968);
or U406 (N_406,In_590,In_356);
nor U407 (N_407,In_206,In_262);
or U408 (N_408,In_803,In_868);
or U409 (N_409,In_644,In_506);
or U410 (N_410,In_488,In_549);
nor U411 (N_411,In_535,In_172);
nor U412 (N_412,In_736,In_127);
nor U413 (N_413,In_93,In_429);
or U414 (N_414,In_306,In_689);
and U415 (N_415,In_59,In_538);
nand U416 (N_416,In_144,In_921);
or U417 (N_417,In_330,In_712);
and U418 (N_418,In_598,In_377);
nand U419 (N_419,In_910,In_345);
nand U420 (N_420,In_809,In_508);
or U421 (N_421,In_851,In_981);
or U422 (N_422,In_473,In_63);
nand U423 (N_423,In_247,In_563);
and U424 (N_424,In_179,In_182);
or U425 (N_425,In_631,In_844);
or U426 (N_426,In_913,In_117);
nand U427 (N_427,In_415,In_700);
or U428 (N_428,In_770,In_515);
and U429 (N_429,In_102,In_622);
or U430 (N_430,In_668,In_456);
or U431 (N_431,In_573,In_228);
nor U432 (N_432,In_50,In_480);
and U433 (N_433,In_582,In_511);
or U434 (N_434,In_56,In_846);
nand U435 (N_435,In_837,In_664);
nor U436 (N_436,In_241,In_19);
or U437 (N_437,In_424,In_841);
or U438 (N_438,In_978,In_717);
nor U439 (N_439,In_789,In_384);
nor U440 (N_440,In_435,In_388);
or U441 (N_441,In_211,In_761);
and U442 (N_442,In_970,In_381);
nand U443 (N_443,In_222,In_606);
and U444 (N_444,In_950,In_811);
nand U445 (N_445,In_321,In_901);
and U446 (N_446,In_335,In_727);
and U447 (N_447,In_29,In_499);
and U448 (N_448,In_507,In_516);
and U449 (N_449,In_299,In_173);
nor U450 (N_450,In_74,In_64);
nand U451 (N_451,In_650,In_580);
nor U452 (N_452,In_277,In_292);
and U453 (N_453,In_363,In_653);
nor U454 (N_454,In_440,In_723);
and U455 (N_455,In_300,In_428);
and U456 (N_456,In_18,In_833);
nand U457 (N_457,In_312,In_866);
nor U458 (N_458,In_763,In_882);
nor U459 (N_459,In_972,In_561);
nand U460 (N_460,In_157,In_85);
and U461 (N_461,In_574,In_246);
nand U462 (N_462,In_876,In_431);
or U463 (N_463,In_401,In_123);
nor U464 (N_464,In_474,In_625);
nor U465 (N_465,In_685,In_44);
and U466 (N_466,In_444,In_265);
nand U467 (N_467,In_0,In_430);
or U468 (N_468,In_272,In_839);
and U469 (N_469,In_533,In_592);
nand U470 (N_470,In_956,In_209);
nor U471 (N_471,In_275,In_203);
or U472 (N_472,In_53,In_858);
or U473 (N_473,In_872,In_77);
and U474 (N_474,In_568,In_378);
nor U475 (N_475,In_519,In_84);
and U476 (N_476,In_531,In_492);
or U477 (N_477,In_261,In_715);
xor U478 (N_478,In_629,In_795);
nor U479 (N_479,In_62,In_617);
and U480 (N_480,In_836,In_297);
or U481 (N_481,In_862,In_663);
nor U482 (N_482,In_856,In_847);
and U483 (N_483,In_139,In_534);
nor U484 (N_484,In_834,In_158);
or U485 (N_485,In_5,In_207);
and U486 (N_486,In_540,In_762);
xnor U487 (N_487,In_677,In_28);
and U488 (N_488,In_89,In_205);
and U489 (N_489,In_714,In_922);
or U490 (N_490,In_767,In_212);
nand U491 (N_491,In_133,In_628);
nor U492 (N_492,In_153,In_453);
nand U493 (N_493,In_926,In_867);
or U494 (N_494,In_565,In_521);
nor U495 (N_495,In_137,In_595);
nor U496 (N_496,In_343,In_835);
and U497 (N_497,In_256,In_419);
nand U498 (N_498,In_999,In_17);
and U499 (N_499,In_562,In_709);
nor U500 (N_500,In_630,In_880);
and U501 (N_501,In_908,In_460);
nor U502 (N_502,In_753,In_304);
nand U503 (N_503,In_915,In_637);
nand U504 (N_504,In_259,In_682);
xnor U505 (N_505,In_76,In_965);
and U506 (N_506,In_604,In_38);
or U507 (N_507,In_594,In_692);
and U508 (N_508,In_493,In_939);
or U509 (N_509,In_312,In_228);
nand U510 (N_510,In_208,In_404);
or U511 (N_511,In_910,In_547);
nor U512 (N_512,In_614,In_932);
nor U513 (N_513,In_385,In_894);
and U514 (N_514,In_639,In_10);
xor U515 (N_515,In_402,In_215);
or U516 (N_516,In_39,In_440);
or U517 (N_517,In_302,In_485);
nand U518 (N_518,In_88,In_814);
or U519 (N_519,In_692,In_926);
nand U520 (N_520,In_878,In_865);
nor U521 (N_521,In_106,In_511);
or U522 (N_522,In_259,In_781);
nor U523 (N_523,In_833,In_850);
nor U524 (N_524,In_270,In_861);
or U525 (N_525,In_902,In_515);
or U526 (N_526,In_990,In_220);
and U527 (N_527,In_586,In_456);
or U528 (N_528,In_279,In_60);
and U529 (N_529,In_957,In_718);
or U530 (N_530,In_545,In_93);
nor U531 (N_531,In_598,In_915);
nor U532 (N_532,In_43,In_17);
or U533 (N_533,In_582,In_920);
and U534 (N_534,In_555,In_599);
nor U535 (N_535,In_870,In_422);
nor U536 (N_536,In_533,In_977);
or U537 (N_537,In_553,In_325);
or U538 (N_538,In_139,In_542);
or U539 (N_539,In_499,In_673);
nor U540 (N_540,In_664,In_540);
or U541 (N_541,In_563,In_227);
nor U542 (N_542,In_691,In_590);
and U543 (N_543,In_26,In_622);
or U544 (N_544,In_385,In_202);
nor U545 (N_545,In_68,In_117);
nand U546 (N_546,In_674,In_228);
and U547 (N_547,In_274,In_271);
nand U548 (N_548,In_828,In_691);
or U549 (N_549,In_886,In_778);
nor U550 (N_550,In_731,In_155);
or U551 (N_551,In_785,In_648);
and U552 (N_552,In_745,In_811);
and U553 (N_553,In_119,In_22);
nand U554 (N_554,In_688,In_907);
nand U555 (N_555,In_666,In_393);
nor U556 (N_556,In_910,In_52);
nor U557 (N_557,In_327,In_640);
and U558 (N_558,In_704,In_408);
or U559 (N_559,In_250,In_349);
nor U560 (N_560,In_478,In_480);
or U561 (N_561,In_214,In_560);
nand U562 (N_562,In_517,In_204);
and U563 (N_563,In_890,In_467);
or U564 (N_564,In_598,In_392);
nor U565 (N_565,In_919,In_540);
or U566 (N_566,In_114,In_318);
nor U567 (N_567,In_987,In_786);
and U568 (N_568,In_20,In_914);
nand U569 (N_569,In_500,In_922);
or U570 (N_570,In_73,In_128);
nand U571 (N_571,In_127,In_405);
nor U572 (N_572,In_554,In_800);
nand U573 (N_573,In_936,In_972);
nor U574 (N_574,In_853,In_389);
nor U575 (N_575,In_270,In_76);
and U576 (N_576,In_819,In_673);
or U577 (N_577,In_561,In_300);
nand U578 (N_578,In_83,In_465);
and U579 (N_579,In_192,In_887);
or U580 (N_580,In_569,In_81);
nand U581 (N_581,In_174,In_601);
and U582 (N_582,In_814,In_956);
or U583 (N_583,In_539,In_429);
nor U584 (N_584,In_220,In_2);
nand U585 (N_585,In_348,In_802);
nor U586 (N_586,In_416,In_271);
nand U587 (N_587,In_59,In_361);
nand U588 (N_588,In_664,In_39);
or U589 (N_589,In_474,In_596);
or U590 (N_590,In_265,In_604);
or U591 (N_591,In_751,In_742);
nor U592 (N_592,In_40,In_357);
nand U593 (N_593,In_236,In_481);
nand U594 (N_594,In_754,In_874);
and U595 (N_595,In_84,In_772);
and U596 (N_596,In_888,In_498);
or U597 (N_597,In_863,In_115);
nand U598 (N_598,In_775,In_999);
or U599 (N_599,In_134,In_845);
or U600 (N_600,In_294,In_106);
and U601 (N_601,In_876,In_784);
and U602 (N_602,In_670,In_137);
or U603 (N_603,In_222,In_439);
nand U604 (N_604,In_572,In_696);
nand U605 (N_605,In_502,In_750);
or U606 (N_606,In_18,In_956);
nand U607 (N_607,In_51,In_725);
nor U608 (N_608,In_959,In_300);
nand U609 (N_609,In_116,In_613);
and U610 (N_610,In_506,In_656);
or U611 (N_611,In_292,In_949);
nor U612 (N_612,In_569,In_928);
or U613 (N_613,In_117,In_336);
nand U614 (N_614,In_630,In_12);
nor U615 (N_615,In_708,In_8);
nand U616 (N_616,In_156,In_416);
nor U617 (N_617,In_628,In_643);
and U618 (N_618,In_630,In_58);
nand U619 (N_619,In_122,In_375);
nand U620 (N_620,In_50,In_988);
nor U621 (N_621,In_301,In_93);
nor U622 (N_622,In_149,In_594);
or U623 (N_623,In_896,In_291);
or U624 (N_624,In_218,In_817);
nor U625 (N_625,In_245,In_235);
and U626 (N_626,In_153,In_512);
nand U627 (N_627,In_930,In_955);
nand U628 (N_628,In_177,In_713);
nor U629 (N_629,In_659,In_506);
nor U630 (N_630,In_871,In_985);
and U631 (N_631,In_245,In_271);
nand U632 (N_632,In_953,In_34);
or U633 (N_633,In_177,In_675);
nor U634 (N_634,In_865,In_592);
nor U635 (N_635,In_928,In_157);
nand U636 (N_636,In_293,In_913);
or U637 (N_637,In_790,In_926);
or U638 (N_638,In_329,In_194);
and U639 (N_639,In_152,In_596);
or U640 (N_640,In_569,In_856);
and U641 (N_641,In_863,In_69);
or U642 (N_642,In_147,In_174);
and U643 (N_643,In_297,In_873);
and U644 (N_644,In_30,In_833);
or U645 (N_645,In_588,In_851);
nand U646 (N_646,In_867,In_374);
or U647 (N_647,In_838,In_328);
or U648 (N_648,In_90,In_74);
nand U649 (N_649,In_485,In_591);
nand U650 (N_650,In_335,In_579);
or U651 (N_651,In_213,In_354);
nor U652 (N_652,In_458,In_317);
and U653 (N_653,In_416,In_444);
xnor U654 (N_654,In_354,In_540);
or U655 (N_655,In_294,In_139);
nor U656 (N_656,In_659,In_693);
or U657 (N_657,In_861,In_427);
or U658 (N_658,In_530,In_204);
nor U659 (N_659,In_791,In_808);
nand U660 (N_660,In_956,In_810);
nor U661 (N_661,In_545,In_478);
and U662 (N_662,In_784,In_203);
and U663 (N_663,In_676,In_45);
or U664 (N_664,In_841,In_364);
nand U665 (N_665,In_767,In_864);
and U666 (N_666,In_725,In_272);
xnor U667 (N_667,In_281,In_293);
xnor U668 (N_668,In_325,In_110);
or U669 (N_669,In_712,In_157);
and U670 (N_670,In_99,In_5);
xnor U671 (N_671,In_476,In_849);
nor U672 (N_672,In_216,In_303);
xor U673 (N_673,In_13,In_824);
xnor U674 (N_674,In_230,In_432);
nand U675 (N_675,In_963,In_408);
and U676 (N_676,In_439,In_724);
or U677 (N_677,In_893,In_189);
xnor U678 (N_678,In_170,In_620);
nand U679 (N_679,In_640,In_902);
nand U680 (N_680,In_486,In_135);
nor U681 (N_681,In_411,In_11);
and U682 (N_682,In_96,In_533);
nor U683 (N_683,In_539,In_382);
or U684 (N_684,In_25,In_477);
or U685 (N_685,In_872,In_118);
and U686 (N_686,In_371,In_906);
nor U687 (N_687,In_334,In_435);
or U688 (N_688,In_460,In_923);
and U689 (N_689,In_924,In_576);
or U690 (N_690,In_337,In_4);
nor U691 (N_691,In_326,In_976);
or U692 (N_692,In_597,In_84);
and U693 (N_693,In_85,In_854);
and U694 (N_694,In_20,In_434);
xor U695 (N_695,In_297,In_554);
and U696 (N_696,In_931,In_537);
nor U697 (N_697,In_659,In_217);
nor U698 (N_698,In_828,In_686);
or U699 (N_699,In_583,In_465);
nor U700 (N_700,In_593,In_386);
nand U701 (N_701,In_16,In_412);
nand U702 (N_702,In_823,In_439);
nor U703 (N_703,In_687,In_754);
nor U704 (N_704,In_20,In_968);
or U705 (N_705,In_300,In_433);
nand U706 (N_706,In_497,In_279);
nand U707 (N_707,In_508,In_16);
nand U708 (N_708,In_700,In_666);
nor U709 (N_709,In_541,In_713);
or U710 (N_710,In_818,In_72);
nor U711 (N_711,In_920,In_857);
nor U712 (N_712,In_24,In_253);
nor U713 (N_713,In_605,In_300);
nand U714 (N_714,In_968,In_182);
nand U715 (N_715,In_665,In_120);
and U716 (N_716,In_539,In_887);
or U717 (N_717,In_768,In_231);
and U718 (N_718,In_125,In_112);
or U719 (N_719,In_465,In_288);
or U720 (N_720,In_48,In_75);
and U721 (N_721,In_522,In_476);
xnor U722 (N_722,In_92,In_162);
and U723 (N_723,In_751,In_932);
nand U724 (N_724,In_277,In_637);
or U725 (N_725,In_679,In_0);
nand U726 (N_726,In_137,In_857);
nand U727 (N_727,In_790,In_966);
nand U728 (N_728,In_279,In_391);
nor U729 (N_729,In_516,In_287);
nor U730 (N_730,In_657,In_679);
nand U731 (N_731,In_977,In_129);
nand U732 (N_732,In_929,In_687);
nor U733 (N_733,In_478,In_670);
nand U734 (N_734,In_829,In_20);
nand U735 (N_735,In_821,In_762);
nand U736 (N_736,In_81,In_456);
or U737 (N_737,In_221,In_473);
nand U738 (N_738,In_910,In_13);
or U739 (N_739,In_399,In_331);
nand U740 (N_740,In_485,In_338);
nand U741 (N_741,In_113,In_985);
nand U742 (N_742,In_64,In_168);
nor U743 (N_743,In_63,In_615);
and U744 (N_744,In_306,In_265);
or U745 (N_745,In_281,In_329);
nor U746 (N_746,In_928,In_302);
or U747 (N_747,In_222,In_329);
nand U748 (N_748,In_67,In_144);
and U749 (N_749,In_305,In_463);
or U750 (N_750,In_653,In_989);
or U751 (N_751,In_753,In_712);
and U752 (N_752,In_435,In_556);
or U753 (N_753,In_332,In_157);
nor U754 (N_754,In_791,In_872);
nor U755 (N_755,In_781,In_756);
nand U756 (N_756,In_849,In_919);
and U757 (N_757,In_885,In_584);
or U758 (N_758,In_948,In_747);
or U759 (N_759,In_124,In_384);
and U760 (N_760,In_142,In_867);
and U761 (N_761,In_878,In_930);
nand U762 (N_762,In_568,In_418);
nand U763 (N_763,In_106,In_203);
and U764 (N_764,In_261,In_796);
and U765 (N_765,In_717,In_99);
and U766 (N_766,In_626,In_23);
nor U767 (N_767,In_469,In_988);
nor U768 (N_768,In_109,In_249);
nand U769 (N_769,In_90,In_15);
or U770 (N_770,In_404,In_386);
nand U771 (N_771,In_162,In_277);
nand U772 (N_772,In_558,In_192);
nor U773 (N_773,In_205,In_171);
nand U774 (N_774,In_342,In_895);
and U775 (N_775,In_437,In_363);
nor U776 (N_776,In_846,In_642);
nand U777 (N_777,In_686,In_776);
or U778 (N_778,In_518,In_418);
and U779 (N_779,In_135,In_290);
and U780 (N_780,In_171,In_63);
and U781 (N_781,In_45,In_930);
and U782 (N_782,In_821,In_211);
nand U783 (N_783,In_382,In_84);
nor U784 (N_784,In_799,In_88);
nand U785 (N_785,In_116,In_699);
or U786 (N_786,In_819,In_364);
nand U787 (N_787,In_255,In_757);
or U788 (N_788,In_13,In_589);
or U789 (N_789,In_379,In_617);
and U790 (N_790,In_957,In_715);
or U791 (N_791,In_680,In_793);
and U792 (N_792,In_141,In_978);
nor U793 (N_793,In_927,In_80);
or U794 (N_794,In_812,In_899);
and U795 (N_795,In_512,In_174);
and U796 (N_796,In_409,In_878);
nand U797 (N_797,In_425,In_558);
nor U798 (N_798,In_784,In_96);
nor U799 (N_799,In_570,In_798);
nor U800 (N_800,In_556,In_116);
and U801 (N_801,In_354,In_400);
nor U802 (N_802,In_169,In_733);
nor U803 (N_803,In_330,In_497);
nand U804 (N_804,In_883,In_595);
and U805 (N_805,In_419,In_347);
nor U806 (N_806,In_833,In_605);
nor U807 (N_807,In_525,In_682);
or U808 (N_808,In_973,In_509);
nand U809 (N_809,In_525,In_88);
or U810 (N_810,In_410,In_943);
or U811 (N_811,In_251,In_128);
and U812 (N_812,In_330,In_397);
xnor U813 (N_813,In_54,In_863);
nand U814 (N_814,In_100,In_708);
nor U815 (N_815,In_456,In_691);
and U816 (N_816,In_26,In_173);
nand U817 (N_817,In_435,In_305);
nor U818 (N_818,In_584,In_708);
and U819 (N_819,In_845,In_433);
and U820 (N_820,In_298,In_610);
and U821 (N_821,In_84,In_5);
or U822 (N_822,In_934,In_574);
and U823 (N_823,In_746,In_190);
or U824 (N_824,In_97,In_418);
and U825 (N_825,In_857,In_249);
and U826 (N_826,In_674,In_849);
nand U827 (N_827,In_201,In_824);
nor U828 (N_828,In_769,In_427);
or U829 (N_829,In_116,In_948);
nand U830 (N_830,In_553,In_8);
and U831 (N_831,In_260,In_124);
and U832 (N_832,In_521,In_865);
nand U833 (N_833,In_48,In_423);
nand U834 (N_834,In_839,In_178);
nand U835 (N_835,In_359,In_462);
nand U836 (N_836,In_648,In_520);
or U837 (N_837,In_626,In_328);
and U838 (N_838,In_60,In_72);
or U839 (N_839,In_968,In_9);
nor U840 (N_840,In_815,In_38);
or U841 (N_841,In_157,In_792);
or U842 (N_842,In_112,In_362);
nand U843 (N_843,In_529,In_838);
xor U844 (N_844,In_311,In_742);
and U845 (N_845,In_294,In_652);
nand U846 (N_846,In_952,In_232);
nor U847 (N_847,In_538,In_258);
nor U848 (N_848,In_993,In_157);
or U849 (N_849,In_654,In_370);
or U850 (N_850,In_610,In_814);
nor U851 (N_851,In_988,In_367);
nor U852 (N_852,In_198,In_958);
or U853 (N_853,In_950,In_798);
or U854 (N_854,In_867,In_245);
and U855 (N_855,In_619,In_396);
nor U856 (N_856,In_201,In_547);
or U857 (N_857,In_531,In_433);
and U858 (N_858,In_916,In_45);
and U859 (N_859,In_216,In_603);
nand U860 (N_860,In_410,In_760);
and U861 (N_861,In_912,In_742);
or U862 (N_862,In_264,In_32);
nor U863 (N_863,In_255,In_645);
or U864 (N_864,In_137,In_518);
or U865 (N_865,In_813,In_803);
nor U866 (N_866,In_331,In_934);
and U867 (N_867,In_205,In_65);
and U868 (N_868,In_147,In_97);
nand U869 (N_869,In_854,In_923);
nand U870 (N_870,In_605,In_460);
nor U871 (N_871,In_358,In_553);
nand U872 (N_872,In_467,In_844);
and U873 (N_873,In_13,In_947);
nand U874 (N_874,In_80,In_188);
nand U875 (N_875,In_100,In_440);
or U876 (N_876,In_777,In_976);
and U877 (N_877,In_698,In_304);
or U878 (N_878,In_90,In_273);
nand U879 (N_879,In_375,In_754);
or U880 (N_880,In_418,In_948);
nand U881 (N_881,In_309,In_99);
and U882 (N_882,In_928,In_646);
nand U883 (N_883,In_720,In_332);
nor U884 (N_884,In_529,In_101);
nand U885 (N_885,In_189,In_928);
nand U886 (N_886,In_906,In_387);
nor U887 (N_887,In_101,In_240);
nand U888 (N_888,In_10,In_783);
or U889 (N_889,In_239,In_961);
and U890 (N_890,In_271,In_760);
or U891 (N_891,In_478,In_552);
and U892 (N_892,In_700,In_274);
or U893 (N_893,In_638,In_899);
nor U894 (N_894,In_961,In_280);
and U895 (N_895,In_58,In_328);
nand U896 (N_896,In_665,In_795);
or U897 (N_897,In_465,In_537);
or U898 (N_898,In_20,In_166);
nand U899 (N_899,In_817,In_767);
or U900 (N_900,In_71,In_247);
nor U901 (N_901,In_242,In_94);
nand U902 (N_902,In_140,In_862);
and U903 (N_903,In_785,In_523);
or U904 (N_904,In_39,In_550);
nor U905 (N_905,In_867,In_208);
nand U906 (N_906,In_106,In_219);
nand U907 (N_907,In_671,In_496);
or U908 (N_908,In_738,In_72);
nand U909 (N_909,In_992,In_420);
nand U910 (N_910,In_982,In_374);
nand U911 (N_911,In_798,In_231);
nand U912 (N_912,In_762,In_403);
or U913 (N_913,In_899,In_16);
or U914 (N_914,In_280,In_428);
and U915 (N_915,In_968,In_301);
and U916 (N_916,In_796,In_709);
and U917 (N_917,In_70,In_663);
nor U918 (N_918,In_629,In_56);
nand U919 (N_919,In_108,In_619);
or U920 (N_920,In_880,In_156);
nor U921 (N_921,In_643,In_266);
nand U922 (N_922,In_96,In_524);
nor U923 (N_923,In_528,In_536);
and U924 (N_924,In_505,In_701);
or U925 (N_925,In_536,In_743);
nor U926 (N_926,In_163,In_650);
nand U927 (N_927,In_560,In_877);
nand U928 (N_928,In_151,In_254);
and U929 (N_929,In_403,In_301);
or U930 (N_930,In_131,In_484);
nand U931 (N_931,In_552,In_885);
xnor U932 (N_932,In_550,In_109);
nand U933 (N_933,In_747,In_27);
and U934 (N_934,In_134,In_838);
and U935 (N_935,In_137,In_459);
or U936 (N_936,In_517,In_964);
and U937 (N_937,In_743,In_926);
nand U938 (N_938,In_113,In_339);
nor U939 (N_939,In_49,In_130);
nor U940 (N_940,In_280,In_966);
and U941 (N_941,In_451,In_720);
and U942 (N_942,In_368,In_937);
and U943 (N_943,In_942,In_947);
nor U944 (N_944,In_44,In_272);
nand U945 (N_945,In_655,In_714);
nand U946 (N_946,In_269,In_17);
nand U947 (N_947,In_696,In_680);
nand U948 (N_948,In_933,In_52);
nor U949 (N_949,In_246,In_705);
nand U950 (N_950,In_309,In_642);
and U951 (N_951,In_226,In_356);
nor U952 (N_952,In_857,In_531);
nor U953 (N_953,In_748,In_706);
or U954 (N_954,In_635,In_700);
and U955 (N_955,In_265,In_989);
or U956 (N_956,In_62,In_359);
or U957 (N_957,In_983,In_982);
nor U958 (N_958,In_870,In_625);
and U959 (N_959,In_767,In_602);
or U960 (N_960,In_816,In_215);
nand U961 (N_961,In_63,In_689);
and U962 (N_962,In_2,In_604);
nand U963 (N_963,In_343,In_139);
or U964 (N_964,In_793,In_434);
and U965 (N_965,In_103,In_550);
and U966 (N_966,In_797,In_741);
xor U967 (N_967,In_664,In_221);
and U968 (N_968,In_582,In_418);
nor U969 (N_969,In_908,In_113);
and U970 (N_970,In_402,In_756);
or U971 (N_971,In_411,In_986);
nor U972 (N_972,In_117,In_141);
nor U973 (N_973,In_626,In_834);
or U974 (N_974,In_768,In_789);
nand U975 (N_975,In_135,In_591);
nand U976 (N_976,In_941,In_1);
or U977 (N_977,In_363,In_559);
nor U978 (N_978,In_23,In_510);
nor U979 (N_979,In_432,In_776);
and U980 (N_980,In_76,In_847);
or U981 (N_981,In_721,In_718);
nand U982 (N_982,In_444,In_208);
nor U983 (N_983,In_935,In_446);
nand U984 (N_984,In_724,In_395);
or U985 (N_985,In_492,In_261);
nand U986 (N_986,In_563,In_535);
nand U987 (N_987,In_723,In_809);
or U988 (N_988,In_56,In_837);
nand U989 (N_989,In_984,In_785);
and U990 (N_990,In_893,In_194);
or U991 (N_991,In_40,In_163);
nor U992 (N_992,In_672,In_955);
or U993 (N_993,In_449,In_314);
nand U994 (N_994,In_797,In_230);
nand U995 (N_995,In_243,In_75);
nor U996 (N_996,In_556,In_105);
and U997 (N_997,In_627,In_397);
nor U998 (N_998,In_821,In_39);
and U999 (N_999,In_957,In_8);
nor U1000 (N_1000,In_466,In_796);
or U1001 (N_1001,In_189,In_507);
nor U1002 (N_1002,In_995,In_300);
nand U1003 (N_1003,In_363,In_615);
nand U1004 (N_1004,In_230,In_831);
nand U1005 (N_1005,In_201,In_71);
nand U1006 (N_1006,In_100,In_585);
xnor U1007 (N_1007,In_497,In_644);
nor U1008 (N_1008,In_422,In_997);
or U1009 (N_1009,In_137,In_657);
and U1010 (N_1010,In_181,In_995);
nor U1011 (N_1011,In_147,In_145);
or U1012 (N_1012,In_637,In_523);
nor U1013 (N_1013,In_933,In_212);
or U1014 (N_1014,In_66,In_427);
or U1015 (N_1015,In_984,In_165);
or U1016 (N_1016,In_384,In_788);
or U1017 (N_1017,In_706,In_547);
nand U1018 (N_1018,In_344,In_213);
nor U1019 (N_1019,In_709,In_177);
nor U1020 (N_1020,In_196,In_880);
nand U1021 (N_1021,In_770,In_605);
nor U1022 (N_1022,In_116,In_16);
or U1023 (N_1023,In_483,In_642);
nand U1024 (N_1024,In_570,In_88);
or U1025 (N_1025,In_517,In_674);
or U1026 (N_1026,In_420,In_889);
nand U1027 (N_1027,In_787,In_993);
nand U1028 (N_1028,In_397,In_621);
or U1029 (N_1029,In_234,In_370);
and U1030 (N_1030,In_78,In_211);
and U1031 (N_1031,In_371,In_437);
nor U1032 (N_1032,In_398,In_945);
and U1033 (N_1033,In_720,In_836);
nor U1034 (N_1034,In_766,In_175);
and U1035 (N_1035,In_999,In_889);
nor U1036 (N_1036,In_628,In_314);
or U1037 (N_1037,In_941,In_185);
nand U1038 (N_1038,In_841,In_451);
nor U1039 (N_1039,In_925,In_480);
and U1040 (N_1040,In_680,In_587);
or U1041 (N_1041,In_299,In_131);
and U1042 (N_1042,In_14,In_85);
and U1043 (N_1043,In_948,In_798);
nor U1044 (N_1044,In_303,In_523);
nor U1045 (N_1045,In_58,In_953);
nor U1046 (N_1046,In_830,In_208);
and U1047 (N_1047,In_174,In_372);
nor U1048 (N_1048,In_387,In_620);
xor U1049 (N_1049,In_30,In_275);
and U1050 (N_1050,In_289,In_452);
nor U1051 (N_1051,In_768,In_529);
or U1052 (N_1052,In_628,In_732);
nor U1053 (N_1053,In_179,In_85);
nand U1054 (N_1054,In_533,In_230);
and U1055 (N_1055,In_886,In_807);
and U1056 (N_1056,In_480,In_939);
nand U1057 (N_1057,In_996,In_217);
and U1058 (N_1058,In_555,In_422);
nand U1059 (N_1059,In_313,In_670);
nor U1060 (N_1060,In_278,In_25);
or U1061 (N_1061,In_34,In_218);
or U1062 (N_1062,In_484,In_106);
nand U1063 (N_1063,In_692,In_72);
nand U1064 (N_1064,In_851,In_866);
or U1065 (N_1065,In_168,In_909);
nand U1066 (N_1066,In_949,In_719);
nor U1067 (N_1067,In_907,In_957);
nand U1068 (N_1068,In_696,In_494);
or U1069 (N_1069,In_933,In_800);
and U1070 (N_1070,In_342,In_518);
and U1071 (N_1071,In_541,In_49);
and U1072 (N_1072,In_503,In_809);
and U1073 (N_1073,In_907,In_542);
nand U1074 (N_1074,In_752,In_932);
nor U1075 (N_1075,In_286,In_576);
nor U1076 (N_1076,In_605,In_739);
and U1077 (N_1077,In_316,In_568);
xor U1078 (N_1078,In_711,In_354);
or U1079 (N_1079,In_456,In_320);
or U1080 (N_1080,In_204,In_749);
nand U1081 (N_1081,In_586,In_731);
nand U1082 (N_1082,In_24,In_840);
or U1083 (N_1083,In_193,In_146);
nand U1084 (N_1084,In_865,In_926);
nor U1085 (N_1085,In_811,In_965);
xnor U1086 (N_1086,In_880,In_268);
or U1087 (N_1087,In_150,In_744);
and U1088 (N_1088,In_959,In_28);
nor U1089 (N_1089,In_945,In_961);
or U1090 (N_1090,In_144,In_677);
nand U1091 (N_1091,In_650,In_883);
or U1092 (N_1092,In_132,In_634);
or U1093 (N_1093,In_175,In_325);
nor U1094 (N_1094,In_196,In_409);
or U1095 (N_1095,In_169,In_647);
nor U1096 (N_1096,In_231,In_637);
and U1097 (N_1097,In_31,In_78);
or U1098 (N_1098,In_824,In_502);
nor U1099 (N_1099,In_903,In_667);
or U1100 (N_1100,In_107,In_556);
nor U1101 (N_1101,In_641,In_299);
nor U1102 (N_1102,In_585,In_594);
nor U1103 (N_1103,In_401,In_599);
or U1104 (N_1104,In_995,In_916);
nor U1105 (N_1105,In_142,In_594);
and U1106 (N_1106,In_78,In_12);
nor U1107 (N_1107,In_531,In_285);
and U1108 (N_1108,In_12,In_227);
and U1109 (N_1109,In_768,In_389);
nand U1110 (N_1110,In_966,In_180);
nor U1111 (N_1111,In_667,In_478);
and U1112 (N_1112,In_107,In_564);
and U1113 (N_1113,In_3,In_172);
nand U1114 (N_1114,In_622,In_686);
nand U1115 (N_1115,In_348,In_785);
nand U1116 (N_1116,In_617,In_647);
nor U1117 (N_1117,In_784,In_831);
nand U1118 (N_1118,In_718,In_578);
and U1119 (N_1119,In_970,In_476);
nor U1120 (N_1120,In_390,In_541);
nand U1121 (N_1121,In_232,In_227);
nand U1122 (N_1122,In_849,In_216);
nor U1123 (N_1123,In_368,In_235);
nor U1124 (N_1124,In_288,In_974);
nand U1125 (N_1125,In_32,In_602);
nand U1126 (N_1126,In_958,In_110);
nand U1127 (N_1127,In_100,In_896);
and U1128 (N_1128,In_928,In_966);
or U1129 (N_1129,In_48,In_46);
or U1130 (N_1130,In_393,In_525);
nand U1131 (N_1131,In_646,In_492);
nand U1132 (N_1132,In_249,In_887);
nor U1133 (N_1133,In_908,In_706);
nand U1134 (N_1134,In_463,In_368);
nor U1135 (N_1135,In_133,In_693);
nand U1136 (N_1136,In_621,In_159);
nand U1137 (N_1137,In_220,In_734);
nand U1138 (N_1138,In_571,In_439);
and U1139 (N_1139,In_774,In_609);
nor U1140 (N_1140,In_279,In_825);
nor U1141 (N_1141,In_201,In_805);
nor U1142 (N_1142,In_0,In_175);
and U1143 (N_1143,In_253,In_880);
nor U1144 (N_1144,In_719,In_44);
nor U1145 (N_1145,In_405,In_492);
or U1146 (N_1146,In_700,In_575);
and U1147 (N_1147,In_98,In_797);
and U1148 (N_1148,In_627,In_848);
or U1149 (N_1149,In_208,In_175);
and U1150 (N_1150,In_678,In_371);
or U1151 (N_1151,In_348,In_127);
or U1152 (N_1152,In_19,In_217);
or U1153 (N_1153,In_567,In_429);
and U1154 (N_1154,In_688,In_323);
nand U1155 (N_1155,In_680,In_236);
nand U1156 (N_1156,In_588,In_517);
nand U1157 (N_1157,In_120,In_271);
nor U1158 (N_1158,In_238,In_237);
nor U1159 (N_1159,In_552,In_674);
nor U1160 (N_1160,In_10,In_422);
and U1161 (N_1161,In_97,In_496);
and U1162 (N_1162,In_594,In_925);
or U1163 (N_1163,In_267,In_914);
nand U1164 (N_1164,In_534,In_952);
or U1165 (N_1165,In_334,In_610);
nand U1166 (N_1166,In_311,In_216);
nand U1167 (N_1167,In_825,In_516);
nor U1168 (N_1168,In_457,In_854);
nand U1169 (N_1169,In_315,In_938);
nor U1170 (N_1170,In_300,In_227);
nor U1171 (N_1171,In_187,In_388);
and U1172 (N_1172,In_259,In_964);
or U1173 (N_1173,In_306,In_897);
and U1174 (N_1174,In_580,In_586);
nand U1175 (N_1175,In_99,In_30);
nor U1176 (N_1176,In_7,In_319);
nand U1177 (N_1177,In_383,In_262);
nand U1178 (N_1178,In_417,In_800);
nor U1179 (N_1179,In_402,In_147);
and U1180 (N_1180,In_985,In_353);
and U1181 (N_1181,In_907,In_547);
nor U1182 (N_1182,In_704,In_211);
and U1183 (N_1183,In_300,In_766);
nand U1184 (N_1184,In_317,In_510);
nand U1185 (N_1185,In_19,In_467);
and U1186 (N_1186,In_720,In_309);
and U1187 (N_1187,In_914,In_765);
nand U1188 (N_1188,In_927,In_783);
nor U1189 (N_1189,In_167,In_857);
and U1190 (N_1190,In_104,In_896);
nand U1191 (N_1191,In_685,In_731);
nor U1192 (N_1192,In_686,In_110);
nand U1193 (N_1193,In_724,In_72);
nor U1194 (N_1194,In_585,In_382);
nand U1195 (N_1195,In_757,In_890);
nor U1196 (N_1196,In_948,In_194);
or U1197 (N_1197,In_673,In_501);
nor U1198 (N_1198,In_744,In_877);
nor U1199 (N_1199,In_331,In_306);
nor U1200 (N_1200,In_784,In_418);
nand U1201 (N_1201,In_67,In_315);
nand U1202 (N_1202,In_366,In_413);
nand U1203 (N_1203,In_111,In_106);
and U1204 (N_1204,In_353,In_756);
or U1205 (N_1205,In_372,In_669);
or U1206 (N_1206,In_306,In_225);
nand U1207 (N_1207,In_492,In_159);
or U1208 (N_1208,In_347,In_133);
nor U1209 (N_1209,In_180,In_974);
nor U1210 (N_1210,In_23,In_5);
nand U1211 (N_1211,In_814,In_576);
and U1212 (N_1212,In_600,In_191);
nand U1213 (N_1213,In_742,In_281);
or U1214 (N_1214,In_18,In_553);
or U1215 (N_1215,In_659,In_28);
or U1216 (N_1216,In_816,In_267);
or U1217 (N_1217,In_372,In_821);
nor U1218 (N_1218,In_939,In_899);
nand U1219 (N_1219,In_751,In_948);
nand U1220 (N_1220,In_883,In_132);
or U1221 (N_1221,In_894,In_196);
nor U1222 (N_1222,In_112,In_634);
or U1223 (N_1223,In_926,In_165);
or U1224 (N_1224,In_768,In_352);
nand U1225 (N_1225,In_355,In_144);
or U1226 (N_1226,In_775,In_401);
nor U1227 (N_1227,In_748,In_130);
and U1228 (N_1228,In_679,In_847);
nand U1229 (N_1229,In_668,In_956);
nand U1230 (N_1230,In_382,In_905);
nor U1231 (N_1231,In_825,In_933);
and U1232 (N_1232,In_459,In_290);
nand U1233 (N_1233,In_898,In_494);
and U1234 (N_1234,In_933,In_727);
or U1235 (N_1235,In_374,In_476);
or U1236 (N_1236,In_27,In_190);
nor U1237 (N_1237,In_616,In_757);
and U1238 (N_1238,In_897,In_848);
nand U1239 (N_1239,In_112,In_818);
nand U1240 (N_1240,In_201,In_959);
nor U1241 (N_1241,In_450,In_974);
and U1242 (N_1242,In_764,In_375);
or U1243 (N_1243,In_88,In_837);
and U1244 (N_1244,In_556,In_200);
or U1245 (N_1245,In_209,In_447);
and U1246 (N_1246,In_502,In_329);
or U1247 (N_1247,In_865,In_278);
nand U1248 (N_1248,In_759,In_6);
or U1249 (N_1249,In_926,In_164);
or U1250 (N_1250,In_483,In_388);
and U1251 (N_1251,In_145,In_835);
or U1252 (N_1252,In_318,In_739);
or U1253 (N_1253,In_154,In_84);
nand U1254 (N_1254,In_39,In_595);
nand U1255 (N_1255,In_362,In_381);
nand U1256 (N_1256,In_239,In_786);
nand U1257 (N_1257,In_878,In_991);
nand U1258 (N_1258,In_850,In_860);
and U1259 (N_1259,In_905,In_174);
nand U1260 (N_1260,In_99,In_523);
or U1261 (N_1261,In_658,In_568);
nand U1262 (N_1262,In_282,In_488);
nand U1263 (N_1263,In_198,In_941);
and U1264 (N_1264,In_169,In_531);
and U1265 (N_1265,In_715,In_803);
nor U1266 (N_1266,In_158,In_714);
or U1267 (N_1267,In_181,In_129);
and U1268 (N_1268,In_957,In_473);
or U1269 (N_1269,In_517,In_808);
or U1270 (N_1270,In_392,In_729);
or U1271 (N_1271,In_79,In_421);
nand U1272 (N_1272,In_399,In_724);
and U1273 (N_1273,In_249,In_64);
or U1274 (N_1274,In_991,In_435);
xnor U1275 (N_1275,In_298,In_152);
and U1276 (N_1276,In_576,In_556);
nand U1277 (N_1277,In_334,In_187);
nand U1278 (N_1278,In_668,In_441);
nor U1279 (N_1279,In_617,In_858);
and U1280 (N_1280,In_929,In_765);
and U1281 (N_1281,In_962,In_385);
nand U1282 (N_1282,In_388,In_456);
and U1283 (N_1283,In_660,In_783);
or U1284 (N_1284,In_275,In_118);
nor U1285 (N_1285,In_798,In_458);
or U1286 (N_1286,In_754,In_351);
or U1287 (N_1287,In_400,In_912);
and U1288 (N_1288,In_678,In_103);
or U1289 (N_1289,In_62,In_840);
nand U1290 (N_1290,In_496,In_119);
nor U1291 (N_1291,In_841,In_259);
and U1292 (N_1292,In_885,In_427);
nor U1293 (N_1293,In_892,In_586);
nor U1294 (N_1294,In_164,In_981);
nor U1295 (N_1295,In_962,In_595);
or U1296 (N_1296,In_954,In_732);
nor U1297 (N_1297,In_992,In_105);
and U1298 (N_1298,In_477,In_629);
and U1299 (N_1299,In_354,In_140);
nand U1300 (N_1300,In_89,In_452);
nand U1301 (N_1301,In_716,In_108);
or U1302 (N_1302,In_7,In_735);
nand U1303 (N_1303,In_322,In_104);
or U1304 (N_1304,In_730,In_965);
or U1305 (N_1305,In_31,In_477);
nand U1306 (N_1306,In_795,In_119);
or U1307 (N_1307,In_15,In_214);
or U1308 (N_1308,In_81,In_101);
nor U1309 (N_1309,In_679,In_598);
nor U1310 (N_1310,In_565,In_910);
and U1311 (N_1311,In_56,In_302);
or U1312 (N_1312,In_360,In_801);
nor U1313 (N_1313,In_86,In_951);
or U1314 (N_1314,In_186,In_61);
and U1315 (N_1315,In_49,In_996);
nor U1316 (N_1316,In_20,In_154);
nor U1317 (N_1317,In_164,In_416);
or U1318 (N_1318,In_373,In_575);
or U1319 (N_1319,In_146,In_119);
nand U1320 (N_1320,In_383,In_99);
and U1321 (N_1321,In_38,In_759);
and U1322 (N_1322,In_275,In_4);
nand U1323 (N_1323,In_707,In_791);
nand U1324 (N_1324,In_924,In_993);
nor U1325 (N_1325,In_909,In_569);
and U1326 (N_1326,In_340,In_224);
or U1327 (N_1327,In_229,In_895);
nand U1328 (N_1328,In_726,In_352);
nand U1329 (N_1329,In_37,In_106);
nand U1330 (N_1330,In_913,In_513);
or U1331 (N_1331,In_287,In_538);
nand U1332 (N_1332,In_632,In_821);
or U1333 (N_1333,In_641,In_116);
or U1334 (N_1334,In_140,In_398);
and U1335 (N_1335,In_251,In_969);
and U1336 (N_1336,In_241,In_25);
nor U1337 (N_1337,In_750,In_375);
and U1338 (N_1338,In_369,In_599);
and U1339 (N_1339,In_597,In_665);
nand U1340 (N_1340,In_160,In_453);
nand U1341 (N_1341,In_702,In_405);
nor U1342 (N_1342,In_496,In_847);
nand U1343 (N_1343,In_591,In_495);
and U1344 (N_1344,In_825,In_327);
nand U1345 (N_1345,In_350,In_359);
nor U1346 (N_1346,In_211,In_900);
nand U1347 (N_1347,In_361,In_189);
or U1348 (N_1348,In_861,In_148);
or U1349 (N_1349,In_208,In_255);
nor U1350 (N_1350,In_487,In_895);
or U1351 (N_1351,In_617,In_662);
or U1352 (N_1352,In_962,In_660);
or U1353 (N_1353,In_783,In_292);
or U1354 (N_1354,In_567,In_214);
nand U1355 (N_1355,In_786,In_88);
and U1356 (N_1356,In_643,In_570);
nand U1357 (N_1357,In_939,In_537);
or U1358 (N_1358,In_415,In_73);
nand U1359 (N_1359,In_664,In_319);
nand U1360 (N_1360,In_559,In_440);
or U1361 (N_1361,In_436,In_829);
xnor U1362 (N_1362,In_870,In_656);
nand U1363 (N_1363,In_398,In_58);
nand U1364 (N_1364,In_398,In_456);
nand U1365 (N_1365,In_551,In_282);
nand U1366 (N_1366,In_145,In_377);
xnor U1367 (N_1367,In_52,In_484);
or U1368 (N_1368,In_904,In_262);
and U1369 (N_1369,In_949,In_165);
or U1370 (N_1370,In_311,In_526);
or U1371 (N_1371,In_569,In_622);
nand U1372 (N_1372,In_239,In_369);
and U1373 (N_1373,In_239,In_689);
nor U1374 (N_1374,In_98,In_614);
or U1375 (N_1375,In_912,In_852);
and U1376 (N_1376,In_702,In_107);
nor U1377 (N_1377,In_718,In_728);
or U1378 (N_1378,In_994,In_599);
or U1379 (N_1379,In_324,In_97);
or U1380 (N_1380,In_168,In_281);
or U1381 (N_1381,In_291,In_853);
or U1382 (N_1382,In_553,In_216);
nand U1383 (N_1383,In_646,In_896);
nand U1384 (N_1384,In_100,In_40);
and U1385 (N_1385,In_616,In_881);
and U1386 (N_1386,In_514,In_984);
or U1387 (N_1387,In_906,In_106);
and U1388 (N_1388,In_422,In_320);
nand U1389 (N_1389,In_1,In_975);
nor U1390 (N_1390,In_382,In_876);
nand U1391 (N_1391,In_120,In_393);
or U1392 (N_1392,In_249,In_936);
nand U1393 (N_1393,In_222,In_992);
nand U1394 (N_1394,In_593,In_993);
and U1395 (N_1395,In_54,In_913);
nand U1396 (N_1396,In_340,In_257);
nand U1397 (N_1397,In_302,In_717);
or U1398 (N_1398,In_973,In_975);
nand U1399 (N_1399,In_577,In_654);
and U1400 (N_1400,In_189,In_164);
nor U1401 (N_1401,In_167,In_911);
xor U1402 (N_1402,In_911,In_665);
and U1403 (N_1403,In_773,In_28);
nor U1404 (N_1404,In_683,In_730);
nand U1405 (N_1405,In_643,In_551);
or U1406 (N_1406,In_125,In_620);
or U1407 (N_1407,In_51,In_281);
nor U1408 (N_1408,In_159,In_151);
or U1409 (N_1409,In_301,In_454);
nor U1410 (N_1410,In_588,In_291);
or U1411 (N_1411,In_760,In_234);
nor U1412 (N_1412,In_731,In_323);
nor U1413 (N_1413,In_974,In_964);
nand U1414 (N_1414,In_916,In_520);
or U1415 (N_1415,In_231,In_111);
and U1416 (N_1416,In_617,In_768);
or U1417 (N_1417,In_393,In_387);
nor U1418 (N_1418,In_237,In_201);
nand U1419 (N_1419,In_212,In_682);
and U1420 (N_1420,In_598,In_948);
or U1421 (N_1421,In_148,In_825);
and U1422 (N_1422,In_26,In_306);
nor U1423 (N_1423,In_367,In_99);
nand U1424 (N_1424,In_308,In_664);
nor U1425 (N_1425,In_7,In_193);
or U1426 (N_1426,In_679,In_237);
nor U1427 (N_1427,In_183,In_466);
nor U1428 (N_1428,In_245,In_580);
and U1429 (N_1429,In_493,In_125);
nand U1430 (N_1430,In_146,In_700);
and U1431 (N_1431,In_119,In_109);
nor U1432 (N_1432,In_215,In_572);
nand U1433 (N_1433,In_941,In_694);
and U1434 (N_1434,In_952,In_16);
xnor U1435 (N_1435,In_39,In_51);
or U1436 (N_1436,In_754,In_37);
nand U1437 (N_1437,In_448,In_653);
nand U1438 (N_1438,In_496,In_489);
or U1439 (N_1439,In_682,In_471);
and U1440 (N_1440,In_994,In_535);
or U1441 (N_1441,In_299,In_951);
and U1442 (N_1442,In_825,In_275);
or U1443 (N_1443,In_327,In_621);
and U1444 (N_1444,In_466,In_84);
or U1445 (N_1445,In_343,In_967);
nand U1446 (N_1446,In_282,In_398);
nor U1447 (N_1447,In_934,In_449);
or U1448 (N_1448,In_485,In_816);
and U1449 (N_1449,In_118,In_413);
nor U1450 (N_1450,In_212,In_24);
nor U1451 (N_1451,In_781,In_834);
nor U1452 (N_1452,In_747,In_760);
nand U1453 (N_1453,In_679,In_411);
nand U1454 (N_1454,In_552,In_916);
nor U1455 (N_1455,In_840,In_956);
and U1456 (N_1456,In_38,In_810);
nor U1457 (N_1457,In_413,In_462);
and U1458 (N_1458,In_889,In_399);
nand U1459 (N_1459,In_143,In_442);
xnor U1460 (N_1460,In_593,In_279);
nor U1461 (N_1461,In_753,In_240);
nor U1462 (N_1462,In_524,In_943);
nand U1463 (N_1463,In_18,In_840);
and U1464 (N_1464,In_91,In_559);
and U1465 (N_1465,In_844,In_887);
nor U1466 (N_1466,In_634,In_181);
or U1467 (N_1467,In_310,In_726);
nand U1468 (N_1468,In_332,In_57);
or U1469 (N_1469,In_105,In_575);
nor U1470 (N_1470,In_99,In_154);
and U1471 (N_1471,In_129,In_393);
nand U1472 (N_1472,In_938,In_360);
nand U1473 (N_1473,In_482,In_926);
or U1474 (N_1474,In_215,In_454);
or U1475 (N_1475,In_672,In_451);
nor U1476 (N_1476,In_542,In_443);
nand U1477 (N_1477,In_393,In_479);
or U1478 (N_1478,In_980,In_868);
nand U1479 (N_1479,In_8,In_31);
nor U1480 (N_1480,In_521,In_972);
and U1481 (N_1481,In_329,In_356);
nor U1482 (N_1482,In_623,In_99);
and U1483 (N_1483,In_965,In_636);
or U1484 (N_1484,In_63,In_117);
nor U1485 (N_1485,In_856,In_190);
nor U1486 (N_1486,In_756,In_574);
and U1487 (N_1487,In_390,In_385);
or U1488 (N_1488,In_593,In_461);
or U1489 (N_1489,In_20,In_138);
and U1490 (N_1490,In_389,In_855);
or U1491 (N_1491,In_854,In_307);
or U1492 (N_1492,In_707,In_857);
nor U1493 (N_1493,In_864,In_269);
nand U1494 (N_1494,In_17,In_40);
and U1495 (N_1495,In_684,In_677);
or U1496 (N_1496,In_104,In_637);
nand U1497 (N_1497,In_806,In_520);
and U1498 (N_1498,In_922,In_317);
or U1499 (N_1499,In_862,In_605);
or U1500 (N_1500,In_592,In_637);
nor U1501 (N_1501,In_300,In_440);
or U1502 (N_1502,In_274,In_588);
nor U1503 (N_1503,In_99,In_634);
nand U1504 (N_1504,In_153,In_328);
nand U1505 (N_1505,In_526,In_233);
nor U1506 (N_1506,In_539,In_550);
nand U1507 (N_1507,In_878,In_46);
nor U1508 (N_1508,In_916,In_925);
nor U1509 (N_1509,In_27,In_226);
or U1510 (N_1510,In_508,In_247);
or U1511 (N_1511,In_454,In_879);
nand U1512 (N_1512,In_777,In_953);
nor U1513 (N_1513,In_851,In_948);
or U1514 (N_1514,In_495,In_935);
and U1515 (N_1515,In_767,In_280);
and U1516 (N_1516,In_251,In_199);
and U1517 (N_1517,In_854,In_39);
nand U1518 (N_1518,In_693,In_642);
nor U1519 (N_1519,In_419,In_503);
and U1520 (N_1520,In_430,In_818);
and U1521 (N_1521,In_223,In_985);
and U1522 (N_1522,In_511,In_177);
and U1523 (N_1523,In_886,In_147);
nand U1524 (N_1524,In_889,In_85);
or U1525 (N_1525,In_193,In_307);
nand U1526 (N_1526,In_31,In_206);
or U1527 (N_1527,In_442,In_953);
and U1528 (N_1528,In_105,In_124);
or U1529 (N_1529,In_632,In_861);
or U1530 (N_1530,In_582,In_207);
nor U1531 (N_1531,In_850,In_472);
nor U1532 (N_1532,In_438,In_49);
or U1533 (N_1533,In_473,In_112);
or U1534 (N_1534,In_716,In_832);
nor U1535 (N_1535,In_826,In_528);
nor U1536 (N_1536,In_248,In_820);
nor U1537 (N_1537,In_181,In_641);
or U1538 (N_1538,In_168,In_125);
nand U1539 (N_1539,In_320,In_356);
and U1540 (N_1540,In_508,In_746);
and U1541 (N_1541,In_257,In_419);
or U1542 (N_1542,In_192,In_560);
nor U1543 (N_1543,In_191,In_851);
nand U1544 (N_1544,In_764,In_130);
nor U1545 (N_1545,In_829,In_128);
nor U1546 (N_1546,In_857,In_235);
nor U1547 (N_1547,In_104,In_185);
nor U1548 (N_1548,In_383,In_797);
nand U1549 (N_1549,In_682,In_686);
nor U1550 (N_1550,In_604,In_213);
and U1551 (N_1551,In_330,In_998);
xnor U1552 (N_1552,In_511,In_869);
nand U1553 (N_1553,In_513,In_650);
nor U1554 (N_1554,In_269,In_287);
nand U1555 (N_1555,In_457,In_542);
nor U1556 (N_1556,In_889,In_718);
and U1557 (N_1557,In_476,In_197);
or U1558 (N_1558,In_668,In_235);
or U1559 (N_1559,In_678,In_160);
nand U1560 (N_1560,In_28,In_712);
and U1561 (N_1561,In_597,In_134);
or U1562 (N_1562,In_986,In_764);
nand U1563 (N_1563,In_8,In_839);
nor U1564 (N_1564,In_5,In_934);
and U1565 (N_1565,In_977,In_413);
nand U1566 (N_1566,In_155,In_214);
and U1567 (N_1567,In_266,In_601);
nand U1568 (N_1568,In_30,In_715);
nand U1569 (N_1569,In_273,In_628);
nand U1570 (N_1570,In_82,In_81);
or U1571 (N_1571,In_151,In_147);
nand U1572 (N_1572,In_707,In_344);
nand U1573 (N_1573,In_862,In_832);
nor U1574 (N_1574,In_658,In_897);
or U1575 (N_1575,In_389,In_813);
nor U1576 (N_1576,In_473,In_680);
nor U1577 (N_1577,In_348,In_147);
and U1578 (N_1578,In_311,In_338);
and U1579 (N_1579,In_147,In_927);
or U1580 (N_1580,In_66,In_384);
or U1581 (N_1581,In_66,In_616);
nand U1582 (N_1582,In_783,In_892);
or U1583 (N_1583,In_181,In_242);
and U1584 (N_1584,In_396,In_82);
or U1585 (N_1585,In_305,In_852);
and U1586 (N_1586,In_612,In_971);
nor U1587 (N_1587,In_424,In_379);
and U1588 (N_1588,In_333,In_166);
nand U1589 (N_1589,In_19,In_754);
and U1590 (N_1590,In_534,In_766);
and U1591 (N_1591,In_370,In_927);
nor U1592 (N_1592,In_576,In_647);
nor U1593 (N_1593,In_589,In_421);
and U1594 (N_1594,In_826,In_738);
nor U1595 (N_1595,In_632,In_423);
or U1596 (N_1596,In_78,In_261);
and U1597 (N_1597,In_583,In_712);
or U1598 (N_1598,In_967,In_914);
or U1599 (N_1599,In_562,In_168);
xnor U1600 (N_1600,In_934,In_910);
or U1601 (N_1601,In_509,In_315);
nor U1602 (N_1602,In_514,In_215);
and U1603 (N_1603,In_452,In_991);
or U1604 (N_1604,In_229,In_887);
nand U1605 (N_1605,In_820,In_478);
nand U1606 (N_1606,In_728,In_156);
nand U1607 (N_1607,In_599,In_389);
or U1608 (N_1608,In_968,In_726);
nand U1609 (N_1609,In_166,In_298);
nor U1610 (N_1610,In_680,In_664);
nor U1611 (N_1611,In_647,In_962);
or U1612 (N_1612,In_97,In_668);
nor U1613 (N_1613,In_656,In_582);
nand U1614 (N_1614,In_195,In_702);
and U1615 (N_1615,In_708,In_663);
and U1616 (N_1616,In_385,In_491);
and U1617 (N_1617,In_344,In_847);
xor U1618 (N_1618,In_85,In_640);
nand U1619 (N_1619,In_437,In_852);
or U1620 (N_1620,In_957,In_645);
and U1621 (N_1621,In_308,In_820);
nor U1622 (N_1622,In_195,In_745);
nor U1623 (N_1623,In_890,In_2);
nor U1624 (N_1624,In_103,In_222);
nand U1625 (N_1625,In_449,In_300);
or U1626 (N_1626,In_632,In_999);
nor U1627 (N_1627,In_984,In_324);
or U1628 (N_1628,In_759,In_942);
and U1629 (N_1629,In_252,In_422);
or U1630 (N_1630,In_417,In_285);
and U1631 (N_1631,In_69,In_656);
xnor U1632 (N_1632,In_303,In_327);
and U1633 (N_1633,In_8,In_445);
and U1634 (N_1634,In_129,In_973);
and U1635 (N_1635,In_34,In_648);
and U1636 (N_1636,In_499,In_962);
nor U1637 (N_1637,In_518,In_467);
or U1638 (N_1638,In_812,In_137);
or U1639 (N_1639,In_535,In_899);
and U1640 (N_1640,In_855,In_256);
nand U1641 (N_1641,In_992,In_354);
nand U1642 (N_1642,In_277,In_504);
nor U1643 (N_1643,In_969,In_115);
nor U1644 (N_1644,In_57,In_618);
nand U1645 (N_1645,In_465,In_494);
xnor U1646 (N_1646,In_8,In_848);
nand U1647 (N_1647,In_790,In_139);
or U1648 (N_1648,In_330,In_568);
nor U1649 (N_1649,In_369,In_871);
nand U1650 (N_1650,In_574,In_60);
nor U1651 (N_1651,In_422,In_743);
or U1652 (N_1652,In_263,In_308);
and U1653 (N_1653,In_999,In_321);
nand U1654 (N_1654,In_82,In_402);
nor U1655 (N_1655,In_225,In_554);
or U1656 (N_1656,In_675,In_18);
and U1657 (N_1657,In_611,In_920);
nand U1658 (N_1658,In_461,In_711);
nand U1659 (N_1659,In_166,In_769);
xnor U1660 (N_1660,In_10,In_996);
or U1661 (N_1661,In_109,In_625);
nand U1662 (N_1662,In_267,In_811);
nor U1663 (N_1663,In_115,In_647);
xnor U1664 (N_1664,In_349,In_525);
or U1665 (N_1665,In_7,In_524);
or U1666 (N_1666,In_834,In_268);
nand U1667 (N_1667,In_247,In_51);
nor U1668 (N_1668,In_604,In_580);
and U1669 (N_1669,In_346,In_510);
nand U1670 (N_1670,In_217,In_137);
or U1671 (N_1671,In_439,In_462);
and U1672 (N_1672,In_909,In_984);
nor U1673 (N_1673,In_841,In_843);
or U1674 (N_1674,In_763,In_784);
or U1675 (N_1675,In_617,In_840);
nor U1676 (N_1676,In_203,In_156);
nor U1677 (N_1677,In_154,In_815);
nand U1678 (N_1678,In_513,In_317);
nor U1679 (N_1679,In_539,In_447);
nor U1680 (N_1680,In_162,In_238);
nand U1681 (N_1681,In_407,In_616);
xor U1682 (N_1682,In_986,In_923);
nand U1683 (N_1683,In_371,In_99);
nor U1684 (N_1684,In_766,In_42);
xnor U1685 (N_1685,In_835,In_902);
and U1686 (N_1686,In_461,In_473);
nand U1687 (N_1687,In_25,In_868);
nand U1688 (N_1688,In_828,In_54);
nor U1689 (N_1689,In_315,In_491);
or U1690 (N_1690,In_604,In_882);
nand U1691 (N_1691,In_827,In_323);
nor U1692 (N_1692,In_342,In_715);
nand U1693 (N_1693,In_129,In_242);
nand U1694 (N_1694,In_422,In_563);
nand U1695 (N_1695,In_715,In_84);
or U1696 (N_1696,In_230,In_767);
nand U1697 (N_1697,In_332,In_265);
and U1698 (N_1698,In_605,In_74);
and U1699 (N_1699,In_786,In_722);
or U1700 (N_1700,In_161,In_141);
and U1701 (N_1701,In_345,In_116);
and U1702 (N_1702,In_850,In_177);
nor U1703 (N_1703,In_928,In_887);
nor U1704 (N_1704,In_709,In_834);
or U1705 (N_1705,In_166,In_152);
or U1706 (N_1706,In_477,In_75);
and U1707 (N_1707,In_30,In_285);
nand U1708 (N_1708,In_708,In_966);
and U1709 (N_1709,In_31,In_53);
or U1710 (N_1710,In_196,In_367);
or U1711 (N_1711,In_529,In_823);
nor U1712 (N_1712,In_998,In_431);
and U1713 (N_1713,In_103,In_297);
or U1714 (N_1714,In_826,In_165);
or U1715 (N_1715,In_189,In_99);
and U1716 (N_1716,In_479,In_639);
nor U1717 (N_1717,In_703,In_323);
nand U1718 (N_1718,In_385,In_270);
and U1719 (N_1719,In_777,In_37);
xnor U1720 (N_1720,In_884,In_450);
and U1721 (N_1721,In_98,In_151);
nor U1722 (N_1722,In_544,In_165);
and U1723 (N_1723,In_821,In_60);
or U1724 (N_1724,In_973,In_447);
nand U1725 (N_1725,In_303,In_174);
and U1726 (N_1726,In_217,In_481);
nor U1727 (N_1727,In_24,In_743);
nand U1728 (N_1728,In_423,In_520);
nor U1729 (N_1729,In_424,In_658);
and U1730 (N_1730,In_136,In_933);
or U1731 (N_1731,In_719,In_263);
nand U1732 (N_1732,In_929,In_974);
and U1733 (N_1733,In_229,In_523);
and U1734 (N_1734,In_909,In_60);
nand U1735 (N_1735,In_400,In_853);
nand U1736 (N_1736,In_463,In_385);
nor U1737 (N_1737,In_576,In_934);
or U1738 (N_1738,In_72,In_690);
and U1739 (N_1739,In_831,In_578);
and U1740 (N_1740,In_978,In_115);
or U1741 (N_1741,In_196,In_854);
and U1742 (N_1742,In_391,In_586);
nand U1743 (N_1743,In_75,In_634);
nand U1744 (N_1744,In_522,In_245);
and U1745 (N_1745,In_9,In_227);
nand U1746 (N_1746,In_6,In_979);
nor U1747 (N_1747,In_953,In_707);
nor U1748 (N_1748,In_256,In_122);
nor U1749 (N_1749,In_12,In_896);
nand U1750 (N_1750,In_494,In_51);
nor U1751 (N_1751,In_7,In_914);
nand U1752 (N_1752,In_840,In_161);
nand U1753 (N_1753,In_937,In_701);
or U1754 (N_1754,In_103,In_182);
and U1755 (N_1755,In_932,In_318);
nor U1756 (N_1756,In_282,In_991);
and U1757 (N_1757,In_697,In_708);
nor U1758 (N_1758,In_639,In_831);
or U1759 (N_1759,In_438,In_986);
or U1760 (N_1760,In_488,In_738);
nor U1761 (N_1761,In_67,In_537);
and U1762 (N_1762,In_877,In_181);
or U1763 (N_1763,In_936,In_94);
nor U1764 (N_1764,In_720,In_599);
and U1765 (N_1765,In_396,In_225);
nor U1766 (N_1766,In_709,In_125);
nand U1767 (N_1767,In_401,In_780);
nand U1768 (N_1768,In_342,In_26);
or U1769 (N_1769,In_834,In_459);
or U1770 (N_1770,In_699,In_506);
or U1771 (N_1771,In_933,In_373);
and U1772 (N_1772,In_639,In_394);
nand U1773 (N_1773,In_913,In_447);
or U1774 (N_1774,In_690,In_579);
and U1775 (N_1775,In_220,In_967);
nor U1776 (N_1776,In_453,In_978);
nor U1777 (N_1777,In_932,In_27);
nand U1778 (N_1778,In_579,In_210);
or U1779 (N_1779,In_35,In_585);
and U1780 (N_1780,In_325,In_739);
nor U1781 (N_1781,In_996,In_401);
or U1782 (N_1782,In_44,In_861);
and U1783 (N_1783,In_883,In_244);
nor U1784 (N_1784,In_712,In_333);
nor U1785 (N_1785,In_773,In_885);
or U1786 (N_1786,In_534,In_54);
nor U1787 (N_1787,In_120,In_73);
or U1788 (N_1788,In_172,In_954);
nor U1789 (N_1789,In_101,In_527);
or U1790 (N_1790,In_465,In_649);
and U1791 (N_1791,In_582,In_733);
nor U1792 (N_1792,In_429,In_589);
nor U1793 (N_1793,In_982,In_323);
and U1794 (N_1794,In_403,In_366);
and U1795 (N_1795,In_249,In_374);
nand U1796 (N_1796,In_891,In_615);
and U1797 (N_1797,In_687,In_250);
nor U1798 (N_1798,In_33,In_596);
or U1799 (N_1799,In_96,In_793);
or U1800 (N_1800,In_874,In_914);
and U1801 (N_1801,In_87,In_814);
nor U1802 (N_1802,In_598,In_436);
and U1803 (N_1803,In_797,In_530);
and U1804 (N_1804,In_126,In_936);
nand U1805 (N_1805,In_25,In_372);
and U1806 (N_1806,In_911,In_32);
nor U1807 (N_1807,In_850,In_828);
nor U1808 (N_1808,In_809,In_854);
nor U1809 (N_1809,In_520,In_591);
nand U1810 (N_1810,In_304,In_823);
or U1811 (N_1811,In_271,In_168);
nor U1812 (N_1812,In_395,In_951);
or U1813 (N_1813,In_88,In_470);
nand U1814 (N_1814,In_862,In_278);
or U1815 (N_1815,In_94,In_46);
and U1816 (N_1816,In_815,In_473);
xnor U1817 (N_1817,In_773,In_827);
or U1818 (N_1818,In_487,In_516);
and U1819 (N_1819,In_470,In_789);
nor U1820 (N_1820,In_196,In_412);
and U1821 (N_1821,In_338,In_758);
and U1822 (N_1822,In_27,In_949);
nand U1823 (N_1823,In_975,In_394);
nor U1824 (N_1824,In_442,In_376);
nor U1825 (N_1825,In_473,In_41);
or U1826 (N_1826,In_983,In_389);
or U1827 (N_1827,In_199,In_847);
nand U1828 (N_1828,In_841,In_248);
nor U1829 (N_1829,In_600,In_548);
and U1830 (N_1830,In_564,In_686);
and U1831 (N_1831,In_629,In_245);
or U1832 (N_1832,In_753,In_376);
nor U1833 (N_1833,In_528,In_626);
nor U1834 (N_1834,In_856,In_767);
nand U1835 (N_1835,In_821,In_615);
nor U1836 (N_1836,In_871,In_474);
or U1837 (N_1837,In_724,In_386);
nand U1838 (N_1838,In_966,In_453);
or U1839 (N_1839,In_232,In_294);
nand U1840 (N_1840,In_541,In_166);
or U1841 (N_1841,In_682,In_492);
and U1842 (N_1842,In_799,In_105);
nand U1843 (N_1843,In_597,In_636);
or U1844 (N_1844,In_643,In_736);
and U1845 (N_1845,In_581,In_514);
nand U1846 (N_1846,In_59,In_206);
nor U1847 (N_1847,In_941,In_759);
nand U1848 (N_1848,In_644,In_686);
nor U1849 (N_1849,In_55,In_210);
nor U1850 (N_1850,In_23,In_19);
nor U1851 (N_1851,In_523,In_969);
nor U1852 (N_1852,In_963,In_139);
nor U1853 (N_1853,In_890,In_107);
or U1854 (N_1854,In_626,In_111);
and U1855 (N_1855,In_90,In_884);
and U1856 (N_1856,In_669,In_107);
and U1857 (N_1857,In_604,In_215);
nand U1858 (N_1858,In_440,In_26);
nor U1859 (N_1859,In_638,In_770);
nand U1860 (N_1860,In_366,In_443);
and U1861 (N_1861,In_208,In_475);
or U1862 (N_1862,In_581,In_120);
and U1863 (N_1863,In_541,In_114);
and U1864 (N_1864,In_947,In_486);
nand U1865 (N_1865,In_264,In_424);
or U1866 (N_1866,In_87,In_742);
nor U1867 (N_1867,In_547,In_843);
nand U1868 (N_1868,In_380,In_573);
nor U1869 (N_1869,In_714,In_828);
or U1870 (N_1870,In_845,In_566);
nor U1871 (N_1871,In_605,In_999);
nand U1872 (N_1872,In_541,In_262);
and U1873 (N_1873,In_652,In_911);
nand U1874 (N_1874,In_367,In_827);
and U1875 (N_1875,In_599,In_675);
or U1876 (N_1876,In_421,In_263);
or U1877 (N_1877,In_458,In_795);
nand U1878 (N_1878,In_727,In_520);
and U1879 (N_1879,In_863,In_346);
or U1880 (N_1880,In_208,In_676);
nand U1881 (N_1881,In_733,In_453);
or U1882 (N_1882,In_427,In_690);
nand U1883 (N_1883,In_519,In_798);
nor U1884 (N_1884,In_889,In_818);
or U1885 (N_1885,In_821,In_552);
nor U1886 (N_1886,In_486,In_857);
or U1887 (N_1887,In_750,In_658);
nor U1888 (N_1888,In_377,In_430);
nor U1889 (N_1889,In_659,In_7);
nor U1890 (N_1890,In_13,In_387);
and U1891 (N_1891,In_550,In_715);
nand U1892 (N_1892,In_991,In_76);
nor U1893 (N_1893,In_821,In_703);
nor U1894 (N_1894,In_30,In_854);
nor U1895 (N_1895,In_610,In_964);
nand U1896 (N_1896,In_146,In_965);
or U1897 (N_1897,In_866,In_697);
nand U1898 (N_1898,In_247,In_324);
and U1899 (N_1899,In_675,In_484);
or U1900 (N_1900,In_795,In_740);
or U1901 (N_1901,In_605,In_609);
or U1902 (N_1902,In_666,In_837);
or U1903 (N_1903,In_210,In_90);
and U1904 (N_1904,In_678,In_596);
nand U1905 (N_1905,In_575,In_164);
nand U1906 (N_1906,In_531,In_422);
nor U1907 (N_1907,In_919,In_837);
nor U1908 (N_1908,In_693,In_23);
or U1909 (N_1909,In_319,In_879);
or U1910 (N_1910,In_732,In_65);
nand U1911 (N_1911,In_363,In_344);
nor U1912 (N_1912,In_753,In_559);
or U1913 (N_1913,In_875,In_244);
nor U1914 (N_1914,In_686,In_643);
and U1915 (N_1915,In_43,In_153);
or U1916 (N_1916,In_960,In_692);
nand U1917 (N_1917,In_516,In_127);
and U1918 (N_1918,In_337,In_130);
nand U1919 (N_1919,In_782,In_469);
and U1920 (N_1920,In_623,In_786);
and U1921 (N_1921,In_176,In_840);
nor U1922 (N_1922,In_83,In_268);
or U1923 (N_1923,In_512,In_119);
and U1924 (N_1924,In_769,In_659);
nand U1925 (N_1925,In_114,In_836);
or U1926 (N_1926,In_68,In_904);
and U1927 (N_1927,In_849,In_236);
nand U1928 (N_1928,In_45,In_217);
nor U1929 (N_1929,In_858,In_712);
or U1930 (N_1930,In_801,In_965);
and U1931 (N_1931,In_832,In_931);
nor U1932 (N_1932,In_601,In_800);
or U1933 (N_1933,In_501,In_592);
or U1934 (N_1934,In_583,In_627);
nand U1935 (N_1935,In_990,In_531);
nor U1936 (N_1936,In_573,In_127);
nand U1937 (N_1937,In_331,In_684);
or U1938 (N_1938,In_302,In_753);
or U1939 (N_1939,In_971,In_393);
nor U1940 (N_1940,In_180,In_708);
and U1941 (N_1941,In_387,In_133);
and U1942 (N_1942,In_424,In_810);
nor U1943 (N_1943,In_764,In_258);
or U1944 (N_1944,In_779,In_74);
and U1945 (N_1945,In_995,In_397);
nor U1946 (N_1946,In_157,In_887);
or U1947 (N_1947,In_483,In_985);
or U1948 (N_1948,In_5,In_307);
or U1949 (N_1949,In_583,In_944);
or U1950 (N_1950,In_343,In_585);
or U1951 (N_1951,In_238,In_272);
nor U1952 (N_1952,In_824,In_789);
or U1953 (N_1953,In_876,In_247);
nand U1954 (N_1954,In_883,In_213);
and U1955 (N_1955,In_68,In_707);
or U1956 (N_1956,In_545,In_385);
or U1957 (N_1957,In_520,In_272);
and U1958 (N_1958,In_51,In_262);
and U1959 (N_1959,In_973,In_549);
or U1960 (N_1960,In_434,In_138);
nand U1961 (N_1961,In_978,In_348);
and U1962 (N_1962,In_546,In_560);
and U1963 (N_1963,In_463,In_453);
nand U1964 (N_1964,In_109,In_430);
or U1965 (N_1965,In_965,In_289);
and U1966 (N_1966,In_774,In_332);
nand U1967 (N_1967,In_895,In_868);
nand U1968 (N_1968,In_162,In_775);
nor U1969 (N_1969,In_720,In_371);
nand U1970 (N_1970,In_645,In_170);
nor U1971 (N_1971,In_642,In_563);
nand U1972 (N_1972,In_787,In_412);
nor U1973 (N_1973,In_415,In_107);
or U1974 (N_1974,In_905,In_197);
and U1975 (N_1975,In_409,In_365);
and U1976 (N_1976,In_876,In_456);
and U1977 (N_1977,In_897,In_354);
nor U1978 (N_1978,In_777,In_551);
or U1979 (N_1979,In_286,In_866);
xor U1980 (N_1980,In_260,In_77);
nand U1981 (N_1981,In_100,In_590);
and U1982 (N_1982,In_169,In_812);
nor U1983 (N_1983,In_89,In_519);
nor U1984 (N_1984,In_299,In_509);
nor U1985 (N_1985,In_445,In_680);
nor U1986 (N_1986,In_450,In_930);
nor U1987 (N_1987,In_387,In_124);
or U1988 (N_1988,In_234,In_262);
and U1989 (N_1989,In_377,In_341);
nand U1990 (N_1990,In_322,In_614);
and U1991 (N_1991,In_421,In_867);
or U1992 (N_1992,In_233,In_549);
or U1993 (N_1993,In_182,In_863);
nand U1994 (N_1994,In_729,In_812);
or U1995 (N_1995,In_352,In_651);
or U1996 (N_1996,In_829,In_737);
and U1997 (N_1997,In_213,In_700);
or U1998 (N_1998,In_451,In_331);
or U1999 (N_1999,In_102,In_799);
nor U2000 (N_2000,In_18,In_516);
nor U2001 (N_2001,In_287,In_993);
or U2002 (N_2002,In_187,In_290);
nor U2003 (N_2003,In_635,In_334);
nand U2004 (N_2004,In_730,In_623);
nand U2005 (N_2005,In_741,In_893);
nor U2006 (N_2006,In_356,In_371);
nor U2007 (N_2007,In_336,In_839);
or U2008 (N_2008,In_205,In_671);
nor U2009 (N_2009,In_313,In_721);
nand U2010 (N_2010,In_799,In_468);
and U2011 (N_2011,In_159,In_221);
or U2012 (N_2012,In_694,In_45);
nor U2013 (N_2013,In_898,In_558);
nor U2014 (N_2014,In_354,In_228);
nor U2015 (N_2015,In_382,In_412);
and U2016 (N_2016,In_287,In_320);
and U2017 (N_2017,In_175,In_134);
nor U2018 (N_2018,In_182,In_429);
nor U2019 (N_2019,In_401,In_689);
or U2020 (N_2020,In_870,In_292);
or U2021 (N_2021,In_435,In_456);
nor U2022 (N_2022,In_716,In_928);
and U2023 (N_2023,In_738,In_778);
nor U2024 (N_2024,In_819,In_225);
nor U2025 (N_2025,In_96,In_313);
or U2026 (N_2026,In_663,In_210);
or U2027 (N_2027,In_130,In_922);
or U2028 (N_2028,In_921,In_572);
nand U2029 (N_2029,In_298,In_10);
nand U2030 (N_2030,In_498,In_471);
or U2031 (N_2031,In_282,In_490);
nand U2032 (N_2032,In_901,In_964);
or U2033 (N_2033,In_803,In_421);
and U2034 (N_2034,In_167,In_163);
or U2035 (N_2035,In_893,In_537);
xor U2036 (N_2036,In_328,In_392);
nor U2037 (N_2037,In_969,In_947);
nor U2038 (N_2038,In_687,In_599);
or U2039 (N_2039,In_495,In_168);
xnor U2040 (N_2040,In_25,In_725);
nor U2041 (N_2041,In_214,In_128);
nand U2042 (N_2042,In_573,In_625);
and U2043 (N_2043,In_68,In_123);
and U2044 (N_2044,In_967,In_953);
or U2045 (N_2045,In_981,In_350);
nor U2046 (N_2046,In_271,In_95);
and U2047 (N_2047,In_965,In_67);
or U2048 (N_2048,In_676,In_129);
and U2049 (N_2049,In_825,In_399);
xnor U2050 (N_2050,In_772,In_785);
nand U2051 (N_2051,In_805,In_313);
and U2052 (N_2052,In_531,In_527);
or U2053 (N_2053,In_161,In_366);
nand U2054 (N_2054,In_505,In_926);
nor U2055 (N_2055,In_37,In_136);
nor U2056 (N_2056,In_322,In_714);
or U2057 (N_2057,In_6,In_437);
nand U2058 (N_2058,In_472,In_841);
nor U2059 (N_2059,In_548,In_623);
and U2060 (N_2060,In_717,In_556);
nor U2061 (N_2061,In_383,In_459);
and U2062 (N_2062,In_73,In_186);
nor U2063 (N_2063,In_234,In_206);
or U2064 (N_2064,In_303,In_794);
nor U2065 (N_2065,In_527,In_255);
nor U2066 (N_2066,In_654,In_80);
or U2067 (N_2067,In_342,In_918);
or U2068 (N_2068,In_275,In_342);
and U2069 (N_2069,In_542,In_632);
nor U2070 (N_2070,In_203,In_849);
and U2071 (N_2071,In_700,In_954);
nand U2072 (N_2072,In_861,In_331);
or U2073 (N_2073,In_240,In_497);
nand U2074 (N_2074,In_659,In_968);
nand U2075 (N_2075,In_333,In_520);
nor U2076 (N_2076,In_228,In_451);
nand U2077 (N_2077,In_553,In_515);
or U2078 (N_2078,In_276,In_673);
or U2079 (N_2079,In_31,In_118);
or U2080 (N_2080,In_944,In_691);
and U2081 (N_2081,In_389,In_616);
nand U2082 (N_2082,In_688,In_786);
nand U2083 (N_2083,In_216,In_485);
or U2084 (N_2084,In_493,In_398);
nand U2085 (N_2085,In_741,In_163);
or U2086 (N_2086,In_114,In_969);
or U2087 (N_2087,In_696,In_151);
and U2088 (N_2088,In_114,In_743);
nand U2089 (N_2089,In_162,In_102);
nand U2090 (N_2090,In_745,In_645);
nor U2091 (N_2091,In_782,In_976);
or U2092 (N_2092,In_625,In_651);
or U2093 (N_2093,In_726,In_101);
nor U2094 (N_2094,In_387,In_509);
or U2095 (N_2095,In_841,In_193);
nand U2096 (N_2096,In_629,In_739);
and U2097 (N_2097,In_125,In_440);
nor U2098 (N_2098,In_531,In_932);
and U2099 (N_2099,In_753,In_572);
nor U2100 (N_2100,In_170,In_71);
or U2101 (N_2101,In_726,In_542);
or U2102 (N_2102,In_199,In_272);
nor U2103 (N_2103,In_378,In_835);
or U2104 (N_2104,In_773,In_858);
or U2105 (N_2105,In_921,In_384);
nand U2106 (N_2106,In_85,In_44);
or U2107 (N_2107,In_315,In_918);
and U2108 (N_2108,In_926,In_370);
nor U2109 (N_2109,In_423,In_815);
and U2110 (N_2110,In_820,In_399);
nand U2111 (N_2111,In_353,In_373);
and U2112 (N_2112,In_537,In_510);
xor U2113 (N_2113,In_989,In_112);
or U2114 (N_2114,In_152,In_597);
or U2115 (N_2115,In_971,In_11);
nand U2116 (N_2116,In_279,In_750);
xor U2117 (N_2117,In_757,In_878);
and U2118 (N_2118,In_758,In_106);
and U2119 (N_2119,In_44,In_624);
and U2120 (N_2120,In_369,In_539);
and U2121 (N_2121,In_27,In_348);
nor U2122 (N_2122,In_711,In_944);
or U2123 (N_2123,In_186,In_924);
and U2124 (N_2124,In_343,In_78);
and U2125 (N_2125,In_659,In_352);
or U2126 (N_2126,In_806,In_696);
and U2127 (N_2127,In_497,In_416);
xor U2128 (N_2128,In_697,In_497);
or U2129 (N_2129,In_479,In_79);
nor U2130 (N_2130,In_153,In_776);
or U2131 (N_2131,In_455,In_410);
nand U2132 (N_2132,In_149,In_87);
or U2133 (N_2133,In_777,In_511);
nor U2134 (N_2134,In_753,In_828);
nor U2135 (N_2135,In_585,In_402);
nor U2136 (N_2136,In_391,In_115);
nand U2137 (N_2137,In_365,In_494);
and U2138 (N_2138,In_806,In_238);
nand U2139 (N_2139,In_617,In_786);
and U2140 (N_2140,In_719,In_420);
nand U2141 (N_2141,In_37,In_436);
nand U2142 (N_2142,In_859,In_208);
nand U2143 (N_2143,In_781,In_96);
nand U2144 (N_2144,In_855,In_950);
nor U2145 (N_2145,In_935,In_984);
nand U2146 (N_2146,In_502,In_840);
nor U2147 (N_2147,In_467,In_966);
and U2148 (N_2148,In_79,In_746);
nor U2149 (N_2149,In_197,In_955);
nand U2150 (N_2150,In_100,In_284);
xor U2151 (N_2151,In_696,In_322);
xnor U2152 (N_2152,In_972,In_588);
and U2153 (N_2153,In_752,In_623);
nor U2154 (N_2154,In_346,In_672);
and U2155 (N_2155,In_312,In_693);
and U2156 (N_2156,In_832,In_306);
or U2157 (N_2157,In_448,In_860);
nor U2158 (N_2158,In_441,In_86);
nor U2159 (N_2159,In_446,In_858);
nand U2160 (N_2160,In_885,In_942);
nor U2161 (N_2161,In_823,In_382);
nor U2162 (N_2162,In_14,In_799);
nor U2163 (N_2163,In_530,In_194);
nand U2164 (N_2164,In_142,In_211);
or U2165 (N_2165,In_705,In_167);
nor U2166 (N_2166,In_197,In_614);
nor U2167 (N_2167,In_465,In_613);
or U2168 (N_2168,In_166,In_537);
or U2169 (N_2169,In_119,In_11);
or U2170 (N_2170,In_991,In_631);
and U2171 (N_2171,In_629,In_147);
and U2172 (N_2172,In_258,In_273);
nor U2173 (N_2173,In_879,In_89);
and U2174 (N_2174,In_505,In_873);
nor U2175 (N_2175,In_488,In_777);
or U2176 (N_2176,In_966,In_488);
or U2177 (N_2177,In_479,In_82);
and U2178 (N_2178,In_77,In_512);
or U2179 (N_2179,In_264,In_861);
nor U2180 (N_2180,In_299,In_89);
nor U2181 (N_2181,In_972,In_971);
and U2182 (N_2182,In_598,In_271);
and U2183 (N_2183,In_232,In_464);
and U2184 (N_2184,In_141,In_167);
and U2185 (N_2185,In_878,In_846);
nor U2186 (N_2186,In_675,In_578);
nand U2187 (N_2187,In_618,In_368);
and U2188 (N_2188,In_687,In_605);
and U2189 (N_2189,In_636,In_337);
nand U2190 (N_2190,In_430,In_869);
or U2191 (N_2191,In_542,In_765);
or U2192 (N_2192,In_845,In_711);
and U2193 (N_2193,In_352,In_730);
and U2194 (N_2194,In_819,In_588);
nor U2195 (N_2195,In_463,In_533);
nor U2196 (N_2196,In_210,In_380);
nor U2197 (N_2197,In_166,In_98);
or U2198 (N_2198,In_654,In_805);
nor U2199 (N_2199,In_489,In_946);
nand U2200 (N_2200,In_741,In_424);
and U2201 (N_2201,In_14,In_209);
and U2202 (N_2202,In_126,In_878);
and U2203 (N_2203,In_549,In_977);
nand U2204 (N_2204,In_225,In_298);
and U2205 (N_2205,In_171,In_283);
nand U2206 (N_2206,In_586,In_576);
nand U2207 (N_2207,In_61,In_732);
or U2208 (N_2208,In_339,In_569);
or U2209 (N_2209,In_271,In_453);
nor U2210 (N_2210,In_929,In_150);
nor U2211 (N_2211,In_542,In_943);
and U2212 (N_2212,In_840,In_511);
and U2213 (N_2213,In_418,In_48);
and U2214 (N_2214,In_925,In_802);
or U2215 (N_2215,In_658,In_678);
nor U2216 (N_2216,In_690,In_555);
nor U2217 (N_2217,In_659,In_354);
or U2218 (N_2218,In_789,In_606);
and U2219 (N_2219,In_72,In_637);
nand U2220 (N_2220,In_920,In_934);
nand U2221 (N_2221,In_985,In_970);
or U2222 (N_2222,In_603,In_899);
nor U2223 (N_2223,In_955,In_727);
nor U2224 (N_2224,In_629,In_654);
nand U2225 (N_2225,In_754,In_207);
nand U2226 (N_2226,In_129,In_383);
nor U2227 (N_2227,In_191,In_460);
nand U2228 (N_2228,In_330,In_417);
or U2229 (N_2229,In_116,In_441);
or U2230 (N_2230,In_469,In_84);
nand U2231 (N_2231,In_199,In_912);
and U2232 (N_2232,In_85,In_896);
nand U2233 (N_2233,In_238,In_566);
and U2234 (N_2234,In_369,In_80);
nand U2235 (N_2235,In_999,In_416);
nor U2236 (N_2236,In_369,In_508);
or U2237 (N_2237,In_711,In_908);
or U2238 (N_2238,In_613,In_230);
and U2239 (N_2239,In_663,In_609);
or U2240 (N_2240,In_621,In_425);
and U2241 (N_2241,In_647,In_545);
nor U2242 (N_2242,In_286,In_354);
nor U2243 (N_2243,In_119,In_587);
and U2244 (N_2244,In_432,In_703);
or U2245 (N_2245,In_575,In_919);
nor U2246 (N_2246,In_966,In_764);
nor U2247 (N_2247,In_743,In_38);
nand U2248 (N_2248,In_436,In_911);
or U2249 (N_2249,In_397,In_422);
and U2250 (N_2250,In_622,In_179);
and U2251 (N_2251,In_984,In_171);
and U2252 (N_2252,In_151,In_536);
xnor U2253 (N_2253,In_58,In_106);
nand U2254 (N_2254,In_404,In_296);
or U2255 (N_2255,In_563,In_120);
nand U2256 (N_2256,In_502,In_662);
or U2257 (N_2257,In_414,In_462);
or U2258 (N_2258,In_778,In_894);
nand U2259 (N_2259,In_237,In_698);
nor U2260 (N_2260,In_306,In_867);
and U2261 (N_2261,In_295,In_431);
and U2262 (N_2262,In_712,In_111);
nor U2263 (N_2263,In_415,In_847);
and U2264 (N_2264,In_845,In_64);
nor U2265 (N_2265,In_184,In_795);
and U2266 (N_2266,In_858,In_635);
and U2267 (N_2267,In_912,In_105);
nor U2268 (N_2268,In_566,In_928);
or U2269 (N_2269,In_995,In_271);
or U2270 (N_2270,In_312,In_330);
or U2271 (N_2271,In_266,In_302);
or U2272 (N_2272,In_89,In_160);
nor U2273 (N_2273,In_869,In_65);
and U2274 (N_2274,In_620,In_385);
nand U2275 (N_2275,In_529,In_385);
nand U2276 (N_2276,In_507,In_486);
or U2277 (N_2277,In_947,In_387);
nand U2278 (N_2278,In_442,In_899);
or U2279 (N_2279,In_90,In_500);
and U2280 (N_2280,In_15,In_459);
and U2281 (N_2281,In_872,In_448);
and U2282 (N_2282,In_287,In_679);
nand U2283 (N_2283,In_447,In_139);
nand U2284 (N_2284,In_257,In_991);
and U2285 (N_2285,In_126,In_103);
or U2286 (N_2286,In_29,In_653);
or U2287 (N_2287,In_615,In_43);
or U2288 (N_2288,In_206,In_9);
and U2289 (N_2289,In_735,In_551);
nand U2290 (N_2290,In_736,In_783);
or U2291 (N_2291,In_711,In_658);
and U2292 (N_2292,In_133,In_846);
nand U2293 (N_2293,In_359,In_836);
nor U2294 (N_2294,In_546,In_190);
and U2295 (N_2295,In_985,In_318);
nand U2296 (N_2296,In_249,In_175);
nand U2297 (N_2297,In_887,In_292);
and U2298 (N_2298,In_423,In_181);
and U2299 (N_2299,In_5,In_677);
nor U2300 (N_2300,In_711,In_611);
and U2301 (N_2301,In_430,In_265);
and U2302 (N_2302,In_329,In_279);
nand U2303 (N_2303,In_662,In_987);
nor U2304 (N_2304,In_533,In_434);
nand U2305 (N_2305,In_861,In_883);
and U2306 (N_2306,In_436,In_641);
nand U2307 (N_2307,In_782,In_435);
nor U2308 (N_2308,In_882,In_699);
and U2309 (N_2309,In_815,In_772);
xnor U2310 (N_2310,In_672,In_408);
or U2311 (N_2311,In_177,In_945);
and U2312 (N_2312,In_701,In_317);
and U2313 (N_2313,In_551,In_652);
and U2314 (N_2314,In_438,In_109);
or U2315 (N_2315,In_773,In_888);
nor U2316 (N_2316,In_613,In_952);
and U2317 (N_2317,In_628,In_570);
nor U2318 (N_2318,In_758,In_26);
nand U2319 (N_2319,In_669,In_958);
nor U2320 (N_2320,In_113,In_478);
nor U2321 (N_2321,In_830,In_943);
or U2322 (N_2322,In_887,In_84);
nand U2323 (N_2323,In_559,In_1);
and U2324 (N_2324,In_277,In_39);
or U2325 (N_2325,In_233,In_79);
and U2326 (N_2326,In_704,In_140);
and U2327 (N_2327,In_626,In_518);
and U2328 (N_2328,In_368,In_574);
nor U2329 (N_2329,In_748,In_936);
and U2330 (N_2330,In_224,In_227);
nor U2331 (N_2331,In_952,In_468);
and U2332 (N_2332,In_291,In_435);
nand U2333 (N_2333,In_986,In_397);
nand U2334 (N_2334,In_273,In_820);
nor U2335 (N_2335,In_303,In_620);
nand U2336 (N_2336,In_197,In_490);
xor U2337 (N_2337,In_140,In_79);
and U2338 (N_2338,In_186,In_45);
nor U2339 (N_2339,In_107,In_246);
nor U2340 (N_2340,In_967,In_186);
or U2341 (N_2341,In_0,In_121);
nand U2342 (N_2342,In_5,In_64);
or U2343 (N_2343,In_762,In_439);
and U2344 (N_2344,In_927,In_932);
and U2345 (N_2345,In_209,In_412);
nand U2346 (N_2346,In_352,In_898);
nor U2347 (N_2347,In_639,In_494);
nor U2348 (N_2348,In_965,In_237);
and U2349 (N_2349,In_743,In_948);
nor U2350 (N_2350,In_16,In_87);
nor U2351 (N_2351,In_489,In_861);
and U2352 (N_2352,In_933,In_271);
nand U2353 (N_2353,In_975,In_325);
nand U2354 (N_2354,In_72,In_625);
nand U2355 (N_2355,In_784,In_637);
nor U2356 (N_2356,In_955,In_854);
and U2357 (N_2357,In_122,In_331);
or U2358 (N_2358,In_317,In_940);
nor U2359 (N_2359,In_824,In_319);
and U2360 (N_2360,In_302,In_793);
or U2361 (N_2361,In_449,In_491);
nor U2362 (N_2362,In_388,In_528);
and U2363 (N_2363,In_284,In_643);
nor U2364 (N_2364,In_375,In_831);
or U2365 (N_2365,In_274,In_698);
nand U2366 (N_2366,In_162,In_70);
nor U2367 (N_2367,In_643,In_437);
nand U2368 (N_2368,In_41,In_735);
nand U2369 (N_2369,In_502,In_961);
nor U2370 (N_2370,In_598,In_314);
nand U2371 (N_2371,In_908,In_203);
nor U2372 (N_2372,In_340,In_141);
and U2373 (N_2373,In_611,In_84);
and U2374 (N_2374,In_464,In_962);
and U2375 (N_2375,In_268,In_518);
or U2376 (N_2376,In_871,In_579);
nand U2377 (N_2377,In_234,In_578);
nor U2378 (N_2378,In_958,In_194);
nand U2379 (N_2379,In_685,In_368);
nor U2380 (N_2380,In_901,In_846);
nor U2381 (N_2381,In_515,In_365);
or U2382 (N_2382,In_489,In_391);
or U2383 (N_2383,In_918,In_472);
and U2384 (N_2384,In_219,In_73);
nor U2385 (N_2385,In_30,In_604);
or U2386 (N_2386,In_468,In_515);
nor U2387 (N_2387,In_765,In_467);
or U2388 (N_2388,In_963,In_648);
nand U2389 (N_2389,In_815,In_487);
and U2390 (N_2390,In_242,In_42);
or U2391 (N_2391,In_256,In_541);
or U2392 (N_2392,In_816,In_90);
or U2393 (N_2393,In_518,In_26);
and U2394 (N_2394,In_942,In_323);
or U2395 (N_2395,In_435,In_705);
and U2396 (N_2396,In_787,In_461);
nor U2397 (N_2397,In_564,In_419);
nand U2398 (N_2398,In_78,In_186);
and U2399 (N_2399,In_234,In_249);
and U2400 (N_2400,In_436,In_247);
nand U2401 (N_2401,In_744,In_369);
nand U2402 (N_2402,In_921,In_250);
nand U2403 (N_2403,In_17,In_551);
and U2404 (N_2404,In_699,In_694);
or U2405 (N_2405,In_141,In_724);
nand U2406 (N_2406,In_143,In_729);
nor U2407 (N_2407,In_959,In_182);
or U2408 (N_2408,In_429,In_683);
nand U2409 (N_2409,In_154,In_846);
nand U2410 (N_2410,In_478,In_301);
nand U2411 (N_2411,In_726,In_137);
and U2412 (N_2412,In_40,In_893);
or U2413 (N_2413,In_117,In_782);
nand U2414 (N_2414,In_434,In_152);
nand U2415 (N_2415,In_506,In_932);
nor U2416 (N_2416,In_870,In_561);
or U2417 (N_2417,In_782,In_928);
nor U2418 (N_2418,In_344,In_642);
nand U2419 (N_2419,In_481,In_685);
nor U2420 (N_2420,In_300,In_462);
or U2421 (N_2421,In_938,In_830);
nand U2422 (N_2422,In_718,In_539);
or U2423 (N_2423,In_284,In_406);
or U2424 (N_2424,In_136,In_287);
nand U2425 (N_2425,In_834,In_209);
nor U2426 (N_2426,In_414,In_211);
and U2427 (N_2427,In_878,In_234);
or U2428 (N_2428,In_492,In_171);
or U2429 (N_2429,In_40,In_234);
nand U2430 (N_2430,In_821,In_50);
nand U2431 (N_2431,In_448,In_356);
and U2432 (N_2432,In_834,In_474);
or U2433 (N_2433,In_675,In_986);
nand U2434 (N_2434,In_553,In_961);
nor U2435 (N_2435,In_811,In_427);
or U2436 (N_2436,In_266,In_564);
or U2437 (N_2437,In_749,In_109);
or U2438 (N_2438,In_8,In_951);
nand U2439 (N_2439,In_781,In_638);
nor U2440 (N_2440,In_543,In_662);
nor U2441 (N_2441,In_456,In_801);
or U2442 (N_2442,In_371,In_154);
nor U2443 (N_2443,In_981,In_677);
nor U2444 (N_2444,In_685,In_587);
nand U2445 (N_2445,In_975,In_424);
and U2446 (N_2446,In_105,In_378);
and U2447 (N_2447,In_186,In_682);
nand U2448 (N_2448,In_349,In_141);
or U2449 (N_2449,In_147,In_648);
or U2450 (N_2450,In_100,In_954);
and U2451 (N_2451,In_319,In_553);
nand U2452 (N_2452,In_474,In_905);
and U2453 (N_2453,In_302,In_67);
nor U2454 (N_2454,In_88,In_748);
nand U2455 (N_2455,In_970,In_918);
and U2456 (N_2456,In_312,In_309);
or U2457 (N_2457,In_549,In_57);
nand U2458 (N_2458,In_387,In_872);
or U2459 (N_2459,In_378,In_682);
nor U2460 (N_2460,In_122,In_589);
nor U2461 (N_2461,In_770,In_374);
nor U2462 (N_2462,In_855,In_504);
or U2463 (N_2463,In_792,In_377);
nand U2464 (N_2464,In_461,In_370);
nand U2465 (N_2465,In_466,In_692);
and U2466 (N_2466,In_859,In_75);
or U2467 (N_2467,In_531,In_789);
nor U2468 (N_2468,In_33,In_575);
and U2469 (N_2469,In_467,In_731);
or U2470 (N_2470,In_92,In_662);
nor U2471 (N_2471,In_929,In_206);
nor U2472 (N_2472,In_781,In_321);
or U2473 (N_2473,In_884,In_985);
nand U2474 (N_2474,In_110,In_106);
or U2475 (N_2475,In_346,In_424);
nor U2476 (N_2476,In_620,In_403);
nand U2477 (N_2477,In_974,In_468);
and U2478 (N_2478,In_282,In_766);
nand U2479 (N_2479,In_153,In_276);
nor U2480 (N_2480,In_868,In_197);
or U2481 (N_2481,In_333,In_419);
nand U2482 (N_2482,In_2,In_863);
or U2483 (N_2483,In_972,In_480);
or U2484 (N_2484,In_698,In_867);
nand U2485 (N_2485,In_290,In_912);
and U2486 (N_2486,In_880,In_258);
or U2487 (N_2487,In_435,In_174);
nand U2488 (N_2488,In_658,In_761);
nor U2489 (N_2489,In_432,In_744);
nand U2490 (N_2490,In_793,In_919);
or U2491 (N_2491,In_337,In_79);
and U2492 (N_2492,In_960,In_418);
nor U2493 (N_2493,In_230,In_167);
nand U2494 (N_2494,In_239,In_746);
nand U2495 (N_2495,In_757,In_646);
nand U2496 (N_2496,In_6,In_837);
and U2497 (N_2497,In_857,In_985);
nand U2498 (N_2498,In_206,In_210);
or U2499 (N_2499,In_546,In_447);
nor U2500 (N_2500,N_744,N_1481);
and U2501 (N_2501,N_706,N_936);
and U2502 (N_2502,N_630,N_32);
and U2503 (N_2503,N_599,N_2472);
nor U2504 (N_2504,N_1501,N_608);
and U2505 (N_2505,N_180,N_1827);
nor U2506 (N_2506,N_492,N_1524);
or U2507 (N_2507,N_831,N_1960);
and U2508 (N_2508,N_1895,N_1076);
nor U2509 (N_2509,N_2491,N_1318);
nor U2510 (N_2510,N_484,N_2165);
or U2511 (N_2511,N_1543,N_591);
nor U2512 (N_2512,N_600,N_1366);
or U2513 (N_2513,N_355,N_1836);
nor U2514 (N_2514,N_987,N_1450);
nor U2515 (N_2515,N_682,N_2328);
nor U2516 (N_2516,N_895,N_19);
nand U2517 (N_2517,N_1986,N_2419);
nand U2518 (N_2518,N_1376,N_1518);
or U2519 (N_2519,N_2348,N_293);
nor U2520 (N_2520,N_2015,N_1843);
or U2521 (N_2521,N_1673,N_2313);
and U2522 (N_2522,N_269,N_1298);
nand U2523 (N_2523,N_977,N_2321);
or U2524 (N_2524,N_704,N_899);
or U2525 (N_2525,N_1891,N_1958);
nor U2526 (N_2526,N_2042,N_673);
nand U2527 (N_2527,N_954,N_2143);
and U2528 (N_2528,N_1175,N_1597);
and U2529 (N_2529,N_65,N_637);
and U2530 (N_2530,N_2260,N_2254);
nor U2531 (N_2531,N_2232,N_585);
nor U2532 (N_2532,N_1754,N_1005);
and U2533 (N_2533,N_399,N_73);
nor U2534 (N_2534,N_1092,N_1688);
or U2535 (N_2535,N_175,N_1896);
nor U2536 (N_2536,N_295,N_2392);
and U2537 (N_2537,N_549,N_2197);
and U2538 (N_2538,N_1401,N_938);
or U2539 (N_2539,N_2410,N_2019);
nand U2540 (N_2540,N_2294,N_788);
nor U2541 (N_2541,N_2344,N_2102);
nand U2542 (N_2542,N_1874,N_1581);
and U2543 (N_2543,N_315,N_618);
or U2544 (N_2544,N_441,N_2479);
or U2545 (N_2545,N_2371,N_1806);
or U2546 (N_2546,N_1341,N_2293);
or U2547 (N_2547,N_955,N_243);
nor U2548 (N_2548,N_2481,N_2338);
nand U2549 (N_2549,N_826,N_834);
nand U2550 (N_2550,N_991,N_1040);
nor U2551 (N_2551,N_1147,N_1582);
or U2552 (N_2552,N_2257,N_613);
nor U2553 (N_2553,N_932,N_359);
or U2554 (N_2554,N_1232,N_2107);
nor U2555 (N_2555,N_402,N_222);
nor U2556 (N_2556,N_1657,N_1238);
nand U2557 (N_2557,N_1864,N_1662);
or U2558 (N_2558,N_1235,N_1844);
and U2559 (N_2559,N_2450,N_229);
nor U2560 (N_2560,N_1505,N_2098);
and U2561 (N_2561,N_661,N_153);
or U2562 (N_2562,N_2246,N_2306);
nor U2563 (N_2563,N_660,N_1104);
nor U2564 (N_2564,N_483,N_1113);
nor U2565 (N_2565,N_2224,N_1568);
nor U2566 (N_2566,N_343,N_964);
nand U2567 (N_2567,N_2092,N_2394);
and U2568 (N_2568,N_1344,N_2498);
nand U2569 (N_2569,N_2148,N_1796);
nand U2570 (N_2570,N_780,N_2453);
nor U2571 (N_2571,N_1359,N_1017);
and U2572 (N_2572,N_835,N_183);
or U2573 (N_2573,N_78,N_240);
and U2574 (N_2574,N_2298,N_1773);
nand U2575 (N_2575,N_1456,N_2071);
and U2576 (N_2576,N_635,N_1669);
or U2577 (N_2577,N_284,N_373);
nand U2578 (N_2578,N_2324,N_1852);
or U2579 (N_2579,N_1496,N_793);
nand U2580 (N_2580,N_1752,N_2047);
nor U2581 (N_2581,N_1508,N_2168);
nand U2582 (N_2582,N_1762,N_832);
and U2583 (N_2583,N_409,N_2242);
nand U2584 (N_2584,N_442,N_513);
or U2585 (N_2585,N_809,N_461);
or U2586 (N_2586,N_1382,N_843);
or U2587 (N_2587,N_1025,N_700);
and U2588 (N_2588,N_514,N_1275);
nand U2589 (N_2589,N_2393,N_733);
and U2590 (N_2590,N_2438,N_499);
and U2591 (N_2591,N_1075,N_1815);
or U2592 (N_2592,N_361,N_686);
nor U2593 (N_2593,N_49,N_1732);
nand U2594 (N_2594,N_703,N_322);
nand U2595 (N_2595,N_2170,N_259);
and U2596 (N_2596,N_1443,N_1941);
and U2597 (N_2597,N_1194,N_1234);
nand U2598 (N_2598,N_1853,N_176);
and U2599 (N_2599,N_2327,N_2243);
or U2600 (N_2600,N_420,N_1408);
nor U2601 (N_2601,N_1247,N_1107);
and U2602 (N_2602,N_2449,N_206);
nor U2603 (N_2603,N_2196,N_1438);
and U2604 (N_2604,N_453,N_1008);
and U2605 (N_2605,N_1070,N_2354);
nand U2606 (N_2606,N_1161,N_2191);
and U2607 (N_2607,N_1979,N_1294);
nor U2608 (N_2608,N_2401,N_965);
or U2609 (N_2609,N_401,N_2139);
nand U2610 (N_2610,N_1830,N_1621);
or U2611 (N_2611,N_2404,N_1368);
nand U2612 (N_2612,N_160,N_2346);
or U2613 (N_2613,N_1934,N_1845);
nand U2614 (N_2614,N_1073,N_1525);
nand U2615 (N_2615,N_1930,N_1677);
or U2616 (N_2616,N_852,N_2110);
nand U2617 (N_2617,N_552,N_1411);
or U2618 (N_2618,N_2012,N_893);
nand U2619 (N_2619,N_2146,N_1586);
nand U2620 (N_2620,N_2446,N_111);
or U2621 (N_2621,N_2462,N_15);
nor U2622 (N_2622,N_1851,N_156);
or U2623 (N_2623,N_1856,N_533);
nor U2624 (N_2624,N_953,N_1010);
or U2625 (N_2625,N_507,N_1530);
nor U2626 (N_2626,N_2417,N_1559);
nand U2627 (N_2627,N_1015,N_550);
nand U2628 (N_2628,N_2087,N_1417);
nor U2629 (N_2629,N_999,N_597);
and U2630 (N_2630,N_594,N_314);
and U2631 (N_2631,N_134,N_1223);
nand U2632 (N_2632,N_1094,N_2266);
or U2633 (N_2633,N_625,N_676);
nor U2634 (N_2634,N_864,N_1336);
nand U2635 (N_2635,N_2433,N_1221);
nor U2636 (N_2636,N_1445,N_1317);
or U2637 (N_2637,N_2355,N_350);
nand U2638 (N_2638,N_927,N_2290);
or U2639 (N_2639,N_1935,N_2383);
nand U2640 (N_2640,N_2362,N_288);
nand U2641 (N_2641,N_447,N_2264);
nand U2642 (N_2642,N_1486,N_726);
nand U2643 (N_2643,N_1548,N_285);
or U2644 (N_2644,N_567,N_2089);
or U2645 (N_2645,N_1579,N_779);
or U2646 (N_2646,N_1848,N_140);
nor U2647 (N_2647,N_1982,N_1605);
or U2648 (N_2648,N_980,N_523);
nand U2649 (N_2649,N_918,N_1499);
nand U2650 (N_2650,N_2311,N_1434);
and U2651 (N_2651,N_1129,N_553);
nor U2652 (N_2652,N_556,N_1765);
nor U2653 (N_2653,N_769,N_1829);
nand U2654 (N_2654,N_2268,N_2238);
or U2655 (N_2655,N_376,N_1573);
nand U2656 (N_2656,N_1013,N_2085);
nand U2657 (N_2657,N_1420,N_2125);
and U2658 (N_2658,N_577,N_1239);
or U2659 (N_2659,N_2063,N_1196);
nand U2660 (N_2660,N_2276,N_202);
nand U2661 (N_2661,N_52,N_1976);
nand U2662 (N_2662,N_425,N_2229);
and U2663 (N_2663,N_1159,N_2323);
nor U2664 (N_2664,N_854,N_79);
nand U2665 (N_2665,N_609,N_1280);
nor U2666 (N_2666,N_1465,N_1000);
nor U2667 (N_2667,N_1973,N_2499);
nand U2668 (N_2668,N_1691,N_2209);
nor U2669 (N_2669,N_1031,N_422);
nand U2670 (N_2670,N_1060,N_2486);
or U2671 (N_2671,N_667,N_1333);
nor U2672 (N_2672,N_1687,N_1213);
and U2673 (N_2673,N_2384,N_1813);
nand U2674 (N_2674,N_1674,N_1590);
nor U2675 (N_2675,N_1780,N_297);
and U2676 (N_2676,N_966,N_997);
or U2677 (N_2677,N_2008,N_1698);
and U2678 (N_2678,N_1176,N_1255);
and U2679 (N_2679,N_712,N_735);
nor U2680 (N_2680,N_164,N_708);
nand U2681 (N_2681,N_1968,N_1470);
or U2682 (N_2682,N_1216,N_396);
or U2683 (N_2683,N_127,N_2342);
or U2684 (N_2684,N_1718,N_2090);
nor U2685 (N_2685,N_2072,N_477);
nor U2686 (N_2686,N_2195,N_626);
nand U2687 (N_2687,N_325,N_1068);
or U2688 (N_2688,N_272,N_1711);
nor U2689 (N_2689,N_2253,N_2334);
nor U2690 (N_2690,N_945,N_2333);
nand U2691 (N_2691,N_346,N_1198);
and U2692 (N_2692,N_471,N_1328);
or U2693 (N_2693,N_18,N_1775);
and U2694 (N_2694,N_981,N_825);
or U2695 (N_2695,N_531,N_2112);
nor U2696 (N_2696,N_1746,N_97);
nand U2697 (N_2697,N_1870,N_1978);
or U2698 (N_2698,N_1915,N_1314);
nor U2699 (N_2699,N_1115,N_118);
nor U2700 (N_2700,N_659,N_1609);
and U2701 (N_2701,N_1670,N_743);
nand U2702 (N_2702,N_1144,N_2002);
or U2703 (N_2703,N_1566,N_1759);
nor U2704 (N_2704,N_1479,N_1360);
nor U2705 (N_2705,N_0,N_569);
nand U2706 (N_2706,N_1347,N_1146);
nor U2707 (N_2707,N_1410,N_12);
nor U2708 (N_2708,N_639,N_2034);
nand U2709 (N_2709,N_1660,N_536);
or U2710 (N_2710,N_1527,N_1028);
and U2711 (N_2711,N_1682,N_1584);
nor U2712 (N_2712,N_1984,N_1576);
nor U2713 (N_2713,N_518,N_2303);
nor U2714 (N_2714,N_790,N_254);
and U2715 (N_2715,N_683,N_227);
xor U2716 (N_2716,N_896,N_1975);
nor U2717 (N_2717,N_1804,N_1021);
and U2718 (N_2718,N_707,N_935);
and U2719 (N_2719,N_1556,N_302);
and U2720 (N_2720,N_2483,N_873);
or U2721 (N_2721,N_730,N_1257);
or U2722 (N_2722,N_200,N_1515);
or U2723 (N_2723,N_2415,N_1211);
and U2724 (N_2724,N_2045,N_1872);
nor U2725 (N_2725,N_1425,N_846);
nand U2726 (N_2726,N_1447,N_2183);
and U2727 (N_2727,N_1051,N_1517);
or U2728 (N_2728,N_1545,N_1835);
xor U2729 (N_2729,N_1335,N_737);
nor U2730 (N_2730,N_96,N_604);
nor U2731 (N_2731,N_1920,N_332);
nand U2732 (N_2732,N_146,N_908);
and U2733 (N_2733,N_891,N_1610);
or U2734 (N_2734,N_474,N_887);
and U2735 (N_2735,N_2007,N_1735);
nor U2736 (N_2736,N_1909,N_1353);
or U2737 (N_2737,N_612,N_239);
and U2738 (N_2738,N_1743,N_281);
nor U2739 (N_2739,N_1726,N_890);
nor U2740 (N_2740,N_1081,N_1418);
nand U2741 (N_2741,N_654,N_656);
or U2742 (N_2742,N_1854,N_674);
and U2743 (N_2743,N_405,N_729);
nor U2744 (N_2744,N_1435,N_798);
and U2745 (N_2745,N_2021,N_414);
nand U2746 (N_2746,N_506,N_219);
and U2747 (N_2747,N_113,N_1277);
nor U2748 (N_2748,N_1840,N_2167);
and U2749 (N_2749,N_1331,N_1055);
and U2750 (N_2750,N_287,N_1308);
nor U2751 (N_2751,N_970,N_2162);
nor U2752 (N_2752,N_1062,N_2339);
nor U2753 (N_2753,N_473,N_1220);
or U2754 (N_2754,N_1903,N_1391);
and U2755 (N_2755,N_329,N_1322);
nand U2756 (N_2756,N_1444,N_1282);
and U2757 (N_2757,N_889,N_27);
nand U2758 (N_2758,N_9,N_1596);
nand U2759 (N_2759,N_1689,N_944);
nor U2760 (N_2760,N_386,N_2035);
nand U2761 (N_2761,N_1003,N_273);
nor U2762 (N_2762,N_1064,N_1024);
or U2763 (N_2763,N_1266,N_2128);
nand U2764 (N_2764,N_2458,N_2077);
and U2765 (N_2765,N_923,N_276);
nor U2766 (N_2766,N_2285,N_1699);
xnor U2767 (N_2767,N_387,N_1777);
nand U2768 (N_2768,N_1925,N_1230);
nor U2769 (N_2769,N_641,N_1821);
nand U2770 (N_2770,N_1324,N_100);
or U2771 (N_2771,N_2274,N_398);
or U2772 (N_2772,N_275,N_1338);
or U2773 (N_2773,N_86,N_1589);
or U2774 (N_2774,N_241,N_1065);
nand U2775 (N_2775,N_2140,N_1702);
and U2776 (N_2776,N_481,N_1912);
nor U2777 (N_2777,N_1138,N_1188);
nand U2778 (N_2778,N_1833,N_898);
and U2779 (N_2779,N_452,N_1936);
or U2780 (N_2780,N_23,N_1858);
nor U2781 (N_2781,N_721,N_1798);
nand U2782 (N_2782,N_872,N_855);
and U2783 (N_2783,N_1602,N_2105);
nand U2784 (N_2784,N_2043,N_1069);
and U2785 (N_2785,N_321,N_1953);
nor U2786 (N_2786,N_371,N_636);
nand U2787 (N_2787,N_2241,N_963);
nand U2788 (N_2788,N_1634,N_2225);
and U2789 (N_2789,N_677,N_1439);
and U2790 (N_2790,N_1174,N_1728);
nor U2791 (N_2791,N_2441,N_267);
nand U2792 (N_2792,N_362,N_1371);
and U2793 (N_2793,N_2489,N_464);
and U2794 (N_2794,N_1259,N_413);
nand U2795 (N_2795,N_764,N_38);
nand U2796 (N_2796,N_1863,N_39);
nor U2797 (N_2797,N_958,N_1473);
nand U2798 (N_2798,N_2316,N_713);
or U2799 (N_2799,N_985,N_21);
or U2800 (N_2800,N_2261,N_1822);
nor U2801 (N_2801,N_1016,N_763);
nand U2802 (N_2802,N_313,N_1367);
and U2803 (N_2803,N_1949,N_861);
nor U2804 (N_2804,N_973,N_1717);
and U2805 (N_2805,N_2397,N_2070);
and U2806 (N_2806,N_2374,N_2149);
nand U2807 (N_2807,N_959,N_1957);
nand U2808 (N_2808,N_1433,N_1767);
or U2809 (N_2809,N_1977,N_2385);
nand U2810 (N_2810,N_1913,N_1938);
nand U2811 (N_2811,N_1562,N_906);
and U2812 (N_2812,N_1170,N_388);
nor U2813 (N_2813,N_1440,N_1380);
and U2814 (N_2814,N_66,N_2388);
and U2815 (N_2815,N_142,N_178);
nor U2816 (N_2816,N_1379,N_505);
and U2817 (N_2817,N_2343,N_653);
nor U2818 (N_2818,N_2381,N_1084);
nor U2819 (N_2819,N_2061,N_722);
or U2820 (N_2820,N_586,N_853);
or U2821 (N_2821,N_2469,N_2065);
nor U2822 (N_2822,N_1637,N_1036);
or U2823 (N_2823,N_574,N_2424);
nor U2824 (N_2824,N_463,N_1477);
nor U2825 (N_2825,N_1183,N_2192);
and U2826 (N_2826,N_1210,N_2447);
nor U2827 (N_2827,N_642,N_2492);
nand U2828 (N_2828,N_1659,N_572);
or U2829 (N_2829,N_949,N_1607);
or U2830 (N_2830,N_128,N_266);
or U2831 (N_2831,N_2208,N_379);
nor U2832 (N_2832,N_2411,N_1177);
nor U2833 (N_2833,N_177,N_1424);
nand U2834 (N_2834,N_1831,N_231);
nor U2835 (N_2835,N_2138,N_516);
or U2836 (N_2836,N_1727,N_415);
or U2837 (N_2837,N_1719,N_1880);
nand U2838 (N_2838,N_2091,N_2423);
and U2839 (N_2839,N_40,N_2006);
and U2840 (N_2840,N_1661,N_1948);
and U2841 (N_2841,N_1878,N_1514);
nor U2842 (N_2842,N_228,N_1561);
nor U2843 (N_2843,N_1990,N_205);
and U2844 (N_2844,N_1722,N_521);
and U2845 (N_2845,N_669,N_294);
nand U2846 (N_2846,N_2050,N_1544);
nand U2847 (N_2847,N_1100,N_1180);
or U2848 (N_2848,N_139,N_539);
and U2849 (N_2849,N_1665,N_2456);
and U2850 (N_2850,N_360,N_1120);
nand U2851 (N_2851,N_1816,N_2004);
or U2852 (N_2852,N_1416,N_2184);
or U2853 (N_2853,N_147,N_1828);
or U2854 (N_2854,N_1027,N_1488);
nor U2855 (N_2855,N_1291,N_2101);
or U2856 (N_2856,N_1205,N_2312);
nand U2857 (N_2857,N_1599,N_2391);
or U2858 (N_2858,N_3,N_2439);
nand U2859 (N_2859,N_2283,N_2096);
and U2860 (N_2860,N_1970,N_995);
nor U2861 (N_2861,N_1469,N_1739);
and U2862 (N_2862,N_848,N_1315);
nor U2863 (N_2863,N_2451,N_1857);
xor U2864 (N_2864,N_1906,N_76);
nand U2865 (N_2865,N_335,N_2194);
nor U2866 (N_2866,N_496,N_1537);
nand U2867 (N_2867,N_6,N_2088);
and U2868 (N_2868,N_270,N_559);
or U2869 (N_2869,N_644,N_529);
and U2870 (N_2870,N_1114,N_1683);
nor U2871 (N_2871,N_232,N_2273);
xnor U2872 (N_2872,N_1241,N_1252);
and U2873 (N_2873,N_880,N_876);
nor U2874 (N_2874,N_1904,N_976);
and U2875 (N_2875,N_69,N_1348);
and U2876 (N_2876,N_462,N_479);
nand U2877 (N_2877,N_458,N_1074);
and U2878 (N_2878,N_211,N_470);
nand U2879 (N_2879,N_851,N_1243);
nand U2880 (N_2880,N_2382,N_61);
nor U2881 (N_2881,N_1914,N_26);
nand U2882 (N_2882,N_1458,N_1928);
or U2883 (N_2883,N_582,N_1924);
nand U2884 (N_2884,N_2444,N_1145);
nand U2885 (N_2885,N_2173,N_102);
nand U2886 (N_2886,N_487,N_1538);
and U2887 (N_2887,N_2267,N_1459);
or U2888 (N_2888,N_690,N_878);
nand U2889 (N_2889,N_323,N_571);
xor U2890 (N_2890,N_2048,N_2027);
and U2891 (N_2891,N_2062,N_2074);
and U2892 (N_2892,N_55,N_799);
nand U2893 (N_2893,N_565,N_2305);
nor U2894 (N_2894,N_2188,N_2059);
nor U2895 (N_2895,N_347,N_260);
and U2896 (N_2896,N_1088,N_969);
and U2897 (N_2897,N_397,N_226);
and U2898 (N_2898,N_1231,N_519);
or U2899 (N_2899,N_1419,N_1510);
nor U2900 (N_2900,N_1867,N_1721);
nor U2901 (N_2901,N_620,N_647);
nand U2902 (N_2902,N_2127,N_187);
or U2903 (N_2903,N_1681,N_165);
nand U2904 (N_2904,N_2473,N_1403);
or U2905 (N_2905,N_687,N_377);
nand U2906 (N_2906,N_2161,N_2198);
and U2907 (N_2907,N_1849,N_740);
xnor U2908 (N_2908,N_290,N_913);
nor U2909 (N_2909,N_1006,N_1395);
nand U2910 (N_2910,N_1884,N_1736);
nor U2911 (N_2911,N_759,N_874);
nor U2912 (N_2912,N_385,N_1492);
nor U2913 (N_2913,N_237,N_334);
nand U2914 (N_2914,N_509,N_617);
or U2915 (N_2915,N_1785,N_1786);
and U2916 (N_2916,N_917,N_2420);
and U2917 (N_2917,N_451,N_1431);
and U2918 (N_2918,N_418,N_190);
nor U2919 (N_2919,N_1731,N_31);
and U2920 (N_2920,N_924,N_1133);
or U2921 (N_2921,N_548,N_540);
or U2922 (N_2922,N_527,N_1185);
and U2923 (N_2923,N_2475,N_104);
nand U2924 (N_2924,N_1894,N_291);
and U2925 (N_2925,N_1554,N_1327);
or U2926 (N_2926,N_1952,N_1105);
nor U2927 (N_2927,N_108,N_2428);
and U2928 (N_2928,N_1511,N_1811);
or U2929 (N_2929,N_2322,N_1781);
and U2930 (N_2930,N_1415,N_392);
or U2931 (N_2931,N_1766,N_668);
nand U2932 (N_2932,N_2020,N_207);
xor U2933 (N_2933,N_1041,N_2069);
nor U2934 (N_2934,N_2277,N_1955);
nor U2935 (N_2935,N_1276,N_221);
and U2936 (N_2936,N_184,N_1883);
or U2937 (N_2937,N_1404,N_590);
nand U2938 (N_2938,N_1377,N_1149);
or U2939 (N_2939,N_2250,N_498);
nand U2940 (N_2940,N_497,N_106);
nand U2941 (N_2941,N_828,N_2289);
nand U2942 (N_2942,N_311,N_246);
nor U2943 (N_2943,N_892,N_638);
nor U2944 (N_2944,N_1564,N_1755);
and U2945 (N_2945,N_67,N_2078);
or U2946 (N_2946,N_2024,N_2304);
and U2947 (N_2947,N_2117,N_670);
nand U2948 (N_2948,N_2465,N_979);
or U2949 (N_2949,N_2398,N_1892);
nand U2950 (N_2950,N_2129,N_1209);
or U2951 (N_2951,N_542,N_17);
nand U2952 (N_2952,N_717,N_665);
and U2953 (N_2953,N_82,N_1504);
and U2954 (N_2954,N_367,N_1897);
nand U2955 (N_2955,N_640,N_1300);
nor U2956 (N_2956,N_1242,N_450);
or U2957 (N_2957,N_437,N_2054);
nor U2958 (N_2958,N_1623,N_1922);
and U2959 (N_2959,N_2206,N_99);
and U2960 (N_2960,N_2,N_1558);
or U2961 (N_2961,N_2134,N_2278);
and U2962 (N_2962,N_1110,N_1640);
nand U2963 (N_2963,N_528,N_598);
nor U2964 (N_2964,N_837,N_1182);
or U2965 (N_2965,N_947,N_2459);
nor U2966 (N_2966,N_172,N_169);
and U2967 (N_2967,N_1267,N_1725);
or U2968 (N_2968,N_1449,N_824);
nor U2969 (N_2969,N_1436,N_1741);
or U2970 (N_2970,N_1394,N_1509);
nand U2971 (N_2971,N_1224,N_1421);
or U2972 (N_2972,N_2335,N_2309);
and U2973 (N_2973,N_1671,N_10);
nor U2974 (N_2974,N_1099,N_72);
nor U2975 (N_2975,N_576,N_986);
nor U2976 (N_2976,N_1685,N_1124);
nor U2977 (N_2977,N_1162,N_1289);
or U2978 (N_2978,N_1042,N_1624);
nand U2979 (N_2979,N_1153,N_2288);
and U2980 (N_2980,N_2297,N_1818);
nand U2981 (N_2981,N_1292,N_561);
nor U2982 (N_2982,N_1690,N_1279);
nand U2983 (N_2983,N_2467,N_300);
and U2984 (N_2984,N_1026,N_131);
nand U2985 (N_2985,N_1046,N_1414);
nand U2986 (N_2986,N_107,N_2057);
or U2987 (N_2987,N_1052,N_1567);
or U2988 (N_2988,N_1842,N_7);
and U2989 (N_2989,N_2314,N_1030);
nor U2990 (N_2990,N_1893,N_150);
nand U2991 (N_2991,N_356,N_2113);
nand U2992 (N_2992,N_1283,N_2186);
nor U2993 (N_2993,N_2023,N_1575);
nand U2994 (N_2994,N_1810,N_204);
nor U2995 (N_2995,N_797,N_711);
xnor U2996 (N_2996,N_2119,N_1776);
and U2997 (N_2997,N_265,N_1071);
nand U2998 (N_2998,N_491,N_2056);
nand U2999 (N_2999,N_59,N_1812);
nand U3000 (N_3000,N_2443,N_2395);
nor U3001 (N_3001,N_51,N_1078);
and U3002 (N_3002,N_731,N_2426);
or U3003 (N_3003,N_1150,N_784);
nor U3004 (N_3004,N_1983,N_1119);
or U3005 (N_3005,N_1190,N_132);
or U3006 (N_3006,N_666,N_2211);
nand U3007 (N_3007,N_766,N_709);
nand U3008 (N_3008,N_1422,N_882);
and U3009 (N_3009,N_1601,N_2222);
or U3010 (N_3010,N_1466,N_1233);
or U3011 (N_3011,N_1516,N_616);
nand U3012 (N_3012,N_1201,N_217);
nand U3013 (N_3013,N_57,N_960);
nand U3014 (N_3014,N_2099,N_905);
or U3015 (N_3015,N_1463,N_2227);
nand U3016 (N_3016,N_24,N_1364);
nor U3017 (N_3017,N_366,N_2234);
or U3018 (N_3018,N_1532,N_2178);
nand U3019 (N_3019,N_1061,N_1716);
nand U3020 (N_3020,N_304,N_1167);
or U3021 (N_3021,N_1014,N_930);
nor U3022 (N_3022,N_2142,N_25);
nand U3023 (N_3023,N_500,N_1142);
nor U3024 (N_3024,N_1089,N_672);
nor U3025 (N_3025,N_624,N_504);
nand U3026 (N_3026,N_1917,N_1506);
or U3027 (N_3027,N_1552,N_428);
nor U3028 (N_3028,N_1963,N_1820);
nand U3029 (N_3029,N_723,N_2082);
or U3030 (N_3030,N_490,N_167);
or U3031 (N_3031,N_233,N_1409);
and U3032 (N_3032,N_2060,N_120);
nand U3033 (N_3033,N_305,N_1093);
and U3034 (N_3034,N_1549,N_1423);
and U3035 (N_3035,N_727,N_956);
and U3036 (N_3036,N_1495,N_847);
nor U3037 (N_3037,N_1097,N_279);
nor U3038 (N_3038,N_2478,N_166);
or U3039 (N_3039,N_2247,N_517);
and U3040 (N_3040,N_2413,N_2133);
nand U3041 (N_3041,N_2380,N_2172);
nor U3042 (N_3042,N_1109,N_1012);
nand U3043 (N_3043,N_1163,N_812);
nand U3044 (N_3044,N_2095,N_2097);
nand U3045 (N_3045,N_454,N_137);
and U3046 (N_3046,N_901,N_789);
or U3047 (N_3047,N_35,N_773);
nor U3048 (N_3048,N_130,N_1859);
or U3049 (N_3049,N_1826,N_1877);
and U3050 (N_3050,N_1989,N_278);
nand U3051 (N_3051,N_1919,N_1855);
nor U3052 (N_3052,N_555,N_2270);
nor U3053 (N_3053,N_2080,N_982);
and U3054 (N_3054,N_1019,N_940);
and U3055 (N_3055,N_1079,N_884);
or U3056 (N_3056,N_1969,N_494);
nand U3057 (N_3057,N_145,N_1058);
or U3058 (N_3058,N_2185,N_319);
or U3059 (N_3059,N_881,N_754);
and U3060 (N_3060,N_2470,N_1219);
nand U3061 (N_3061,N_1988,N_1285);
or U3062 (N_3062,N_1926,N_978);
nand U3063 (N_3063,N_679,N_1521);
nor U3064 (N_3064,N_1313,N_1888);
and U3065 (N_3065,N_1155,N_1937);
nor U3066 (N_3066,N_1037,N_1825);
and U3067 (N_3067,N_1879,N_1303);
nand U3068 (N_3068,N_1135,N_1199);
or U3069 (N_3069,N_501,N_1032);
nor U3070 (N_3070,N_1157,N_251);
or U3071 (N_3071,N_2040,N_596);
nor U3072 (N_3072,N_1222,N_342);
nor U3073 (N_3073,N_250,N_1441);
or U3074 (N_3074,N_1761,N_2269);
and U3075 (N_3075,N_602,N_1009);
nor U3076 (N_3076,N_2436,N_1372);
nor U3077 (N_3077,N_2352,N_475);
nand U3078 (N_3078,N_1090,N_946);
nor U3079 (N_3079,N_1744,N_2177);
nor U3080 (N_3080,N_2408,N_1817);
or U3081 (N_3081,N_1381,N_1966);
nand U3082 (N_3082,N_2480,N_286);
nand U3083 (N_3083,N_2068,N_1954);
nand U3084 (N_3084,N_2412,N_2474);
nand U3085 (N_3085,N_951,N_83);
nand U3086 (N_3086,N_306,N_1992);
nand U3087 (N_3087,N_109,N_2152);
nor U3088 (N_3088,N_1742,N_1302);
nand U3089 (N_3089,N_1656,N_2076);
nand U3090 (N_3090,N_1866,N_416);
and U3091 (N_3091,N_431,N_971);
or U3092 (N_3092,N_1373,N_94);
or U3093 (N_3093,N_421,N_114);
and U3094 (N_3094,N_1063,N_696);
nor U3095 (N_3095,N_651,N_1972);
nand U3096 (N_3096,N_752,N_532);
and U3097 (N_3097,N_2175,N_445);
nand U3098 (N_3098,N_1868,N_728);
or U3099 (N_3099,N_58,N_1165);
nand U3100 (N_3100,N_2226,N_1140);
nor U3101 (N_3101,N_2329,N_564);
and U3102 (N_3102,N_1043,N_2440);
or U3103 (N_3103,N_1965,N_2476);
nor U3104 (N_3104,N_2256,N_2240);
or U3105 (N_3105,N_1272,N_1595);
and U3106 (N_3106,N_64,N_406);
and U3107 (N_3107,N_2151,N_374);
nand U3108 (N_3108,N_400,N_144);
or U3109 (N_3109,N_1655,N_2135);
nand U3110 (N_3110,N_2364,N_262);
or U3111 (N_3111,N_296,N_2400);
nand U3112 (N_3112,N_510,N_8);
nand U3113 (N_3113,N_870,N_389);
or U3114 (N_3114,N_50,N_466);
nand U3115 (N_3115,N_1999,N_345);
xnor U3116 (N_3116,N_327,N_2490);
nor U3117 (N_3117,N_393,N_22);
and U3118 (N_3118,N_1723,N_544);
and U3119 (N_3119,N_1981,N_1551);
or U3120 (N_3120,N_2330,N_1002);
and U3121 (N_3121,N_1933,N_1116);
xor U3122 (N_3122,N_1405,N_842);
nor U3123 (N_3123,N_2028,N_280);
nand U3124 (N_3124,N_1204,N_283);
and U3125 (N_3125,N_903,N_2421);
nand U3126 (N_3126,N_560,N_2493);
and U3127 (N_3127,N_257,N_629);
nand U3128 (N_3128,N_1795,N_1323);
nand U3129 (N_3129,N_996,N_1782);
nor U3130 (N_3130,N_1748,N_5);
and U3131 (N_3131,N_1998,N_354);
and U3132 (N_3132,N_28,N_1374);
nor U3133 (N_3133,N_1784,N_2109);
nor U3134 (N_3134,N_154,N_745);
nor U3135 (N_3135,N_2210,N_472);
or U3136 (N_3136,N_2442,N_363);
or U3137 (N_3137,N_214,N_380);
and U3138 (N_3138,N_1350,N_328);
or U3139 (N_3139,N_1225,N_1365);
nand U3140 (N_3140,N_1383,N_1393);
nor U3141 (N_3141,N_526,N_192);
or U3142 (N_3142,N_2118,N_435);
and U3143 (N_3143,N_316,N_1342);
nor U3144 (N_3144,N_897,N_2286);
and U3145 (N_3145,N_2214,N_1178);
nand U3146 (N_3146,N_1160,N_1797);
xor U3147 (N_3147,N_1668,N_950);
nand U3148 (N_3148,N_829,N_838);
nand U3149 (N_3149,N_1361,N_1236);
nand U3150 (N_3150,N_860,N_1207);
and U3151 (N_3151,N_2052,N_365);
nand U3152 (N_3152,N_720,N_1098);
nor U3153 (N_3153,N_827,N_1898);
nor U3154 (N_3154,N_2407,N_46);
nor U3155 (N_3155,N_2181,N_216);
nor U3156 (N_3156,N_1571,N_242);
and U3157 (N_3157,N_1158,N_1494);
nand U3158 (N_3158,N_607,N_1771);
and U3159 (N_3159,N_1663,N_1942);
or U3160 (N_3160,N_1264,N_2216);
and U3161 (N_3161,N_2049,N_983);
nand U3162 (N_3162,N_1646,N_1077);
nor U3163 (N_3163,N_649,N_1121);
nor U3164 (N_3164,N_919,N_143);
nor U3165 (N_3165,N_783,N_1334);
or U3166 (N_3166,N_1993,N_423);
and U3167 (N_3167,N_2132,N_2379);
xor U3168 (N_3168,N_318,N_1697);
and U3169 (N_3169,N_48,N_777);
nand U3170 (N_3170,N_2308,N_1059);
and U3171 (N_3171,N_98,N_1018);
nor U3172 (N_3172,N_136,N_440);
and U3173 (N_3173,N_480,N_126);
nor U3174 (N_3174,N_2204,N_1929);
or U3175 (N_3175,N_62,N_2340);
and U3176 (N_3176,N_2307,N_593);
and U3177 (N_3177,N_1442,N_253);
nor U3178 (N_3178,N_2466,N_1526);
and U3179 (N_3179,N_815,N_2010);
and U3180 (N_3180,N_681,N_554);
nand U3181 (N_3181,N_1750,N_1096);
nand U3182 (N_3182,N_2389,N_42);
nand U3183 (N_3183,N_2066,N_1995);
nor U3184 (N_3184,N_395,N_408);
or U3185 (N_3185,N_914,N_331);
or U3186 (N_3186,N_1067,N_716);
and U3187 (N_3187,N_1500,N_2484);
nand U3188 (N_3188,N_1512,N_2252);
or U3189 (N_3189,N_1263,N_904);
or U3190 (N_3190,N_515,N_2084);
nor U3191 (N_3191,N_1057,N_975);
nand U3192 (N_3192,N_1004,N_822);
and U3193 (N_3193,N_1799,N_2000);
and U3194 (N_3194,N_210,N_839);
or U3195 (N_3195,N_757,N_1284);
and U3196 (N_3196,N_2136,N_1462);
nor U3197 (N_3197,N_942,N_2349);
nor U3198 (N_3198,N_2284,N_1507);
nor U3199 (N_3199,N_1764,N_1370);
nor U3200 (N_3200,N_2201,N_129);
nor U3201 (N_3201,N_357,N_580);
or U3202 (N_3202,N_1033,N_2347);
nand U3203 (N_3203,N_1102,N_2231);
and U3204 (N_3204,N_1519,N_758);
and U3205 (N_3205,N_1029,N_1357);
and U3206 (N_3206,N_802,N_2016);
and U3207 (N_3207,N_1541,N_2263);
and U3208 (N_3208,N_1356,N_121);
and U3209 (N_3209,N_112,N_1397);
nand U3210 (N_3210,N_63,N_1457);
and U3211 (N_3211,N_1358,N_71);
and U3212 (N_3212,N_2153,N_805);
and U3213 (N_3213,N_2299,N_1181);
nand U3214 (N_3214,N_819,N_1604);
and U3215 (N_3215,N_771,N_911);
or U3216 (N_3216,N_1132,N_2300);
and U3217 (N_3217,N_547,N_1756);
nor U3218 (N_3218,N_1701,N_37);
nand U3219 (N_3219,N_2150,N_2120);
and U3220 (N_3220,N_1876,N_750);
nor U3221 (N_3221,N_1916,N_1900);
nor U3222 (N_3222,N_1838,N_900);
nand U3223 (N_3223,N_2448,N_836);
nand U3224 (N_3224,N_753,N_1106);
and U3225 (N_3225,N_1217,N_1485);
nor U3226 (N_3226,N_1483,N_1319);
nor U3227 (N_3227,N_1841,N_91);
or U3228 (N_3228,N_2230,N_2432);
nand U3229 (N_3229,N_934,N_36);
nor U3230 (N_3230,N_1808,N_1641);
or U3231 (N_3231,N_738,N_268);
nand U3232 (N_3232,N_957,N_810);
or U3233 (N_3233,N_236,N_1715);
nand U3234 (N_3234,N_213,N_337);
or U3235 (N_3235,N_1740,N_1570);
nand U3236 (N_3236,N_719,N_1326);
or U3237 (N_3237,N_990,N_230);
nand U3238 (N_3238,N_1249,N_1528);
or U3239 (N_3239,N_235,N_1664);
nor U3240 (N_3240,N_2171,N_1964);
or U3241 (N_3241,N_1617,N_1996);
or U3242 (N_3242,N_2452,N_662);
nor U3243 (N_3243,N_289,N_2488);
nand U3244 (N_3244,N_330,N_1390);
or U3245 (N_3245,N_2009,N_1426);
xor U3246 (N_3246,N_524,N_163);
nand U3247 (N_3247,N_2001,N_1339);
and U3248 (N_3248,N_1269,N_2390);
nand U3249 (N_3249,N_545,N_1908);
nor U3250 (N_3250,N_2190,N_2025);
and U3251 (N_3251,N_601,N_338);
nor U3252 (N_3252,N_1638,N_1675);
or U3253 (N_3253,N_245,N_1907);
and U3254 (N_3254,N_1228,N_271);
nor U3255 (N_3255,N_44,N_1631);
nor U3256 (N_3256,N_862,N_1846);
nand U3257 (N_3257,N_258,N_457);
nand U3258 (N_3258,N_875,N_2337);
nand U3259 (N_3259,N_2468,N_1720);
nand U3260 (N_3260,N_2031,N_2287);
or U3261 (N_3261,N_2176,N_1034);
or U3262 (N_3262,N_1398,N_135);
nand U3263 (N_3263,N_1700,N_1861);
nand U3264 (N_3264,N_910,N_530);
nand U3265 (N_3265,N_1536,N_2367);
nand U3266 (N_3266,N_1237,N_2386);
and U3267 (N_3267,N_1206,N_1402);
nand U3268 (N_3268,N_1520,N_606);
or U3269 (N_3269,N_695,N_383);
nand U3270 (N_3270,N_170,N_1108);
or U3271 (N_3271,N_1305,N_664);
nor U3272 (N_3272,N_2282,N_2032);
nand U3273 (N_3273,N_101,N_103);
nand U3274 (N_3274,N_833,N_1295);
and U3275 (N_3275,N_1734,N_701);
nor U3276 (N_3276,N_1650,N_2245);
nand U3277 (N_3277,N_443,N_2044);
nor U3278 (N_3278,N_2361,N_391);
nand U3279 (N_3279,N_1974,N_252);
and U3280 (N_3280,N_2244,N_1783);
nand U3281 (N_3281,N_926,N_1152);
or U3282 (N_3282,N_1166,N_1355);
nor U3283 (N_3283,N_1921,N_2122);
nand U3284 (N_3284,N_1956,N_93);
and U3285 (N_3285,N_1184,N_2039);
or U3286 (N_3286,N_2199,N_718);
xor U3287 (N_3287,N_2496,N_2180);
nand U3288 (N_3288,N_1887,N_952);
nor U3289 (N_3289,N_1250,N_1794);
and U3290 (N_3290,N_1658,N_1139);
xor U3291 (N_3291,N_247,N_1406);
nand U3292 (N_3292,N_1281,N_426);
and U3293 (N_3293,N_2378,N_1585);
and U3294 (N_3294,N_2058,N_117);
or U3295 (N_3295,N_663,N_1600);
nor U3296 (N_3296,N_1299,N_816);
and U3297 (N_3297,N_171,N_1778);
and U3298 (N_3298,N_2372,N_698);
or U3299 (N_3299,N_724,N_381);
nor U3300 (N_3300,N_2038,N_2158);
and U3301 (N_3301,N_749,N_1703);
and U3302 (N_3302,N_1136,N_535);
nor U3303 (N_3303,N_1048,N_2014);
nor U3304 (N_3304,N_1918,N_920);
nor U3305 (N_3305,N_1569,N_2221);
nor U3306 (N_3306,N_520,N_961);
or U3307 (N_3307,N_1886,N_2471);
nor U3308 (N_3308,N_1980,N_592);
or U3309 (N_3309,N_1375,N_2202);
xor U3310 (N_3310,N_622,N_191);
or U3311 (N_3311,N_1636,N_558);
and U3312 (N_3312,N_174,N_1478);
nor U3313 (N_3313,N_1684,N_77);
and U3314 (N_3314,N_148,N_215);
nor U3315 (N_3315,N_1572,N_1871);
or U3316 (N_3316,N_430,N_1187);
nor U3317 (N_3317,N_1385,N_2457);
nand U3318 (N_3318,N_1148,N_1212);
or U3319 (N_3319,N_785,N_1083);
and U3320 (N_3320,N_2166,N_1437);
and U3321 (N_3321,N_1608,N_2425);
nand U3322 (N_3322,N_1707,N_336);
or U3323 (N_3323,N_1522,N_1407);
or U3324 (N_3324,N_1215,N_1297);
nand U3325 (N_3325,N_1901,N_310);
and U3326 (N_3326,N_88,N_741);
and U3327 (N_3327,N_2189,N_248);
or U3328 (N_3328,N_185,N_2159);
nor U3329 (N_3329,N_261,N_1770);
and U3330 (N_3330,N_2046,N_1620);
or U3331 (N_3331,N_449,N_1542);
and U3332 (N_3332,N_2434,N_1007);
nor U3333 (N_3333,N_652,N_525);
nor U3334 (N_3334,N_1270,N_1363);
nor U3335 (N_3335,N_1265,N_1672);
nand U3336 (N_3336,N_2123,N_2373);
xnor U3337 (N_3337,N_1193,N_34);
or U3338 (N_3338,N_1709,N_863);
or U3339 (N_3339,N_1612,N_1310);
or U3340 (N_3340,N_369,N_1189);
or U3341 (N_3341,N_1378,N_1902);
nand U3342 (N_3342,N_1045,N_1399);
or U3343 (N_3343,N_792,N_1274);
and U3344 (N_3344,N_85,N_675);
or U3345 (N_3345,N_1332,N_1246);
and U3346 (N_3346,N_1679,N_1923);
nor U3347 (N_3347,N_2455,N_1349);
nand U3348 (N_3348,N_158,N_1192);
nand U3349 (N_3349,N_715,N_1400);
nor U3350 (N_3350,N_684,N_1022);
nand U3351 (N_3351,N_1753,N_886);
and U3352 (N_3352,N_775,N_962);
nand U3353 (N_3353,N_2207,N_1630);
and U3354 (N_3354,N_2163,N_2350);
nor U3355 (N_3355,N_433,N_2387);
nor U3356 (N_3356,N_1680,N_1351);
and U3357 (N_3357,N_2037,N_925);
nand U3358 (N_3358,N_1118,N_244);
and U3359 (N_3359,N_1890,N_844);
nand U3360 (N_3360,N_493,N_1304);
nand U3361 (N_3361,N_584,N_1550);
or U3362 (N_3362,N_1557,N_768);
nand U3363 (N_3363,N_1819,N_1593);
nand U3364 (N_3364,N_1534,N_29);
nor U3365 (N_3365,N_2017,N_1446);
nor U3366 (N_3366,N_1490,N_218);
and U3367 (N_3367,N_1329,N_404);
nor U3368 (N_3368,N_1625,N_1248);
nand U3369 (N_3369,N_351,N_1268);
nor U3370 (N_3370,N_989,N_761);
nor U3371 (N_3371,N_1117,N_2358);
and U3372 (N_3372,N_469,N_1943);
and U3373 (N_3373,N_444,N_2033);
nand U3374 (N_3374,N_152,N_224);
nor U3375 (N_3375,N_2402,N_1747);
and U3376 (N_3376,N_1678,N_11);
and U3377 (N_3377,N_648,N_81);
nand U3378 (N_3378,N_671,N_1633);
nor U3379 (N_3379,N_692,N_16);
and U3380 (N_3380,N_2160,N_1997);
nand U3381 (N_3381,N_1218,N_201);
or U3382 (N_3382,N_2051,N_2094);
or U3383 (N_3383,N_1714,N_2233);
nand U3384 (N_3384,N_1389,N_615);
and U3385 (N_3385,N_736,N_888);
nor U3386 (N_3386,N_794,N_2124);
nand U3387 (N_3387,N_312,N_883);
nor U3388 (N_3388,N_1050,N_748);
or U3389 (N_3389,N_358,N_2366);
nand U3390 (N_3390,N_2325,N_857);
or U3391 (N_3391,N_2259,N_1768);
or U3392 (N_3392,N_811,N_1056);
nor U3393 (N_3393,N_1503,N_476);
or U3394 (N_3394,N_2018,N_2292);
nand U3395 (N_3395,N_1468,N_1513);
or U3396 (N_3396,N_931,N_1172);
nor U3397 (N_3397,N_1927,N_1386);
or U3398 (N_3398,N_588,N_1911);
or U3399 (N_3399,N_489,N_1278);
or U3400 (N_3400,N_1643,N_693);
and U3401 (N_3401,N_1760,N_1606);
xor U3402 (N_3402,N_1862,N_1580);
nor U3403 (N_3403,N_486,N_89);
or U3404 (N_3404,N_116,N_1345);
nor U3405 (N_3405,N_292,N_2235);
and U3406 (N_3406,N_403,N_1622);
nor U3407 (N_3407,N_534,N_2405);
and U3408 (N_3408,N_631,N_2005);
nand U3409 (N_3409,N_1772,N_238);
and U3410 (N_3410,N_162,N_188);
or U3411 (N_3411,N_1792,N_2103);
nor U3412 (N_3412,N_467,N_658);
or U3413 (N_3413,N_1001,N_427);
nand U3414 (N_3414,N_522,N_2317);
and U3415 (N_3415,N_43,N_821);
nand U3416 (N_3416,N_581,N_1791);
nand U3417 (N_3417,N_1286,N_1692);
and U3418 (N_3418,N_1154,N_1649);
and U3419 (N_3419,N_1244,N_1875);
or U3420 (N_3420,N_448,N_2310);
and U3421 (N_3421,N_2365,N_998);
nand U3422 (N_3422,N_1020,N_2073);
nand U3423 (N_3423,N_1137,N_849);
or U3424 (N_3424,N_691,N_308);
and U3425 (N_3425,N_1082,N_1256);
nor U3426 (N_3426,N_119,N_1758);
or U3427 (N_3427,N_655,N_2251);
nand U3428 (N_3428,N_390,N_1498);
nand U3429 (N_3429,N_2104,N_1273);
nand U3430 (N_3430,N_503,N_994);
or U3431 (N_3431,N_1202,N_1834);
and U3432 (N_3432,N_1325,N_419);
or U3433 (N_3433,N_1644,N_2318);
nand U3434 (N_3434,N_2296,N_1392);
or U3435 (N_3435,N_1947,N_1985);
nand U3436 (N_3436,N_80,N_92);
nor U3437 (N_3437,N_657,N_1337);
or U3438 (N_3438,N_2418,N_1645);
nor U3439 (N_3439,N_340,N_1460);
or U3440 (N_3440,N_1,N_2108);
nand U3441 (N_3441,N_1774,N_885);
and U3442 (N_3442,N_138,N_1309);
nor U3443 (N_3443,N_541,N_1944);
and U3444 (N_3444,N_866,N_573);
and U3445 (N_3445,N_867,N_2279);
nor U3446 (N_3446,N_2141,N_2215);
and U3447 (N_3447,N_610,N_1724);
nand U3448 (N_3448,N_2414,N_595);
nand U3449 (N_3449,N_2193,N_353);
nor U3450 (N_3450,N_537,N_303);
and U3451 (N_3451,N_1362,N_344);
nand U3452 (N_3452,N_1533,N_929);
or U3453 (N_3453,N_1384,N_1293);
or U3454 (N_3454,N_2126,N_1491);
nand U3455 (N_3455,N_125,N_767);
nand U3456 (N_3456,N_1540,N_2275);
nor U3457 (N_3457,N_87,N_578);
or U3458 (N_3458,N_1112,N_2182);
nor U3459 (N_3459,N_364,N_1253);
xor U3460 (N_3460,N_1598,N_1803);
and U3461 (N_3461,N_2147,N_2326);
and U3462 (N_3462,N_1467,N_557);
or U3463 (N_3463,N_155,N_1432);
or U3464 (N_3464,N_2086,N_90);
and U3465 (N_3465,N_937,N_324);
and U3466 (N_3466,N_2248,N_189);
nor U3467 (N_3467,N_968,N_182);
or U3468 (N_3468,N_2429,N_1429);
and U3469 (N_3469,N_1635,N_1751);
nor U3470 (N_3470,N_1648,N_2011);
and U3471 (N_3471,N_2271,N_1704);
nand U3472 (N_3472,N_568,N_511);
nor U3473 (N_3473,N_587,N_2187);
and U3474 (N_3474,N_1693,N_1769);
nor U3475 (N_3475,N_299,N_603);
nor U3476 (N_3476,N_928,N_14);
or U3477 (N_3477,N_333,N_1618);
and U3478 (N_3478,N_772,N_865);
and U3479 (N_3479,N_678,N_1713);
and U3480 (N_3480,N_756,N_566);
and U3481 (N_3481,N_209,N_2156);
nand U3482 (N_3482,N_868,N_75);
and U3483 (N_3483,N_1860,N_2482);
and U3484 (N_3484,N_1497,N_1251);
or U3485 (N_3485,N_2205,N_916);
nand U3486 (N_3486,N_234,N_485);
or U3487 (N_3487,N_1583,N_2218);
or U3488 (N_3488,N_776,N_543);
and U3489 (N_3489,N_264,N_220);
and U3490 (N_3490,N_877,N_1951);
or U3491 (N_3491,N_307,N_2359);
or U3492 (N_3492,N_702,N_320);
nor U3493 (N_3493,N_1484,N_412);
or U3494 (N_3494,N_1730,N_1430);
and U3495 (N_3495,N_424,N_2075);
and U3496 (N_3496,N_1628,N_2315);
nor U3497 (N_3497,N_1652,N_223);
and U3498 (N_3498,N_1340,N_1696);
nand U3499 (N_3499,N_122,N_1413);
and U3500 (N_3500,N_806,N_1164);
and U3501 (N_3501,N_755,N_2360);
nand U3502 (N_3502,N_563,N_841);
and U3503 (N_3503,N_1647,N_1560);
or U3504 (N_3504,N_2217,N_2368);
nor U3505 (N_3505,N_943,N_575);
nand U3506 (N_3506,N_1654,N_1695);
and U3507 (N_3507,N_2494,N_1788);
and U3508 (N_3508,N_95,N_1186);
and U3509 (N_3509,N_621,N_1987);
nor U3510 (N_3510,N_179,N_298);
nor U3511 (N_3511,N_2036,N_781);
nor U3512 (N_3512,N_611,N_2106);
nand U3513 (N_3513,N_2154,N_770);
nor U3514 (N_3514,N_800,N_2427);
nand U3515 (N_3515,N_1143,N_1850);
nand U3516 (N_3516,N_1653,N_1832);
nor U3517 (N_3517,N_2375,N_196);
or U3518 (N_3518,N_2155,N_1290);
nor U3519 (N_3519,N_538,N_70);
or U3520 (N_3520,N_2003,N_1616);
or U3521 (N_3521,N_786,N_2376);
nand U3522 (N_3522,N_1312,N_1047);
or U3523 (N_3523,N_1950,N_742);
and U3524 (N_3524,N_478,N_2406);
nand U3525 (N_3525,N_2236,N_1959);
nand U3526 (N_3526,N_1260,N_801);
nor U3527 (N_3527,N_1553,N_2137);
nor U3528 (N_3528,N_2295,N_688);
nor U3529 (N_3529,N_1594,N_1480);
or U3530 (N_3530,N_2064,N_1072);
and U3531 (N_3531,N_705,N_645);
and U3532 (N_3532,N_1539,N_850);
or U3533 (N_3533,N_1086,N_1712);
nor U3534 (N_3534,N_407,N_1787);
nor U3535 (N_3535,N_2093,N_1651);
nand U3536 (N_3536,N_2341,N_370);
or U3537 (N_3537,N_1125,N_912);
and U3538 (N_3538,N_326,N_1369);
nand U3539 (N_3539,N_195,N_13);
or U3540 (N_3540,N_41,N_1169);
nand U3541 (N_3541,N_840,N_2356);
nand U3542 (N_3542,N_1330,N_1103);
and U3543 (N_3543,N_2220,N_984);
or U3544 (N_3544,N_1961,N_1789);
nor U3545 (N_3545,N_168,N_1316);
and U3546 (N_3546,N_1626,N_614);
or U3547 (N_3547,N_1200,N_680);
or U3548 (N_3548,N_2437,N_2055);
nand U3549 (N_3549,N_394,N_1023);
and U3550 (N_3550,N_685,N_348);
nor U3551 (N_3551,N_1049,N_439);
or U3552 (N_3552,N_68,N_2219);
or U3553 (N_3553,N_1271,N_84);
nor U3554 (N_3554,N_747,N_1611);
nand U3555 (N_3555,N_2203,N_1940);
and U3556 (N_3556,N_2363,N_1301);
and U3557 (N_3557,N_149,N_2320);
and U3558 (N_3558,N_2081,N_1111);
nand U3559 (N_3559,N_1311,N_1547);
or U3560 (N_3560,N_1448,N_2336);
nand U3561 (N_3561,N_746,N_133);
nand U3562 (N_3562,N_2302,N_1296);
or U3563 (N_3563,N_2083,N_54);
or U3564 (N_3564,N_1095,N_1011);
nor U3565 (N_3565,N_1666,N_1502);
nor U3566 (N_3566,N_1171,N_2223);
or U3567 (N_3567,N_1214,N_1168);
nand U3568 (N_3568,N_845,N_823);
and U3569 (N_3569,N_1686,N_1307);
and U3570 (N_3570,N_627,N_1619);
nand U3571 (N_3571,N_1472,N_1885);
nand U3572 (N_3572,N_1134,N_45);
and U3573 (N_3573,N_2369,N_1208);
and U3574 (N_3574,N_1869,N_2200);
nor U3575 (N_3575,N_349,N_1130);
nor U3576 (N_3576,N_546,N_341);
and U3577 (N_3577,N_56,N_632);
and U3578 (N_3578,N_2485,N_2164);
nor U3579 (N_3579,N_1474,N_410);
nand U3580 (N_3580,N_1126,N_110);
or U3581 (N_3581,N_1493,N_1195);
nand U3582 (N_3582,N_2237,N_1035);
or U3583 (N_3583,N_1603,N_2351);
or U3584 (N_3584,N_508,N_760);
or U3585 (N_3585,N_765,N_762);
and U3586 (N_3586,N_436,N_193);
nand U3587 (N_3587,N_817,N_1039);
or U3588 (N_3588,N_1946,N_1388);
nand U3589 (N_3589,N_1054,N_198);
nand U3590 (N_3590,N_915,N_2121);
nand U3591 (N_3591,N_1615,N_1800);
or U3592 (N_3592,N_2497,N_1412);
and U3593 (N_3593,N_384,N_710);
nand U3594 (N_3594,N_871,N_2041);
or U3595 (N_3595,N_2319,N_1592);
and U3596 (N_3596,N_1476,N_33);
nand U3597 (N_3597,N_1523,N_2454);
and U3598 (N_3598,N_1489,N_1101);
or U3599 (N_3599,N_1461,N_808);
or U3600 (N_3600,N_255,N_1814);
and U3601 (N_3601,N_778,N_856);
or U3602 (N_3602,N_974,N_1577);
nor U3603 (N_3603,N_194,N_1710);
nand U3604 (N_3604,N_739,N_1354);
and U3605 (N_3605,N_1546,N_2430);
or U3606 (N_3606,N_2157,N_909);
and U3607 (N_3607,N_972,N_2174);
and U3608 (N_3608,N_1080,N_468);
nand U3609 (N_3609,N_1931,N_787);
nor U3610 (N_3610,N_199,N_1091);
nor U3611 (N_3611,N_382,N_208);
nand U3612 (N_3612,N_804,N_1453);
and U3613 (N_3613,N_2131,N_225);
or U3614 (N_3614,N_830,N_921);
or U3615 (N_3615,N_1066,N_161);
nand U3616 (N_3616,N_432,N_605);
or U3617 (N_3617,N_482,N_795);
and U3618 (N_3618,N_2114,N_807);
and U3619 (N_3619,N_1258,N_1173);
nor U3620 (N_3620,N_646,N_375);
nor U3621 (N_3621,N_317,N_309);
or U3622 (N_3622,N_1128,N_1971);
nand U3623 (N_3623,N_1288,N_1254);
or U3624 (N_3624,N_2262,N_1287);
nand U3625 (N_3625,N_301,N_2280);
nand U3626 (N_3626,N_1262,N_1531);
nor U3627 (N_3627,N_2291,N_1667);
and U3628 (N_3628,N_1705,N_502);
or U3629 (N_3629,N_123,N_1226);
and U3630 (N_3630,N_60,N_181);
or U3631 (N_3631,N_495,N_879);
and U3632 (N_3632,N_1706,N_459);
or U3633 (N_3633,N_2169,N_411);
nand U3634 (N_3634,N_1087,N_2030);
nor U3635 (N_3635,N_1487,N_818);
nand U3636 (N_3636,N_4,N_282);
nand U3637 (N_3637,N_697,N_1464);
nand U3638 (N_3638,N_619,N_2022);
nor U3639 (N_3639,N_643,N_186);
nand U3640 (N_3640,N_2249,N_2100);
nand U3641 (N_3641,N_2396,N_1793);
nor U3642 (N_3642,N_734,N_1809);
nand U3643 (N_3643,N_157,N_1749);
or U3644 (N_3644,N_1127,N_967);
or U3645 (N_3645,N_339,N_2464);
and U3646 (N_3646,N_2179,N_988);
or U3647 (N_3647,N_1482,N_1801);
and U3648 (N_3648,N_1882,N_465);
nor U3649 (N_3649,N_429,N_446);
or U3650 (N_3650,N_2332,N_2460);
and U3651 (N_3651,N_1873,N_197);
nand U3652 (N_3652,N_1428,N_803);
or U3653 (N_3653,N_1141,N_2145);
or U3654 (N_3654,N_1823,N_1805);
and U3655 (N_3655,N_47,N_796);
and U3656 (N_3656,N_1346,N_941);
nand U3657 (N_3657,N_1708,N_699);
and U3658 (N_3658,N_1471,N_813);
nand U3659 (N_3659,N_1591,N_1191);
or U3660 (N_3660,N_115,N_1085);
and U3661 (N_3661,N_2067,N_2353);
nand U3662 (N_3662,N_894,N_1563);
and U3663 (N_3663,N_1131,N_1945);
or U3664 (N_3664,N_212,N_1627);
nand U3665 (N_3665,N_1320,N_1967);
nand U3666 (N_3666,N_939,N_714);
or U3667 (N_3667,N_1587,N_2370);
nor U3668 (N_3668,N_2116,N_1574);
and U3669 (N_3669,N_2403,N_2399);
nor U3670 (N_3670,N_589,N_1053);
nor U3671 (N_3671,N_1991,N_623);
and U3672 (N_3672,N_434,N_105);
nor U3673 (N_3673,N_1745,N_2228);
nor U3674 (N_3674,N_1122,N_173);
nand U3675 (N_3675,N_141,N_633);
nand U3676 (N_3676,N_2079,N_2144);
or U3677 (N_3677,N_858,N_438);
and U3678 (N_3678,N_2357,N_2212);
and U3679 (N_3679,N_372,N_512);
or U3680 (N_3680,N_74,N_2477);
nand U3681 (N_3681,N_30,N_456);
nor U3682 (N_3682,N_1455,N_277);
nor U3683 (N_3683,N_1451,N_782);
nand U3684 (N_3684,N_1738,N_368);
nand U3685 (N_3685,N_2301,N_1729);
or U3686 (N_3686,N_751,N_562);
and U3687 (N_3687,N_1962,N_2461);
xnor U3688 (N_3688,N_948,N_2422);
or U3689 (N_3689,N_2026,N_1847);
nand U3690 (N_3690,N_1837,N_2281);
or U3691 (N_3691,N_1387,N_2053);
and U3692 (N_3692,N_1807,N_1905);
or U3693 (N_3693,N_203,N_2487);
nand U3694 (N_3694,N_2029,N_650);
nand U3695 (N_3695,N_2272,N_2495);
nor U3696 (N_3696,N_1427,N_1452);
and U3697 (N_3697,N_1578,N_2115);
or U3698 (N_3698,N_2331,N_1321);
nor U3699 (N_3699,N_1779,N_570);
nand U3700 (N_3700,N_263,N_1629);
nor U3701 (N_3701,N_417,N_460);
nor U3702 (N_3702,N_1994,N_922);
or U3703 (N_3703,N_1261,N_1588);
nor U3704 (N_3704,N_2130,N_1639);
nand U3705 (N_3705,N_902,N_992);
nand U3706 (N_3706,N_2409,N_1565);
nor U3707 (N_3707,N_869,N_1839);
or U3708 (N_3708,N_1475,N_551);
nand U3709 (N_3709,N_2013,N_159);
and U3710 (N_3710,N_1613,N_1454);
or U3711 (N_3711,N_1203,N_725);
or U3712 (N_3712,N_1757,N_2345);
nand U3713 (N_3713,N_1763,N_2416);
and U3714 (N_3714,N_1352,N_1889);
nor U3715 (N_3715,N_1632,N_1642);
and U3716 (N_3716,N_579,N_1535);
nand U3717 (N_3717,N_1737,N_933);
nor U3718 (N_3718,N_1614,N_1227);
nor U3719 (N_3719,N_20,N_1802);
or U3720 (N_3720,N_1824,N_628);
nand U3721 (N_3721,N_352,N_1396);
or U3722 (N_3722,N_124,N_2377);
or U3723 (N_3723,N_2431,N_634);
nand U3724 (N_3724,N_2239,N_907);
and U3725 (N_3725,N_791,N_2111);
nor U3726 (N_3726,N_993,N_1197);
or U3727 (N_3727,N_1733,N_1044);
or U3728 (N_3728,N_859,N_1229);
nor U3729 (N_3729,N_2435,N_1306);
nand U3730 (N_3730,N_1343,N_814);
nand U3731 (N_3731,N_2255,N_1240);
and U3732 (N_3732,N_1790,N_774);
nor U3733 (N_3733,N_249,N_2265);
and U3734 (N_3734,N_820,N_274);
and U3735 (N_3735,N_256,N_1939);
nor U3736 (N_3736,N_1123,N_1932);
nand U3737 (N_3737,N_1179,N_2213);
and U3738 (N_3738,N_583,N_689);
nand U3739 (N_3739,N_455,N_1910);
nand U3740 (N_3740,N_694,N_2258);
nand U3741 (N_3741,N_2463,N_1151);
nor U3742 (N_3742,N_1245,N_53);
nand U3743 (N_3743,N_1156,N_488);
or U3744 (N_3744,N_1676,N_1038);
or U3745 (N_3745,N_1881,N_1865);
nor U3746 (N_3746,N_1899,N_1529);
and U3747 (N_3747,N_1694,N_1555);
and U3748 (N_3748,N_2445,N_378);
nand U3749 (N_3749,N_732,N_151);
or U3750 (N_3750,N_881,N_35);
and U3751 (N_3751,N_1331,N_2009);
nor U3752 (N_3752,N_1066,N_1181);
nand U3753 (N_3753,N_1820,N_732);
or U3754 (N_3754,N_615,N_843);
nor U3755 (N_3755,N_1236,N_983);
nand U3756 (N_3756,N_417,N_1480);
and U3757 (N_3757,N_2073,N_669);
nor U3758 (N_3758,N_1079,N_1073);
nor U3759 (N_3759,N_2090,N_2344);
and U3760 (N_3760,N_680,N_1531);
nand U3761 (N_3761,N_276,N_435);
and U3762 (N_3762,N_240,N_852);
nor U3763 (N_3763,N_385,N_2181);
nor U3764 (N_3764,N_24,N_1079);
nor U3765 (N_3765,N_1384,N_2422);
nand U3766 (N_3766,N_912,N_843);
or U3767 (N_3767,N_1509,N_1597);
nor U3768 (N_3768,N_650,N_98);
nand U3769 (N_3769,N_1904,N_1913);
and U3770 (N_3770,N_1506,N_1570);
nor U3771 (N_3771,N_2328,N_1347);
or U3772 (N_3772,N_387,N_1988);
or U3773 (N_3773,N_1116,N_2137);
and U3774 (N_3774,N_929,N_2010);
or U3775 (N_3775,N_1782,N_1727);
nor U3776 (N_3776,N_373,N_909);
and U3777 (N_3777,N_2057,N_2235);
nand U3778 (N_3778,N_556,N_2197);
nor U3779 (N_3779,N_1943,N_1705);
nand U3780 (N_3780,N_2414,N_2381);
and U3781 (N_3781,N_1718,N_1295);
nand U3782 (N_3782,N_868,N_2359);
nor U3783 (N_3783,N_994,N_63);
or U3784 (N_3784,N_2242,N_1311);
and U3785 (N_3785,N_929,N_1096);
or U3786 (N_3786,N_768,N_1245);
nor U3787 (N_3787,N_1428,N_1019);
or U3788 (N_3788,N_281,N_1020);
nor U3789 (N_3789,N_1276,N_1545);
or U3790 (N_3790,N_1960,N_1061);
nand U3791 (N_3791,N_2116,N_1550);
nand U3792 (N_3792,N_1361,N_2073);
nor U3793 (N_3793,N_558,N_1663);
and U3794 (N_3794,N_794,N_1409);
nor U3795 (N_3795,N_2211,N_1247);
or U3796 (N_3796,N_2253,N_2367);
nand U3797 (N_3797,N_437,N_443);
and U3798 (N_3798,N_1319,N_1439);
and U3799 (N_3799,N_2181,N_1365);
nand U3800 (N_3800,N_1487,N_1087);
xor U3801 (N_3801,N_2070,N_12);
and U3802 (N_3802,N_1905,N_1157);
or U3803 (N_3803,N_2175,N_365);
nor U3804 (N_3804,N_2131,N_2047);
nand U3805 (N_3805,N_1421,N_1517);
nor U3806 (N_3806,N_1914,N_2113);
or U3807 (N_3807,N_2310,N_2079);
nand U3808 (N_3808,N_1939,N_2203);
nor U3809 (N_3809,N_1919,N_1958);
nor U3810 (N_3810,N_7,N_731);
nor U3811 (N_3811,N_33,N_1071);
nand U3812 (N_3812,N_2167,N_2189);
or U3813 (N_3813,N_2370,N_1642);
or U3814 (N_3814,N_1641,N_790);
nand U3815 (N_3815,N_465,N_298);
or U3816 (N_3816,N_21,N_39);
and U3817 (N_3817,N_296,N_139);
or U3818 (N_3818,N_2010,N_2152);
nor U3819 (N_3819,N_458,N_968);
or U3820 (N_3820,N_480,N_1853);
and U3821 (N_3821,N_813,N_1579);
or U3822 (N_3822,N_2473,N_1158);
nand U3823 (N_3823,N_509,N_819);
nand U3824 (N_3824,N_1861,N_674);
and U3825 (N_3825,N_2110,N_1422);
and U3826 (N_3826,N_12,N_1712);
nor U3827 (N_3827,N_128,N_1670);
xnor U3828 (N_3828,N_1585,N_733);
nand U3829 (N_3829,N_1913,N_2080);
nor U3830 (N_3830,N_1300,N_438);
nand U3831 (N_3831,N_1621,N_277);
or U3832 (N_3832,N_101,N_829);
nand U3833 (N_3833,N_1101,N_1432);
or U3834 (N_3834,N_447,N_628);
xor U3835 (N_3835,N_625,N_1605);
nor U3836 (N_3836,N_1174,N_1904);
and U3837 (N_3837,N_1688,N_641);
or U3838 (N_3838,N_1352,N_215);
or U3839 (N_3839,N_699,N_2334);
or U3840 (N_3840,N_1717,N_337);
and U3841 (N_3841,N_1094,N_1900);
and U3842 (N_3842,N_280,N_1003);
and U3843 (N_3843,N_1750,N_809);
and U3844 (N_3844,N_2004,N_2086);
nand U3845 (N_3845,N_671,N_1175);
nor U3846 (N_3846,N_1040,N_2278);
nor U3847 (N_3847,N_1185,N_1558);
or U3848 (N_3848,N_554,N_1390);
nand U3849 (N_3849,N_1413,N_1954);
or U3850 (N_3850,N_81,N_336);
or U3851 (N_3851,N_289,N_1252);
nand U3852 (N_3852,N_1070,N_1781);
or U3853 (N_3853,N_789,N_975);
or U3854 (N_3854,N_1942,N_1854);
and U3855 (N_3855,N_176,N_1126);
or U3856 (N_3856,N_892,N_1826);
and U3857 (N_3857,N_1971,N_2100);
and U3858 (N_3858,N_897,N_485);
or U3859 (N_3859,N_2030,N_883);
nor U3860 (N_3860,N_205,N_1059);
or U3861 (N_3861,N_535,N_1117);
nand U3862 (N_3862,N_1879,N_698);
and U3863 (N_3863,N_1815,N_2114);
or U3864 (N_3864,N_306,N_875);
nand U3865 (N_3865,N_883,N_1349);
nand U3866 (N_3866,N_1827,N_1619);
nand U3867 (N_3867,N_852,N_1798);
nor U3868 (N_3868,N_1085,N_760);
nor U3869 (N_3869,N_818,N_1283);
nor U3870 (N_3870,N_529,N_1473);
and U3871 (N_3871,N_688,N_2154);
nand U3872 (N_3872,N_511,N_1013);
or U3873 (N_3873,N_1149,N_79);
or U3874 (N_3874,N_516,N_728);
nor U3875 (N_3875,N_2129,N_2076);
nand U3876 (N_3876,N_54,N_246);
nor U3877 (N_3877,N_1114,N_1555);
nand U3878 (N_3878,N_801,N_1895);
and U3879 (N_3879,N_489,N_1578);
or U3880 (N_3880,N_745,N_2046);
and U3881 (N_3881,N_2480,N_803);
and U3882 (N_3882,N_1479,N_2359);
or U3883 (N_3883,N_1560,N_240);
nand U3884 (N_3884,N_2078,N_811);
or U3885 (N_3885,N_1459,N_748);
nor U3886 (N_3886,N_1392,N_1524);
nand U3887 (N_3887,N_46,N_1130);
nor U3888 (N_3888,N_25,N_1712);
nor U3889 (N_3889,N_398,N_2320);
and U3890 (N_3890,N_1699,N_2266);
nor U3891 (N_3891,N_800,N_301);
nor U3892 (N_3892,N_1651,N_2013);
and U3893 (N_3893,N_1430,N_2028);
nand U3894 (N_3894,N_2189,N_864);
and U3895 (N_3895,N_1016,N_1263);
nor U3896 (N_3896,N_593,N_2486);
and U3897 (N_3897,N_1551,N_1206);
nor U3898 (N_3898,N_1590,N_207);
nand U3899 (N_3899,N_954,N_158);
nor U3900 (N_3900,N_528,N_1576);
nor U3901 (N_3901,N_1031,N_1844);
or U3902 (N_3902,N_1969,N_1280);
nand U3903 (N_3903,N_2122,N_385);
nand U3904 (N_3904,N_537,N_1998);
nand U3905 (N_3905,N_1502,N_353);
or U3906 (N_3906,N_1364,N_22);
nor U3907 (N_3907,N_1455,N_448);
nor U3908 (N_3908,N_19,N_657);
nor U3909 (N_3909,N_22,N_808);
nand U3910 (N_3910,N_680,N_354);
or U3911 (N_3911,N_1257,N_620);
and U3912 (N_3912,N_2375,N_55);
nand U3913 (N_3913,N_1548,N_459);
nand U3914 (N_3914,N_111,N_2214);
nor U3915 (N_3915,N_1529,N_1704);
nor U3916 (N_3916,N_625,N_1734);
and U3917 (N_3917,N_1740,N_1733);
nor U3918 (N_3918,N_809,N_1181);
nand U3919 (N_3919,N_1467,N_1964);
and U3920 (N_3920,N_2332,N_702);
or U3921 (N_3921,N_1823,N_190);
and U3922 (N_3922,N_123,N_258);
nor U3923 (N_3923,N_2258,N_963);
nor U3924 (N_3924,N_2409,N_1479);
nand U3925 (N_3925,N_882,N_34);
nor U3926 (N_3926,N_2030,N_370);
nor U3927 (N_3927,N_2476,N_2045);
or U3928 (N_3928,N_1069,N_460);
nor U3929 (N_3929,N_2124,N_1552);
or U3930 (N_3930,N_2302,N_1559);
nor U3931 (N_3931,N_163,N_385);
and U3932 (N_3932,N_1858,N_988);
nor U3933 (N_3933,N_652,N_1316);
or U3934 (N_3934,N_117,N_1099);
nor U3935 (N_3935,N_844,N_432);
nor U3936 (N_3936,N_2086,N_1606);
and U3937 (N_3937,N_2360,N_2047);
and U3938 (N_3938,N_593,N_986);
and U3939 (N_3939,N_2095,N_1206);
or U3940 (N_3940,N_1442,N_1195);
and U3941 (N_3941,N_870,N_876);
or U3942 (N_3942,N_986,N_610);
nand U3943 (N_3943,N_1632,N_1510);
nor U3944 (N_3944,N_839,N_931);
or U3945 (N_3945,N_1916,N_902);
nor U3946 (N_3946,N_1082,N_1886);
nor U3947 (N_3947,N_1058,N_1509);
and U3948 (N_3948,N_2129,N_1962);
nand U3949 (N_3949,N_1328,N_2171);
nand U3950 (N_3950,N_2254,N_2066);
or U3951 (N_3951,N_2065,N_2254);
nor U3952 (N_3952,N_2275,N_541);
or U3953 (N_3953,N_1305,N_377);
nand U3954 (N_3954,N_1849,N_786);
or U3955 (N_3955,N_1993,N_1308);
xnor U3956 (N_3956,N_1567,N_131);
nor U3957 (N_3957,N_353,N_543);
nor U3958 (N_3958,N_535,N_1277);
nor U3959 (N_3959,N_2289,N_938);
or U3960 (N_3960,N_671,N_1739);
and U3961 (N_3961,N_686,N_1128);
and U3962 (N_3962,N_919,N_2298);
nand U3963 (N_3963,N_1429,N_2016);
nand U3964 (N_3964,N_1360,N_354);
nand U3965 (N_3965,N_1151,N_1868);
or U3966 (N_3966,N_1031,N_1965);
nand U3967 (N_3967,N_1490,N_187);
nand U3968 (N_3968,N_1320,N_1852);
nor U3969 (N_3969,N_1261,N_1891);
nor U3970 (N_3970,N_1340,N_2202);
nor U3971 (N_3971,N_946,N_49);
or U3972 (N_3972,N_1290,N_29);
and U3973 (N_3973,N_975,N_261);
and U3974 (N_3974,N_44,N_875);
nand U3975 (N_3975,N_809,N_1887);
nor U3976 (N_3976,N_841,N_748);
xnor U3977 (N_3977,N_1575,N_943);
or U3978 (N_3978,N_2410,N_1102);
or U3979 (N_3979,N_676,N_225);
nor U3980 (N_3980,N_457,N_1588);
or U3981 (N_3981,N_341,N_904);
nand U3982 (N_3982,N_1591,N_2418);
nor U3983 (N_3983,N_2327,N_421);
or U3984 (N_3984,N_2119,N_33);
nor U3985 (N_3985,N_855,N_66);
nor U3986 (N_3986,N_907,N_601);
nand U3987 (N_3987,N_2360,N_2018);
and U3988 (N_3988,N_2479,N_1347);
nor U3989 (N_3989,N_59,N_313);
nand U3990 (N_3990,N_1037,N_1779);
and U3991 (N_3991,N_659,N_2082);
or U3992 (N_3992,N_1283,N_1996);
nand U3993 (N_3993,N_1279,N_465);
and U3994 (N_3994,N_1288,N_1603);
nor U3995 (N_3995,N_2401,N_1712);
nand U3996 (N_3996,N_1846,N_891);
nand U3997 (N_3997,N_2337,N_672);
nor U3998 (N_3998,N_1075,N_528);
nor U3999 (N_3999,N_812,N_176);
and U4000 (N_4000,N_380,N_918);
and U4001 (N_4001,N_1393,N_930);
and U4002 (N_4002,N_66,N_195);
nor U4003 (N_4003,N_1293,N_1098);
or U4004 (N_4004,N_64,N_1420);
nand U4005 (N_4005,N_2131,N_2266);
nor U4006 (N_4006,N_825,N_1295);
and U4007 (N_4007,N_506,N_36);
nand U4008 (N_4008,N_2153,N_984);
or U4009 (N_4009,N_1589,N_1411);
and U4010 (N_4010,N_2075,N_664);
and U4011 (N_4011,N_2151,N_841);
and U4012 (N_4012,N_122,N_95);
nor U4013 (N_4013,N_787,N_1261);
nand U4014 (N_4014,N_1934,N_1345);
nor U4015 (N_4015,N_536,N_81);
and U4016 (N_4016,N_2484,N_176);
or U4017 (N_4017,N_520,N_2194);
nor U4018 (N_4018,N_176,N_2206);
and U4019 (N_4019,N_589,N_1089);
or U4020 (N_4020,N_728,N_1051);
or U4021 (N_4021,N_2287,N_1888);
nand U4022 (N_4022,N_1365,N_1114);
nor U4023 (N_4023,N_2430,N_2081);
and U4024 (N_4024,N_1142,N_724);
and U4025 (N_4025,N_1326,N_1876);
or U4026 (N_4026,N_195,N_427);
or U4027 (N_4027,N_2084,N_2281);
nor U4028 (N_4028,N_96,N_914);
nor U4029 (N_4029,N_21,N_1412);
nor U4030 (N_4030,N_517,N_2481);
and U4031 (N_4031,N_74,N_115);
nor U4032 (N_4032,N_1410,N_639);
or U4033 (N_4033,N_947,N_1205);
nand U4034 (N_4034,N_1477,N_1467);
or U4035 (N_4035,N_1335,N_988);
and U4036 (N_4036,N_738,N_188);
nand U4037 (N_4037,N_2103,N_1770);
nand U4038 (N_4038,N_1750,N_734);
nor U4039 (N_4039,N_1084,N_831);
or U4040 (N_4040,N_1067,N_651);
and U4041 (N_4041,N_575,N_638);
and U4042 (N_4042,N_726,N_1157);
nor U4043 (N_4043,N_1232,N_785);
nor U4044 (N_4044,N_1890,N_971);
and U4045 (N_4045,N_334,N_566);
nand U4046 (N_4046,N_5,N_1497);
and U4047 (N_4047,N_66,N_1318);
nor U4048 (N_4048,N_1356,N_539);
and U4049 (N_4049,N_1080,N_2208);
nor U4050 (N_4050,N_90,N_1599);
nand U4051 (N_4051,N_543,N_1005);
and U4052 (N_4052,N_306,N_148);
and U4053 (N_4053,N_814,N_1971);
nor U4054 (N_4054,N_429,N_2433);
nand U4055 (N_4055,N_673,N_1063);
nor U4056 (N_4056,N_1620,N_919);
and U4057 (N_4057,N_1160,N_2063);
nor U4058 (N_4058,N_153,N_1486);
nand U4059 (N_4059,N_1162,N_45);
or U4060 (N_4060,N_898,N_2044);
nand U4061 (N_4061,N_1950,N_2148);
or U4062 (N_4062,N_275,N_831);
nand U4063 (N_4063,N_1446,N_1985);
nor U4064 (N_4064,N_1298,N_34);
and U4065 (N_4065,N_289,N_2424);
or U4066 (N_4066,N_1137,N_2214);
nand U4067 (N_4067,N_948,N_1035);
nand U4068 (N_4068,N_1889,N_714);
and U4069 (N_4069,N_619,N_2355);
nand U4070 (N_4070,N_756,N_492);
nand U4071 (N_4071,N_1121,N_2263);
nand U4072 (N_4072,N_127,N_405);
nor U4073 (N_4073,N_621,N_1096);
nor U4074 (N_4074,N_435,N_1085);
nand U4075 (N_4075,N_2182,N_1183);
and U4076 (N_4076,N_418,N_334);
nand U4077 (N_4077,N_1031,N_1914);
and U4078 (N_4078,N_802,N_272);
nand U4079 (N_4079,N_737,N_422);
nor U4080 (N_4080,N_1491,N_2014);
or U4081 (N_4081,N_829,N_815);
or U4082 (N_4082,N_2450,N_1476);
nand U4083 (N_4083,N_896,N_2478);
nand U4084 (N_4084,N_1549,N_755);
nor U4085 (N_4085,N_1207,N_2246);
nand U4086 (N_4086,N_630,N_755);
or U4087 (N_4087,N_1167,N_1704);
or U4088 (N_4088,N_1529,N_953);
nor U4089 (N_4089,N_1750,N_592);
nor U4090 (N_4090,N_2313,N_128);
nand U4091 (N_4091,N_51,N_2336);
nand U4092 (N_4092,N_223,N_1210);
or U4093 (N_4093,N_2109,N_257);
or U4094 (N_4094,N_1183,N_2082);
nor U4095 (N_4095,N_486,N_2438);
nor U4096 (N_4096,N_253,N_1419);
or U4097 (N_4097,N_1103,N_89);
and U4098 (N_4098,N_2332,N_1054);
nor U4099 (N_4099,N_1124,N_2125);
nor U4100 (N_4100,N_1938,N_1397);
and U4101 (N_4101,N_1323,N_488);
or U4102 (N_4102,N_1050,N_2006);
nand U4103 (N_4103,N_2139,N_1816);
and U4104 (N_4104,N_226,N_969);
nand U4105 (N_4105,N_585,N_1856);
nand U4106 (N_4106,N_1373,N_119);
or U4107 (N_4107,N_789,N_2474);
and U4108 (N_4108,N_1735,N_2349);
and U4109 (N_4109,N_408,N_521);
and U4110 (N_4110,N_929,N_272);
nand U4111 (N_4111,N_581,N_1907);
or U4112 (N_4112,N_1526,N_818);
and U4113 (N_4113,N_811,N_1308);
nand U4114 (N_4114,N_1384,N_811);
nor U4115 (N_4115,N_774,N_758);
and U4116 (N_4116,N_968,N_143);
nor U4117 (N_4117,N_2441,N_495);
or U4118 (N_4118,N_339,N_67);
and U4119 (N_4119,N_1541,N_1701);
or U4120 (N_4120,N_2460,N_2139);
and U4121 (N_4121,N_2313,N_928);
and U4122 (N_4122,N_846,N_418);
and U4123 (N_4123,N_1057,N_1704);
and U4124 (N_4124,N_109,N_2012);
or U4125 (N_4125,N_1313,N_1783);
or U4126 (N_4126,N_426,N_466);
nor U4127 (N_4127,N_811,N_2204);
or U4128 (N_4128,N_749,N_1908);
nand U4129 (N_4129,N_2049,N_1750);
and U4130 (N_4130,N_699,N_860);
and U4131 (N_4131,N_1163,N_2347);
xnor U4132 (N_4132,N_2112,N_2018);
nand U4133 (N_4133,N_555,N_975);
or U4134 (N_4134,N_299,N_1876);
nand U4135 (N_4135,N_1953,N_1979);
and U4136 (N_4136,N_2406,N_2196);
nor U4137 (N_4137,N_1038,N_361);
nand U4138 (N_4138,N_2107,N_849);
or U4139 (N_4139,N_1031,N_865);
and U4140 (N_4140,N_870,N_1044);
nand U4141 (N_4141,N_107,N_1968);
and U4142 (N_4142,N_2227,N_2085);
nor U4143 (N_4143,N_1772,N_1324);
and U4144 (N_4144,N_443,N_1971);
xor U4145 (N_4145,N_197,N_473);
nor U4146 (N_4146,N_1276,N_2486);
nand U4147 (N_4147,N_2262,N_2496);
nor U4148 (N_4148,N_2081,N_2277);
and U4149 (N_4149,N_890,N_2443);
nand U4150 (N_4150,N_1075,N_1525);
nand U4151 (N_4151,N_1239,N_1879);
and U4152 (N_4152,N_1516,N_362);
and U4153 (N_4153,N_1949,N_2123);
and U4154 (N_4154,N_783,N_2370);
and U4155 (N_4155,N_1562,N_966);
or U4156 (N_4156,N_328,N_1700);
and U4157 (N_4157,N_2160,N_1911);
or U4158 (N_4158,N_1566,N_195);
nand U4159 (N_4159,N_724,N_217);
and U4160 (N_4160,N_1458,N_500);
or U4161 (N_4161,N_564,N_1633);
nand U4162 (N_4162,N_1465,N_1339);
and U4163 (N_4163,N_1124,N_1799);
or U4164 (N_4164,N_2034,N_457);
or U4165 (N_4165,N_721,N_2006);
and U4166 (N_4166,N_1435,N_861);
and U4167 (N_4167,N_1270,N_2383);
or U4168 (N_4168,N_454,N_1922);
nand U4169 (N_4169,N_2013,N_529);
nand U4170 (N_4170,N_2066,N_1980);
and U4171 (N_4171,N_702,N_1579);
nand U4172 (N_4172,N_1107,N_333);
nand U4173 (N_4173,N_2324,N_542);
and U4174 (N_4174,N_48,N_1796);
or U4175 (N_4175,N_1385,N_2078);
nor U4176 (N_4176,N_407,N_1617);
nand U4177 (N_4177,N_1340,N_173);
nand U4178 (N_4178,N_1120,N_1434);
and U4179 (N_4179,N_429,N_998);
nor U4180 (N_4180,N_110,N_925);
and U4181 (N_4181,N_541,N_569);
xnor U4182 (N_4182,N_2462,N_146);
and U4183 (N_4183,N_1783,N_172);
nand U4184 (N_4184,N_1900,N_660);
nand U4185 (N_4185,N_767,N_1264);
nand U4186 (N_4186,N_118,N_92);
and U4187 (N_4187,N_1241,N_1197);
nand U4188 (N_4188,N_46,N_993);
nand U4189 (N_4189,N_333,N_1525);
nor U4190 (N_4190,N_2021,N_1916);
and U4191 (N_4191,N_82,N_2014);
and U4192 (N_4192,N_2482,N_2069);
nand U4193 (N_4193,N_405,N_106);
or U4194 (N_4194,N_804,N_1855);
and U4195 (N_4195,N_1789,N_1175);
or U4196 (N_4196,N_1103,N_2296);
and U4197 (N_4197,N_814,N_1112);
nor U4198 (N_4198,N_1659,N_1003);
or U4199 (N_4199,N_1946,N_1244);
and U4200 (N_4200,N_1464,N_1338);
nand U4201 (N_4201,N_2451,N_1261);
or U4202 (N_4202,N_381,N_1781);
or U4203 (N_4203,N_1014,N_1430);
and U4204 (N_4204,N_1605,N_56);
or U4205 (N_4205,N_2126,N_2351);
and U4206 (N_4206,N_1492,N_2150);
nand U4207 (N_4207,N_2303,N_712);
nand U4208 (N_4208,N_2461,N_2018);
nor U4209 (N_4209,N_2175,N_1965);
and U4210 (N_4210,N_2287,N_2340);
nor U4211 (N_4211,N_2344,N_1222);
and U4212 (N_4212,N_736,N_742);
nand U4213 (N_4213,N_159,N_898);
nand U4214 (N_4214,N_1284,N_1852);
nand U4215 (N_4215,N_2384,N_1758);
and U4216 (N_4216,N_1054,N_109);
nor U4217 (N_4217,N_1889,N_1668);
or U4218 (N_4218,N_1958,N_1523);
and U4219 (N_4219,N_1980,N_2077);
nor U4220 (N_4220,N_307,N_1679);
nand U4221 (N_4221,N_741,N_1737);
nor U4222 (N_4222,N_1277,N_212);
or U4223 (N_4223,N_1624,N_461);
or U4224 (N_4224,N_296,N_1085);
nor U4225 (N_4225,N_79,N_285);
or U4226 (N_4226,N_194,N_1779);
or U4227 (N_4227,N_1572,N_11);
and U4228 (N_4228,N_845,N_1637);
nor U4229 (N_4229,N_1193,N_1000);
nor U4230 (N_4230,N_2486,N_545);
or U4231 (N_4231,N_167,N_1171);
nor U4232 (N_4232,N_774,N_1223);
nor U4233 (N_4233,N_618,N_1320);
nand U4234 (N_4234,N_364,N_846);
and U4235 (N_4235,N_250,N_1616);
nor U4236 (N_4236,N_1167,N_191);
nand U4237 (N_4237,N_2081,N_2309);
nand U4238 (N_4238,N_263,N_951);
nand U4239 (N_4239,N_1386,N_470);
and U4240 (N_4240,N_113,N_1828);
or U4241 (N_4241,N_1810,N_2364);
nor U4242 (N_4242,N_1779,N_167);
or U4243 (N_4243,N_2275,N_307);
nor U4244 (N_4244,N_854,N_94);
nand U4245 (N_4245,N_2456,N_1380);
nor U4246 (N_4246,N_1331,N_421);
and U4247 (N_4247,N_1837,N_305);
nand U4248 (N_4248,N_419,N_1120);
nand U4249 (N_4249,N_650,N_2366);
nor U4250 (N_4250,N_976,N_429);
xnor U4251 (N_4251,N_1796,N_55);
nor U4252 (N_4252,N_1724,N_1888);
nand U4253 (N_4253,N_323,N_1698);
nor U4254 (N_4254,N_1815,N_2492);
and U4255 (N_4255,N_2236,N_927);
nor U4256 (N_4256,N_1847,N_1595);
nand U4257 (N_4257,N_178,N_674);
and U4258 (N_4258,N_278,N_1207);
or U4259 (N_4259,N_1953,N_181);
or U4260 (N_4260,N_1033,N_1832);
nor U4261 (N_4261,N_106,N_214);
nand U4262 (N_4262,N_2231,N_973);
and U4263 (N_4263,N_2388,N_1069);
or U4264 (N_4264,N_2033,N_1997);
nand U4265 (N_4265,N_549,N_1501);
nor U4266 (N_4266,N_690,N_315);
nand U4267 (N_4267,N_949,N_2144);
or U4268 (N_4268,N_315,N_999);
and U4269 (N_4269,N_2141,N_65);
and U4270 (N_4270,N_174,N_2070);
xnor U4271 (N_4271,N_2471,N_362);
and U4272 (N_4272,N_2417,N_1115);
and U4273 (N_4273,N_1342,N_749);
or U4274 (N_4274,N_115,N_2458);
or U4275 (N_4275,N_1629,N_1232);
and U4276 (N_4276,N_1970,N_563);
nand U4277 (N_4277,N_37,N_1575);
nor U4278 (N_4278,N_1248,N_848);
nand U4279 (N_4279,N_481,N_650);
and U4280 (N_4280,N_1841,N_1118);
and U4281 (N_4281,N_2016,N_967);
or U4282 (N_4282,N_2490,N_2220);
nor U4283 (N_4283,N_1728,N_2316);
xnor U4284 (N_4284,N_949,N_2086);
and U4285 (N_4285,N_1008,N_238);
and U4286 (N_4286,N_1153,N_1085);
nand U4287 (N_4287,N_1342,N_455);
and U4288 (N_4288,N_1639,N_1573);
and U4289 (N_4289,N_719,N_1662);
nor U4290 (N_4290,N_1336,N_1944);
or U4291 (N_4291,N_805,N_1529);
and U4292 (N_4292,N_28,N_2130);
nor U4293 (N_4293,N_2228,N_862);
or U4294 (N_4294,N_787,N_1965);
and U4295 (N_4295,N_872,N_2447);
and U4296 (N_4296,N_2011,N_2202);
and U4297 (N_4297,N_1533,N_1236);
xnor U4298 (N_4298,N_1327,N_1370);
and U4299 (N_4299,N_1422,N_1240);
or U4300 (N_4300,N_1418,N_1562);
nor U4301 (N_4301,N_1737,N_1574);
nand U4302 (N_4302,N_1530,N_31);
nand U4303 (N_4303,N_2464,N_3);
nand U4304 (N_4304,N_966,N_1890);
or U4305 (N_4305,N_2148,N_767);
nor U4306 (N_4306,N_99,N_401);
or U4307 (N_4307,N_369,N_772);
xor U4308 (N_4308,N_2245,N_86);
nor U4309 (N_4309,N_2312,N_1215);
and U4310 (N_4310,N_1011,N_568);
or U4311 (N_4311,N_733,N_1002);
and U4312 (N_4312,N_1700,N_1703);
or U4313 (N_4313,N_1107,N_754);
nand U4314 (N_4314,N_1236,N_1292);
nor U4315 (N_4315,N_108,N_614);
and U4316 (N_4316,N_1392,N_1428);
nor U4317 (N_4317,N_1534,N_1003);
and U4318 (N_4318,N_168,N_417);
nor U4319 (N_4319,N_2451,N_1529);
and U4320 (N_4320,N_28,N_231);
nor U4321 (N_4321,N_1118,N_2057);
and U4322 (N_4322,N_1084,N_416);
or U4323 (N_4323,N_264,N_962);
and U4324 (N_4324,N_715,N_1491);
or U4325 (N_4325,N_2394,N_2380);
and U4326 (N_4326,N_902,N_2156);
or U4327 (N_4327,N_2441,N_1730);
or U4328 (N_4328,N_242,N_1553);
and U4329 (N_4329,N_326,N_976);
nor U4330 (N_4330,N_212,N_556);
nor U4331 (N_4331,N_310,N_68);
nor U4332 (N_4332,N_1523,N_2366);
nand U4333 (N_4333,N_2094,N_2460);
nand U4334 (N_4334,N_394,N_1439);
or U4335 (N_4335,N_2121,N_1841);
nor U4336 (N_4336,N_1758,N_1311);
nor U4337 (N_4337,N_175,N_2340);
nand U4338 (N_4338,N_2,N_1175);
nand U4339 (N_4339,N_1485,N_859);
or U4340 (N_4340,N_134,N_640);
nor U4341 (N_4341,N_1132,N_2293);
nor U4342 (N_4342,N_985,N_2087);
and U4343 (N_4343,N_1100,N_175);
nor U4344 (N_4344,N_101,N_914);
nand U4345 (N_4345,N_204,N_522);
xnor U4346 (N_4346,N_1474,N_157);
and U4347 (N_4347,N_662,N_1539);
nor U4348 (N_4348,N_1531,N_2221);
nand U4349 (N_4349,N_1840,N_1248);
nand U4350 (N_4350,N_1298,N_2400);
nor U4351 (N_4351,N_2119,N_396);
nor U4352 (N_4352,N_576,N_1896);
nor U4353 (N_4353,N_2186,N_1269);
or U4354 (N_4354,N_2094,N_724);
and U4355 (N_4355,N_812,N_2456);
or U4356 (N_4356,N_2189,N_410);
or U4357 (N_4357,N_839,N_903);
and U4358 (N_4358,N_2131,N_1911);
nor U4359 (N_4359,N_45,N_478);
or U4360 (N_4360,N_595,N_1729);
nand U4361 (N_4361,N_571,N_232);
or U4362 (N_4362,N_881,N_2118);
or U4363 (N_4363,N_669,N_1059);
nand U4364 (N_4364,N_1219,N_695);
or U4365 (N_4365,N_1466,N_1934);
or U4366 (N_4366,N_1240,N_2391);
or U4367 (N_4367,N_1089,N_1312);
nand U4368 (N_4368,N_1089,N_2126);
nor U4369 (N_4369,N_1716,N_870);
or U4370 (N_4370,N_710,N_1024);
nand U4371 (N_4371,N_558,N_2362);
nand U4372 (N_4372,N_647,N_1046);
and U4373 (N_4373,N_466,N_2269);
nand U4374 (N_4374,N_1266,N_293);
nor U4375 (N_4375,N_2156,N_1197);
nor U4376 (N_4376,N_1831,N_835);
or U4377 (N_4377,N_1355,N_2119);
nand U4378 (N_4378,N_715,N_2251);
nor U4379 (N_4379,N_910,N_2132);
and U4380 (N_4380,N_2253,N_2441);
nor U4381 (N_4381,N_2378,N_2359);
or U4382 (N_4382,N_2363,N_1897);
and U4383 (N_4383,N_1587,N_1321);
and U4384 (N_4384,N_110,N_635);
nand U4385 (N_4385,N_2386,N_1607);
and U4386 (N_4386,N_1248,N_21);
nor U4387 (N_4387,N_804,N_284);
nor U4388 (N_4388,N_1075,N_273);
nor U4389 (N_4389,N_182,N_1272);
nor U4390 (N_4390,N_447,N_2254);
and U4391 (N_4391,N_339,N_2131);
nand U4392 (N_4392,N_729,N_1349);
and U4393 (N_4393,N_1827,N_124);
nor U4394 (N_4394,N_1450,N_525);
and U4395 (N_4395,N_1247,N_118);
or U4396 (N_4396,N_971,N_2045);
nor U4397 (N_4397,N_559,N_1024);
nand U4398 (N_4398,N_2016,N_856);
nor U4399 (N_4399,N_214,N_1282);
and U4400 (N_4400,N_98,N_1777);
and U4401 (N_4401,N_692,N_1902);
or U4402 (N_4402,N_59,N_1068);
and U4403 (N_4403,N_1329,N_1664);
and U4404 (N_4404,N_721,N_1631);
nor U4405 (N_4405,N_469,N_145);
nor U4406 (N_4406,N_1509,N_795);
nor U4407 (N_4407,N_1644,N_619);
or U4408 (N_4408,N_795,N_578);
and U4409 (N_4409,N_2207,N_147);
and U4410 (N_4410,N_2056,N_1684);
and U4411 (N_4411,N_2372,N_1218);
nand U4412 (N_4412,N_1466,N_1605);
nand U4413 (N_4413,N_419,N_2048);
nand U4414 (N_4414,N_2012,N_1408);
and U4415 (N_4415,N_2036,N_1819);
nor U4416 (N_4416,N_1368,N_2385);
or U4417 (N_4417,N_1198,N_1756);
and U4418 (N_4418,N_1075,N_1932);
or U4419 (N_4419,N_1899,N_847);
nand U4420 (N_4420,N_1069,N_538);
and U4421 (N_4421,N_2157,N_2164);
and U4422 (N_4422,N_2158,N_470);
or U4423 (N_4423,N_2465,N_597);
and U4424 (N_4424,N_2471,N_2077);
nand U4425 (N_4425,N_754,N_1259);
nand U4426 (N_4426,N_111,N_1149);
nor U4427 (N_4427,N_394,N_2107);
nand U4428 (N_4428,N_932,N_984);
or U4429 (N_4429,N_1594,N_744);
or U4430 (N_4430,N_1888,N_2060);
nand U4431 (N_4431,N_523,N_708);
and U4432 (N_4432,N_2042,N_588);
nand U4433 (N_4433,N_474,N_246);
and U4434 (N_4434,N_1374,N_2290);
nand U4435 (N_4435,N_2021,N_2287);
nand U4436 (N_4436,N_179,N_527);
nor U4437 (N_4437,N_1873,N_970);
nand U4438 (N_4438,N_1155,N_2040);
or U4439 (N_4439,N_1700,N_2435);
nand U4440 (N_4440,N_2142,N_341);
or U4441 (N_4441,N_2066,N_994);
or U4442 (N_4442,N_35,N_163);
or U4443 (N_4443,N_134,N_160);
nor U4444 (N_4444,N_2255,N_265);
or U4445 (N_4445,N_1571,N_75);
and U4446 (N_4446,N_1251,N_674);
nand U4447 (N_4447,N_1002,N_368);
nand U4448 (N_4448,N_1551,N_1711);
nor U4449 (N_4449,N_2239,N_1800);
or U4450 (N_4450,N_1781,N_491);
or U4451 (N_4451,N_2065,N_234);
and U4452 (N_4452,N_1994,N_2207);
nand U4453 (N_4453,N_2135,N_2167);
and U4454 (N_4454,N_1832,N_681);
and U4455 (N_4455,N_1962,N_1384);
and U4456 (N_4456,N_219,N_2295);
or U4457 (N_4457,N_544,N_1377);
and U4458 (N_4458,N_501,N_2324);
or U4459 (N_4459,N_2027,N_1530);
or U4460 (N_4460,N_990,N_1021);
nand U4461 (N_4461,N_1172,N_2019);
and U4462 (N_4462,N_1162,N_1048);
nand U4463 (N_4463,N_1935,N_171);
and U4464 (N_4464,N_75,N_2227);
nor U4465 (N_4465,N_307,N_1335);
nor U4466 (N_4466,N_768,N_650);
nor U4467 (N_4467,N_251,N_1824);
nand U4468 (N_4468,N_1387,N_155);
or U4469 (N_4469,N_1477,N_1450);
or U4470 (N_4470,N_1552,N_1649);
or U4471 (N_4471,N_2192,N_298);
nor U4472 (N_4472,N_1783,N_2370);
and U4473 (N_4473,N_1158,N_1140);
and U4474 (N_4474,N_112,N_593);
nor U4475 (N_4475,N_274,N_389);
nor U4476 (N_4476,N_231,N_1667);
or U4477 (N_4477,N_1443,N_2136);
or U4478 (N_4478,N_73,N_1718);
or U4479 (N_4479,N_990,N_370);
or U4480 (N_4480,N_699,N_115);
nor U4481 (N_4481,N_426,N_2106);
or U4482 (N_4482,N_1116,N_388);
nor U4483 (N_4483,N_674,N_1945);
nand U4484 (N_4484,N_292,N_2206);
and U4485 (N_4485,N_1673,N_2448);
nand U4486 (N_4486,N_2029,N_1045);
nand U4487 (N_4487,N_2473,N_212);
nor U4488 (N_4488,N_429,N_1692);
nor U4489 (N_4489,N_1786,N_1678);
and U4490 (N_4490,N_221,N_324);
and U4491 (N_4491,N_876,N_1524);
nand U4492 (N_4492,N_997,N_80);
nand U4493 (N_4493,N_1097,N_2357);
or U4494 (N_4494,N_127,N_1645);
or U4495 (N_4495,N_1672,N_2436);
or U4496 (N_4496,N_1283,N_1447);
and U4497 (N_4497,N_968,N_197);
and U4498 (N_4498,N_594,N_877);
nand U4499 (N_4499,N_1861,N_1167);
nor U4500 (N_4500,N_2210,N_21);
and U4501 (N_4501,N_876,N_925);
or U4502 (N_4502,N_880,N_899);
xnor U4503 (N_4503,N_331,N_1086);
or U4504 (N_4504,N_370,N_2489);
nor U4505 (N_4505,N_130,N_2034);
and U4506 (N_4506,N_2430,N_1187);
nand U4507 (N_4507,N_1403,N_172);
nand U4508 (N_4508,N_83,N_2068);
nand U4509 (N_4509,N_1303,N_1429);
nor U4510 (N_4510,N_689,N_1543);
or U4511 (N_4511,N_544,N_1894);
or U4512 (N_4512,N_1984,N_2188);
nor U4513 (N_4513,N_306,N_63);
or U4514 (N_4514,N_1245,N_279);
nand U4515 (N_4515,N_1212,N_1089);
nor U4516 (N_4516,N_2352,N_2440);
and U4517 (N_4517,N_784,N_2468);
nor U4518 (N_4518,N_1343,N_2441);
nand U4519 (N_4519,N_789,N_2131);
nand U4520 (N_4520,N_1494,N_1042);
and U4521 (N_4521,N_117,N_2095);
nand U4522 (N_4522,N_2233,N_1291);
nand U4523 (N_4523,N_2372,N_627);
or U4524 (N_4524,N_1418,N_952);
and U4525 (N_4525,N_1413,N_1891);
or U4526 (N_4526,N_339,N_2182);
and U4527 (N_4527,N_2442,N_1111);
nand U4528 (N_4528,N_1120,N_238);
nor U4529 (N_4529,N_1699,N_2291);
or U4530 (N_4530,N_1834,N_822);
or U4531 (N_4531,N_1080,N_1500);
xor U4532 (N_4532,N_447,N_2377);
and U4533 (N_4533,N_70,N_1048);
or U4534 (N_4534,N_1511,N_1051);
and U4535 (N_4535,N_1116,N_2291);
nand U4536 (N_4536,N_564,N_1376);
nand U4537 (N_4537,N_312,N_2458);
nand U4538 (N_4538,N_188,N_1187);
nor U4539 (N_4539,N_2398,N_269);
or U4540 (N_4540,N_504,N_1304);
nand U4541 (N_4541,N_589,N_44);
nor U4542 (N_4542,N_872,N_306);
nor U4543 (N_4543,N_955,N_1704);
and U4544 (N_4544,N_1298,N_1860);
nand U4545 (N_4545,N_220,N_115);
and U4546 (N_4546,N_1078,N_2072);
or U4547 (N_4547,N_1654,N_2019);
and U4548 (N_4548,N_1241,N_1899);
and U4549 (N_4549,N_149,N_21);
nor U4550 (N_4550,N_325,N_597);
nand U4551 (N_4551,N_400,N_2261);
nor U4552 (N_4552,N_1426,N_2100);
and U4553 (N_4553,N_385,N_2424);
nand U4554 (N_4554,N_1010,N_1967);
nor U4555 (N_4555,N_123,N_640);
and U4556 (N_4556,N_1897,N_1782);
or U4557 (N_4557,N_661,N_1392);
or U4558 (N_4558,N_1940,N_1968);
or U4559 (N_4559,N_2258,N_53);
nor U4560 (N_4560,N_283,N_553);
nand U4561 (N_4561,N_2370,N_1959);
nand U4562 (N_4562,N_714,N_111);
nand U4563 (N_4563,N_1749,N_2453);
nor U4564 (N_4564,N_1971,N_1400);
or U4565 (N_4565,N_1678,N_2357);
nand U4566 (N_4566,N_1494,N_2455);
and U4567 (N_4567,N_2218,N_1190);
nor U4568 (N_4568,N_339,N_551);
nand U4569 (N_4569,N_1629,N_904);
nand U4570 (N_4570,N_1064,N_2030);
nor U4571 (N_4571,N_2349,N_555);
and U4572 (N_4572,N_6,N_1031);
or U4573 (N_4573,N_1673,N_1993);
nand U4574 (N_4574,N_509,N_2322);
nand U4575 (N_4575,N_1142,N_2393);
and U4576 (N_4576,N_846,N_999);
nor U4577 (N_4577,N_719,N_97);
or U4578 (N_4578,N_2382,N_1870);
and U4579 (N_4579,N_696,N_1378);
and U4580 (N_4580,N_984,N_107);
nor U4581 (N_4581,N_1159,N_2228);
nand U4582 (N_4582,N_2059,N_1939);
nor U4583 (N_4583,N_1737,N_762);
nand U4584 (N_4584,N_2372,N_246);
nor U4585 (N_4585,N_212,N_2332);
and U4586 (N_4586,N_1277,N_2112);
nand U4587 (N_4587,N_712,N_2410);
or U4588 (N_4588,N_1466,N_1968);
nor U4589 (N_4589,N_1259,N_1738);
and U4590 (N_4590,N_611,N_104);
or U4591 (N_4591,N_1958,N_2269);
and U4592 (N_4592,N_2064,N_1076);
nand U4593 (N_4593,N_667,N_2012);
nor U4594 (N_4594,N_613,N_2354);
or U4595 (N_4595,N_862,N_1587);
or U4596 (N_4596,N_1502,N_2403);
and U4597 (N_4597,N_1003,N_2053);
nor U4598 (N_4598,N_895,N_1599);
or U4599 (N_4599,N_2483,N_1395);
or U4600 (N_4600,N_1320,N_1420);
nor U4601 (N_4601,N_1984,N_1505);
nand U4602 (N_4602,N_930,N_2221);
or U4603 (N_4603,N_181,N_1484);
nor U4604 (N_4604,N_1511,N_851);
nor U4605 (N_4605,N_1784,N_1219);
nand U4606 (N_4606,N_1040,N_853);
or U4607 (N_4607,N_1078,N_2362);
or U4608 (N_4608,N_1950,N_942);
or U4609 (N_4609,N_1356,N_1202);
nor U4610 (N_4610,N_1759,N_700);
nor U4611 (N_4611,N_111,N_1206);
nand U4612 (N_4612,N_2095,N_458);
nand U4613 (N_4613,N_1384,N_655);
nand U4614 (N_4614,N_1208,N_2120);
and U4615 (N_4615,N_215,N_1426);
nor U4616 (N_4616,N_1485,N_61);
or U4617 (N_4617,N_1234,N_878);
and U4618 (N_4618,N_1290,N_2148);
or U4619 (N_4619,N_1053,N_351);
and U4620 (N_4620,N_1220,N_1921);
or U4621 (N_4621,N_99,N_2192);
xor U4622 (N_4622,N_743,N_755);
nor U4623 (N_4623,N_1711,N_1200);
nand U4624 (N_4624,N_1559,N_1193);
and U4625 (N_4625,N_2273,N_10);
or U4626 (N_4626,N_2254,N_1910);
nand U4627 (N_4627,N_2390,N_165);
nor U4628 (N_4628,N_1392,N_528);
nand U4629 (N_4629,N_2358,N_910);
and U4630 (N_4630,N_2420,N_1825);
or U4631 (N_4631,N_2129,N_1909);
nand U4632 (N_4632,N_1034,N_1814);
nor U4633 (N_4633,N_585,N_2189);
nor U4634 (N_4634,N_869,N_1947);
nand U4635 (N_4635,N_512,N_1291);
nor U4636 (N_4636,N_275,N_1196);
nor U4637 (N_4637,N_1270,N_2346);
nor U4638 (N_4638,N_138,N_835);
nor U4639 (N_4639,N_1773,N_518);
or U4640 (N_4640,N_2448,N_707);
and U4641 (N_4641,N_200,N_1188);
and U4642 (N_4642,N_1009,N_903);
nor U4643 (N_4643,N_1170,N_2126);
and U4644 (N_4644,N_1089,N_1971);
or U4645 (N_4645,N_2258,N_1439);
nand U4646 (N_4646,N_1361,N_1898);
and U4647 (N_4647,N_99,N_372);
nor U4648 (N_4648,N_369,N_1937);
nand U4649 (N_4649,N_1399,N_1303);
or U4650 (N_4650,N_1648,N_768);
nor U4651 (N_4651,N_1980,N_1116);
nor U4652 (N_4652,N_2169,N_2260);
nand U4653 (N_4653,N_968,N_1688);
nor U4654 (N_4654,N_278,N_1600);
or U4655 (N_4655,N_1321,N_712);
nor U4656 (N_4656,N_1261,N_593);
and U4657 (N_4657,N_1418,N_458);
and U4658 (N_4658,N_2171,N_2256);
nand U4659 (N_4659,N_464,N_416);
nand U4660 (N_4660,N_1936,N_1422);
or U4661 (N_4661,N_1869,N_526);
or U4662 (N_4662,N_1153,N_2350);
nor U4663 (N_4663,N_1428,N_1659);
nor U4664 (N_4664,N_1944,N_1338);
or U4665 (N_4665,N_580,N_1235);
or U4666 (N_4666,N_629,N_60);
and U4667 (N_4667,N_1631,N_2353);
nor U4668 (N_4668,N_653,N_2180);
nor U4669 (N_4669,N_1321,N_740);
or U4670 (N_4670,N_2075,N_736);
nor U4671 (N_4671,N_461,N_1485);
and U4672 (N_4672,N_1951,N_1302);
nor U4673 (N_4673,N_298,N_1495);
or U4674 (N_4674,N_865,N_1611);
or U4675 (N_4675,N_742,N_1805);
and U4676 (N_4676,N_899,N_2440);
or U4677 (N_4677,N_767,N_353);
and U4678 (N_4678,N_417,N_2092);
and U4679 (N_4679,N_1476,N_1468);
nor U4680 (N_4680,N_2312,N_2354);
and U4681 (N_4681,N_2115,N_2218);
nand U4682 (N_4682,N_1240,N_2041);
nor U4683 (N_4683,N_1769,N_255);
nand U4684 (N_4684,N_1796,N_1280);
or U4685 (N_4685,N_983,N_1697);
and U4686 (N_4686,N_1148,N_1621);
nor U4687 (N_4687,N_2262,N_2323);
or U4688 (N_4688,N_81,N_1898);
nand U4689 (N_4689,N_232,N_566);
nand U4690 (N_4690,N_1540,N_942);
nor U4691 (N_4691,N_1127,N_1793);
nand U4692 (N_4692,N_422,N_199);
nor U4693 (N_4693,N_1044,N_1335);
nand U4694 (N_4694,N_258,N_1981);
or U4695 (N_4695,N_627,N_574);
or U4696 (N_4696,N_1340,N_1335);
or U4697 (N_4697,N_235,N_1560);
nand U4698 (N_4698,N_872,N_1637);
nor U4699 (N_4699,N_69,N_9);
or U4700 (N_4700,N_353,N_335);
or U4701 (N_4701,N_2091,N_1087);
or U4702 (N_4702,N_2408,N_681);
or U4703 (N_4703,N_1987,N_1583);
nand U4704 (N_4704,N_62,N_1449);
or U4705 (N_4705,N_651,N_1229);
nor U4706 (N_4706,N_1711,N_2144);
nor U4707 (N_4707,N_402,N_11);
or U4708 (N_4708,N_907,N_1417);
nand U4709 (N_4709,N_2283,N_1755);
nor U4710 (N_4710,N_1986,N_2084);
and U4711 (N_4711,N_782,N_2036);
or U4712 (N_4712,N_782,N_686);
nand U4713 (N_4713,N_562,N_2457);
or U4714 (N_4714,N_1576,N_1905);
nand U4715 (N_4715,N_1734,N_1224);
nand U4716 (N_4716,N_370,N_335);
or U4717 (N_4717,N_2470,N_1463);
and U4718 (N_4718,N_919,N_2164);
nor U4719 (N_4719,N_1328,N_399);
and U4720 (N_4720,N_173,N_478);
xnor U4721 (N_4721,N_130,N_572);
nor U4722 (N_4722,N_357,N_43);
nor U4723 (N_4723,N_1831,N_2495);
nor U4724 (N_4724,N_1582,N_241);
and U4725 (N_4725,N_1409,N_120);
and U4726 (N_4726,N_1638,N_1958);
nand U4727 (N_4727,N_994,N_1081);
nand U4728 (N_4728,N_1404,N_60);
nor U4729 (N_4729,N_406,N_542);
and U4730 (N_4730,N_1428,N_605);
nor U4731 (N_4731,N_332,N_1032);
nand U4732 (N_4732,N_1399,N_560);
nor U4733 (N_4733,N_290,N_1462);
xnor U4734 (N_4734,N_242,N_2047);
nand U4735 (N_4735,N_628,N_2245);
nand U4736 (N_4736,N_2003,N_360);
nand U4737 (N_4737,N_780,N_1782);
xor U4738 (N_4738,N_1530,N_2196);
nor U4739 (N_4739,N_1322,N_1239);
and U4740 (N_4740,N_1505,N_1212);
or U4741 (N_4741,N_1148,N_1131);
nor U4742 (N_4742,N_629,N_660);
xnor U4743 (N_4743,N_979,N_1652);
nor U4744 (N_4744,N_1793,N_499);
and U4745 (N_4745,N_1198,N_627);
and U4746 (N_4746,N_362,N_1142);
and U4747 (N_4747,N_781,N_155);
or U4748 (N_4748,N_1826,N_2202);
and U4749 (N_4749,N_1274,N_2488);
and U4750 (N_4750,N_1955,N_199);
nor U4751 (N_4751,N_301,N_1613);
nor U4752 (N_4752,N_284,N_2414);
and U4753 (N_4753,N_608,N_593);
and U4754 (N_4754,N_1625,N_957);
or U4755 (N_4755,N_84,N_511);
nor U4756 (N_4756,N_641,N_1278);
or U4757 (N_4757,N_594,N_1960);
nand U4758 (N_4758,N_60,N_713);
nor U4759 (N_4759,N_1098,N_2420);
nand U4760 (N_4760,N_1942,N_1351);
and U4761 (N_4761,N_328,N_87);
and U4762 (N_4762,N_894,N_1449);
nand U4763 (N_4763,N_552,N_1526);
or U4764 (N_4764,N_969,N_2264);
or U4765 (N_4765,N_1093,N_1948);
or U4766 (N_4766,N_1064,N_1967);
and U4767 (N_4767,N_13,N_465);
nor U4768 (N_4768,N_1332,N_523);
nand U4769 (N_4769,N_1109,N_758);
nor U4770 (N_4770,N_471,N_1299);
and U4771 (N_4771,N_1876,N_21);
and U4772 (N_4772,N_2349,N_1028);
or U4773 (N_4773,N_502,N_884);
and U4774 (N_4774,N_204,N_39);
nor U4775 (N_4775,N_2128,N_2475);
or U4776 (N_4776,N_2221,N_1270);
or U4777 (N_4777,N_1079,N_1501);
nor U4778 (N_4778,N_1981,N_1689);
nand U4779 (N_4779,N_1919,N_1394);
nor U4780 (N_4780,N_241,N_2025);
and U4781 (N_4781,N_2351,N_168);
nand U4782 (N_4782,N_1253,N_1869);
or U4783 (N_4783,N_2057,N_873);
nand U4784 (N_4784,N_2482,N_1596);
or U4785 (N_4785,N_1458,N_691);
nor U4786 (N_4786,N_30,N_627);
and U4787 (N_4787,N_1,N_1164);
and U4788 (N_4788,N_1811,N_2320);
nor U4789 (N_4789,N_2264,N_1735);
or U4790 (N_4790,N_862,N_1420);
nor U4791 (N_4791,N_118,N_1894);
or U4792 (N_4792,N_472,N_1424);
nor U4793 (N_4793,N_264,N_1237);
and U4794 (N_4794,N_1474,N_1400);
and U4795 (N_4795,N_553,N_1297);
or U4796 (N_4796,N_451,N_1300);
nand U4797 (N_4797,N_2179,N_368);
nand U4798 (N_4798,N_18,N_2169);
and U4799 (N_4799,N_265,N_1321);
nand U4800 (N_4800,N_909,N_1466);
nand U4801 (N_4801,N_2485,N_1643);
and U4802 (N_4802,N_1488,N_548);
and U4803 (N_4803,N_2228,N_31);
nand U4804 (N_4804,N_1309,N_1502);
or U4805 (N_4805,N_356,N_686);
nor U4806 (N_4806,N_704,N_1289);
and U4807 (N_4807,N_613,N_2139);
nor U4808 (N_4808,N_136,N_960);
nand U4809 (N_4809,N_985,N_596);
nor U4810 (N_4810,N_1515,N_299);
or U4811 (N_4811,N_998,N_2469);
nor U4812 (N_4812,N_2300,N_5);
and U4813 (N_4813,N_1116,N_250);
and U4814 (N_4814,N_987,N_2406);
or U4815 (N_4815,N_1351,N_2182);
nor U4816 (N_4816,N_648,N_2319);
nor U4817 (N_4817,N_859,N_830);
and U4818 (N_4818,N_2446,N_1394);
nor U4819 (N_4819,N_1375,N_2063);
nor U4820 (N_4820,N_584,N_2377);
and U4821 (N_4821,N_283,N_638);
nor U4822 (N_4822,N_1112,N_647);
nor U4823 (N_4823,N_2137,N_2055);
nand U4824 (N_4824,N_977,N_2123);
and U4825 (N_4825,N_2304,N_436);
nand U4826 (N_4826,N_414,N_1051);
or U4827 (N_4827,N_408,N_2460);
or U4828 (N_4828,N_1594,N_119);
nand U4829 (N_4829,N_1321,N_1811);
or U4830 (N_4830,N_577,N_2291);
nor U4831 (N_4831,N_23,N_1532);
and U4832 (N_4832,N_1291,N_876);
nand U4833 (N_4833,N_584,N_1854);
and U4834 (N_4834,N_340,N_661);
nand U4835 (N_4835,N_2221,N_556);
xnor U4836 (N_4836,N_1099,N_2018);
and U4837 (N_4837,N_1999,N_434);
nand U4838 (N_4838,N_1385,N_1471);
and U4839 (N_4839,N_878,N_2150);
xor U4840 (N_4840,N_336,N_177);
and U4841 (N_4841,N_2245,N_2492);
or U4842 (N_4842,N_1531,N_780);
and U4843 (N_4843,N_1457,N_2464);
or U4844 (N_4844,N_1240,N_1740);
nand U4845 (N_4845,N_448,N_1504);
nor U4846 (N_4846,N_1623,N_819);
nor U4847 (N_4847,N_471,N_185);
and U4848 (N_4848,N_154,N_939);
and U4849 (N_4849,N_1645,N_683);
nand U4850 (N_4850,N_2003,N_68);
or U4851 (N_4851,N_2389,N_50);
nand U4852 (N_4852,N_2026,N_964);
nand U4853 (N_4853,N_664,N_1325);
nor U4854 (N_4854,N_1206,N_705);
nand U4855 (N_4855,N_859,N_1591);
nand U4856 (N_4856,N_2495,N_1318);
nor U4857 (N_4857,N_1740,N_356);
and U4858 (N_4858,N_2158,N_2082);
or U4859 (N_4859,N_929,N_736);
and U4860 (N_4860,N_2113,N_1100);
nand U4861 (N_4861,N_1554,N_1689);
nor U4862 (N_4862,N_2442,N_2226);
nand U4863 (N_4863,N_1276,N_2228);
nor U4864 (N_4864,N_9,N_1997);
nor U4865 (N_4865,N_1244,N_1293);
nand U4866 (N_4866,N_226,N_2470);
nor U4867 (N_4867,N_1629,N_2034);
xor U4868 (N_4868,N_286,N_603);
and U4869 (N_4869,N_623,N_427);
or U4870 (N_4870,N_1179,N_381);
nor U4871 (N_4871,N_1892,N_1435);
nand U4872 (N_4872,N_78,N_2414);
xor U4873 (N_4873,N_1266,N_1629);
and U4874 (N_4874,N_443,N_499);
nand U4875 (N_4875,N_1482,N_315);
nor U4876 (N_4876,N_1023,N_1228);
and U4877 (N_4877,N_589,N_1798);
or U4878 (N_4878,N_1153,N_689);
nand U4879 (N_4879,N_835,N_2162);
nor U4880 (N_4880,N_729,N_334);
nand U4881 (N_4881,N_2427,N_602);
and U4882 (N_4882,N_2103,N_1763);
and U4883 (N_4883,N_489,N_1664);
nand U4884 (N_4884,N_1647,N_1259);
nand U4885 (N_4885,N_8,N_1569);
nand U4886 (N_4886,N_207,N_458);
nor U4887 (N_4887,N_140,N_748);
nor U4888 (N_4888,N_1685,N_2218);
and U4889 (N_4889,N_2089,N_2085);
and U4890 (N_4890,N_771,N_1913);
and U4891 (N_4891,N_1069,N_1442);
nand U4892 (N_4892,N_1165,N_1559);
nand U4893 (N_4893,N_1797,N_730);
and U4894 (N_4894,N_452,N_2104);
or U4895 (N_4895,N_29,N_794);
and U4896 (N_4896,N_478,N_1647);
nand U4897 (N_4897,N_485,N_1436);
nand U4898 (N_4898,N_2107,N_2344);
or U4899 (N_4899,N_2248,N_1273);
and U4900 (N_4900,N_1677,N_1579);
and U4901 (N_4901,N_2024,N_523);
or U4902 (N_4902,N_1162,N_1987);
and U4903 (N_4903,N_55,N_2094);
nor U4904 (N_4904,N_1889,N_1254);
nand U4905 (N_4905,N_358,N_1408);
or U4906 (N_4906,N_904,N_1748);
nand U4907 (N_4907,N_1098,N_1947);
nand U4908 (N_4908,N_1117,N_1859);
or U4909 (N_4909,N_2205,N_212);
nand U4910 (N_4910,N_2164,N_41);
or U4911 (N_4911,N_1612,N_1165);
and U4912 (N_4912,N_1477,N_1034);
and U4913 (N_4913,N_167,N_911);
and U4914 (N_4914,N_1379,N_607);
nand U4915 (N_4915,N_1441,N_849);
or U4916 (N_4916,N_89,N_918);
nand U4917 (N_4917,N_894,N_1909);
and U4918 (N_4918,N_189,N_1683);
xnor U4919 (N_4919,N_728,N_1429);
nor U4920 (N_4920,N_1167,N_2416);
and U4921 (N_4921,N_361,N_2135);
nand U4922 (N_4922,N_338,N_493);
or U4923 (N_4923,N_1913,N_906);
nor U4924 (N_4924,N_1010,N_1095);
nor U4925 (N_4925,N_2105,N_1183);
and U4926 (N_4926,N_781,N_1445);
or U4927 (N_4927,N_1331,N_1828);
nor U4928 (N_4928,N_1081,N_248);
nor U4929 (N_4929,N_1835,N_1396);
or U4930 (N_4930,N_2362,N_2122);
or U4931 (N_4931,N_1323,N_14);
or U4932 (N_4932,N_1965,N_2222);
and U4933 (N_4933,N_2241,N_1586);
or U4934 (N_4934,N_525,N_2044);
or U4935 (N_4935,N_722,N_1025);
nor U4936 (N_4936,N_124,N_2130);
or U4937 (N_4937,N_901,N_1073);
nor U4938 (N_4938,N_541,N_944);
and U4939 (N_4939,N_455,N_1386);
or U4940 (N_4940,N_2045,N_299);
and U4941 (N_4941,N_367,N_327);
and U4942 (N_4942,N_707,N_1447);
nor U4943 (N_4943,N_1482,N_712);
nor U4944 (N_4944,N_456,N_2347);
nand U4945 (N_4945,N_619,N_1960);
nor U4946 (N_4946,N_1934,N_1882);
nor U4947 (N_4947,N_962,N_970);
nor U4948 (N_4948,N_2499,N_2385);
or U4949 (N_4949,N_147,N_1723);
and U4950 (N_4950,N_473,N_47);
nand U4951 (N_4951,N_780,N_2386);
and U4952 (N_4952,N_1125,N_345);
and U4953 (N_4953,N_285,N_1214);
nor U4954 (N_4954,N_2336,N_1091);
nor U4955 (N_4955,N_1476,N_2477);
and U4956 (N_4956,N_1523,N_1753);
nor U4957 (N_4957,N_2102,N_266);
nand U4958 (N_4958,N_2398,N_1197);
or U4959 (N_4959,N_1879,N_2219);
nor U4960 (N_4960,N_1530,N_1276);
nor U4961 (N_4961,N_892,N_1538);
nor U4962 (N_4962,N_1041,N_1537);
or U4963 (N_4963,N_2104,N_110);
xor U4964 (N_4964,N_926,N_1145);
nand U4965 (N_4965,N_905,N_185);
and U4966 (N_4966,N_2172,N_1938);
nor U4967 (N_4967,N_738,N_2244);
nor U4968 (N_4968,N_1617,N_1063);
or U4969 (N_4969,N_1353,N_77);
nand U4970 (N_4970,N_415,N_1726);
nor U4971 (N_4971,N_2188,N_2423);
nand U4972 (N_4972,N_50,N_696);
nor U4973 (N_4973,N_1970,N_993);
nand U4974 (N_4974,N_761,N_1336);
nand U4975 (N_4975,N_848,N_679);
nand U4976 (N_4976,N_1083,N_1193);
and U4977 (N_4977,N_2434,N_1511);
and U4978 (N_4978,N_2398,N_1329);
and U4979 (N_4979,N_1133,N_1012);
nand U4980 (N_4980,N_1109,N_1174);
nand U4981 (N_4981,N_470,N_2394);
nand U4982 (N_4982,N_968,N_1760);
nor U4983 (N_4983,N_237,N_2196);
or U4984 (N_4984,N_75,N_986);
nor U4985 (N_4985,N_287,N_2033);
or U4986 (N_4986,N_2393,N_2277);
or U4987 (N_4987,N_253,N_554);
nand U4988 (N_4988,N_2295,N_2321);
xnor U4989 (N_4989,N_1685,N_519);
and U4990 (N_4990,N_1511,N_799);
nand U4991 (N_4991,N_245,N_1157);
nor U4992 (N_4992,N_777,N_2398);
and U4993 (N_4993,N_2212,N_1403);
nor U4994 (N_4994,N_2277,N_340);
and U4995 (N_4995,N_624,N_721);
nor U4996 (N_4996,N_1796,N_1952);
nand U4997 (N_4997,N_2155,N_409);
and U4998 (N_4998,N_1991,N_1327);
and U4999 (N_4999,N_2001,N_1477);
and U5000 (N_5000,N_3951,N_4125);
and U5001 (N_5001,N_3713,N_3282);
nand U5002 (N_5002,N_2896,N_3477);
nor U5003 (N_5003,N_4470,N_3409);
and U5004 (N_5004,N_3950,N_3649);
nand U5005 (N_5005,N_4006,N_2936);
and U5006 (N_5006,N_4372,N_3820);
nand U5007 (N_5007,N_3944,N_2579);
nand U5008 (N_5008,N_4968,N_4082);
or U5009 (N_5009,N_2775,N_3485);
or U5010 (N_5010,N_2857,N_4616);
nor U5011 (N_5011,N_3965,N_4702);
and U5012 (N_5012,N_4270,N_3032);
or U5013 (N_5013,N_3515,N_4199);
nand U5014 (N_5014,N_3229,N_3019);
nand U5015 (N_5015,N_4031,N_4770);
and U5016 (N_5016,N_4340,N_4212);
nor U5017 (N_5017,N_4876,N_4570);
or U5018 (N_5018,N_2517,N_3058);
nand U5019 (N_5019,N_4257,N_4840);
and U5020 (N_5020,N_3131,N_2767);
and U5021 (N_5021,N_2625,N_3446);
and U5022 (N_5022,N_4800,N_3440);
or U5023 (N_5023,N_3768,N_3194);
and U5024 (N_5024,N_4777,N_3373);
nor U5025 (N_5025,N_4015,N_3895);
or U5026 (N_5026,N_2679,N_4453);
and U5027 (N_5027,N_4419,N_3272);
and U5028 (N_5028,N_4630,N_3645);
and U5029 (N_5029,N_3821,N_2808);
and U5030 (N_5030,N_4473,N_4053);
nand U5031 (N_5031,N_2923,N_3925);
and U5032 (N_5032,N_4640,N_3223);
and U5033 (N_5033,N_4107,N_3494);
or U5034 (N_5034,N_3694,N_4239);
nor U5035 (N_5035,N_2878,N_4818);
nand U5036 (N_5036,N_3149,N_2649);
or U5037 (N_5037,N_4292,N_4900);
nor U5038 (N_5038,N_4195,N_2774);
nor U5039 (N_5039,N_4917,N_2846);
or U5040 (N_5040,N_4138,N_4303);
nand U5041 (N_5041,N_4454,N_2590);
and U5042 (N_5042,N_4606,N_2897);
nand U5043 (N_5043,N_3604,N_2550);
and U5044 (N_5044,N_4209,N_4124);
or U5045 (N_5045,N_2950,N_3263);
nor U5046 (N_5046,N_3743,N_4431);
nor U5047 (N_5047,N_2593,N_4515);
nor U5048 (N_5048,N_4830,N_4423);
nor U5049 (N_5049,N_4821,N_4106);
nand U5050 (N_5050,N_3523,N_4699);
and U5051 (N_5051,N_4156,N_3901);
nand U5052 (N_5052,N_3598,N_3383);
nor U5053 (N_5053,N_4399,N_4507);
nor U5054 (N_5054,N_3259,N_2752);
or U5055 (N_5055,N_3453,N_3359);
nor U5056 (N_5056,N_3000,N_4673);
and U5057 (N_5057,N_3558,N_4398);
or U5058 (N_5058,N_2570,N_3309);
and U5059 (N_5059,N_3844,N_3335);
nand U5060 (N_5060,N_2829,N_4761);
nand U5061 (N_5061,N_3854,N_3980);
or U5062 (N_5062,N_3143,N_3184);
nor U5063 (N_5063,N_2639,N_4690);
or U5064 (N_5064,N_4835,N_3336);
and U5065 (N_5065,N_3405,N_3260);
nor U5066 (N_5066,N_4854,N_3419);
xnor U5067 (N_5067,N_3812,N_4997);
or U5068 (N_5068,N_4281,N_3614);
nand U5069 (N_5069,N_3512,N_4576);
or U5070 (N_5070,N_3356,N_2680);
nand U5071 (N_5071,N_3848,N_4300);
and U5072 (N_5072,N_4058,N_4801);
nor U5073 (N_5073,N_3176,N_4963);
and U5074 (N_5074,N_3095,N_2854);
nand U5075 (N_5075,N_4809,N_3006);
nor U5076 (N_5076,N_3702,N_4946);
nor U5077 (N_5077,N_4989,N_4127);
nor U5078 (N_5078,N_4574,N_4462);
and U5079 (N_5079,N_3817,N_2841);
nand U5080 (N_5080,N_3370,N_4554);
or U5081 (N_5081,N_3119,N_3536);
nor U5082 (N_5082,N_3639,N_4725);
and U5083 (N_5083,N_2844,N_2665);
nand U5084 (N_5084,N_3305,N_2515);
nand U5085 (N_5085,N_2778,N_4126);
nor U5086 (N_5086,N_3436,N_3894);
and U5087 (N_5087,N_3150,N_4223);
nand U5088 (N_5088,N_2801,N_3246);
or U5089 (N_5089,N_4000,N_4162);
and U5090 (N_5090,N_4406,N_4157);
and U5091 (N_5091,N_4544,N_4390);
or U5092 (N_5092,N_2540,N_2969);
or U5093 (N_5093,N_4084,N_2693);
and U5094 (N_5094,N_3703,N_4421);
and U5095 (N_5095,N_2733,N_3715);
and U5096 (N_5096,N_4683,N_3550);
nor U5097 (N_5097,N_2911,N_3306);
nor U5098 (N_5098,N_2973,N_3544);
nor U5099 (N_5099,N_2553,N_4524);
nand U5100 (N_5100,N_3947,N_4135);
xor U5101 (N_5101,N_2521,N_2994);
nand U5102 (N_5102,N_4776,N_4420);
nor U5103 (N_5103,N_3746,N_2949);
nor U5104 (N_5104,N_2859,N_4693);
nand U5105 (N_5105,N_3255,N_3066);
or U5106 (N_5106,N_3672,N_4905);
nor U5107 (N_5107,N_4095,N_2974);
nor U5108 (N_5108,N_3172,N_3799);
nor U5109 (N_5109,N_4437,N_3545);
and U5110 (N_5110,N_3532,N_4150);
or U5111 (N_5111,N_4033,N_3624);
and U5112 (N_5112,N_3090,N_3287);
nand U5113 (N_5113,N_3943,N_3392);
nor U5114 (N_5114,N_2556,N_4247);
nand U5115 (N_5115,N_3843,N_2934);
nor U5116 (N_5116,N_3926,N_4101);
nand U5117 (N_5117,N_4768,N_4733);
or U5118 (N_5118,N_4996,N_3683);
nor U5119 (N_5119,N_2605,N_4594);
and U5120 (N_5120,N_4704,N_4021);
and U5121 (N_5121,N_3455,N_4207);
nand U5122 (N_5122,N_3295,N_3525);
or U5123 (N_5123,N_3687,N_4526);
or U5124 (N_5124,N_2781,N_4951);
nand U5125 (N_5125,N_3480,N_4650);
nor U5126 (N_5126,N_3736,N_4653);
and U5127 (N_5127,N_4678,N_3810);
nor U5128 (N_5128,N_4986,N_3101);
or U5129 (N_5129,N_2700,N_3004);
and U5130 (N_5130,N_3625,N_4277);
or U5131 (N_5131,N_2863,N_4228);
or U5132 (N_5132,N_4294,N_4430);
and U5133 (N_5133,N_3922,N_3721);
nand U5134 (N_5134,N_4852,N_2996);
nor U5135 (N_5135,N_4903,N_3372);
and U5136 (N_5136,N_3358,N_4141);
nand U5137 (N_5137,N_2618,N_4050);
or U5138 (N_5138,N_2601,N_2559);
nor U5139 (N_5139,N_3406,N_3399);
nand U5140 (N_5140,N_3958,N_3533);
nor U5141 (N_5141,N_2821,N_4767);
or U5142 (N_5142,N_2581,N_2770);
or U5143 (N_5143,N_3754,N_4792);
nand U5144 (N_5144,N_4395,N_3834);
nand U5145 (N_5145,N_3072,N_4932);
nand U5146 (N_5146,N_4560,N_3668);
nor U5147 (N_5147,N_3977,N_4295);
and U5148 (N_5148,N_3781,N_3479);
or U5149 (N_5149,N_4930,N_2648);
and U5150 (N_5150,N_2864,N_2732);
and U5151 (N_5151,N_4758,N_3775);
nand U5152 (N_5152,N_3278,N_2787);
nand U5153 (N_5153,N_4347,N_3915);
and U5154 (N_5154,N_4875,N_4374);
nor U5155 (N_5155,N_3568,N_4323);
and U5156 (N_5156,N_3934,N_4729);
nor U5157 (N_5157,N_2756,N_4279);
nor U5158 (N_5158,N_4692,N_3562);
nand U5159 (N_5159,N_4566,N_3851);
nor U5160 (N_5160,N_2734,N_4320);
or U5161 (N_5161,N_3232,N_3966);
or U5162 (N_5162,N_2908,N_3648);
and U5163 (N_5163,N_4788,N_4737);
and U5164 (N_5164,N_4086,N_3644);
nor U5165 (N_5165,N_4363,N_4427);
nor U5166 (N_5166,N_3474,N_4966);
nor U5167 (N_5167,N_3053,N_3055);
nand U5168 (N_5168,N_2573,N_4056);
or U5169 (N_5169,N_4856,N_3155);
nor U5170 (N_5170,N_3199,N_3449);
nor U5171 (N_5171,N_3876,N_4943);
and U5172 (N_5172,N_3829,N_2607);
or U5173 (N_5173,N_3941,N_2873);
nor U5174 (N_5174,N_3164,N_4880);
or U5175 (N_5175,N_4319,N_3783);
and U5176 (N_5176,N_2834,N_2771);
nor U5177 (N_5177,N_3909,N_4253);
and U5178 (N_5178,N_4085,N_3113);
and U5179 (N_5179,N_3145,N_4909);
and U5180 (N_5180,N_2571,N_3320);
nand U5181 (N_5181,N_4497,N_3945);
or U5182 (N_5182,N_4397,N_4271);
nand U5183 (N_5183,N_3470,N_2503);
and U5184 (N_5184,N_3240,N_3798);
nor U5185 (N_5185,N_4208,N_4036);
and U5186 (N_5186,N_3547,N_3122);
nor U5187 (N_5187,N_3201,N_3226);
nand U5188 (N_5188,N_4328,N_4112);
nand U5189 (N_5189,N_2592,N_4565);
nor U5190 (N_5190,N_3008,N_3501);
and U5191 (N_5191,N_2913,N_4002);
nand U5192 (N_5192,N_2688,N_3187);
nand U5193 (N_5193,N_3062,N_2504);
xnor U5194 (N_5194,N_2621,N_3478);
nor U5195 (N_5195,N_2837,N_3039);
and U5196 (N_5196,N_2850,N_4781);
nand U5197 (N_5197,N_4111,N_3230);
nand U5198 (N_5198,N_4218,N_3565);
or U5199 (N_5199,N_2509,N_3106);
or U5200 (N_5200,N_3621,N_3613);
nand U5201 (N_5201,N_3967,N_4795);
or U5202 (N_5202,N_3160,N_4578);
and U5203 (N_5203,N_4636,N_3068);
or U5204 (N_5204,N_4433,N_4703);
nand U5205 (N_5205,N_4684,N_2710);
xnor U5206 (N_5206,N_3144,N_2663);
nor U5207 (N_5207,N_4227,N_3081);
and U5208 (N_5208,N_2696,N_3350);
and U5209 (N_5209,N_4592,N_3815);
or U5210 (N_5210,N_4695,N_4358);
and U5211 (N_5211,N_2669,N_4225);
nand U5212 (N_5212,N_3836,N_4635);
or U5213 (N_5213,N_3636,N_4059);
nor U5214 (N_5214,N_2622,N_3650);
nand U5215 (N_5215,N_4008,N_4786);
nand U5216 (N_5216,N_4129,N_3602);
nor U5217 (N_5217,N_2662,N_4102);
nor U5218 (N_5218,N_2714,N_4409);
or U5219 (N_5219,N_3369,N_3714);
and U5220 (N_5220,N_3773,N_4958);
nor U5221 (N_5221,N_3337,N_4742);
and U5222 (N_5222,N_3756,N_2769);
xor U5223 (N_5223,N_4045,N_3590);
or U5224 (N_5224,N_3609,N_4083);
and U5225 (N_5225,N_3589,N_3196);
and U5226 (N_5226,N_4765,N_4003);
and U5227 (N_5227,N_3498,N_3040);
and U5228 (N_5228,N_2788,N_4663);
nor U5229 (N_5229,N_3744,N_4625);
and U5230 (N_5230,N_4133,N_4463);
or U5231 (N_5231,N_4476,N_4747);
or U5232 (N_5232,N_4422,N_2800);
and U5233 (N_5233,N_2904,N_3802);
nor U5234 (N_5234,N_3010,N_2968);
and U5235 (N_5235,N_4763,N_4146);
nand U5236 (N_5236,N_3513,N_3200);
nand U5237 (N_5237,N_3686,N_4120);
nor U5238 (N_5238,N_3992,N_4456);
nor U5239 (N_5239,N_3957,N_4534);
nand U5240 (N_5240,N_3415,N_4886);
or U5241 (N_5241,N_4491,N_2704);
nand U5242 (N_5242,N_3450,N_3174);
nor U5243 (N_5243,N_2624,N_4233);
nand U5244 (N_5244,N_4140,N_3911);
nand U5245 (N_5245,N_4642,N_3796);
and U5246 (N_5246,N_3816,N_4672);
nor U5247 (N_5247,N_4243,N_4244);
nand U5248 (N_5248,N_2914,N_4097);
or U5249 (N_5249,N_3688,N_4410);
nand U5250 (N_5250,N_4912,N_3036);
or U5251 (N_5251,N_4438,N_3161);
xnor U5252 (N_5252,N_4849,N_4487);
nand U5253 (N_5253,N_4154,N_4334);
nand U5254 (N_5254,N_3031,N_3803);
or U5255 (N_5255,N_4190,N_4632);
and U5256 (N_5256,N_2548,N_3924);
xor U5257 (N_5257,N_4877,N_3469);
nor U5258 (N_5258,N_4501,N_2925);
nor U5259 (N_5259,N_2554,N_4400);
nand U5260 (N_5260,N_2742,N_4152);
nor U5261 (N_5261,N_3740,N_4687);
nand U5262 (N_5262,N_4482,N_3711);
nor U5263 (N_5263,N_2749,N_4317);
nand U5264 (N_5264,N_4131,N_4307);
nand U5265 (N_5265,N_2839,N_4339);
and U5266 (N_5266,N_4285,N_4711);
and U5267 (N_5267,N_3659,N_2884);
nand U5268 (N_5268,N_2790,N_3779);
or U5269 (N_5269,N_4315,N_2764);
or U5270 (N_5270,N_4739,N_4735);
nor U5271 (N_5271,N_4477,N_2776);
nand U5272 (N_5272,N_4386,N_3871);
or U5273 (N_5273,N_4119,N_3363);
and U5274 (N_5274,N_4913,N_3927);
nor U5275 (N_5275,N_4068,N_4364);
nand U5276 (N_5276,N_4807,N_3452);
or U5277 (N_5277,N_3211,N_3573);
nor U5278 (N_5278,N_2674,N_3929);
nor U5279 (N_5279,N_2617,N_2532);
nor U5280 (N_5280,N_3353,N_4745);
nand U5281 (N_5281,N_3013,N_2920);
and U5282 (N_5282,N_4426,N_3734);
nor U5283 (N_5283,N_3151,N_3458);
and U5284 (N_5284,N_4604,N_4705);
and U5285 (N_5285,N_4853,N_3873);
or U5286 (N_5286,N_4936,N_3236);
nor U5287 (N_5287,N_4682,N_3462);
nor U5288 (N_5288,N_3352,N_4603);
nor U5289 (N_5289,N_3430,N_3572);
nor U5290 (N_5290,N_4744,N_4288);
or U5291 (N_5291,N_3724,N_4669);
nand U5292 (N_5292,N_4266,N_4143);
xnor U5293 (N_5293,N_4910,N_4441);
nand U5294 (N_5294,N_4783,N_4325);
nand U5295 (N_5295,N_4757,N_3638);
nand U5296 (N_5296,N_4383,N_3351);
or U5297 (N_5297,N_2651,N_3365);
and U5298 (N_5298,N_3988,N_4301);
nand U5299 (N_5299,N_4823,N_3376);
or U5300 (N_5300,N_2522,N_3280);
nor U5301 (N_5301,N_4024,N_4485);
and U5302 (N_5302,N_3412,N_4953);
or U5303 (N_5303,N_3719,N_4858);
and U5304 (N_5304,N_4037,N_3972);
or U5305 (N_5305,N_4612,N_2826);
nor U5306 (N_5306,N_4774,N_4287);
nand U5307 (N_5307,N_3561,N_4210);
nand U5308 (N_5308,N_3043,N_3075);
nand U5309 (N_5309,N_4429,N_3481);
xor U5310 (N_5310,N_2927,N_4911);
nand U5311 (N_5311,N_2825,N_2664);
and U5312 (N_5312,N_2538,N_2594);
or U5313 (N_5313,N_2615,N_4706);
nor U5314 (N_5314,N_3134,N_3026);
and U5315 (N_5315,N_2574,N_4543);
and U5316 (N_5316,N_4975,N_4698);
nand U5317 (N_5317,N_2811,N_2791);
or U5318 (N_5318,N_3884,N_3869);
nor U5319 (N_5319,N_3761,N_2585);
and U5320 (N_5320,N_3265,N_4845);
or U5321 (N_5321,N_4896,N_4012);
nand U5322 (N_5322,N_4860,N_2613);
nand U5323 (N_5323,N_3003,N_4797);
or U5324 (N_5324,N_4289,N_3887);
or U5325 (N_5325,N_4256,N_2557);
nand U5326 (N_5326,N_2758,N_3794);
nand U5327 (N_5327,N_4960,N_3204);
and U5328 (N_5328,N_3770,N_3181);
or U5329 (N_5329,N_3998,N_3738);
and U5330 (N_5330,N_4848,N_4661);
nand U5331 (N_5331,N_4343,N_3413);
nand U5332 (N_5332,N_3690,N_2792);
nor U5333 (N_5333,N_4892,N_4035);
and U5334 (N_5334,N_3697,N_3125);
nor U5335 (N_5335,N_2836,N_3165);
and U5336 (N_5336,N_4028,N_3749);
nand U5337 (N_5337,N_2508,N_2833);
nand U5338 (N_5338,N_4581,N_4030);
nor U5339 (N_5339,N_3655,N_3661);
nor U5340 (N_5340,N_2616,N_3167);
and U5341 (N_5341,N_4802,N_4488);
nor U5342 (N_5342,N_4633,N_3764);
nor U5343 (N_5343,N_2902,N_4567);
and U5344 (N_5344,N_4392,N_4327);
or U5345 (N_5345,N_4691,N_3942);
and U5346 (N_5346,N_2804,N_3669);
nor U5347 (N_5347,N_2715,N_2985);
or U5348 (N_5348,N_4957,N_3986);
or U5349 (N_5349,N_3243,N_4504);
nor U5350 (N_5350,N_4622,N_4424);
or U5351 (N_5351,N_3130,N_2546);
and U5352 (N_5352,N_2806,N_2589);
or U5353 (N_5353,N_4824,N_3234);
nand U5354 (N_5354,N_4144,N_4571);
nand U5355 (N_5355,N_4722,N_4959);
and U5356 (N_5356,N_3978,N_3023);
and U5357 (N_5357,N_3235,N_2683);
nor U5358 (N_5358,N_3939,N_3033);
nand U5359 (N_5359,N_3197,N_2793);
nand U5360 (N_5360,N_2886,N_3519);
and U5361 (N_5361,N_4659,N_3382);
nor U5362 (N_5362,N_4866,N_3098);
nand U5363 (N_5363,N_2561,N_2917);
or U5364 (N_5364,N_3463,N_2919);
and U5365 (N_5365,N_4440,N_3838);
nand U5366 (N_5366,N_2865,N_3554);
xor U5367 (N_5367,N_3451,N_4513);
nand U5368 (N_5368,N_3671,N_2910);
and U5369 (N_5369,N_3386,N_2513);
nand U5370 (N_5370,N_2830,N_4309);
and U5371 (N_5371,N_3607,N_2888);
or U5372 (N_5372,N_3667,N_2741);
nand U5373 (N_5373,N_4075,N_4925);
nor U5374 (N_5374,N_2860,N_4505);
and U5375 (N_5375,N_4443,N_2952);
or U5376 (N_5376,N_3218,N_3616);
and U5377 (N_5377,N_4893,N_4754);
and U5378 (N_5378,N_4922,N_3707);
or U5379 (N_5379,N_3185,N_3586);
nor U5380 (N_5380,N_2653,N_2726);
nand U5381 (N_5381,N_4486,N_4775);
or U5382 (N_5382,N_3782,N_2529);
or U5383 (N_5383,N_4335,N_4004);
nor U5384 (N_5384,N_3631,N_2737);
or U5385 (N_5385,N_3366,N_3805);
nand U5386 (N_5386,N_2525,N_4381);
or U5387 (N_5387,N_3492,N_3227);
or U5388 (N_5388,N_4274,N_3107);
nand U5389 (N_5389,N_3526,N_3921);
nor U5390 (N_5390,N_4182,N_3955);
and U5391 (N_5391,N_3587,N_2772);
nor U5392 (N_5392,N_4793,N_4707);
nor U5393 (N_5393,N_4471,N_4656);
or U5394 (N_5394,N_4623,N_4621);
nand U5395 (N_5395,N_4538,N_3504);
nor U5396 (N_5396,N_3261,N_4286);
nor U5397 (N_5397,N_3932,N_4013);
nand U5398 (N_5398,N_3421,N_4018);
nor U5399 (N_5399,N_2956,N_4874);
and U5400 (N_5400,N_3179,N_2835);
nor U5401 (N_5401,N_3049,N_4819);
xor U5402 (N_5402,N_4573,N_4627);
nor U5403 (N_5403,N_4718,N_3441);
or U5404 (N_5404,N_4407,N_3156);
and U5405 (N_5405,N_4738,N_4155);
and U5406 (N_5406,N_2626,N_4916);
and U5407 (N_5407,N_3431,N_2939);
or U5408 (N_5408,N_3250,N_2721);
nand U5409 (N_5409,N_2640,N_4153);
or U5410 (N_5410,N_2641,N_3057);
and U5411 (N_5411,N_3009,N_4826);
or U5412 (N_5412,N_3038,N_3030);
nor U5413 (N_5413,N_2729,N_3269);
and U5414 (N_5414,N_4479,N_2799);
and U5415 (N_5415,N_2785,N_2610);
and U5416 (N_5416,N_2814,N_4549);
nor U5417 (N_5417,N_3074,N_3933);
nor U5418 (N_5418,N_3379,N_2988);
nor U5419 (N_5419,N_4982,N_3946);
xor U5420 (N_5420,N_3847,N_4638);
nand U5421 (N_5421,N_4961,N_4483);
or U5422 (N_5422,N_3785,N_3345);
or U5423 (N_5423,N_4361,N_3658);
nand U5424 (N_5424,N_3126,N_3765);
and U5425 (N_5425,N_3078,N_3475);
nand U5426 (N_5426,N_4785,N_4356);
or U5427 (N_5427,N_3028,N_3618);
nand U5428 (N_5428,N_4847,N_2536);
or U5429 (N_5429,N_4694,N_4679);
nand U5430 (N_5430,N_3949,N_4278);
and U5431 (N_5431,N_4947,N_3476);
or U5432 (N_5432,N_3315,N_3456);
and U5433 (N_5433,N_4316,N_2630);
and U5434 (N_5434,N_3330,N_4168);
nor U5435 (N_5435,N_2684,N_2718);
nand U5436 (N_5436,N_2713,N_4177);
or U5437 (N_5437,N_4898,N_4685);
nor U5438 (N_5438,N_3005,N_3818);
nor U5439 (N_5439,N_3891,N_3825);
and U5440 (N_5440,N_3600,N_3076);
nand U5441 (N_5441,N_4188,N_2849);
nand U5442 (N_5442,N_3401,N_2856);
and U5443 (N_5443,N_2677,N_4416);
nor U5444 (N_5444,N_4889,N_4926);
and U5445 (N_5445,N_4841,N_4379);
nand U5446 (N_5446,N_2894,N_4639);
nor U5447 (N_5447,N_3642,N_4391);
or U5448 (N_5448,N_2728,N_3983);
nand U5449 (N_5449,N_3880,N_3534);
and U5450 (N_5450,N_4585,N_3402);
or U5451 (N_5451,N_4403,N_3675);
and U5452 (N_5452,N_4969,N_4235);
nand U5453 (N_5453,N_3666,N_2541);
or U5454 (N_5454,N_3699,N_3698);
or U5455 (N_5455,N_3814,N_3940);
or U5456 (N_5456,N_2646,N_3205);
nor U5457 (N_5457,N_4324,N_3605);
xnor U5458 (N_5458,N_2523,N_2588);
or U5459 (N_5459,N_2586,N_2526);
and U5460 (N_5460,N_2828,N_4562);
nand U5461 (N_5461,N_4796,N_3222);
or U5462 (N_5462,N_3042,N_4336);
nor U5463 (N_5463,N_4995,N_3637);
and U5464 (N_5464,N_2689,N_4248);
and U5465 (N_5465,N_4670,N_2962);
nor U5466 (N_5466,N_4353,N_3276);
nand U5467 (N_5467,N_4194,N_4128);
and U5468 (N_5468,N_4956,N_4401);
nand U5469 (N_5469,N_2603,N_2924);
nor U5470 (N_5470,N_3391,N_4665);
nand U5471 (N_5471,N_3321,N_3024);
nor U5472 (N_5472,N_4655,N_3270);
nand U5473 (N_5473,N_3312,N_2966);
nor U5474 (N_5474,N_3571,N_4350);
nor U5475 (N_5475,N_4791,N_4557);
nor U5476 (N_5476,N_2572,N_4475);
or U5477 (N_5477,N_4832,N_3712);
nand U5478 (N_5478,N_2995,N_2568);
or U5479 (N_5479,N_3262,N_2634);
and U5480 (N_5480,N_4697,N_3990);
nand U5481 (N_5481,N_2890,N_4628);
and U5482 (N_5482,N_3396,N_4165);
or U5483 (N_5483,N_3855,N_2569);
and U5484 (N_5484,N_3375,N_3676);
and U5485 (N_5485,N_4547,N_2880);
nand U5486 (N_5486,N_4686,N_2595);
and U5487 (N_5487,N_4749,N_3508);
and U5488 (N_5488,N_3466,N_3541);
or U5489 (N_5489,N_3035,N_3173);
and U5490 (N_5490,N_4550,N_3302);
and U5491 (N_5491,N_2543,N_3867);
or U5492 (N_5492,N_2701,N_3393);
or U5493 (N_5493,N_3289,N_3152);
or U5494 (N_5494,N_3537,N_3828);
nand U5495 (N_5495,N_3546,N_3082);
and U5496 (N_5496,N_3423,N_3178);
nand U5497 (N_5497,N_3583,N_3408);
nand U5498 (N_5498,N_4262,N_3670);
and U5499 (N_5499,N_3716,N_2843);
nor U5500 (N_5500,N_4260,N_4552);
nand U5501 (N_5501,N_4298,N_2944);
or U5502 (N_5502,N_2755,N_2964);
and U5503 (N_5503,N_3245,N_3182);
nor U5504 (N_5504,N_4032,N_3296);
nand U5505 (N_5505,N_4367,N_3215);
or U5506 (N_5506,N_2943,N_4093);
or U5507 (N_5507,N_2552,N_4326);
nand U5508 (N_5508,N_3883,N_3538);
or U5509 (N_5509,N_3678,N_3486);
nor U5510 (N_5510,N_3959,N_2960);
and U5511 (N_5511,N_4322,N_3656);
or U5512 (N_5512,N_4634,N_3051);
and U5513 (N_5513,N_4283,N_3139);
nor U5514 (N_5514,N_4404,N_4688);
and U5515 (N_5515,N_2816,N_3091);
and U5516 (N_5516,N_2817,N_4945);
nor U5517 (N_5517,N_4313,N_2692);
nand U5518 (N_5518,N_4297,N_3827);
nor U5519 (N_5519,N_4902,N_4933);
nand U5520 (N_5520,N_3432,N_4109);
or U5521 (N_5521,N_3256,N_3870);
and U5522 (N_5522,N_2932,N_4178);
or U5523 (N_5523,N_3136,N_2891);
or U5524 (N_5524,N_3212,N_4306);
or U5525 (N_5525,N_4701,N_3427);
or U5526 (N_5526,N_3180,N_3443);
nand U5527 (N_5527,N_3071,N_2931);
nand U5528 (N_5528,N_4643,N_4206);
nor U5529 (N_5529,N_2845,N_4939);
nand U5530 (N_5530,N_4829,N_3696);
nor U5531 (N_5531,N_4520,N_4034);
or U5532 (N_5532,N_4159,N_4872);
and U5533 (N_5533,N_3239,N_2519);
nor U5534 (N_5534,N_4412,N_3511);
and U5535 (N_5535,N_4500,N_2597);
nor U5536 (N_5536,N_3790,N_4333);
and U5537 (N_5537,N_3468,N_3237);
and U5538 (N_5538,N_3046,N_3646);
nand U5539 (N_5539,N_2980,N_4089);
or U5540 (N_5540,N_2868,N_4329);
nand U5541 (N_5541,N_3268,N_3700);
nor U5542 (N_5542,N_3835,N_2802);
nand U5543 (N_5543,N_4985,N_2537);
and U5544 (N_5544,N_4114,N_2906);
and U5545 (N_5545,N_3603,N_4827);
nand U5546 (N_5546,N_3326,N_2716);
nand U5547 (N_5547,N_4349,N_3093);
nor U5548 (N_5548,N_3021,N_4553);
nand U5549 (N_5549,N_4435,N_3570);
or U5550 (N_5550,N_4907,N_4528);
and U5551 (N_5551,N_4869,N_4580);
and U5552 (N_5552,N_3329,N_4668);
and U5553 (N_5553,N_2652,N_4981);
nor U5554 (N_5554,N_4662,N_4771);
nor U5555 (N_5555,N_3069,N_3387);
and U5556 (N_5556,N_3811,N_3241);
and U5557 (N_5557,N_4980,N_4493);
and U5558 (N_5558,N_3209,N_4202);
nor U5559 (N_5559,N_3629,N_3857);
nor U5560 (N_5560,N_2697,N_4555);
and U5561 (N_5561,N_4806,N_2668);
nor U5562 (N_5562,N_3530,N_3001);
and U5563 (N_5563,N_3643,N_4066);
or U5564 (N_5564,N_4755,N_2892);
nand U5565 (N_5565,N_3045,N_4312);
or U5566 (N_5566,N_2997,N_3555);
nor U5567 (N_5567,N_3953,N_2867);
or U5568 (N_5568,N_3448,N_2794);
or U5569 (N_5569,N_3758,N_3993);
nor U5570 (N_5570,N_4252,N_2803);
nor U5571 (N_5571,N_4070,N_4756);
nand U5572 (N_5572,N_4530,N_4589);
nand U5573 (N_5573,N_3984,N_4752);
and U5574 (N_5574,N_3338,N_4360);
nor U5575 (N_5575,N_4291,N_2922);
or U5576 (N_5576,N_4280,N_4232);
nand U5577 (N_5577,N_4503,N_4600);
nand U5578 (N_5578,N_4496,N_3496);
and U5579 (N_5579,N_4063,N_4241);
or U5580 (N_5580,N_4782,N_3283);
and U5581 (N_5581,N_3022,N_4414);
nand U5582 (N_5582,N_4719,N_4716);
nor U5583 (N_5583,N_4044,N_4769);
or U5584 (N_5584,N_3244,N_2895);
nor U5585 (N_5585,N_4870,N_4310);
nand U5586 (N_5586,N_4545,N_4814);
nand U5587 (N_5587,N_3706,N_3778);
xnor U5588 (N_5588,N_3495,N_4803);
nor U5589 (N_5589,N_2612,N_2879);
and U5590 (N_5590,N_3679,N_4929);
and U5591 (N_5591,N_4103,N_3394);
or U5592 (N_5592,N_3833,N_3739);
or U5593 (N_5593,N_4425,N_4088);
or U5594 (N_5594,N_4941,N_4411);
or U5595 (N_5595,N_4556,N_2882);
and U5596 (N_5596,N_3727,N_3653);
nor U5597 (N_5597,N_4394,N_3813);
nor U5598 (N_5598,N_3923,N_2604);
nor U5599 (N_5599,N_4736,N_4055);
and U5600 (N_5600,N_3665,N_4773);
nor U5601 (N_5601,N_4813,N_4010);
and U5602 (N_5602,N_4020,N_4027);
nand U5603 (N_5603,N_4535,N_4048);
nor U5604 (N_5604,N_4561,N_3824);
or U5605 (N_5605,N_3088,N_2720);
and U5606 (N_5606,N_3788,N_4467);
nand U5607 (N_5607,N_3822,N_4741);
or U5608 (N_5608,N_3969,N_4130);
nor U5609 (N_5609,N_4047,N_4817);
or U5610 (N_5610,N_3318,N_3271);
or U5611 (N_5611,N_4950,N_2875);
and U5612 (N_5612,N_4879,N_4836);
and U5613 (N_5613,N_4901,N_4993);
nand U5614 (N_5614,N_3556,N_4839);
nand U5615 (N_5615,N_2738,N_3029);
or U5616 (N_5616,N_4618,N_4664);
nand U5617 (N_5617,N_2930,N_4022);
and U5618 (N_5618,N_4890,N_2866);
or U5619 (N_5619,N_3433,N_4548);
and U5620 (N_5620,N_2635,N_2636);
nor U5621 (N_5621,N_4091,N_4115);
and U5622 (N_5622,N_4546,N_4049);
nor U5623 (N_5623,N_4644,N_3733);
nand U5624 (N_5624,N_3612,N_4991);
nor U5625 (N_5625,N_3214,N_3175);
and U5626 (N_5626,N_4891,N_3169);
or U5627 (N_5627,N_2656,N_2685);
nand U5628 (N_5628,N_4979,N_3286);
and U5629 (N_5629,N_3016,N_2754);
and U5630 (N_5630,N_4999,N_3528);
nor U5631 (N_5631,N_2609,N_3221);
nor U5632 (N_5632,N_2591,N_3860);
nor U5633 (N_5633,N_3722,N_4459);
nand U5634 (N_5634,N_3192,N_3277);
and U5635 (N_5635,N_4224,N_4885);
nand U5636 (N_5636,N_3954,N_4163);
nand U5637 (N_5637,N_4305,N_3520);
and U5638 (N_5638,N_4038,N_3809);
or U5639 (N_5639,N_3725,N_4708);
nand U5640 (N_5640,N_3973,N_2723);
nand U5641 (N_5641,N_3417,N_3875);
nand U5642 (N_5642,N_4564,N_4284);
nand U5643 (N_5643,N_4365,N_3484);
nand U5644 (N_5644,N_3473,N_4213);
nand U5645 (N_5645,N_4834,N_2655);
or U5646 (N_5646,N_4746,N_3132);
and U5647 (N_5647,N_2858,N_3140);
and U5648 (N_5648,N_3238,N_3989);
nand U5649 (N_5649,N_4185,N_4180);
nand U5650 (N_5650,N_4850,N_4042);
nand U5651 (N_5651,N_3109,N_3889);
or U5652 (N_5652,N_3213,N_4490);
nor U5653 (N_5653,N_4290,N_2958);
and U5654 (N_5654,N_3750,N_4994);
and U5655 (N_5655,N_3841,N_4551);
nor U5656 (N_5656,N_3216,N_4965);
nor U5657 (N_5657,N_4894,N_3348);
xor U5658 (N_5658,N_3410,N_2823);
xnor U5659 (N_5659,N_4434,N_4584);
nor U5660 (N_5660,N_2903,N_4368);
nand U5661 (N_5661,N_3792,N_4007);
and U5662 (N_5662,N_2987,N_3886);
and U5663 (N_5663,N_4734,N_4935);
nand U5664 (N_5664,N_2978,N_3293);
or U5665 (N_5665,N_3327,N_3385);
nor U5666 (N_5666,N_3588,N_3987);
or U5667 (N_5667,N_4652,N_4468);
nor U5668 (N_5668,N_3349,N_4387);
nor U5669 (N_5669,N_3866,N_2549);
or U5670 (N_5670,N_3411,N_3507);
or U5671 (N_5671,N_3355,N_3837);
or U5672 (N_5672,N_4937,N_4822);
and U5673 (N_5673,N_3594,N_3414);
or U5674 (N_5674,N_3251,N_4204);
nor U5675 (N_5675,N_4342,N_4231);
xor U5676 (N_5676,N_3219,N_4983);
or U5677 (N_5677,N_3500,N_3503);
or U5678 (N_5678,N_3444,N_2516);
nand U5679 (N_5679,N_2584,N_4214);
or U5680 (N_5680,N_4709,N_4611);
nand U5681 (N_5681,N_4132,N_4521);
nor U5682 (N_5682,N_4229,N_2847);
or U5683 (N_5683,N_4236,N_4099);
nand U5684 (N_5684,N_3100,N_4681);
nor U5685 (N_5685,N_4710,N_2598);
or U5686 (N_5686,N_3114,N_3680);
nand U5687 (N_5687,N_2578,N_4620);
and U5688 (N_5688,N_3012,N_4559);
nor U5689 (N_5689,N_4226,N_4617);
and U5690 (N_5690,N_3807,N_3709);
nor U5691 (N_5691,N_3892,N_4428);
and U5692 (N_5692,N_4954,N_2731);
nor U5693 (N_5693,N_3483,N_3996);
or U5694 (N_5694,N_3354,N_3731);
nor U5695 (N_5695,N_4439,N_3457);
or U5696 (N_5696,N_2992,N_2507);
or U5697 (N_5697,N_3317,N_3388);
or U5698 (N_5698,N_3755,N_2813);
nand U5699 (N_5699,N_4160,N_4184);
and U5700 (N_5700,N_4081,N_4311);
or U5701 (N_5701,N_3831,N_3682);
and U5702 (N_5702,N_3582,N_4494);
xnor U5703 (N_5703,N_2945,N_3341);
nand U5704 (N_5704,N_3418,N_2807);
nor U5705 (N_5705,N_3020,N_4940);
and U5706 (N_5706,N_4527,N_2563);
or U5707 (N_5707,N_2970,N_3472);
or U5708 (N_5708,N_3730,N_3054);
or U5709 (N_5709,N_4646,N_4275);
or U5710 (N_5710,N_4949,N_3897);
nand U5711 (N_5711,N_3623,N_3628);
nand U5712 (N_5712,N_4460,N_4838);
nand U5713 (N_5713,N_4465,N_2511);
and U5714 (N_5714,N_3313,N_3908);
or U5715 (N_5715,N_2562,N_3395);
or U5716 (N_5716,N_3094,N_4001);
and U5717 (N_5717,N_4029,N_3830);
nand U5718 (N_5718,N_3918,N_4464);
nor U5719 (N_5719,N_2938,N_4810);
nand U5720 (N_5720,N_4450,N_3902);
xor U5721 (N_5721,N_4273,N_4987);
or U5722 (N_5722,N_4077,N_2533);
and U5723 (N_5723,N_2993,N_3509);
or U5724 (N_5724,N_3859,N_3685);
nand U5725 (N_5725,N_4648,N_4651);
nor U5726 (N_5726,N_2976,N_4258);
nor U5727 (N_5727,N_3663,N_3840);
and U5728 (N_5728,N_3279,N_4740);
and U5729 (N_5729,N_3963,N_3753);
or U5730 (N_5730,N_4192,N_4812);
nor U5731 (N_5731,N_4215,N_4723);
nor U5732 (N_5732,N_4341,N_3931);
or U5733 (N_5733,N_3460,N_4370);
and U5734 (N_5734,N_3027,N_4171);
nor U5735 (N_5735,N_2855,N_4474);
and U5736 (N_5736,N_4523,N_3163);
or U5737 (N_5737,N_4815,N_3874);
or U5738 (N_5738,N_4990,N_4675);
xnor U5739 (N_5739,N_4308,N_2687);
or U5740 (N_5740,N_2575,N_3910);
or U5741 (N_5741,N_3704,N_3117);
and U5742 (N_5742,N_4509,N_4043);
nand U5743 (N_5743,N_4844,N_2824);
nand U5744 (N_5744,N_4016,N_3129);
and U5745 (N_5745,N_4512,N_4624);
or U5746 (N_5746,N_4355,N_3189);
and U5747 (N_5747,N_4862,N_2901);
or U5748 (N_5748,N_2761,N_4591);
and U5749 (N_5749,N_4216,N_2972);
nor U5750 (N_5750,N_3542,N_3879);
or U5751 (N_5751,N_3077,N_3170);
or U5752 (N_5752,N_3872,N_4220);
and U5753 (N_5753,N_2633,N_4388);
and U5754 (N_5754,N_4667,N_4100);
or U5755 (N_5755,N_3751,N_3059);
nor U5756 (N_5756,N_3228,N_4366);
nand U5757 (N_5757,N_2673,N_4867);
or U5758 (N_5758,N_4117,N_4948);
and U5759 (N_5759,N_4345,N_3487);
nor U5760 (N_5760,N_2582,N_3303);
or U5761 (N_5761,N_4110,N_2818);
and U5762 (N_5762,N_4899,N_3784);
nor U5763 (N_5763,N_2905,N_3800);
nand U5764 (N_5764,N_4302,N_3202);
or U5765 (N_5765,N_4234,N_4931);
and U5766 (N_5766,N_4522,N_4452);
or U5767 (N_5767,N_3995,N_2660);
nor U5768 (N_5768,N_4906,N_4318);
or U5769 (N_5769,N_4671,N_4448);
and U5770 (N_5770,N_3708,N_2999);
and U5771 (N_5771,N_2501,N_4700);
or U5772 (N_5772,N_4378,N_3741);
and U5773 (N_5773,N_3593,N_3397);
nor U5774 (N_5774,N_3428,N_2822);
or U5775 (N_5775,N_2783,N_4579);
and U5776 (N_5776,N_4293,N_3971);
nor U5777 (N_5777,N_4105,N_3491);
and U5778 (N_5778,N_4843,N_4457);
and U5779 (N_5779,N_3377,N_4714);
nand U5780 (N_5780,N_3566,N_2645);
nor U5781 (N_5781,N_3521,N_4338);
nor U5782 (N_5782,N_3217,N_3171);
nand U5783 (N_5783,N_4362,N_3177);
nor U5784 (N_5784,N_3297,N_4970);
and U5785 (N_5785,N_3757,N_2647);
nand U5786 (N_5786,N_4415,N_2502);
and U5787 (N_5787,N_4502,N_4158);
or U5788 (N_5788,N_4161,N_2907);
or U5789 (N_5789,N_2848,N_4944);
nand U5790 (N_5790,N_3735,N_2768);
or U5791 (N_5791,N_3579,N_3611);
nand U5792 (N_5792,N_4730,N_3342);
nor U5793 (N_5793,N_2740,N_4299);
nand U5794 (N_5794,N_2643,N_3264);
and U5795 (N_5795,N_4607,N_4481);
nand U5796 (N_5796,N_4221,N_3527);
and U5797 (N_5797,N_2819,N_2815);
or U5798 (N_5798,N_4382,N_3762);
nor U5799 (N_5799,N_2518,N_4458);
nor U5800 (N_5800,N_4590,N_2887);
nand U5801 (N_5801,N_3339,N_3158);
nand U5802 (N_5802,N_3047,N_4189);
and U5803 (N_5803,N_2676,N_4780);
and U5804 (N_5804,N_4861,N_4080);
nor U5805 (N_5805,N_3975,N_2961);
nor U5806 (N_5806,N_3242,N_2990);
nand U5807 (N_5807,N_4721,N_3898);
nand U5808 (N_5808,N_3291,N_2608);
or U5809 (N_5809,N_3193,N_3328);
nor U5810 (N_5810,N_3632,N_3347);
or U5811 (N_5811,N_3195,N_3332);
or U5812 (N_5812,N_4510,N_3524);
and U5813 (N_5813,N_4921,N_3083);
or U5814 (N_5814,N_4436,N_4799);
or U5815 (N_5815,N_4998,N_2916);
and U5816 (N_5816,N_3493,N_3808);
nand U5817 (N_5817,N_3539,N_3266);
or U5818 (N_5818,N_3804,N_3745);
nor U5819 (N_5819,N_4385,N_2762);
nor U5820 (N_5820,N_4637,N_2717);
nor U5821 (N_5821,N_3850,N_4868);
and U5822 (N_5822,N_2531,N_3063);
or U5823 (N_5823,N_3574,N_2743);
nand U5824 (N_5824,N_3080,N_4952);
or U5825 (N_5825,N_3207,N_3371);
nand U5826 (N_5826,N_3273,N_3384);
or U5827 (N_5827,N_4614,N_2547);
nor U5828 (N_5828,N_4172,N_2505);
and U5829 (N_5829,N_3445,N_3797);
and U5830 (N_5830,N_3858,N_4629);
nand U5831 (N_5831,N_3569,N_2935);
nor U5832 (N_5832,N_2694,N_3064);
or U5833 (N_5833,N_3052,N_4451);
and U5834 (N_5834,N_4025,N_4615);
or U5835 (N_5835,N_2951,N_4587);
and U5836 (N_5836,N_4787,N_4794);
nand U5837 (N_5837,N_2838,N_4373);
nor U5838 (N_5838,N_3619,N_2606);
or U5839 (N_5839,N_4654,N_4240);
nand U5840 (N_5840,N_2942,N_2915);
and U5841 (N_5841,N_4597,N_3426);
and U5842 (N_5842,N_2940,N_4139);
and U5843 (N_5843,N_3720,N_4492);
nor U5844 (N_5844,N_4569,N_3087);
or U5845 (N_5845,N_2675,N_4851);
nor U5846 (N_5846,N_4601,N_4732);
and U5847 (N_5847,N_4914,N_3135);
nand U5848 (N_5848,N_3208,N_2928);
and U5849 (N_5849,N_4657,N_3592);
or U5850 (N_5850,N_4789,N_3461);
or U5851 (N_5851,N_3017,N_4717);
or U5852 (N_5852,N_2599,N_4820);
nor U5853 (N_5853,N_4121,N_3563);
nand U5854 (N_5854,N_3903,N_3105);
and U5855 (N_5855,N_3999,N_4712);
or U5856 (N_5856,N_4542,N_3323);
nor U5857 (N_5857,N_4766,N_2706);
xor U5858 (N_5858,N_3488,N_3183);
nand U5859 (N_5859,N_3505,N_3729);
nor U5860 (N_5860,N_3767,N_4014);
nand U5861 (N_5861,N_4396,N_4658);
or U5862 (N_5862,N_4825,N_2998);
and U5863 (N_5863,N_4517,N_3845);
and U5864 (N_5864,N_3826,N_3007);
or U5865 (N_5865,N_3935,N_3307);
xnor U5866 (N_5866,N_4201,N_4645);
nor U5867 (N_5867,N_3529,N_2707);
or U5868 (N_5868,N_3842,N_3275);
nand U5869 (N_5869,N_3249,N_3115);
or U5870 (N_5870,N_3747,N_4246);
nand U5871 (N_5871,N_3956,N_2989);
or U5872 (N_5872,N_3960,N_4784);
and U5873 (N_5873,N_4314,N_3919);
or U5874 (N_5874,N_4472,N_3695);
nor U5875 (N_5875,N_3248,N_4113);
and U5876 (N_5876,N_3111,N_2670);
or U5877 (N_5877,N_3224,N_3118);
nand U5878 (N_5878,N_3400,N_2948);
nor U5879 (N_5879,N_4026,N_4237);
or U5880 (N_5880,N_4883,N_2810);
and U5881 (N_5881,N_3673,N_3560);
nand U5882 (N_5882,N_3374,N_3878);
and U5883 (N_5883,N_4882,N_3112);
xor U5884 (N_5884,N_2667,N_4674);
and U5885 (N_5885,N_4855,N_2565);
nand U5886 (N_5886,N_3979,N_2971);
or U5887 (N_5887,N_2889,N_3920);
nor U5888 (N_5888,N_3168,N_2534);
nand U5889 (N_5889,N_3552,N_3333);
and U5890 (N_5890,N_3937,N_4072);
nor U5891 (N_5891,N_3849,N_2746);
and U5892 (N_5892,N_3308,N_2921);
or U5893 (N_5893,N_3634,N_3490);
or U5894 (N_5894,N_2883,N_4480);
nand U5895 (N_5895,N_4242,N_3220);
and U5896 (N_5896,N_2535,N_3793);
nor U5897 (N_5897,N_3780,N_4136);
or U5898 (N_5898,N_3801,N_4857);
and U5899 (N_5899,N_4586,N_4748);
nor U5900 (N_5900,N_4173,N_2893);
nor U5901 (N_5901,N_4296,N_4065);
or U5902 (N_5902,N_4039,N_4149);
and U5903 (N_5903,N_2524,N_3976);
nand U5904 (N_5904,N_4696,N_2954);
nor U5905 (N_5905,N_4608,N_3516);
nor U5906 (N_5906,N_2709,N_3123);
nor U5907 (N_5907,N_2957,N_2745);
nand U5908 (N_5908,N_4137,N_3206);
and U5909 (N_5909,N_2644,N_2909);
or U5910 (N_5910,N_4918,N_3567);
or U5911 (N_5911,N_4384,N_3422);
nor U5912 (N_5912,N_3994,N_3437);
nand U5913 (N_5913,N_4864,N_4134);
and U5914 (N_5914,N_2661,N_2619);
nand U5915 (N_5915,N_3557,N_4599);
nand U5916 (N_5916,N_4978,N_4508);
nor U5917 (N_5917,N_2991,N_2853);
or U5918 (N_5918,N_2686,N_2520);
or U5919 (N_5919,N_3786,N_3599);
nand U5920 (N_5920,N_3073,N_3948);
nand U5921 (N_5921,N_2983,N_3693);
nor U5922 (N_5922,N_3564,N_3856);
nor U5923 (N_5923,N_4666,N_4238);
or U5924 (N_5924,N_3300,N_4005);
nand U5925 (N_5925,N_4304,N_4357);
or U5926 (N_5926,N_4887,N_4245);
or U5927 (N_5927,N_2777,N_3641);
and U5928 (N_5928,N_3108,N_4532);
nand U5929 (N_5929,N_4753,N_4052);
nor U5930 (N_5930,N_4575,N_3997);
nor U5931 (N_5931,N_3502,N_4351);
nand U5932 (N_5932,N_3597,N_2861);
and U5933 (N_5933,N_4540,N_3647);
and U5934 (N_5934,N_4563,N_4393);
or U5935 (N_5935,N_2539,N_3882);
or U5936 (N_5936,N_4539,N_4495);
xnor U5937 (N_5937,N_4069,N_2870);
xor U5938 (N_5938,N_2654,N_4588);
or U5939 (N_5939,N_3015,N_4167);
nand U5940 (N_5940,N_3056,N_2695);
and U5941 (N_5941,N_3065,N_2699);
nor U5942 (N_5942,N_2735,N_3522);
nor U5943 (N_5943,N_3772,N_2929);
or U5944 (N_5944,N_2596,N_4598);
or U5945 (N_5945,N_2500,N_3465);
nor U5946 (N_5946,N_3585,N_4380);
nor U5947 (N_5947,N_2698,N_3718);
or U5948 (N_5948,N_2827,N_3635);
nor U5949 (N_5949,N_3548,N_3002);
nand U5950 (N_5950,N_3258,N_4726);
and U5951 (N_5951,N_3128,N_4371);
and U5952 (N_5952,N_4352,N_4461);
nor U5953 (N_5953,N_2666,N_4613);
nand U5954 (N_5954,N_3316,N_3930);
and U5955 (N_5955,N_3769,N_3439);
or U5956 (N_5956,N_2986,N_4727);
or U5957 (N_5957,N_3198,N_3404);
nand U5958 (N_5958,N_4267,N_3578);
nor U5959 (N_5959,N_2842,N_3343);
nand U5960 (N_5960,N_4449,N_4145);
and U5961 (N_5961,N_2805,N_4331);
nand U5962 (N_5962,N_3677,N_2881);
and U5963 (N_5963,N_3247,N_3633);
or U5964 (N_5964,N_4724,N_3506);
nor U5965 (N_5965,N_3832,N_3346);
and U5966 (N_5966,N_4750,N_4054);
and U5967 (N_5967,N_2620,N_4166);
nand U5968 (N_5968,N_3846,N_2631);
nand U5969 (N_5969,N_2730,N_2979);
nor U5970 (N_5970,N_4609,N_3962);
and U5971 (N_5971,N_3759,N_2751);
nor U5972 (N_5972,N_3914,N_4418);
or U5973 (N_5973,N_4631,N_3159);
nand U5974 (N_5974,N_2678,N_4187);
and U5975 (N_5975,N_4506,N_4837);
and U5976 (N_5976,N_3281,N_3340);
or U5977 (N_5977,N_3325,N_4098);
and U5978 (N_5978,N_3116,N_3257);
nand U5979 (N_5979,N_3018,N_2566);
or U5980 (N_5980,N_3674,N_4205);
nor U5981 (N_5981,N_3086,N_2766);
nor U5982 (N_5982,N_4321,N_3806);
nand U5983 (N_5983,N_4865,N_3543);
or U5984 (N_5984,N_4442,N_4276);
nand U5985 (N_5985,N_3888,N_4096);
nand U5986 (N_5986,N_4023,N_3692);
nand U5987 (N_5987,N_3596,N_3952);
and U5988 (N_5988,N_4582,N_3079);
nand U5989 (N_5989,N_4219,N_4516);
and U5990 (N_5990,N_4489,N_4605);
or U5991 (N_5991,N_2506,N_4610);
and U5992 (N_5992,N_3447,N_3067);
and U5993 (N_5993,N_3916,N_2900);
or U5994 (N_5994,N_2862,N_3622);
or U5995 (N_5995,N_2926,N_2898);
nand U5996 (N_5996,N_3489,N_4122);
or U5997 (N_5997,N_4169,N_2941);
nor U5998 (N_5998,N_3120,N_2765);
nand U5999 (N_5999,N_3981,N_4344);
and U6000 (N_6000,N_3938,N_3763);
nor U6001 (N_6001,N_4976,N_4375);
nand U6002 (N_6002,N_3274,N_4179);
nand U6003 (N_6003,N_4760,N_3760);
nand U6004 (N_6004,N_4282,N_4593);
and U6005 (N_6005,N_4191,N_4873);
and U6006 (N_6006,N_3360,N_3459);
nor U6007 (N_6007,N_3864,N_3893);
nand U6008 (N_6008,N_4779,N_3334);
nor U6009 (N_6009,N_2623,N_2796);
or U6010 (N_6010,N_2748,N_4263);
nor U6011 (N_6011,N_4060,N_2690);
and U6012 (N_6012,N_4715,N_2977);
and U6013 (N_6013,N_3299,N_3723);
and U6014 (N_6014,N_2551,N_4148);
nand U6015 (N_6015,N_3319,N_3454);
or U6016 (N_6016,N_2657,N_3575);
and U6017 (N_6017,N_4924,N_2852);
and U6018 (N_6018,N_4529,N_3133);
or U6019 (N_6019,N_4897,N_3041);
and U6020 (N_6020,N_3304,N_4079);
nor U6021 (N_6021,N_4583,N_4051);
xor U6022 (N_6022,N_3791,N_4498);
nand U6023 (N_6023,N_3789,N_3654);
and U6024 (N_6024,N_2851,N_3025);
or U6025 (N_6025,N_3434,N_4074);
nor U6026 (N_6026,N_4831,N_3991);
nor U6027 (N_6027,N_2779,N_3777);
nand U6028 (N_6028,N_4369,N_3231);
nand U6029 (N_6029,N_4846,N_3288);
nor U6030 (N_6030,N_3551,N_4484);
or U6031 (N_6031,N_2946,N_4046);
or U6032 (N_6032,N_3514,N_2782);
nand U6033 (N_6033,N_3497,N_3580);
nor U6034 (N_6034,N_3154,N_4677);
or U6035 (N_6035,N_4743,N_2682);
nand U6036 (N_6036,N_3190,N_3210);
or U6037 (N_6037,N_3435,N_4222);
nand U6038 (N_6038,N_3162,N_3774);
nor U6039 (N_6039,N_4332,N_3917);
or U6040 (N_6040,N_4176,N_3085);
nand U6041 (N_6041,N_3060,N_4759);
nand U6042 (N_6042,N_3651,N_3689);
nand U6043 (N_6043,N_2576,N_2614);
nor U6044 (N_6044,N_3885,N_4164);
nor U6045 (N_6045,N_3471,N_2872);
nand U6046 (N_6046,N_4988,N_4040);
or U6047 (N_6047,N_3252,N_4011);
or U6048 (N_6048,N_2627,N_4720);
nor U6049 (N_6049,N_4123,N_4626);
nand U6050 (N_6050,N_3092,N_2567);
or U6051 (N_6051,N_3153,N_4972);
or U6052 (N_6052,N_2671,N_4798);
and U6053 (N_6053,N_4731,N_4595);
or U6054 (N_6054,N_4888,N_4170);
nand U6055 (N_6055,N_3146,N_4881);
nor U6056 (N_6056,N_3398,N_2602);
nor U6057 (N_6057,N_3968,N_4525);
and U6058 (N_6058,N_4272,N_4778);
nor U6059 (N_6059,N_4919,N_4268);
or U6060 (N_6060,N_2784,N_3576);
or U6061 (N_6061,N_3416,N_3141);
and U6062 (N_6062,N_3627,N_2797);
nand U6063 (N_6063,N_3253,N_4203);
or U6064 (N_6064,N_3852,N_4511);
and U6065 (N_6065,N_4964,N_3862);
or U6066 (N_6066,N_3233,N_4151);
nand U6067 (N_6067,N_2786,N_4444);
nor U6068 (N_6068,N_3225,N_4230);
nand U6069 (N_6069,N_2812,N_4076);
xnor U6070 (N_6070,N_4478,N_4408);
and U6071 (N_6071,N_4974,N_3906);
nand U6072 (N_6072,N_4649,N_3974);
nand U6073 (N_6073,N_4863,N_3913);
nor U6074 (N_6074,N_2953,N_3517);
nand U6075 (N_6075,N_4250,N_4017);
and U6076 (N_6076,N_3011,N_4977);
nor U6077 (N_6077,N_3839,N_3099);
nor U6078 (N_6078,N_2659,N_3577);
xnor U6079 (N_6079,N_3014,N_3381);
nand U6080 (N_6080,N_4536,N_2832);
or U6081 (N_6081,N_3823,N_2871);
or U6082 (N_6082,N_3203,N_3595);
nor U6083 (N_6083,N_2583,N_4904);
nand U6084 (N_6084,N_3037,N_4255);
or U6085 (N_6085,N_4186,N_3652);
or U6086 (N_6086,N_2708,N_4647);
and U6087 (N_6087,N_4211,N_3110);
or U6088 (N_6088,N_3368,N_2918);
and U6089 (N_6089,N_2544,N_4377);
nand U6090 (N_6090,N_2580,N_3467);
nor U6091 (N_6091,N_3549,N_4923);
xnor U6092 (N_6092,N_2681,N_3899);
and U6093 (N_6093,N_4962,N_3601);
or U6094 (N_6094,N_3766,N_4446);
nand U6095 (N_6095,N_4641,N_3732);
or U6096 (N_6096,N_4108,N_3752);
nor U6097 (N_6097,N_4389,N_3324);
or U6098 (N_6098,N_2727,N_4264);
nor U6099 (N_6099,N_4596,N_3717);
nor U6100 (N_6100,N_3936,N_3344);
nand U6101 (N_6101,N_3861,N_3362);
nand U6102 (N_6102,N_2722,N_3787);
nor U6103 (N_6103,N_4660,N_3403);
nor U6104 (N_6104,N_3626,N_2874);
nor U6105 (N_6105,N_3900,N_2763);
or U6106 (N_6106,N_4920,N_3499);
and U6107 (N_6107,N_4541,N_3853);
and U6108 (N_6108,N_3664,N_3657);
nor U6109 (N_6109,N_4198,N_2747);
nand U6110 (N_6110,N_4938,N_3660);
nor U6111 (N_6111,N_2789,N_2975);
nand U6112 (N_6112,N_3584,N_2965);
and U6113 (N_6113,N_4261,N_4533);
nand U6114 (N_6114,N_3142,N_3254);
and U6115 (N_6115,N_4118,N_3429);
and U6116 (N_6116,N_3905,N_2545);
nand U6117 (N_6117,N_2629,N_3284);
or U6118 (N_6118,N_4090,N_2955);
nor U6119 (N_6119,N_2947,N_3662);
nand U6120 (N_6120,N_2724,N_2542);
nand U6121 (N_6121,N_2658,N_3890);
nor U6122 (N_6122,N_4064,N_3314);
or U6123 (N_6123,N_3186,N_4073);
nand U6124 (N_6124,N_4259,N_3877);
nor U6125 (N_6125,N_4413,N_3617);
and U6126 (N_6126,N_2820,N_4354);
and U6127 (N_6127,N_3138,N_4619);
nand U6128 (N_6128,N_2840,N_3581);
or U6129 (N_6129,N_2912,N_3701);
or U6130 (N_6130,N_4346,N_4984);
and U6131 (N_6131,N_3819,N_3640);
nor U6132 (N_6132,N_3390,N_3050);
nand U6133 (N_6133,N_3147,N_2899);
and U6134 (N_6134,N_3310,N_4871);
and U6135 (N_6135,N_4895,N_2650);
or U6136 (N_6136,N_2632,N_2959);
nand U6137 (N_6137,N_4249,N_4915);
or U6138 (N_6138,N_4676,N_3610);
nor U6139 (N_6139,N_3559,N_3705);
xor U6140 (N_6140,N_3907,N_3089);
nand U6141 (N_6141,N_3322,N_4445);
nor U6142 (N_6142,N_3608,N_3970);
nor U6143 (N_6143,N_4196,N_3928);
and U6144 (N_6144,N_4175,N_3510);
nand U6145 (N_6145,N_2744,N_2725);
nor U6146 (N_6146,N_4337,N_4197);
or U6147 (N_6147,N_4751,N_4842);
or U6148 (N_6148,N_3389,N_2711);
nand U6149 (N_6149,N_4811,N_4078);
nor U6150 (N_6150,N_4992,N_4804);
and U6151 (N_6151,N_3364,N_2528);
nor U6152 (N_6152,N_2869,N_3912);
nand U6153 (N_6153,N_3863,N_3361);
and U6154 (N_6154,N_3367,N_4348);
nand U6155 (N_6155,N_4104,N_2560);
nand U6156 (N_6156,N_4019,N_3540);
nor U6157 (N_6157,N_3420,N_4041);
and U6158 (N_6158,N_4805,N_4934);
nand U6159 (N_6159,N_3425,N_4828);
nand U6160 (N_6160,N_2795,N_3121);
nor U6161 (N_6161,N_4833,N_4537);
nor U6162 (N_6162,N_2512,N_3881);
and U6163 (N_6163,N_4514,N_4174);
nor U6164 (N_6164,N_4859,N_4062);
or U6165 (N_6165,N_3726,N_2933);
or U6166 (N_6166,N_3606,N_3267);
nand U6167 (N_6167,N_3531,N_4181);
nand U6168 (N_6168,N_2982,N_3034);
or U6169 (N_6169,N_3084,N_2798);
nand U6170 (N_6170,N_4577,N_4568);
nand U6171 (N_6171,N_2527,N_3137);
nand U6172 (N_6172,N_4764,N_2877);
or U6173 (N_6173,N_2984,N_4955);
or U6174 (N_6174,N_4518,N_4927);
nand U6175 (N_6175,N_3407,N_3438);
nor U6176 (N_6176,N_3124,N_3298);
or U6177 (N_6177,N_3166,N_3985);
nor U6178 (N_6178,N_3048,N_3311);
and U6179 (N_6179,N_4689,N_4447);
nor U6180 (N_6180,N_2759,N_2937);
and U6181 (N_6181,N_3964,N_4251);
nand U6182 (N_6182,N_4092,N_2719);
nor U6183 (N_6183,N_2773,N_4908);
nor U6184 (N_6184,N_4967,N_4376);
and U6185 (N_6185,N_4602,N_2611);
or U6186 (N_6186,N_4531,N_3442);
or U6187 (N_6187,N_4402,N_3748);
and U6188 (N_6188,N_4200,N_3127);
nor U6189 (N_6189,N_2691,N_2739);
nor U6190 (N_6190,N_2876,N_3681);
and U6191 (N_6191,N_4142,N_4558);
or U6192 (N_6192,N_2753,N_4466);
nand U6193 (N_6193,N_3104,N_3188);
nor U6194 (N_6194,N_3771,N_2637);
nor U6195 (N_6195,N_4269,N_2558);
nor U6196 (N_6196,N_2600,N_4067);
nor U6197 (N_6197,N_3378,N_4183);
and U6198 (N_6198,N_3070,N_4469);
or U6199 (N_6199,N_3630,N_3868);
or U6200 (N_6200,N_4057,N_2642);
and U6201 (N_6201,N_2510,N_2750);
nor U6202 (N_6202,N_4455,N_2702);
nor U6203 (N_6203,N_3357,N_2885);
nand U6204 (N_6204,N_4432,N_3096);
and U6205 (N_6205,N_4519,N_2809);
and U6206 (N_6206,N_3795,N_2577);
nor U6207 (N_6207,N_2780,N_3380);
nand U6208 (N_6208,N_2703,N_3865);
nand U6209 (N_6209,N_3061,N_3464);
nor U6210 (N_6210,N_4772,N_4884);
or U6211 (N_6211,N_4790,N_3482);
nand U6212 (N_6212,N_4971,N_4928);
or U6213 (N_6213,N_4405,N_3742);
and U6214 (N_6214,N_3157,N_4193);
nand U6215 (N_6215,N_2530,N_3097);
nor U6216 (N_6216,N_3148,N_3710);
nand U6217 (N_6217,N_3535,N_4359);
nor U6218 (N_6218,N_3191,N_4680);
and U6219 (N_6219,N_3691,N_3301);
or U6220 (N_6220,N_4816,N_3961);
and U6221 (N_6221,N_4265,N_3620);
nand U6222 (N_6222,N_3044,N_3776);
nor U6223 (N_6223,N_4061,N_3591);
nand U6224 (N_6224,N_2760,N_2967);
nand U6225 (N_6225,N_4808,N_2514);
nand U6226 (N_6226,N_3737,N_2963);
and U6227 (N_6227,N_4147,N_2638);
or U6228 (N_6228,N_3103,N_3518);
nor U6229 (N_6229,N_3285,N_2705);
nor U6230 (N_6230,N_4973,N_3615);
or U6231 (N_6231,N_4071,N_2564);
or U6232 (N_6232,N_4878,N_3553);
and U6233 (N_6233,N_3331,N_4116);
or U6234 (N_6234,N_4572,N_4330);
nor U6235 (N_6235,N_3102,N_3896);
or U6236 (N_6236,N_4094,N_2736);
or U6237 (N_6237,N_4713,N_2981);
or U6238 (N_6238,N_3982,N_4217);
and U6239 (N_6239,N_2555,N_3424);
or U6240 (N_6240,N_3684,N_2757);
and U6241 (N_6241,N_3728,N_4254);
nor U6242 (N_6242,N_2712,N_4417);
and U6243 (N_6243,N_4762,N_4087);
or U6244 (N_6244,N_3904,N_2831);
and U6245 (N_6245,N_4009,N_4728);
and U6246 (N_6246,N_2628,N_3292);
and U6247 (N_6247,N_3290,N_2587);
nand U6248 (N_6248,N_3294,N_2672);
nand U6249 (N_6249,N_4942,N_4499);
and U6250 (N_6250,N_3671,N_4447);
nor U6251 (N_6251,N_4602,N_4085);
or U6252 (N_6252,N_3566,N_4872);
nor U6253 (N_6253,N_3733,N_2721);
and U6254 (N_6254,N_4852,N_4174);
nor U6255 (N_6255,N_3662,N_2531);
nor U6256 (N_6256,N_3639,N_3322);
nand U6257 (N_6257,N_4661,N_4186);
or U6258 (N_6258,N_4679,N_3476);
nor U6259 (N_6259,N_4656,N_2564);
or U6260 (N_6260,N_2519,N_2648);
and U6261 (N_6261,N_3250,N_3678);
nor U6262 (N_6262,N_4245,N_3625);
and U6263 (N_6263,N_4793,N_3212);
nand U6264 (N_6264,N_3251,N_3548);
or U6265 (N_6265,N_3556,N_3944);
or U6266 (N_6266,N_3588,N_2533);
or U6267 (N_6267,N_2728,N_4535);
and U6268 (N_6268,N_4014,N_2754);
or U6269 (N_6269,N_4798,N_4907);
nand U6270 (N_6270,N_2928,N_3792);
and U6271 (N_6271,N_3742,N_4144);
or U6272 (N_6272,N_4935,N_4747);
nand U6273 (N_6273,N_2971,N_3800);
and U6274 (N_6274,N_4930,N_3506);
nand U6275 (N_6275,N_2626,N_4759);
nand U6276 (N_6276,N_2939,N_3766);
nand U6277 (N_6277,N_3758,N_3246);
or U6278 (N_6278,N_3846,N_4667);
or U6279 (N_6279,N_3627,N_4202);
or U6280 (N_6280,N_3651,N_3980);
or U6281 (N_6281,N_2698,N_3441);
nor U6282 (N_6282,N_2866,N_2788);
nand U6283 (N_6283,N_3753,N_3591);
nor U6284 (N_6284,N_3131,N_4163);
or U6285 (N_6285,N_3013,N_3806);
and U6286 (N_6286,N_4940,N_3189);
and U6287 (N_6287,N_4552,N_3567);
or U6288 (N_6288,N_2679,N_4958);
nor U6289 (N_6289,N_2790,N_4411);
xor U6290 (N_6290,N_4266,N_4377);
nand U6291 (N_6291,N_3107,N_3518);
or U6292 (N_6292,N_2539,N_2761);
nor U6293 (N_6293,N_2599,N_3389);
nor U6294 (N_6294,N_2997,N_3306);
or U6295 (N_6295,N_3476,N_4456);
or U6296 (N_6296,N_4759,N_2871);
nor U6297 (N_6297,N_4451,N_3249);
nand U6298 (N_6298,N_4995,N_3869);
and U6299 (N_6299,N_2816,N_3468);
and U6300 (N_6300,N_3836,N_4713);
nor U6301 (N_6301,N_4568,N_2563);
nor U6302 (N_6302,N_4951,N_4735);
nand U6303 (N_6303,N_4230,N_3261);
nand U6304 (N_6304,N_4150,N_3297);
nand U6305 (N_6305,N_3378,N_4920);
and U6306 (N_6306,N_4875,N_4329);
or U6307 (N_6307,N_2533,N_4928);
nor U6308 (N_6308,N_3866,N_3815);
or U6309 (N_6309,N_4981,N_4216);
nor U6310 (N_6310,N_2561,N_4798);
nor U6311 (N_6311,N_2980,N_2818);
or U6312 (N_6312,N_2920,N_4268);
and U6313 (N_6313,N_4941,N_4432);
nand U6314 (N_6314,N_3195,N_4774);
nand U6315 (N_6315,N_2804,N_3454);
nand U6316 (N_6316,N_2991,N_3310);
and U6317 (N_6317,N_3031,N_3484);
nand U6318 (N_6318,N_3500,N_3280);
nor U6319 (N_6319,N_3862,N_4304);
nand U6320 (N_6320,N_4041,N_2904);
or U6321 (N_6321,N_4964,N_4523);
nor U6322 (N_6322,N_3681,N_2652);
and U6323 (N_6323,N_3870,N_3528);
or U6324 (N_6324,N_3936,N_4181);
nand U6325 (N_6325,N_2677,N_4602);
or U6326 (N_6326,N_2695,N_3890);
and U6327 (N_6327,N_2565,N_4987);
or U6328 (N_6328,N_3875,N_4133);
or U6329 (N_6329,N_3675,N_3388);
or U6330 (N_6330,N_2664,N_3201);
or U6331 (N_6331,N_4160,N_2701);
or U6332 (N_6332,N_2683,N_4899);
nand U6333 (N_6333,N_4181,N_2781);
nor U6334 (N_6334,N_3307,N_3916);
nand U6335 (N_6335,N_3206,N_3953);
or U6336 (N_6336,N_4735,N_4595);
nor U6337 (N_6337,N_4827,N_3379);
and U6338 (N_6338,N_2636,N_3347);
nand U6339 (N_6339,N_3619,N_4632);
nand U6340 (N_6340,N_3963,N_4737);
or U6341 (N_6341,N_4299,N_3078);
and U6342 (N_6342,N_4148,N_3018);
nor U6343 (N_6343,N_3484,N_3215);
and U6344 (N_6344,N_3191,N_3019);
and U6345 (N_6345,N_3637,N_4348);
xor U6346 (N_6346,N_3370,N_3214);
or U6347 (N_6347,N_3623,N_4317);
nand U6348 (N_6348,N_4683,N_3051);
nand U6349 (N_6349,N_4501,N_2910);
xor U6350 (N_6350,N_4403,N_3842);
and U6351 (N_6351,N_4295,N_2852);
nor U6352 (N_6352,N_2683,N_3229);
or U6353 (N_6353,N_3495,N_3391);
and U6354 (N_6354,N_4062,N_4951);
or U6355 (N_6355,N_3482,N_3848);
nand U6356 (N_6356,N_2714,N_4588);
and U6357 (N_6357,N_3018,N_4276);
nor U6358 (N_6358,N_3026,N_4618);
nand U6359 (N_6359,N_3814,N_4615);
or U6360 (N_6360,N_4859,N_3495);
nor U6361 (N_6361,N_3067,N_3844);
and U6362 (N_6362,N_4168,N_2626);
nand U6363 (N_6363,N_4871,N_3678);
or U6364 (N_6364,N_3799,N_4624);
or U6365 (N_6365,N_3812,N_2700);
nor U6366 (N_6366,N_3100,N_3156);
nand U6367 (N_6367,N_4830,N_4229);
and U6368 (N_6368,N_3474,N_4751);
nand U6369 (N_6369,N_3999,N_4929);
nand U6370 (N_6370,N_3703,N_3590);
and U6371 (N_6371,N_4626,N_3029);
nor U6372 (N_6372,N_3878,N_4674);
and U6373 (N_6373,N_4936,N_4731);
or U6374 (N_6374,N_3465,N_3686);
nand U6375 (N_6375,N_2915,N_2820);
nor U6376 (N_6376,N_3133,N_3763);
nor U6377 (N_6377,N_3673,N_2640);
nand U6378 (N_6378,N_3122,N_3701);
or U6379 (N_6379,N_3649,N_4399);
nor U6380 (N_6380,N_2612,N_3950);
nor U6381 (N_6381,N_3621,N_4450);
nand U6382 (N_6382,N_3801,N_3891);
or U6383 (N_6383,N_2785,N_4978);
nand U6384 (N_6384,N_3589,N_3444);
or U6385 (N_6385,N_3436,N_4838);
and U6386 (N_6386,N_2654,N_3829);
nand U6387 (N_6387,N_4101,N_4904);
or U6388 (N_6388,N_3792,N_3445);
nand U6389 (N_6389,N_3889,N_4633);
or U6390 (N_6390,N_2971,N_4122);
nand U6391 (N_6391,N_4470,N_4861);
nand U6392 (N_6392,N_3236,N_3000);
and U6393 (N_6393,N_4169,N_3750);
or U6394 (N_6394,N_4854,N_4094);
and U6395 (N_6395,N_3934,N_4078);
and U6396 (N_6396,N_2654,N_4762);
nor U6397 (N_6397,N_4169,N_4491);
xor U6398 (N_6398,N_3566,N_3267);
and U6399 (N_6399,N_3725,N_3376);
and U6400 (N_6400,N_4505,N_3382);
nand U6401 (N_6401,N_3365,N_3851);
or U6402 (N_6402,N_4056,N_3802);
and U6403 (N_6403,N_3207,N_4466);
and U6404 (N_6404,N_3009,N_2631);
nor U6405 (N_6405,N_4265,N_2578);
and U6406 (N_6406,N_4403,N_3490);
xnor U6407 (N_6407,N_4163,N_4668);
nand U6408 (N_6408,N_4055,N_4365);
or U6409 (N_6409,N_4591,N_2917);
and U6410 (N_6410,N_3231,N_2687);
and U6411 (N_6411,N_4205,N_2636);
nand U6412 (N_6412,N_3056,N_4979);
nor U6413 (N_6413,N_4713,N_4155);
nor U6414 (N_6414,N_2518,N_4409);
or U6415 (N_6415,N_3359,N_4265);
and U6416 (N_6416,N_3429,N_3276);
and U6417 (N_6417,N_4748,N_4710);
nor U6418 (N_6418,N_3437,N_4002);
nor U6419 (N_6419,N_4800,N_4834);
or U6420 (N_6420,N_3495,N_2847);
or U6421 (N_6421,N_3535,N_4951);
or U6422 (N_6422,N_4498,N_4276);
and U6423 (N_6423,N_2810,N_3846);
or U6424 (N_6424,N_3663,N_4770);
or U6425 (N_6425,N_4399,N_3112);
nand U6426 (N_6426,N_3788,N_4613);
and U6427 (N_6427,N_4876,N_2850);
xnor U6428 (N_6428,N_3831,N_3392);
or U6429 (N_6429,N_2813,N_4921);
nor U6430 (N_6430,N_4060,N_3179);
nor U6431 (N_6431,N_4089,N_4674);
or U6432 (N_6432,N_4445,N_3909);
and U6433 (N_6433,N_4271,N_3614);
or U6434 (N_6434,N_3541,N_3577);
or U6435 (N_6435,N_4649,N_4095);
nand U6436 (N_6436,N_2638,N_4369);
and U6437 (N_6437,N_2874,N_3097);
nor U6438 (N_6438,N_3123,N_4126);
or U6439 (N_6439,N_3902,N_4979);
or U6440 (N_6440,N_4510,N_3618);
and U6441 (N_6441,N_2936,N_4526);
nand U6442 (N_6442,N_2782,N_4445);
and U6443 (N_6443,N_3645,N_3516);
and U6444 (N_6444,N_2712,N_4902);
or U6445 (N_6445,N_4271,N_3901);
nor U6446 (N_6446,N_3504,N_3979);
nand U6447 (N_6447,N_3734,N_3996);
nand U6448 (N_6448,N_3113,N_2969);
nand U6449 (N_6449,N_4340,N_3311);
nor U6450 (N_6450,N_3568,N_3546);
nand U6451 (N_6451,N_2508,N_4694);
nand U6452 (N_6452,N_3147,N_4564);
nand U6453 (N_6453,N_2538,N_3665);
nand U6454 (N_6454,N_3323,N_4377);
nand U6455 (N_6455,N_4270,N_2795);
nand U6456 (N_6456,N_3940,N_3350);
and U6457 (N_6457,N_3856,N_4149);
nor U6458 (N_6458,N_4517,N_3927);
xor U6459 (N_6459,N_3687,N_3071);
xor U6460 (N_6460,N_2592,N_3869);
nor U6461 (N_6461,N_4227,N_3091);
or U6462 (N_6462,N_4453,N_3277);
xor U6463 (N_6463,N_4903,N_4341);
nand U6464 (N_6464,N_3300,N_3401);
nand U6465 (N_6465,N_2528,N_4625);
nand U6466 (N_6466,N_4345,N_3076);
nor U6467 (N_6467,N_3745,N_4116);
or U6468 (N_6468,N_4009,N_2576);
nor U6469 (N_6469,N_3275,N_4140);
or U6470 (N_6470,N_2722,N_2639);
nand U6471 (N_6471,N_3821,N_4199);
or U6472 (N_6472,N_3363,N_4120);
nand U6473 (N_6473,N_3617,N_4792);
and U6474 (N_6474,N_4396,N_2528);
and U6475 (N_6475,N_4763,N_4769);
nand U6476 (N_6476,N_3631,N_3938);
nand U6477 (N_6477,N_3248,N_4641);
or U6478 (N_6478,N_4711,N_3663);
nand U6479 (N_6479,N_4236,N_3815);
nand U6480 (N_6480,N_3303,N_4498);
and U6481 (N_6481,N_2971,N_4727);
or U6482 (N_6482,N_3998,N_3844);
or U6483 (N_6483,N_2599,N_3586);
nand U6484 (N_6484,N_3161,N_4060);
and U6485 (N_6485,N_2754,N_4488);
and U6486 (N_6486,N_3789,N_4050);
nand U6487 (N_6487,N_4317,N_3227);
and U6488 (N_6488,N_4908,N_4942);
or U6489 (N_6489,N_4933,N_2536);
and U6490 (N_6490,N_4064,N_3351);
nand U6491 (N_6491,N_3336,N_4632);
or U6492 (N_6492,N_2738,N_3695);
nand U6493 (N_6493,N_2628,N_3780);
or U6494 (N_6494,N_4410,N_4830);
nor U6495 (N_6495,N_4282,N_4118);
nor U6496 (N_6496,N_2701,N_4241);
and U6497 (N_6497,N_4755,N_4305);
or U6498 (N_6498,N_2697,N_2715);
nand U6499 (N_6499,N_3630,N_3260);
and U6500 (N_6500,N_4684,N_3325);
and U6501 (N_6501,N_3274,N_4846);
nand U6502 (N_6502,N_4371,N_3089);
and U6503 (N_6503,N_2993,N_2924);
or U6504 (N_6504,N_4441,N_2624);
nand U6505 (N_6505,N_4358,N_4150);
xnor U6506 (N_6506,N_3329,N_3030);
nor U6507 (N_6507,N_2779,N_3009);
nor U6508 (N_6508,N_4514,N_2618);
and U6509 (N_6509,N_3835,N_2839);
or U6510 (N_6510,N_3477,N_3609);
nand U6511 (N_6511,N_3320,N_3907);
nor U6512 (N_6512,N_3211,N_4958);
or U6513 (N_6513,N_2610,N_4586);
or U6514 (N_6514,N_4865,N_2510);
nand U6515 (N_6515,N_4826,N_3213);
nor U6516 (N_6516,N_2766,N_2791);
nand U6517 (N_6517,N_4580,N_4030);
or U6518 (N_6518,N_4819,N_2922);
nand U6519 (N_6519,N_3183,N_4413);
nor U6520 (N_6520,N_4568,N_3284);
nand U6521 (N_6521,N_2903,N_3406);
nand U6522 (N_6522,N_4089,N_3724);
or U6523 (N_6523,N_2543,N_2780);
nand U6524 (N_6524,N_4639,N_3238);
and U6525 (N_6525,N_4335,N_4353);
and U6526 (N_6526,N_2741,N_4911);
or U6527 (N_6527,N_4733,N_2825);
nand U6528 (N_6528,N_3910,N_3442);
or U6529 (N_6529,N_4524,N_3304);
nor U6530 (N_6530,N_4681,N_3118);
or U6531 (N_6531,N_4975,N_3336);
nand U6532 (N_6532,N_4889,N_3893);
nand U6533 (N_6533,N_3537,N_4135);
nand U6534 (N_6534,N_4189,N_3871);
and U6535 (N_6535,N_2880,N_3167);
nand U6536 (N_6536,N_2921,N_4916);
and U6537 (N_6537,N_3500,N_3586);
nand U6538 (N_6538,N_2856,N_3194);
xor U6539 (N_6539,N_4281,N_3285);
or U6540 (N_6540,N_4605,N_4442);
nor U6541 (N_6541,N_3376,N_2709);
and U6542 (N_6542,N_3659,N_3660);
nand U6543 (N_6543,N_3206,N_4879);
nor U6544 (N_6544,N_4912,N_3711);
and U6545 (N_6545,N_4073,N_2534);
or U6546 (N_6546,N_3295,N_4284);
nor U6547 (N_6547,N_2745,N_4035);
nand U6548 (N_6548,N_3990,N_2985);
nor U6549 (N_6549,N_4674,N_3183);
nor U6550 (N_6550,N_3893,N_4710);
nor U6551 (N_6551,N_4716,N_4465);
or U6552 (N_6552,N_4105,N_3811);
or U6553 (N_6553,N_3411,N_4706);
nor U6554 (N_6554,N_4173,N_2572);
nor U6555 (N_6555,N_2517,N_4766);
nand U6556 (N_6556,N_4855,N_4717);
nor U6557 (N_6557,N_4183,N_3517);
and U6558 (N_6558,N_4082,N_4349);
nor U6559 (N_6559,N_3651,N_2560);
and U6560 (N_6560,N_2566,N_4288);
and U6561 (N_6561,N_2858,N_2962);
or U6562 (N_6562,N_4739,N_3141);
nand U6563 (N_6563,N_4947,N_3153);
or U6564 (N_6564,N_2779,N_2529);
nand U6565 (N_6565,N_3167,N_2801);
nand U6566 (N_6566,N_4653,N_3773);
nor U6567 (N_6567,N_4307,N_4377);
nand U6568 (N_6568,N_4823,N_2859);
nand U6569 (N_6569,N_4027,N_4197);
nor U6570 (N_6570,N_4320,N_2701);
nand U6571 (N_6571,N_3774,N_2502);
nand U6572 (N_6572,N_3542,N_3500);
or U6573 (N_6573,N_4721,N_2528);
nor U6574 (N_6574,N_3610,N_4996);
or U6575 (N_6575,N_4538,N_4136);
nand U6576 (N_6576,N_4086,N_3221);
nand U6577 (N_6577,N_3036,N_3469);
nor U6578 (N_6578,N_4036,N_3072);
or U6579 (N_6579,N_4625,N_2871);
or U6580 (N_6580,N_3361,N_3519);
nor U6581 (N_6581,N_3828,N_2833);
nor U6582 (N_6582,N_3719,N_4541);
or U6583 (N_6583,N_4328,N_3032);
or U6584 (N_6584,N_3374,N_2550);
and U6585 (N_6585,N_2617,N_3446);
nor U6586 (N_6586,N_3281,N_3082);
or U6587 (N_6587,N_3489,N_2656);
and U6588 (N_6588,N_4638,N_3057);
and U6589 (N_6589,N_3651,N_4863);
nand U6590 (N_6590,N_2778,N_3687);
or U6591 (N_6591,N_3249,N_2721);
nand U6592 (N_6592,N_4415,N_4660);
and U6593 (N_6593,N_3731,N_3933);
nand U6594 (N_6594,N_3475,N_4101);
or U6595 (N_6595,N_3482,N_4649);
and U6596 (N_6596,N_3802,N_4982);
nand U6597 (N_6597,N_4961,N_4388);
nor U6598 (N_6598,N_4860,N_2581);
and U6599 (N_6599,N_4243,N_2872);
and U6600 (N_6600,N_4562,N_4208);
nor U6601 (N_6601,N_4336,N_3149);
nand U6602 (N_6602,N_3394,N_2589);
nor U6603 (N_6603,N_4343,N_4604);
nand U6604 (N_6604,N_3809,N_3608);
nor U6605 (N_6605,N_2509,N_3756);
nor U6606 (N_6606,N_4924,N_4160);
nor U6607 (N_6607,N_4614,N_3814);
nand U6608 (N_6608,N_3872,N_3504);
nand U6609 (N_6609,N_3494,N_3354);
nand U6610 (N_6610,N_4804,N_3793);
nand U6611 (N_6611,N_4611,N_3491);
and U6612 (N_6612,N_2725,N_4130);
nand U6613 (N_6613,N_3254,N_2777);
nand U6614 (N_6614,N_3332,N_2831);
nand U6615 (N_6615,N_4916,N_3859);
nor U6616 (N_6616,N_3323,N_3372);
or U6617 (N_6617,N_4882,N_3690);
or U6618 (N_6618,N_2700,N_4130);
and U6619 (N_6619,N_3553,N_4253);
or U6620 (N_6620,N_3414,N_2828);
or U6621 (N_6621,N_4878,N_3329);
nand U6622 (N_6622,N_3593,N_3470);
nand U6623 (N_6623,N_4635,N_3157);
or U6624 (N_6624,N_3397,N_3342);
and U6625 (N_6625,N_3349,N_4674);
and U6626 (N_6626,N_4736,N_3307);
nor U6627 (N_6627,N_3159,N_3284);
or U6628 (N_6628,N_3821,N_4689);
or U6629 (N_6629,N_3583,N_3382);
nand U6630 (N_6630,N_4746,N_3501);
and U6631 (N_6631,N_4953,N_2915);
or U6632 (N_6632,N_4782,N_4081);
nand U6633 (N_6633,N_3680,N_3268);
or U6634 (N_6634,N_3020,N_4438);
nand U6635 (N_6635,N_4422,N_4309);
nor U6636 (N_6636,N_4660,N_4011);
nor U6637 (N_6637,N_2518,N_4168);
and U6638 (N_6638,N_4553,N_4552);
nor U6639 (N_6639,N_3228,N_3966);
and U6640 (N_6640,N_4288,N_3853);
nor U6641 (N_6641,N_4406,N_4720);
nor U6642 (N_6642,N_3726,N_3491);
and U6643 (N_6643,N_3036,N_3339);
or U6644 (N_6644,N_4611,N_4232);
nor U6645 (N_6645,N_3447,N_3500);
nor U6646 (N_6646,N_3028,N_3692);
nand U6647 (N_6647,N_4780,N_3134);
and U6648 (N_6648,N_3027,N_2633);
or U6649 (N_6649,N_3701,N_3903);
and U6650 (N_6650,N_2791,N_3392);
xor U6651 (N_6651,N_4972,N_2612);
nor U6652 (N_6652,N_4327,N_3423);
nor U6653 (N_6653,N_3402,N_3569);
nor U6654 (N_6654,N_3417,N_2541);
nor U6655 (N_6655,N_4292,N_2968);
or U6656 (N_6656,N_4092,N_4627);
or U6657 (N_6657,N_3143,N_3278);
nor U6658 (N_6658,N_2954,N_2862);
or U6659 (N_6659,N_3917,N_4866);
nor U6660 (N_6660,N_3661,N_4610);
nand U6661 (N_6661,N_3307,N_4586);
or U6662 (N_6662,N_3156,N_3051);
or U6663 (N_6663,N_2886,N_2673);
nor U6664 (N_6664,N_2986,N_3498);
and U6665 (N_6665,N_4663,N_3438);
and U6666 (N_6666,N_3646,N_3210);
or U6667 (N_6667,N_4826,N_2703);
or U6668 (N_6668,N_3471,N_3439);
nor U6669 (N_6669,N_2769,N_4515);
nor U6670 (N_6670,N_4066,N_3498);
and U6671 (N_6671,N_3846,N_4977);
nor U6672 (N_6672,N_3760,N_3662);
nand U6673 (N_6673,N_2707,N_2618);
and U6674 (N_6674,N_3440,N_4014);
or U6675 (N_6675,N_3791,N_4750);
or U6676 (N_6676,N_3532,N_3837);
and U6677 (N_6677,N_4429,N_2667);
and U6678 (N_6678,N_4980,N_3098);
nor U6679 (N_6679,N_4732,N_3374);
or U6680 (N_6680,N_3263,N_4118);
and U6681 (N_6681,N_2601,N_3409);
or U6682 (N_6682,N_4086,N_3953);
and U6683 (N_6683,N_4670,N_2860);
or U6684 (N_6684,N_4714,N_3664);
nor U6685 (N_6685,N_3974,N_4757);
or U6686 (N_6686,N_3404,N_3617);
and U6687 (N_6687,N_4561,N_2693);
nand U6688 (N_6688,N_3885,N_4991);
or U6689 (N_6689,N_4182,N_3922);
nor U6690 (N_6690,N_2652,N_4046);
nand U6691 (N_6691,N_2662,N_2843);
and U6692 (N_6692,N_4460,N_2706);
nand U6693 (N_6693,N_4666,N_4169);
nand U6694 (N_6694,N_3068,N_4011);
and U6695 (N_6695,N_4953,N_3060);
and U6696 (N_6696,N_4114,N_3267);
or U6697 (N_6697,N_4908,N_4383);
nand U6698 (N_6698,N_2551,N_3688);
nor U6699 (N_6699,N_4000,N_3282);
nor U6700 (N_6700,N_4247,N_3372);
nand U6701 (N_6701,N_3747,N_4581);
and U6702 (N_6702,N_4027,N_3007);
or U6703 (N_6703,N_3004,N_2639);
and U6704 (N_6704,N_3481,N_4732);
and U6705 (N_6705,N_3117,N_3550);
nor U6706 (N_6706,N_4251,N_3352);
nand U6707 (N_6707,N_3742,N_4194);
nand U6708 (N_6708,N_4175,N_3299);
and U6709 (N_6709,N_2599,N_3867);
nor U6710 (N_6710,N_4629,N_3407);
nor U6711 (N_6711,N_4627,N_4708);
nand U6712 (N_6712,N_4905,N_3337);
and U6713 (N_6713,N_3854,N_3613);
or U6714 (N_6714,N_3915,N_3720);
and U6715 (N_6715,N_3566,N_3729);
or U6716 (N_6716,N_4878,N_4477);
or U6717 (N_6717,N_3944,N_3687);
nor U6718 (N_6718,N_2855,N_4812);
nor U6719 (N_6719,N_4425,N_3953);
nor U6720 (N_6720,N_3134,N_3632);
nor U6721 (N_6721,N_4596,N_3373);
and U6722 (N_6722,N_3835,N_3761);
or U6723 (N_6723,N_2570,N_4127);
nand U6724 (N_6724,N_3768,N_3728);
nand U6725 (N_6725,N_4969,N_2899);
or U6726 (N_6726,N_4178,N_4159);
or U6727 (N_6727,N_3017,N_3946);
and U6728 (N_6728,N_3129,N_3290);
nor U6729 (N_6729,N_2704,N_3494);
nor U6730 (N_6730,N_4003,N_3217);
nor U6731 (N_6731,N_3144,N_4527);
xnor U6732 (N_6732,N_3935,N_4788);
nand U6733 (N_6733,N_3569,N_3259);
or U6734 (N_6734,N_3661,N_3677);
xor U6735 (N_6735,N_3346,N_3605);
or U6736 (N_6736,N_3206,N_3149);
nand U6737 (N_6737,N_4423,N_4113);
nor U6738 (N_6738,N_4456,N_4897);
nand U6739 (N_6739,N_4016,N_4716);
or U6740 (N_6740,N_4296,N_2766);
nand U6741 (N_6741,N_3641,N_4630);
or U6742 (N_6742,N_4470,N_4332);
and U6743 (N_6743,N_4658,N_4698);
nand U6744 (N_6744,N_2597,N_3156);
nand U6745 (N_6745,N_2687,N_3842);
and U6746 (N_6746,N_2850,N_4124);
nand U6747 (N_6747,N_4479,N_4838);
nor U6748 (N_6748,N_3341,N_2895);
or U6749 (N_6749,N_3975,N_4839);
nand U6750 (N_6750,N_4774,N_4918);
and U6751 (N_6751,N_2753,N_2915);
nand U6752 (N_6752,N_4728,N_3634);
and U6753 (N_6753,N_4136,N_4763);
nor U6754 (N_6754,N_3308,N_2932);
nand U6755 (N_6755,N_3837,N_3561);
and U6756 (N_6756,N_2536,N_4302);
and U6757 (N_6757,N_4496,N_3574);
nor U6758 (N_6758,N_4190,N_3397);
nand U6759 (N_6759,N_3462,N_3785);
nand U6760 (N_6760,N_3580,N_4404);
nor U6761 (N_6761,N_4825,N_2980);
nor U6762 (N_6762,N_3755,N_4866);
nand U6763 (N_6763,N_4667,N_4090);
nor U6764 (N_6764,N_4237,N_3930);
nand U6765 (N_6765,N_3853,N_3087);
nand U6766 (N_6766,N_2927,N_4366);
nand U6767 (N_6767,N_3087,N_3071);
nor U6768 (N_6768,N_4224,N_3056);
nand U6769 (N_6769,N_4613,N_2941);
nand U6770 (N_6770,N_4205,N_3244);
or U6771 (N_6771,N_4768,N_3110);
or U6772 (N_6772,N_3390,N_2513);
and U6773 (N_6773,N_4618,N_2837);
nand U6774 (N_6774,N_4212,N_3880);
and U6775 (N_6775,N_3498,N_3043);
or U6776 (N_6776,N_3266,N_3477);
or U6777 (N_6777,N_2601,N_3655);
and U6778 (N_6778,N_2712,N_2940);
nor U6779 (N_6779,N_4430,N_4617);
nor U6780 (N_6780,N_4239,N_3954);
and U6781 (N_6781,N_4665,N_3968);
and U6782 (N_6782,N_2914,N_4656);
and U6783 (N_6783,N_3770,N_3021);
nand U6784 (N_6784,N_3860,N_3516);
nor U6785 (N_6785,N_4560,N_3234);
and U6786 (N_6786,N_3601,N_3481);
nor U6787 (N_6787,N_4741,N_4568);
or U6788 (N_6788,N_4522,N_4912);
and U6789 (N_6789,N_2813,N_4599);
nor U6790 (N_6790,N_2909,N_3264);
nor U6791 (N_6791,N_3194,N_4066);
nand U6792 (N_6792,N_2572,N_4231);
or U6793 (N_6793,N_2866,N_2668);
nand U6794 (N_6794,N_2619,N_3888);
and U6795 (N_6795,N_4887,N_4821);
or U6796 (N_6796,N_3506,N_4471);
nor U6797 (N_6797,N_3856,N_3035);
and U6798 (N_6798,N_4260,N_3951);
nand U6799 (N_6799,N_3247,N_4322);
and U6800 (N_6800,N_3248,N_2547);
or U6801 (N_6801,N_3585,N_3507);
nor U6802 (N_6802,N_3612,N_3083);
or U6803 (N_6803,N_4334,N_4088);
nand U6804 (N_6804,N_3247,N_4898);
nor U6805 (N_6805,N_4718,N_4150);
or U6806 (N_6806,N_2921,N_4200);
nand U6807 (N_6807,N_3302,N_4641);
and U6808 (N_6808,N_2956,N_4460);
and U6809 (N_6809,N_4168,N_3597);
or U6810 (N_6810,N_4472,N_3938);
nand U6811 (N_6811,N_3270,N_4329);
nand U6812 (N_6812,N_3215,N_2779);
or U6813 (N_6813,N_2692,N_3095);
nand U6814 (N_6814,N_4699,N_4254);
or U6815 (N_6815,N_2966,N_4577);
or U6816 (N_6816,N_4066,N_2669);
or U6817 (N_6817,N_4103,N_2853);
nor U6818 (N_6818,N_4559,N_4330);
nor U6819 (N_6819,N_2772,N_3118);
or U6820 (N_6820,N_4761,N_3501);
and U6821 (N_6821,N_4041,N_2902);
and U6822 (N_6822,N_3882,N_3445);
nand U6823 (N_6823,N_2608,N_2797);
nand U6824 (N_6824,N_2931,N_3737);
nand U6825 (N_6825,N_4705,N_3021);
and U6826 (N_6826,N_4280,N_3146);
nand U6827 (N_6827,N_3009,N_4209);
and U6828 (N_6828,N_3581,N_3997);
or U6829 (N_6829,N_4765,N_4671);
nor U6830 (N_6830,N_4978,N_2999);
nor U6831 (N_6831,N_3945,N_4665);
nand U6832 (N_6832,N_3456,N_4246);
nor U6833 (N_6833,N_3332,N_4289);
nor U6834 (N_6834,N_4994,N_4818);
nand U6835 (N_6835,N_3547,N_3298);
or U6836 (N_6836,N_3427,N_4564);
or U6837 (N_6837,N_4546,N_4024);
or U6838 (N_6838,N_3790,N_3318);
nand U6839 (N_6839,N_3290,N_3840);
nor U6840 (N_6840,N_4879,N_4380);
nand U6841 (N_6841,N_2808,N_2738);
and U6842 (N_6842,N_3430,N_4603);
nor U6843 (N_6843,N_4344,N_3051);
nand U6844 (N_6844,N_2817,N_4785);
or U6845 (N_6845,N_4685,N_3447);
nand U6846 (N_6846,N_3658,N_3415);
or U6847 (N_6847,N_3800,N_3304);
or U6848 (N_6848,N_2600,N_3491);
nand U6849 (N_6849,N_4497,N_4605);
or U6850 (N_6850,N_3984,N_4071);
or U6851 (N_6851,N_2573,N_4098);
and U6852 (N_6852,N_4617,N_3126);
nand U6853 (N_6853,N_3964,N_3356);
or U6854 (N_6854,N_3199,N_2978);
or U6855 (N_6855,N_3360,N_2795);
and U6856 (N_6856,N_4829,N_4615);
xnor U6857 (N_6857,N_3091,N_4864);
and U6858 (N_6858,N_3193,N_4938);
nor U6859 (N_6859,N_2911,N_3091);
or U6860 (N_6860,N_4274,N_4255);
and U6861 (N_6861,N_4056,N_4754);
nor U6862 (N_6862,N_2817,N_4108);
nand U6863 (N_6863,N_4219,N_3093);
nand U6864 (N_6864,N_3474,N_4731);
nor U6865 (N_6865,N_3942,N_4235);
nand U6866 (N_6866,N_3569,N_4978);
and U6867 (N_6867,N_4801,N_3993);
nor U6868 (N_6868,N_4183,N_3583);
or U6869 (N_6869,N_2827,N_3415);
nor U6870 (N_6870,N_2858,N_3112);
nand U6871 (N_6871,N_3342,N_3791);
and U6872 (N_6872,N_3207,N_4509);
nand U6873 (N_6873,N_4249,N_4090);
nor U6874 (N_6874,N_3965,N_3719);
and U6875 (N_6875,N_2836,N_2749);
or U6876 (N_6876,N_3815,N_4001);
or U6877 (N_6877,N_4876,N_4259);
and U6878 (N_6878,N_3742,N_3078);
nand U6879 (N_6879,N_3256,N_4224);
nand U6880 (N_6880,N_4154,N_3577);
nor U6881 (N_6881,N_4530,N_2683);
or U6882 (N_6882,N_4193,N_4446);
or U6883 (N_6883,N_2702,N_2851);
and U6884 (N_6884,N_3697,N_3305);
and U6885 (N_6885,N_4744,N_3984);
nand U6886 (N_6886,N_2762,N_3553);
or U6887 (N_6887,N_3922,N_2889);
nor U6888 (N_6888,N_2755,N_4499);
or U6889 (N_6889,N_3970,N_3818);
and U6890 (N_6890,N_3370,N_4709);
nor U6891 (N_6891,N_3602,N_4789);
or U6892 (N_6892,N_3803,N_3744);
nor U6893 (N_6893,N_3544,N_3472);
nand U6894 (N_6894,N_4906,N_2938);
or U6895 (N_6895,N_2725,N_3687);
and U6896 (N_6896,N_3269,N_4739);
nand U6897 (N_6897,N_3787,N_4535);
nand U6898 (N_6898,N_2984,N_2753);
nor U6899 (N_6899,N_4264,N_4260);
nand U6900 (N_6900,N_4650,N_3778);
or U6901 (N_6901,N_3205,N_4987);
and U6902 (N_6902,N_3472,N_2771);
nand U6903 (N_6903,N_4489,N_3997);
xnor U6904 (N_6904,N_4608,N_4753);
nor U6905 (N_6905,N_2832,N_2578);
or U6906 (N_6906,N_3909,N_3261);
or U6907 (N_6907,N_4119,N_3163);
nand U6908 (N_6908,N_4377,N_4689);
nand U6909 (N_6909,N_3474,N_2879);
and U6910 (N_6910,N_3431,N_4976);
and U6911 (N_6911,N_4310,N_3793);
and U6912 (N_6912,N_3329,N_3261);
and U6913 (N_6913,N_3647,N_3889);
nand U6914 (N_6914,N_2566,N_3521);
nor U6915 (N_6915,N_4534,N_3875);
nor U6916 (N_6916,N_3566,N_4142);
nor U6917 (N_6917,N_4379,N_4179);
or U6918 (N_6918,N_3555,N_2990);
or U6919 (N_6919,N_3355,N_4818);
nor U6920 (N_6920,N_3328,N_3293);
and U6921 (N_6921,N_2582,N_2687);
and U6922 (N_6922,N_3114,N_2818);
and U6923 (N_6923,N_3632,N_3894);
nor U6924 (N_6924,N_3639,N_3061);
nand U6925 (N_6925,N_3646,N_2549);
or U6926 (N_6926,N_2689,N_3242);
nand U6927 (N_6927,N_3757,N_3852);
or U6928 (N_6928,N_3764,N_3273);
nand U6929 (N_6929,N_2717,N_3253);
and U6930 (N_6930,N_4367,N_4583);
and U6931 (N_6931,N_4134,N_3229);
or U6932 (N_6932,N_3231,N_3745);
xor U6933 (N_6933,N_2986,N_4416);
nand U6934 (N_6934,N_3948,N_4043);
or U6935 (N_6935,N_4555,N_3251);
nand U6936 (N_6936,N_3966,N_3057);
and U6937 (N_6937,N_3683,N_3714);
and U6938 (N_6938,N_3057,N_4101);
or U6939 (N_6939,N_2812,N_3794);
nand U6940 (N_6940,N_4562,N_2612);
nor U6941 (N_6941,N_4884,N_4845);
nor U6942 (N_6942,N_4651,N_4623);
nand U6943 (N_6943,N_3247,N_2569);
and U6944 (N_6944,N_4529,N_4385);
nand U6945 (N_6945,N_4571,N_3287);
nor U6946 (N_6946,N_2914,N_4378);
nand U6947 (N_6947,N_4750,N_3254);
nand U6948 (N_6948,N_3000,N_4754);
nor U6949 (N_6949,N_3859,N_3932);
nor U6950 (N_6950,N_3157,N_2655);
nor U6951 (N_6951,N_3639,N_3634);
nand U6952 (N_6952,N_2630,N_4798);
nor U6953 (N_6953,N_3490,N_3839);
nand U6954 (N_6954,N_3004,N_2844);
nand U6955 (N_6955,N_3064,N_4509);
and U6956 (N_6956,N_4178,N_4999);
nand U6957 (N_6957,N_3684,N_4184);
nand U6958 (N_6958,N_4106,N_4690);
nor U6959 (N_6959,N_3377,N_3246);
nand U6960 (N_6960,N_3826,N_3331);
nor U6961 (N_6961,N_3187,N_3488);
or U6962 (N_6962,N_3065,N_3751);
and U6963 (N_6963,N_4198,N_4072);
nand U6964 (N_6964,N_3046,N_3865);
and U6965 (N_6965,N_2832,N_4424);
nor U6966 (N_6966,N_2636,N_4796);
nand U6967 (N_6967,N_3461,N_4447);
nor U6968 (N_6968,N_4624,N_4472);
nand U6969 (N_6969,N_3665,N_4177);
or U6970 (N_6970,N_2564,N_4115);
nand U6971 (N_6971,N_3180,N_3246);
nand U6972 (N_6972,N_3717,N_3813);
and U6973 (N_6973,N_4471,N_4472);
or U6974 (N_6974,N_3741,N_4599);
and U6975 (N_6975,N_3260,N_4670);
and U6976 (N_6976,N_3150,N_3143);
and U6977 (N_6977,N_2836,N_3154);
nand U6978 (N_6978,N_4956,N_2868);
nand U6979 (N_6979,N_3569,N_3187);
nand U6980 (N_6980,N_3206,N_3359);
or U6981 (N_6981,N_4538,N_3978);
or U6982 (N_6982,N_4587,N_4469);
and U6983 (N_6983,N_3759,N_3307);
nor U6984 (N_6984,N_4558,N_3249);
nand U6985 (N_6985,N_3447,N_2734);
nor U6986 (N_6986,N_4134,N_3626);
or U6987 (N_6987,N_4379,N_3053);
or U6988 (N_6988,N_4043,N_2702);
nand U6989 (N_6989,N_3119,N_4167);
and U6990 (N_6990,N_3007,N_2753);
nand U6991 (N_6991,N_3535,N_4931);
or U6992 (N_6992,N_3364,N_3917);
and U6993 (N_6993,N_3490,N_3087);
nand U6994 (N_6994,N_4774,N_2948);
or U6995 (N_6995,N_3346,N_3187);
nor U6996 (N_6996,N_3655,N_3329);
or U6997 (N_6997,N_3344,N_3882);
and U6998 (N_6998,N_2874,N_3564);
or U6999 (N_6999,N_4966,N_2588);
and U7000 (N_7000,N_4685,N_2684);
and U7001 (N_7001,N_4138,N_3494);
nor U7002 (N_7002,N_4364,N_3806);
and U7003 (N_7003,N_4984,N_3062);
and U7004 (N_7004,N_4575,N_4671);
or U7005 (N_7005,N_3384,N_4548);
and U7006 (N_7006,N_4018,N_4934);
nand U7007 (N_7007,N_2766,N_4678);
nand U7008 (N_7008,N_4112,N_2778);
nor U7009 (N_7009,N_3677,N_4504);
or U7010 (N_7010,N_3446,N_3505);
nand U7011 (N_7011,N_3806,N_2919);
and U7012 (N_7012,N_4184,N_3774);
nand U7013 (N_7013,N_3764,N_4028);
nand U7014 (N_7014,N_2716,N_4453);
nand U7015 (N_7015,N_2721,N_3299);
nor U7016 (N_7016,N_3097,N_2787);
nor U7017 (N_7017,N_2694,N_2885);
or U7018 (N_7018,N_3130,N_3844);
and U7019 (N_7019,N_3720,N_2592);
nand U7020 (N_7020,N_2863,N_3424);
nand U7021 (N_7021,N_4292,N_3799);
and U7022 (N_7022,N_4139,N_3681);
nor U7023 (N_7023,N_4262,N_2993);
nor U7024 (N_7024,N_3973,N_4888);
and U7025 (N_7025,N_3274,N_4931);
nor U7026 (N_7026,N_4004,N_3437);
xor U7027 (N_7027,N_3211,N_2762);
or U7028 (N_7028,N_2899,N_2775);
nor U7029 (N_7029,N_3945,N_4579);
nand U7030 (N_7030,N_4266,N_2664);
nand U7031 (N_7031,N_3315,N_3679);
or U7032 (N_7032,N_2973,N_2814);
nor U7033 (N_7033,N_4127,N_2697);
nor U7034 (N_7034,N_4315,N_3801);
nand U7035 (N_7035,N_4977,N_2863);
nand U7036 (N_7036,N_4265,N_3236);
or U7037 (N_7037,N_4520,N_4953);
nor U7038 (N_7038,N_2940,N_3533);
nand U7039 (N_7039,N_4092,N_4463);
nand U7040 (N_7040,N_2590,N_2909);
nand U7041 (N_7041,N_4234,N_3203);
or U7042 (N_7042,N_2914,N_2622);
or U7043 (N_7043,N_3523,N_3169);
or U7044 (N_7044,N_3158,N_4262);
and U7045 (N_7045,N_4465,N_4969);
nor U7046 (N_7046,N_2635,N_4942);
nand U7047 (N_7047,N_3644,N_2846);
nor U7048 (N_7048,N_3202,N_4585);
nand U7049 (N_7049,N_3972,N_3081);
nor U7050 (N_7050,N_3031,N_4076);
or U7051 (N_7051,N_4544,N_4641);
and U7052 (N_7052,N_2718,N_3117);
nor U7053 (N_7053,N_4724,N_4393);
and U7054 (N_7054,N_4067,N_4684);
or U7055 (N_7055,N_3266,N_3918);
nor U7056 (N_7056,N_4460,N_4761);
or U7057 (N_7057,N_3332,N_4888);
or U7058 (N_7058,N_3042,N_2750);
nor U7059 (N_7059,N_3809,N_4968);
and U7060 (N_7060,N_3930,N_3236);
nor U7061 (N_7061,N_4705,N_2748);
nand U7062 (N_7062,N_4463,N_4816);
and U7063 (N_7063,N_4222,N_3765);
nand U7064 (N_7064,N_4620,N_3219);
or U7065 (N_7065,N_3639,N_2729);
nand U7066 (N_7066,N_4586,N_3992);
nand U7067 (N_7067,N_3211,N_3861);
nor U7068 (N_7068,N_4395,N_4060);
and U7069 (N_7069,N_3075,N_3778);
or U7070 (N_7070,N_3146,N_4865);
or U7071 (N_7071,N_3215,N_3771);
or U7072 (N_7072,N_3054,N_4911);
and U7073 (N_7073,N_3127,N_3070);
or U7074 (N_7074,N_4854,N_3048);
and U7075 (N_7075,N_3050,N_3883);
and U7076 (N_7076,N_4263,N_4131);
and U7077 (N_7077,N_2871,N_4905);
nor U7078 (N_7078,N_3655,N_4479);
and U7079 (N_7079,N_4994,N_4680);
nand U7080 (N_7080,N_2546,N_3810);
nor U7081 (N_7081,N_4693,N_4856);
nor U7082 (N_7082,N_3211,N_3035);
nor U7083 (N_7083,N_2508,N_4955);
nand U7084 (N_7084,N_4350,N_3856);
and U7085 (N_7085,N_3769,N_3698);
nand U7086 (N_7086,N_3778,N_3115);
and U7087 (N_7087,N_3168,N_3760);
nand U7088 (N_7088,N_3324,N_2793);
nor U7089 (N_7089,N_2765,N_4754);
and U7090 (N_7090,N_3001,N_3499);
or U7091 (N_7091,N_3858,N_3995);
nor U7092 (N_7092,N_3356,N_3211);
and U7093 (N_7093,N_4853,N_4786);
nor U7094 (N_7094,N_2732,N_3338);
and U7095 (N_7095,N_4780,N_3265);
nor U7096 (N_7096,N_3693,N_4171);
nand U7097 (N_7097,N_3184,N_4916);
nor U7098 (N_7098,N_3147,N_3088);
and U7099 (N_7099,N_4856,N_4314);
nor U7100 (N_7100,N_3969,N_4332);
or U7101 (N_7101,N_2894,N_4550);
or U7102 (N_7102,N_4971,N_3454);
nor U7103 (N_7103,N_2640,N_3643);
or U7104 (N_7104,N_4206,N_3505);
or U7105 (N_7105,N_4099,N_4459);
and U7106 (N_7106,N_3574,N_4879);
nand U7107 (N_7107,N_4703,N_2857);
nor U7108 (N_7108,N_4540,N_3944);
nor U7109 (N_7109,N_4006,N_4302);
nor U7110 (N_7110,N_4256,N_2651);
and U7111 (N_7111,N_2888,N_3669);
nand U7112 (N_7112,N_2581,N_4954);
nor U7113 (N_7113,N_4575,N_4415);
nand U7114 (N_7114,N_2529,N_2773);
and U7115 (N_7115,N_3773,N_3435);
and U7116 (N_7116,N_3763,N_2803);
or U7117 (N_7117,N_2722,N_4594);
nor U7118 (N_7118,N_4862,N_3590);
xor U7119 (N_7119,N_3506,N_3806);
or U7120 (N_7120,N_2666,N_4376);
or U7121 (N_7121,N_4046,N_3773);
nand U7122 (N_7122,N_2911,N_2993);
or U7123 (N_7123,N_4788,N_3426);
or U7124 (N_7124,N_3792,N_4238);
and U7125 (N_7125,N_3208,N_3008);
and U7126 (N_7126,N_4325,N_2792);
or U7127 (N_7127,N_4677,N_3061);
or U7128 (N_7128,N_3914,N_3383);
or U7129 (N_7129,N_3411,N_3542);
nor U7130 (N_7130,N_4018,N_2847);
nand U7131 (N_7131,N_4723,N_2762);
nor U7132 (N_7132,N_4182,N_3179);
and U7133 (N_7133,N_4267,N_4678);
nor U7134 (N_7134,N_2500,N_3298);
nor U7135 (N_7135,N_3202,N_3497);
or U7136 (N_7136,N_4437,N_3359);
or U7137 (N_7137,N_3312,N_3603);
and U7138 (N_7138,N_3332,N_3772);
nand U7139 (N_7139,N_3342,N_3035);
or U7140 (N_7140,N_3870,N_3031);
nor U7141 (N_7141,N_2799,N_3550);
nand U7142 (N_7142,N_3791,N_3276);
nor U7143 (N_7143,N_4470,N_2774);
nor U7144 (N_7144,N_3591,N_4567);
nand U7145 (N_7145,N_3526,N_4808);
or U7146 (N_7146,N_4926,N_3573);
and U7147 (N_7147,N_3643,N_4610);
nor U7148 (N_7148,N_4446,N_4062);
or U7149 (N_7149,N_4091,N_4634);
and U7150 (N_7150,N_3205,N_3430);
nor U7151 (N_7151,N_2557,N_3269);
nand U7152 (N_7152,N_2899,N_2709);
or U7153 (N_7153,N_4770,N_2940);
and U7154 (N_7154,N_2885,N_4103);
and U7155 (N_7155,N_2895,N_3364);
and U7156 (N_7156,N_2931,N_2927);
nand U7157 (N_7157,N_4842,N_2731);
and U7158 (N_7158,N_4293,N_3505);
and U7159 (N_7159,N_4739,N_3131);
or U7160 (N_7160,N_3530,N_4935);
xor U7161 (N_7161,N_3232,N_4721);
or U7162 (N_7162,N_4713,N_3236);
nand U7163 (N_7163,N_3141,N_3173);
and U7164 (N_7164,N_4670,N_3449);
nand U7165 (N_7165,N_4699,N_4480);
nor U7166 (N_7166,N_2983,N_3134);
nor U7167 (N_7167,N_2712,N_2744);
and U7168 (N_7168,N_2570,N_3997);
or U7169 (N_7169,N_3938,N_4879);
nand U7170 (N_7170,N_2570,N_3805);
and U7171 (N_7171,N_3605,N_4978);
nor U7172 (N_7172,N_4029,N_3533);
nor U7173 (N_7173,N_3145,N_3664);
or U7174 (N_7174,N_4610,N_3840);
nand U7175 (N_7175,N_4331,N_4184);
nor U7176 (N_7176,N_4597,N_4118);
and U7177 (N_7177,N_4898,N_2720);
and U7178 (N_7178,N_3803,N_3806);
nor U7179 (N_7179,N_4447,N_4238);
xnor U7180 (N_7180,N_3713,N_4509);
or U7181 (N_7181,N_3744,N_2744);
nor U7182 (N_7182,N_4842,N_2881);
nand U7183 (N_7183,N_3266,N_3833);
nor U7184 (N_7184,N_3476,N_2867);
nand U7185 (N_7185,N_2587,N_3763);
nor U7186 (N_7186,N_3157,N_3977);
nor U7187 (N_7187,N_4627,N_4652);
or U7188 (N_7188,N_3381,N_4932);
nor U7189 (N_7189,N_4846,N_4076);
or U7190 (N_7190,N_3082,N_4577);
nor U7191 (N_7191,N_3853,N_4491);
nor U7192 (N_7192,N_3972,N_2608);
nand U7193 (N_7193,N_3612,N_2958);
or U7194 (N_7194,N_4762,N_3586);
or U7195 (N_7195,N_4633,N_2604);
or U7196 (N_7196,N_4170,N_4106);
nor U7197 (N_7197,N_3658,N_3032);
nor U7198 (N_7198,N_3904,N_4505);
nor U7199 (N_7199,N_2841,N_4651);
or U7200 (N_7200,N_4234,N_4469);
and U7201 (N_7201,N_3247,N_3524);
and U7202 (N_7202,N_4630,N_3143);
nand U7203 (N_7203,N_4965,N_3908);
or U7204 (N_7204,N_3271,N_3993);
and U7205 (N_7205,N_4916,N_3707);
nor U7206 (N_7206,N_3393,N_3010);
nor U7207 (N_7207,N_3582,N_3506);
nor U7208 (N_7208,N_4539,N_3414);
nand U7209 (N_7209,N_4560,N_3173);
nand U7210 (N_7210,N_3218,N_3159);
or U7211 (N_7211,N_4941,N_4026);
nor U7212 (N_7212,N_3557,N_4191);
nand U7213 (N_7213,N_4861,N_2839);
and U7214 (N_7214,N_3794,N_3908);
and U7215 (N_7215,N_2771,N_4121);
nor U7216 (N_7216,N_2796,N_4724);
and U7217 (N_7217,N_3671,N_3589);
or U7218 (N_7218,N_4627,N_3083);
or U7219 (N_7219,N_4915,N_4657);
and U7220 (N_7220,N_3072,N_4135);
and U7221 (N_7221,N_3247,N_3991);
and U7222 (N_7222,N_4005,N_4143);
or U7223 (N_7223,N_4806,N_4265);
and U7224 (N_7224,N_4477,N_4676);
and U7225 (N_7225,N_4950,N_2686);
nand U7226 (N_7226,N_3128,N_3434);
xor U7227 (N_7227,N_4003,N_4165);
or U7228 (N_7228,N_4441,N_4643);
xnor U7229 (N_7229,N_3153,N_3796);
or U7230 (N_7230,N_3605,N_4069);
or U7231 (N_7231,N_4024,N_3742);
nor U7232 (N_7232,N_4600,N_4034);
nand U7233 (N_7233,N_3353,N_2754);
and U7234 (N_7234,N_4193,N_4688);
and U7235 (N_7235,N_4373,N_4089);
or U7236 (N_7236,N_4034,N_4501);
and U7237 (N_7237,N_3837,N_2907);
nor U7238 (N_7238,N_4345,N_3782);
nand U7239 (N_7239,N_4729,N_3582);
nor U7240 (N_7240,N_4291,N_2855);
and U7241 (N_7241,N_2500,N_3713);
and U7242 (N_7242,N_4360,N_4768);
or U7243 (N_7243,N_3003,N_3391);
nor U7244 (N_7244,N_4385,N_3503);
and U7245 (N_7245,N_4031,N_4496);
or U7246 (N_7246,N_4249,N_4229);
and U7247 (N_7247,N_3345,N_4052);
and U7248 (N_7248,N_4667,N_2800);
nor U7249 (N_7249,N_3082,N_3264);
or U7250 (N_7250,N_3336,N_4468);
and U7251 (N_7251,N_3870,N_2673);
or U7252 (N_7252,N_2772,N_4027);
nand U7253 (N_7253,N_4446,N_4389);
or U7254 (N_7254,N_4525,N_3167);
or U7255 (N_7255,N_3891,N_2982);
nor U7256 (N_7256,N_3474,N_3254);
or U7257 (N_7257,N_3823,N_4541);
nand U7258 (N_7258,N_4597,N_4514);
or U7259 (N_7259,N_3477,N_3259);
nor U7260 (N_7260,N_3632,N_3329);
or U7261 (N_7261,N_4092,N_4743);
and U7262 (N_7262,N_4083,N_4471);
nand U7263 (N_7263,N_3908,N_2956);
and U7264 (N_7264,N_4304,N_3906);
and U7265 (N_7265,N_3412,N_3938);
nor U7266 (N_7266,N_3875,N_3890);
and U7267 (N_7267,N_3635,N_3887);
nand U7268 (N_7268,N_2886,N_3498);
or U7269 (N_7269,N_3522,N_4193);
nand U7270 (N_7270,N_4556,N_3578);
nand U7271 (N_7271,N_2844,N_3122);
and U7272 (N_7272,N_2821,N_3549);
nand U7273 (N_7273,N_3900,N_2906);
and U7274 (N_7274,N_3613,N_4394);
or U7275 (N_7275,N_4225,N_2618);
xnor U7276 (N_7276,N_3772,N_4405);
and U7277 (N_7277,N_4309,N_4529);
or U7278 (N_7278,N_4221,N_3332);
and U7279 (N_7279,N_2607,N_4592);
or U7280 (N_7280,N_4411,N_2899);
or U7281 (N_7281,N_2536,N_4056);
or U7282 (N_7282,N_4895,N_2951);
or U7283 (N_7283,N_4885,N_3001);
nor U7284 (N_7284,N_3381,N_3296);
or U7285 (N_7285,N_3578,N_3109);
and U7286 (N_7286,N_4543,N_3094);
and U7287 (N_7287,N_3310,N_4575);
and U7288 (N_7288,N_3251,N_3535);
nor U7289 (N_7289,N_3464,N_2651);
or U7290 (N_7290,N_4650,N_4211);
or U7291 (N_7291,N_4289,N_3842);
and U7292 (N_7292,N_2738,N_3399);
nand U7293 (N_7293,N_3316,N_4548);
and U7294 (N_7294,N_4070,N_4281);
or U7295 (N_7295,N_4787,N_4404);
and U7296 (N_7296,N_4503,N_3426);
nor U7297 (N_7297,N_3030,N_3497);
and U7298 (N_7298,N_2555,N_4611);
nand U7299 (N_7299,N_4219,N_2933);
and U7300 (N_7300,N_4018,N_3047);
nand U7301 (N_7301,N_3871,N_3136);
or U7302 (N_7302,N_4170,N_2630);
nor U7303 (N_7303,N_4263,N_3325);
nor U7304 (N_7304,N_2886,N_3150);
nand U7305 (N_7305,N_4737,N_4255);
nor U7306 (N_7306,N_4123,N_2599);
nor U7307 (N_7307,N_4395,N_3721);
nor U7308 (N_7308,N_4053,N_4146);
nor U7309 (N_7309,N_4588,N_3913);
and U7310 (N_7310,N_4142,N_3102);
nand U7311 (N_7311,N_4352,N_2522);
nand U7312 (N_7312,N_3768,N_4488);
nor U7313 (N_7313,N_3749,N_3867);
and U7314 (N_7314,N_2903,N_4628);
and U7315 (N_7315,N_4041,N_2635);
or U7316 (N_7316,N_3757,N_3668);
and U7317 (N_7317,N_4243,N_4652);
or U7318 (N_7318,N_2737,N_3203);
nand U7319 (N_7319,N_4507,N_4932);
and U7320 (N_7320,N_3730,N_4689);
and U7321 (N_7321,N_4241,N_2594);
and U7322 (N_7322,N_2821,N_3323);
and U7323 (N_7323,N_3218,N_4015);
nor U7324 (N_7324,N_2643,N_4738);
nand U7325 (N_7325,N_2948,N_3542);
nor U7326 (N_7326,N_4618,N_3164);
nor U7327 (N_7327,N_3738,N_4269);
nor U7328 (N_7328,N_3806,N_3891);
nand U7329 (N_7329,N_4450,N_3433);
or U7330 (N_7330,N_4837,N_4447);
and U7331 (N_7331,N_3284,N_2556);
nor U7332 (N_7332,N_3772,N_3260);
nand U7333 (N_7333,N_4372,N_4769);
or U7334 (N_7334,N_3413,N_4166);
or U7335 (N_7335,N_3763,N_3901);
or U7336 (N_7336,N_2706,N_3574);
nor U7337 (N_7337,N_3561,N_3184);
nor U7338 (N_7338,N_3645,N_3499);
and U7339 (N_7339,N_4043,N_2706);
or U7340 (N_7340,N_3016,N_4355);
and U7341 (N_7341,N_3773,N_3844);
and U7342 (N_7342,N_4114,N_4428);
nor U7343 (N_7343,N_4313,N_4946);
nor U7344 (N_7344,N_2657,N_3466);
or U7345 (N_7345,N_3951,N_4843);
and U7346 (N_7346,N_3388,N_4849);
or U7347 (N_7347,N_2678,N_2796);
and U7348 (N_7348,N_4676,N_4513);
nor U7349 (N_7349,N_4016,N_3048);
or U7350 (N_7350,N_4147,N_2516);
nor U7351 (N_7351,N_3173,N_3831);
nand U7352 (N_7352,N_3232,N_3787);
and U7353 (N_7353,N_4550,N_3168);
nor U7354 (N_7354,N_4269,N_3546);
nand U7355 (N_7355,N_4175,N_3604);
nand U7356 (N_7356,N_4726,N_3774);
nor U7357 (N_7357,N_2973,N_4883);
nor U7358 (N_7358,N_3174,N_2551);
nor U7359 (N_7359,N_4386,N_4853);
and U7360 (N_7360,N_3076,N_4696);
and U7361 (N_7361,N_2853,N_4934);
nor U7362 (N_7362,N_4244,N_3136);
and U7363 (N_7363,N_4901,N_3166);
nor U7364 (N_7364,N_4120,N_4997);
or U7365 (N_7365,N_4891,N_2918);
and U7366 (N_7366,N_2793,N_4094);
or U7367 (N_7367,N_2694,N_4284);
or U7368 (N_7368,N_4109,N_3143);
or U7369 (N_7369,N_3906,N_2654);
or U7370 (N_7370,N_2819,N_3704);
or U7371 (N_7371,N_2651,N_4434);
or U7372 (N_7372,N_2860,N_4291);
nor U7373 (N_7373,N_3299,N_4974);
or U7374 (N_7374,N_2932,N_2573);
and U7375 (N_7375,N_4345,N_2847);
or U7376 (N_7376,N_2736,N_4377);
and U7377 (N_7377,N_2741,N_3061);
or U7378 (N_7378,N_3970,N_4071);
nand U7379 (N_7379,N_3348,N_3519);
or U7380 (N_7380,N_4732,N_4724);
nor U7381 (N_7381,N_4121,N_4041);
or U7382 (N_7382,N_3525,N_4052);
and U7383 (N_7383,N_3630,N_4389);
or U7384 (N_7384,N_3103,N_4222);
or U7385 (N_7385,N_3530,N_2805);
or U7386 (N_7386,N_4423,N_4332);
or U7387 (N_7387,N_4151,N_3770);
nand U7388 (N_7388,N_4801,N_2877);
nor U7389 (N_7389,N_2864,N_4464);
nand U7390 (N_7390,N_4415,N_2646);
and U7391 (N_7391,N_2806,N_3918);
nor U7392 (N_7392,N_4449,N_3543);
and U7393 (N_7393,N_4305,N_3753);
or U7394 (N_7394,N_3050,N_4624);
nor U7395 (N_7395,N_4926,N_3572);
nand U7396 (N_7396,N_4496,N_4769);
nand U7397 (N_7397,N_3934,N_3871);
nor U7398 (N_7398,N_4299,N_4363);
nand U7399 (N_7399,N_3769,N_3778);
nor U7400 (N_7400,N_2720,N_2949);
nand U7401 (N_7401,N_4320,N_3461);
nor U7402 (N_7402,N_3350,N_4703);
xnor U7403 (N_7403,N_4730,N_3753);
nand U7404 (N_7404,N_2929,N_3159);
or U7405 (N_7405,N_3521,N_4154);
or U7406 (N_7406,N_3546,N_2741);
nand U7407 (N_7407,N_3000,N_3318);
nand U7408 (N_7408,N_2731,N_3217);
and U7409 (N_7409,N_4037,N_4570);
nand U7410 (N_7410,N_3217,N_4133);
or U7411 (N_7411,N_3604,N_3463);
nor U7412 (N_7412,N_4419,N_3024);
nor U7413 (N_7413,N_2927,N_2920);
nor U7414 (N_7414,N_2679,N_4655);
nor U7415 (N_7415,N_2885,N_3291);
and U7416 (N_7416,N_4083,N_4224);
nor U7417 (N_7417,N_2888,N_2637);
or U7418 (N_7418,N_4809,N_4639);
nor U7419 (N_7419,N_3630,N_3328);
nand U7420 (N_7420,N_4894,N_2543);
xor U7421 (N_7421,N_3049,N_4710);
nor U7422 (N_7422,N_2967,N_3692);
or U7423 (N_7423,N_3773,N_4094);
nor U7424 (N_7424,N_2665,N_4892);
nor U7425 (N_7425,N_3561,N_2602);
nand U7426 (N_7426,N_3274,N_3300);
or U7427 (N_7427,N_3011,N_4951);
or U7428 (N_7428,N_3423,N_3524);
nor U7429 (N_7429,N_3051,N_3100);
nor U7430 (N_7430,N_3648,N_4834);
or U7431 (N_7431,N_3109,N_4264);
xnor U7432 (N_7432,N_3898,N_4185);
and U7433 (N_7433,N_3741,N_3040);
or U7434 (N_7434,N_4755,N_2900);
or U7435 (N_7435,N_4885,N_4293);
and U7436 (N_7436,N_4086,N_2897);
or U7437 (N_7437,N_3017,N_4818);
or U7438 (N_7438,N_3030,N_3793);
or U7439 (N_7439,N_3741,N_3739);
nand U7440 (N_7440,N_4012,N_3252);
nand U7441 (N_7441,N_3889,N_3907);
or U7442 (N_7442,N_4290,N_4736);
and U7443 (N_7443,N_4216,N_4831);
or U7444 (N_7444,N_2509,N_2661);
nor U7445 (N_7445,N_3194,N_3461);
nor U7446 (N_7446,N_3029,N_4677);
xor U7447 (N_7447,N_4956,N_3455);
nor U7448 (N_7448,N_2892,N_4290);
nand U7449 (N_7449,N_4684,N_3360);
or U7450 (N_7450,N_4205,N_2988);
nor U7451 (N_7451,N_4043,N_2819);
and U7452 (N_7452,N_4834,N_2753);
nand U7453 (N_7453,N_4418,N_2846);
or U7454 (N_7454,N_3875,N_3726);
nor U7455 (N_7455,N_2902,N_2896);
and U7456 (N_7456,N_4868,N_4758);
or U7457 (N_7457,N_4876,N_4133);
nand U7458 (N_7458,N_2918,N_3107);
or U7459 (N_7459,N_3118,N_4143);
nor U7460 (N_7460,N_2964,N_4268);
nor U7461 (N_7461,N_4903,N_4207);
or U7462 (N_7462,N_3776,N_3758);
nand U7463 (N_7463,N_4601,N_3702);
nand U7464 (N_7464,N_4818,N_2895);
or U7465 (N_7465,N_4154,N_3160);
nor U7466 (N_7466,N_4465,N_4803);
nand U7467 (N_7467,N_3048,N_3314);
and U7468 (N_7468,N_2931,N_4257);
and U7469 (N_7469,N_4489,N_3126);
nand U7470 (N_7470,N_3753,N_3535);
or U7471 (N_7471,N_3655,N_4236);
or U7472 (N_7472,N_3894,N_4032);
nor U7473 (N_7473,N_4193,N_4426);
or U7474 (N_7474,N_4997,N_4125);
or U7475 (N_7475,N_3884,N_3481);
and U7476 (N_7476,N_3402,N_4792);
nand U7477 (N_7477,N_3715,N_2857);
or U7478 (N_7478,N_3827,N_3337);
nand U7479 (N_7479,N_2549,N_3247);
nor U7480 (N_7480,N_4086,N_4336);
and U7481 (N_7481,N_4927,N_3047);
nand U7482 (N_7482,N_3416,N_2774);
nor U7483 (N_7483,N_3180,N_3893);
nand U7484 (N_7484,N_3905,N_4524);
and U7485 (N_7485,N_3580,N_2628);
and U7486 (N_7486,N_3555,N_4309);
nor U7487 (N_7487,N_4985,N_3926);
or U7488 (N_7488,N_4901,N_4703);
and U7489 (N_7489,N_4533,N_3714);
or U7490 (N_7490,N_3212,N_3421);
nand U7491 (N_7491,N_2666,N_3109);
or U7492 (N_7492,N_4527,N_3577);
or U7493 (N_7493,N_4945,N_4645);
and U7494 (N_7494,N_3912,N_3802);
nor U7495 (N_7495,N_4612,N_4014);
or U7496 (N_7496,N_2976,N_3817);
nand U7497 (N_7497,N_3040,N_2540);
and U7498 (N_7498,N_3046,N_4299);
nand U7499 (N_7499,N_3358,N_4583);
xnor U7500 (N_7500,N_5856,N_6871);
xor U7501 (N_7501,N_6034,N_5857);
and U7502 (N_7502,N_5181,N_6905);
nand U7503 (N_7503,N_5158,N_5116);
nor U7504 (N_7504,N_6669,N_5866);
nor U7505 (N_7505,N_5802,N_6341);
and U7506 (N_7506,N_5677,N_7276);
and U7507 (N_7507,N_5728,N_6052);
nor U7508 (N_7508,N_6105,N_5597);
nand U7509 (N_7509,N_5273,N_7200);
nor U7510 (N_7510,N_7039,N_6569);
or U7511 (N_7511,N_6759,N_6789);
or U7512 (N_7512,N_5548,N_7082);
and U7513 (N_7513,N_5893,N_7202);
or U7514 (N_7514,N_5163,N_6324);
nand U7515 (N_7515,N_6302,N_5274);
or U7516 (N_7516,N_5456,N_7259);
or U7517 (N_7517,N_6749,N_7454);
nor U7518 (N_7518,N_5926,N_6387);
and U7519 (N_7519,N_7499,N_5519);
and U7520 (N_7520,N_6217,N_5780);
and U7521 (N_7521,N_6991,N_6157);
nor U7522 (N_7522,N_6875,N_6608);
or U7523 (N_7523,N_6014,N_5094);
or U7524 (N_7524,N_5422,N_5304);
and U7525 (N_7525,N_6045,N_7497);
and U7526 (N_7526,N_6584,N_6778);
nor U7527 (N_7527,N_7262,N_5712);
and U7528 (N_7528,N_7461,N_6076);
nand U7529 (N_7529,N_5336,N_6472);
and U7530 (N_7530,N_6912,N_5298);
or U7531 (N_7531,N_6420,N_5371);
or U7532 (N_7532,N_5377,N_5930);
nor U7533 (N_7533,N_6786,N_5753);
and U7534 (N_7534,N_5560,N_7065);
or U7535 (N_7535,N_5318,N_6475);
nand U7536 (N_7536,N_6412,N_6171);
or U7537 (N_7537,N_7296,N_7046);
or U7538 (N_7538,N_6868,N_5536);
and U7539 (N_7539,N_6444,N_5195);
and U7540 (N_7540,N_6974,N_7165);
nor U7541 (N_7541,N_5529,N_6518);
or U7542 (N_7542,N_5632,N_7184);
and U7543 (N_7543,N_5769,N_6048);
nor U7544 (N_7544,N_5933,N_7058);
and U7545 (N_7545,N_5767,N_7033);
and U7546 (N_7546,N_6941,N_6292);
and U7547 (N_7547,N_5807,N_5287);
nor U7548 (N_7548,N_6657,N_5007);
nor U7549 (N_7549,N_7164,N_5290);
nand U7550 (N_7550,N_7224,N_5027);
nand U7551 (N_7551,N_5004,N_5967);
nand U7552 (N_7552,N_6476,N_7087);
and U7553 (N_7553,N_6561,N_7193);
and U7554 (N_7554,N_5420,N_5858);
nand U7555 (N_7555,N_6655,N_6506);
nor U7556 (N_7556,N_6768,N_5294);
and U7557 (N_7557,N_6590,N_5894);
or U7558 (N_7558,N_6918,N_6524);
or U7559 (N_7559,N_7206,N_5948);
and U7560 (N_7560,N_5830,N_5014);
nand U7561 (N_7561,N_6581,N_6451);
xor U7562 (N_7562,N_6046,N_6252);
and U7563 (N_7563,N_6445,N_6139);
nor U7564 (N_7564,N_6194,N_6234);
and U7565 (N_7565,N_6520,N_6049);
and U7566 (N_7566,N_5144,N_5434);
nand U7567 (N_7567,N_6887,N_5212);
nand U7568 (N_7568,N_7068,N_6044);
nand U7569 (N_7569,N_6151,N_5929);
nand U7570 (N_7570,N_6062,N_7061);
and U7571 (N_7571,N_5036,N_7270);
nand U7572 (N_7572,N_6714,N_6345);
nand U7573 (N_7573,N_5480,N_5887);
and U7574 (N_7574,N_6943,N_7094);
nor U7575 (N_7575,N_7089,N_6240);
or U7576 (N_7576,N_7234,N_7322);
and U7577 (N_7577,N_5576,N_5556);
and U7578 (N_7578,N_6056,N_5716);
nor U7579 (N_7579,N_5917,N_7097);
nor U7580 (N_7580,N_7182,N_6270);
or U7581 (N_7581,N_6334,N_7060);
nand U7582 (N_7582,N_6167,N_5414);
and U7583 (N_7583,N_7249,N_6266);
and U7584 (N_7584,N_7319,N_7080);
nand U7585 (N_7585,N_5932,N_6253);
nor U7586 (N_7586,N_6419,N_7291);
or U7587 (N_7587,N_6214,N_6884);
nand U7588 (N_7588,N_7205,N_6588);
nor U7589 (N_7589,N_6104,N_5341);
nand U7590 (N_7590,N_5906,N_5310);
nor U7591 (N_7591,N_5477,N_5628);
nand U7592 (N_7592,N_7473,N_5847);
and U7593 (N_7593,N_7337,N_5166);
and U7594 (N_7594,N_5111,N_6114);
nand U7595 (N_7595,N_5385,N_7051);
and U7596 (N_7596,N_6528,N_5380);
or U7597 (N_7597,N_5312,N_6067);
or U7598 (N_7598,N_5331,N_6374);
and U7599 (N_7599,N_6946,N_5621);
and U7600 (N_7600,N_7154,N_5538);
and U7601 (N_7601,N_6275,N_7000);
and U7602 (N_7602,N_6615,N_6351);
and U7603 (N_7603,N_5271,N_7382);
nand U7604 (N_7604,N_5794,N_6957);
and U7605 (N_7605,N_5759,N_5810);
nor U7606 (N_7606,N_6913,N_5539);
nor U7607 (N_7607,N_6935,N_5194);
nor U7608 (N_7608,N_5708,N_7278);
and U7609 (N_7609,N_6764,N_5622);
or U7610 (N_7610,N_5224,N_6425);
nor U7611 (N_7611,N_6478,N_6304);
and U7612 (N_7612,N_5461,N_6666);
nor U7613 (N_7613,N_7323,N_6002);
and U7614 (N_7614,N_5695,N_6646);
nor U7615 (N_7615,N_7367,N_5132);
nor U7616 (N_7616,N_6070,N_5394);
nor U7617 (N_7617,N_6068,N_7196);
or U7618 (N_7618,N_5077,N_6720);
nor U7619 (N_7619,N_5600,N_5988);
nor U7620 (N_7620,N_7340,N_7242);
nand U7621 (N_7621,N_5282,N_6822);
or U7622 (N_7622,N_5201,N_6687);
nor U7623 (N_7623,N_5900,N_6522);
nor U7624 (N_7624,N_7434,N_6592);
and U7625 (N_7625,N_5444,N_6810);
or U7626 (N_7626,N_5185,N_5500);
nand U7627 (N_7627,N_5903,N_5247);
nor U7628 (N_7628,N_7239,N_5923);
or U7629 (N_7629,N_7045,N_6161);
and U7630 (N_7630,N_5675,N_6402);
and U7631 (N_7631,N_5211,N_6496);
nor U7632 (N_7632,N_6814,N_5521);
and U7633 (N_7633,N_5925,N_5100);
and U7634 (N_7634,N_7062,N_6315);
nand U7635 (N_7635,N_7431,N_6342);
nand U7636 (N_7636,N_6670,N_7130);
nand U7637 (N_7637,N_7019,N_7448);
nor U7638 (N_7638,N_6075,N_6724);
or U7639 (N_7639,N_6087,N_5286);
nor U7640 (N_7640,N_5293,N_6298);
nor U7641 (N_7641,N_7118,N_5882);
or U7642 (N_7642,N_5612,N_6256);
nand U7643 (N_7643,N_6538,N_6272);
nor U7644 (N_7644,N_5751,N_6683);
nand U7645 (N_7645,N_6664,N_5474);
nor U7646 (N_7646,N_5797,N_5245);
or U7647 (N_7647,N_6812,N_5075);
nor U7648 (N_7648,N_6083,N_5868);
nor U7649 (N_7649,N_5848,N_5180);
nand U7650 (N_7650,N_7447,N_7251);
or U7651 (N_7651,N_5179,N_6689);
and U7652 (N_7652,N_6771,N_6368);
xor U7653 (N_7653,N_6785,N_7144);
or U7654 (N_7654,N_7308,N_6774);
and U7655 (N_7655,N_5637,N_5469);
nor U7656 (N_7656,N_5955,N_5426);
nand U7657 (N_7657,N_6096,N_5233);
nand U7658 (N_7658,N_6550,N_5827);
nor U7659 (N_7659,N_5066,N_6951);
and U7660 (N_7660,N_7160,N_5186);
and U7661 (N_7661,N_5470,N_6848);
and U7662 (N_7662,N_5995,N_6316);
nor U7663 (N_7663,N_5513,N_5392);
or U7664 (N_7664,N_6441,N_7336);
nand U7665 (N_7665,N_5042,N_6995);
nand U7666 (N_7666,N_6880,N_6635);
nand U7667 (N_7667,N_6416,N_7283);
nor U7668 (N_7668,N_5402,N_6755);
nor U7669 (N_7669,N_6955,N_7198);
and U7670 (N_7670,N_5162,N_5819);
or U7671 (N_7671,N_5611,N_7096);
and U7672 (N_7672,N_6211,N_6858);
and U7673 (N_7673,N_6611,N_5199);
and U7674 (N_7674,N_6001,N_5197);
nor U7675 (N_7675,N_6806,N_7493);
or U7676 (N_7676,N_5129,N_6127);
nand U7677 (N_7677,N_5815,N_5733);
nor U7678 (N_7678,N_7083,N_6949);
nand U7679 (N_7679,N_6403,N_5373);
and U7680 (N_7680,N_6996,N_5326);
nand U7681 (N_7681,N_6357,N_5095);
nand U7682 (N_7682,N_6066,N_6968);
nor U7683 (N_7683,N_7360,N_7380);
nand U7684 (N_7684,N_5320,N_6264);
or U7685 (N_7685,N_7158,N_7100);
nand U7686 (N_7686,N_7248,N_7405);
nor U7687 (N_7687,N_6366,N_5241);
or U7688 (N_7688,N_6484,N_5124);
nor U7689 (N_7689,N_7150,N_5289);
and U7690 (N_7690,N_6643,N_5172);
or U7691 (N_7691,N_5410,N_5169);
nand U7692 (N_7692,N_6313,N_6100);
nor U7693 (N_7693,N_5656,N_7174);
nand U7694 (N_7694,N_5142,N_6805);
nor U7695 (N_7695,N_6371,N_6906);
nor U7696 (N_7696,N_7294,N_6542);
or U7697 (N_7697,N_5861,N_7432);
nor U7698 (N_7698,N_5641,N_6291);
nand U7699 (N_7699,N_5306,N_5024);
and U7700 (N_7700,N_5540,N_6598);
nand U7701 (N_7701,N_6808,N_5037);
nand U7702 (N_7702,N_7298,N_6874);
or U7703 (N_7703,N_5704,N_6121);
nor U7704 (N_7704,N_5873,N_6709);
nor U7705 (N_7705,N_5001,N_5419);
or U7706 (N_7706,N_5453,N_6492);
nor U7707 (N_7707,N_7002,N_7371);
nor U7708 (N_7708,N_6944,N_6978);
or U7709 (N_7709,N_5798,N_6556);
nand U7710 (N_7710,N_5601,N_6471);
nand U7711 (N_7711,N_5821,N_6861);
and U7712 (N_7712,N_5030,N_6244);
and U7713 (N_7713,N_6959,N_5292);
nor U7714 (N_7714,N_6443,N_5565);
nor U7715 (N_7715,N_5936,N_7456);
and U7716 (N_7716,N_6470,N_5046);
or U7717 (N_7717,N_6525,N_5697);
nor U7718 (N_7718,N_5329,N_5057);
nor U7719 (N_7719,N_7467,N_6006);
and U7720 (N_7720,N_6748,N_5911);
nor U7721 (N_7721,N_6367,N_7219);
nor U7722 (N_7722,N_7304,N_6932);
nor U7723 (N_7723,N_5105,N_5221);
nor U7724 (N_7724,N_6558,N_7166);
nor U7725 (N_7725,N_5796,N_5460);
or U7726 (N_7726,N_7204,N_6747);
and U7727 (N_7727,N_6889,N_7085);
or U7728 (N_7728,N_5690,N_6450);
and U7729 (N_7729,N_7066,N_5491);
or U7730 (N_7730,N_6767,N_5942);
nor U7731 (N_7731,N_6411,N_5840);
nor U7732 (N_7732,N_7269,N_5227);
or U7733 (N_7733,N_7250,N_5526);
nand U7734 (N_7734,N_5964,N_6656);
and U7735 (N_7735,N_7403,N_6204);
or U7736 (N_7736,N_6094,N_5515);
nor U7737 (N_7737,N_6365,N_7318);
nor U7738 (N_7738,N_7077,N_5891);
nand U7739 (N_7739,N_5897,N_6220);
and U7740 (N_7740,N_6653,N_5455);
nand U7741 (N_7741,N_5492,N_5525);
nand U7742 (N_7742,N_5191,N_5358);
or U7743 (N_7743,N_6277,N_5645);
and U7744 (N_7744,N_7314,N_5725);
nor U7745 (N_7745,N_6756,N_6997);
nor U7746 (N_7746,N_5533,N_6933);
or U7747 (N_7747,N_7346,N_6973);
or U7748 (N_7748,N_7284,N_5164);
or U7749 (N_7749,N_7306,N_5761);
and U7750 (N_7750,N_6809,N_5123);
nor U7751 (N_7751,N_5086,N_5019);
nand U7752 (N_7752,N_5251,N_6110);
nand U7753 (N_7753,N_5741,N_5720);
nand U7754 (N_7754,N_6072,N_6576);
nor U7755 (N_7755,N_5334,N_5136);
nand U7756 (N_7756,N_6945,N_7411);
or U7757 (N_7757,N_5583,N_5333);
nor U7758 (N_7758,N_5701,N_5018);
or U7759 (N_7759,N_7307,N_5008);
or U7760 (N_7760,N_7013,N_6084);
nor U7761 (N_7761,N_5584,N_6318);
and U7762 (N_7762,N_6773,N_5451);
or U7763 (N_7763,N_7420,N_5048);
nor U7764 (N_7764,N_5825,N_5087);
nand U7765 (N_7765,N_6727,N_7135);
and U7766 (N_7766,N_5564,N_6007);
or U7767 (N_7767,N_7483,N_6831);
and U7768 (N_7768,N_6119,N_5770);
nor U7769 (N_7769,N_5698,N_5888);
nor U7770 (N_7770,N_6845,N_5514);
or U7771 (N_7771,N_5412,N_6591);
nor U7772 (N_7772,N_5442,N_5726);
nand U7773 (N_7773,N_6852,N_5907);
nor U7774 (N_7774,N_5052,N_7071);
nor U7775 (N_7775,N_6925,N_5384);
nor U7776 (N_7776,N_7084,N_5330);
nor U7777 (N_7777,N_7098,N_5416);
or U7778 (N_7778,N_7417,N_7407);
and U7779 (N_7779,N_5188,N_7038);
nor U7780 (N_7780,N_5051,N_5649);
nor U7781 (N_7781,N_6866,N_5535);
or U7782 (N_7782,N_6940,N_5204);
nor U7783 (N_7783,N_5634,N_6661);
nand U7784 (N_7784,N_5029,N_6029);
and U7785 (N_7785,N_7067,N_5060);
or U7786 (N_7786,N_5317,N_6468);
and U7787 (N_7787,N_6827,N_5844);
and U7788 (N_7788,N_7101,N_5122);
nand U7789 (N_7789,N_5603,N_6983);
or U7790 (N_7790,N_5192,N_6409);
nor U7791 (N_7791,N_5763,N_6290);
nand U7792 (N_7792,N_6490,N_5680);
or U7793 (N_7793,N_5393,N_6899);
and U7794 (N_7794,N_5218,N_7173);
nand U7795 (N_7795,N_6516,N_5619);
nor U7796 (N_7796,N_6872,N_7063);
or U7797 (N_7797,N_7175,N_6566);
nor U7798 (N_7798,N_6849,N_5272);
nor U7799 (N_7799,N_6249,N_5776);
and U7800 (N_7800,N_5939,N_7436);
or U7801 (N_7801,N_5719,N_5731);
and U7802 (N_7802,N_7147,N_5240);
nor U7803 (N_7803,N_6429,N_6833);
and U7804 (N_7804,N_6385,N_6065);
or U7805 (N_7805,N_6461,N_5730);
nand U7806 (N_7806,N_5744,N_7243);
nand U7807 (N_7807,N_6855,N_6553);
or U7808 (N_7808,N_6843,N_5604);
nor U7809 (N_7809,N_5285,N_6937);
nand U7810 (N_7810,N_6711,N_5035);
nor U7811 (N_7811,N_5448,N_6869);
or U7812 (N_7812,N_5015,N_5345);
nand U7813 (N_7813,N_5954,N_5626);
or U7814 (N_7814,N_5703,N_5774);
nor U7815 (N_7815,N_5465,N_5280);
and U7816 (N_7816,N_5022,N_6015);
nor U7817 (N_7817,N_7273,N_6606);
nand U7818 (N_7818,N_7469,N_7415);
or U7819 (N_7819,N_5013,N_6297);
nand U7820 (N_7820,N_5616,N_5457);
and U7821 (N_7821,N_5112,N_6514);
nor U7822 (N_7822,N_7492,N_5588);
nor U7823 (N_7823,N_6099,N_6281);
nand U7824 (N_7824,N_5752,N_5546);
or U7825 (N_7825,N_5629,N_6354);
and U7826 (N_7826,N_5459,N_5278);
nand U7827 (N_7827,N_5405,N_7124);
xnor U7828 (N_7828,N_6010,N_6609);
and U7829 (N_7829,N_7229,N_6642);
and U7830 (N_7830,N_5106,N_5440);
and U7831 (N_7831,N_6457,N_6688);
and U7832 (N_7832,N_6469,N_7095);
and U7833 (N_7833,N_6307,N_7169);
or U7834 (N_7834,N_5579,N_5828);
nor U7835 (N_7835,N_5625,N_5507);
or U7836 (N_7836,N_7120,N_5950);
and U7837 (N_7837,N_6430,N_6740);
nand U7838 (N_7838,N_5544,N_5149);
nand U7839 (N_7839,N_5554,N_6488);
nor U7840 (N_7840,N_5322,N_6265);
nor U7841 (N_7841,N_6706,N_5337);
and U7842 (N_7842,N_6090,N_6859);
nand U7843 (N_7843,N_6624,N_6942);
or U7844 (N_7844,N_6662,N_7451);
nand U7845 (N_7845,N_5391,N_7444);
nand U7846 (N_7846,N_6465,N_6107);
or U7847 (N_7847,N_7455,N_7064);
and U7848 (N_7848,N_5362,N_7321);
nand U7849 (N_7849,N_7352,N_6156);
nand U7850 (N_7850,N_7127,N_5458);
or U7851 (N_7851,N_7297,N_6552);
nand U7852 (N_7852,N_6260,N_5313);
or U7853 (N_7853,N_7238,N_5646);
or U7854 (N_7854,N_6971,N_5934);
nor U7855 (N_7855,N_6452,N_6735);
nor U7856 (N_7856,N_5792,N_5928);
nor U7857 (N_7857,N_5432,N_7470);
and U7858 (N_7858,N_5811,N_7464);
nand U7859 (N_7859,N_5660,N_5998);
and U7860 (N_7860,N_5779,N_6545);
nand U7861 (N_7861,N_6219,N_6464);
or U7862 (N_7862,N_6819,N_5973);
and U7863 (N_7863,N_6563,N_6703);
and U7864 (N_7864,N_7342,N_6400);
nor U7865 (N_7865,N_6381,N_7138);
nor U7866 (N_7866,N_6574,N_6562);
nand U7867 (N_7867,N_5679,N_6477);
and U7868 (N_7868,N_5231,N_6881);
and U7869 (N_7869,N_5396,N_5184);
and U7870 (N_7870,N_6614,N_7264);
nand U7871 (N_7871,N_5356,N_5376);
nor U7872 (N_7872,N_6329,N_6212);
nand U7873 (N_7873,N_7438,N_7237);
nor U7874 (N_7874,N_6877,N_6434);
nor U7875 (N_7875,N_6684,N_5167);
or U7876 (N_7876,N_7156,N_6305);
and U7877 (N_7877,N_5147,N_6972);
and U7878 (N_7878,N_6123,N_5746);
or U7879 (N_7879,N_5642,N_5002);
and U7880 (N_7880,N_5667,N_5239);
or U7881 (N_7881,N_7358,N_7162);
nor U7882 (N_7882,N_6440,N_5993);
and U7883 (N_7883,N_6388,N_6082);
or U7884 (N_7884,N_5153,N_5053);
nor U7885 (N_7885,N_7222,N_5640);
and U7886 (N_7886,N_6725,N_5319);
and U7887 (N_7887,N_6557,N_6987);
or U7888 (N_7888,N_6141,N_6456);
nand U7889 (N_7889,N_5814,N_6485);
nand U7890 (N_7890,N_6190,N_7212);
nor U7891 (N_7891,N_7384,N_7365);
nand U7892 (N_7892,N_5068,N_6251);
or U7893 (N_7893,N_6707,N_6186);
or U7894 (N_7894,N_7208,N_6311);
nand U7895 (N_7895,N_6481,N_7379);
or U7896 (N_7896,N_7295,N_5791);
nor U7897 (N_7897,N_7446,N_6101);
nor U7898 (N_7898,N_5812,N_6746);
or U7899 (N_7899,N_5784,N_5824);
and U7900 (N_7900,N_6020,N_5837);
or U7901 (N_7901,N_7285,N_7134);
and U7902 (N_7902,N_5764,N_7481);
nor U7903 (N_7903,N_7290,N_6989);
nor U7904 (N_7904,N_7163,N_5501);
nand U7905 (N_7905,N_7011,N_5665);
nor U7906 (N_7906,N_5269,N_5177);
nand U7907 (N_7907,N_6549,N_5034);
nor U7908 (N_7908,N_5388,N_6081);
or U7909 (N_7909,N_6799,N_6701);
nor U7910 (N_7910,N_5284,N_6055);
nor U7911 (N_7911,N_5476,N_5938);
and U7912 (N_7912,N_5099,N_6384);
nor U7913 (N_7913,N_7378,N_5982);
nor U7914 (N_7914,N_6348,N_5056);
or U7915 (N_7915,N_6137,N_7474);
or U7916 (N_7916,N_6405,N_6353);
or U7917 (N_7917,N_5482,N_6836);
nor U7918 (N_7918,N_6061,N_5131);
nor U7919 (N_7919,N_6829,N_6031);
and U7920 (N_7920,N_6763,N_6572);
nor U7921 (N_7921,N_6271,N_6954);
or U7922 (N_7922,N_5101,N_6734);
nor U7923 (N_7923,N_7133,N_5570);
or U7924 (N_7924,N_6335,N_5441);
xor U7925 (N_7925,N_7075,N_5209);
nand U7926 (N_7926,N_7494,N_6494);
nor U7927 (N_7927,N_6640,N_5527);
and U7928 (N_7928,N_5109,N_5510);
and U7929 (N_7929,N_6089,N_5061);
nor U7930 (N_7930,N_5499,N_5424);
nor U7931 (N_7931,N_5838,N_7197);
or U7932 (N_7932,N_6507,N_5026);
or U7933 (N_7933,N_5816,N_6617);
nand U7934 (N_7934,N_5081,N_6998);
nand U7935 (N_7935,N_7185,N_7201);
nor U7936 (N_7936,N_6395,N_7139);
and U7937 (N_7937,N_6308,N_6603);
and U7938 (N_7938,N_6926,N_5003);
nor U7939 (N_7939,N_7400,N_5021);
nor U7940 (N_7940,N_5038,N_6482);
and U7941 (N_7941,N_7374,N_5648);
nand U7942 (N_7942,N_5479,N_5425);
and U7943 (N_7943,N_6043,N_6179);
and U7944 (N_7944,N_7149,N_5531);
nor U7945 (N_7945,N_5495,N_5586);
and U7946 (N_7946,N_6969,N_7361);
nor U7947 (N_7947,N_7181,N_6191);
or U7948 (N_7948,N_7031,N_5437);
nor U7949 (N_7949,N_6312,N_6599);
or U7950 (N_7950,N_6363,N_6509);
nor U7951 (N_7951,N_6605,N_6399);
or U7952 (N_7952,N_5745,N_6948);
and U7953 (N_7953,N_6792,N_6300);
and U7954 (N_7954,N_5781,N_5578);
or U7955 (N_7955,N_6261,N_7034);
or U7956 (N_7956,N_6559,N_5711);
nand U7957 (N_7957,N_6144,N_6633);
nand U7958 (N_7958,N_5655,N_5864);
and U7959 (N_7959,N_6442,N_6543);
or U7960 (N_7960,N_7091,N_6970);
or U7961 (N_7961,N_5407,N_6723);
nand U7962 (N_7962,N_6934,N_6436);
and U7963 (N_7963,N_6761,N_6344);
and U7964 (N_7964,N_5859,N_5598);
nor U7965 (N_7965,N_5567,N_6691);
nand U7966 (N_7966,N_6659,N_6589);
nand U7967 (N_7967,N_6473,N_6920);
nor U7968 (N_7968,N_6663,N_6333);
and U7969 (N_7969,N_6517,N_5126);
nor U7970 (N_7970,N_6890,N_7328);
and U7971 (N_7971,N_5562,N_7110);
and U7972 (N_7972,N_5127,N_7332);
and U7973 (N_7973,N_5108,N_7073);
and U7974 (N_7974,N_6393,N_5252);
or U7975 (N_7975,N_6169,N_7217);
nand U7976 (N_7976,N_7114,N_5069);
nor U7977 (N_7977,N_7305,N_5876);
and U7978 (N_7978,N_5276,N_5497);
and U7979 (N_7979,N_6648,N_6676);
nand U7980 (N_7980,N_7123,N_5987);
or U7981 (N_7981,N_6057,N_5691);
nand U7982 (N_7982,N_7443,N_5755);
nand U7983 (N_7983,N_7107,N_6960);
or U7984 (N_7984,N_6188,N_6967);
nor U7985 (N_7985,N_6437,N_7427);
xor U7986 (N_7986,N_7194,N_6654);
or U7987 (N_7987,N_6459,N_7035);
nand U7988 (N_7988,N_7300,N_6246);
nand U7989 (N_7989,N_5210,N_7442);
and U7990 (N_7990,N_5074,N_7122);
nand U7991 (N_7991,N_5113,N_6607);
or U7992 (N_7992,N_7070,N_5820);
or U7993 (N_7993,N_6327,N_5503);
nor U7994 (N_7994,N_5589,N_7007);
nor U7995 (N_7995,N_6779,N_5267);
or U7996 (N_7996,N_6821,N_6573);
nor U7997 (N_7997,N_6794,N_6879);
and U7998 (N_7998,N_5238,N_5735);
nand U7999 (N_7999,N_5960,N_6206);
nand U8000 (N_8000,N_7195,N_5010);
nand U8001 (N_8001,N_6856,N_7396);
or U8002 (N_8002,N_6894,N_5742);
nor U8003 (N_8003,N_5846,N_6751);
or U8004 (N_8004,N_5110,N_6565);
and U8005 (N_8005,N_5165,N_5257);
nand U8006 (N_8006,N_7188,N_5624);
nand U8007 (N_8007,N_5323,N_5545);
and U8008 (N_8008,N_6233,N_5722);
nand U8009 (N_8009,N_7449,N_5765);
and U8010 (N_8010,N_5591,N_5534);
or U8011 (N_8011,N_6752,N_7490);
nand U8012 (N_8012,N_6975,N_5650);
and U8013 (N_8013,N_5307,N_5549);
nand U8014 (N_8014,N_5009,N_6842);
nor U8015 (N_8015,N_6458,N_5653);
or U8016 (N_8016,N_6702,N_7445);
or U8017 (N_8017,N_7260,N_7406);
nor U8018 (N_8018,N_5343,N_7236);
and U8019 (N_8019,N_5085,N_7151);
and U8020 (N_8020,N_6375,N_6804);
nand U8021 (N_8021,N_5399,N_7303);
or U8022 (N_8022,N_6143,N_5528);
or U8023 (N_8023,N_6873,N_7496);
or U8024 (N_8024,N_5615,N_5990);
or U8025 (N_8025,N_7186,N_5740);
and U8026 (N_8026,N_5732,N_5446);
or U8027 (N_8027,N_6404,N_5404);
and U8028 (N_8028,N_5854,N_6626);
nand U8029 (N_8029,N_7111,N_5901);
nor U8030 (N_8030,N_7301,N_6762);
nor U8031 (N_8031,N_5978,N_6146);
nor U8032 (N_8032,N_5058,N_6377);
nor U8033 (N_8033,N_6343,N_6225);
nor U8034 (N_8034,N_6467,N_7310);
nor U8035 (N_8035,N_6373,N_7488);
nor U8036 (N_8036,N_6278,N_5793);
nand U8037 (N_8037,N_5915,N_6340);
nand U8038 (N_8038,N_7440,N_6355);
or U8039 (N_8039,N_6575,N_7430);
nand U8040 (N_8040,N_6346,N_5193);
nand U8041 (N_8041,N_5134,N_6314);
nor U8042 (N_8042,N_5871,N_5916);
nor U8043 (N_8043,N_7183,N_5135);
nand U8044 (N_8044,N_6596,N_7159);
or U8045 (N_8045,N_5486,N_6039);
nor U8046 (N_8046,N_7463,N_7281);
nor U8047 (N_8047,N_5032,N_7452);
and U8048 (N_8048,N_6394,N_5115);
nor U8049 (N_8049,N_6782,N_5630);
nor U8050 (N_8050,N_6455,N_5788);
or U8051 (N_8051,N_6585,N_6284);
nor U8052 (N_8052,N_7274,N_5870);
and U8053 (N_8053,N_7362,N_6736);
and U8054 (N_8054,N_5639,N_7267);
and U8055 (N_8055,N_6199,N_5305);
nor U8056 (N_8056,N_7213,N_5509);
nor U8057 (N_8057,N_5994,N_5524);
and U8058 (N_8058,N_6111,N_6447);
nand U8059 (N_8059,N_5372,N_7040);
nand U8060 (N_8060,N_5488,N_6147);
or U8061 (N_8061,N_7105,N_6628);
nor U8062 (N_8062,N_5920,N_5965);
nor U8063 (N_8063,N_5582,N_5547);
nand U8064 (N_8064,N_6036,N_5299);
nand U8065 (N_8065,N_6548,N_6232);
nand U8066 (N_8066,N_7252,N_5705);
nor U8067 (N_8067,N_6904,N_6699);
nand U8068 (N_8068,N_6780,N_5574);
or U8069 (N_8069,N_6356,N_7112);
nand U8070 (N_8070,N_5980,N_5706);
nor U8071 (N_8071,N_5359,N_5614);
or U8072 (N_8072,N_7155,N_5205);
nor U8073 (N_8073,N_7228,N_6248);
and U8074 (N_8074,N_5092,N_7121);
or U8075 (N_8075,N_5747,N_5300);
nor U8076 (N_8076,N_5504,N_5062);
nand U8077 (N_8077,N_5071,N_5606);
and U8078 (N_8078,N_5572,N_6929);
nor U8079 (N_8079,N_6237,N_5349);
nand U8080 (N_8080,N_7137,N_6433);
or U8081 (N_8081,N_7235,N_6682);
nor U8082 (N_8082,N_7117,N_6531);
nor U8083 (N_8083,N_6483,N_6163);
and U8084 (N_8084,N_6888,N_6729);
or U8085 (N_8085,N_7171,N_7435);
nand U8086 (N_8086,N_5610,N_6336);
nor U8087 (N_8087,N_7218,N_5734);
or U8088 (N_8088,N_5198,N_5281);
and U8089 (N_8089,N_6332,N_5502);
nor U8090 (N_8090,N_6936,N_5674);
nand U8091 (N_8091,N_6176,N_7475);
nor U8092 (N_8092,N_6982,N_7081);
nor U8093 (N_8093,N_7126,N_5321);
nand U8094 (N_8094,N_7349,N_6037);
or U8095 (N_8095,N_5023,N_6113);
nand U8096 (N_8096,N_5558,N_5693);
or U8097 (N_8097,N_6919,N_5736);
and U8098 (N_8098,N_5104,N_5945);
nor U8099 (N_8099,N_6921,N_6988);
nor U8100 (N_8100,N_5575,N_6361);
nand U8101 (N_8101,N_7412,N_6835);
nor U8102 (N_8102,N_5800,N_6577);
and U8103 (N_8103,N_7227,N_5910);
and U8104 (N_8104,N_6915,N_5909);
or U8105 (N_8105,N_5485,N_6612);
or U8106 (N_8106,N_6604,N_7458);
and U8107 (N_8107,N_6178,N_6675);
or U8108 (N_8108,N_6641,N_6813);
nor U8109 (N_8109,N_7231,N_6857);
nor U8110 (N_8110,N_6694,N_5832);
nand U8111 (N_8111,N_5213,N_5662);
and U8112 (N_8112,N_6309,N_5750);
nand U8113 (N_8113,N_6226,N_5768);
nand U8114 (N_8114,N_7498,N_5072);
or U8115 (N_8115,N_5130,N_5151);
xor U8116 (N_8116,N_7210,N_7277);
or U8117 (N_8117,N_5225,N_6287);
nor U8118 (N_8118,N_7468,N_5354);
or U8119 (N_8119,N_6508,N_5064);
nor U8120 (N_8120,N_6816,N_5946);
nor U8121 (N_8121,N_5831,N_5511);
nor U8122 (N_8122,N_6024,N_7399);
or U8123 (N_8123,N_7178,N_5039);
or U8124 (N_8124,N_5643,N_7076);
and U8125 (N_8125,N_6028,N_6513);
or U8126 (N_8126,N_6622,N_5481);
nand U8127 (N_8127,N_5638,N_6793);
or U8128 (N_8128,N_5427,N_5872);
nor U8129 (N_8129,N_6644,N_7240);
nand U8130 (N_8130,N_5729,N_6033);
nand U8131 (N_8131,N_6776,N_6910);
nor U8132 (N_8132,N_6985,N_6184);
nor U8133 (N_8133,N_5879,N_6601);
and U8134 (N_8134,N_6680,N_7153);
nand U8135 (N_8135,N_6560,N_6022);
nor U8136 (N_8136,N_5076,N_7041);
nor U8137 (N_8137,N_5080,N_6370);
or U8138 (N_8138,N_6850,N_5707);
nand U8139 (N_8139,N_5363,N_7049);
and U8140 (N_8140,N_5737,N_6645);
nand U8141 (N_8141,N_6864,N_7140);
and U8142 (N_8142,N_6902,N_5230);
nor U8143 (N_8143,N_5397,N_5120);
or U8144 (N_8144,N_6170,N_7422);
or U8145 (N_8145,N_7258,N_5943);
and U8146 (N_8146,N_6268,N_5260);
and U8147 (N_8147,N_7008,N_6928);
or U8148 (N_8148,N_7450,N_6132);
nand U8149 (N_8149,N_5222,N_6841);
and U8150 (N_8150,N_7026,N_6222);
and U8151 (N_8151,N_5357,N_5417);
or U8152 (N_8152,N_7282,N_7372);
and U8153 (N_8153,N_6958,N_6532);
or U8154 (N_8154,N_7053,N_6059);
nor U8155 (N_8155,N_5754,N_7132);
or U8156 (N_8156,N_5862,N_5974);
nor U8157 (N_8157,N_5970,N_5244);
and U8158 (N_8158,N_5067,N_6286);
nor U8159 (N_8159,N_5786,N_7480);
or U8160 (N_8160,N_5258,N_6678);
nor U8161 (N_8161,N_6784,N_5670);
or U8162 (N_8162,N_6448,N_5467);
nand U8163 (N_8163,N_7225,N_5904);
and U8164 (N_8164,N_5775,N_6738);
nand U8165 (N_8165,N_6192,N_6515);
nor U8166 (N_8166,N_6423,N_7429);
nor U8167 (N_8167,N_7292,N_5471);
or U8168 (N_8168,N_5408,N_6262);
or U8169 (N_8169,N_7409,N_5922);
or U8170 (N_8170,N_5874,N_6386);
or U8171 (N_8171,N_5364,N_6851);
or U8172 (N_8172,N_7418,N_5082);
and U8173 (N_8173,N_7402,N_5000);
and U8174 (N_8174,N_7102,N_6610);
nand U8175 (N_8175,N_6732,N_5992);
and U8176 (N_8176,N_5220,N_5671);
and U8177 (N_8177,N_6038,N_5756);
and U8178 (N_8178,N_5999,N_7072);
nor U8179 (N_8179,N_7090,N_6435);
nand U8180 (N_8180,N_7223,N_6963);
or U8181 (N_8181,N_5369,N_6086);
and U8182 (N_8182,N_5595,N_6672);
or U8183 (N_8183,N_6103,N_5202);
or U8184 (N_8184,N_6674,N_6840);
nor U8185 (N_8185,N_6964,N_6745);
nor U8186 (N_8186,N_5098,N_6180);
and U8187 (N_8187,N_7309,N_6911);
and U8188 (N_8188,N_5869,N_5883);
nor U8189 (N_8189,N_5543,N_6040);
nand U8190 (N_8190,N_5117,N_5395);
and U8191 (N_8191,N_6229,N_5979);
or U8192 (N_8192,N_5975,N_7226);
and U8193 (N_8193,N_6885,N_6085);
nor U8194 (N_8194,N_6255,N_5107);
and U8195 (N_8195,N_5070,N_5818);
or U8196 (N_8196,N_5040,N_6896);
and U8197 (N_8197,N_5789,N_7143);
nor U8198 (N_8198,N_6317,N_5353);
nor U8199 (N_8199,N_6414,N_6173);
nand U8200 (N_8200,N_5571,N_5183);
nand U8201 (N_8201,N_5012,N_7428);
or U8202 (N_8202,N_6990,N_5283);
and U8203 (N_8203,N_7466,N_5718);
or U8204 (N_8204,N_7383,N_6236);
nor U8205 (N_8205,N_6131,N_6753);
nand U8206 (N_8206,N_7376,N_5483);
nor U8207 (N_8207,N_7024,N_5150);
or U8208 (N_8208,N_7330,N_7353);
nor U8209 (N_8209,N_7131,N_5439);
nand U8210 (N_8210,N_6631,N_5905);
nor U8211 (N_8211,N_5413,N_5016);
or U8212 (N_8212,N_5664,N_5133);
nand U8213 (N_8213,N_5841,N_6153);
and U8214 (N_8214,N_5762,N_6710);
and U8215 (N_8215,N_6526,N_6122);
nor U8216 (N_8216,N_7368,N_6125);
and U8217 (N_8217,N_5968,N_7245);
nor U8218 (N_8218,N_6213,N_7016);
nand U8219 (N_8219,N_6218,N_6401);
nand U8220 (N_8220,N_6331,N_7388);
or U8221 (N_8221,N_5913,N_6021);
nor U8222 (N_8222,N_5494,N_7324);
nand U8223 (N_8223,N_6818,N_6726);
or U8224 (N_8224,N_5160,N_6986);
nand U8225 (N_8225,N_6116,N_6979);
nand U8226 (N_8226,N_5297,N_7478);
or U8227 (N_8227,N_6825,N_6202);
nor U8228 (N_8228,N_5618,N_5496);
or U8229 (N_8229,N_6977,N_5644);
or U8230 (N_8230,N_7241,N_6965);
nor U8231 (N_8231,N_5277,N_7017);
nor U8232 (N_8232,N_6060,N_6993);
or U8233 (N_8233,N_5447,N_5073);
nand U8234 (N_8234,N_5328,N_5803);
or U8235 (N_8235,N_5991,N_6091);
nor U8236 (N_8236,N_6108,N_6432);
and U8237 (N_8237,N_6296,N_7426);
and U8238 (N_8238,N_7385,N_6183);
and U8239 (N_8239,N_6294,N_6984);
xnor U8240 (N_8240,N_6600,N_6274);
or U8241 (N_8241,N_5555,N_7489);
or U8242 (N_8242,N_5383,N_5723);
nor U8243 (N_8243,N_5977,N_7393);
xor U8244 (N_8244,N_5102,N_7472);
and U8245 (N_8245,N_5498,N_7148);
or U8246 (N_8246,N_6129,N_6454);
nor U8247 (N_8247,N_6077,N_6397);
nor U8248 (N_8248,N_6823,N_5976);
nor U8249 (N_8249,N_6013,N_5242);
nor U8250 (N_8250,N_7354,N_6892);
and U8251 (N_8251,N_6330,N_6939);
nor U8252 (N_8252,N_7037,N_5785);
or U8253 (N_8253,N_6883,N_7268);
nand U8254 (N_8254,N_6900,N_6426);
nor U8255 (N_8255,N_5344,N_7462);
and U8256 (N_8256,N_6580,N_7356);
or U8257 (N_8257,N_5512,N_5599);
nor U8258 (N_8258,N_5466,N_6673);
or U8259 (N_8259,N_6269,N_7395);
or U8260 (N_8260,N_5896,N_5801);
nor U8261 (N_8261,N_5464,N_5229);
nand U8262 (N_8262,N_6372,N_5523);
nand U8263 (N_8263,N_5669,N_5663);
or U8264 (N_8264,N_7042,N_5563);
nand U8265 (N_8265,N_5760,N_6660);
nor U8266 (N_8266,N_5682,N_6695);
nor U8267 (N_8267,N_6930,N_5338);
nor U8268 (N_8268,N_7214,N_7404);
nand U8269 (N_8269,N_5489,N_6306);
nor U8270 (N_8270,N_5219,N_7054);
or U8271 (N_8271,N_5683,N_5717);
nand U8272 (N_8272,N_5161,N_5374);
nand U8273 (N_8273,N_7043,N_6112);
nor U8274 (N_8274,N_6757,N_6830);
or U8275 (N_8275,N_6529,N_5381);
and U8276 (N_8276,N_6787,N_7471);
nor U8277 (N_8277,N_5315,N_6462);
or U8278 (N_8278,N_6158,N_7167);
nor U8279 (N_8279,N_6693,N_6408);
nor U8280 (N_8280,N_5182,N_5462);
and U8281 (N_8281,N_6358,N_7299);
or U8282 (N_8282,N_5790,N_6895);
or U8283 (N_8283,N_6554,N_5079);
nand U8284 (N_8284,N_6733,N_6847);
nor U8285 (N_8285,N_7093,N_6898);
nor U8286 (N_8286,N_7347,N_7476);
or U8287 (N_8287,N_6231,N_6797);
and U8288 (N_8288,N_7311,N_5687);
nor U8289 (N_8289,N_5055,N_6257);
nor U8290 (N_8290,N_6530,N_6613);
nand U8291 (N_8291,N_6832,N_5216);
nor U8292 (N_8292,N_5647,N_5566);
nor U8293 (N_8293,N_5924,N_5232);
nand U8294 (N_8294,N_5365,N_6295);
nor U8295 (N_8295,N_5889,N_6181);
nand U8296 (N_8296,N_5050,N_6512);
or U8297 (N_8297,N_5516,N_6692);
nand U8298 (N_8298,N_6731,N_7326);
and U8299 (N_8299,N_5047,N_5593);
nand U8300 (N_8300,N_6078,N_5823);
nand U8301 (N_8301,N_6621,N_5743);
nor U8302 (N_8302,N_5958,N_5686);
nand U8303 (N_8303,N_7413,N_5813);
and U8304 (N_8304,N_5947,N_7338);
nor U8305 (N_8305,N_6254,N_7215);
nor U8306 (N_8306,N_6539,N_5997);
nand U8307 (N_8307,N_6853,N_6369);
or U8308 (N_8308,N_5137,N_5403);
nand U8309 (N_8309,N_6555,N_7433);
nor U8310 (N_8310,N_6000,N_5678);
nand U8311 (N_8311,N_7387,N_6593);
and U8312 (N_8312,N_6215,N_7484);
and U8313 (N_8313,N_5884,N_6495);
and U8314 (N_8314,N_5806,N_5592);
and U8315 (N_8315,N_5981,N_7177);
nand U8316 (N_8316,N_5379,N_6074);
and U8317 (N_8317,N_5672,N_6534);
and U8318 (N_8318,N_5291,N_6339);
or U8319 (N_8319,N_5187,N_6389);
nand U8320 (N_8320,N_7255,N_5937);
nor U8321 (N_8321,N_6474,N_5028);
or U8322 (N_8322,N_6966,N_5829);
nor U8323 (N_8323,N_5308,N_7119);
nand U8324 (N_8324,N_5011,N_6259);
nand U8325 (N_8325,N_6424,N_6950);
nor U8326 (N_8326,N_6410,N_7261);
and U8327 (N_8327,N_7423,N_5843);
nand U8328 (N_8328,N_5296,N_5627);
nand U8329 (N_8329,N_6962,N_6088);
nor U8330 (N_8330,N_6493,N_5215);
nand U8331 (N_8331,N_5772,N_6198);
or U8332 (N_8332,N_5355,N_7486);
or U8333 (N_8333,N_6200,N_5809);
nand U8334 (N_8334,N_5585,N_6207);
nand U8335 (N_8335,N_7253,N_6058);
or U8336 (N_8336,N_5522,N_5506);
or U8337 (N_8337,N_6421,N_7003);
and U8338 (N_8338,N_6803,N_7263);
or U8339 (N_8339,N_6054,N_7317);
nor U8340 (N_8340,N_5757,N_6499);
nand U8341 (N_8341,N_6953,N_6728);
or U8342 (N_8342,N_6338,N_6698);
or U8343 (N_8343,N_5207,N_5853);
nand U8344 (N_8344,N_6705,N_6276);
and U8345 (N_8345,N_7048,N_5454);
nor U8346 (N_8346,N_5551,N_5121);
and U8347 (N_8347,N_7477,N_7022);
nor U8348 (N_8348,N_5895,N_7397);
nor U8349 (N_8349,N_7088,N_5594);
and U8350 (N_8350,N_7329,N_6159);
or U8351 (N_8351,N_5152,N_6148);
nor U8352 (N_8352,N_6069,N_7271);
nor U8353 (N_8353,N_5368,N_5661);
nand U8354 (N_8354,N_7312,N_5951);
nand U8355 (N_8355,N_7348,N_7424);
nor U8356 (N_8356,N_5433,N_6398);
and U8357 (N_8357,N_7230,N_6790);
and U8358 (N_8358,N_6193,N_6019);
and U8359 (N_8359,N_5468,N_5435);
and U8360 (N_8360,N_5097,N_6788);
nand U8361 (N_8361,N_7146,N_5478);
nand U8362 (N_8362,N_7453,N_5766);
or U8363 (N_8363,N_5253,N_5596);
or U8364 (N_8364,N_5899,N_6690);
nor U8365 (N_8365,N_5366,N_5063);
and U8366 (N_8366,N_7345,N_5143);
or U8367 (N_8367,N_6413,N_7289);
and U8368 (N_8368,N_7232,N_6364);
and U8369 (N_8369,N_5835,N_6671);
or U8370 (N_8370,N_7044,N_6152);
and U8371 (N_8371,N_5332,N_6722);
or U8372 (N_8372,N_6632,N_7364);
nor U8373 (N_8373,N_5739,N_7014);
and U8374 (N_8374,N_7288,N_6638);
or U8375 (N_8375,N_6500,N_5475);
nand U8376 (N_8376,N_5941,N_6649);
or U8377 (N_8377,N_6981,N_5635);
nor U8378 (N_8378,N_6223,N_5141);
and U8379 (N_8379,N_6582,N_6187);
or U8380 (N_8380,N_6182,N_6025);
and U8381 (N_8381,N_6051,N_7279);
and U8382 (N_8382,N_6134,N_5389);
nor U8383 (N_8383,N_5573,N_5748);
and U8384 (N_8384,N_5953,N_5049);
and U8385 (N_8385,N_5263,N_7125);
nor U8386 (N_8386,N_7052,N_5944);
nor U8387 (N_8387,N_6079,N_5378);
and U8388 (N_8388,N_6639,N_6303);
and U8389 (N_8389,N_5264,N_7092);
or U8390 (N_8390,N_5912,N_6623);
or U8391 (N_8391,N_6498,N_5771);
nor U8392 (N_8392,N_5956,N_5541);
and U8393 (N_8393,N_6824,N_5940);
and U8394 (N_8394,N_7333,N_5658);
nand U8395 (N_8395,N_6716,N_6783);
nand U8396 (N_8396,N_6120,N_6619);
or U8397 (N_8397,N_7398,N_6130);
and U8398 (N_8398,N_6063,N_5314);
or U8399 (N_8399,N_6901,N_5303);
nor U8400 (N_8400,N_5436,N_5236);
nand U8401 (N_8401,N_5487,N_6390);
or U8402 (N_8402,N_5268,N_5156);
nor U8403 (N_8403,N_7390,N_6396);
nor U8404 (N_8404,N_6630,N_6647);
and U8405 (N_8405,N_5602,N_5892);
nand U8406 (N_8406,N_6760,N_6730);
xor U8407 (N_8407,N_6133,N_5025);
and U8408 (N_8408,N_5804,N_7009);
and U8409 (N_8409,N_5580,N_5302);
and U8410 (N_8410,N_7203,N_5325);
nand U8411 (N_8411,N_5484,N_6704);
and U8412 (N_8412,N_7401,N_5983);
and U8413 (N_8413,N_7047,N_6870);
nand U8414 (N_8414,N_6016,N_5059);
or U8415 (N_8415,N_5139,N_5890);
and U8416 (N_8416,N_7216,N_5044);
nand U8417 (N_8417,N_7099,N_5927);
xnor U8418 (N_8418,N_5902,N_6721);
nand U8419 (N_8419,N_7439,N_6289);
nand U8420 (N_8420,N_5346,N_6422);
nor U8421 (N_8421,N_5266,N_7010);
nor U8422 (N_8422,N_5985,N_7421);
and U8423 (N_8423,N_6406,N_5119);
nand U8424 (N_8424,N_5189,N_6844);
and U8425 (N_8425,N_5713,N_7355);
or U8426 (N_8426,N_5652,N_6681);
and U8427 (N_8427,N_6064,N_7086);
xor U8428 (N_8428,N_6828,N_6568);
and U8429 (N_8429,N_6677,N_6634);
or U8430 (N_8430,N_6863,N_5919);
nor U8431 (N_8431,N_6009,N_6035);
or U8432 (N_8432,N_6003,N_5681);
and U8433 (N_8433,N_6205,N_6865);
nor U8434 (N_8434,N_6597,N_6322);
and U8435 (N_8435,N_6503,N_7161);
nand U8436 (N_8436,N_6536,N_5493);
and U8437 (N_8437,N_7341,N_5262);
nand U8438 (N_8438,N_7190,N_6579);
and U8439 (N_8439,N_5256,N_5452);
nand U8440 (N_8440,N_6770,N_5398);
and U8441 (N_8441,N_6427,N_5155);
nor U8442 (N_8442,N_7113,N_5851);
and U8443 (N_8443,N_6897,N_6650);
nand U8444 (N_8444,N_6168,N_5145);
and U8445 (N_8445,N_7359,N_6544);
xor U8446 (N_8446,N_5709,N_7377);
nand U8447 (N_8447,N_5367,N_6501);
nand U8448 (N_8448,N_6636,N_5962);
nor U8449 (N_8449,N_6418,N_5250);
or U8450 (N_8450,N_6992,N_5581);
xnor U8451 (N_8451,N_6382,N_5311);
or U8452 (N_8452,N_5834,N_5347);
nor U8453 (N_8453,N_6050,N_6801);
nor U8454 (N_8454,N_7275,N_5702);
and U8455 (N_8455,N_5200,N_6004);
nor U8456 (N_8456,N_5324,N_5608);
nand U8457 (N_8457,N_6041,N_6376);
and U8458 (N_8458,N_5190,N_5532);
nand U8459 (N_8459,N_6224,N_5852);
and U8460 (N_8460,N_7257,N_5045);
or U8461 (N_8461,N_6030,N_7018);
or U8462 (N_8462,N_5443,N_6876);
and U8463 (N_8463,N_5817,N_7020);
or U8464 (N_8464,N_7386,N_6325);
nand U8465 (N_8465,N_6781,N_5959);
nor U8466 (N_8466,N_5617,N_7343);
or U8467 (N_8467,N_7036,N_5174);
nand U8468 (N_8468,N_6438,N_6150);
or U8469 (N_8469,N_5850,N_5382);
and U8470 (N_8470,N_7023,N_5727);
nor U8471 (N_8471,N_5808,N_6098);
nor U8472 (N_8472,N_5918,N_6867);
or U8473 (N_8473,N_7172,N_6719);
and U8474 (N_8474,N_5623,N_5096);
or U8475 (N_8475,N_6023,N_6359);
and U8476 (N_8476,N_5083,N_7313);
nor U8477 (N_8477,N_7168,N_6209);
and U8478 (N_8478,N_6228,N_7187);
xnor U8479 (N_8479,N_5265,N_7115);
and U8480 (N_8480,N_5865,N_7389);
nor U8481 (N_8481,N_6208,N_6798);
nor U8482 (N_8482,N_6195,N_6846);
nand U8483 (N_8483,N_6258,N_6775);
nor U8484 (N_8484,N_6097,N_7059);
nand U8485 (N_8485,N_6106,N_6011);
and U8486 (N_8486,N_6802,N_6922);
nand U8487 (N_8487,N_5684,N_5657);
and U8488 (N_8488,N_7001,N_6012);
or U8489 (N_8489,N_7331,N_5569);
and U8490 (N_8490,N_6018,N_7482);
nand U8491 (N_8491,N_7460,N_6535);
nand U8492 (N_8492,N_6570,N_6337);
nor U8493 (N_8493,N_5472,N_7176);
nand U8494 (N_8494,N_5327,N_5140);
nor U8495 (N_8495,N_6280,N_6466);
nand U8496 (N_8496,N_5093,N_6505);
nor U8497 (N_8497,N_6511,N_6347);
nor U8498 (N_8498,N_5214,N_6310);
nand U8499 (N_8499,N_6026,N_7392);
nor U8500 (N_8500,N_5561,N_5091);
and U8501 (N_8501,N_5223,N_5996);
and U8502 (N_8502,N_6017,N_5375);
and U8503 (N_8503,N_5898,N_7074);
or U8504 (N_8504,N_5966,N_7152);
and U8505 (N_8505,N_6602,N_5849);
nor U8506 (N_8506,N_6658,N_5103);
nand U8507 (N_8507,N_5401,N_6428);
and U8508 (N_8508,N_7170,N_6267);
nand U8509 (N_8509,N_6651,N_7191);
nand U8510 (N_8510,N_6293,N_6080);
and U8511 (N_8511,N_6301,N_5673);
nand U8512 (N_8512,N_7425,N_6480);
nor U8513 (N_8513,N_5914,N_7320);
nand U8514 (N_8514,N_7459,N_7485);
or U8515 (N_8515,N_5517,N_6891);
and U8516 (N_8516,N_7479,N_7272);
nand U8517 (N_8517,N_5590,N_5360);
nand U8518 (N_8518,N_6360,N_6135);
or U8519 (N_8519,N_5568,N_7015);
nor U8520 (N_8520,N_6595,N_5406);
nand U8521 (N_8521,N_6328,N_7351);
nand U8522 (N_8522,N_5778,N_7391);
nor U8523 (N_8523,N_5931,N_5288);
nand U8524 (N_8524,N_5342,N_6742);
nor U8525 (N_8525,N_5146,N_5553);
nand U8526 (N_8526,N_7491,N_6449);
nand U8527 (N_8527,N_6177,N_5986);
or U8528 (N_8528,N_6238,N_6239);
nand U8529 (N_8529,N_5508,N_6138);
nor U8530 (N_8530,N_5175,N_5885);
or U8531 (N_8531,N_5351,N_6439);
or U8532 (N_8532,N_5390,N_5316);
nand U8533 (N_8533,N_6166,N_5138);
or U8534 (N_8534,N_5839,N_5777);
and U8535 (N_8535,N_5633,N_5078);
nor U8536 (N_8536,N_5352,N_5243);
nor U8537 (N_8537,N_5114,N_5275);
or U8538 (N_8538,N_6765,N_5415);
and U8539 (N_8539,N_7316,N_6578);
nand U8540 (N_8540,N_6820,N_6652);
and U8541 (N_8541,N_7266,N_5430);
nor U8542 (N_8542,N_5335,N_6118);
nand U8543 (N_8543,N_6140,N_7366);
and U8544 (N_8544,N_7050,N_6583);
nand U8545 (N_8545,N_5217,N_5031);
and U8546 (N_8546,N_5787,N_6914);
nor U8547 (N_8547,N_6826,N_5721);
and U8548 (N_8548,N_5339,N_5043);
nand U8549 (N_8549,N_5088,N_5971);
and U8550 (N_8550,N_7029,N_6321);
or U8551 (N_8551,N_6288,N_6750);
nand U8552 (N_8552,N_5694,N_6460);
and U8553 (N_8553,N_5715,N_5431);
nand U8554 (N_8554,N_7128,N_5963);
nor U8555 (N_8555,N_5921,N_6124);
nor U8556 (N_8556,N_7408,N_5270);
nor U8557 (N_8557,N_7028,N_5587);
nand U8558 (N_8558,N_6350,N_5688);
nand U8559 (N_8559,N_6283,N_5878);
and U8560 (N_8560,N_5090,N_6758);
nand U8561 (N_8561,N_6189,N_6379);
nand U8562 (N_8562,N_5411,N_6718);
nand U8563 (N_8563,N_5033,N_6665);
nand U8564 (N_8564,N_7247,N_6564);
nor U8565 (N_8565,N_7021,N_6279);
or U8566 (N_8566,N_5157,N_5877);
nor U8567 (N_8567,N_6754,N_6947);
and U8568 (N_8568,N_6042,N_5989);
nand U8569 (N_8569,N_5159,N_5370);
nand U8570 (N_8570,N_5961,N_7106);
and U8571 (N_8571,N_6362,N_5668);
nor U8572 (N_8572,N_6128,N_5309);
nor U8573 (N_8573,N_6093,N_6893);
nor U8574 (N_8574,N_6586,N_6145);
nor U8575 (N_8575,N_6142,N_5881);
or U8576 (N_8576,N_5738,N_7220);
nand U8577 (N_8577,N_7057,N_6453);
or U8578 (N_8578,N_6952,N_6860);
nor U8579 (N_8579,N_6685,N_6587);
nand U8580 (N_8580,N_5783,N_7357);
and U8581 (N_8581,N_5170,N_6837);
and U8582 (N_8582,N_5607,N_6743);
and U8583 (N_8583,N_6210,N_7414);
or U8584 (N_8584,N_5387,N_7286);
and U8585 (N_8585,N_6109,N_6160);
nand U8586 (N_8586,N_5842,N_5176);
or U8587 (N_8587,N_5171,N_7344);
and U8588 (N_8588,N_5248,N_6807);
or U8589 (N_8589,N_6717,N_6618);
or U8590 (N_8590,N_5255,N_6032);
nand U8591 (N_8591,N_7280,N_7381);
nor U8592 (N_8592,N_6916,N_5542);
and U8593 (N_8593,N_5836,N_7416);
and U8594 (N_8594,N_6547,N_6744);
or U8595 (N_8595,N_6245,N_6489);
or U8596 (N_8596,N_6909,N_6319);
nor U8597 (N_8597,N_6629,N_6491);
or U8598 (N_8598,N_6766,N_5423);
nand U8599 (N_8599,N_6027,N_6504);
nor U8600 (N_8600,N_5125,N_5935);
nor U8601 (N_8601,N_6811,N_6567);
and U8602 (N_8602,N_7032,N_7339);
nor U8603 (N_8603,N_7141,N_6102);
nand U8604 (N_8604,N_5348,N_5041);
or U8605 (N_8605,N_6541,N_5054);
or U8606 (N_8606,N_5428,N_6154);
nand U8607 (N_8607,N_5065,N_6903);
and U8608 (N_8608,N_6571,N_6737);
nor U8609 (N_8609,N_6175,N_7373);
nand U8610 (N_8610,N_5128,N_6216);
or U8611 (N_8611,N_5254,N_7350);
nor U8612 (N_8612,N_6882,N_6697);
nor U8613 (N_8613,N_5350,N_5886);
or U8614 (N_8614,N_6243,N_6800);
nand U8615 (N_8615,N_7157,N_6136);
nand U8616 (N_8616,N_7056,N_6497);
or U8617 (N_8617,N_6834,N_6938);
nor U8618 (N_8618,N_6071,N_6241);
and U8619 (N_8619,N_5651,N_5620);
and U8620 (N_8620,N_5445,N_7363);
nor U8621 (N_8621,N_6155,N_7370);
or U8622 (N_8622,N_6923,N_5429);
nand U8623 (N_8623,N_6908,N_5845);
nor U8624 (N_8624,N_5880,N_7457);
nor U8625 (N_8625,N_5636,N_6616);
nor U8626 (N_8626,N_6620,N_5386);
and U8627 (N_8627,N_5700,N_7079);
and U8628 (N_8628,N_6715,N_7180);
and U8629 (N_8629,N_6839,N_7293);
or U8630 (N_8630,N_5400,N_6927);
and U8631 (N_8631,N_6712,N_7004);
nor U8632 (N_8632,N_6980,N_5984);
and U8633 (N_8633,N_6352,N_5006);
xnor U8634 (N_8634,N_6594,N_7375);
and U8635 (N_8635,N_6221,N_6185);
nor U8636 (N_8636,N_6796,N_5969);
or U8637 (N_8637,N_6479,N_5795);
nor U8638 (N_8638,N_6349,N_5609);
or U8639 (N_8639,N_7441,N_5676);
or U8640 (N_8640,N_7325,N_7221);
and U8641 (N_8641,N_5295,N_6815);
nand U8642 (N_8642,N_5228,N_5875);
nor U8643 (N_8643,N_5463,N_6795);
nand U8644 (N_8644,N_5301,N_5577);
and U8645 (N_8645,N_5654,N_6917);
nand U8646 (N_8646,N_5689,N_6095);
or U8647 (N_8647,N_7335,N_7394);
or U8648 (N_8648,N_6772,N_5908);
or U8649 (N_8649,N_5237,N_6174);
nand U8650 (N_8650,N_7334,N_6502);
or U8651 (N_8651,N_6708,N_6886);
nor U8652 (N_8652,N_5234,N_6519);
nand U8653 (N_8653,N_7254,N_5557);
and U8654 (N_8654,N_6924,N_6627);
or U8655 (N_8655,N_6247,N_6679);
nand U8656 (N_8656,N_6383,N_6999);
nand U8657 (N_8657,N_5017,N_7078);
nor U8658 (N_8658,N_5685,N_5409);
and U8659 (N_8659,N_6273,N_6487);
nor U8660 (N_8660,N_5490,N_7287);
nand U8661 (N_8661,N_6053,N_7302);
nor U8662 (N_8662,N_6961,N_6115);
nor U8663 (N_8663,N_5118,N_5505);
nand U8664 (N_8664,N_6527,N_5235);
and U8665 (N_8665,N_5168,N_5089);
and U8666 (N_8666,N_6378,N_7006);
or U8667 (N_8667,N_6907,N_6878);
and U8668 (N_8668,N_7315,N_6203);
nand U8669 (N_8669,N_6117,N_7145);
nor U8670 (N_8670,N_5418,N_7189);
nor U8671 (N_8671,N_5666,N_5208);
xor U8672 (N_8672,N_5148,N_5340);
or U8673 (N_8673,N_5552,N_7129);
and U8674 (N_8674,N_5799,N_7487);
nand U8675 (N_8675,N_5421,N_6463);
nand U8676 (N_8676,N_6230,N_6196);
nand U8677 (N_8677,N_6739,N_5261);
or U8678 (N_8678,N_6126,N_7327);
and U8679 (N_8679,N_5692,N_5972);
nand U8680 (N_8680,N_6320,N_6637);
and U8681 (N_8681,N_6073,N_6299);
or U8682 (N_8682,N_5659,N_6521);
nand U8683 (N_8683,N_5203,N_6235);
and U8684 (N_8684,N_7233,N_6242);
nand U8685 (N_8685,N_5782,N_5826);
or U8686 (N_8686,N_5696,N_5520);
nor U8687 (N_8687,N_6282,N_6197);
or U8688 (N_8688,N_5952,N_7256);
and U8689 (N_8689,N_5559,N_6486);
nor U8690 (N_8690,N_7179,N_6047);
or U8691 (N_8691,N_6431,N_7005);
nor U8692 (N_8692,N_7108,N_7136);
nand U8693 (N_8693,N_6741,N_6092);
nor U8694 (N_8694,N_6523,N_6668);
or U8695 (N_8695,N_5714,N_6380);
nor U8696 (N_8696,N_6931,N_7103);
and U8697 (N_8697,N_6713,N_6667);
nand U8698 (N_8698,N_5020,N_5005);
nand U8699 (N_8699,N_6546,N_6700);
or U8700 (N_8700,N_7104,N_6817);
or U8701 (N_8701,N_5710,N_6956);
and U8702 (N_8702,N_5226,N_5259);
and U8703 (N_8703,N_5833,N_6994);
or U8704 (N_8704,N_6164,N_6407);
or U8705 (N_8705,N_5631,N_7369);
nor U8706 (N_8706,N_6165,N_6540);
nand U8707 (N_8707,N_5530,N_5084);
and U8708 (N_8708,N_5537,N_6008);
or U8709 (N_8709,N_6862,N_5758);
nor U8710 (N_8710,N_7419,N_6777);
nor U8711 (N_8711,N_5613,N_7437);
or U8712 (N_8712,N_6446,N_7495);
or U8713 (N_8713,N_6323,N_6005);
or U8714 (N_8714,N_5279,N_5246);
nor U8715 (N_8715,N_7211,N_6533);
nand U8716 (N_8716,N_6162,N_7025);
nor U8717 (N_8717,N_5154,N_6510);
nand U8718 (N_8718,N_5249,N_5773);
and U8719 (N_8719,N_7055,N_6791);
or U8720 (N_8720,N_7207,N_5855);
nand U8721 (N_8721,N_5438,N_7142);
and U8722 (N_8722,N_5863,N_6769);
nor U8723 (N_8723,N_7246,N_6838);
and U8724 (N_8724,N_5178,N_7012);
nor U8725 (N_8725,N_5805,N_6551);
and U8726 (N_8726,N_5173,N_7244);
or U8727 (N_8727,N_5196,N_5957);
or U8728 (N_8728,N_5724,N_7069);
or U8729 (N_8729,N_5518,N_7199);
nand U8730 (N_8730,N_5949,N_6537);
nand U8731 (N_8731,N_7116,N_6625);
nand U8732 (N_8732,N_6172,N_7109);
nor U8733 (N_8733,N_7030,N_7410);
or U8734 (N_8734,N_5867,N_7265);
nand U8735 (N_8735,N_6149,N_5699);
nor U8736 (N_8736,N_5860,N_5749);
nand U8737 (N_8737,N_6415,N_5449);
nor U8738 (N_8738,N_6686,N_6976);
nand U8739 (N_8739,N_6417,N_5473);
nor U8740 (N_8740,N_7465,N_5550);
nand U8741 (N_8741,N_5822,N_6201);
or U8742 (N_8742,N_7192,N_7209);
nand U8743 (N_8743,N_5450,N_5605);
or U8744 (N_8744,N_6696,N_6392);
or U8745 (N_8745,N_6854,N_7027);
nand U8746 (N_8746,N_5206,N_5361);
nor U8747 (N_8747,N_6391,N_6250);
nor U8748 (N_8748,N_6227,N_6263);
nor U8749 (N_8749,N_6326,N_6285);
nand U8750 (N_8750,N_6532,N_5737);
and U8751 (N_8751,N_6185,N_5939);
or U8752 (N_8752,N_6962,N_6974);
nand U8753 (N_8753,N_5053,N_5443);
and U8754 (N_8754,N_5535,N_6353);
nand U8755 (N_8755,N_6721,N_6797);
or U8756 (N_8756,N_6370,N_7261);
nand U8757 (N_8757,N_6771,N_7433);
and U8758 (N_8758,N_7044,N_5504);
nor U8759 (N_8759,N_6523,N_6320);
nand U8760 (N_8760,N_5533,N_6876);
nor U8761 (N_8761,N_7427,N_5977);
nand U8762 (N_8762,N_5583,N_5937);
or U8763 (N_8763,N_6791,N_5336);
or U8764 (N_8764,N_5790,N_6438);
and U8765 (N_8765,N_7367,N_5392);
or U8766 (N_8766,N_6736,N_6520);
nor U8767 (N_8767,N_6039,N_6395);
and U8768 (N_8768,N_7283,N_5421);
nor U8769 (N_8769,N_5380,N_5450);
nand U8770 (N_8770,N_5710,N_6110);
and U8771 (N_8771,N_6412,N_5228);
and U8772 (N_8772,N_5953,N_6273);
and U8773 (N_8773,N_6729,N_7202);
and U8774 (N_8774,N_6053,N_5826);
nor U8775 (N_8775,N_6726,N_5944);
nor U8776 (N_8776,N_5187,N_6722);
nand U8777 (N_8777,N_5959,N_6757);
and U8778 (N_8778,N_6711,N_5745);
nor U8779 (N_8779,N_7343,N_5106);
or U8780 (N_8780,N_7192,N_5543);
nand U8781 (N_8781,N_5319,N_7156);
nand U8782 (N_8782,N_7341,N_5040);
and U8783 (N_8783,N_7221,N_5182);
or U8784 (N_8784,N_5446,N_6389);
nand U8785 (N_8785,N_6989,N_6539);
nor U8786 (N_8786,N_6063,N_5077);
or U8787 (N_8787,N_5906,N_5452);
or U8788 (N_8788,N_6263,N_6978);
and U8789 (N_8789,N_6988,N_5952);
nor U8790 (N_8790,N_5122,N_7383);
nand U8791 (N_8791,N_5674,N_7180);
or U8792 (N_8792,N_5595,N_5013);
nor U8793 (N_8793,N_7484,N_5206);
or U8794 (N_8794,N_7186,N_6729);
nand U8795 (N_8795,N_5805,N_7460);
or U8796 (N_8796,N_5075,N_5944);
nor U8797 (N_8797,N_6230,N_7059);
nor U8798 (N_8798,N_6262,N_5427);
nand U8799 (N_8799,N_5304,N_6257);
nor U8800 (N_8800,N_7462,N_6844);
nand U8801 (N_8801,N_7469,N_7197);
or U8802 (N_8802,N_6676,N_6217);
nor U8803 (N_8803,N_5575,N_5322);
or U8804 (N_8804,N_6299,N_7125);
and U8805 (N_8805,N_5245,N_7181);
nor U8806 (N_8806,N_5015,N_7302);
or U8807 (N_8807,N_6373,N_6529);
or U8808 (N_8808,N_6350,N_5393);
nor U8809 (N_8809,N_5056,N_6191);
nand U8810 (N_8810,N_6249,N_5856);
or U8811 (N_8811,N_5283,N_6699);
nand U8812 (N_8812,N_5127,N_5368);
or U8813 (N_8813,N_5719,N_6189);
nor U8814 (N_8814,N_6012,N_5407);
nor U8815 (N_8815,N_6693,N_7003);
nand U8816 (N_8816,N_6764,N_7070);
or U8817 (N_8817,N_7219,N_5072);
and U8818 (N_8818,N_7355,N_5567);
nor U8819 (N_8819,N_5762,N_7455);
and U8820 (N_8820,N_5813,N_7005);
nor U8821 (N_8821,N_5156,N_7083);
nand U8822 (N_8822,N_6025,N_5064);
nand U8823 (N_8823,N_5867,N_5275);
nand U8824 (N_8824,N_6121,N_5736);
nand U8825 (N_8825,N_7475,N_5318);
nand U8826 (N_8826,N_6003,N_6558);
nor U8827 (N_8827,N_7103,N_5211);
nand U8828 (N_8828,N_5263,N_5839);
and U8829 (N_8829,N_6556,N_5150);
nor U8830 (N_8830,N_6750,N_7055);
or U8831 (N_8831,N_6124,N_6016);
nand U8832 (N_8832,N_5600,N_5696);
nor U8833 (N_8833,N_6379,N_7468);
and U8834 (N_8834,N_5339,N_6773);
or U8835 (N_8835,N_5425,N_6740);
xnor U8836 (N_8836,N_6617,N_6838);
or U8837 (N_8837,N_6217,N_6301);
or U8838 (N_8838,N_7095,N_6420);
and U8839 (N_8839,N_7180,N_5927);
nor U8840 (N_8840,N_5865,N_6094);
nor U8841 (N_8841,N_5481,N_5763);
and U8842 (N_8842,N_6112,N_5771);
or U8843 (N_8843,N_6048,N_6559);
nor U8844 (N_8844,N_6886,N_7004);
xor U8845 (N_8845,N_6321,N_6109);
nand U8846 (N_8846,N_6481,N_5331);
or U8847 (N_8847,N_7234,N_7249);
nand U8848 (N_8848,N_6333,N_7468);
nor U8849 (N_8849,N_6531,N_6701);
or U8850 (N_8850,N_5261,N_6954);
or U8851 (N_8851,N_6288,N_7255);
nor U8852 (N_8852,N_5549,N_5161);
and U8853 (N_8853,N_5863,N_6971);
nand U8854 (N_8854,N_7108,N_5299);
or U8855 (N_8855,N_6096,N_5211);
nor U8856 (N_8856,N_7257,N_6782);
and U8857 (N_8857,N_7406,N_5708);
and U8858 (N_8858,N_6915,N_5389);
xnor U8859 (N_8859,N_5930,N_5778);
nor U8860 (N_8860,N_6848,N_5647);
and U8861 (N_8861,N_7113,N_5974);
and U8862 (N_8862,N_5024,N_7439);
or U8863 (N_8863,N_6668,N_7421);
nor U8864 (N_8864,N_6823,N_6461);
nand U8865 (N_8865,N_5947,N_7089);
nor U8866 (N_8866,N_7478,N_5653);
nand U8867 (N_8867,N_5563,N_5726);
or U8868 (N_8868,N_5041,N_6094);
and U8869 (N_8869,N_6313,N_5846);
nand U8870 (N_8870,N_6013,N_5207);
or U8871 (N_8871,N_5931,N_5644);
or U8872 (N_8872,N_5752,N_6979);
or U8873 (N_8873,N_6254,N_5265);
nand U8874 (N_8874,N_6561,N_5788);
nand U8875 (N_8875,N_6105,N_5435);
and U8876 (N_8876,N_5977,N_7070);
or U8877 (N_8877,N_5829,N_5470);
and U8878 (N_8878,N_7249,N_6000);
nand U8879 (N_8879,N_5690,N_5035);
nand U8880 (N_8880,N_5720,N_6629);
and U8881 (N_8881,N_5535,N_5889);
xnor U8882 (N_8882,N_7224,N_5531);
and U8883 (N_8883,N_5767,N_6528);
nand U8884 (N_8884,N_6688,N_7207);
or U8885 (N_8885,N_6367,N_5323);
nand U8886 (N_8886,N_7025,N_6262);
and U8887 (N_8887,N_6036,N_5621);
nor U8888 (N_8888,N_7264,N_7187);
or U8889 (N_8889,N_5204,N_5392);
nand U8890 (N_8890,N_6475,N_5636);
nand U8891 (N_8891,N_5142,N_5394);
nand U8892 (N_8892,N_6647,N_6370);
nor U8893 (N_8893,N_7434,N_6142);
nand U8894 (N_8894,N_6933,N_5185);
nand U8895 (N_8895,N_5685,N_5303);
or U8896 (N_8896,N_5382,N_5411);
and U8897 (N_8897,N_6461,N_5617);
nor U8898 (N_8898,N_5314,N_7074);
nor U8899 (N_8899,N_6960,N_6841);
and U8900 (N_8900,N_6164,N_6084);
nor U8901 (N_8901,N_7483,N_6307);
and U8902 (N_8902,N_6951,N_7405);
and U8903 (N_8903,N_6065,N_6902);
nor U8904 (N_8904,N_5731,N_7458);
and U8905 (N_8905,N_6581,N_7391);
or U8906 (N_8906,N_7411,N_5174);
nor U8907 (N_8907,N_5280,N_6219);
and U8908 (N_8908,N_6155,N_7168);
nor U8909 (N_8909,N_7023,N_7261);
nand U8910 (N_8910,N_6347,N_5457);
or U8911 (N_8911,N_7287,N_7416);
nand U8912 (N_8912,N_6280,N_5493);
nand U8913 (N_8913,N_5192,N_5738);
and U8914 (N_8914,N_6415,N_7172);
nor U8915 (N_8915,N_6257,N_6892);
nor U8916 (N_8916,N_6470,N_7292);
nand U8917 (N_8917,N_6431,N_7074);
or U8918 (N_8918,N_5329,N_7239);
or U8919 (N_8919,N_5302,N_7147);
and U8920 (N_8920,N_6663,N_5909);
nor U8921 (N_8921,N_5148,N_7437);
and U8922 (N_8922,N_5915,N_6877);
or U8923 (N_8923,N_6302,N_5086);
or U8924 (N_8924,N_6487,N_5616);
nand U8925 (N_8925,N_6709,N_6839);
and U8926 (N_8926,N_5090,N_6365);
nor U8927 (N_8927,N_7492,N_6580);
or U8928 (N_8928,N_6963,N_7390);
nor U8929 (N_8929,N_5039,N_5984);
and U8930 (N_8930,N_6648,N_6420);
or U8931 (N_8931,N_5376,N_7319);
and U8932 (N_8932,N_5397,N_7345);
nand U8933 (N_8933,N_6616,N_5494);
nand U8934 (N_8934,N_6024,N_5990);
and U8935 (N_8935,N_5150,N_5712);
nand U8936 (N_8936,N_6558,N_7253);
or U8937 (N_8937,N_5786,N_5385);
nand U8938 (N_8938,N_5640,N_7063);
nand U8939 (N_8939,N_6271,N_6238);
and U8940 (N_8940,N_5572,N_7009);
nand U8941 (N_8941,N_5898,N_5354);
nand U8942 (N_8942,N_6761,N_6613);
nand U8943 (N_8943,N_6495,N_7374);
or U8944 (N_8944,N_6213,N_5450);
and U8945 (N_8945,N_6541,N_7042);
nand U8946 (N_8946,N_5002,N_5261);
nand U8947 (N_8947,N_6977,N_5896);
nor U8948 (N_8948,N_5624,N_5185);
or U8949 (N_8949,N_7402,N_7485);
or U8950 (N_8950,N_5185,N_7458);
or U8951 (N_8951,N_5696,N_5433);
nor U8952 (N_8952,N_5554,N_7082);
or U8953 (N_8953,N_6311,N_6211);
nor U8954 (N_8954,N_6556,N_6613);
nor U8955 (N_8955,N_5139,N_5405);
or U8956 (N_8956,N_6469,N_6581);
and U8957 (N_8957,N_7341,N_7146);
or U8958 (N_8958,N_6652,N_6341);
and U8959 (N_8959,N_7216,N_6333);
nand U8960 (N_8960,N_7082,N_5536);
and U8961 (N_8961,N_5977,N_6421);
nor U8962 (N_8962,N_6648,N_6694);
and U8963 (N_8963,N_7467,N_5946);
or U8964 (N_8964,N_7136,N_7225);
nor U8965 (N_8965,N_6739,N_6928);
or U8966 (N_8966,N_6814,N_7340);
and U8967 (N_8967,N_5573,N_6674);
and U8968 (N_8968,N_5682,N_5734);
or U8969 (N_8969,N_5623,N_5546);
and U8970 (N_8970,N_7322,N_6114);
and U8971 (N_8971,N_5348,N_7036);
nand U8972 (N_8972,N_5604,N_5738);
or U8973 (N_8973,N_7181,N_6452);
nor U8974 (N_8974,N_5053,N_5014);
nand U8975 (N_8975,N_5064,N_6389);
and U8976 (N_8976,N_5418,N_6523);
nor U8977 (N_8977,N_6790,N_7170);
or U8978 (N_8978,N_6117,N_7087);
and U8979 (N_8979,N_6371,N_5554);
nor U8980 (N_8980,N_7477,N_5243);
and U8981 (N_8981,N_6520,N_6876);
nand U8982 (N_8982,N_6050,N_6726);
and U8983 (N_8983,N_6872,N_6823);
nand U8984 (N_8984,N_5048,N_5900);
nand U8985 (N_8985,N_6192,N_6379);
and U8986 (N_8986,N_6998,N_5371);
nand U8987 (N_8987,N_7389,N_6295);
nand U8988 (N_8988,N_6786,N_5850);
nand U8989 (N_8989,N_6009,N_5299);
nand U8990 (N_8990,N_6113,N_5904);
nor U8991 (N_8991,N_7036,N_6709);
nor U8992 (N_8992,N_6353,N_6225);
or U8993 (N_8993,N_6415,N_7146);
or U8994 (N_8994,N_7034,N_7411);
nand U8995 (N_8995,N_5865,N_6714);
and U8996 (N_8996,N_7236,N_6031);
nand U8997 (N_8997,N_7192,N_6832);
nor U8998 (N_8998,N_5915,N_6297);
and U8999 (N_8999,N_6699,N_5733);
nand U9000 (N_9000,N_5273,N_6759);
nor U9001 (N_9001,N_7239,N_6659);
or U9002 (N_9002,N_7468,N_5852);
nor U9003 (N_9003,N_7026,N_5459);
nor U9004 (N_9004,N_5907,N_5473);
nand U9005 (N_9005,N_7281,N_5450);
nand U9006 (N_9006,N_6765,N_5121);
nand U9007 (N_9007,N_7184,N_5276);
nor U9008 (N_9008,N_6130,N_5881);
nor U9009 (N_9009,N_5106,N_6631);
and U9010 (N_9010,N_5995,N_5109);
nand U9011 (N_9011,N_6359,N_7412);
nor U9012 (N_9012,N_7048,N_5817);
and U9013 (N_9013,N_5724,N_5572);
and U9014 (N_9014,N_6376,N_5280);
or U9015 (N_9015,N_5110,N_5768);
or U9016 (N_9016,N_7144,N_5877);
and U9017 (N_9017,N_7015,N_5302);
nor U9018 (N_9018,N_5976,N_7015);
or U9019 (N_9019,N_7082,N_5960);
nand U9020 (N_9020,N_5949,N_5092);
and U9021 (N_9021,N_6256,N_5618);
nor U9022 (N_9022,N_7126,N_6336);
nor U9023 (N_9023,N_6159,N_5784);
and U9024 (N_9024,N_6190,N_7360);
and U9025 (N_9025,N_6704,N_6660);
nor U9026 (N_9026,N_6608,N_5052);
nor U9027 (N_9027,N_6933,N_5553);
nor U9028 (N_9028,N_5288,N_5920);
or U9029 (N_9029,N_5129,N_5620);
nor U9030 (N_9030,N_5686,N_5758);
nor U9031 (N_9031,N_6886,N_7017);
or U9032 (N_9032,N_6159,N_6314);
nand U9033 (N_9033,N_5428,N_7029);
or U9034 (N_9034,N_6363,N_6109);
or U9035 (N_9035,N_5747,N_5941);
and U9036 (N_9036,N_6032,N_5073);
nand U9037 (N_9037,N_5557,N_5412);
and U9038 (N_9038,N_7284,N_5941);
or U9039 (N_9039,N_6209,N_5271);
or U9040 (N_9040,N_5748,N_7089);
or U9041 (N_9041,N_5259,N_5669);
nand U9042 (N_9042,N_5469,N_5246);
nor U9043 (N_9043,N_6398,N_6890);
and U9044 (N_9044,N_5169,N_5396);
or U9045 (N_9045,N_5471,N_7388);
or U9046 (N_9046,N_6906,N_5037);
nand U9047 (N_9047,N_5883,N_6171);
nor U9048 (N_9048,N_7049,N_5143);
nor U9049 (N_9049,N_5383,N_7338);
and U9050 (N_9050,N_5887,N_6613);
nand U9051 (N_9051,N_5068,N_7356);
nor U9052 (N_9052,N_7027,N_6151);
or U9053 (N_9053,N_7400,N_6215);
nor U9054 (N_9054,N_5210,N_5488);
nor U9055 (N_9055,N_5614,N_6272);
nor U9056 (N_9056,N_7353,N_5669);
or U9057 (N_9057,N_5914,N_5287);
and U9058 (N_9058,N_5396,N_6222);
or U9059 (N_9059,N_6140,N_5352);
nor U9060 (N_9060,N_7254,N_5047);
nand U9061 (N_9061,N_5164,N_5377);
and U9062 (N_9062,N_5463,N_5575);
and U9063 (N_9063,N_6278,N_6066);
nand U9064 (N_9064,N_6577,N_5117);
nor U9065 (N_9065,N_5592,N_6475);
nand U9066 (N_9066,N_5325,N_7125);
xnor U9067 (N_9067,N_5196,N_6774);
or U9068 (N_9068,N_6769,N_5469);
and U9069 (N_9069,N_6756,N_5047);
nand U9070 (N_9070,N_7005,N_5927);
nand U9071 (N_9071,N_6629,N_5421);
and U9072 (N_9072,N_6885,N_7031);
xnor U9073 (N_9073,N_7307,N_6922);
nand U9074 (N_9074,N_6669,N_5073);
or U9075 (N_9075,N_6709,N_6898);
nand U9076 (N_9076,N_6208,N_5607);
and U9077 (N_9077,N_7329,N_5145);
and U9078 (N_9078,N_5905,N_6483);
or U9079 (N_9079,N_5886,N_6768);
or U9080 (N_9080,N_5696,N_6946);
nor U9081 (N_9081,N_7472,N_5097);
nand U9082 (N_9082,N_7088,N_5420);
or U9083 (N_9083,N_5619,N_6740);
nor U9084 (N_9084,N_6466,N_5916);
and U9085 (N_9085,N_5582,N_5406);
and U9086 (N_9086,N_7377,N_7479);
nand U9087 (N_9087,N_5501,N_5284);
nor U9088 (N_9088,N_6588,N_6486);
or U9089 (N_9089,N_5073,N_6247);
or U9090 (N_9090,N_5170,N_5707);
nor U9091 (N_9091,N_5583,N_6490);
and U9092 (N_9092,N_7272,N_6991);
or U9093 (N_9093,N_5875,N_6823);
nor U9094 (N_9094,N_5421,N_6120);
or U9095 (N_9095,N_5615,N_6590);
xor U9096 (N_9096,N_5369,N_6608);
and U9097 (N_9097,N_6480,N_5029);
and U9098 (N_9098,N_5971,N_6760);
nor U9099 (N_9099,N_5986,N_5709);
nand U9100 (N_9100,N_5469,N_6670);
or U9101 (N_9101,N_5133,N_5660);
xnor U9102 (N_9102,N_6028,N_5004);
and U9103 (N_9103,N_6559,N_5687);
or U9104 (N_9104,N_5749,N_7491);
nand U9105 (N_9105,N_5173,N_6257);
nand U9106 (N_9106,N_6238,N_7190);
or U9107 (N_9107,N_5802,N_5768);
nand U9108 (N_9108,N_6653,N_6229);
nand U9109 (N_9109,N_6215,N_5899);
and U9110 (N_9110,N_5709,N_6036);
and U9111 (N_9111,N_6628,N_5748);
nor U9112 (N_9112,N_5112,N_6397);
nand U9113 (N_9113,N_5021,N_5604);
xnor U9114 (N_9114,N_7489,N_7370);
and U9115 (N_9115,N_5509,N_6120);
nor U9116 (N_9116,N_7222,N_5253);
and U9117 (N_9117,N_5934,N_6474);
nor U9118 (N_9118,N_6904,N_6016);
or U9119 (N_9119,N_6259,N_5140);
and U9120 (N_9120,N_6201,N_6682);
nand U9121 (N_9121,N_7243,N_6935);
nor U9122 (N_9122,N_7103,N_6808);
and U9123 (N_9123,N_5130,N_7054);
nor U9124 (N_9124,N_6379,N_6112);
or U9125 (N_9125,N_5543,N_6579);
or U9126 (N_9126,N_6434,N_7173);
and U9127 (N_9127,N_5265,N_6717);
nor U9128 (N_9128,N_6512,N_6099);
nand U9129 (N_9129,N_5396,N_7325);
nor U9130 (N_9130,N_6529,N_5115);
nand U9131 (N_9131,N_7203,N_7260);
nor U9132 (N_9132,N_6746,N_5031);
and U9133 (N_9133,N_6943,N_5632);
or U9134 (N_9134,N_5299,N_5879);
and U9135 (N_9135,N_6741,N_6224);
nor U9136 (N_9136,N_5985,N_5929);
or U9137 (N_9137,N_6529,N_6041);
nor U9138 (N_9138,N_5300,N_5144);
and U9139 (N_9139,N_6233,N_5888);
or U9140 (N_9140,N_7416,N_6443);
nand U9141 (N_9141,N_6149,N_5165);
nor U9142 (N_9142,N_7176,N_5487);
nand U9143 (N_9143,N_7382,N_5227);
nor U9144 (N_9144,N_5672,N_6717);
nor U9145 (N_9145,N_5199,N_6698);
and U9146 (N_9146,N_6760,N_6080);
or U9147 (N_9147,N_5888,N_5490);
nand U9148 (N_9148,N_7263,N_7092);
nand U9149 (N_9149,N_7002,N_6642);
and U9150 (N_9150,N_6400,N_6114);
nand U9151 (N_9151,N_5352,N_5891);
nor U9152 (N_9152,N_6478,N_7376);
and U9153 (N_9153,N_5012,N_6507);
and U9154 (N_9154,N_6162,N_5919);
nand U9155 (N_9155,N_5067,N_7118);
or U9156 (N_9156,N_6361,N_6265);
or U9157 (N_9157,N_5178,N_7227);
or U9158 (N_9158,N_6904,N_6794);
nand U9159 (N_9159,N_6460,N_6721);
or U9160 (N_9160,N_5138,N_7126);
nor U9161 (N_9161,N_5800,N_5533);
and U9162 (N_9162,N_5060,N_5961);
and U9163 (N_9163,N_6026,N_7139);
nor U9164 (N_9164,N_6535,N_6397);
nor U9165 (N_9165,N_7200,N_6725);
and U9166 (N_9166,N_7069,N_7021);
nor U9167 (N_9167,N_5311,N_5622);
nand U9168 (N_9168,N_5835,N_5644);
nand U9169 (N_9169,N_6668,N_6591);
nand U9170 (N_9170,N_7479,N_5113);
or U9171 (N_9171,N_5163,N_5016);
nor U9172 (N_9172,N_6405,N_6429);
and U9173 (N_9173,N_7173,N_6167);
and U9174 (N_9174,N_6854,N_5836);
and U9175 (N_9175,N_5599,N_5422);
nand U9176 (N_9176,N_6464,N_6003);
nor U9177 (N_9177,N_7047,N_5345);
and U9178 (N_9178,N_7469,N_6060);
nand U9179 (N_9179,N_7336,N_7245);
and U9180 (N_9180,N_6067,N_5235);
and U9181 (N_9181,N_7261,N_5348);
and U9182 (N_9182,N_5976,N_6182);
or U9183 (N_9183,N_6318,N_5604);
or U9184 (N_9184,N_5426,N_6510);
or U9185 (N_9185,N_5290,N_7042);
and U9186 (N_9186,N_6639,N_6459);
nand U9187 (N_9187,N_6373,N_5479);
nand U9188 (N_9188,N_7080,N_6054);
or U9189 (N_9189,N_6517,N_5291);
and U9190 (N_9190,N_5482,N_6443);
nand U9191 (N_9191,N_7494,N_6525);
nor U9192 (N_9192,N_5627,N_5047);
and U9193 (N_9193,N_7176,N_7103);
or U9194 (N_9194,N_5711,N_6522);
and U9195 (N_9195,N_6169,N_5006);
nand U9196 (N_9196,N_7301,N_6999);
or U9197 (N_9197,N_6582,N_5460);
and U9198 (N_9198,N_6256,N_6650);
or U9199 (N_9199,N_5057,N_7182);
nor U9200 (N_9200,N_6371,N_7288);
nor U9201 (N_9201,N_5689,N_5141);
nand U9202 (N_9202,N_5607,N_5167);
and U9203 (N_9203,N_5634,N_5691);
nand U9204 (N_9204,N_6490,N_7425);
and U9205 (N_9205,N_6549,N_6295);
nor U9206 (N_9206,N_5831,N_6005);
nor U9207 (N_9207,N_7214,N_5077);
and U9208 (N_9208,N_5629,N_5498);
nor U9209 (N_9209,N_5076,N_7435);
nor U9210 (N_9210,N_6885,N_5412);
nand U9211 (N_9211,N_5398,N_6599);
and U9212 (N_9212,N_5825,N_6181);
and U9213 (N_9213,N_7012,N_6948);
or U9214 (N_9214,N_6305,N_7376);
or U9215 (N_9215,N_6702,N_6683);
nand U9216 (N_9216,N_6224,N_5006);
nand U9217 (N_9217,N_5617,N_5504);
and U9218 (N_9218,N_7170,N_6202);
or U9219 (N_9219,N_7116,N_6025);
nand U9220 (N_9220,N_5567,N_5576);
nor U9221 (N_9221,N_5906,N_5868);
xor U9222 (N_9222,N_5150,N_6772);
nor U9223 (N_9223,N_6869,N_5795);
and U9224 (N_9224,N_6030,N_5659);
nand U9225 (N_9225,N_5985,N_6423);
nand U9226 (N_9226,N_5904,N_6007);
and U9227 (N_9227,N_5151,N_6999);
nand U9228 (N_9228,N_6167,N_6887);
or U9229 (N_9229,N_6362,N_5473);
or U9230 (N_9230,N_5449,N_5985);
or U9231 (N_9231,N_7142,N_6511);
nand U9232 (N_9232,N_6506,N_5324);
and U9233 (N_9233,N_6922,N_6364);
nand U9234 (N_9234,N_6708,N_5063);
or U9235 (N_9235,N_7244,N_6023);
or U9236 (N_9236,N_5196,N_7142);
nor U9237 (N_9237,N_6972,N_6564);
nand U9238 (N_9238,N_5109,N_6993);
or U9239 (N_9239,N_5053,N_5263);
nor U9240 (N_9240,N_5395,N_5774);
and U9241 (N_9241,N_5097,N_5185);
and U9242 (N_9242,N_6094,N_6011);
nor U9243 (N_9243,N_5085,N_5658);
nand U9244 (N_9244,N_5307,N_5170);
and U9245 (N_9245,N_5974,N_5586);
and U9246 (N_9246,N_6965,N_5199);
or U9247 (N_9247,N_7067,N_5616);
or U9248 (N_9248,N_5292,N_7028);
nor U9249 (N_9249,N_5885,N_6385);
nand U9250 (N_9250,N_6484,N_5873);
and U9251 (N_9251,N_5272,N_6886);
and U9252 (N_9252,N_6541,N_5529);
nand U9253 (N_9253,N_7173,N_5634);
nand U9254 (N_9254,N_5195,N_5326);
or U9255 (N_9255,N_5172,N_6927);
nor U9256 (N_9256,N_5047,N_7251);
nand U9257 (N_9257,N_7256,N_5191);
or U9258 (N_9258,N_7462,N_6616);
nand U9259 (N_9259,N_6455,N_7427);
nand U9260 (N_9260,N_6098,N_6521);
and U9261 (N_9261,N_5449,N_6133);
nor U9262 (N_9262,N_5164,N_7263);
nor U9263 (N_9263,N_5662,N_5557);
nor U9264 (N_9264,N_5982,N_6811);
and U9265 (N_9265,N_6108,N_6036);
or U9266 (N_9266,N_5279,N_5288);
nor U9267 (N_9267,N_5655,N_5094);
or U9268 (N_9268,N_5251,N_6616);
and U9269 (N_9269,N_5344,N_6467);
nand U9270 (N_9270,N_5113,N_5869);
and U9271 (N_9271,N_6556,N_6084);
nand U9272 (N_9272,N_6591,N_6223);
and U9273 (N_9273,N_6747,N_6423);
and U9274 (N_9274,N_7270,N_7148);
nor U9275 (N_9275,N_5834,N_6594);
and U9276 (N_9276,N_6633,N_6768);
or U9277 (N_9277,N_6061,N_5204);
nor U9278 (N_9278,N_5687,N_6440);
nand U9279 (N_9279,N_5112,N_6816);
nor U9280 (N_9280,N_6011,N_7026);
nand U9281 (N_9281,N_5903,N_7089);
and U9282 (N_9282,N_7082,N_5507);
and U9283 (N_9283,N_6170,N_6638);
nand U9284 (N_9284,N_5421,N_6794);
and U9285 (N_9285,N_5472,N_5198);
nor U9286 (N_9286,N_6913,N_6804);
or U9287 (N_9287,N_7027,N_6893);
nor U9288 (N_9288,N_5611,N_5254);
and U9289 (N_9289,N_5209,N_5349);
nand U9290 (N_9290,N_5064,N_5648);
or U9291 (N_9291,N_5009,N_5639);
or U9292 (N_9292,N_5051,N_7494);
and U9293 (N_9293,N_7243,N_6732);
and U9294 (N_9294,N_6234,N_6982);
or U9295 (N_9295,N_5981,N_5101);
and U9296 (N_9296,N_7171,N_6151);
or U9297 (N_9297,N_6946,N_6196);
or U9298 (N_9298,N_6785,N_5704);
and U9299 (N_9299,N_5597,N_7011);
or U9300 (N_9300,N_6760,N_7172);
nor U9301 (N_9301,N_5966,N_5795);
and U9302 (N_9302,N_7381,N_6227);
nor U9303 (N_9303,N_5823,N_7312);
nand U9304 (N_9304,N_6508,N_6317);
nand U9305 (N_9305,N_6724,N_6565);
or U9306 (N_9306,N_5557,N_7236);
nand U9307 (N_9307,N_6269,N_6660);
nand U9308 (N_9308,N_6245,N_7148);
and U9309 (N_9309,N_5001,N_6384);
xor U9310 (N_9310,N_5595,N_5528);
nor U9311 (N_9311,N_6121,N_5363);
nand U9312 (N_9312,N_6718,N_7418);
and U9313 (N_9313,N_7270,N_6678);
nand U9314 (N_9314,N_5368,N_7252);
and U9315 (N_9315,N_5479,N_5652);
nor U9316 (N_9316,N_6099,N_6443);
nor U9317 (N_9317,N_5542,N_7436);
nand U9318 (N_9318,N_5428,N_6428);
nor U9319 (N_9319,N_5847,N_7044);
nor U9320 (N_9320,N_6321,N_5018);
nand U9321 (N_9321,N_5340,N_6602);
or U9322 (N_9322,N_7460,N_5568);
and U9323 (N_9323,N_5437,N_5058);
nand U9324 (N_9324,N_6478,N_6735);
nand U9325 (N_9325,N_6767,N_6229);
nor U9326 (N_9326,N_6628,N_7255);
nand U9327 (N_9327,N_6890,N_7308);
and U9328 (N_9328,N_6944,N_7368);
nor U9329 (N_9329,N_6122,N_5771);
and U9330 (N_9330,N_6818,N_6093);
nor U9331 (N_9331,N_6221,N_7090);
nor U9332 (N_9332,N_5043,N_5869);
and U9333 (N_9333,N_5311,N_5094);
and U9334 (N_9334,N_6579,N_6346);
or U9335 (N_9335,N_6568,N_6335);
nor U9336 (N_9336,N_6666,N_6236);
nand U9337 (N_9337,N_5628,N_5590);
and U9338 (N_9338,N_6542,N_6187);
or U9339 (N_9339,N_5217,N_5215);
and U9340 (N_9340,N_5843,N_7123);
nand U9341 (N_9341,N_6501,N_6127);
and U9342 (N_9342,N_7219,N_6610);
and U9343 (N_9343,N_6087,N_5987);
or U9344 (N_9344,N_5965,N_6043);
and U9345 (N_9345,N_6803,N_5824);
nor U9346 (N_9346,N_5528,N_5174);
xor U9347 (N_9347,N_6889,N_6832);
nand U9348 (N_9348,N_7429,N_7419);
or U9349 (N_9349,N_6879,N_5432);
nor U9350 (N_9350,N_5220,N_6316);
nor U9351 (N_9351,N_6676,N_5315);
and U9352 (N_9352,N_7303,N_7183);
and U9353 (N_9353,N_6403,N_7012);
nand U9354 (N_9354,N_5300,N_6050);
or U9355 (N_9355,N_7028,N_6956);
and U9356 (N_9356,N_6816,N_6838);
nand U9357 (N_9357,N_6132,N_5762);
xnor U9358 (N_9358,N_7246,N_7288);
or U9359 (N_9359,N_5913,N_5506);
nor U9360 (N_9360,N_6490,N_6417);
and U9361 (N_9361,N_6706,N_5912);
nand U9362 (N_9362,N_5759,N_6404);
nor U9363 (N_9363,N_5609,N_6010);
nor U9364 (N_9364,N_5610,N_5901);
and U9365 (N_9365,N_6707,N_7140);
or U9366 (N_9366,N_5466,N_7329);
and U9367 (N_9367,N_6413,N_5534);
or U9368 (N_9368,N_6313,N_6750);
and U9369 (N_9369,N_6634,N_7031);
and U9370 (N_9370,N_6740,N_7318);
and U9371 (N_9371,N_6628,N_5606);
or U9372 (N_9372,N_6623,N_5942);
and U9373 (N_9373,N_6486,N_5447);
nand U9374 (N_9374,N_6727,N_7179);
xor U9375 (N_9375,N_7238,N_6892);
nand U9376 (N_9376,N_5253,N_6066);
or U9377 (N_9377,N_6624,N_5087);
or U9378 (N_9378,N_5640,N_5954);
and U9379 (N_9379,N_7074,N_5897);
nor U9380 (N_9380,N_6899,N_6443);
nor U9381 (N_9381,N_6976,N_5461);
and U9382 (N_9382,N_6791,N_7395);
nand U9383 (N_9383,N_7188,N_7448);
nand U9384 (N_9384,N_6484,N_6127);
nand U9385 (N_9385,N_6843,N_5781);
and U9386 (N_9386,N_5401,N_5683);
and U9387 (N_9387,N_6707,N_5124);
nand U9388 (N_9388,N_5223,N_7099);
or U9389 (N_9389,N_5958,N_5967);
and U9390 (N_9390,N_7284,N_6342);
nor U9391 (N_9391,N_7267,N_5238);
nand U9392 (N_9392,N_5144,N_6523);
or U9393 (N_9393,N_6380,N_5927);
and U9394 (N_9394,N_6998,N_6358);
nor U9395 (N_9395,N_7042,N_5494);
and U9396 (N_9396,N_6075,N_5922);
and U9397 (N_9397,N_7183,N_5439);
nand U9398 (N_9398,N_7192,N_6411);
and U9399 (N_9399,N_5694,N_5308);
nor U9400 (N_9400,N_5160,N_5677);
or U9401 (N_9401,N_5888,N_7292);
nor U9402 (N_9402,N_5997,N_5735);
and U9403 (N_9403,N_5605,N_5121);
nor U9404 (N_9404,N_7102,N_6425);
or U9405 (N_9405,N_7414,N_6289);
and U9406 (N_9406,N_7098,N_5600);
nor U9407 (N_9407,N_6073,N_6453);
nand U9408 (N_9408,N_6295,N_7095);
nor U9409 (N_9409,N_5582,N_7346);
nor U9410 (N_9410,N_7401,N_5346);
nand U9411 (N_9411,N_7030,N_7014);
or U9412 (N_9412,N_7405,N_6891);
nor U9413 (N_9413,N_6643,N_5916);
or U9414 (N_9414,N_5596,N_6326);
nor U9415 (N_9415,N_5116,N_6815);
and U9416 (N_9416,N_6572,N_6968);
nor U9417 (N_9417,N_5121,N_6606);
nand U9418 (N_9418,N_6054,N_6405);
or U9419 (N_9419,N_6387,N_6907);
and U9420 (N_9420,N_7052,N_6831);
and U9421 (N_9421,N_6989,N_6811);
nor U9422 (N_9422,N_5745,N_5586);
nor U9423 (N_9423,N_5363,N_5564);
and U9424 (N_9424,N_6359,N_7216);
xnor U9425 (N_9425,N_6638,N_5188);
nand U9426 (N_9426,N_5549,N_6073);
nor U9427 (N_9427,N_5330,N_6436);
nor U9428 (N_9428,N_7358,N_6411);
nor U9429 (N_9429,N_6527,N_7238);
or U9430 (N_9430,N_7330,N_6829);
nor U9431 (N_9431,N_6286,N_5073);
nand U9432 (N_9432,N_5052,N_6857);
or U9433 (N_9433,N_6714,N_7060);
or U9434 (N_9434,N_5320,N_7340);
or U9435 (N_9435,N_6852,N_6161);
or U9436 (N_9436,N_5886,N_5288);
or U9437 (N_9437,N_5705,N_7203);
nand U9438 (N_9438,N_6631,N_6652);
and U9439 (N_9439,N_7259,N_5010);
nor U9440 (N_9440,N_5275,N_7112);
and U9441 (N_9441,N_5471,N_5077);
and U9442 (N_9442,N_5676,N_5463);
nand U9443 (N_9443,N_6880,N_7363);
or U9444 (N_9444,N_6503,N_5705);
and U9445 (N_9445,N_5603,N_7419);
or U9446 (N_9446,N_7268,N_5694);
nor U9447 (N_9447,N_6429,N_5295);
or U9448 (N_9448,N_7326,N_5583);
nor U9449 (N_9449,N_5219,N_5536);
nor U9450 (N_9450,N_5167,N_5125);
nand U9451 (N_9451,N_5098,N_6771);
or U9452 (N_9452,N_7312,N_6732);
or U9453 (N_9453,N_5385,N_6402);
nand U9454 (N_9454,N_5488,N_5520);
nor U9455 (N_9455,N_7244,N_5159);
nand U9456 (N_9456,N_5991,N_5285);
and U9457 (N_9457,N_6065,N_5573);
and U9458 (N_9458,N_5361,N_5063);
nor U9459 (N_9459,N_5640,N_5964);
nor U9460 (N_9460,N_5667,N_6113);
or U9461 (N_9461,N_5973,N_7135);
and U9462 (N_9462,N_6538,N_5214);
nor U9463 (N_9463,N_5736,N_6677);
or U9464 (N_9464,N_7097,N_6856);
nor U9465 (N_9465,N_6182,N_5843);
nor U9466 (N_9466,N_7019,N_6491);
and U9467 (N_9467,N_5173,N_5886);
nand U9468 (N_9468,N_6501,N_5073);
nand U9469 (N_9469,N_7306,N_6384);
and U9470 (N_9470,N_5677,N_6708);
nor U9471 (N_9471,N_6306,N_5723);
or U9472 (N_9472,N_5101,N_6624);
xnor U9473 (N_9473,N_6207,N_6164);
nand U9474 (N_9474,N_6883,N_5353);
nand U9475 (N_9475,N_7043,N_6065);
and U9476 (N_9476,N_6416,N_5687);
nor U9477 (N_9477,N_5131,N_6892);
and U9478 (N_9478,N_5854,N_6830);
or U9479 (N_9479,N_6461,N_6679);
nand U9480 (N_9480,N_6560,N_6813);
nand U9481 (N_9481,N_7470,N_7064);
or U9482 (N_9482,N_6106,N_7248);
and U9483 (N_9483,N_6639,N_6680);
nand U9484 (N_9484,N_6834,N_7242);
nand U9485 (N_9485,N_6808,N_6743);
nor U9486 (N_9486,N_5821,N_5770);
and U9487 (N_9487,N_6109,N_5040);
or U9488 (N_9488,N_5716,N_5356);
or U9489 (N_9489,N_5492,N_5854);
nor U9490 (N_9490,N_6972,N_5301);
nor U9491 (N_9491,N_6279,N_6583);
nand U9492 (N_9492,N_5766,N_5587);
or U9493 (N_9493,N_7147,N_6488);
and U9494 (N_9494,N_6532,N_5807);
or U9495 (N_9495,N_6434,N_6401);
nor U9496 (N_9496,N_5425,N_6974);
and U9497 (N_9497,N_7186,N_6178);
nand U9498 (N_9498,N_5063,N_7078);
and U9499 (N_9499,N_6898,N_7073);
or U9500 (N_9500,N_5791,N_5678);
nand U9501 (N_9501,N_6346,N_5669);
nand U9502 (N_9502,N_6177,N_6990);
and U9503 (N_9503,N_6740,N_6815);
and U9504 (N_9504,N_5630,N_5759);
nor U9505 (N_9505,N_6090,N_6270);
nand U9506 (N_9506,N_5087,N_6330);
or U9507 (N_9507,N_6290,N_5572);
or U9508 (N_9508,N_7176,N_7210);
and U9509 (N_9509,N_5613,N_6631);
or U9510 (N_9510,N_5963,N_5551);
or U9511 (N_9511,N_6985,N_5871);
nor U9512 (N_9512,N_5503,N_5497);
nand U9513 (N_9513,N_6029,N_7185);
and U9514 (N_9514,N_6602,N_6860);
nor U9515 (N_9515,N_6431,N_7451);
nor U9516 (N_9516,N_5195,N_6158);
or U9517 (N_9517,N_6474,N_5054);
nand U9518 (N_9518,N_6944,N_6475);
nor U9519 (N_9519,N_6080,N_6928);
or U9520 (N_9520,N_6442,N_6378);
nand U9521 (N_9521,N_5136,N_6656);
or U9522 (N_9522,N_5960,N_6705);
or U9523 (N_9523,N_6265,N_6653);
nand U9524 (N_9524,N_6135,N_7142);
nand U9525 (N_9525,N_5373,N_6463);
nor U9526 (N_9526,N_5956,N_6719);
nor U9527 (N_9527,N_6659,N_7378);
nor U9528 (N_9528,N_5517,N_5129);
nand U9529 (N_9529,N_5457,N_5193);
and U9530 (N_9530,N_7253,N_5338);
and U9531 (N_9531,N_5011,N_7085);
and U9532 (N_9532,N_6157,N_7343);
nor U9533 (N_9533,N_7446,N_5115);
and U9534 (N_9534,N_5077,N_6027);
and U9535 (N_9535,N_6959,N_5684);
and U9536 (N_9536,N_6462,N_7400);
or U9537 (N_9537,N_5380,N_6915);
or U9538 (N_9538,N_7226,N_5664);
nand U9539 (N_9539,N_6425,N_5549);
and U9540 (N_9540,N_6389,N_5676);
and U9541 (N_9541,N_5960,N_5797);
nor U9542 (N_9542,N_7195,N_6053);
nand U9543 (N_9543,N_6648,N_7133);
and U9544 (N_9544,N_6670,N_5134);
and U9545 (N_9545,N_6746,N_7465);
nand U9546 (N_9546,N_6227,N_7370);
and U9547 (N_9547,N_5674,N_6390);
or U9548 (N_9548,N_5191,N_6471);
and U9549 (N_9549,N_6041,N_6893);
nand U9550 (N_9550,N_6762,N_6494);
or U9551 (N_9551,N_5528,N_5004);
or U9552 (N_9552,N_6462,N_5945);
and U9553 (N_9553,N_7006,N_5010);
and U9554 (N_9554,N_7224,N_7094);
nor U9555 (N_9555,N_7295,N_7082);
nor U9556 (N_9556,N_6310,N_5023);
and U9557 (N_9557,N_7156,N_5504);
or U9558 (N_9558,N_6451,N_5049);
nand U9559 (N_9559,N_6458,N_5660);
nand U9560 (N_9560,N_6625,N_7375);
and U9561 (N_9561,N_6574,N_6643);
and U9562 (N_9562,N_5287,N_5024);
and U9563 (N_9563,N_6647,N_6611);
or U9564 (N_9564,N_7411,N_5282);
or U9565 (N_9565,N_7062,N_6252);
nand U9566 (N_9566,N_5824,N_7208);
nand U9567 (N_9567,N_6087,N_5676);
nor U9568 (N_9568,N_6311,N_5929);
nand U9569 (N_9569,N_5609,N_5483);
and U9570 (N_9570,N_6725,N_7349);
and U9571 (N_9571,N_7012,N_5762);
nand U9572 (N_9572,N_7344,N_5858);
and U9573 (N_9573,N_6512,N_6858);
or U9574 (N_9574,N_5899,N_6985);
and U9575 (N_9575,N_5194,N_6671);
nor U9576 (N_9576,N_5737,N_7425);
and U9577 (N_9577,N_6150,N_5644);
nand U9578 (N_9578,N_7037,N_6400);
and U9579 (N_9579,N_7000,N_6922);
and U9580 (N_9580,N_5339,N_5172);
or U9581 (N_9581,N_6970,N_6389);
nor U9582 (N_9582,N_7247,N_5501);
nand U9583 (N_9583,N_5353,N_7151);
or U9584 (N_9584,N_5508,N_5244);
and U9585 (N_9585,N_6286,N_6418);
xnor U9586 (N_9586,N_7301,N_6740);
and U9587 (N_9587,N_5648,N_6341);
and U9588 (N_9588,N_6284,N_5504);
nand U9589 (N_9589,N_5997,N_7446);
and U9590 (N_9590,N_5613,N_7352);
or U9591 (N_9591,N_7359,N_5049);
or U9592 (N_9592,N_6173,N_7351);
or U9593 (N_9593,N_6035,N_5561);
or U9594 (N_9594,N_6088,N_6315);
or U9595 (N_9595,N_6136,N_5247);
xor U9596 (N_9596,N_5401,N_6063);
nor U9597 (N_9597,N_5774,N_5064);
nor U9598 (N_9598,N_6797,N_5446);
and U9599 (N_9599,N_5626,N_6968);
nand U9600 (N_9600,N_6858,N_6319);
nor U9601 (N_9601,N_6685,N_6471);
nor U9602 (N_9602,N_5048,N_5182);
or U9603 (N_9603,N_7132,N_6817);
and U9604 (N_9604,N_6085,N_5671);
or U9605 (N_9605,N_6167,N_5143);
nor U9606 (N_9606,N_6464,N_6842);
or U9607 (N_9607,N_6833,N_6559);
nand U9608 (N_9608,N_6001,N_6984);
and U9609 (N_9609,N_7425,N_5939);
and U9610 (N_9610,N_6715,N_5870);
or U9611 (N_9611,N_6836,N_6017);
nand U9612 (N_9612,N_6274,N_6909);
and U9613 (N_9613,N_7191,N_7276);
nand U9614 (N_9614,N_6827,N_7414);
or U9615 (N_9615,N_6537,N_7414);
xor U9616 (N_9616,N_5975,N_6595);
or U9617 (N_9617,N_5060,N_6138);
nand U9618 (N_9618,N_5654,N_5157);
nor U9619 (N_9619,N_5758,N_5849);
and U9620 (N_9620,N_5429,N_5440);
and U9621 (N_9621,N_7461,N_7420);
nand U9622 (N_9622,N_5034,N_6284);
nand U9623 (N_9623,N_6192,N_7158);
and U9624 (N_9624,N_5728,N_5470);
nor U9625 (N_9625,N_5161,N_6031);
and U9626 (N_9626,N_5969,N_6474);
nand U9627 (N_9627,N_6273,N_6280);
or U9628 (N_9628,N_5293,N_6342);
nand U9629 (N_9629,N_5672,N_5682);
nand U9630 (N_9630,N_5047,N_6218);
nor U9631 (N_9631,N_6231,N_5691);
or U9632 (N_9632,N_7235,N_6795);
and U9633 (N_9633,N_6985,N_5851);
and U9634 (N_9634,N_6912,N_6129);
or U9635 (N_9635,N_6974,N_6207);
or U9636 (N_9636,N_5106,N_7238);
nand U9637 (N_9637,N_5285,N_6921);
and U9638 (N_9638,N_6542,N_5858);
nand U9639 (N_9639,N_5330,N_5531);
nor U9640 (N_9640,N_5842,N_5236);
nor U9641 (N_9641,N_6329,N_6286);
nand U9642 (N_9642,N_5921,N_6648);
or U9643 (N_9643,N_6065,N_6253);
nor U9644 (N_9644,N_5632,N_5401);
nor U9645 (N_9645,N_5711,N_5610);
nor U9646 (N_9646,N_5766,N_7164);
nor U9647 (N_9647,N_5153,N_6569);
nor U9648 (N_9648,N_5246,N_7038);
and U9649 (N_9649,N_6098,N_5929);
nand U9650 (N_9650,N_5673,N_5497);
and U9651 (N_9651,N_7164,N_6791);
nand U9652 (N_9652,N_5983,N_5265);
or U9653 (N_9653,N_6092,N_7428);
nand U9654 (N_9654,N_6971,N_5686);
nand U9655 (N_9655,N_7001,N_6606);
or U9656 (N_9656,N_6822,N_7095);
nor U9657 (N_9657,N_5573,N_6989);
nand U9658 (N_9658,N_5183,N_5146);
nor U9659 (N_9659,N_6873,N_7188);
and U9660 (N_9660,N_7376,N_5661);
and U9661 (N_9661,N_5732,N_6804);
and U9662 (N_9662,N_5459,N_7116);
or U9663 (N_9663,N_5455,N_6044);
nor U9664 (N_9664,N_5161,N_5885);
nor U9665 (N_9665,N_7301,N_6067);
and U9666 (N_9666,N_6823,N_6006);
or U9667 (N_9667,N_7307,N_6075);
and U9668 (N_9668,N_5693,N_6968);
nand U9669 (N_9669,N_6222,N_5656);
nand U9670 (N_9670,N_6763,N_7361);
and U9671 (N_9671,N_5743,N_6726);
nor U9672 (N_9672,N_7497,N_6981);
and U9673 (N_9673,N_5563,N_6800);
nand U9674 (N_9674,N_5950,N_5200);
and U9675 (N_9675,N_6269,N_6197);
nand U9676 (N_9676,N_5692,N_6574);
or U9677 (N_9677,N_5586,N_6286);
nand U9678 (N_9678,N_5467,N_6491);
or U9679 (N_9679,N_6517,N_6877);
and U9680 (N_9680,N_5744,N_6209);
and U9681 (N_9681,N_7089,N_7166);
and U9682 (N_9682,N_5224,N_5806);
nand U9683 (N_9683,N_6521,N_7480);
or U9684 (N_9684,N_5828,N_6428);
nand U9685 (N_9685,N_7256,N_6644);
nor U9686 (N_9686,N_5021,N_6891);
nor U9687 (N_9687,N_5420,N_7045);
nand U9688 (N_9688,N_6899,N_5006);
nor U9689 (N_9689,N_5865,N_5530);
nand U9690 (N_9690,N_6019,N_5291);
or U9691 (N_9691,N_7224,N_5413);
nor U9692 (N_9692,N_6813,N_5999);
or U9693 (N_9693,N_5836,N_6557);
and U9694 (N_9694,N_6108,N_6767);
nand U9695 (N_9695,N_5159,N_6937);
and U9696 (N_9696,N_6061,N_5105);
and U9697 (N_9697,N_5735,N_6435);
and U9698 (N_9698,N_6863,N_7244);
and U9699 (N_9699,N_6917,N_7166);
and U9700 (N_9700,N_7418,N_6246);
and U9701 (N_9701,N_7454,N_6858);
nor U9702 (N_9702,N_6558,N_5836);
and U9703 (N_9703,N_7120,N_5354);
nand U9704 (N_9704,N_6582,N_6730);
and U9705 (N_9705,N_5341,N_5745);
nor U9706 (N_9706,N_7246,N_5098);
or U9707 (N_9707,N_5732,N_5540);
or U9708 (N_9708,N_6060,N_6990);
nor U9709 (N_9709,N_5529,N_7305);
nand U9710 (N_9710,N_6834,N_5973);
nand U9711 (N_9711,N_5864,N_5646);
nor U9712 (N_9712,N_7037,N_7088);
nand U9713 (N_9713,N_5346,N_6658);
or U9714 (N_9714,N_6300,N_5571);
and U9715 (N_9715,N_7484,N_7123);
and U9716 (N_9716,N_6064,N_5161);
nor U9717 (N_9717,N_6256,N_6218);
and U9718 (N_9718,N_5427,N_7348);
nor U9719 (N_9719,N_5890,N_6168);
or U9720 (N_9720,N_5774,N_6079);
nand U9721 (N_9721,N_5906,N_5723);
or U9722 (N_9722,N_6003,N_5448);
or U9723 (N_9723,N_6542,N_7279);
and U9724 (N_9724,N_6727,N_6001);
nor U9725 (N_9725,N_7170,N_6109);
or U9726 (N_9726,N_5982,N_6275);
or U9727 (N_9727,N_5625,N_7184);
nor U9728 (N_9728,N_5778,N_7201);
or U9729 (N_9729,N_6247,N_6091);
nor U9730 (N_9730,N_6419,N_7290);
and U9731 (N_9731,N_5805,N_5888);
nand U9732 (N_9732,N_7007,N_5949);
nor U9733 (N_9733,N_6076,N_5702);
and U9734 (N_9734,N_6748,N_7073);
and U9735 (N_9735,N_6145,N_5522);
nand U9736 (N_9736,N_6768,N_6308);
nor U9737 (N_9737,N_6964,N_5199);
or U9738 (N_9738,N_5350,N_6232);
or U9739 (N_9739,N_6278,N_6916);
nand U9740 (N_9740,N_7426,N_6477);
and U9741 (N_9741,N_7173,N_6547);
nand U9742 (N_9742,N_6627,N_7078);
nor U9743 (N_9743,N_5515,N_6102);
nand U9744 (N_9744,N_6179,N_5572);
nor U9745 (N_9745,N_5109,N_7455);
or U9746 (N_9746,N_6106,N_5586);
nor U9747 (N_9747,N_5143,N_7095);
xnor U9748 (N_9748,N_5538,N_6738);
nand U9749 (N_9749,N_7216,N_5078);
and U9750 (N_9750,N_5747,N_6150);
or U9751 (N_9751,N_6181,N_5022);
nand U9752 (N_9752,N_5098,N_7396);
or U9753 (N_9753,N_6016,N_5727);
nand U9754 (N_9754,N_5375,N_5089);
xnor U9755 (N_9755,N_5508,N_7091);
nand U9756 (N_9756,N_5632,N_5088);
and U9757 (N_9757,N_6140,N_5077);
nand U9758 (N_9758,N_5070,N_5580);
nand U9759 (N_9759,N_7115,N_6370);
nor U9760 (N_9760,N_5703,N_6254);
or U9761 (N_9761,N_5741,N_7176);
nand U9762 (N_9762,N_5352,N_7311);
and U9763 (N_9763,N_6717,N_6391);
and U9764 (N_9764,N_6742,N_5846);
and U9765 (N_9765,N_5926,N_6447);
nand U9766 (N_9766,N_7034,N_6341);
or U9767 (N_9767,N_6264,N_6238);
nand U9768 (N_9768,N_6591,N_5494);
nor U9769 (N_9769,N_7398,N_5157);
nor U9770 (N_9770,N_5729,N_5153);
nand U9771 (N_9771,N_6130,N_6650);
or U9772 (N_9772,N_7456,N_6021);
or U9773 (N_9773,N_6890,N_5114);
nor U9774 (N_9774,N_5938,N_5272);
nand U9775 (N_9775,N_5973,N_6792);
nand U9776 (N_9776,N_5661,N_5788);
and U9777 (N_9777,N_6008,N_6312);
nand U9778 (N_9778,N_6274,N_7375);
and U9779 (N_9779,N_7113,N_7331);
nand U9780 (N_9780,N_6876,N_5606);
nor U9781 (N_9781,N_5671,N_7393);
and U9782 (N_9782,N_7019,N_7140);
and U9783 (N_9783,N_6635,N_7489);
or U9784 (N_9784,N_7305,N_5002);
and U9785 (N_9785,N_5732,N_7114);
nand U9786 (N_9786,N_6696,N_5166);
and U9787 (N_9787,N_6116,N_6551);
nand U9788 (N_9788,N_6012,N_5505);
and U9789 (N_9789,N_6389,N_5883);
or U9790 (N_9790,N_5149,N_7114);
or U9791 (N_9791,N_5357,N_6469);
or U9792 (N_9792,N_6649,N_7111);
nor U9793 (N_9793,N_5474,N_6314);
nor U9794 (N_9794,N_7381,N_6857);
or U9795 (N_9795,N_5064,N_7250);
nor U9796 (N_9796,N_6476,N_6284);
nor U9797 (N_9797,N_7454,N_5728);
or U9798 (N_9798,N_5949,N_5688);
or U9799 (N_9799,N_6794,N_5927);
nand U9800 (N_9800,N_5318,N_5122);
or U9801 (N_9801,N_6736,N_7077);
and U9802 (N_9802,N_6753,N_5281);
or U9803 (N_9803,N_5273,N_6831);
nand U9804 (N_9804,N_5467,N_5904);
nor U9805 (N_9805,N_5048,N_6220);
or U9806 (N_9806,N_6098,N_6755);
or U9807 (N_9807,N_5652,N_5571);
nand U9808 (N_9808,N_5113,N_5903);
and U9809 (N_9809,N_6150,N_5977);
nand U9810 (N_9810,N_5996,N_6007);
or U9811 (N_9811,N_6506,N_5614);
or U9812 (N_9812,N_7229,N_6361);
nor U9813 (N_9813,N_6438,N_6632);
nand U9814 (N_9814,N_5306,N_5659);
and U9815 (N_9815,N_5092,N_5293);
nor U9816 (N_9816,N_6434,N_6735);
or U9817 (N_9817,N_7132,N_5287);
or U9818 (N_9818,N_5498,N_5123);
nand U9819 (N_9819,N_5462,N_6407);
nand U9820 (N_9820,N_6136,N_7111);
nand U9821 (N_9821,N_5775,N_6644);
or U9822 (N_9822,N_6482,N_5664);
nor U9823 (N_9823,N_5150,N_7385);
nand U9824 (N_9824,N_5516,N_7037);
or U9825 (N_9825,N_5699,N_6194);
nor U9826 (N_9826,N_6820,N_7050);
and U9827 (N_9827,N_6947,N_7305);
nor U9828 (N_9828,N_6944,N_6209);
nor U9829 (N_9829,N_5899,N_6062);
and U9830 (N_9830,N_7088,N_7239);
nor U9831 (N_9831,N_5848,N_5967);
nand U9832 (N_9832,N_6407,N_6916);
nand U9833 (N_9833,N_6860,N_5599);
nand U9834 (N_9834,N_6501,N_5364);
nor U9835 (N_9835,N_5178,N_6321);
nand U9836 (N_9836,N_5611,N_5071);
nand U9837 (N_9837,N_6413,N_7111);
or U9838 (N_9838,N_5633,N_7199);
or U9839 (N_9839,N_6870,N_5890);
or U9840 (N_9840,N_6214,N_5331);
or U9841 (N_9841,N_5640,N_5510);
nand U9842 (N_9842,N_5813,N_5593);
nand U9843 (N_9843,N_6268,N_5894);
nor U9844 (N_9844,N_6642,N_6362);
xor U9845 (N_9845,N_6312,N_6103);
or U9846 (N_9846,N_5097,N_5152);
and U9847 (N_9847,N_5080,N_5888);
or U9848 (N_9848,N_5439,N_7224);
or U9849 (N_9849,N_5530,N_5323);
nor U9850 (N_9850,N_6414,N_6227);
nand U9851 (N_9851,N_6673,N_5950);
nor U9852 (N_9852,N_7396,N_7495);
nand U9853 (N_9853,N_6346,N_6132);
and U9854 (N_9854,N_5240,N_6315);
nand U9855 (N_9855,N_6476,N_5238);
or U9856 (N_9856,N_6999,N_5828);
or U9857 (N_9857,N_7221,N_6544);
nor U9858 (N_9858,N_6949,N_5666);
or U9859 (N_9859,N_5807,N_5737);
or U9860 (N_9860,N_5660,N_6623);
nand U9861 (N_9861,N_7351,N_5263);
nand U9862 (N_9862,N_5925,N_5350);
or U9863 (N_9863,N_5687,N_5814);
nor U9864 (N_9864,N_6050,N_6532);
nor U9865 (N_9865,N_5829,N_6948);
nor U9866 (N_9866,N_5144,N_6862);
and U9867 (N_9867,N_6142,N_6392);
or U9868 (N_9868,N_7180,N_6903);
nor U9869 (N_9869,N_6891,N_6161);
nor U9870 (N_9870,N_7209,N_5704);
and U9871 (N_9871,N_7351,N_7209);
nand U9872 (N_9872,N_6480,N_6373);
nor U9873 (N_9873,N_6398,N_5741);
nand U9874 (N_9874,N_5664,N_6961);
or U9875 (N_9875,N_5268,N_5482);
or U9876 (N_9876,N_7369,N_6559);
nor U9877 (N_9877,N_7479,N_7236);
nand U9878 (N_9878,N_7451,N_6086);
and U9879 (N_9879,N_5729,N_6816);
nand U9880 (N_9880,N_6716,N_6664);
or U9881 (N_9881,N_6914,N_6745);
or U9882 (N_9882,N_6549,N_5124);
nand U9883 (N_9883,N_5801,N_7008);
and U9884 (N_9884,N_6451,N_6109);
and U9885 (N_9885,N_6268,N_5765);
or U9886 (N_9886,N_5728,N_5567);
nand U9887 (N_9887,N_6702,N_6863);
or U9888 (N_9888,N_6182,N_7416);
and U9889 (N_9889,N_5368,N_7281);
nor U9890 (N_9890,N_6626,N_7005);
nand U9891 (N_9891,N_5748,N_6595);
or U9892 (N_9892,N_5361,N_5943);
xor U9893 (N_9893,N_5409,N_6833);
or U9894 (N_9894,N_6732,N_6202);
nor U9895 (N_9895,N_5605,N_7117);
nor U9896 (N_9896,N_6976,N_5799);
nor U9897 (N_9897,N_6015,N_6288);
and U9898 (N_9898,N_6059,N_5515);
nor U9899 (N_9899,N_6819,N_5180);
nor U9900 (N_9900,N_5805,N_7052);
nand U9901 (N_9901,N_6904,N_7122);
and U9902 (N_9902,N_6025,N_5826);
nand U9903 (N_9903,N_5474,N_6741);
nand U9904 (N_9904,N_5287,N_6971);
or U9905 (N_9905,N_6998,N_6144);
or U9906 (N_9906,N_6744,N_6086);
nor U9907 (N_9907,N_7342,N_5377);
nor U9908 (N_9908,N_6298,N_5970);
or U9909 (N_9909,N_5900,N_5599);
xnor U9910 (N_9910,N_5543,N_6637);
nand U9911 (N_9911,N_7443,N_5240);
or U9912 (N_9912,N_6715,N_5130);
and U9913 (N_9913,N_7050,N_6923);
or U9914 (N_9914,N_7438,N_6477);
nor U9915 (N_9915,N_5800,N_6390);
nor U9916 (N_9916,N_5720,N_6415);
nor U9917 (N_9917,N_6659,N_5131);
nor U9918 (N_9918,N_5717,N_6982);
and U9919 (N_9919,N_6158,N_5095);
nand U9920 (N_9920,N_6469,N_6018);
nor U9921 (N_9921,N_6517,N_5184);
and U9922 (N_9922,N_6263,N_6870);
or U9923 (N_9923,N_6113,N_7191);
nand U9924 (N_9924,N_5176,N_7192);
nand U9925 (N_9925,N_5147,N_6284);
xnor U9926 (N_9926,N_7234,N_7006);
nor U9927 (N_9927,N_6630,N_6662);
or U9928 (N_9928,N_6902,N_5921);
nor U9929 (N_9929,N_5917,N_6755);
nand U9930 (N_9930,N_6759,N_6937);
nand U9931 (N_9931,N_6154,N_5242);
nand U9932 (N_9932,N_6944,N_6381);
and U9933 (N_9933,N_6877,N_5636);
nand U9934 (N_9934,N_5212,N_7105);
and U9935 (N_9935,N_6207,N_7343);
nand U9936 (N_9936,N_6868,N_7154);
nor U9937 (N_9937,N_6952,N_6861);
nand U9938 (N_9938,N_5272,N_7092);
and U9939 (N_9939,N_7338,N_7445);
and U9940 (N_9940,N_5506,N_6081);
or U9941 (N_9941,N_5058,N_7489);
or U9942 (N_9942,N_7089,N_5886);
nor U9943 (N_9943,N_7107,N_6903);
or U9944 (N_9944,N_5617,N_6095);
nand U9945 (N_9945,N_5405,N_7169);
or U9946 (N_9946,N_5542,N_7290);
nor U9947 (N_9947,N_6012,N_6113);
nor U9948 (N_9948,N_7482,N_5074);
nor U9949 (N_9949,N_6594,N_6687);
or U9950 (N_9950,N_5132,N_6982);
nand U9951 (N_9951,N_5122,N_5591);
nor U9952 (N_9952,N_5337,N_6215);
or U9953 (N_9953,N_6786,N_6018);
and U9954 (N_9954,N_6444,N_6059);
nand U9955 (N_9955,N_7232,N_7010);
or U9956 (N_9956,N_5872,N_7160);
nand U9957 (N_9957,N_5013,N_7073);
nand U9958 (N_9958,N_5359,N_5446);
or U9959 (N_9959,N_6843,N_7397);
or U9960 (N_9960,N_6307,N_5994);
and U9961 (N_9961,N_6541,N_5971);
and U9962 (N_9962,N_5593,N_5681);
and U9963 (N_9963,N_6103,N_5678);
nand U9964 (N_9964,N_7064,N_5713);
and U9965 (N_9965,N_6378,N_5163);
or U9966 (N_9966,N_5926,N_5645);
and U9967 (N_9967,N_5687,N_7245);
nand U9968 (N_9968,N_7364,N_6113);
or U9969 (N_9969,N_5970,N_6398);
nor U9970 (N_9970,N_6131,N_7108);
nor U9971 (N_9971,N_6948,N_5900);
or U9972 (N_9972,N_7099,N_7309);
xnor U9973 (N_9973,N_7033,N_6662);
nand U9974 (N_9974,N_6476,N_6023);
nand U9975 (N_9975,N_5660,N_7428);
or U9976 (N_9976,N_6994,N_5590);
nand U9977 (N_9977,N_6217,N_7238);
nand U9978 (N_9978,N_5785,N_7258);
and U9979 (N_9979,N_6703,N_7344);
or U9980 (N_9980,N_5378,N_5954);
or U9981 (N_9981,N_5574,N_5953);
nand U9982 (N_9982,N_7201,N_6844);
or U9983 (N_9983,N_7426,N_5457);
nand U9984 (N_9984,N_6156,N_5452);
or U9985 (N_9985,N_6016,N_5297);
nor U9986 (N_9986,N_6467,N_5645);
nor U9987 (N_9987,N_5011,N_6343);
nand U9988 (N_9988,N_6115,N_5901);
or U9989 (N_9989,N_6785,N_5406);
nor U9990 (N_9990,N_5790,N_5265);
and U9991 (N_9991,N_5066,N_6759);
nor U9992 (N_9992,N_7120,N_7276);
or U9993 (N_9993,N_5888,N_6764);
nand U9994 (N_9994,N_6697,N_6767);
nand U9995 (N_9995,N_6448,N_5887);
or U9996 (N_9996,N_5577,N_6948);
and U9997 (N_9997,N_5710,N_5702);
nor U9998 (N_9998,N_7120,N_6323);
and U9999 (N_9999,N_7256,N_5142);
nand UO_0 (O_0,N_8839,N_8582);
nor UO_1 (O_1,N_8745,N_8938);
nand UO_2 (O_2,N_8836,N_8030);
nand UO_3 (O_3,N_8845,N_9609);
and UO_4 (O_4,N_8342,N_9413);
nor UO_5 (O_5,N_9541,N_9838);
or UO_6 (O_6,N_7581,N_9367);
or UO_7 (O_7,N_9555,N_9973);
and UO_8 (O_8,N_9300,N_7868);
or UO_9 (O_9,N_9060,N_8795);
nand UO_10 (O_10,N_9497,N_9680);
and UO_11 (O_11,N_8132,N_8639);
and UO_12 (O_12,N_8599,N_9959);
or UO_13 (O_13,N_7927,N_7904);
nand UO_14 (O_14,N_8310,N_8256);
nor UO_15 (O_15,N_8637,N_8065);
nor UO_16 (O_16,N_9032,N_8859);
nand UO_17 (O_17,N_7801,N_7632);
nor UO_18 (O_18,N_8482,N_8224);
nor UO_19 (O_19,N_8192,N_9692);
nor UO_20 (O_20,N_9711,N_7620);
nand UO_21 (O_21,N_8759,N_9518);
and UO_22 (O_22,N_8411,N_9850);
nand UO_23 (O_23,N_9050,N_9107);
nor UO_24 (O_24,N_8855,N_9172);
nand UO_25 (O_25,N_9411,N_8661);
nand UO_26 (O_26,N_8327,N_9767);
or UO_27 (O_27,N_8353,N_9179);
nor UO_28 (O_28,N_9800,N_8138);
or UO_29 (O_29,N_9905,N_9092);
or UO_30 (O_30,N_8079,N_7876);
nand UO_31 (O_31,N_9448,N_9823);
nand UO_32 (O_32,N_9424,N_9807);
or UO_33 (O_33,N_8468,N_7624);
nand UO_34 (O_34,N_9126,N_9952);
nor UO_35 (O_35,N_7901,N_8526);
nor UO_36 (O_36,N_9094,N_8470);
and UO_37 (O_37,N_8767,N_9849);
or UO_38 (O_38,N_7948,N_8788);
nor UO_39 (O_39,N_7995,N_8766);
and UO_40 (O_40,N_8010,N_8055);
nand UO_41 (O_41,N_9827,N_9420);
and UO_42 (O_42,N_8469,N_8674);
and UO_43 (O_43,N_8155,N_7764);
and UO_44 (O_44,N_9073,N_8241);
or UO_45 (O_45,N_8508,N_8518);
or UO_46 (O_46,N_8198,N_9370);
and UO_47 (O_47,N_8507,N_8997);
nor UO_48 (O_48,N_8877,N_8301);
nand UO_49 (O_49,N_9922,N_9347);
or UO_50 (O_50,N_9855,N_8764);
nand UO_51 (O_51,N_9858,N_8294);
nor UO_52 (O_52,N_9842,N_8513);
or UO_53 (O_53,N_8169,N_8045);
nor UO_54 (O_54,N_8874,N_8221);
and UO_55 (O_55,N_9998,N_9070);
or UO_56 (O_56,N_7880,N_7798);
or UO_57 (O_57,N_9241,N_9319);
and UO_58 (O_58,N_8897,N_9771);
or UO_59 (O_59,N_7780,N_9691);
and UO_60 (O_60,N_7735,N_7902);
nor UO_61 (O_61,N_8087,N_9787);
nand UO_62 (O_62,N_7794,N_8512);
nor UO_63 (O_63,N_9699,N_8796);
nand UO_64 (O_64,N_8243,N_9949);
and UO_65 (O_65,N_7922,N_9100);
nor UO_66 (O_66,N_8977,N_8509);
and UO_67 (O_67,N_7743,N_7938);
and UO_68 (O_68,N_9893,N_9540);
nand UO_69 (O_69,N_8696,N_8946);
nand UO_70 (O_70,N_8188,N_7918);
nand UO_71 (O_71,N_8817,N_8704);
nor UO_72 (O_72,N_7592,N_7903);
nand UO_73 (O_73,N_8016,N_8925);
and UO_74 (O_74,N_7627,N_8762);
nor UO_75 (O_75,N_8731,N_8664);
and UO_76 (O_76,N_7828,N_9221);
nand UO_77 (O_77,N_9613,N_7593);
and UO_78 (O_78,N_8950,N_9324);
nand UO_79 (O_79,N_8370,N_8211);
or UO_80 (O_80,N_7680,N_8751);
nand UO_81 (O_81,N_8690,N_8868);
nand UO_82 (O_82,N_9753,N_9415);
or UO_83 (O_83,N_9023,N_7830);
and UO_84 (O_84,N_8364,N_8746);
nand UO_85 (O_85,N_7838,N_9496);
and UO_86 (O_86,N_8414,N_9174);
nor UO_87 (O_87,N_8734,N_8500);
nand UO_88 (O_88,N_8214,N_9789);
nand UO_89 (O_89,N_8075,N_8604);
and UO_90 (O_90,N_8572,N_7991);
nor UO_91 (O_91,N_8929,N_8015);
and UO_92 (O_92,N_7808,N_8275);
nand UO_93 (O_93,N_7961,N_8164);
and UO_94 (O_94,N_8653,N_9610);
and UO_95 (O_95,N_7879,N_9469);
nand UO_96 (O_96,N_7944,N_9351);
nand UO_97 (O_97,N_8412,N_8565);
and UO_98 (O_98,N_7651,N_9472);
nand UO_99 (O_99,N_7863,N_8799);
or UO_100 (O_100,N_9397,N_8625);
and UO_101 (O_101,N_7689,N_9586);
nor UO_102 (O_102,N_9095,N_9218);
and UO_103 (O_103,N_7869,N_8154);
nand UO_104 (O_104,N_9658,N_8820);
nand UO_105 (O_105,N_8095,N_8144);
and UO_106 (O_106,N_8430,N_7841);
nor UO_107 (O_107,N_7625,N_8854);
and UO_108 (O_108,N_7534,N_7742);
and UO_109 (O_109,N_8419,N_8876);
nor UO_110 (O_110,N_9794,N_8388);
nand UO_111 (O_111,N_9272,N_9607);
nand UO_112 (O_112,N_9734,N_9573);
or UO_113 (O_113,N_9403,N_8418);
nand UO_114 (O_114,N_9080,N_8880);
nor UO_115 (O_115,N_8392,N_8161);
or UO_116 (O_116,N_8094,N_7820);
nand UO_117 (O_117,N_9890,N_9649);
or UO_118 (O_118,N_9662,N_8752);
or UO_119 (O_119,N_8398,N_7628);
nand UO_120 (O_120,N_9685,N_8521);
nand UO_121 (O_121,N_9962,N_9234);
and UO_122 (O_122,N_8922,N_8023);
nand UO_123 (O_123,N_8076,N_8628);
or UO_124 (O_124,N_8748,N_9048);
nand UO_125 (O_125,N_7762,N_9034);
nor UO_126 (O_126,N_9236,N_7595);
nor UO_127 (O_127,N_7616,N_8505);
nand UO_128 (O_128,N_7555,N_7776);
and UO_129 (O_129,N_9731,N_9512);
nor UO_130 (O_130,N_9097,N_7635);
nand UO_131 (O_131,N_9908,N_7512);
and UO_132 (O_132,N_8683,N_9372);
nor UO_133 (O_133,N_9406,N_9686);
nor UO_134 (O_134,N_8973,N_8601);
and UO_135 (O_135,N_8197,N_7516);
nor UO_136 (O_136,N_9741,N_9620);
nor UO_137 (O_137,N_9345,N_9943);
or UO_138 (O_138,N_9309,N_8099);
and UO_139 (O_139,N_9334,N_9166);
nand UO_140 (O_140,N_7818,N_9918);
and UO_141 (O_141,N_9726,N_7973);
nor UO_142 (O_142,N_9804,N_7727);
nand UO_143 (O_143,N_9005,N_9932);
nand UO_144 (O_144,N_9368,N_9493);
or UO_145 (O_145,N_7972,N_8082);
nor UO_146 (O_146,N_9453,N_9839);
nand UO_147 (O_147,N_9862,N_7898);
and UO_148 (O_148,N_9043,N_9957);
nand UO_149 (O_149,N_9875,N_7993);
nand UO_150 (O_150,N_9615,N_9207);
nand UO_151 (O_151,N_8088,N_9733);
nand UO_152 (O_152,N_8904,N_7572);
nand UO_153 (O_153,N_8806,N_9052);
nor UO_154 (O_154,N_7761,N_9260);
and UO_155 (O_155,N_9841,N_9900);
nand UO_156 (O_156,N_7747,N_9116);
nand UO_157 (O_157,N_7521,N_9441);
nor UO_158 (O_158,N_7967,N_9478);
or UO_159 (O_159,N_9251,N_8575);
or UO_160 (O_160,N_9944,N_8047);
or UO_161 (O_161,N_9579,N_9990);
nor UO_162 (O_162,N_8570,N_9145);
nor UO_163 (O_163,N_8589,N_8586);
nand UO_164 (O_164,N_7782,N_8288);
nor UO_165 (O_165,N_7577,N_9676);
or UO_166 (O_166,N_9399,N_9056);
nor UO_167 (O_167,N_9750,N_8264);
nand UO_168 (O_168,N_7951,N_8375);
or UO_169 (O_169,N_7923,N_9114);
or UO_170 (O_170,N_7525,N_7655);
nor UO_171 (O_171,N_9795,N_7607);
or UO_172 (O_172,N_9027,N_7936);
nor UO_173 (O_173,N_7988,N_9119);
or UO_174 (O_174,N_8728,N_9860);
nor UO_175 (O_175,N_7849,N_9854);
nand UO_176 (O_176,N_9373,N_7781);
nand UO_177 (O_177,N_9972,N_7544);
nand UO_178 (O_178,N_7935,N_8598);
xnor UO_179 (O_179,N_9778,N_9171);
or UO_180 (O_180,N_9481,N_9267);
or UO_181 (O_181,N_7891,N_8506);
nor UO_182 (O_182,N_7603,N_8822);
nand UO_183 (O_183,N_8835,N_9679);
and UO_184 (O_184,N_7515,N_7677);
and UO_185 (O_185,N_7738,N_8052);
nor UO_186 (O_186,N_8557,N_8810);
or UO_187 (O_187,N_8544,N_7746);
and UO_188 (O_188,N_8891,N_9987);
or UO_189 (O_189,N_9813,N_9316);
or UO_190 (O_190,N_9906,N_8449);
and UO_191 (O_191,N_8270,N_8133);
nand UO_192 (O_192,N_9970,N_9008);
nor UO_193 (O_193,N_9786,N_9099);
nor UO_194 (O_194,N_9700,N_9640);
or UO_195 (O_195,N_8818,N_8816);
nand UO_196 (O_196,N_9417,N_7752);
nand UO_197 (O_197,N_9035,N_8062);
or UO_198 (O_198,N_7709,N_9825);
and UO_199 (O_199,N_9999,N_8051);
nor UO_200 (O_200,N_8407,N_7569);
nor UO_201 (O_201,N_8149,N_7562);
and UO_202 (O_202,N_9889,N_7598);
or UO_203 (O_203,N_9561,N_7688);
and UO_204 (O_204,N_8669,N_9728);
or UO_205 (O_205,N_8383,N_7609);
or UO_206 (O_206,N_9069,N_9661);
and UO_207 (O_207,N_7817,N_8479);
nand UO_208 (O_208,N_8417,N_9047);
nor UO_209 (O_209,N_8665,N_7653);
nand UO_210 (O_210,N_9516,N_8536);
or UO_211 (O_211,N_7864,N_9200);
and UO_212 (O_212,N_7896,N_8714);
nor UO_213 (O_213,N_8970,N_9104);
nor UO_214 (O_214,N_7714,N_8381);
or UO_215 (O_215,N_8178,N_9020);
nor UO_216 (O_216,N_8534,N_9393);
nand UO_217 (O_217,N_9337,N_8223);
or UO_218 (O_218,N_9756,N_9562);
nor UO_219 (O_219,N_8120,N_8231);
and UO_220 (O_220,N_7588,N_9625);
nand UO_221 (O_221,N_8140,N_9395);
or UO_222 (O_222,N_7882,N_8940);
nand UO_223 (O_223,N_8056,N_8332);
or UO_224 (O_224,N_9296,N_9899);
nand UO_225 (O_225,N_9852,N_9582);
and UO_226 (O_226,N_9101,N_8083);
nor UO_227 (O_227,N_8860,N_9301);
nor UO_228 (O_228,N_8899,N_9567);
and UO_229 (O_229,N_9435,N_9216);
nand UO_230 (O_230,N_9278,N_9210);
nand UO_231 (O_231,N_7905,N_8190);
and UO_232 (O_232,N_9773,N_8048);
or UO_233 (O_233,N_7510,N_7899);
and UO_234 (O_234,N_9519,N_9531);
nand UO_235 (O_235,N_9202,N_7968);
and UO_236 (O_236,N_8488,N_8237);
or UO_237 (O_237,N_9530,N_7622);
nand UO_238 (O_238,N_9643,N_9239);
and UO_239 (O_239,N_9678,N_8576);
nand UO_240 (O_240,N_9856,N_9590);
nor UO_241 (O_241,N_8283,N_7731);
nand UO_242 (O_242,N_9327,N_8801);
nand UO_243 (O_243,N_7543,N_8614);
or UO_244 (O_244,N_8424,N_8898);
and UO_245 (O_245,N_8335,N_8196);
or UO_246 (O_246,N_9230,N_7802);
or UO_247 (O_247,N_9792,N_8141);
nand UO_248 (O_248,N_8720,N_8152);
and UO_249 (O_249,N_8621,N_9380);
nor UO_250 (O_250,N_8260,N_9112);
nand UO_251 (O_251,N_9712,N_8394);
and UO_252 (O_252,N_8176,N_7590);
and UO_253 (O_253,N_8890,N_9134);
or UO_254 (O_254,N_9359,N_8632);
or UO_255 (O_255,N_9132,N_9802);
nand UO_256 (O_256,N_9705,N_9559);
and UO_257 (O_257,N_8921,N_9198);
nand UO_258 (O_258,N_9798,N_8969);
and UO_259 (O_259,N_7816,N_7987);
nor UO_260 (O_260,N_7770,N_9709);
nand UO_261 (O_261,N_8692,N_9664);
xnor UO_262 (O_262,N_9204,N_8109);
and UO_263 (O_263,N_9211,N_8773);
nand UO_264 (O_264,N_8914,N_9294);
or UO_265 (O_265,N_8432,N_9365);
or UO_266 (O_266,N_7528,N_7943);
nand UO_267 (O_267,N_7806,N_7872);
nand UO_268 (O_268,N_8368,N_7832);
and UO_269 (O_269,N_8213,N_7698);
nor UO_270 (O_270,N_9464,N_9102);
or UO_271 (O_271,N_9332,N_9755);
or UO_272 (O_272,N_8131,N_7647);
and UO_273 (O_273,N_7504,N_8778);
nand UO_274 (O_274,N_8957,N_8805);
or UO_275 (O_275,N_8996,N_7757);
nand UO_276 (O_276,N_8910,N_7812);
and UO_277 (O_277,N_9475,N_8815);
or UO_278 (O_278,N_9015,N_8971);
or UO_279 (O_279,N_8261,N_8620);
and UO_280 (O_280,N_9488,N_9244);
and UO_281 (O_281,N_9517,N_9085);
or UO_282 (O_282,N_9446,N_7545);
and UO_283 (O_283,N_9730,N_8587);
nand UO_284 (O_284,N_9660,N_8091);
or UO_285 (O_285,N_7795,N_8017);
and UO_286 (O_286,N_7921,N_9279);
or UO_287 (O_287,N_8093,N_8299);
nor UO_288 (O_288,N_8504,N_7969);
nand UO_289 (O_289,N_9322,N_9898);
nor UO_290 (O_290,N_8841,N_8548);
and UO_291 (O_291,N_9532,N_8069);
or UO_292 (O_292,N_7733,N_9877);
and UO_293 (O_293,N_7845,N_9407);
or UO_294 (O_294,N_8790,N_9500);
nand UO_295 (O_295,N_9729,N_7977);
and UO_296 (O_296,N_7884,N_9865);
nor UO_297 (O_297,N_8619,N_9414);
nand UO_298 (O_298,N_8349,N_8077);
and UO_299 (O_299,N_7700,N_8749);
nor UO_300 (O_300,N_8351,N_8225);
nand UO_301 (O_301,N_9556,N_8769);
and UO_302 (O_302,N_9298,N_7835);
nor UO_303 (O_303,N_7566,N_9748);
or UO_304 (O_304,N_7759,N_9977);
or UO_305 (O_305,N_9285,N_9317);
nand UO_306 (O_306,N_7576,N_8054);
and UO_307 (O_307,N_9096,N_7906);
nor UO_308 (O_308,N_7621,N_9287);
nor UO_309 (O_309,N_9809,N_9781);
or UO_310 (O_310,N_9539,N_9017);
nor UO_311 (O_311,N_8926,N_8286);
and UO_312 (O_312,N_7914,N_7631);
nand UO_313 (O_313,N_7767,N_8654);
or UO_314 (O_314,N_9156,N_9992);
nand UO_315 (O_315,N_8687,N_7537);
nand UO_316 (O_316,N_8732,N_9024);
or UO_317 (O_317,N_7791,N_8360);
nand UO_318 (O_318,N_9895,N_9391);
or UO_319 (O_319,N_8166,N_7763);
or UO_320 (O_320,N_8736,N_9923);
and UO_321 (O_321,N_9945,N_9969);
and UO_322 (O_322,N_7813,N_9003);
and UO_323 (O_323,N_9161,N_9378);
nor UO_324 (O_324,N_8964,N_9338);
and UO_325 (O_325,N_8501,N_9468);
nand UO_326 (O_326,N_9265,N_8340);
nor UO_327 (O_327,N_9398,N_7568);
and UO_328 (O_328,N_7716,N_8523);
nand UO_329 (O_329,N_9713,N_7619);
nand UO_330 (O_330,N_7549,N_8535);
or UO_331 (O_331,N_9892,N_8333);
and UO_332 (O_332,N_9656,N_9921);
nor UO_333 (O_333,N_8563,N_8948);
or UO_334 (O_334,N_8629,N_9249);
and UO_335 (O_335,N_8165,N_9946);
nor UO_336 (O_336,N_9245,N_8952);
or UO_337 (O_337,N_7586,N_8702);
or UO_338 (O_338,N_9188,N_9057);
nand UO_339 (O_339,N_8935,N_9571);
and UO_340 (O_340,N_9641,N_8027);
nand UO_341 (O_341,N_8640,N_9311);
and UO_342 (O_342,N_8362,N_9450);
and UO_343 (O_343,N_9292,N_9308);
and UO_344 (O_344,N_8551,N_8843);
nor UO_345 (O_345,N_9340,N_9833);
nor UO_346 (O_346,N_8255,N_7976);
nand UO_347 (O_347,N_9157,N_9612);
nor UO_348 (O_348,N_8331,N_9264);
nand UO_349 (O_349,N_7613,N_7721);
xor UO_350 (O_350,N_8495,N_7821);
or UO_351 (O_351,N_7583,N_7966);
nand UO_352 (O_352,N_8905,N_9626);
or UO_353 (O_353,N_9525,N_8652);
and UO_354 (O_354,N_7711,N_7657);
and UO_355 (O_355,N_8579,N_9247);
and UO_356 (O_356,N_9843,N_7686);
nor UO_357 (O_357,N_7908,N_7513);
and UO_358 (O_358,N_8445,N_8057);
nand UO_359 (O_359,N_8480,N_8485);
nand UO_360 (O_360,N_7826,N_7777);
nand UO_361 (O_361,N_8760,N_9192);
or UO_362 (O_362,N_8262,N_9873);
nand UO_363 (O_363,N_9966,N_9173);
and UO_364 (O_364,N_7929,N_9832);
nand UO_365 (O_365,N_8300,N_8909);
and UO_366 (O_366,N_9884,N_9288);
nor UO_367 (O_367,N_9507,N_9688);
nand UO_368 (O_368,N_8343,N_9927);
nor UO_369 (O_369,N_7636,N_7732);
or UO_370 (O_370,N_8643,N_9036);
nand UO_371 (O_371,N_9979,N_7754);
nor UO_372 (O_372,N_8537,N_9683);
or UO_373 (O_373,N_8797,N_8234);
and UO_374 (O_374,N_9277,N_9784);
and UO_375 (O_375,N_7584,N_8872);
and UO_376 (O_376,N_8033,N_9543);
nand UO_377 (O_377,N_7811,N_9769);
and UO_378 (O_378,N_8217,N_9668);
and UO_379 (O_379,N_8827,N_8402);
and UO_380 (O_380,N_8514,N_9593);
and UO_381 (O_381,N_8167,N_9268);
or UO_382 (O_382,N_7894,N_7810);
or UO_383 (O_383,N_8000,N_9082);
or UO_384 (O_384,N_8583,N_8987);
nand UO_385 (O_385,N_7654,N_7797);
or UO_386 (O_386,N_8058,N_9901);
or UO_387 (O_387,N_7666,N_8812);
nor UO_388 (O_388,N_8185,N_9628);
xnor UO_389 (O_389,N_8274,N_9982);
xor UO_390 (O_390,N_9019,N_8588);
or UO_391 (O_391,N_8029,N_8346);
or UO_392 (O_392,N_7582,N_9595);
and UO_393 (O_393,N_8416,N_8577);
nand UO_394 (O_394,N_7708,N_8866);
and UO_395 (O_395,N_9390,N_9714);
nand UO_396 (O_396,N_9419,N_9576);
nor UO_397 (O_397,N_9721,N_9928);
nand UO_398 (O_398,N_7520,N_8980);
and UO_399 (O_399,N_9814,N_9563);
and UO_400 (O_400,N_7717,N_9046);
or UO_401 (O_401,N_8556,N_8547);
and UO_402 (O_402,N_9569,N_8528);
or UO_403 (O_403,N_9164,N_9243);
and UO_404 (O_404,N_8159,N_7524);
nand UO_405 (O_405,N_9907,N_8697);
xor UO_406 (O_406,N_9229,N_8756);
and UO_407 (O_407,N_9090,N_9275);
nor UO_408 (O_408,N_8560,N_8089);
or UO_409 (O_409,N_8953,N_9209);
nor UO_410 (O_410,N_8887,N_7726);
nor UO_411 (O_411,N_8122,N_9109);
nand UO_412 (O_412,N_9749,N_9055);
or UO_413 (O_413,N_8113,N_8794);
and UO_414 (O_414,N_8981,N_8330);
nand UO_415 (O_415,N_9695,N_7669);
nand UO_416 (O_416,N_8390,N_9396);
nor UO_417 (O_417,N_7643,N_9759);
and UO_418 (O_418,N_9283,N_8642);
and UO_419 (O_419,N_7508,N_9635);
nor UO_420 (O_420,N_9152,N_9031);
and UO_421 (O_421,N_7843,N_8956);
nor UO_422 (O_422,N_7786,N_9502);
nor UO_423 (O_423,N_8434,N_8889);
and UO_424 (O_424,N_9624,N_9371);
nor UO_425 (O_425,N_8781,N_8129);
or UO_426 (O_426,N_9697,N_8990);
nand UO_427 (O_427,N_7602,N_9909);
and UO_428 (O_428,N_8063,N_9670);
nor UO_429 (O_429,N_9760,N_9696);
nor UO_430 (O_430,N_9293,N_8061);
or UO_431 (O_431,N_8338,N_9203);
or UO_432 (O_432,N_8823,N_7842);
nor UO_433 (O_433,N_8531,N_8934);
nand UO_434 (O_434,N_8684,N_8391);
nor UO_435 (O_435,N_9953,N_7829);
nor UO_436 (O_436,N_8596,N_7678);
nand UO_437 (O_437,N_7611,N_8457);
or UO_438 (O_438,N_8311,N_9425);
nand UO_439 (O_439,N_9124,N_8266);
nand UO_440 (O_440,N_8290,N_7889);
nand UO_441 (O_441,N_9986,N_9273);
nor UO_442 (O_442,N_9837,N_9560);
nand UO_443 (O_443,N_9834,N_9698);
and UO_444 (O_444,N_9471,N_9483);
and UO_445 (O_445,N_9818,N_9363);
nand UO_446 (O_446,N_9639,N_8968);
or UO_447 (O_447,N_8972,N_7629);
xnor UO_448 (O_448,N_8933,N_8871);
or UO_449 (O_449,N_9106,N_9515);
nand UO_450 (O_450,N_9514,N_8263);
nand UO_451 (O_451,N_9180,N_8606);
or UO_452 (O_452,N_8422,N_8829);
nand UO_453 (O_453,N_7874,N_9710);
nor UO_454 (O_454,N_9150,N_8828);
nor UO_455 (O_455,N_8481,N_9851);
and UO_456 (O_456,N_7949,N_8670);
nor UO_457 (O_457,N_9473,N_8830);
nand UO_458 (O_458,N_7550,N_9993);
and UO_459 (O_459,N_8902,N_8673);
and UO_460 (O_460,N_8517,N_9439);
or UO_461 (O_461,N_9328,N_7996);
or UO_462 (O_462,N_8888,N_8114);
or UO_463 (O_463,N_9742,N_9524);
nor UO_464 (O_464,N_8676,N_9355);
nor UO_465 (O_465,N_9330,N_9788);
nor UO_466 (O_466,N_9829,N_8584);
or UO_467 (O_467,N_8372,N_7979);
nor UO_468 (O_468,N_8918,N_7684);
or UO_469 (O_469,N_9259,N_8142);
nor UO_470 (O_470,N_7507,N_8292);
and UO_471 (O_471,N_9079,N_8376);
nand UO_472 (O_472,N_8867,N_8305);
nand UO_473 (O_473,N_8706,N_9401);
nand UO_474 (O_474,N_9940,N_8228);
nor UO_475 (O_475,N_9476,N_7793);
and UO_476 (O_476,N_7502,N_9605);
or UO_477 (O_477,N_8497,N_7911);
nand UO_478 (O_478,N_9616,N_8156);
or UO_479 (O_479,N_9964,N_8807);
and UO_480 (O_480,N_9182,N_9785);
nor UO_481 (O_481,N_8126,N_7950);
nor UO_482 (O_482,N_7725,N_9400);
nor UO_483 (O_483,N_9470,N_9989);
nor UO_484 (O_484,N_9968,N_9690);
nor UO_485 (O_485,N_8833,N_9689);
nor UO_486 (O_486,N_8207,N_8757);
xnor UO_487 (O_487,N_9436,N_9580);
and UO_488 (O_488,N_8648,N_7751);
nand UO_489 (O_489,N_9651,N_9168);
or UO_490 (O_490,N_9904,N_9147);
and UO_491 (O_491,N_9657,N_7790);
nand UO_492 (O_492,N_8123,N_8246);
nor UO_493 (O_493,N_9339,N_7985);
nand UO_494 (O_494,N_9888,N_8277);
nand UO_495 (O_495,N_9026,N_9550);
or UO_496 (O_496,N_8718,N_9504);
and UO_497 (O_497,N_7933,N_7740);
and UO_498 (O_498,N_9083,N_9647);
or UO_499 (O_499,N_7695,N_8205);
nor UO_500 (O_500,N_8296,N_8307);
nand UO_501 (O_501,N_7859,N_9376);
nand UO_502 (O_502,N_7873,N_8289);
nand UO_503 (O_503,N_9603,N_8382);
or UO_504 (O_504,N_7693,N_9675);
nand UO_505 (O_505,N_8433,N_8559);
and UO_506 (O_506,N_7980,N_8153);
or UO_507 (O_507,N_9533,N_8993);
and UO_508 (O_508,N_8252,N_7753);
nor UO_509 (O_509,N_9871,N_7660);
and UO_510 (O_510,N_9310,N_9763);
and UO_511 (O_511,N_9482,N_9066);
or UO_512 (O_512,N_9103,N_9146);
or UO_513 (O_513,N_7964,N_8285);
nor UO_514 (O_514,N_9521,N_8369);
nor UO_515 (O_515,N_9868,N_9346);
nand UO_516 (O_516,N_9752,N_8117);
nor UO_517 (O_517,N_8239,N_7608);
and UO_518 (O_518,N_8216,N_8863);
or UO_519 (O_519,N_7511,N_9280);
and UO_520 (O_520,N_9044,N_9037);
and UO_521 (O_521,N_8150,N_7837);
nand UO_522 (O_522,N_9447,N_8429);
nor UO_523 (O_523,N_7649,N_8963);
nor UO_524 (O_524,N_7887,N_8195);
nand UO_525 (O_525,N_9725,N_8838);
or UO_526 (O_526,N_9226,N_8883);
or UO_527 (O_527,N_9410,N_8139);
nor UO_528 (O_528,N_9021,N_9242);
nor UO_529 (O_529,N_7604,N_8202);
or UO_530 (O_530,N_8553,N_9879);
nor UO_531 (O_531,N_7928,N_8721);
and UO_532 (O_532,N_9232,N_9583);
nand UO_533 (O_533,N_9961,N_8735);
or UO_534 (O_534,N_9078,N_9950);
or UO_535 (O_535,N_9349,N_8847);
or UO_536 (O_536,N_8194,N_8102);
or UO_537 (O_537,N_8989,N_8724);
nand UO_538 (O_538,N_7634,N_9030);
nor UO_539 (O_539,N_9876,N_8592);
nand UO_540 (O_540,N_9754,N_9354);
nand UO_541 (O_541,N_9937,N_8406);
or UO_542 (O_542,N_8611,N_8688);
and UO_543 (O_543,N_9882,N_9768);
and UO_544 (O_544,N_9246,N_9806);
nor UO_545 (O_545,N_9071,N_9520);
nor UO_546 (O_546,N_9594,N_8064);
or UO_547 (O_547,N_8538,N_8121);
nand UO_548 (O_548,N_8808,N_7825);
nor UO_549 (O_549,N_7926,N_9029);
nor UO_550 (O_550,N_9503,N_7529);
or UO_551 (O_551,N_9304,N_8915);
or UO_552 (O_552,N_8656,N_7854);
or UO_553 (O_553,N_8409,N_9976);
nor UO_554 (O_554,N_8693,N_7834);
nand UO_555 (O_555,N_8750,N_8529);
nand UO_556 (O_556,N_9313,N_9958);
and UO_557 (O_557,N_9575,N_7990);
and UO_558 (O_558,N_8677,N_8276);
and UO_559 (O_559,N_7518,N_9191);
or UO_560 (O_560,N_8522,N_8415);
and UO_561 (O_561,N_8679,N_7707);
nand UO_562 (O_562,N_7663,N_9666);
and UO_563 (O_563,N_9065,N_9591);
and UO_564 (O_564,N_7807,N_9648);
nand UO_565 (O_565,N_9585,N_8135);
nor UO_566 (O_566,N_9329,N_7858);
nor UO_567 (O_567,N_7683,N_9331);
nor UO_568 (O_568,N_8105,N_9886);
nand UO_569 (O_569,N_8715,N_8110);
or UO_570 (O_570,N_9796,N_8744);
or UO_571 (O_571,N_9006,N_8727);
nand UO_572 (O_572,N_7803,N_9931);
or UO_573 (O_573,N_8374,N_7941);
nand UO_574 (O_574,N_9859,N_8212);
nand UO_575 (O_575,N_8431,N_8613);
nand UO_576 (O_576,N_9926,N_9258);
and UO_577 (O_577,N_8026,N_9033);
nor UO_578 (O_578,N_8494,N_8612);
xor UO_579 (O_579,N_8966,N_9341);
and UO_580 (O_580,N_8784,N_8344);
nand UO_581 (O_581,N_9038,N_8282);
or UO_582 (O_582,N_9263,N_8594);
nor UO_583 (O_583,N_9115,N_7561);
nor UO_584 (O_584,N_9291,N_9526);
and UO_585 (O_585,N_8019,N_8259);
and UO_586 (O_586,N_8561,N_9684);
nand UO_587 (O_587,N_8758,N_8917);
or UO_588 (O_588,N_9938,N_8651);
nor UO_589 (O_589,N_9614,N_8503);
and UO_590 (O_590,N_7667,N_9764);
and UO_591 (O_591,N_9087,N_8976);
nand UO_592 (O_592,N_8363,N_9219);
nor UO_593 (O_593,N_8486,N_8322);
nor UO_594 (O_594,N_7954,N_8984);
or UO_595 (O_595,N_8148,N_9392);
nor UO_596 (O_596,N_8249,N_8334);
and UO_597 (O_597,N_8175,N_8303);
nand UO_598 (O_598,N_8199,N_9528);
nand UO_599 (O_599,N_9163,N_8425);
and UO_600 (O_600,N_7737,N_8708);
xor UO_601 (O_601,N_8861,N_8722);
xnor UO_602 (O_602,N_9974,N_8886);
nor UO_603 (O_603,N_9223,N_8472);
nand UO_604 (O_604,N_9960,N_8385);
and UO_605 (O_605,N_9387,N_9894);
or UO_606 (O_606,N_8779,N_8137);
nor UO_607 (O_607,N_9627,N_8180);
or UO_608 (O_608,N_8662,N_8882);
and UO_609 (O_609,N_8073,N_9381);
nand UO_610 (O_610,N_7850,N_9845);
nand UO_611 (O_611,N_8869,N_9431);
and UO_612 (O_612,N_8786,N_7917);
and UO_613 (O_613,N_8009,N_7618);
nor UO_614 (O_614,N_9140,N_7591);
and UO_615 (O_615,N_9707,N_9819);
nor UO_616 (O_616,N_9176,N_8473);
nor UO_617 (O_617,N_9237,N_9255);
and UO_618 (O_618,N_9201,N_9529);
and UO_619 (O_619,N_9004,N_8413);
nor UO_620 (O_620,N_9059,N_8074);
or UO_621 (O_621,N_8581,N_8371);
and UO_622 (O_622,N_8819,N_7893);
or UO_623 (O_623,N_7652,N_9633);
nor UO_624 (O_624,N_7633,N_9250);
nand UO_625 (O_625,N_8490,N_9477);
and UO_626 (O_626,N_8493,N_9669);
nor UO_627 (O_627,N_8272,N_8770);
or UO_628 (O_628,N_9634,N_9404);
and UO_629 (O_629,N_7750,N_8302);
nand UO_630 (O_630,N_7648,N_9091);
nor UO_631 (O_631,N_9857,N_7664);
nand UO_632 (O_632,N_7913,N_8295);
or UO_633 (O_633,N_8885,N_8320);
or UO_634 (O_634,N_7642,N_7855);
nand UO_635 (O_635,N_7533,N_8478);
nand UO_636 (O_636,N_8403,N_8265);
and UO_637 (O_637,N_9505,N_8242);
nor UO_638 (O_638,N_8170,N_7594);
nand UO_639 (O_639,N_9599,N_8999);
or UO_640 (O_640,N_7851,N_8096);
nor UO_641 (O_641,N_8663,N_9307);
and UO_642 (O_642,N_9377,N_8315);
or UO_643 (O_643,N_9016,N_9454);
or UO_644 (O_644,N_8590,N_8568);
and UO_645 (O_645,N_8840,N_9914);
nand UO_646 (O_646,N_8725,N_7600);
or UO_647 (O_647,N_8824,N_8862);
nor UO_648 (O_648,N_9214,N_9199);
and UO_649 (O_649,N_8354,N_8813);
nand UO_650 (O_650,N_9508,N_9025);
nand UO_651 (O_651,N_9416,N_7745);
and UO_652 (O_652,N_8284,N_9693);
and UO_653 (O_653,N_8396,N_7559);
nor UO_654 (O_654,N_9405,N_8555);
or UO_655 (O_655,N_9565,N_9830);
or UO_656 (O_656,N_9261,N_8814);
and UO_657 (O_657,N_8901,N_8550);
and UO_658 (O_658,N_9547,N_8240);
or UO_659 (O_659,N_7527,N_9618);
nor UO_660 (O_660,N_8864,N_7823);
nor UO_661 (O_661,N_8022,N_7570);
nand UO_662 (O_662,N_8181,N_9956);
or UO_663 (O_663,N_8608,N_8097);
nor UO_664 (O_664,N_9501,N_9121);
nand UO_665 (O_665,N_9394,N_7857);
and UO_666 (O_666,N_9389,N_7637);
nand UO_667 (O_667,N_8499,N_8644);
or UO_668 (O_668,N_9743,N_8037);
or UO_669 (O_669,N_9584,N_7871);
or UO_670 (O_670,N_9797,N_9185);
nor UO_671 (O_671,N_8842,N_8118);
nor UO_672 (O_672,N_8558,N_9941);
or UO_673 (O_673,N_9929,N_8787);
or UO_674 (O_674,N_7981,N_8378);
nand UO_675 (O_675,N_8326,N_8456);
nand UO_676 (O_676,N_9262,N_9604);
and UO_677 (O_677,N_8798,N_9238);
nor UO_678 (O_678,N_8616,N_7610);
nor UO_679 (O_679,N_9269,N_8399);
and UO_680 (O_680,N_8610,N_9333);
nor UO_681 (O_681,N_9222,N_9010);
nor UO_682 (O_682,N_9361,N_9650);
and UO_683 (O_683,N_9426,N_8130);
and UO_684 (O_684,N_9352,N_8461);
nand UO_685 (O_685,N_8081,N_9175);
nand UO_686 (O_686,N_9215,N_8597);
or UO_687 (O_687,N_9652,N_9682);
and UO_688 (O_688,N_7724,N_7682);
nand UO_689 (O_689,N_9732,N_9418);
and UO_690 (O_690,N_9637,N_9636);
nand UO_691 (O_691,N_9064,N_8271);
or UO_692 (O_692,N_8435,N_9133);
nor UO_693 (O_693,N_9870,N_9994);
or UO_694 (O_694,N_8358,N_7580);
nor UO_695 (O_695,N_8287,N_7558);
nand UO_696 (O_696,N_8230,N_9887);
and UO_697 (O_697,N_9835,N_9617);
or UO_698 (O_698,N_8567,N_8747);
or UO_699 (O_699,N_8967,N_8541);
and UO_700 (O_700,N_8477,N_8783);
or UO_701 (O_701,N_7641,N_9129);
and UO_702 (O_702,N_9284,N_9362);
nor UO_703 (O_703,N_8519,N_9622);
xnor UO_704 (O_704,N_8622,N_7907);
or UO_705 (O_705,N_9409,N_8903);
nand UO_706 (O_706,N_9924,N_9303);
and UO_707 (O_707,N_9193,N_8200);
nor UO_708 (O_708,N_9139,N_9552);
xor UO_709 (O_709,N_8459,N_8066);
and UO_710 (O_710,N_7661,N_8046);
and UO_711 (O_711,N_9939,N_8631);
and UO_712 (O_712,N_9089,N_8660);
or UO_713 (O_713,N_7992,N_9169);
and UO_714 (O_714,N_7623,N_9703);
or UO_715 (O_715,N_9254,N_7937);
nand UO_716 (O_716,N_7659,N_9910);
nor UO_717 (O_717,N_8119,N_8578);
nand UO_718 (O_718,N_8014,N_9149);
and UO_719 (O_719,N_8269,N_9646);
nor UO_720 (O_720,N_8179,N_9659);
and UO_721 (O_721,N_7784,N_9916);
nor UO_722 (O_722,N_7567,N_8730);
nand UO_723 (O_723,N_8668,N_9777);
or UO_724 (O_724,N_8441,N_8884);
or UO_725 (O_725,N_9930,N_9452);
and UO_726 (O_726,N_9935,N_9815);
or UO_727 (O_727,N_9654,N_8008);
and UO_728 (O_728,N_9704,N_9965);
nor UO_729 (O_729,N_7547,N_8100);
and UO_730 (O_730,N_8658,N_8982);
nand UO_731 (O_731,N_8626,N_9276);
and UO_732 (O_732,N_9444,N_8229);
and UO_733 (O_733,N_8455,N_9326);
or UO_734 (O_734,N_8080,N_8540);
and UO_735 (O_735,N_8496,N_7691);
nor UO_736 (O_736,N_8319,N_8532);
nor UO_737 (O_737,N_7617,N_9708);
nand UO_738 (O_738,N_9863,N_9499);
or UO_739 (O_739,N_8965,N_8428);
nor UO_740 (O_740,N_8947,N_9846);
or UO_741 (O_741,N_8844,N_7982);
and UO_742 (O_742,N_9779,N_9318);
nor UO_743 (O_743,N_8498,N_8995);
or UO_744 (O_744,N_8339,N_8401);
and UO_745 (O_745,N_8705,N_8647);
nor UO_746 (O_746,N_7909,N_9118);
and UO_747 (O_747,N_9486,N_9736);
and UO_748 (O_748,N_7779,N_9379);
and UO_749 (O_749,N_7703,N_7959);
nor UO_750 (O_750,N_9706,N_7564);
or UO_751 (O_751,N_8857,N_9342);
nor UO_752 (O_752,N_8451,N_8437);
nor UO_753 (O_753,N_8681,N_7963);
or UO_754 (O_754,N_7956,N_9480);
or UO_755 (O_755,N_8680,N_8979);
nand UO_756 (O_756,N_8892,N_9861);
nor UO_757 (O_757,N_8580,N_9217);
nand UO_758 (O_758,N_8106,N_7554);
nand UO_759 (O_759,N_7694,N_8395);
nand UO_760 (O_760,N_7997,N_9256);
nand UO_761 (O_761,N_9527,N_9891);
or UO_762 (O_762,N_8994,N_8635);
nor UO_763 (O_763,N_8936,N_8895);
nor UO_764 (O_764,N_8615,N_9925);
and UO_765 (O_765,N_9782,N_7563);
nor UO_766 (O_766,N_9490,N_8251);
or UO_767 (O_767,N_8552,N_7640);
nand UO_768 (O_768,N_8021,N_8233);
nand UO_769 (O_769,N_8881,N_9653);
and UO_770 (O_770,N_7526,N_9805);
nor UO_771 (O_771,N_7895,N_9997);
nand UO_772 (O_772,N_8003,N_9063);
or UO_773 (O_773,N_7994,N_9186);
or UO_774 (O_774,N_9144,N_8694);
nand UO_775 (O_775,N_9716,N_9902);
and UO_776 (O_776,N_8618,N_9062);
or UO_777 (O_777,N_8005,N_8278);
nand UO_778 (O_778,N_8800,N_9160);
and UO_779 (O_779,N_8209,N_7939);
nor UO_780 (O_780,N_7946,N_8851);
nand UO_781 (O_781,N_9224,N_7706);
nand UO_782 (O_782,N_8780,N_8304);
or UO_783 (O_783,N_9111,N_7940);
nand UO_784 (O_784,N_8633,N_8682);
nor UO_785 (O_785,N_9681,N_9810);
and UO_786 (O_786,N_8108,N_8236);
nand UO_787 (O_787,N_9880,N_8743);
or UO_788 (O_788,N_8328,N_9915);
or UO_789 (O_789,N_9984,N_9105);
nand UO_790 (O_790,N_7540,N_8894);
and UO_791 (O_791,N_8357,N_9600);
nor UO_792 (O_792,N_9715,N_8204);
nor UO_793 (O_793,N_9386,N_7553);
nand UO_794 (O_794,N_9382,N_8039);
nand UO_795 (O_795,N_9587,N_7734);
or UO_796 (O_796,N_8244,N_9821);
nand UO_797 (O_797,N_8423,N_9432);
and UO_798 (O_798,N_8831,N_9305);
and UO_799 (O_799,N_8685,N_7712);
nor UO_800 (O_800,N_7931,N_8667);
nor UO_801 (O_801,N_9739,N_8931);
nand UO_802 (O_802,N_7836,N_9995);
and UO_803 (O_803,N_9009,N_9282);
or UO_804 (O_804,N_8329,N_8226);
or UO_805 (O_805,N_8527,N_7890);
or UO_806 (O_806,N_8280,N_9434);
or UO_807 (O_807,N_9538,N_9808);
nor UO_808 (O_808,N_8267,N_7542);
or UO_809 (O_809,N_8317,N_8324);
nor UO_810 (O_810,N_9745,N_8609);
nor UO_811 (O_811,N_9606,N_9803);
nor UO_812 (O_812,N_8695,N_9122);
or UO_813 (O_813,N_8410,N_8049);
nand UO_814 (O_814,N_8450,N_9542);
nand UO_815 (O_815,N_9154,N_9878);
nand UO_816 (O_816,N_8489,N_9457);
nor UO_817 (O_817,N_7986,N_7862);
nor UO_818 (O_818,N_9597,N_8007);
and UO_819 (O_819,N_8564,N_9744);
and UO_820 (O_820,N_8060,N_8711);
and UO_821 (O_821,N_8440,N_8098);
and UO_822 (O_822,N_8991,N_7719);
or UO_823 (O_823,N_7844,N_7744);
nand UO_824 (O_824,N_9384,N_9874);
nand UO_825 (O_825,N_8562,N_9012);
nand UO_826 (O_826,N_9257,N_9638);
nor UO_827 (O_827,N_8763,N_9335);
and UO_828 (O_828,N_8365,N_7692);
nand UO_829 (O_829,N_8134,N_9975);
and UO_830 (O_830,N_8738,N_9167);
nand UO_831 (O_831,N_8397,N_7919);
nand UO_832 (O_832,N_9177,N_9848);
nor UO_833 (O_833,N_7589,N_9336);
or UO_834 (O_834,N_8458,N_8465);
and UO_835 (O_835,N_7536,N_9045);
nand UO_836 (O_836,N_8928,N_8649);
or UO_837 (O_837,N_8878,N_9551);
nand UO_838 (O_838,N_9534,N_7500);
and UO_839 (O_839,N_8254,N_9151);
and UO_840 (O_840,N_7514,N_7883);
nor UO_841 (O_841,N_9770,N_9357);
nor UO_842 (O_842,N_9314,N_8943);
or UO_843 (O_843,N_8992,N_9955);
and UO_844 (O_844,N_7505,N_9451);
or UO_845 (O_845,N_9445,N_9840);
nand UO_846 (O_846,N_9001,N_9988);
nor UO_847 (O_847,N_7670,N_7551);
nand UO_848 (O_848,N_8157,N_9737);
nor UO_849 (O_849,N_7535,N_9479);
or UO_850 (O_850,N_8443,N_9295);
nor UO_851 (O_851,N_9068,N_9302);
or UO_852 (O_852,N_7953,N_9536);
and UO_853 (O_853,N_9195,N_8215);
or UO_854 (O_854,N_8913,N_8442);
or UO_855 (O_855,N_9220,N_8247);
nand UO_856 (O_856,N_8492,N_8316);
and UO_857 (O_857,N_8811,N_7789);
nand UO_858 (O_858,N_8222,N_7773);
and UO_859 (O_859,N_8739,N_9934);
and UO_860 (O_860,N_7853,N_8421);
nor UO_861 (O_861,N_8937,N_7962);
or UO_862 (O_862,N_7847,N_9942);
and UO_863 (O_863,N_7614,N_9812);
or UO_864 (O_864,N_9912,N_9919);
and UO_865 (O_865,N_8678,N_7690);
or UO_866 (O_866,N_8268,N_8951);
nor UO_867 (O_867,N_8998,N_9466);
nand UO_868 (O_868,N_8802,N_9013);
and UO_869 (O_869,N_9816,N_9847);
and UO_870 (O_870,N_8092,N_9438);
nand UO_871 (O_871,N_9343,N_8516);
or UO_872 (O_872,N_9724,N_9954);
xor UO_873 (O_873,N_9225,N_9374);
nor UO_874 (O_874,N_7606,N_9801);
nand UO_875 (O_875,N_9353,N_8768);
or UO_876 (O_876,N_8539,N_9645);
nand UO_877 (O_877,N_9677,N_9674);
and UO_878 (O_878,N_8203,N_8774);
nand UO_879 (O_879,N_7814,N_9040);
and UO_880 (O_880,N_8930,N_9162);
nand UO_881 (O_881,N_8025,N_8041);
nand UO_882 (O_882,N_9811,N_7897);
nand UO_883 (O_883,N_7952,N_8659);
nand UO_884 (O_884,N_8923,N_9983);
nand UO_885 (O_885,N_8716,N_8467);
or UO_886 (O_886,N_9189,N_8291);
nand UO_887 (O_887,N_9135,N_9963);
nand UO_888 (O_888,N_7596,N_7886);
or UO_889 (O_889,N_9920,N_8776);
nor UO_890 (O_890,N_9197,N_8723);
and UO_891 (O_891,N_9170,N_8958);
and UO_892 (O_892,N_9491,N_9213);
nor UO_893 (O_893,N_9981,N_8900);
and UO_894 (O_894,N_8191,N_8825);
nand UO_895 (O_895,N_8312,N_9817);
or UO_896 (O_896,N_8955,N_9233);
or UO_897 (O_897,N_8235,N_8177);
nand UO_898 (O_898,N_8771,N_9235);
nor UO_899 (O_899,N_8107,N_8848);
nor UO_900 (O_900,N_9535,N_9844);
and UO_901 (O_901,N_9369,N_7910);
or UO_902 (O_902,N_8245,N_9673);
and UO_903 (O_903,N_7892,N_9776);
and UO_904 (O_904,N_9751,N_7925);
nor UO_905 (O_905,N_8151,N_8530);
nand UO_906 (O_906,N_8427,N_9049);
or UO_907 (O_907,N_8373,N_7668);
or UO_908 (O_908,N_8638,N_8717);
and UO_909 (O_909,N_9783,N_9465);
and UO_910 (O_910,N_7599,N_9665);
and UO_911 (O_911,N_8983,N_8031);
nor UO_912 (O_912,N_9306,N_8438);
nand UO_913 (O_913,N_7679,N_9131);
nor UO_914 (O_914,N_8765,N_9885);
nor UO_915 (O_915,N_8941,N_8852);
nor UO_916 (O_916,N_9510,N_8006);
nand UO_917 (O_917,N_9205,N_7650);
nand UO_918 (O_918,N_7681,N_8792);
nor UO_919 (O_919,N_8932,N_8059);
nor UO_920 (O_920,N_9554,N_8115);
and UO_921 (O_921,N_8032,N_8605);
and UO_922 (O_922,N_9281,N_9159);
nor UO_923 (O_923,N_8361,N_7519);
nand UO_924 (O_924,N_7878,N_7702);
nor UO_925 (O_925,N_9631,N_8487);
and UO_926 (O_926,N_8510,N_7771);
and UO_927 (O_927,N_8471,N_8873);
and UO_928 (O_928,N_8193,N_9086);
nor UO_929 (O_929,N_8018,N_8545);
or UO_930 (O_930,N_7626,N_8593);
nand UO_931 (O_931,N_7965,N_9774);
and UO_932 (O_932,N_9948,N_9110);
and UO_933 (O_933,N_9971,N_7704);
nor UO_934 (O_934,N_8085,N_7605);
and UO_935 (O_935,N_8090,N_8707);
nand UO_936 (O_936,N_8542,N_9826);
nor UO_937 (O_937,N_8420,N_9853);
nand UO_938 (O_938,N_8853,N_8125);
or UO_939 (O_939,N_9917,N_9117);
nand UO_940 (O_940,N_7866,N_8961);
nor UO_941 (O_941,N_8617,N_8879);
or UO_942 (O_942,N_9081,N_7815);
or UO_943 (O_943,N_8761,N_9793);
nor UO_944 (O_944,N_8162,N_9592);
or UO_945 (O_945,N_8035,N_8084);
nor UO_946 (O_946,N_9828,N_8184);
nor UO_947 (O_947,N_7509,N_8308);
nor UO_948 (O_948,N_7539,N_8258);
nor UO_949 (O_949,N_8549,N_8960);
or UO_950 (O_950,N_7792,N_9084);
xnor UO_951 (O_951,N_9671,N_9822);
nand UO_952 (O_952,N_7728,N_8741);
nand UO_953 (O_953,N_9061,N_9375);
nand UO_954 (O_954,N_9897,N_8436);
and UO_955 (O_955,N_8986,N_7718);
and UO_956 (O_956,N_8389,N_7597);
nand UO_957 (O_957,N_9428,N_9772);
or UO_958 (O_958,N_8591,N_8248);
nand UO_959 (O_959,N_9667,N_9740);
or UO_960 (O_960,N_7556,N_7676);
nand UO_961 (O_961,N_7701,N_8043);
nor UO_962 (O_962,N_8366,N_8067);
nand UO_963 (O_963,N_9422,N_8484);
nand UO_964 (O_964,N_7870,N_7772);
nor UO_965 (O_965,N_7852,N_8975);
nor UO_966 (O_966,N_8210,N_7575);
nand UO_967 (O_967,N_8740,N_7785);
nand UO_968 (O_968,N_8384,N_9467);
and UO_969 (O_969,N_8112,N_9274);
and UO_970 (O_970,N_8068,N_9022);
nand UO_971 (O_971,N_7665,N_8463);
and UO_972 (O_972,N_7856,N_9108);
nand UO_973 (O_973,N_8826,N_9596);
and UO_974 (O_974,N_7824,N_8775);
nand UO_975 (O_975,N_8293,N_8004);
nand UO_976 (O_976,N_8742,N_8250);
nor UO_977 (O_977,N_7827,N_8712);
and UO_978 (O_978,N_9933,N_8036);
nand UO_979 (O_979,N_7720,N_9544);
or UO_980 (O_980,N_9437,N_9702);
or UO_981 (O_981,N_9589,N_8858);
nand UO_982 (O_982,N_7673,N_8636);
nand UO_983 (O_983,N_7697,N_7885);
and UO_984 (O_984,N_8646,N_7819);
nand UO_985 (O_985,N_8754,N_8359);
xor UO_986 (O_986,N_8171,N_9630);
and UO_987 (O_987,N_9443,N_9548);
or UO_988 (O_988,N_8924,N_7778);
and UO_989 (O_989,N_9672,N_9208);
nand UO_990 (O_990,N_9323,N_9557);
nand UO_991 (O_991,N_9042,N_7912);
nor UO_992 (O_992,N_8585,N_7920);
nand UO_993 (O_993,N_8404,N_8942);
or UO_994 (O_994,N_9184,N_9663);
and UO_995 (O_995,N_7999,N_7800);
nor UO_996 (O_996,N_8772,N_7805);
nor UO_997 (O_997,N_8367,N_7579);
or UO_998 (O_998,N_9315,N_9570);
nor UO_999 (O_999,N_8675,N_9632);
or UO_1000 (O_1000,N_7538,N_9687);
or UO_1001 (O_1001,N_8172,N_7865);
nand UO_1002 (O_1002,N_9545,N_9252);
and UO_1003 (O_1003,N_9412,N_9385);
nor UO_1004 (O_1004,N_9461,N_7739);
and UO_1005 (O_1005,N_7560,N_7875);
nor UO_1006 (O_1006,N_8219,N_8183);
nor UO_1007 (O_1007,N_9522,N_7671);
and UO_1008 (O_1008,N_9206,N_8974);
nor UO_1009 (O_1009,N_7517,N_7881);
nand UO_1010 (O_1010,N_9350,N_8020);
nand UO_1011 (O_1011,N_9722,N_9460);
and UO_1012 (O_1012,N_9358,N_9271);
xnor UO_1013 (O_1013,N_8044,N_8447);
and UO_1014 (O_1014,N_8462,N_8569);
nand UO_1015 (O_1015,N_7960,N_8086);
nor UO_1016 (O_1016,N_7531,N_8474);
nand UO_1017 (O_1017,N_8733,N_7506);
and UO_1018 (O_1018,N_9717,N_9000);
and UO_1019 (O_1019,N_7984,N_8387);
nor UO_1020 (O_1020,N_8634,N_9187);
and UO_1021 (O_1021,N_8554,N_9137);
nor UO_1022 (O_1022,N_9067,N_8515);
and UO_1023 (O_1023,N_7672,N_7839);
nor UO_1024 (O_1024,N_9143,N_8253);
and UO_1025 (O_1025,N_8949,N_9494);
nand UO_1026 (O_1026,N_9623,N_8911);
nand UO_1027 (O_1027,N_9869,N_7915);
nor UO_1028 (O_1028,N_8726,N_8448);
and UO_1029 (O_1029,N_8386,N_7675);
nor UO_1030 (O_1030,N_9051,N_7833);
and UO_1031 (O_1031,N_7958,N_9158);
or UO_1032 (O_1032,N_8908,N_9799);
nand UO_1033 (O_1033,N_8954,N_8350);
and UO_1034 (O_1034,N_9611,N_7775);
or UO_1035 (O_1035,N_9181,N_9896);
nand UO_1036 (O_1036,N_9120,N_7530);
nor UO_1037 (O_1037,N_7974,N_9388);
nor UO_1038 (O_1038,N_9459,N_8719);
and UO_1039 (O_1039,N_9492,N_9455);
or UO_1040 (O_1040,N_7848,N_8919);
and UO_1041 (O_1041,N_9598,N_9240);
nor UO_1042 (O_1042,N_9088,N_8446);
or UO_1043 (O_1043,N_8189,N_7646);
and UO_1044 (O_1044,N_8689,N_9286);
nand UO_1045 (O_1045,N_8273,N_8671);
nand UO_1046 (O_1046,N_9568,N_8145);
or UO_1047 (O_1047,N_8837,N_8700);
xnor UO_1048 (O_1048,N_7523,N_8571);
nor UO_1049 (O_1049,N_7552,N_7769);
and UO_1050 (O_1050,N_9790,N_8945);
or UO_1051 (O_1051,N_7831,N_9723);
nor UO_1052 (O_1052,N_8078,N_8336);
nor UO_1053 (O_1053,N_9765,N_8101);
and UO_1054 (O_1054,N_9383,N_8452);
and UO_1055 (O_1055,N_8962,N_9549);
and UO_1056 (O_1056,N_9462,N_9621);
nor UO_1057 (O_1057,N_9746,N_8988);
nor UO_1058 (O_1058,N_7730,N_8408);
nor UO_1059 (O_1059,N_9967,N_9608);
or UO_1060 (O_1060,N_8475,N_9075);
nor UO_1061 (O_1061,N_9153,N_8657);
and UO_1062 (O_1062,N_9098,N_8050);
or UO_1063 (O_1063,N_9947,N_7501);
nor UO_1064 (O_1064,N_8001,N_7638);
nor UO_1065 (O_1065,N_9430,N_9423);
and UO_1066 (O_1066,N_9442,N_9867);
nor UO_1067 (O_1067,N_7796,N_9719);
nor UO_1068 (O_1068,N_8978,N_9190);
nand UO_1069 (O_1069,N_9644,N_9619);
nand UO_1070 (O_1070,N_8566,N_8377);
nand UO_1071 (O_1071,N_7741,N_7696);
nor UO_1072 (O_1072,N_7787,N_9196);
nand UO_1073 (O_1073,N_9820,N_7924);
nor UO_1074 (O_1074,N_8201,N_7989);
or UO_1075 (O_1075,N_7900,N_8920);
nand UO_1076 (O_1076,N_7729,N_9913);
and UO_1077 (O_1077,N_8454,N_9701);
nand UO_1078 (O_1078,N_8147,N_8220);
nor UO_1079 (O_1079,N_8168,N_7503);
and UO_1080 (O_1080,N_8476,N_8453);
nor UO_1081 (O_1081,N_8160,N_9655);
or UO_1082 (O_1082,N_7978,N_9128);
or UO_1083 (O_1083,N_8856,N_8116);
or UO_1084 (O_1084,N_9433,N_9440);
nand UO_1085 (O_1085,N_8355,N_8182);
nand UO_1086 (O_1086,N_9578,N_8187);
and UO_1087 (O_1087,N_9402,N_8103);
nand UO_1088 (O_1088,N_7783,N_8111);
or UO_1089 (O_1089,N_9178,N_7645);
or UO_1090 (O_1090,N_9978,N_8380);
or UO_1091 (O_1091,N_8186,N_7970);
nand UO_1092 (O_1092,N_8753,N_8701);
or UO_1093 (O_1093,N_9408,N_7788);
nor UO_1094 (O_1094,N_9018,N_9911);
nor UO_1095 (O_1095,N_9054,N_9588);
and UO_1096 (O_1096,N_8865,N_8944);
nand UO_1097 (O_1097,N_9155,N_8511);
nand UO_1098 (O_1098,N_9558,N_8325);
or UO_1099 (O_1099,N_7765,N_9881);
nand UO_1100 (O_1100,N_7942,N_9290);
and UO_1101 (O_1101,N_8042,N_9523);
nor UO_1102 (O_1102,N_8703,N_7916);
and UO_1103 (O_1103,N_8206,N_9757);
and UO_1104 (O_1104,N_8912,N_8146);
nand UO_1105 (O_1105,N_9720,N_8136);
nand UO_1106 (O_1106,N_9231,N_9325);
nor UO_1107 (O_1107,N_8729,N_9125);
nand UO_1108 (O_1108,N_9364,N_8699);
nor UO_1109 (O_1109,N_8002,N_8607);
or UO_1110 (O_1110,N_7945,N_9297);
nor UO_1111 (O_1111,N_9489,N_8318);
nor UO_1112 (O_1112,N_9513,N_8208);
and UO_1113 (O_1113,N_9546,N_8846);
or UO_1114 (O_1114,N_7932,N_7755);
and UO_1115 (O_1115,N_9506,N_7578);
nand UO_1116 (O_1116,N_9498,N_8238);
xor UO_1117 (O_1117,N_8907,N_7723);
or UO_1118 (O_1118,N_7574,N_8012);
nand UO_1119 (O_1119,N_9344,N_7804);
or UO_1120 (O_1120,N_7760,N_9076);
nor UO_1121 (O_1121,N_9566,N_7656);
and UO_1122 (O_1122,N_8655,N_9996);
nor UO_1123 (O_1123,N_7546,N_8313);
or UO_1124 (O_1124,N_8174,N_9072);
nand UO_1125 (O_1125,N_9572,N_9227);
or UO_1126 (O_1126,N_9694,N_9348);
nor UO_1127 (O_1127,N_7860,N_7888);
and UO_1128 (O_1128,N_8737,N_9142);
or UO_1129 (O_1129,N_9581,N_8939);
or UO_1130 (O_1130,N_9718,N_8053);
nand UO_1131 (O_1131,N_9824,N_9761);
nor UO_1132 (O_1132,N_9735,N_9866);
nand UO_1133 (O_1133,N_7799,N_9356);
nand UO_1134 (O_1134,N_8849,N_8832);
nor UO_1135 (O_1135,N_7822,N_8257);
or UO_1136 (O_1136,N_9495,N_8672);
nand UO_1137 (O_1137,N_8281,N_7955);
and UO_1138 (O_1138,N_7840,N_8279);
and UO_1139 (O_1139,N_8789,N_8124);
and UO_1140 (O_1140,N_7699,N_9011);
nor UO_1141 (O_1141,N_9136,N_9762);
nor UO_1142 (O_1142,N_9127,N_8710);
xor UO_1143 (O_1143,N_9747,N_7573);
or UO_1144 (O_1144,N_9936,N_9312);
or UO_1145 (O_1145,N_9775,N_9791);
or UO_1146 (O_1146,N_8483,N_8777);
or UO_1147 (O_1147,N_8623,N_8791);
or UO_1148 (O_1148,N_8627,N_9058);
or UO_1149 (O_1149,N_7998,N_9864);
nand UO_1150 (O_1150,N_8959,N_8543);
or UO_1151 (O_1151,N_9456,N_9951);
nor UO_1152 (O_1152,N_8347,N_9077);
or UO_1153 (O_1153,N_8306,N_8337);
nand UO_1154 (O_1154,N_8071,N_9474);
nor UO_1155 (O_1155,N_7930,N_8875);
or UO_1156 (O_1156,N_7644,N_8323);
nand UO_1157 (O_1157,N_8218,N_9509);
nand UO_1158 (O_1158,N_9007,N_8533);
or UO_1159 (O_1159,N_7685,N_8502);
nand UO_1160 (O_1160,N_8040,N_7749);
nor UO_1161 (O_1161,N_9727,N_8602);
nand UO_1162 (O_1162,N_8603,N_9074);
nand UO_1163 (O_1163,N_7971,N_8525);
nor UO_1164 (O_1164,N_9028,N_9053);
nor UO_1165 (O_1165,N_8400,N_9553);
or UO_1166 (O_1166,N_8352,N_7722);
nor UO_1167 (O_1167,N_9485,N_8298);
or UO_1168 (O_1168,N_8072,N_8803);
nand UO_1169 (O_1169,N_7748,N_7877);
or UO_1170 (O_1170,N_8524,N_8439);
and UO_1171 (O_1171,N_8624,N_8520);
or UO_1172 (O_1172,N_8297,N_7809);
nor UO_1173 (O_1173,N_8793,N_9360);
nand UO_1174 (O_1174,N_8128,N_8024);
nor UO_1175 (O_1175,N_8906,N_8650);
nor UO_1176 (O_1176,N_8070,N_9429);
nand UO_1177 (O_1177,N_8158,N_7861);
nor UO_1178 (O_1178,N_8405,N_8028);
or UO_1179 (O_1179,N_8709,N_9449);
and UO_1180 (O_1180,N_9836,N_8600);
or UO_1181 (O_1181,N_7557,N_8645);
and UO_1182 (O_1182,N_8821,N_7585);
or UO_1183 (O_1183,N_8630,N_9165);
and UO_1184 (O_1184,N_8321,N_9039);
and UO_1185 (O_1185,N_9991,N_7846);
nand UO_1186 (O_1186,N_8916,N_9564);
nor UO_1187 (O_1187,N_8686,N_8834);
nor UO_1188 (O_1188,N_7522,N_8426);
or UO_1189 (O_1189,N_9484,N_8698);
or UO_1190 (O_1190,N_7768,N_7758);
nor UO_1191 (O_1191,N_8356,N_9141);
nand UO_1192 (O_1192,N_9642,N_9738);
or UO_1193 (O_1193,N_9537,N_8034);
nor UO_1194 (O_1194,N_9427,N_9758);
and UO_1195 (O_1195,N_9980,N_9299);
and UO_1196 (O_1196,N_8011,N_8870);
nand UO_1197 (O_1197,N_9041,N_8491);
nor UO_1198 (O_1198,N_9321,N_7532);
and UO_1199 (O_1199,N_8309,N_8345);
or UO_1200 (O_1200,N_8163,N_7736);
nor UO_1201 (O_1201,N_9123,N_7639);
nand UO_1202 (O_1202,N_8393,N_9872);
and UO_1203 (O_1203,N_9248,N_8348);
and UO_1204 (O_1204,N_8038,N_9629);
and UO_1205 (O_1205,N_9093,N_8755);
and UO_1206 (O_1206,N_7565,N_9903);
nor UO_1207 (O_1207,N_7934,N_8896);
nor UO_1208 (O_1208,N_9883,N_7630);
nand UO_1209 (O_1209,N_8546,N_9320);
nand UO_1210 (O_1210,N_7710,N_8691);
and UO_1211 (O_1211,N_8013,N_7587);
xor UO_1212 (O_1212,N_9780,N_7867);
nor UO_1213 (O_1213,N_8641,N_9602);
nand UO_1214 (O_1214,N_9212,N_8927);
nor UO_1215 (O_1215,N_7658,N_7541);
and UO_1216 (O_1216,N_7756,N_9766);
and UO_1217 (O_1217,N_8379,N_7612);
and UO_1218 (O_1218,N_8143,N_9577);
or UO_1219 (O_1219,N_9463,N_8574);
nand UO_1220 (O_1220,N_7715,N_7705);
nor UO_1221 (O_1221,N_9511,N_7601);
or UO_1222 (O_1222,N_9366,N_9985);
or UO_1223 (O_1223,N_7983,N_8985);
nor UO_1224 (O_1224,N_9421,N_7774);
nand UO_1225 (O_1225,N_7548,N_7571);
or UO_1226 (O_1226,N_8104,N_8782);
or UO_1227 (O_1227,N_9002,N_7947);
nor UO_1228 (O_1228,N_8466,N_7615);
nor UO_1229 (O_1229,N_8573,N_8232);
xnor UO_1230 (O_1230,N_9487,N_8227);
nand UO_1231 (O_1231,N_8341,N_9253);
and UO_1232 (O_1232,N_9228,N_7957);
or UO_1233 (O_1233,N_9183,N_8464);
nand UO_1234 (O_1234,N_7674,N_9270);
nor UO_1235 (O_1235,N_9458,N_7687);
or UO_1236 (O_1236,N_8804,N_9113);
or UO_1237 (O_1237,N_9148,N_8595);
or UO_1238 (O_1238,N_8460,N_9138);
nor UO_1239 (O_1239,N_8893,N_8785);
nand UO_1240 (O_1240,N_9130,N_8444);
nor UO_1241 (O_1241,N_8173,N_7766);
and UO_1242 (O_1242,N_7662,N_8713);
and UO_1243 (O_1243,N_9266,N_9831);
nor UO_1244 (O_1244,N_8666,N_7975);
or UO_1245 (O_1245,N_9574,N_7713);
or UO_1246 (O_1246,N_9014,N_8809);
nand UO_1247 (O_1247,N_8850,N_9601);
or UO_1248 (O_1248,N_9194,N_8127);
nor UO_1249 (O_1249,N_9289,N_8314);
or UO_1250 (O_1250,N_8157,N_7567);
nor UO_1251 (O_1251,N_9479,N_9433);
and UO_1252 (O_1252,N_8148,N_9646);
xor UO_1253 (O_1253,N_8661,N_9630);
and UO_1254 (O_1254,N_9657,N_9514);
or UO_1255 (O_1255,N_8633,N_9341);
nor UO_1256 (O_1256,N_7927,N_8393);
or UO_1257 (O_1257,N_7743,N_8833);
nand UO_1258 (O_1258,N_9330,N_8774);
or UO_1259 (O_1259,N_8448,N_9495);
or UO_1260 (O_1260,N_8155,N_8165);
or UO_1261 (O_1261,N_7956,N_7916);
and UO_1262 (O_1262,N_8259,N_7873);
or UO_1263 (O_1263,N_7969,N_9291);
nor UO_1264 (O_1264,N_9264,N_8472);
xor UO_1265 (O_1265,N_9229,N_9930);
nor UO_1266 (O_1266,N_8951,N_7819);
or UO_1267 (O_1267,N_8935,N_8383);
nand UO_1268 (O_1268,N_7958,N_7931);
nand UO_1269 (O_1269,N_8322,N_9162);
and UO_1270 (O_1270,N_8411,N_8311);
nor UO_1271 (O_1271,N_9435,N_7690);
nand UO_1272 (O_1272,N_7841,N_7637);
or UO_1273 (O_1273,N_8435,N_9709);
or UO_1274 (O_1274,N_8383,N_8461);
and UO_1275 (O_1275,N_8668,N_9119);
or UO_1276 (O_1276,N_8009,N_8462);
or UO_1277 (O_1277,N_8406,N_9772);
nor UO_1278 (O_1278,N_8142,N_9333);
nand UO_1279 (O_1279,N_8750,N_9870);
nor UO_1280 (O_1280,N_7623,N_8249);
nand UO_1281 (O_1281,N_8753,N_7713);
or UO_1282 (O_1282,N_9647,N_8116);
nor UO_1283 (O_1283,N_7714,N_9550);
or UO_1284 (O_1284,N_9179,N_9205);
or UO_1285 (O_1285,N_8380,N_9021);
nor UO_1286 (O_1286,N_9871,N_7812);
or UO_1287 (O_1287,N_8011,N_8102);
nand UO_1288 (O_1288,N_8198,N_7928);
nor UO_1289 (O_1289,N_9281,N_8263);
and UO_1290 (O_1290,N_8038,N_8922);
or UO_1291 (O_1291,N_8214,N_8680);
nand UO_1292 (O_1292,N_8198,N_8902);
and UO_1293 (O_1293,N_9141,N_8967);
nand UO_1294 (O_1294,N_9433,N_9571);
nor UO_1295 (O_1295,N_7645,N_9818);
and UO_1296 (O_1296,N_9851,N_7532);
or UO_1297 (O_1297,N_8705,N_9065);
nor UO_1298 (O_1298,N_8068,N_8789);
or UO_1299 (O_1299,N_9522,N_7882);
nand UO_1300 (O_1300,N_8338,N_7695);
and UO_1301 (O_1301,N_7520,N_8725);
nand UO_1302 (O_1302,N_9537,N_9526);
nand UO_1303 (O_1303,N_9023,N_9131);
nand UO_1304 (O_1304,N_7602,N_7822);
or UO_1305 (O_1305,N_9817,N_9577);
nor UO_1306 (O_1306,N_9395,N_9300);
or UO_1307 (O_1307,N_9555,N_8463);
and UO_1308 (O_1308,N_8316,N_9425);
or UO_1309 (O_1309,N_8022,N_7868);
and UO_1310 (O_1310,N_9321,N_7900);
nor UO_1311 (O_1311,N_9016,N_7637);
nand UO_1312 (O_1312,N_8276,N_7530);
nor UO_1313 (O_1313,N_7845,N_9421);
nand UO_1314 (O_1314,N_7955,N_7850);
or UO_1315 (O_1315,N_9809,N_9981);
nand UO_1316 (O_1316,N_8682,N_8765);
and UO_1317 (O_1317,N_8386,N_8646);
and UO_1318 (O_1318,N_8880,N_9785);
or UO_1319 (O_1319,N_9447,N_8935);
nand UO_1320 (O_1320,N_8202,N_9342);
nor UO_1321 (O_1321,N_8483,N_9168);
and UO_1322 (O_1322,N_9624,N_9469);
nand UO_1323 (O_1323,N_8084,N_8783);
nor UO_1324 (O_1324,N_8453,N_7712);
and UO_1325 (O_1325,N_8987,N_8140);
or UO_1326 (O_1326,N_9302,N_9714);
and UO_1327 (O_1327,N_8418,N_9870);
nor UO_1328 (O_1328,N_7886,N_9411);
and UO_1329 (O_1329,N_9869,N_9223);
nand UO_1330 (O_1330,N_7907,N_8511);
nand UO_1331 (O_1331,N_8899,N_9823);
or UO_1332 (O_1332,N_9816,N_8726);
and UO_1333 (O_1333,N_9782,N_9343);
and UO_1334 (O_1334,N_7868,N_9581);
and UO_1335 (O_1335,N_8792,N_9450);
or UO_1336 (O_1336,N_8717,N_8937);
or UO_1337 (O_1337,N_8043,N_9883);
nor UO_1338 (O_1338,N_7842,N_9249);
or UO_1339 (O_1339,N_8955,N_8564);
and UO_1340 (O_1340,N_9986,N_9343);
nand UO_1341 (O_1341,N_8279,N_9509);
and UO_1342 (O_1342,N_8777,N_9493);
nor UO_1343 (O_1343,N_9866,N_8135);
or UO_1344 (O_1344,N_7860,N_9765);
nor UO_1345 (O_1345,N_7991,N_8123);
and UO_1346 (O_1346,N_8265,N_9483);
nand UO_1347 (O_1347,N_7538,N_8743);
and UO_1348 (O_1348,N_9196,N_9338);
nand UO_1349 (O_1349,N_8467,N_9687);
or UO_1350 (O_1350,N_8861,N_9071);
or UO_1351 (O_1351,N_8093,N_7737);
and UO_1352 (O_1352,N_9833,N_8468);
and UO_1353 (O_1353,N_9368,N_9856);
nand UO_1354 (O_1354,N_9800,N_8350);
or UO_1355 (O_1355,N_8066,N_8886);
nand UO_1356 (O_1356,N_9581,N_8066);
nor UO_1357 (O_1357,N_9672,N_9865);
and UO_1358 (O_1358,N_9573,N_8688);
nor UO_1359 (O_1359,N_9906,N_8041);
or UO_1360 (O_1360,N_9828,N_8743);
nor UO_1361 (O_1361,N_8545,N_7788);
nand UO_1362 (O_1362,N_9695,N_8042);
nor UO_1363 (O_1363,N_9228,N_7881);
or UO_1364 (O_1364,N_8341,N_8885);
and UO_1365 (O_1365,N_9433,N_8430);
nand UO_1366 (O_1366,N_7801,N_9482);
nor UO_1367 (O_1367,N_8977,N_9518);
nand UO_1368 (O_1368,N_7895,N_8944);
and UO_1369 (O_1369,N_9886,N_8995);
nand UO_1370 (O_1370,N_8785,N_9187);
or UO_1371 (O_1371,N_8266,N_9393);
nand UO_1372 (O_1372,N_7617,N_8807);
or UO_1373 (O_1373,N_9711,N_9208);
nor UO_1374 (O_1374,N_9751,N_8140);
or UO_1375 (O_1375,N_8849,N_8790);
nand UO_1376 (O_1376,N_8516,N_8013);
nor UO_1377 (O_1377,N_8017,N_7519);
nor UO_1378 (O_1378,N_8162,N_8719);
nor UO_1379 (O_1379,N_9342,N_9210);
nand UO_1380 (O_1380,N_7819,N_8175);
and UO_1381 (O_1381,N_9101,N_8930);
or UO_1382 (O_1382,N_7928,N_8942);
and UO_1383 (O_1383,N_9745,N_8346);
nor UO_1384 (O_1384,N_8127,N_8588);
nand UO_1385 (O_1385,N_7766,N_7518);
and UO_1386 (O_1386,N_7767,N_9215);
and UO_1387 (O_1387,N_7784,N_8876);
or UO_1388 (O_1388,N_9156,N_7558);
and UO_1389 (O_1389,N_9482,N_8573);
nor UO_1390 (O_1390,N_7523,N_8743);
nor UO_1391 (O_1391,N_9648,N_9142);
xnor UO_1392 (O_1392,N_9949,N_7561);
and UO_1393 (O_1393,N_8374,N_9674);
nand UO_1394 (O_1394,N_9021,N_9012);
and UO_1395 (O_1395,N_9631,N_7987);
or UO_1396 (O_1396,N_9761,N_8666);
nor UO_1397 (O_1397,N_7857,N_7747);
or UO_1398 (O_1398,N_8799,N_7584);
nand UO_1399 (O_1399,N_9499,N_9173);
nor UO_1400 (O_1400,N_9070,N_8206);
or UO_1401 (O_1401,N_8968,N_8604);
nor UO_1402 (O_1402,N_8938,N_7974);
and UO_1403 (O_1403,N_7720,N_9720);
and UO_1404 (O_1404,N_9013,N_7903);
nor UO_1405 (O_1405,N_7616,N_9180);
or UO_1406 (O_1406,N_7710,N_8501);
and UO_1407 (O_1407,N_7665,N_8757);
and UO_1408 (O_1408,N_9174,N_8673);
or UO_1409 (O_1409,N_9310,N_7691);
xnor UO_1410 (O_1410,N_8291,N_8232);
nor UO_1411 (O_1411,N_7555,N_9597);
nor UO_1412 (O_1412,N_8041,N_8202);
nand UO_1413 (O_1413,N_9517,N_9969);
nor UO_1414 (O_1414,N_9453,N_7765);
or UO_1415 (O_1415,N_8588,N_9626);
or UO_1416 (O_1416,N_7818,N_7898);
nand UO_1417 (O_1417,N_7827,N_9789);
or UO_1418 (O_1418,N_9866,N_8239);
nor UO_1419 (O_1419,N_7703,N_9704);
nand UO_1420 (O_1420,N_9172,N_7600);
nand UO_1421 (O_1421,N_9210,N_8976);
or UO_1422 (O_1422,N_9971,N_7848);
and UO_1423 (O_1423,N_9804,N_8839);
or UO_1424 (O_1424,N_9486,N_9744);
or UO_1425 (O_1425,N_8256,N_9665);
and UO_1426 (O_1426,N_9623,N_9414);
nand UO_1427 (O_1427,N_7644,N_8319);
and UO_1428 (O_1428,N_7927,N_9928);
or UO_1429 (O_1429,N_9060,N_8298);
nor UO_1430 (O_1430,N_9779,N_7969);
nand UO_1431 (O_1431,N_8358,N_8385);
or UO_1432 (O_1432,N_8071,N_7931);
or UO_1433 (O_1433,N_9636,N_7626);
nand UO_1434 (O_1434,N_9953,N_7838);
or UO_1435 (O_1435,N_8282,N_9822);
nor UO_1436 (O_1436,N_8291,N_8498);
or UO_1437 (O_1437,N_8104,N_7570);
and UO_1438 (O_1438,N_9161,N_7987);
or UO_1439 (O_1439,N_9392,N_8587);
or UO_1440 (O_1440,N_9574,N_7956);
nor UO_1441 (O_1441,N_9107,N_7968);
or UO_1442 (O_1442,N_7808,N_8203);
nand UO_1443 (O_1443,N_8841,N_7500);
nand UO_1444 (O_1444,N_8191,N_7655);
nor UO_1445 (O_1445,N_8946,N_8776);
nor UO_1446 (O_1446,N_9495,N_7720);
nand UO_1447 (O_1447,N_8533,N_8607);
nand UO_1448 (O_1448,N_7521,N_9783);
nor UO_1449 (O_1449,N_7916,N_8921);
nand UO_1450 (O_1450,N_8500,N_9812);
nand UO_1451 (O_1451,N_9395,N_9262);
nor UO_1452 (O_1452,N_8571,N_8961);
or UO_1453 (O_1453,N_8540,N_9126);
nor UO_1454 (O_1454,N_8276,N_7568);
or UO_1455 (O_1455,N_9983,N_8589);
or UO_1456 (O_1456,N_7774,N_8778);
nor UO_1457 (O_1457,N_8322,N_9412);
nor UO_1458 (O_1458,N_7729,N_9211);
nand UO_1459 (O_1459,N_7545,N_9157);
nand UO_1460 (O_1460,N_8540,N_9720);
nand UO_1461 (O_1461,N_7892,N_8333);
nand UO_1462 (O_1462,N_9141,N_9069);
or UO_1463 (O_1463,N_7673,N_8793);
or UO_1464 (O_1464,N_7570,N_7664);
and UO_1465 (O_1465,N_7825,N_9275);
nor UO_1466 (O_1466,N_9136,N_7998);
or UO_1467 (O_1467,N_7809,N_7982);
nand UO_1468 (O_1468,N_7936,N_8474);
nand UO_1469 (O_1469,N_8195,N_8870);
nand UO_1470 (O_1470,N_8192,N_9290);
nand UO_1471 (O_1471,N_9585,N_9291);
nand UO_1472 (O_1472,N_9284,N_8847);
nor UO_1473 (O_1473,N_8114,N_8163);
nor UO_1474 (O_1474,N_7919,N_9881);
or UO_1475 (O_1475,N_9522,N_8555);
nand UO_1476 (O_1476,N_9441,N_8877);
nor UO_1477 (O_1477,N_9275,N_9974);
nand UO_1478 (O_1478,N_9645,N_9099);
nand UO_1479 (O_1479,N_8323,N_7582);
or UO_1480 (O_1480,N_7809,N_7674);
or UO_1481 (O_1481,N_8839,N_9346);
or UO_1482 (O_1482,N_9745,N_8217);
nand UO_1483 (O_1483,N_9150,N_8509);
and UO_1484 (O_1484,N_9001,N_8349);
and UO_1485 (O_1485,N_9725,N_7760);
nand UO_1486 (O_1486,N_8000,N_8264);
and UO_1487 (O_1487,N_9805,N_9894);
xor UO_1488 (O_1488,N_9097,N_9359);
nor UO_1489 (O_1489,N_7913,N_8014);
nor UO_1490 (O_1490,N_9946,N_8266);
and UO_1491 (O_1491,N_8955,N_9512);
nand UO_1492 (O_1492,N_8887,N_7590);
and UO_1493 (O_1493,N_7506,N_9951);
nor UO_1494 (O_1494,N_9435,N_7544);
nand UO_1495 (O_1495,N_8628,N_9716);
and UO_1496 (O_1496,N_8681,N_9447);
or UO_1497 (O_1497,N_9083,N_9397);
or UO_1498 (O_1498,N_7836,N_7977);
nor UO_1499 (O_1499,N_9946,N_8016);
endmodule