module basic_2500_25000_3000_5_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1776,In_1771);
nor U1 (N_1,In_2166,In_124);
nor U2 (N_2,In_1149,In_1673);
nor U3 (N_3,In_943,In_1219);
or U4 (N_4,In_1848,In_1971);
nor U5 (N_5,In_940,In_508);
nand U6 (N_6,In_889,In_853);
or U7 (N_7,In_66,In_1871);
nor U8 (N_8,In_1765,In_2405);
and U9 (N_9,In_161,In_1066);
nor U10 (N_10,In_1596,In_2499);
nand U11 (N_11,In_752,In_974);
nand U12 (N_12,In_152,In_1387);
and U13 (N_13,In_166,In_181);
nor U14 (N_14,In_2056,In_798);
or U15 (N_15,In_302,In_680);
nor U16 (N_16,In_311,In_756);
and U17 (N_17,In_592,In_670);
nand U18 (N_18,In_268,In_1227);
nor U19 (N_19,In_2101,In_2346);
or U20 (N_20,In_2171,In_1630);
or U21 (N_21,In_1130,In_704);
nand U22 (N_22,In_1942,In_1054);
nor U23 (N_23,In_1716,In_952);
and U24 (N_24,In_2277,In_1518);
and U25 (N_25,In_532,In_2469);
or U26 (N_26,In_1124,In_621);
and U27 (N_27,In_1178,In_1413);
xnor U28 (N_28,In_771,In_1141);
and U29 (N_29,In_2282,In_1660);
or U30 (N_30,In_1175,In_1183);
nand U31 (N_31,In_1273,In_226);
or U32 (N_32,In_2480,In_1969);
nand U33 (N_33,In_369,In_1921);
or U34 (N_34,In_1010,In_1880);
and U35 (N_35,In_1912,In_1424);
or U36 (N_36,In_1843,In_30);
nor U37 (N_37,In_103,In_1333);
xnor U38 (N_38,In_1624,In_923);
and U39 (N_39,In_1829,In_1464);
or U40 (N_40,In_1091,In_389);
nor U41 (N_41,In_1080,In_1634);
nor U42 (N_42,In_1063,In_368);
or U43 (N_43,In_998,In_1537);
xor U44 (N_44,In_214,In_1523);
nand U45 (N_45,In_457,In_2017);
nand U46 (N_46,In_1000,In_1437);
nand U47 (N_47,In_238,In_295);
or U48 (N_48,In_2260,In_2200);
and U49 (N_49,In_785,In_1929);
and U50 (N_50,In_2250,In_1743);
nor U51 (N_51,In_783,In_292);
xor U52 (N_52,In_394,In_1348);
nor U53 (N_53,In_1043,In_1497);
nand U54 (N_54,In_672,In_1128);
nor U55 (N_55,In_958,In_1650);
and U56 (N_56,In_1255,In_40);
nor U57 (N_57,In_2394,In_1571);
nor U58 (N_58,In_1306,In_2124);
nor U59 (N_59,In_1747,In_936);
nand U60 (N_60,In_945,In_135);
or U61 (N_61,In_1269,In_1234);
nor U62 (N_62,In_875,In_1590);
or U63 (N_63,In_1990,In_1356);
nor U64 (N_64,In_1636,In_1807);
or U65 (N_65,In_240,In_1996);
xnor U66 (N_66,In_458,In_819);
and U67 (N_67,In_2107,In_1198);
nor U68 (N_68,In_797,In_754);
nand U69 (N_69,In_1613,In_1231);
xnor U70 (N_70,In_938,In_1465);
and U71 (N_71,In_2284,In_1194);
or U72 (N_72,In_779,In_435);
nor U73 (N_73,In_1642,In_1296);
nand U74 (N_74,In_2345,In_398);
and U75 (N_75,In_1378,In_362);
nor U76 (N_76,In_2073,In_1079);
nand U77 (N_77,In_542,In_858);
or U78 (N_78,In_2093,In_1385);
xnor U79 (N_79,In_782,In_1480);
or U80 (N_80,In_1827,In_980);
nor U81 (N_81,In_984,In_1867);
or U82 (N_82,In_873,In_1013);
and U83 (N_83,In_2266,In_207);
nor U84 (N_84,In_477,In_1312);
xnor U85 (N_85,In_1617,In_2371);
xor U86 (N_86,In_106,In_1386);
nor U87 (N_87,In_1560,In_916);
nand U88 (N_88,In_999,In_44);
nand U89 (N_89,In_1671,In_19);
nand U90 (N_90,In_2011,In_2026);
or U91 (N_91,In_628,In_1648);
nand U92 (N_92,In_48,In_461);
or U93 (N_93,In_299,In_2215);
and U94 (N_94,In_1811,In_267);
xnor U95 (N_95,In_1467,In_1979);
and U96 (N_96,In_1210,In_598);
nor U97 (N_97,In_2397,In_1574);
nor U98 (N_98,In_1801,In_23);
or U99 (N_99,In_582,In_1429);
nand U100 (N_100,In_63,In_1318);
nand U101 (N_101,In_313,In_57);
and U102 (N_102,In_212,In_352);
and U103 (N_103,In_511,In_564);
and U104 (N_104,In_1045,In_1721);
and U105 (N_105,In_820,In_1770);
and U106 (N_106,In_1111,In_538);
nand U107 (N_107,In_550,In_1007);
and U108 (N_108,In_2417,In_1478);
and U109 (N_109,In_288,In_1939);
or U110 (N_110,In_440,In_2204);
xor U111 (N_111,In_1311,In_2079);
nor U112 (N_112,In_1557,In_1153);
and U113 (N_113,In_1719,In_417);
and U114 (N_114,In_1620,In_1099);
or U115 (N_115,In_1932,In_846);
nand U116 (N_116,In_2339,In_713);
or U117 (N_117,In_922,In_514);
and U118 (N_118,In_344,In_963);
nor U119 (N_119,In_1443,In_824);
nand U120 (N_120,In_823,In_371);
or U121 (N_121,In_2237,In_775);
nor U122 (N_122,In_2433,In_1872);
nand U123 (N_123,In_1678,In_685);
nor U124 (N_124,In_1439,In_2210);
nor U125 (N_125,In_2172,In_1191);
or U126 (N_126,In_147,In_423);
nor U127 (N_127,In_2470,In_2475);
or U128 (N_128,In_1949,In_338);
and U129 (N_129,In_992,In_2140);
nor U130 (N_130,In_2238,In_2476);
nand U131 (N_131,In_2029,In_50);
xor U132 (N_132,In_1181,In_2445);
nand U133 (N_133,In_1305,In_2316);
or U134 (N_134,In_1694,In_2141);
or U135 (N_135,In_1883,In_16);
nand U136 (N_136,In_1758,In_1082);
nand U137 (N_137,In_911,In_574);
nor U138 (N_138,In_1566,In_125);
xnor U139 (N_139,In_1899,In_2412);
and U140 (N_140,In_1316,In_1391);
and U141 (N_141,In_1024,In_1358);
and U142 (N_142,In_1221,In_1334);
xor U143 (N_143,In_1328,In_657);
nor U144 (N_144,In_2183,In_4);
nand U145 (N_145,In_773,In_2488);
or U146 (N_146,In_615,In_24);
and U147 (N_147,In_364,In_1607);
nand U148 (N_148,In_460,In_2311);
or U149 (N_149,In_1274,In_6);
nand U150 (N_150,In_2449,In_312);
nor U151 (N_151,In_223,In_193);
and U152 (N_152,In_1362,In_690);
xnor U153 (N_153,In_1120,In_2437);
nor U154 (N_154,In_780,In_2203);
or U155 (N_155,In_1220,In_1762);
and U156 (N_156,In_1185,In_720);
and U157 (N_157,In_410,In_1197);
nor U158 (N_158,In_202,In_1174);
nor U159 (N_159,In_251,In_235);
nor U160 (N_160,In_8,In_1856);
nor U161 (N_161,In_1886,In_2032);
nand U162 (N_162,In_2464,In_1299);
and U163 (N_163,In_1987,In_2111);
or U164 (N_164,In_1044,In_1182);
nor U165 (N_165,In_1235,In_1171);
or U166 (N_166,In_336,In_1554);
or U167 (N_167,In_932,In_744);
nand U168 (N_168,In_2130,In_2361);
and U169 (N_169,In_1798,In_904);
nand U170 (N_170,In_492,In_1692);
nor U171 (N_171,In_1831,In_272);
nand U172 (N_172,In_178,In_2465);
or U173 (N_173,In_224,In_1240);
or U174 (N_174,In_218,In_1857);
nor U175 (N_175,In_1340,In_1610);
nand U176 (N_176,In_2393,In_957);
and U177 (N_177,In_1879,In_1331);
or U178 (N_178,In_1276,In_1307);
nor U179 (N_179,In_1631,In_1520);
nand U180 (N_180,In_883,In_2078);
nor U181 (N_181,In_590,In_979);
nand U182 (N_182,In_2187,In_1127);
xor U183 (N_183,In_1202,In_1972);
nand U184 (N_184,In_290,In_600);
or U185 (N_185,In_427,In_328);
and U186 (N_186,In_80,In_99);
nor U187 (N_187,In_1001,In_517);
nand U188 (N_188,In_201,In_120);
nand U189 (N_189,In_1584,In_79);
nor U190 (N_190,In_342,In_1917);
and U191 (N_191,In_2424,In_521);
xor U192 (N_192,In_206,In_835);
nor U193 (N_193,In_1053,In_512);
or U194 (N_194,In_1753,In_839);
nand U195 (N_195,In_1304,In_885);
and U196 (N_196,In_2342,In_2427);
or U197 (N_197,In_795,In_1058);
nor U198 (N_198,In_1789,In_1196);
or U199 (N_199,In_2122,In_35);
nand U200 (N_200,In_1676,In_1579);
and U201 (N_201,In_1261,In_494);
or U202 (N_202,In_1794,In_1346);
nor U203 (N_203,In_1492,In_62);
nand U204 (N_204,In_1687,In_169);
or U205 (N_205,In_122,In_863);
and U206 (N_206,In_675,In_2217);
and U207 (N_207,In_231,In_894);
or U208 (N_208,In_2106,In_154);
and U209 (N_209,In_1207,In_973);
nand U210 (N_210,In_1160,In_2149);
nand U211 (N_211,In_2420,In_2483);
and U212 (N_212,In_324,In_21);
nand U213 (N_213,In_809,In_1322);
nor U214 (N_214,In_1420,In_1495);
and U215 (N_215,In_1992,In_2223);
or U216 (N_216,In_1513,In_1368);
nor U217 (N_217,In_1956,In_1578);
nand U218 (N_218,In_1375,In_996);
or U219 (N_219,In_699,In_1587);
and U220 (N_220,In_1682,In_480);
and U221 (N_221,In_919,In_1618);
xor U222 (N_222,In_2207,In_1115);
nor U223 (N_223,In_2466,In_840);
and U224 (N_224,In_56,In_363);
or U225 (N_225,In_374,In_1760);
nor U226 (N_226,In_482,In_2481);
nor U227 (N_227,In_306,In_1050);
nand U228 (N_228,In_642,In_2010);
and U229 (N_229,In_1994,In_102);
nor U230 (N_230,In_2389,In_614);
and U231 (N_231,In_1840,In_2060);
nand U232 (N_232,In_553,In_1301);
nand U233 (N_233,In_948,In_523);
nand U234 (N_234,In_2162,In_1874);
and U235 (N_235,In_49,In_1715);
nand U236 (N_236,In_1597,In_1940);
and U237 (N_237,In_1282,In_715);
or U238 (N_238,In_537,In_1906);
and U239 (N_239,In_1549,In_351);
nand U240 (N_240,In_2391,In_1611);
and U241 (N_241,In_1498,In_2357);
and U242 (N_242,In_705,In_2461);
xnor U243 (N_243,In_1473,In_585);
and U244 (N_244,In_641,In_396);
and U245 (N_245,In_1270,In_865);
or U246 (N_246,In_2062,In_1695);
and U247 (N_247,In_887,In_740);
nor U248 (N_248,In_1034,In_730);
nand U249 (N_249,In_1913,In_384);
nand U250 (N_250,In_1842,In_1486);
or U251 (N_251,In_880,In_107);
nand U252 (N_252,In_725,In_991);
and U253 (N_253,In_2247,In_695);
and U254 (N_254,In_465,In_1825);
and U255 (N_255,In_228,In_1187);
and U256 (N_256,In_997,In_2471);
or U257 (N_257,In_1657,In_1895);
nor U258 (N_258,In_82,In_700);
nand U259 (N_259,In_276,In_2377);
and U260 (N_260,In_1190,In_770);
or U261 (N_261,In_866,In_800);
and U262 (N_262,In_1793,In_518);
and U263 (N_263,In_366,In_1105);
nand U264 (N_264,In_1173,In_1014);
xor U265 (N_265,In_620,In_2186);
and U266 (N_266,In_320,In_2309);
and U267 (N_267,In_0,In_441);
nand U268 (N_268,In_1780,In_581);
nor U269 (N_269,In_2194,In_1705);
nor U270 (N_270,In_1315,In_10);
and U271 (N_271,In_330,In_2047);
xnor U272 (N_272,In_192,In_1514);
nor U273 (N_273,In_1752,In_2334);
nor U274 (N_274,In_386,In_2096);
nor U275 (N_275,In_1628,In_1217);
xor U276 (N_276,In_815,In_1446);
and U277 (N_277,In_506,In_1106);
nand U278 (N_278,In_1057,In_1891);
xor U279 (N_279,In_1922,In_1774);
and U280 (N_280,In_2281,In_660);
nor U281 (N_281,In_2315,In_26);
or U282 (N_282,In_1077,In_456);
or U283 (N_283,In_1935,In_1188);
nor U284 (N_284,In_2262,In_2151);
nand U285 (N_285,In_1452,In_1909);
nor U286 (N_286,In_2132,In_432);
or U287 (N_287,In_1409,In_1865);
nand U288 (N_288,In_25,In_222);
xnor U289 (N_289,In_2232,In_2103);
and U290 (N_290,In_1675,In_1545);
nand U291 (N_291,In_297,In_1086);
nand U292 (N_292,In_2416,In_2409);
or U293 (N_293,In_867,In_339);
or U294 (N_294,In_1728,In_2369);
and U295 (N_295,In_2014,In_210);
nand U296 (N_296,In_227,In_2312);
nand U297 (N_297,In_1302,In_803);
nand U298 (N_298,In_2155,In_1820);
nand U299 (N_299,In_2045,In_1816);
or U300 (N_300,In_1565,In_179);
and U301 (N_301,In_53,In_332);
nor U302 (N_302,In_486,In_59);
and U303 (N_303,In_12,In_647);
nor U304 (N_304,In_1354,In_1928);
xnor U305 (N_305,In_28,In_544);
and U306 (N_306,In_665,In_2372);
nand U307 (N_307,In_1543,In_94);
or U308 (N_308,In_2478,In_1468);
and U309 (N_309,In_1941,In_879);
nor U310 (N_310,In_649,In_2362);
nand U311 (N_311,In_644,In_2125);
nor U312 (N_312,In_1748,In_2450);
nor U313 (N_313,In_2325,In_503);
nor U314 (N_314,In_2374,In_850);
nor U315 (N_315,In_2330,In_408);
nor U316 (N_316,In_326,In_1457);
xnor U317 (N_317,In_255,In_2228);
nand U318 (N_318,In_2294,In_886);
or U319 (N_319,In_2307,In_2002);
nor U320 (N_320,In_1140,In_289);
nor U321 (N_321,In_1833,In_2340);
xnor U322 (N_322,In_2050,In_2072);
nand U323 (N_323,In_85,In_1726);
nor U324 (N_324,In_1658,In_1643);
xnor U325 (N_325,In_913,In_668);
nor U326 (N_326,In_110,In_1600);
xor U327 (N_327,In_1944,In_1325);
and U328 (N_328,In_2066,In_909);
nand U329 (N_329,In_2319,In_1417);
nor U330 (N_330,In_1094,In_309);
nor U331 (N_331,In_1622,In_1858);
and U332 (N_332,In_575,In_1766);
xnor U333 (N_333,In_1977,In_2129);
or U334 (N_334,In_2058,In_1162);
nor U335 (N_335,In_2218,In_1646);
nand U336 (N_336,In_187,In_205);
and U337 (N_337,In_490,In_1357);
and U338 (N_338,In_2328,In_462);
and U339 (N_339,In_505,In_1509);
nor U340 (N_340,In_1009,In_2279);
and U341 (N_341,In_1625,In_1238);
and U342 (N_342,In_1364,In_1718);
or U343 (N_343,In_1538,In_116);
xor U344 (N_344,In_749,In_287);
nand U345 (N_345,In_1277,In_925);
nand U346 (N_346,In_1293,In_2095);
nand U347 (N_347,In_694,In_176);
or U348 (N_348,In_758,In_1741);
nand U349 (N_349,In_1143,In_111);
nand U350 (N_350,In_1,In_407);
or U351 (N_351,In_681,In_870);
or U352 (N_352,In_2343,In_421);
nand U353 (N_353,In_18,In_527);
or U354 (N_354,In_682,In_2081);
xor U355 (N_355,In_191,In_1258);
nor U356 (N_356,In_1614,In_1338);
nand U357 (N_357,In_2191,In_2318);
nand U358 (N_358,In_2375,In_2080);
nor U359 (N_359,In_2364,In_818);
nor U360 (N_360,In_2188,In_360);
xor U361 (N_361,In_653,In_1550);
xnor U362 (N_362,In_1696,In_722);
nor U363 (N_363,In_2451,In_579);
nor U364 (N_364,In_661,In_502);
nand U365 (N_365,In_1900,In_807);
nand U366 (N_366,In_1397,In_1796);
or U367 (N_367,In_1121,In_2051);
and U368 (N_368,In_2495,In_1915);
or U369 (N_369,In_2181,In_1846);
nor U370 (N_370,In_2278,In_2182);
nand U371 (N_371,In_1479,In_2335);
xor U372 (N_372,In_2033,In_2244);
xor U373 (N_373,In_1005,In_1575);
nor U374 (N_374,In_1564,In_1224);
and U375 (N_375,In_1243,In_357);
and U376 (N_376,In_1205,In_890);
nor U377 (N_377,In_1866,In_1936);
nor U378 (N_378,In_2021,In_985);
or U379 (N_379,In_1109,In_2486);
or U380 (N_380,In_425,In_42);
and U381 (N_381,In_882,In_1072);
nand U382 (N_382,In_2264,In_844);
nand U383 (N_383,In_1402,In_738);
nand U384 (N_384,In_11,In_584);
nor U385 (N_385,In_1421,In_1419);
xnor U386 (N_386,In_2439,In_1155);
xor U387 (N_387,In_356,In_1161);
or U388 (N_388,In_841,In_591);
and U389 (N_389,In_1916,In_1159);
or U390 (N_390,In_1700,In_655);
and U391 (N_391,In_859,In_721);
and U392 (N_392,In_716,In_2314);
or U393 (N_393,In_118,In_1179);
xnor U394 (N_394,In_2387,In_1740);
nor U395 (N_395,In_519,In_404);
and U396 (N_396,In_257,In_1176);
nor U397 (N_397,In_1986,In_965);
and U398 (N_398,In_445,In_1195);
xor U399 (N_399,In_931,In_1237);
or U400 (N_400,In_1701,In_2399);
nor U401 (N_401,In_378,In_434);
xor U402 (N_402,In_1474,In_220);
xnor U403 (N_403,In_1319,In_133);
nor U404 (N_404,In_856,In_1389);
nand U405 (N_405,In_552,In_2097);
nand U406 (N_406,In_708,In_2295);
nand U407 (N_407,In_1686,In_2378);
nand U408 (N_408,In_1963,In_2268);
xnor U409 (N_409,In_254,In_1755);
nor U410 (N_410,In_1403,In_516);
nand U411 (N_411,In_75,In_1426);
or U412 (N_412,In_373,In_1395);
and U413 (N_413,In_849,In_1707);
or U414 (N_414,In_1681,In_693);
nand U415 (N_415,In_1133,In_243);
nor U416 (N_416,In_724,In_2185);
xor U417 (N_417,In_1084,In_2257);
and U418 (N_418,In_597,In_2429);
or U419 (N_419,In_1892,In_27);
or U420 (N_420,In_1021,In_1369);
xnor U421 (N_421,In_1868,In_1887);
nor U422 (N_422,In_1062,In_258);
nand U423 (N_423,In_651,In_1703);
xnor U424 (N_424,In_1108,In_1323);
and U425 (N_425,In_712,In_489);
and U426 (N_426,In_1924,In_1947);
or U427 (N_427,In_570,In_1134);
or U428 (N_428,In_2484,In_1422);
and U429 (N_429,In_2211,In_1951);
nand U430 (N_430,In_1392,In_2089);
or U431 (N_431,In_2253,In_1309);
nand U432 (N_432,In_1608,In_1107);
nand U433 (N_433,In_1745,In_2161);
nand U434 (N_434,In_84,In_656);
nor U435 (N_435,In_1327,In_761);
and U436 (N_436,In_500,In_189);
nor U437 (N_437,In_1595,In_1905);
nand U438 (N_438,In_1727,In_183);
nand U439 (N_439,In_1247,In_2255);
nand U440 (N_440,In_1476,In_2177);
nand U441 (N_441,In_1408,In_1961);
or U442 (N_442,In_1893,In_1085);
nor U443 (N_443,In_203,In_676);
and U444 (N_444,In_1785,In_348);
or U445 (N_445,In_2440,In_392);
nand U446 (N_446,In_2157,In_1157);
nor U447 (N_447,In_1339,In_2249);
nor U448 (N_448,In_960,In_1100);
and U449 (N_449,In_1551,In_2298);
and U450 (N_450,In_158,In_2);
nand U451 (N_451,In_264,In_170);
xnor U452 (N_452,In_1945,In_580);
or U453 (N_453,In_784,In_616);
or U454 (N_454,In_2441,In_688);
or U455 (N_455,In_2110,In_499);
nor U456 (N_456,In_2115,In_2027);
or U457 (N_457,In_164,In_270);
nand U458 (N_458,In_2384,In_1363);
nor U459 (N_459,In_1493,In_266);
and U460 (N_460,In_1999,In_1029);
and U461 (N_461,In_2327,In_2102);
nand U462 (N_462,In_1097,In_2438);
nand U463 (N_463,In_1954,In_2356);
nand U464 (N_464,In_1666,In_347);
nand U465 (N_465,In_317,In_2165);
nand U466 (N_466,In_148,In_2082);
nand U467 (N_467,In_2270,In_1505);
and U468 (N_468,In_130,In_1022);
and U469 (N_469,In_117,In_2426);
and U470 (N_470,In_1683,In_265);
nand U471 (N_471,In_640,In_2174);
nor U472 (N_472,In_399,In_1329);
or U473 (N_473,In_833,In_159);
nor U474 (N_474,In_1225,In_1399);
nor U475 (N_475,In_150,In_860);
nand U476 (N_476,In_727,In_1964);
nor U477 (N_477,In_194,In_1768);
nor U478 (N_478,In_2313,In_2001);
or U479 (N_479,In_1092,In_2020);
and U480 (N_480,In_403,In_1754);
nor U481 (N_481,In_830,In_1923);
nand U482 (N_482,In_1216,In_349);
nand U483 (N_483,In_2192,In_2071);
xor U484 (N_484,In_1837,In_1347);
nor U485 (N_485,In_1882,In_1616);
nand U486 (N_486,In_821,In_2169);
nand U487 (N_487,In_1263,In_1985);
and U488 (N_488,In_781,In_464);
and U489 (N_489,In_2112,In_1090);
nor U490 (N_490,In_2408,In_622);
or U491 (N_491,In_817,In_556);
xnor U492 (N_492,In_215,In_2022);
nand U493 (N_493,In_1405,In_2413);
and U494 (N_494,In_453,In_1959);
and U495 (N_495,In_1980,In_496);
nor U496 (N_496,In_710,In_1812);
nand U497 (N_497,In_2018,In_1907);
and U498 (N_498,In_734,In_1172);
and U499 (N_499,In_232,In_1734);
nand U500 (N_500,In_455,In_1169);
or U501 (N_501,In_2322,In_1152);
and U502 (N_502,In_2213,In_137);
xor U503 (N_503,In_1724,In_1461);
xor U504 (N_504,In_627,In_2139);
nor U505 (N_505,In_81,In_2428);
xor U506 (N_506,In_1449,In_1808);
nand U507 (N_507,In_1170,In_2292);
nor U508 (N_508,In_229,In_1314);
or U509 (N_509,In_1621,In_1275);
or U510 (N_510,In_2241,In_1502);
and U511 (N_511,In_1067,In_1761);
nand U512 (N_512,In_47,In_1731);
nor U513 (N_513,In_51,In_1265);
or U514 (N_514,In_1836,In_759);
or U515 (N_515,In_1663,In_149);
xor U516 (N_516,In_563,In_1526);
or U517 (N_517,In_1114,In_1573);
and U518 (N_518,In_2134,In_1647);
or U519 (N_519,In_1455,In_36);
or U520 (N_520,In_696,In_969);
and U521 (N_521,In_329,In_1697);
or U522 (N_522,In_95,In_1732);
or U523 (N_523,In_38,In_2236);
or U524 (N_524,In_340,In_1644);
xnor U525 (N_525,In_126,In_2396);
or U526 (N_526,In_100,In_757);
or U527 (N_527,In_2164,In_2076);
nor U528 (N_528,In_567,In_1040);
nor U529 (N_529,In_395,In_1896);
or U530 (N_530,In_139,In_239);
nand U531 (N_531,In_1390,In_1425);
nor U532 (N_532,In_2453,In_249);
or U533 (N_533,In_792,In_843);
and U534 (N_534,In_60,In_1218);
or U535 (N_535,In_1163,In_1568);
nand U536 (N_536,In_528,In_1450);
and U537 (N_537,In_2333,In_1410);
or U538 (N_538,In_659,In_1531);
and U539 (N_539,In_1324,In_1563);
and U540 (N_540,In_296,In_918);
and U541 (N_541,In_128,In_1885);
or U542 (N_542,In_1569,In_1360);
and U543 (N_543,In_2015,In_1239);
xnor U544 (N_544,In_2289,In_2075);
nor U545 (N_545,In_679,In_990);
or U546 (N_546,In_701,In_151);
or U547 (N_547,In_1295,In_986);
and U548 (N_548,In_479,In_1469);
xnor U549 (N_549,In_664,In_476);
or U550 (N_550,In_1065,In_1974);
nor U551 (N_551,In_7,In_2276);
xor U552 (N_552,In_469,In_525);
nand U553 (N_553,In_766,In_852);
nand U554 (N_554,In_613,In_707);
xor U555 (N_555,In_337,In_1581);
nand U556 (N_556,In_1499,In_1943);
or U557 (N_557,In_976,In_2366);
or U558 (N_558,In_806,In_2332);
or U559 (N_559,In_273,In_1637);
nand U560 (N_560,In_2098,In_321);
nor U561 (N_561,In_671,In_1448);
and U562 (N_562,In_32,In_731);
nor U563 (N_563,In_692,In_1477);
nand U564 (N_564,In_2109,In_1393);
or U565 (N_565,In_1381,In_77);
xnor U566 (N_566,In_1997,In_971);
or U567 (N_567,In_1838,In_1792);
or U568 (N_568,In_1791,In_216);
and U569 (N_569,In_1784,In_1343);
and U570 (N_570,In_1805,In_1102);
nand U571 (N_571,In_1285,In_431);
xor U572 (N_572,In_293,In_861);
nand U573 (N_573,In_132,In_1652);
and U574 (N_574,In_109,In_1048);
nand U575 (N_575,In_1436,In_778);
or U576 (N_576,In_2007,In_977);
nand U577 (N_577,In_359,In_2263);
and U578 (N_578,In_1733,In_1713);
nand U579 (N_579,In_2242,In_654);
xnor U580 (N_580,In_1462,In_831);
and U581 (N_581,In_2304,In_1998);
nand U582 (N_582,In_1670,In_375);
or U583 (N_583,In_333,In_586);
nand U584 (N_584,In_691,In_1254);
or U585 (N_585,In_813,In_213);
or U586 (N_586,In_1208,In_2457);
nor U587 (N_587,In_1435,In_2030);
and U588 (N_588,In_1146,In_2305);
or U589 (N_589,In_663,In_1491);
nor U590 (N_590,In_639,In_1246);
nor U591 (N_591,In_1699,In_684);
and U592 (N_592,In_1335,In_1052);
and U593 (N_593,In_558,In_810);
or U594 (N_594,In_1104,In_1504);
xnor U595 (N_595,In_902,In_1407);
and U596 (N_596,In_2400,In_802);
and U597 (N_597,In_2025,In_1380);
nor U598 (N_598,In_2184,In_2430);
nand U599 (N_599,In_2040,In_1788);
or U600 (N_600,In_534,In_531);
or U601 (N_601,In_1326,In_1638);
nor U602 (N_602,In_1918,In_2347);
xnor U603 (N_603,In_1228,In_2105);
or U604 (N_604,In_1962,In_2442);
nand U605 (N_605,In_769,In_2317);
or U606 (N_606,In_1166,In_1136);
nor U607 (N_607,In_673,In_959);
and U608 (N_608,In_1781,In_382);
nand U609 (N_609,In_463,In_2320);
nand U610 (N_610,In_796,In_930);
or U611 (N_611,In_1129,In_334);
xnor U612 (N_612,In_1096,In_454);
and U613 (N_613,In_872,In_411);
or U614 (N_614,In_1308,In_1830);
nand U615 (N_615,In_1189,In_1589);
xor U616 (N_616,In_367,In_529);
or U617 (N_617,In_1125,In_1488);
nor U618 (N_618,In_827,In_593);
or U619 (N_619,In_729,In_987);
and U620 (N_620,In_1763,In_197);
or U621 (N_621,In_127,In_1976);
nor U622 (N_622,In_1680,In_577);
nand U623 (N_623,In_1981,In_1633);
or U624 (N_624,In_101,In_1957);
xnor U625 (N_625,In_252,In_1167);
or U626 (N_626,In_2422,In_646);
and U627 (N_627,In_1342,In_439);
nand U628 (N_628,In_1645,In_915);
or U629 (N_629,In_1931,In_964);
nor U630 (N_630,In_171,In_275);
nand U631 (N_631,In_789,In_2458);
or U632 (N_632,In_2248,In_805);
and U633 (N_633,In_199,In_1475);
and U634 (N_634,In_241,In_74);
xnor U635 (N_635,In_1592,In_1729);
xnor U636 (N_636,In_1859,In_1668);
nand U637 (N_637,In_626,In_388);
nand U638 (N_638,In_1144,In_2064);
or U639 (N_639,In_914,In_857);
nand U640 (N_640,In_1902,In_58);
and U641 (N_641,In_1026,In_1786);
xor U642 (N_642,In_1209,In_1904);
xor U643 (N_643,In_1712,In_1177);
or U644 (N_644,In_1165,In_745);
and U645 (N_645,In_2252,In_1113);
nand U646 (N_646,In_274,In_1484);
and U647 (N_647,In_1524,In_1151);
nand U648 (N_648,In_2494,In_1601);
nor U649 (N_649,In_2159,In_2273);
nor U650 (N_650,In_808,In_1352);
nand U651 (N_651,In_2028,In_1490);
and U652 (N_652,In_1222,In_1003);
xnor U653 (N_653,In_2120,In_2150);
nand U654 (N_654,In_2083,In_1599);
and U655 (N_655,In_131,In_1418);
nand U656 (N_656,In_413,In_895);
or U657 (N_657,In_669,In_269);
nor U658 (N_658,In_41,In_475);
or U659 (N_659,In_698,In_1186);
and U660 (N_660,In_2395,In_1655);
and U661 (N_661,In_2013,In_1824);
nand U662 (N_662,In_2158,In_400);
and U663 (N_663,In_1374,In_1881);
nand U664 (N_664,In_157,In_370);
and U665 (N_665,In_2216,In_2302);
and U666 (N_666,In_554,In_608);
or U667 (N_667,In_636,In_1783);
nor U668 (N_668,In_983,In_2344);
xor U669 (N_669,In_245,In_1877);
nand U670 (N_670,In_2114,In_474);
nand U671 (N_671,In_751,In_1500);
xnor U672 (N_672,In_1736,In_719);
nand U673 (N_673,In_2376,In_1023);
nand U674 (N_674,In_278,In_728);
or U675 (N_675,In_2415,In_225);
nor U676 (N_676,In_946,In_1693);
or U677 (N_677,In_603,In_2491);
xor U678 (N_678,In_888,In_1510);
nor U679 (N_679,In_1145,In_2175);
nand U680 (N_680,In_1822,In_1242);
or U681 (N_681,In_548,In_426);
and U682 (N_682,In_924,In_1561);
and U683 (N_683,In_141,In_1373);
nor U684 (N_684,In_2180,In_1559);
and U685 (N_685,In_1359,In_1441);
or U686 (N_686,In_1995,In_1850);
or U687 (N_687,In_2049,In_259);
and U688 (N_688,In_2406,In_2091);
nor U689 (N_689,In_2163,In_2326);
nor U690 (N_690,In_1416,In_415);
or U691 (N_691,In_1076,In_1456);
nor U692 (N_692,In_2310,In_2303);
nand U693 (N_693,In_804,In_1852);
nand U694 (N_694,In_2154,In_897);
and U695 (N_695,In_767,In_1722);
and U696 (N_696,In_1967,In_1772);
and U697 (N_697,In_559,In_1336);
nand U698 (N_698,In_2354,In_1711);
or U699 (N_699,In_607,In_1290);
nor U700 (N_700,In_755,In_1983);
nand U701 (N_701,In_497,In_1081);
nor U702 (N_702,In_303,In_1394);
nand U703 (N_703,In_1725,In_678);
xor U704 (N_704,In_134,In_735);
nor U705 (N_705,In_436,In_2148);
nand U706 (N_706,In_1083,In_1585);
xor U707 (N_707,In_1201,In_2290);
nor U708 (N_708,In_868,In_551);
nand U709 (N_709,In_71,In_828);
nand U710 (N_710,In_217,In_917);
nor U711 (N_711,In_1496,In_2153);
nand U712 (N_712,In_412,In_448);
nor U713 (N_713,In_928,In_1073);
and U714 (N_714,In_353,In_1317);
or U715 (N_715,In_1677,In_543);
and U716 (N_716,In_1371,In_2275);
xnor U717 (N_717,In_1552,In_711);
and U718 (N_718,In_1423,In_2053);
nor U719 (N_719,In_78,In_633);
and U720 (N_720,In_907,In_2286);
or U721 (N_721,In_1759,In_262);
nor U722 (N_722,In_2337,In_2443);
and U723 (N_723,In_1485,In_2414);
and U724 (N_724,In_136,In_2392);
and U725 (N_725,In_1508,In_2005);
xor U726 (N_726,In_2331,In_718);
or U727 (N_727,In_2460,In_1489);
and U728 (N_728,In_560,In_1016);
xor U729 (N_729,In_1193,In_1006);
nand U730 (N_730,In_331,In_2012);
xor U731 (N_731,In_1773,In_1832);
nor U732 (N_732,In_1011,In_814);
nor U733 (N_733,In_1926,In_2138);
or U734 (N_734,In_829,In_1787);
or U735 (N_735,In_1583,In_934);
and U736 (N_736,In_864,In_1035);
or U737 (N_737,In_995,In_643);
or U738 (N_738,In_847,In_540);
or U739 (N_739,In_1521,In_2136);
nand U740 (N_740,In_2219,In_1609);
nand U741 (N_741,In_507,In_2070);
and U742 (N_742,In_377,In_2057);
nand U743 (N_743,In_935,In_801);
nand U744 (N_744,In_2176,In_1515);
or U745 (N_745,In_774,In_726);
xnor U746 (N_746,In_327,In_2127);
nand U747 (N_747,In_209,In_2035);
xor U748 (N_748,In_1649,In_1087);
nand U749 (N_749,In_450,In_1853);
and U750 (N_750,In_966,In_2487);
nand U751 (N_751,In_1204,In_912);
and U752 (N_752,In_1267,In_5);
nor U753 (N_753,In_1698,In_1903);
xor U754 (N_754,In_2341,In_96);
nand U755 (N_755,In_1993,In_1730);
and U756 (N_756,In_588,In_283);
nor U757 (N_757,In_1570,In_825);
xor U758 (N_758,In_1984,In_2323);
nor U759 (N_759,In_76,In_34);
and U760 (N_760,In_442,In_1028);
or U761 (N_761,In_401,In_390);
xor U762 (N_762,In_1158,In_282);
nand U763 (N_763,In_1946,In_1370);
xnor U764 (N_764,In_1629,In_2447);
or U765 (N_765,In_1401,In_683);
xor U766 (N_766,In_2349,In_2301);
nor U767 (N_767,In_15,In_702);
or U768 (N_768,In_2031,In_1064);
xor U769 (N_769,In_1278,In_1516);
and U770 (N_770,In_162,In_1365);
or U771 (N_771,In_589,In_1025);
or U772 (N_772,In_1555,In_1288);
xor U773 (N_773,In_2363,In_247);
or U774 (N_774,In_1623,In_1139);
and U775 (N_775,In_1869,In_1665);
nor U776 (N_776,In_2368,In_1215);
xnor U777 (N_777,In_1372,In_143);
xor U778 (N_778,In_2365,In_799);
nand U779 (N_779,In_2016,In_1534);
nor U780 (N_780,In_2065,In_155);
nand U781 (N_781,In_1861,In_2477);
or U782 (N_782,In_764,In_2246);
nand U783 (N_783,In_1291,In_2046);
nor U784 (N_784,In_260,In_2462);
nor U785 (N_785,In_70,In_2055);
nand U786 (N_786,In_1015,In_447);
or U787 (N_787,In_1706,In_545);
and U788 (N_788,In_1744,In_746);
nand U789 (N_789,In_68,In_1714);
nor U790 (N_790,In_1672,In_832);
nand U791 (N_791,In_1200,In_811);
nand U792 (N_792,In_1430,In_2459);
xor U793 (N_793,In_1819,In_1870);
nand U794 (N_794,In_1351,In_666);
nand U795 (N_795,In_1937,In_208);
xnor U796 (N_796,In_1349,In_1088);
xor U797 (N_797,In_1810,In_1910);
nand U798 (N_798,In_2173,In_787);
xor U799 (N_799,In_2468,In_658);
and U800 (N_800,In_1075,In_1466);
or U801 (N_801,In_632,In_316);
xor U802 (N_802,In_2054,In_2104);
or U803 (N_803,In_376,In_2170);
and U804 (N_804,In_2145,In_1536);
xor U805 (N_805,In_1547,In_2479);
and U806 (N_806,In_822,In_1864);
nor U807 (N_807,In_1018,In_298);
nand U808 (N_808,In_1232,In_1431);
nand U809 (N_809,In_634,In_2271);
nor U810 (N_810,In_2041,In_1117);
nor U811 (N_811,In_1164,In_2023);
nor U812 (N_812,In_380,In_409);
or U813 (N_813,In_2084,In_576);
and U814 (N_814,In_113,In_468);
nand U815 (N_815,In_419,In_1047);
and U816 (N_816,In_1019,In_2052);
or U817 (N_817,In_2230,In_1150);
nor U818 (N_818,In_104,In_495);
nor U819 (N_819,In_1433,In_1377);
nand U820 (N_820,In_1382,In_2272);
nand U821 (N_821,In_1253,In_105);
and U822 (N_822,In_1262,In_242);
nor U823 (N_823,In_20,In_1619);
nor U824 (N_824,In_1008,In_2493);
or U825 (N_825,In_1519,In_1777);
nand U826 (N_826,In_91,In_186);
and U827 (N_827,In_1717,In_1279);
nand U828 (N_828,In_2259,In_910);
and U829 (N_829,In_355,In_714);
or U830 (N_830,In_1558,In_1684);
and U831 (N_831,In_788,In_1453);
nor U832 (N_832,In_2077,In_1445);
nand U833 (N_833,In_478,In_1546);
nor U834 (N_834,In_650,In_854);
nand U835 (N_835,In_2042,In_504);
nor U836 (N_836,In_772,In_2285);
or U837 (N_837,In_1260,In_2280);
nor U838 (N_838,In_487,In_703);
nand U839 (N_839,In_1782,In_1535);
and U840 (N_840,In_1512,In_1803);
and U841 (N_841,In_1556,In_763);
nand U842 (N_842,In_2118,In_301);
nand U843 (N_843,In_1350,In_509);
xor U844 (N_844,In_112,In_1481);
and U845 (N_845,In_617,In_345);
and U846 (N_846,In_1049,In_623);
nand U847 (N_847,In_851,In_285);
xnor U848 (N_848,In_855,In_165);
xor U849 (N_849,In_687,In_1641);
nor U850 (N_850,In_565,In_204);
nor U851 (N_851,In_140,In_2283);
or U852 (N_852,In_2350,In_1297);
xor U853 (N_853,In_793,In_473);
nor U854 (N_854,In_1103,In_1950);
nor U855 (N_855,In_1203,In_1888);
nor U856 (N_856,In_2160,In_881);
or U857 (N_857,In_978,In_1586);
or U858 (N_858,In_180,In_2231);
nand U859 (N_859,In_901,In_1032);
nand U860 (N_860,In_280,In_1233);
and U861 (N_861,In_184,In_1366);
xor U862 (N_862,In_1427,In_429);
or U863 (N_863,In_1934,In_739);
nand U864 (N_864,In_1635,In_1735);
nand U865 (N_865,In_1991,In_2128);
nor U866 (N_866,In_609,In_156);
or U867 (N_867,In_67,In_604);
and U868 (N_868,In_1933,In_1250);
or U869 (N_869,In_2009,In_2061);
xor U870 (N_870,In_1131,In_845);
and U871 (N_871,In_294,In_899);
and U872 (N_872,In_1415,In_2068);
nand U873 (N_873,In_1398,In_1168);
and U874 (N_874,In_2116,In_1226);
nand U875 (N_875,In_393,In_686);
xnor U876 (N_876,In_524,In_2258);
and U877 (N_877,In_1854,In_2006);
nand U878 (N_878,In_2044,In_1042);
or U879 (N_879,In_1286,In_1135);
and U880 (N_880,In_2472,In_1795);
or U881 (N_881,In_1580,In_1821);
nor U882 (N_882,In_1337,In_1341);
nor U883 (N_883,In_1688,In_2497);
or U884 (N_884,In_2432,In_1321);
and U885 (N_885,In_1664,In_1953);
nand U886 (N_886,In_750,In_1236);
or U887 (N_887,In_536,In_1503);
nand U888 (N_888,In_786,In_2144);
nand U889 (N_889,In_2353,In_1344);
and U890 (N_890,In_286,In_452);
nand U891 (N_891,In_1532,In_596);
or U892 (N_892,In_1494,In_629);
nand U893 (N_893,In_1142,In_1511);
or U894 (N_894,In_1252,In_491);
nand U895 (N_895,In_54,In_291);
or U896 (N_896,In_2297,In_1548);
nor U897 (N_897,In_248,In_1122);
and U898 (N_898,In_2421,In_594);
xnor U899 (N_899,In_522,In_947);
and U900 (N_900,In_1751,In_2206);
or U901 (N_901,In_2074,In_1704);
and U902 (N_902,In_1383,In_325);
and U903 (N_903,In_2099,In_1593);
nand U904 (N_904,In_1463,In_898);
or U905 (N_905,In_1908,In_2467);
and U906 (N_906,In_308,In_619);
nand U907 (N_907,In_571,In_587);
nand U908 (N_908,In_1955,In_405);
xnor U909 (N_909,In_871,In_1444);
and U910 (N_910,In_1482,In_72);
or U911 (N_911,In_195,In_1112);
nor U912 (N_912,In_1442,In_1720);
nand U913 (N_913,In_43,In_1248);
nor U914 (N_914,In_1669,In_1070);
nor U915 (N_915,In_546,In_2269);
nand U916 (N_916,In_595,In_1036);
and U917 (N_917,In_1662,In_2239);
nor U918 (N_918,In_2291,In_1750);
xnor U919 (N_919,In_2212,In_2403);
nand U920 (N_920,In_1860,In_2121);
nand U921 (N_921,In_2198,In_444);
xor U922 (N_922,In_884,In_1598);
nand U923 (N_923,In_2398,In_2224);
and U924 (N_924,In_1839,In_1041);
or U925 (N_925,In_1982,In_1266);
nand U926 (N_926,In_2100,In_1615);
and U927 (N_927,In_13,In_284);
nand U928 (N_928,In_1919,In_848);
and U929 (N_929,In_709,In_1245);
and U930 (N_930,In_1147,In_1211);
nor U931 (N_931,In_1855,In_98);
nor U932 (N_932,In_121,In_196);
nor U933 (N_933,In_956,In_791);
or U934 (N_934,In_1313,In_2452);
nand U935 (N_935,In_1376,In_2431);
and U936 (N_936,In_1890,In_906);
nand U937 (N_937,In_2227,In_219);
and U938 (N_938,In_1320,In_86);
nand U939 (N_939,In_2358,In_2048);
nand U940 (N_940,In_1039,In_2043);
and U941 (N_941,In_424,In_46);
nand U942 (N_942,In_89,In_1004);
nor U943 (N_943,In_547,In_1412);
or U944 (N_944,In_510,In_1823);
nand U945 (N_945,In_662,In_2178);
nand U946 (N_946,In_1797,In_2492);
or U947 (N_947,In_1414,In_17);
nand U948 (N_948,In_485,In_2037);
and U949 (N_949,In_1790,In_611);
nand U950 (N_950,In_138,In_1588);
and U951 (N_951,In_341,In_1817);
or U952 (N_952,In_876,In_549);
nand U953 (N_953,In_573,In_2036);
nor U954 (N_954,In_1017,In_1046);
nand U955 (N_955,In_648,In_318);
or U956 (N_956,In_2090,In_1137);
or U957 (N_957,In_372,In_1757);
nand U958 (N_958,In_1710,In_1257);
nor U959 (N_959,In_271,In_1897);
or U960 (N_960,In_951,In_2063);
or U961 (N_961,In_2038,In_61);
nand U962 (N_962,In_1689,In_1280);
nor U963 (N_963,In_115,In_365);
or U964 (N_964,In_1901,In_1653);
and U965 (N_965,In_1659,In_1685);
and U966 (N_966,In_1702,In_1229);
or U967 (N_967,In_967,In_483);
nor U968 (N_968,In_1212,In_1738);
and U969 (N_969,In_438,In_1154);
and U970 (N_970,In_501,In_921);
or U971 (N_971,In_1938,In_1458);
and U972 (N_972,In_1379,In_237);
and U973 (N_973,In_1542,In_526);
nor U974 (N_974,In_1804,In_2434);
nor U975 (N_975,In_256,In_1739);
nor U976 (N_976,In_812,In_1180);
nor U977 (N_977,In_2388,In_1460);
nand U978 (N_978,In_1268,In_1298);
nor U979 (N_979,In_190,In_2293);
xor U980 (N_980,In_2142,In_667);
nand U981 (N_981,In_2411,In_2008);
and U982 (N_982,In_1294,In_599);
or U983 (N_983,In_2419,In_1068);
nor U984 (N_984,In_1471,In_2137);
or U985 (N_985,In_185,In_2380);
and U986 (N_986,In_533,In_834);
or U987 (N_987,In_129,In_2382);
or U988 (N_988,In_2199,In_776);
or U989 (N_989,In_97,In_2143);
and U990 (N_990,In_1769,In_1925);
nor U991 (N_991,In_188,In_1960);
and U992 (N_992,In_1487,In_498);
xor U993 (N_993,In_2329,In_142);
or U994 (N_994,In_631,In_93);
and U995 (N_995,In_1533,In_878);
nand U996 (N_996,In_1454,In_1428);
or U997 (N_997,In_9,In_2113);
nor U998 (N_998,In_1562,In_606);
and U999 (N_999,In_1800,In_741);
xor U1000 (N_1000,In_114,In_515);
or U1001 (N_1001,In_1849,In_869);
nor U1002 (N_1002,In_777,In_2240);
nand U1003 (N_1003,In_1123,In_1061);
nor U1004 (N_1004,In_2229,In_2373);
nor U1005 (N_1005,In_638,In_530);
or U1006 (N_1006,In_2435,In_397);
and U1007 (N_1007,In_1930,In_2092);
and U1008 (N_1008,In_387,In_1281);
or U1009 (N_1009,In_2463,In_1603);
nand U1010 (N_1010,In_578,In_624);
or U1011 (N_1011,In_836,In_2133);
and U1012 (N_1012,In_45,In_2235);
and U1013 (N_1013,In_905,In_1889);
or U1014 (N_1014,In_234,In_1553);
nor U1015 (N_1015,In_233,In_2402);
or U1016 (N_1016,In_1989,In_1020);
nand U1017 (N_1017,In_689,In_900);
or U1018 (N_1018,In_926,In_314);
nor U1019 (N_1019,In_1292,In_315);
nand U1020 (N_1020,In_1400,In_55);
nand U1021 (N_1021,In_566,In_437);
xor U1022 (N_1022,In_717,In_1271);
and U1023 (N_1023,In_1138,In_652);
and U1024 (N_1024,In_1875,In_145);
or U1025 (N_1025,In_1876,In_2226);
and U1026 (N_1026,In_736,In_1605);
nand U1027 (N_1027,In_87,In_1970);
and U1028 (N_1028,In_385,In_742);
nand U1029 (N_1029,In_1709,In_929);
or U1030 (N_1030,In_319,In_723);
xor U1031 (N_1031,In_304,In_920);
nor U1032 (N_1032,In_961,In_743);
nor U1033 (N_1033,In_354,In_762);
or U1034 (N_1034,In_1300,In_2287);
nand U1035 (N_1035,In_1244,In_625);
and U1036 (N_1036,In_253,In_2267);
nor U1037 (N_1037,In_1156,In_1737);
nor U1038 (N_1038,In_981,In_244);
or U1039 (N_1039,In_2385,In_2108);
or U1040 (N_1040,In_2067,In_1213);
and U1041 (N_1041,In_451,In_1440);
xnor U1042 (N_1042,In_2299,In_605);
nor U1043 (N_1043,In_1958,In_1506);
and U1044 (N_1044,In_433,In_2367);
nor U1045 (N_1045,In_2085,In_941);
and U1046 (N_1046,In_1071,In_2221);
nand U1047 (N_1047,In_1878,In_2205);
xnor U1048 (N_1048,In_1287,In_602);
xnor U1049 (N_1049,In_1640,In_1283);
and U1050 (N_1050,In_1051,In_1256);
or U1051 (N_1051,In_1602,In_2069);
xor U1052 (N_1052,In_1845,In_1690);
or U1053 (N_1053,In_211,In_1632);
or U1054 (N_1054,In_22,In_1223);
nor U1055 (N_1055,In_1651,In_2024);
and U1056 (N_1056,In_381,In_2498);
and U1057 (N_1057,In_2088,In_842);
nand U1058 (N_1058,In_1764,In_1914);
and U1059 (N_1059,In_175,In_903);
nor U1060 (N_1060,In_1529,In_1355);
nand U1061 (N_1061,In_350,In_167);
and U1062 (N_1062,In_1434,In_1767);
nand U1063 (N_1063,In_1184,In_261);
or U1064 (N_1064,In_1577,In_153);
and U1065 (N_1065,In_562,In_645);
nor U1066 (N_1066,In_221,In_2214);
nor U1067 (N_1067,In_2274,In_1708);
nor U1068 (N_1068,In_2386,In_760);
nor U1069 (N_1069,In_119,In_1834);
nor U1070 (N_1070,In_1544,In_1002);
nor U1071 (N_1071,In_2208,In_1038);
and U1072 (N_1072,In_335,In_1799);
nand U1073 (N_1073,In_837,In_2379);
nand U1074 (N_1074,In_449,In_29);
nor U1075 (N_1075,In_635,In_2482);
nand U1076 (N_1076,In_1272,In_1813);
or U1077 (N_1077,In_1027,In_2222);
nor U1078 (N_1078,In_14,In_2034);
and U1079 (N_1079,In_794,In_1345);
or U1080 (N_1080,In_1911,In_2197);
nand U1081 (N_1081,In_2243,In_2156);
xnor U1082 (N_1082,In_1384,In_1654);
xnor U1083 (N_1083,In_2193,In_1828);
nor U1084 (N_1084,In_874,In_470);
and U1085 (N_1085,In_816,In_182);
nor U1086 (N_1086,In_1148,In_1406);
nand U1087 (N_1087,In_583,In_1404);
xor U1088 (N_1088,In_937,In_263);
nor U1089 (N_1089,In_1118,In_33);
nand U1090 (N_1090,In_2179,In_753);
xor U1091 (N_1091,In_630,In_1241);
nor U1092 (N_1092,In_568,In_2485);
nand U1093 (N_1093,In_2251,In_1289);
and U1094 (N_1094,In_535,In_2131);
nand U1095 (N_1095,In_1756,In_1264);
or U1096 (N_1096,In_1078,In_1361);
nor U1097 (N_1097,In_1572,In_1126);
and U1098 (N_1098,In_198,In_1691);
or U1099 (N_1099,In_1411,In_1330);
and U1100 (N_1100,In_1826,In_561);
or U1101 (N_1101,In_674,In_1948);
or U1102 (N_1102,In_1527,In_2019);
xnor U1103 (N_1103,In_2360,In_927);
or U1104 (N_1104,In_230,In_2147);
nand U1105 (N_1105,In_2004,In_677);
nor U1106 (N_1106,In_1396,In_2234);
or U1107 (N_1107,In_305,In_2126);
nand U1108 (N_1108,In_279,In_1841);
or U1109 (N_1109,In_1206,In_2336);
nand U1110 (N_1110,In_1920,In_1517);
nand U1111 (N_1111,In_443,In_1591);
nor U1112 (N_1112,In_1530,In_612);
nand U1113 (N_1113,In_942,In_90);
nand U1114 (N_1114,In_2195,In_2407);
nor U1115 (N_1115,In_1582,In_1056);
nand U1116 (N_1116,In_933,In_601);
and U1117 (N_1117,In_2256,In_1806);
and U1118 (N_1118,In_1470,In_2220);
nor U1119 (N_1119,In_1388,In_1031);
nor U1120 (N_1120,In_988,In_1814);
or U1121 (N_1121,In_1522,In_2410);
nand U1122 (N_1122,In_2324,In_358);
nor U1123 (N_1123,In_2381,In_1069);
and U1124 (N_1124,In_323,In_1447);
or U1125 (N_1125,In_953,In_1862);
nand U1126 (N_1126,In_2135,In_1778);
nand U1127 (N_1127,In_322,In_1230);
and U1128 (N_1128,In_1332,In_484);
and U1129 (N_1129,In_2209,In_1802);
and U1130 (N_1130,In_174,In_467);
and U1131 (N_1131,In_1525,In_2000);
xor U1132 (N_1132,In_732,In_572);
and U1133 (N_1133,In_1353,In_1898);
nand U1134 (N_1134,In_569,In_1098);
or U1135 (N_1135,In_428,In_420);
nor U1136 (N_1136,In_459,In_1541);
and U1137 (N_1137,In_2308,In_1093);
and U1138 (N_1138,In_416,In_539);
and U1139 (N_1139,In_939,In_361);
or U1140 (N_1140,In_610,In_1656);
xor U1141 (N_1141,In_826,In_1679);
nand U1142 (N_1142,In_1459,In_52);
nor U1143 (N_1143,In_1030,In_108);
or U1144 (N_1144,In_346,In_1060);
nand U1145 (N_1145,In_2383,In_1975);
xor U1146 (N_1146,In_414,In_555);
xor U1147 (N_1147,In_513,In_2087);
or U1148 (N_1148,In_446,In_1661);
nand U1149 (N_1149,In_2352,In_144);
nand U1150 (N_1150,In_160,In_83);
xnor U1151 (N_1151,In_2338,In_1952);
xor U1152 (N_1152,In_2003,In_2496);
or U1153 (N_1153,In_1818,In_541);
or U1154 (N_1154,In_92,In_1310);
nor U1155 (N_1155,In_737,In_697);
nor U1156 (N_1156,In_1966,In_893);
nand U1157 (N_1157,In_1775,In_1567);
nand U1158 (N_1158,In_73,In_310);
and U1159 (N_1159,In_1667,In_402);
nand U1160 (N_1160,In_2152,In_2401);
xor U1161 (N_1161,In_1037,In_982);
nand U1162 (N_1162,In_1074,In_2261);
nand U1163 (N_1163,In_520,In_250);
and U1164 (N_1164,In_1101,In_862);
or U1165 (N_1165,In_391,In_970);
or U1166 (N_1166,In_962,In_2490);
or U1167 (N_1167,In_277,In_307);
or U1168 (N_1168,In_2039,In_2436);
nor U1169 (N_1169,In_2189,In_1884);
and U1170 (N_1170,In_1012,In_2167);
or U1171 (N_1171,In_173,In_944);
nand U1172 (N_1172,In_1055,In_1438);
nor U1173 (N_1173,In_1779,In_1674);
nor U1174 (N_1174,In_2094,In_891);
or U1175 (N_1175,In_343,In_1627);
nor U1176 (N_1176,In_493,In_472);
or U1177 (N_1177,In_908,In_1214);
and U1178 (N_1178,In_2245,In_200);
nor U1179 (N_1179,In_2288,In_765);
nand U1180 (N_1180,In_1192,In_2296);
nor U1181 (N_1181,In_949,In_2086);
and U1182 (N_1182,In_65,In_1978);
xnor U1183 (N_1183,In_1367,In_2168);
or U1184 (N_1184,In_2473,In_2146);
and U1185 (N_1185,In_1844,In_406);
nor U1186 (N_1186,In_975,In_968);
and U1187 (N_1187,In_422,In_993);
or U1188 (N_1188,In_2202,In_281);
and U1189 (N_1189,In_2201,In_236);
or U1190 (N_1190,In_2418,In_2233);
nor U1191 (N_1191,In_2425,In_1132);
nand U1192 (N_1192,In_2300,In_1540);
and U1193 (N_1193,In_123,In_1847);
or U1194 (N_1194,In_466,In_1033);
and U1195 (N_1195,In_1199,In_163);
and U1196 (N_1196,In_618,In_1742);
or U1197 (N_1197,In_2225,In_954);
nor U1198 (N_1198,In_1809,In_1251);
nor U1199 (N_1199,In_1451,In_1746);
nand U1200 (N_1200,In_2454,In_1749);
nand U1201 (N_1201,In_1095,In_88);
nand U1202 (N_1202,In_2370,In_177);
nand U1203 (N_1203,In_1723,In_1965);
and U1204 (N_1204,In_2196,In_379);
xnor U1205 (N_1205,In_1815,In_1863);
nand U1206 (N_1206,In_1894,In_989);
nor U1207 (N_1207,In_896,In_1626);
nor U1208 (N_1208,In_2444,In_383);
or U1209 (N_1209,In_1110,In_2455);
nor U1210 (N_1210,In_747,In_1835);
nand U1211 (N_1211,In_2351,In_168);
or U1212 (N_1212,In_2423,In_246);
nor U1213 (N_1213,In_637,In_2474);
and U1214 (N_1214,In_2355,In_1284);
or U1215 (N_1215,In_1259,In_2489);
nor U1216 (N_1216,In_838,In_1973);
xnor U1217 (N_1217,In_471,In_1594);
nand U1218 (N_1218,In_706,In_69);
or U1219 (N_1219,In_2456,In_2390);
nand U1220 (N_1220,In_2359,In_1249);
and U1221 (N_1221,In_3,In_300);
nand U1222 (N_1222,In_2348,In_994);
or U1223 (N_1223,In_2446,In_2190);
nand U1224 (N_1224,In_790,In_1119);
nand U1225 (N_1225,In_488,In_39);
and U1226 (N_1226,In_950,In_418);
nand U1227 (N_1227,In_1472,In_146);
and U1228 (N_1228,In_2059,In_1507);
nor U1229 (N_1229,In_1851,In_1432);
or U1230 (N_1230,In_1059,In_37);
or U1231 (N_1231,In_2117,In_2254);
xnor U1232 (N_1232,In_768,In_2448);
nand U1233 (N_1233,In_1927,In_557);
nor U1234 (N_1234,In_1483,In_1968);
and U1235 (N_1235,In_1116,In_1604);
and U1236 (N_1236,In_1528,In_2123);
and U1237 (N_1237,In_2306,In_1501);
nor U1238 (N_1238,In_1988,In_892);
nor U1239 (N_1239,In_2404,In_955);
and U1240 (N_1240,In_64,In_877);
or U1241 (N_1241,In_1612,In_1089);
or U1242 (N_1242,In_1539,In_2321);
and U1243 (N_1243,In_1639,In_481);
and U1244 (N_1244,In_1576,In_972);
or U1245 (N_1245,In_748,In_1606);
xor U1246 (N_1246,In_733,In_2119);
nand U1247 (N_1247,In_1873,In_430);
or U1248 (N_1248,In_31,In_1303);
nand U1249 (N_1249,In_172,In_2265);
or U1250 (N_1250,In_2373,In_1583);
or U1251 (N_1251,In_223,In_1804);
nand U1252 (N_1252,In_855,In_1618);
xor U1253 (N_1253,In_1529,In_1850);
xor U1254 (N_1254,In_806,In_2436);
nor U1255 (N_1255,In_2024,In_1768);
nor U1256 (N_1256,In_848,In_1851);
nand U1257 (N_1257,In_1087,In_2486);
nand U1258 (N_1258,In_1469,In_2383);
and U1259 (N_1259,In_530,In_486);
nand U1260 (N_1260,In_72,In_451);
and U1261 (N_1261,In_1991,In_603);
nor U1262 (N_1262,In_422,In_2498);
nand U1263 (N_1263,In_1189,In_1915);
nor U1264 (N_1264,In_704,In_2044);
nor U1265 (N_1265,In_477,In_726);
nand U1266 (N_1266,In_678,In_879);
nor U1267 (N_1267,In_766,In_1196);
nor U1268 (N_1268,In_1057,In_1330);
nor U1269 (N_1269,In_2150,In_1718);
nor U1270 (N_1270,In_1665,In_2176);
nand U1271 (N_1271,In_2110,In_2479);
xnor U1272 (N_1272,In_1613,In_850);
and U1273 (N_1273,In_1536,In_336);
nand U1274 (N_1274,In_484,In_784);
nor U1275 (N_1275,In_1393,In_1499);
nand U1276 (N_1276,In_1326,In_1690);
xor U1277 (N_1277,In_873,In_1559);
nor U1278 (N_1278,In_1798,In_1593);
and U1279 (N_1279,In_1842,In_1589);
nand U1280 (N_1280,In_2175,In_1852);
nand U1281 (N_1281,In_1283,In_2106);
or U1282 (N_1282,In_1136,In_1687);
nor U1283 (N_1283,In_1022,In_1658);
nand U1284 (N_1284,In_555,In_2434);
or U1285 (N_1285,In_744,In_150);
nand U1286 (N_1286,In_422,In_2373);
xnor U1287 (N_1287,In_337,In_1210);
or U1288 (N_1288,In_781,In_1998);
and U1289 (N_1289,In_461,In_2357);
and U1290 (N_1290,In_424,In_1377);
or U1291 (N_1291,In_854,In_1372);
or U1292 (N_1292,In_723,In_1532);
and U1293 (N_1293,In_858,In_1715);
nand U1294 (N_1294,In_1958,In_926);
nor U1295 (N_1295,In_1729,In_407);
and U1296 (N_1296,In_721,In_2101);
xnor U1297 (N_1297,In_1313,In_58);
or U1298 (N_1298,In_1201,In_199);
and U1299 (N_1299,In_2205,In_339);
or U1300 (N_1300,In_2242,In_1335);
or U1301 (N_1301,In_2330,In_1830);
nand U1302 (N_1302,In_480,In_1263);
or U1303 (N_1303,In_2067,In_2353);
xnor U1304 (N_1304,In_1394,In_2353);
nor U1305 (N_1305,In_1257,In_1008);
and U1306 (N_1306,In_111,In_184);
nand U1307 (N_1307,In_27,In_681);
and U1308 (N_1308,In_874,In_96);
nand U1309 (N_1309,In_1260,In_265);
or U1310 (N_1310,In_1895,In_972);
nand U1311 (N_1311,In_77,In_574);
and U1312 (N_1312,In_687,In_135);
nor U1313 (N_1313,In_1347,In_1734);
or U1314 (N_1314,In_677,In_1325);
nor U1315 (N_1315,In_1366,In_1057);
nand U1316 (N_1316,In_843,In_1219);
or U1317 (N_1317,In_349,In_1215);
xnor U1318 (N_1318,In_184,In_1331);
and U1319 (N_1319,In_1396,In_1522);
nand U1320 (N_1320,In_1760,In_896);
nor U1321 (N_1321,In_99,In_1146);
and U1322 (N_1322,In_482,In_1510);
or U1323 (N_1323,In_2361,In_1132);
nand U1324 (N_1324,In_1886,In_1908);
or U1325 (N_1325,In_201,In_1674);
nor U1326 (N_1326,In_514,In_1365);
nor U1327 (N_1327,In_177,In_741);
nand U1328 (N_1328,In_1449,In_2131);
nand U1329 (N_1329,In_1725,In_613);
nand U1330 (N_1330,In_424,In_127);
xor U1331 (N_1331,In_568,In_54);
nor U1332 (N_1332,In_1809,In_635);
nor U1333 (N_1333,In_1368,In_1691);
or U1334 (N_1334,In_267,In_1872);
nand U1335 (N_1335,In_1763,In_1056);
and U1336 (N_1336,In_1602,In_2291);
and U1337 (N_1337,In_129,In_2268);
and U1338 (N_1338,In_1383,In_2238);
or U1339 (N_1339,In_437,In_521);
nand U1340 (N_1340,In_904,In_1997);
or U1341 (N_1341,In_1587,In_176);
or U1342 (N_1342,In_1705,In_1071);
nand U1343 (N_1343,In_670,In_801);
or U1344 (N_1344,In_1493,In_18);
and U1345 (N_1345,In_953,In_805);
nor U1346 (N_1346,In_1212,In_1673);
nand U1347 (N_1347,In_176,In_1753);
and U1348 (N_1348,In_220,In_287);
nor U1349 (N_1349,In_1812,In_1377);
or U1350 (N_1350,In_46,In_2365);
xor U1351 (N_1351,In_1450,In_312);
nand U1352 (N_1352,In_1408,In_1308);
nor U1353 (N_1353,In_355,In_1436);
nand U1354 (N_1354,In_1468,In_2334);
nor U1355 (N_1355,In_1879,In_1463);
nor U1356 (N_1356,In_649,In_180);
or U1357 (N_1357,In_699,In_672);
and U1358 (N_1358,In_1869,In_1808);
xor U1359 (N_1359,In_2000,In_1126);
nand U1360 (N_1360,In_1322,In_358);
or U1361 (N_1361,In_1433,In_226);
xor U1362 (N_1362,In_759,In_890);
nand U1363 (N_1363,In_110,In_2187);
xnor U1364 (N_1364,In_2059,In_2400);
nand U1365 (N_1365,In_453,In_1833);
or U1366 (N_1366,In_2418,In_384);
nor U1367 (N_1367,In_1498,In_645);
or U1368 (N_1368,In_450,In_751);
and U1369 (N_1369,In_1071,In_948);
nand U1370 (N_1370,In_1188,In_394);
nand U1371 (N_1371,In_564,In_1850);
nand U1372 (N_1372,In_1558,In_2174);
xor U1373 (N_1373,In_1289,In_689);
or U1374 (N_1374,In_2363,In_1079);
nor U1375 (N_1375,In_1223,In_231);
nor U1376 (N_1376,In_1831,In_1996);
xor U1377 (N_1377,In_2266,In_1404);
nand U1378 (N_1378,In_402,In_804);
or U1379 (N_1379,In_1125,In_2380);
or U1380 (N_1380,In_1638,In_264);
or U1381 (N_1381,In_1079,In_919);
or U1382 (N_1382,In_1776,In_2233);
xnor U1383 (N_1383,In_2336,In_269);
or U1384 (N_1384,In_518,In_1430);
nor U1385 (N_1385,In_2142,In_849);
nor U1386 (N_1386,In_608,In_1704);
or U1387 (N_1387,In_2299,In_420);
and U1388 (N_1388,In_760,In_105);
nor U1389 (N_1389,In_1850,In_74);
nor U1390 (N_1390,In_1249,In_1537);
nor U1391 (N_1391,In_273,In_858);
nor U1392 (N_1392,In_1214,In_1446);
nand U1393 (N_1393,In_152,In_618);
and U1394 (N_1394,In_491,In_1475);
nor U1395 (N_1395,In_347,In_2082);
or U1396 (N_1396,In_2393,In_1941);
nor U1397 (N_1397,In_791,In_1981);
nor U1398 (N_1398,In_575,In_2155);
xor U1399 (N_1399,In_2269,In_459);
or U1400 (N_1400,In_2474,In_1233);
and U1401 (N_1401,In_1038,In_2447);
or U1402 (N_1402,In_440,In_482);
nand U1403 (N_1403,In_1308,In_140);
or U1404 (N_1404,In_1570,In_1277);
nor U1405 (N_1405,In_777,In_360);
nor U1406 (N_1406,In_1089,In_2261);
nand U1407 (N_1407,In_2240,In_1003);
or U1408 (N_1408,In_689,In_369);
or U1409 (N_1409,In_447,In_1685);
nor U1410 (N_1410,In_1371,In_368);
or U1411 (N_1411,In_2310,In_2433);
nor U1412 (N_1412,In_2220,In_1604);
xor U1413 (N_1413,In_2093,In_1121);
nand U1414 (N_1414,In_485,In_39);
nor U1415 (N_1415,In_2010,In_1445);
or U1416 (N_1416,In_878,In_436);
nand U1417 (N_1417,In_760,In_1119);
xor U1418 (N_1418,In_140,In_661);
nand U1419 (N_1419,In_2117,In_1275);
nor U1420 (N_1420,In_67,In_2436);
nand U1421 (N_1421,In_962,In_740);
nand U1422 (N_1422,In_421,In_2323);
and U1423 (N_1423,In_898,In_145);
nand U1424 (N_1424,In_441,In_619);
nor U1425 (N_1425,In_2198,In_1750);
and U1426 (N_1426,In_812,In_240);
and U1427 (N_1427,In_1550,In_1770);
or U1428 (N_1428,In_345,In_780);
nor U1429 (N_1429,In_1177,In_260);
nand U1430 (N_1430,In_2287,In_1029);
and U1431 (N_1431,In_2027,In_1734);
and U1432 (N_1432,In_1716,In_2053);
nor U1433 (N_1433,In_1358,In_1741);
or U1434 (N_1434,In_606,In_854);
nand U1435 (N_1435,In_527,In_2019);
nand U1436 (N_1436,In_291,In_2253);
nor U1437 (N_1437,In_522,In_89);
nor U1438 (N_1438,In_2054,In_288);
and U1439 (N_1439,In_1951,In_1745);
and U1440 (N_1440,In_1039,In_315);
nand U1441 (N_1441,In_1632,In_925);
nor U1442 (N_1442,In_635,In_1214);
nor U1443 (N_1443,In_224,In_332);
or U1444 (N_1444,In_1924,In_2069);
and U1445 (N_1445,In_2312,In_1084);
xor U1446 (N_1446,In_2341,In_2128);
xnor U1447 (N_1447,In_652,In_336);
nand U1448 (N_1448,In_1145,In_608);
or U1449 (N_1449,In_1581,In_2400);
nor U1450 (N_1450,In_851,In_388);
xor U1451 (N_1451,In_959,In_381);
and U1452 (N_1452,In_2217,In_2171);
xnor U1453 (N_1453,In_2426,In_1849);
and U1454 (N_1454,In_986,In_1775);
or U1455 (N_1455,In_1045,In_451);
and U1456 (N_1456,In_1208,In_291);
or U1457 (N_1457,In_2177,In_1564);
nor U1458 (N_1458,In_394,In_2263);
and U1459 (N_1459,In_1041,In_1776);
nand U1460 (N_1460,In_1486,In_984);
nand U1461 (N_1461,In_355,In_2190);
xor U1462 (N_1462,In_1882,In_403);
or U1463 (N_1463,In_2097,In_1845);
nand U1464 (N_1464,In_974,In_784);
nand U1465 (N_1465,In_2319,In_1288);
and U1466 (N_1466,In_1659,In_2425);
nand U1467 (N_1467,In_2430,In_1438);
nand U1468 (N_1468,In_476,In_243);
and U1469 (N_1469,In_335,In_988);
nor U1470 (N_1470,In_840,In_1863);
or U1471 (N_1471,In_706,In_3);
or U1472 (N_1472,In_2206,In_419);
nor U1473 (N_1473,In_1830,In_1105);
and U1474 (N_1474,In_47,In_2492);
nor U1475 (N_1475,In_1722,In_93);
xor U1476 (N_1476,In_2222,In_231);
or U1477 (N_1477,In_1050,In_1900);
nor U1478 (N_1478,In_1425,In_1614);
nand U1479 (N_1479,In_1225,In_2425);
nand U1480 (N_1480,In_2166,In_1122);
nor U1481 (N_1481,In_193,In_790);
nand U1482 (N_1482,In_1899,In_2356);
nand U1483 (N_1483,In_656,In_2472);
and U1484 (N_1484,In_1229,In_2455);
or U1485 (N_1485,In_423,In_1741);
or U1486 (N_1486,In_1780,In_371);
nor U1487 (N_1487,In_1191,In_367);
nor U1488 (N_1488,In_495,In_1662);
or U1489 (N_1489,In_1467,In_2055);
nor U1490 (N_1490,In_1739,In_865);
or U1491 (N_1491,In_1298,In_628);
and U1492 (N_1492,In_786,In_654);
and U1493 (N_1493,In_1019,In_316);
nand U1494 (N_1494,In_100,In_871);
or U1495 (N_1495,In_20,In_1727);
or U1496 (N_1496,In_115,In_1196);
nor U1497 (N_1497,In_363,In_2167);
nand U1498 (N_1498,In_12,In_766);
xor U1499 (N_1499,In_206,In_1844);
xor U1500 (N_1500,In_1161,In_327);
nand U1501 (N_1501,In_1169,In_2023);
nand U1502 (N_1502,In_1262,In_2237);
nor U1503 (N_1503,In_111,In_664);
nand U1504 (N_1504,In_1494,In_1917);
nand U1505 (N_1505,In_1698,In_2414);
or U1506 (N_1506,In_1139,In_852);
nor U1507 (N_1507,In_38,In_75);
or U1508 (N_1508,In_2066,In_2360);
xnor U1509 (N_1509,In_1766,In_1613);
and U1510 (N_1510,In_425,In_2328);
nand U1511 (N_1511,In_625,In_1292);
and U1512 (N_1512,In_1296,In_114);
nor U1513 (N_1513,In_1281,In_1796);
nand U1514 (N_1514,In_1315,In_1899);
and U1515 (N_1515,In_335,In_300);
and U1516 (N_1516,In_141,In_2023);
nor U1517 (N_1517,In_1098,In_938);
and U1518 (N_1518,In_2221,In_2485);
and U1519 (N_1519,In_312,In_428);
nand U1520 (N_1520,In_1179,In_611);
nand U1521 (N_1521,In_233,In_1955);
xnor U1522 (N_1522,In_20,In_800);
or U1523 (N_1523,In_373,In_380);
nand U1524 (N_1524,In_216,In_661);
nor U1525 (N_1525,In_1699,In_1596);
or U1526 (N_1526,In_859,In_2329);
or U1527 (N_1527,In_853,In_2340);
nand U1528 (N_1528,In_1756,In_1979);
and U1529 (N_1529,In_1801,In_1509);
or U1530 (N_1530,In_124,In_1892);
and U1531 (N_1531,In_718,In_2181);
nand U1532 (N_1532,In_1541,In_1209);
nor U1533 (N_1533,In_1281,In_1805);
nand U1534 (N_1534,In_1197,In_390);
nor U1535 (N_1535,In_1068,In_254);
and U1536 (N_1536,In_313,In_892);
xnor U1537 (N_1537,In_1789,In_300);
nor U1538 (N_1538,In_1809,In_956);
or U1539 (N_1539,In_1135,In_667);
nand U1540 (N_1540,In_872,In_2470);
nand U1541 (N_1541,In_589,In_2497);
or U1542 (N_1542,In_18,In_1654);
nor U1543 (N_1543,In_1821,In_1083);
nand U1544 (N_1544,In_912,In_2185);
xnor U1545 (N_1545,In_2064,In_1420);
or U1546 (N_1546,In_824,In_1834);
or U1547 (N_1547,In_74,In_1710);
nand U1548 (N_1548,In_1423,In_2193);
and U1549 (N_1549,In_734,In_1522);
and U1550 (N_1550,In_2073,In_1108);
nor U1551 (N_1551,In_1011,In_1491);
and U1552 (N_1552,In_2249,In_1508);
nor U1553 (N_1553,In_2039,In_45);
nand U1554 (N_1554,In_1511,In_2377);
or U1555 (N_1555,In_2385,In_95);
nand U1556 (N_1556,In_2267,In_763);
xnor U1557 (N_1557,In_1297,In_2067);
or U1558 (N_1558,In_756,In_2368);
and U1559 (N_1559,In_134,In_1218);
nand U1560 (N_1560,In_1387,In_2163);
or U1561 (N_1561,In_438,In_1408);
or U1562 (N_1562,In_2408,In_2483);
nor U1563 (N_1563,In_424,In_1218);
and U1564 (N_1564,In_978,In_1319);
xnor U1565 (N_1565,In_902,In_1831);
xnor U1566 (N_1566,In_201,In_422);
and U1567 (N_1567,In_1484,In_1493);
nor U1568 (N_1568,In_631,In_1219);
nor U1569 (N_1569,In_1618,In_1624);
nand U1570 (N_1570,In_1010,In_1829);
or U1571 (N_1571,In_2153,In_579);
and U1572 (N_1572,In_1248,In_1928);
or U1573 (N_1573,In_807,In_1829);
nor U1574 (N_1574,In_2390,In_602);
nor U1575 (N_1575,In_964,In_2228);
nand U1576 (N_1576,In_1171,In_1115);
nand U1577 (N_1577,In_1870,In_745);
xor U1578 (N_1578,In_1590,In_1784);
xor U1579 (N_1579,In_312,In_97);
xnor U1580 (N_1580,In_1679,In_825);
and U1581 (N_1581,In_1016,In_1509);
nor U1582 (N_1582,In_1468,In_2028);
nor U1583 (N_1583,In_1615,In_676);
or U1584 (N_1584,In_159,In_825);
or U1585 (N_1585,In_2098,In_625);
nor U1586 (N_1586,In_1242,In_1689);
nor U1587 (N_1587,In_1741,In_651);
nand U1588 (N_1588,In_595,In_633);
nand U1589 (N_1589,In_1409,In_775);
xor U1590 (N_1590,In_1981,In_1259);
and U1591 (N_1591,In_1772,In_1604);
or U1592 (N_1592,In_613,In_1730);
nor U1593 (N_1593,In_518,In_389);
nand U1594 (N_1594,In_1926,In_1742);
nand U1595 (N_1595,In_29,In_588);
and U1596 (N_1596,In_2369,In_919);
nand U1597 (N_1597,In_539,In_1659);
and U1598 (N_1598,In_1021,In_410);
nand U1599 (N_1599,In_114,In_943);
nor U1600 (N_1600,In_1886,In_218);
nand U1601 (N_1601,In_2399,In_2369);
nand U1602 (N_1602,In_1453,In_1323);
or U1603 (N_1603,In_604,In_1342);
or U1604 (N_1604,In_1974,In_1108);
nand U1605 (N_1605,In_1535,In_2283);
nor U1606 (N_1606,In_816,In_1172);
nand U1607 (N_1607,In_606,In_1778);
xor U1608 (N_1608,In_1693,In_1528);
nand U1609 (N_1609,In_506,In_280);
nand U1610 (N_1610,In_1021,In_659);
and U1611 (N_1611,In_1922,In_1754);
nand U1612 (N_1612,In_727,In_1498);
nand U1613 (N_1613,In_2222,In_2245);
and U1614 (N_1614,In_2025,In_235);
nand U1615 (N_1615,In_1803,In_2142);
and U1616 (N_1616,In_551,In_341);
nand U1617 (N_1617,In_1594,In_797);
xnor U1618 (N_1618,In_476,In_2057);
or U1619 (N_1619,In_874,In_1940);
nor U1620 (N_1620,In_2147,In_1420);
nor U1621 (N_1621,In_2192,In_1640);
nand U1622 (N_1622,In_2181,In_428);
or U1623 (N_1623,In_1580,In_176);
nand U1624 (N_1624,In_1540,In_1940);
nand U1625 (N_1625,In_427,In_1951);
nand U1626 (N_1626,In_2025,In_948);
nand U1627 (N_1627,In_222,In_40);
nor U1628 (N_1628,In_1336,In_1850);
or U1629 (N_1629,In_2220,In_464);
or U1630 (N_1630,In_2024,In_896);
or U1631 (N_1631,In_2071,In_73);
nand U1632 (N_1632,In_1508,In_1524);
nor U1633 (N_1633,In_1121,In_1223);
nor U1634 (N_1634,In_366,In_1384);
nor U1635 (N_1635,In_360,In_1363);
and U1636 (N_1636,In_1222,In_223);
nor U1637 (N_1637,In_1524,In_2047);
or U1638 (N_1638,In_1383,In_2018);
nor U1639 (N_1639,In_1680,In_1138);
and U1640 (N_1640,In_162,In_1626);
nor U1641 (N_1641,In_190,In_1084);
and U1642 (N_1642,In_1694,In_575);
nor U1643 (N_1643,In_1472,In_296);
and U1644 (N_1644,In_1368,In_1069);
nor U1645 (N_1645,In_7,In_1423);
or U1646 (N_1646,In_1407,In_394);
and U1647 (N_1647,In_2434,In_1388);
xor U1648 (N_1648,In_1330,In_2319);
nor U1649 (N_1649,In_179,In_2162);
or U1650 (N_1650,In_1686,In_8);
nand U1651 (N_1651,In_853,In_1212);
xor U1652 (N_1652,In_2052,In_1986);
and U1653 (N_1653,In_2064,In_1054);
or U1654 (N_1654,In_279,In_2025);
and U1655 (N_1655,In_2138,In_284);
xnor U1656 (N_1656,In_888,In_1777);
nand U1657 (N_1657,In_1033,In_2154);
or U1658 (N_1658,In_2087,In_1352);
xor U1659 (N_1659,In_47,In_1443);
or U1660 (N_1660,In_1678,In_1083);
or U1661 (N_1661,In_761,In_80);
nand U1662 (N_1662,In_1730,In_713);
or U1663 (N_1663,In_1594,In_1495);
nand U1664 (N_1664,In_1459,In_1552);
and U1665 (N_1665,In_460,In_896);
nand U1666 (N_1666,In_408,In_603);
and U1667 (N_1667,In_509,In_567);
nand U1668 (N_1668,In_240,In_1052);
and U1669 (N_1669,In_2476,In_746);
or U1670 (N_1670,In_603,In_1785);
nand U1671 (N_1671,In_2338,In_1369);
xnor U1672 (N_1672,In_2465,In_1226);
nor U1673 (N_1673,In_793,In_1732);
nand U1674 (N_1674,In_795,In_1479);
or U1675 (N_1675,In_2281,In_1345);
and U1676 (N_1676,In_20,In_1143);
nor U1677 (N_1677,In_2207,In_1607);
and U1678 (N_1678,In_896,In_1094);
and U1679 (N_1679,In_441,In_2192);
xnor U1680 (N_1680,In_344,In_1263);
and U1681 (N_1681,In_758,In_1809);
nand U1682 (N_1682,In_2007,In_2243);
nand U1683 (N_1683,In_30,In_2309);
and U1684 (N_1684,In_455,In_1433);
nor U1685 (N_1685,In_1047,In_1602);
nand U1686 (N_1686,In_2238,In_115);
nor U1687 (N_1687,In_502,In_1376);
nor U1688 (N_1688,In_2355,In_2237);
nor U1689 (N_1689,In_1957,In_1020);
or U1690 (N_1690,In_2252,In_372);
nor U1691 (N_1691,In_2339,In_1785);
nand U1692 (N_1692,In_2248,In_2011);
and U1693 (N_1693,In_1564,In_1411);
or U1694 (N_1694,In_1968,In_870);
nand U1695 (N_1695,In_1285,In_561);
xnor U1696 (N_1696,In_1213,In_1302);
nor U1697 (N_1697,In_1385,In_947);
nor U1698 (N_1698,In_2204,In_2304);
and U1699 (N_1699,In_1803,In_958);
or U1700 (N_1700,In_2062,In_1784);
and U1701 (N_1701,In_2295,In_2350);
nor U1702 (N_1702,In_12,In_2278);
and U1703 (N_1703,In_2311,In_1437);
or U1704 (N_1704,In_2075,In_2409);
or U1705 (N_1705,In_302,In_482);
xor U1706 (N_1706,In_693,In_818);
and U1707 (N_1707,In_414,In_2104);
xor U1708 (N_1708,In_660,In_2054);
nand U1709 (N_1709,In_1278,In_541);
or U1710 (N_1710,In_1414,In_832);
and U1711 (N_1711,In_1952,In_917);
nand U1712 (N_1712,In_2173,In_139);
nand U1713 (N_1713,In_1185,In_1562);
and U1714 (N_1714,In_2180,In_1482);
nand U1715 (N_1715,In_271,In_2268);
or U1716 (N_1716,In_276,In_587);
and U1717 (N_1717,In_1878,In_1774);
and U1718 (N_1718,In_1479,In_1930);
and U1719 (N_1719,In_919,In_667);
and U1720 (N_1720,In_730,In_161);
nor U1721 (N_1721,In_1336,In_544);
or U1722 (N_1722,In_167,In_1021);
or U1723 (N_1723,In_565,In_2400);
nand U1724 (N_1724,In_1313,In_866);
nand U1725 (N_1725,In_2275,In_1535);
nand U1726 (N_1726,In_2209,In_2432);
or U1727 (N_1727,In_2433,In_1336);
and U1728 (N_1728,In_1029,In_64);
nor U1729 (N_1729,In_2217,In_773);
nand U1730 (N_1730,In_1079,In_1696);
or U1731 (N_1731,In_877,In_332);
and U1732 (N_1732,In_2398,In_109);
and U1733 (N_1733,In_2427,In_2237);
or U1734 (N_1734,In_618,In_43);
or U1735 (N_1735,In_13,In_819);
nor U1736 (N_1736,In_1352,In_2113);
xor U1737 (N_1737,In_1359,In_231);
or U1738 (N_1738,In_638,In_1302);
or U1739 (N_1739,In_1160,In_1851);
xnor U1740 (N_1740,In_1132,In_1702);
xor U1741 (N_1741,In_39,In_1078);
or U1742 (N_1742,In_316,In_4);
or U1743 (N_1743,In_1029,In_1552);
or U1744 (N_1744,In_4,In_1808);
nand U1745 (N_1745,In_1119,In_375);
xor U1746 (N_1746,In_563,In_646);
or U1747 (N_1747,In_2285,In_219);
xnor U1748 (N_1748,In_2246,In_1861);
or U1749 (N_1749,In_811,In_1306);
xor U1750 (N_1750,In_1156,In_2452);
or U1751 (N_1751,In_2361,In_220);
nand U1752 (N_1752,In_1390,In_911);
and U1753 (N_1753,In_2037,In_324);
nor U1754 (N_1754,In_2359,In_1629);
and U1755 (N_1755,In_2436,In_2048);
nor U1756 (N_1756,In_672,In_512);
nor U1757 (N_1757,In_2268,In_2027);
and U1758 (N_1758,In_1639,In_2273);
nor U1759 (N_1759,In_1769,In_1206);
and U1760 (N_1760,In_1101,In_874);
and U1761 (N_1761,In_806,In_938);
and U1762 (N_1762,In_394,In_1150);
xor U1763 (N_1763,In_1588,In_925);
and U1764 (N_1764,In_2258,In_1721);
nor U1765 (N_1765,In_477,In_200);
or U1766 (N_1766,In_820,In_1397);
and U1767 (N_1767,In_1703,In_397);
xnor U1768 (N_1768,In_85,In_2346);
or U1769 (N_1769,In_2021,In_600);
nor U1770 (N_1770,In_2405,In_1845);
nor U1771 (N_1771,In_1504,In_1126);
nor U1772 (N_1772,In_1258,In_554);
and U1773 (N_1773,In_743,In_1896);
nor U1774 (N_1774,In_984,In_2003);
nor U1775 (N_1775,In_925,In_1994);
nor U1776 (N_1776,In_544,In_1142);
nor U1777 (N_1777,In_126,In_69);
nand U1778 (N_1778,In_1677,In_1153);
or U1779 (N_1779,In_2296,In_96);
nor U1780 (N_1780,In_2226,In_459);
or U1781 (N_1781,In_1575,In_36);
or U1782 (N_1782,In_1537,In_1432);
xnor U1783 (N_1783,In_434,In_869);
nand U1784 (N_1784,In_24,In_2294);
and U1785 (N_1785,In_865,In_1454);
and U1786 (N_1786,In_1616,In_401);
nor U1787 (N_1787,In_1513,In_1839);
and U1788 (N_1788,In_1240,In_1943);
and U1789 (N_1789,In_1256,In_2123);
nor U1790 (N_1790,In_1925,In_525);
or U1791 (N_1791,In_1429,In_2285);
and U1792 (N_1792,In_1677,In_813);
and U1793 (N_1793,In_836,In_1286);
and U1794 (N_1794,In_1731,In_2057);
and U1795 (N_1795,In_1488,In_1759);
nand U1796 (N_1796,In_336,In_1001);
and U1797 (N_1797,In_2224,In_1931);
or U1798 (N_1798,In_2386,In_176);
nand U1799 (N_1799,In_1673,In_1669);
nor U1800 (N_1800,In_769,In_912);
xnor U1801 (N_1801,In_342,In_1000);
nand U1802 (N_1802,In_1274,In_1398);
xor U1803 (N_1803,In_1760,In_1835);
nand U1804 (N_1804,In_544,In_1537);
nand U1805 (N_1805,In_1317,In_2174);
nor U1806 (N_1806,In_2052,In_216);
nor U1807 (N_1807,In_529,In_932);
nand U1808 (N_1808,In_446,In_1656);
nand U1809 (N_1809,In_515,In_115);
nand U1810 (N_1810,In_2241,In_1421);
nor U1811 (N_1811,In_1925,In_635);
nand U1812 (N_1812,In_1552,In_1698);
or U1813 (N_1813,In_2091,In_1607);
nor U1814 (N_1814,In_293,In_260);
xnor U1815 (N_1815,In_649,In_2138);
and U1816 (N_1816,In_230,In_1988);
or U1817 (N_1817,In_2098,In_2371);
nand U1818 (N_1818,In_1550,In_1615);
nor U1819 (N_1819,In_12,In_2068);
nor U1820 (N_1820,In_1078,In_1693);
and U1821 (N_1821,In_2314,In_2393);
nor U1822 (N_1822,In_1464,In_1015);
or U1823 (N_1823,In_99,In_2390);
and U1824 (N_1824,In_1634,In_2478);
xor U1825 (N_1825,In_1301,In_25);
xnor U1826 (N_1826,In_1723,In_1699);
or U1827 (N_1827,In_946,In_1061);
or U1828 (N_1828,In_915,In_1650);
and U1829 (N_1829,In_1171,In_50);
nor U1830 (N_1830,In_1145,In_623);
or U1831 (N_1831,In_2259,In_1567);
or U1832 (N_1832,In_2137,In_1643);
and U1833 (N_1833,In_2292,In_1745);
nor U1834 (N_1834,In_1827,In_1165);
nor U1835 (N_1835,In_247,In_285);
and U1836 (N_1836,In_1507,In_965);
or U1837 (N_1837,In_1517,In_1307);
nor U1838 (N_1838,In_1662,In_535);
nor U1839 (N_1839,In_1286,In_2017);
and U1840 (N_1840,In_1341,In_314);
nor U1841 (N_1841,In_566,In_267);
or U1842 (N_1842,In_673,In_1069);
nor U1843 (N_1843,In_1415,In_102);
and U1844 (N_1844,In_1588,In_621);
or U1845 (N_1845,In_960,In_1450);
nor U1846 (N_1846,In_827,In_96);
nor U1847 (N_1847,In_2212,In_1585);
or U1848 (N_1848,In_322,In_475);
and U1849 (N_1849,In_821,In_2382);
or U1850 (N_1850,In_731,In_1247);
and U1851 (N_1851,In_2129,In_2133);
nor U1852 (N_1852,In_1418,In_1904);
xor U1853 (N_1853,In_2049,In_936);
nand U1854 (N_1854,In_1174,In_422);
nor U1855 (N_1855,In_591,In_632);
nor U1856 (N_1856,In_1919,In_1287);
and U1857 (N_1857,In_1804,In_702);
nand U1858 (N_1858,In_420,In_813);
and U1859 (N_1859,In_1198,In_1937);
xor U1860 (N_1860,In_1895,In_2194);
nand U1861 (N_1861,In_1981,In_619);
nand U1862 (N_1862,In_767,In_2003);
nor U1863 (N_1863,In_2207,In_1372);
nor U1864 (N_1864,In_2101,In_905);
or U1865 (N_1865,In_45,In_452);
nor U1866 (N_1866,In_472,In_1934);
nand U1867 (N_1867,In_1869,In_1879);
and U1868 (N_1868,In_1373,In_767);
nand U1869 (N_1869,In_2398,In_1706);
nor U1870 (N_1870,In_54,In_2345);
or U1871 (N_1871,In_1307,In_756);
nand U1872 (N_1872,In_1648,In_1204);
and U1873 (N_1873,In_281,In_860);
nand U1874 (N_1874,In_2308,In_86);
or U1875 (N_1875,In_147,In_841);
nor U1876 (N_1876,In_1902,In_2246);
or U1877 (N_1877,In_1110,In_2396);
nand U1878 (N_1878,In_1557,In_21);
and U1879 (N_1879,In_2476,In_1288);
and U1880 (N_1880,In_425,In_907);
nor U1881 (N_1881,In_1259,In_831);
or U1882 (N_1882,In_901,In_1750);
and U1883 (N_1883,In_1559,In_1792);
and U1884 (N_1884,In_1065,In_1873);
and U1885 (N_1885,In_1143,In_137);
or U1886 (N_1886,In_1611,In_1495);
or U1887 (N_1887,In_1020,In_1521);
xor U1888 (N_1888,In_1815,In_1731);
or U1889 (N_1889,In_1151,In_885);
and U1890 (N_1890,In_2214,In_1876);
or U1891 (N_1891,In_1823,In_1209);
xor U1892 (N_1892,In_2106,In_850);
nor U1893 (N_1893,In_1123,In_2328);
nand U1894 (N_1894,In_2012,In_1373);
or U1895 (N_1895,In_330,In_341);
and U1896 (N_1896,In_844,In_498);
nand U1897 (N_1897,In_2192,In_950);
xor U1898 (N_1898,In_1349,In_1498);
nor U1899 (N_1899,In_1989,In_1722);
nor U1900 (N_1900,In_2416,In_2187);
nor U1901 (N_1901,In_1427,In_1752);
nor U1902 (N_1902,In_1874,In_1290);
and U1903 (N_1903,In_2364,In_1898);
nor U1904 (N_1904,In_1049,In_1576);
nor U1905 (N_1905,In_1734,In_461);
and U1906 (N_1906,In_1087,In_656);
and U1907 (N_1907,In_1039,In_211);
or U1908 (N_1908,In_969,In_2420);
nor U1909 (N_1909,In_1825,In_2114);
or U1910 (N_1910,In_259,In_2446);
nand U1911 (N_1911,In_969,In_2192);
and U1912 (N_1912,In_1574,In_453);
and U1913 (N_1913,In_177,In_2267);
nand U1914 (N_1914,In_624,In_550);
and U1915 (N_1915,In_770,In_1308);
nor U1916 (N_1916,In_1860,In_2487);
or U1917 (N_1917,In_1980,In_163);
xor U1918 (N_1918,In_647,In_274);
nand U1919 (N_1919,In_263,In_2149);
or U1920 (N_1920,In_454,In_1946);
and U1921 (N_1921,In_629,In_2223);
and U1922 (N_1922,In_1112,In_1828);
nor U1923 (N_1923,In_2349,In_2340);
nor U1924 (N_1924,In_1472,In_827);
nand U1925 (N_1925,In_2199,In_736);
and U1926 (N_1926,In_2262,In_2206);
or U1927 (N_1927,In_2411,In_720);
nand U1928 (N_1928,In_90,In_1917);
xnor U1929 (N_1929,In_1839,In_2488);
nand U1930 (N_1930,In_1646,In_1349);
nand U1931 (N_1931,In_1152,In_404);
nor U1932 (N_1932,In_1621,In_202);
nand U1933 (N_1933,In_1839,In_1037);
or U1934 (N_1934,In_2245,In_278);
xor U1935 (N_1935,In_1746,In_1765);
nand U1936 (N_1936,In_271,In_428);
nor U1937 (N_1937,In_1152,In_1448);
or U1938 (N_1938,In_2319,In_1079);
or U1939 (N_1939,In_1768,In_2464);
xnor U1940 (N_1940,In_1766,In_892);
or U1941 (N_1941,In_227,In_92);
and U1942 (N_1942,In_747,In_2159);
nor U1943 (N_1943,In_589,In_1946);
and U1944 (N_1944,In_2176,In_1411);
nor U1945 (N_1945,In_704,In_1676);
or U1946 (N_1946,In_252,In_296);
and U1947 (N_1947,In_2354,In_878);
nand U1948 (N_1948,In_2490,In_2219);
or U1949 (N_1949,In_1988,In_1757);
or U1950 (N_1950,In_32,In_664);
nor U1951 (N_1951,In_1996,In_1509);
and U1952 (N_1952,In_1106,In_1563);
and U1953 (N_1953,In_2227,In_2062);
and U1954 (N_1954,In_1405,In_1974);
xnor U1955 (N_1955,In_1266,In_1882);
nor U1956 (N_1956,In_2263,In_1493);
or U1957 (N_1957,In_1421,In_1389);
and U1958 (N_1958,In_2346,In_182);
nand U1959 (N_1959,In_1888,In_1963);
nand U1960 (N_1960,In_97,In_1156);
or U1961 (N_1961,In_1282,In_1714);
nand U1962 (N_1962,In_138,In_636);
or U1963 (N_1963,In_1739,In_319);
nor U1964 (N_1964,In_1063,In_1390);
nor U1965 (N_1965,In_270,In_1127);
and U1966 (N_1966,In_819,In_328);
nand U1967 (N_1967,In_411,In_59);
nand U1968 (N_1968,In_425,In_322);
or U1969 (N_1969,In_1390,In_950);
or U1970 (N_1970,In_508,In_997);
or U1971 (N_1971,In_1412,In_1707);
or U1972 (N_1972,In_743,In_725);
xor U1973 (N_1973,In_1831,In_2303);
or U1974 (N_1974,In_2047,In_2145);
nand U1975 (N_1975,In_2217,In_2300);
nand U1976 (N_1976,In_2475,In_1334);
xnor U1977 (N_1977,In_139,In_604);
nor U1978 (N_1978,In_1473,In_1168);
and U1979 (N_1979,In_71,In_693);
and U1980 (N_1980,In_1543,In_2389);
nand U1981 (N_1981,In_113,In_1331);
nor U1982 (N_1982,In_1327,In_2454);
or U1983 (N_1983,In_2351,In_2062);
or U1984 (N_1984,In_1652,In_1928);
or U1985 (N_1985,In_2329,In_924);
or U1986 (N_1986,In_2088,In_1244);
nand U1987 (N_1987,In_1847,In_1136);
or U1988 (N_1988,In_43,In_1715);
xnor U1989 (N_1989,In_882,In_806);
nand U1990 (N_1990,In_1465,In_237);
nand U1991 (N_1991,In_1372,In_1725);
or U1992 (N_1992,In_2464,In_383);
or U1993 (N_1993,In_2206,In_1269);
or U1994 (N_1994,In_1527,In_1322);
and U1995 (N_1995,In_1392,In_2356);
and U1996 (N_1996,In_1289,In_2017);
or U1997 (N_1997,In_2050,In_2350);
or U1998 (N_1998,In_1683,In_1801);
and U1999 (N_1999,In_1546,In_382);
or U2000 (N_2000,In_2147,In_2000);
nand U2001 (N_2001,In_1133,In_350);
nor U2002 (N_2002,In_1726,In_705);
nand U2003 (N_2003,In_1225,In_179);
nand U2004 (N_2004,In_1572,In_1545);
and U2005 (N_2005,In_2074,In_1687);
nand U2006 (N_2006,In_1049,In_330);
nand U2007 (N_2007,In_727,In_55);
and U2008 (N_2008,In_2029,In_160);
xnor U2009 (N_2009,In_2163,In_849);
or U2010 (N_2010,In_1238,In_1033);
nand U2011 (N_2011,In_1049,In_2209);
xor U2012 (N_2012,In_526,In_702);
or U2013 (N_2013,In_2455,In_104);
nand U2014 (N_2014,In_2110,In_543);
or U2015 (N_2015,In_1590,In_2430);
nand U2016 (N_2016,In_835,In_2103);
and U2017 (N_2017,In_2237,In_1328);
or U2018 (N_2018,In_1822,In_941);
and U2019 (N_2019,In_708,In_1767);
or U2020 (N_2020,In_2080,In_1333);
xor U2021 (N_2021,In_1598,In_959);
and U2022 (N_2022,In_351,In_2251);
xnor U2023 (N_2023,In_945,In_1911);
nor U2024 (N_2024,In_1340,In_157);
and U2025 (N_2025,In_2299,In_1510);
and U2026 (N_2026,In_116,In_1701);
and U2027 (N_2027,In_1352,In_723);
xnor U2028 (N_2028,In_1088,In_1396);
nor U2029 (N_2029,In_900,In_2143);
or U2030 (N_2030,In_47,In_828);
and U2031 (N_2031,In_1122,In_839);
nor U2032 (N_2032,In_1419,In_1906);
and U2033 (N_2033,In_2135,In_1821);
xor U2034 (N_2034,In_1247,In_743);
or U2035 (N_2035,In_1337,In_85);
nand U2036 (N_2036,In_1718,In_1767);
nor U2037 (N_2037,In_617,In_31);
and U2038 (N_2038,In_821,In_1250);
nor U2039 (N_2039,In_1877,In_1095);
nand U2040 (N_2040,In_2018,In_1593);
nor U2041 (N_2041,In_1690,In_939);
and U2042 (N_2042,In_944,In_1047);
nor U2043 (N_2043,In_2210,In_1658);
and U2044 (N_2044,In_505,In_2214);
nand U2045 (N_2045,In_515,In_1479);
and U2046 (N_2046,In_1896,In_1213);
nand U2047 (N_2047,In_1962,In_14);
nand U2048 (N_2048,In_1072,In_1329);
nand U2049 (N_2049,In_1655,In_1952);
nor U2050 (N_2050,In_2498,In_2143);
and U2051 (N_2051,In_34,In_1945);
xor U2052 (N_2052,In_1328,In_1704);
nor U2053 (N_2053,In_1539,In_2119);
or U2054 (N_2054,In_2183,In_1856);
or U2055 (N_2055,In_229,In_1431);
xor U2056 (N_2056,In_1865,In_2013);
or U2057 (N_2057,In_1994,In_1850);
nand U2058 (N_2058,In_2223,In_756);
nor U2059 (N_2059,In_296,In_937);
nand U2060 (N_2060,In_152,In_2484);
nand U2061 (N_2061,In_1685,In_344);
or U2062 (N_2062,In_1438,In_1395);
xor U2063 (N_2063,In_1387,In_2270);
or U2064 (N_2064,In_1955,In_166);
or U2065 (N_2065,In_2420,In_1755);
nand U2066 (N_2066,In_1604,In_1374);
and U2067 (N_2067,In_478,In_168);
nor U2068 (N_2068,In_2177,In_2155);
nand U2069 (N_2069,In_818,In_90);
or U2070 (N_2070,In_776,In_1896);
nor U2071 (N_2071,In_1362,In_694);
nor U2072 (N_2072,In_2036,In_1372);
or U2073 (N_2073,In_1780,In_2383);
nor U2074 (N_2074,In_10,In_920);
or U2075 (N_2075,In_1972,In_226);
and U2076 (N_2076,In_2432,In_2479);
nand U2077 (N_2077,In_2136,In_2230);
xnor U2078 (N_2078,In_2232,In_2482);
and U2079 (N_2079,In_830,In_2058);
nand U2080 (N_2080,In_1353,In_2491);
nand U2081 (N_2081,In_1889,In_144);
or U2082 (N_2082,In_2198,In_575);
nand U2083 (N_2083,In_995,In_1136);
nor U2084 (N_2084,In_180,In_820);
and U2085 (N_2085,In_270,In_2455);
nand U2086 (N_2086,In_1491,In_234);
or U2087 (N_2087,In_2020,In_2260);
nand U2088 (N_2088,In_484,In_1076);
and U2089 (N_2089,In_5,In_1148);
and U2090 (N_2090,In_398,In_818);
and U2091 (N_2091,In_959,In_561);
nor U2092 (N_2092,In_240,In_954);
and U2093 (N_2093,In_2436,In_647);
and U2094 (N_2094,In_2067,In_26);
nor U2095 (N_2095,In_1286,In_2306);
or U2096 (N_2096,In_817,In_1085);
and U2097 (N_2097,In_1251,In_2040);
nor U2098 (N_2098,In_1432,In_152);
nand U2099 (N_2099,In_39,In_1378);
and U2100 (N_2100,In_201,In_922);
xnor U2101 (N_2101,In_852,In_84);
and U2102 (N_2102,In_1754,In_1134);
nand U2103 (N_2103,In_2081,In_2214);
nand U2104 (N_2104,In_591,In_1681);
or U2105 (N_2105,In_1614,In_1507);
or U2106 (N_2106,In_1397,In_19);
or U2107 (N_2107,In_828,In_320);
and U2108 (N_2108,In_1368,In_962);
and U2109 (N_2109,In_1835,In_1453);
or U2110 (N_2110,In_1142,In_2014);
or U2111 (N_2111,In_1188,In_495);
nand U2112 (N_2112,In_902,In_1717);
nand U2113 (N_2113,In_800,In_604);
or U2114 (N_2114,In_2177,In_2015);
or U2115 (N_2115,In_2014,In_2340);
nor U2116 (N_2116,In_2399,In_2448);
nor U2117 (N_2117,In_1675,In_1149);
or U2118 (N_2118,In_1138,In_1218);
or U2119 (N_2119,In_668,In_833);
or U2120 (N_2120,In_695,In_906);
and U2121 (N_2121,In_1189,In_2389);
nand U2122 (N_2122,In_392,In_2075);
nor U2123 (N_2123,In_480,In_813);
nor U2124 (N_2124,In_1156,In_729);
nor U2125 (N_2125,In_1955,In_1061);
xnor U2126 (N_2126,In_2471,In_2351);
and U2127 (N_2127,In_507,In_1585);
nor U2128 (N_2128,In_2127,In_2463);
nand U2129 (N_2129,In_63,In_1429);
and U2130 (N_2130,In_2213,In_1265);
and U2131 (N_2131,In_1301,In_1511);
nor U2132 (N_2132,In_1147,In_2325);
xnor U2133 (N_2133,In_137,In_2284);
nor U2134 (N_2134,In_2140,In_984);
nor U2135 (N_2135,In_244,In_1164);
nand U2136 (N_2136,In_477,In_2484);
and U2137 (N_2137,In_650,In_836);
xnor U2138 (N_2138,In_2410,In_729);
or U2139 (N_2139,In_262,In_79);
nor U2140 (N_2140,In_1846,In_371);
and U2141 (N_2141,In_2318,In_817);
xor U2142 (N_2142,In_820,In_1889);
and U2143 (N_2143,In_1464,In_1843);
nor U2144 (N_2144,In_1669,In_948);
xor U2145 (N_2145,In_1952,In_1112);
or U2146 (N_2146,In_1939,In_358);
nor U2147 (N_2147,In_1329,In_43);
nor U2148 (N_2148,In_2215,In_1730);
nand U2149 (N_2149,In_619,In_64);
and U2150 (N_2150,In_2396,In_1318);
nor U2151 (N_2151,In_1356,In_870);
nor U2152 (N_2152,In_289,In_113);
and U2153 (N_2153,In_1131,In_1728);
and U2154 (N_2154,In_1790,In_725);
nor U2155 (N_2155,In_2330,In_275);
xnor U2156 (N_2156,In_490,In_403);
nand U2157 (N_2157,In_1341,In_1191);
or U2158 (N_2158,In_1201,In_1426);
or U2159 (N_2159,In_1697,In_729);
and U2160 (N_2160,In_688,In_730);
nand U2161 (N_2161,In_1622,In_2240);
nand U2162 (N_2162,In_271,In_614);
nand U2163 (N_2163,In_1550,In_1771);
or U2164 (N_2164,In_1447,In_885);
nor U2165 (N_2165,In_2289,In_1803);
or U2166 (N_2166,In_917,In_466);
nand U2167 (N_2167,In_223,In_526);
or U2168 (N_2168,In_2463,In_747);
or U2169 (N_2169,In_2137,In_2222);
nand U2170 (N_2170,In_1346,In_754);
nor U2171 (N_2171,In_1940,In_701);
nand U2172 (N_2172,In_41,In_1971);
xnor U2173 (N_2173,In_1944,In_1054);
and U2174 (N_2174,In_2002,In_2091);
nand U2175 (N_2175,In_2008,In_1888);
nand U2176 (N_2176,In_1003,In_1310);
nand U2177 (N_2177,In_1112,In_781);
and U2178 (N_2178,In_165,In_248);
and U2179 (N_2179,In_1187,In_1381);
and U2180 (N_2180,In_564,In_1789);
or U2181 (N_2181,In_2358,In_2473);
xnor U2182 (N_2182,In_1692,In_434);
nor U2183 (N_2183,In_755,In_1735);
and U2184 (N_2184,In_1374,In_1582);
nor U2185 (N_2185,In_2074,In_1983);
or U2186 (N_2186,In_2131,In_2265);
xor U2187 (N_2187,In_154,In_530);
xnor U2188 (N_2188,In_643,In_1070);
or U2189 (N_2189,In_369,In_538);
and U2190 (N_2190,In_16,In_493);
xnor U2191 (N_2191,In_2444,In_669);
or U2192 (N_2192,In_1258,In_1751);
nor U2193 (N_2193,In_660,In_3);
nor U2194 (N_2194,In_314,In_2064);
nand U2195 (N_2195,In_1289,In_1848);
nand U2196 (N_2196,In_47,In_1516);
or U2197 (N_2197,In_963,In_2264);
nand U2198 (N_2198,In_781,In_240);
and U2199 (N_2199,In_1198,In_262);
and U2200 (N_2200,In_339,In_2008);
nor U2201 (N_2201,In_1045,In_1109);
nand U2202 (N_2202,In_1055,In_1424);
or U2203 (N_2203,In_278,In_1869);
or U2204 (N_2204,In_833,In_1968);
or U2205 (N_2205,In_1891,In_373);
nor U2206 (N_2206,In_1839,In_1025);
nand U2207 (N_2207,In_211,In_935);
nor U2208 (N_2208,In_1631,In_2133);
xor U2209 (N_2209,In_276,In_1374);
nor U2210 (N_2210,In_1044,In_463);
or U2211 (N_2211,In_2342,In_1988);
and U2212 (N_2212,In_94,In_1892);
or U2213 (N_2213,In_1102,In_1360);
nor U2214 (N_2214,In_1640,In_1853);
nand U2215 (N_2215,In_1750,In_29);
and U2216 (N_2216,In_557,In_210);
nor U2217 (N_2217,In_1905,In_475);
nor U2218 (N_2218,In_218,In_519);
nor U2219 (N_2219,In_1037,In_19);
or U2220 (N_2220,In_1856,In_1728);
and U2221 (N_2221,In_420,In_1039);
nand U2222 (N_2222,In_2317,In_556);
and U2223 (N_2223,In_219,In_18);
or U2224 (N_2224,In_1767,In_952);
and U2225 (N_2225,In_785,In_2431);
nand U2226 (N_2226,In_1146,In_2293);
nor U2227 (N_2227,In_1596,In_738);
and U2228 (N_2228,In_560,In_1158);
nor U2229 (N_2229,In_1117,In_1558);
or U2230 (N_2230,In_1671,In_738);
nand U2231 (N_2231,In_1520,In_291);
and U2232 (N_2232,In_470,In_985);
or U2233 (N_2233,In_2498,In_1974);
nand U2234 (N_2234,In_1554,In_717);
or U2235 (N_2235,In_977,In_1234);
nor U2236 (N_2236,In_967,In_1935);
xor U2237 (N_2237,In_1367,In_422);
or U2238 (N_2238,In_418,In_537);
or U2239 (N_2239,In_990,In_868);
or U2240 (N_2240,In_2060,In_2262);
xor U2241 (N_2241,In_1161,In_831);
and U2242 (N_2242,In_1259,In_1321);
nand U2243 (N_2243,In_1304,In_1156);
nor U2244 (N_2244,In_935,In_2135);
xnor U2245 (N_2245,In_349,In_1554);
nor U2246 (N_2246,In_2161,In_2265);
xnor U2247 (N_2247,In_220,In_2118);
nand U2248 (N_2248,In_914,In_1654);
nor U2249 (N_2249,In_1187,In_2087);
nand U2250 (N_2250,In_879,In_649);
and U2251 (N_2251,In_1945,In_2305);
nor U2252 (N_2252,In_1401,In_1194);
nor U2253 (N_2253,In_1286,In_1212);
nor U2254 (N_2254,In_1586,In_1340);
or U2255 (N_2255,In_1442,In_848);
nor U2256 (N_2256,In_1018,In_373);
or U2257 (N_2257,In_1474,In_77);
xnor U2258 (N_2258,In_1464,In_248);
nor U2259 (N_2259,In_587,In_778);
xor U2260 (N_2260,In_2005,In_1107);
or U2261 (N_2261,In_593,In_1311);
and U2262 (N_2262,In_1682,In_724);
or U2263 (N_2263,In_927,In_116);
or U2264 (N_2264,In_1416,In_1299);
or U2265 (N_2265,In_2218,In_2021);
nor U2266 (N_2266,In_1581,In_519);
nand U2267 (N_2267,In_851,In_794);
and U2268 (N_2268,In_1412,In_1713);
or U2269 (N_2269,In_1472,In_735);
nor U2270 (N_2270,In_1027,In_415);
nand U2271 (N_2271,In_2118,In_1578);
nor U2272 (N_2272,In_1903,In_1808);
nor U2273 (N_2273,In_1118,In_1732);
nand U2274 (N_2274,In_910,In_726);
nand U2275 (N_2275,In_1791,In_1316);
nor U2276 (N_2276,In_1075,In_2489);
or U2277 (N_2277,In_571,In_849);
nand U2278 (N_2278,In_1118,In_1830);
or U2279 (N_2279,In_840,In_2046);
nor U2280 (N_2280,In_1874,In_1367);
or U2281 (N_2281,In_1322,In_275);
xnor U2282 (N_2282,In_369,In_1728);
nor U2283 (N_2283,In_63,In_1050);
nor U2284 (N_2284,In_1798,In_2399);
nor U2285 (N_2285,In_1766,In_1963);
and U2286 (N_2286,In_2313,In_1053);
and U2287 (N_2287,In_2418,In_1877);
or U2288 (N_2288,In_573,In_886);
and U2289 (N_2289,In_1428,In_1972);
nor U2290 (N_2290,In_757,In_60);
nor U2291 (N_2291,In_546,In_2038);
nor U2292 (N_2292,In_895,In_2183);
nand U2293 (N_2293,In_1389,In_389);
nand U2294 (N_2294,In_1866,In_2035);
nor U2295 (N_2295,In_2457,In_2313);
nor U2296 (N_2296,In_2349,In_214);
and U2297 (N_2297,In_1384,In_238);
and U2298 (N_2298,In_1555,In_1946);
and U2299 (N_2299,In_986,In_1304);
and U2300 (N_2300,In_1950,In_0);
or U2301 (N_2301,In_1890,In_797);
nor U2302 (N_2302,In_407,In_1427);
and U2303 (N_2303,In_42,In_1777);
or U2304 (N_2304,In_2373,In_1815);
or U2305 (N_2305,In_1731,In_2261);
and U2306 (N_2306,In_1043,In_1828);
and U2307 (N_2307,In_1419,In_2337);
or U2308 (N_2308,In_1328,In_1727);
or U2309 (N_2309,In_1396,In_1552);
nor U2310 (N_2310,In_2345,In_947);
and U2311 (N_2311,In_1643,In_1880);
or U2312 (N_2312,In_698,In_121);
nor U2313 (N_2313,In_69,In_1253);
nand U2314 (N_2314,In_1708,In_1799);
nand U2315 (N_2315,In_1024,In_1053);
and U2316 (N_2316,In_1734,In_667);
and U2317 (N_2317,In_368,In_106);
and U2318 (N_2318,In_765,In_676);
and U2319 (N_2319,In_1739,In_96);
and U2320 (N_2320,In_1614,In_2469);
nor U2321 (N_2321,In_382,In_2401);
nor U2322 (N_2322,In_770,In_2313);
or U2323 (N_2323,In_594,In_605);
or U2324 (N_2324,In_1915,In_2225);
xnor U2325 (N_2325,In_655,In_1840);
nor U2326 (N_2326,In_2289,In_795);
nand U2327 (N_2327,In_1404,In_1365);
nand U2328 (N_2328,In_1890,In_163);
nand U2329 (N_2329,In_310,In_1837);
xnor U2330 (N_2330,In_452,In_439);
or U2331 (N_2331,In_1859,In_2128);
or U2332 (N_2332,In_1834,In_1599);
nand U2333 (N_2333,In_657,In_2186);
nand U2334 (N_2334,In_2073,In_1498);
and U2335 (N_2335,In_901,In_1375);
nand U2336 (N_2336,In_1534,In_2440);
nor U2337 (N_2337,In_1595,In_287);
or U2338 (N_2338,In_1891,In_909);
and U2339 (N_2339,In_1503,In_1394);
nor U2340 (N_2340,In_2069,In_1008);
or U2341 (N_2341,In_2420,In_909);
xnor U2342 (N_2342,In_379,In_1257);
nor U2343 (N_2343,In_215,In_591);
or U2344 (N_2344,In_651,In_2075);
and U2345 (N_2345,In_1994,In_922);
nand U2346 (N_2346,In_1085,In_1089);
or U2347 (N_2347,In_892,In_292);
or U2348 (N_2348,In_1027,In_494);
and U2349 (N_2349,In_757,In_2102);
or U2350 (N_2350,In_1170,In_507);
nand U2351 (N_2351,In_2065,In_672);
and U2352 (N_2352,In_981,In_2263);
or U2353 (N_2353,In_606,In_411);
nor U2354 (N_2354,In_1170,In_1843);
or U2355 (N_2355,In_2452,In_219);
and U2356 (N_2356,In_1100,In_1556);
and U2357 (N_2357,In_574,In_741);
and U2358 (N_2358,In_2297,In_797);
nor U2359 (N_2359,In_1233,In_1746);
nor U2360 (N_2360,In_935,In_1244);
xor U2361 (N_2361,In_690,In_256);
and U2362 (N_2362,In_2490,In_2498);
nor U2363 (N_2363,In_1474,In_542);
nand U2364 (N_2364,In_570,In_411);
xnor U2365 (N_2365,In_2247,In_220);
and U2366 (N_2366,In_1018,In_813);
and U2367 (N_2367,In_302,In_261);
nand U2368 (N_2368,In_1868,In_884);
nand U2369 (N_2369,In_864,In_2464);
nand U2370 (N_2370,In_1492,In_1625);
nor U2371 (N_2371,In_1236,In_679);
or U2372 (N_2372,In_1515,In_58);
or U2373 (N_2373,In_1101,In_2362);
nor U2374 (N_2374,In_2081,In_498);
nor U2375 (N_2375,In_29,In_862);
or U2376 (N_2376,In_2433,In_276);
or U2377 (N_2377,In_1063,In_2404);
and U2378 (N_2378,In_1195,In_920);
nor U2379 (N_2379,In_2208,In_721);
nand U2380 (N_2380,In_104,In_1224);
and U2381 (N_2381,In_1431,In_1040);
and U2382 (N_2382,In_1229,In_693);
nand U2383 (N_2383,In_110,In_308);
and U2384 (N_2384,In_1896,In_2203);
and U2385 (N_2385,In_1329,In_636);
xor U2386 (N_2386,In_426,In_540);
or U2387 (N_2387,In_437,In_1986);
xor U2388 (N_2388,In_569,In_1732);
and U2389 (N_2389,In_100,In_664);
nor U2390 (N_2390,In_1229,In_1769);
nand U2391 (N_2391,In_1253,In_942);
and U2392 (N_2392,In_2304,In_1859);
and U2393 (N_2393,In_1904,In_2318);
and U2394 (N_2394,In_1225,In_183);
or U2395 (N_2395,In_2393,In_1849);
nand U2396 (N_2396,In_872,In_178);
or U2397 (N_2397,In_2182,In_1042);
and U2398 (N_2398,In_441,In_1361);
or U2399 (N_2399,In_454,In_1124);
or U2400 (N_2400,In_483,In_746);
nor U2401 (N_2401,In_44,In_1703);
xnor U2402 (N_2402,In_1486,In_1645);
nor U2403 (N_2403,In_987,In_1284);
nor U2404 (N_2404,In_1535,In_688);
and U2405 (N_2405,In_1324,In_1819);
nand U2406 (N_2406,In_2281,In_1417);
and U2407 (N_2407,In_243,In_1999);
and U2408 (N_2408,In_713,In_2344);
xor U2409 (N_2409,In_1661,In_454);
or U2410 (N_2410,In_1668,In_756);
nand U2411 (N_2411,In_549,In_452);
nor U2412 (N_2412,In_2181,In_1304);
nand U2413 (N_2413,In_856,In_184);
and U2414 (N_2414,In_1944,In_895);
nor U2415 (N_2415,In_2084,In_572);
or U2416 (N_2416,In_1398,In_1409);
nand U2417 (N_2417,In_2372,In_345);
nand U2418 (N_2418,In_1345,In_1007);
or U2419 (N_2419,In_1728,In_424);
xnor U2420 (N_2420,In_200,In_1800);
or U2421 (N_2421,In_1652,In_1989);
xnor U2422 (N_2422,In_651,In_2448);
nand U2423 (N_2423,In_2421,In_1715);
or U2424 (N_2424,In_27,In_252);
or U2425 (N_2425,In_771,In_2017);
and U2426 (N_2426,In_1653,In_660);
xor U2427 (N_2427,In_1042,In_1032);
nor U2428 (N_2428,In_541,In_1021);
nand U2429 (N_2429,In_912,In_1346);
nor U2430 (N_2430,In_509,In_468);
and U2431 (N_2431,In_14,In_2422);
and U2432 (N_2432,In_1931,In_31);
and U2433 (N_2433,In_1681,In_991);
or U2434 (N_2434,In_1095,In_1220);
or U2435 (N_2435,In_132,In_138);
nor U2436 (N_2436,In_595,In_765);
nor U2437 (N_2437,In_1994,In_1869);
and U2438 (N_2438,In_2484,In_481);
xnor U2439 (N_2439,In_1715,In_1408);
nand U2440 (N_2440,In_2303,In_1455);
xnor U2441 (N_2441,In_1112,In_1912);
or U2442 (N_2442,In_543,In_2141);
nand U2443 (N_2443,In_1067,In_1250);
nand U2444 (N_2444,In_1644,In_1197);
or U2445 (N_2445,In_1831,In_1643);
and U2446 (N_2446,In_1482,In_2035);
nor U2447 (N_2447,In_1027,In_1660);
nand U2448 (N_2448,In_2028,In_1283);
nor U2449 (N_2449,In_1883,In_2292);
and U2450 (N_2450,In_93,In_516);
nor U2451 (N_2451,In_1842,In_1237);
nand U2452 (N_2452,In_687,In_2391);
or U2453 (N_2453,In_2494,In_764);
nand U2454 (N_2454,In_295,In_2388);
nand U2455 (N_2455,In_916,In_1262);
nand U2456 (N_2456,In_1693,In_1610);
nand U2457 (N_2457,In_66,In_295);
nand U2458 (N_2458,In_1371,In_507);
or U2459 (N_2459,In_650,In_1014);
and U2460 (N_2460,In_1325,In_29);
nand U2461 (N_2461,In_2312,In_2091);
or U2462 (N_2462,In_2230,In_757);
nor U2463 (N_2463,In_1746,In_1295);
or U2464 (N_2464,In_1658,In_714);
and U2465 (N_2465,In_376,In_1345);
and U2466 (N_2466,In_2273,In_1874);
xor U2467 (N_2467,In_2198,In_1782);
nand U2468 (N_2468,In_294,In_2343);
or U2469 (N_2469,In_1344,In_467);
nand U2470 (N_2470,In_443,In_446);
xor U2471 (N_2471,In_2249,In_289);
nand U2472 (N_2472,In_1111,In_633);
and U2473 (N_2473,In_1901,In_1362);
or U2474 (N_2474,In_650,In_392);
xor U2475 (N_2475,In_2383,In_1216);
or U2476 (N_2476,In_762,In_915);
nand U2477 (N_2477,In_220,In_2369);
nand U2478 (N_2478,In_44,In_1514);
nor U2479 (N_2479,In_2250,In_107);
nor U2480 (N_2480,In_863,In_1281);
and U2481 (N_2481,In_1531,In_1500);
nand U2482 (N_2482,In_913,In_964);
nor U2483 (N_2483,In_838,In_1925);
xor U2484 (N_2484,In_674,In_382);
and U2485 (N_2485,In_1392,In_797);
or U2486 (N_2486,In_1463,In_1980);
and U2487 (N_2487,In_1785,In_77);
and U2488 (N_2488,In_139,In_1322);
or U2489 (N_2489,In_2261,In_2320);
and U2490 (N_2490,In_2416,In_1324);
and U2491 (N_2491,In_1972,In_1118);
and U2492 (N_2492,In_1987,In_2278);
and U2493 (N_2493,In_1780,In_1858);
or U2494 (N_2494,In_664,In_2136);
nor U2495 (N_2495,In_1,In_1999);
nand U2496 (N_2496,In_1585,In_537);
nand U2497 (N_2497,In_275,In_2244);
or U2498 (N_2498,In_1443,In_421);
or U2499 (N_2499,In_1550,In_1188);
or U2500 (N_2500,In_792,In_2376);
nor U2501 (N_2501,In_2122,In_212);
and U2502 (N_2502,In_2138,In_11);
nor U2503 (N_2503,In_1953,In_1378);
or U2504 (N_2504,In_2286,In_599);
nand U2505 (N_2505,In_1196,In_959);
nor U2506 (N_2506,In_252,In_1030);
nor U2507 (N_2507,In_333,In_2322);
nor U2508 (N_2508,In_365,In_2194);
or U2509 (N_2509,In_1212,In_1135);
nand U2510 (N_2510,In_1129,In_1351);
nor U2511 (N_2511,In_1061,In_2426);
xnor U2512 (N_2512,In_1579,In_1012);
or U2513 (N_2513,In_135,In_1176);
nand U2514 (N_2514,In_2396,In_386);
or U2515 (N_2515,In_1228,In_68);
xor U2516 (N_2516,In_1967,In_2319);
nand U2517 (N_2517,In_360,In_528);
or U2518 (N_2518,In_1028,In_1304);
nand U2519 (N_2519,In_170,In_1433);
and U2520 (N_2520,In_588,In_1645);
nor U2521 (N_2521,In_624,In_708);
xnor U2522 (N_2522,In_1917,In_2451);
nor U2523 (N_2523,In_962,In_181);
and U2524 (N_2524,In_474,In_1973);
and U2525 (N_2525,In_124,In_2335);
nor U2526 (N_2526,In_438,In_208);
and U2527 (N_2527,In_2331,In_569);
and U2528 (N_2528,In_248,In_818);
xnor U2529 (N_2529,In_723,In_520);
nor U2530 (N_2530,In_2415,In_1095);
xor U2531 (N_2531,In_486,In_536);
nor U2532 (N_2532,In_1477,In_2250);
or U2533 (N_2533,In_1677,In_2174);
xnor U2534 (N_2534,In_1126,In_1972);
and U2535 (N_2535,In_2183,In_1556);
xnor U2536 (N_2536,In_105,In_37);
and U2537 (N_2537,In_1221,In_1961);
nand U2538 (N_2538,In_1606,In_1798);
or U2539 (N_2539,In_847,In_2464);
nor U2540 (N_2540,In_2480,In_1858);
nor U2541 (N_2541,In_243,In_26);
or U2542 (N_2542,In_2241,In_1036);
or U2543 (N_2543,In_1603,In_1565);
nor U2544 (N_2544,In_879,In_1607);
or U2545 (N_2545,In_191,In_831);
xor U2546 (N_2546,In_1004,In_216);
and U2547 (N_2547,In_1463,In_1679);
nor U2548 (N_2548,In_2360,In_57);
nand U2549 (N_2549,In_786,In_1972);
nor U2550 (N_2550,In_1252,In_1263);
nor U2551 (N_2551,In_1690,In_1505);
nand U2552 (N_2552,In_1691,In_508);
xor U2553 (N_2553,In_1756,In_983);
or U2554 (N_2554,In_997,In_1899);
nor U2555 (N_2555,In_2397,In_450);
or U2556 (N_2556,In_1300,In_361);
nand U2557 (N_2557,In_298,In_1418);
and U2558 (N_2558,In_850,In_103);
or U2559 (N_2559,In_854,In_28);
or U2560 (N_2560,In_418,In_273);
nand U2561 (N_2561,In_69,In_1472);
and U2562 (N_2562,In_878,In_1696);
and U2563 (N_2563,In_740,In_1327);
nor U2564 (N_2564,In_506,In_666);
and U2565 (N_2565,In_1268,In_1591);
xor U2566 (N_2566,In_593,In_1142);
or U2567 (N_2567,In_2319,In_416);
xnor U2568 (N_2568,In_1594,In_1794);
xnor U2569 (N_2569,In_1386,In_2185);
or U2570 (N_2570,In_2436,In_1961);
or U2571 (N_2571,In_2347,In_1983);
nand U2572 (N_2572,In_1144,In_403);
and U2573 (N_2573,In_1557,In_2374);
nor U2574 (N_2574,In_568,In_1618);
and U2575 (N_2575,In_1807,In_1583);
or U2576 (N_2576,In_381,In_1300);
nor U2577 (N_2577,In_1416,In_207);
nor U2578 (N_2578,In_2064,In_1519);
and U2579 (N_2579,In_836,In_607);
or U2580 (N_2580,In_893,In_1007);
and U2581 (N_2581,In_471,In_854);
nand U2582 (N_2582,In_2460,In_1441);
nand U2583 (N_2583,In_811,In_1210);
nor U2584 (N_2584,In_292,In_281);
and U2585 (N_2585,In_1141,In_1934);
or U2586 (N_2586,In_1878,In_1888);
or U2587 (N_2587,In_94,In_1214);
nand U2588 (N_2588,In_1235,In_135);
or U2589 (N_2589,In_1231,In_1003);
xnor U2590 (N_2590,In_2098,In_2318);
nor U2591 (N_2591,In_19,In_760);
nor U2592 (N_2592,In_1465,In_1115);
nand U2593 (N_2593,In_2100,In_323);
nand U2594 (N_2594,In_1633,In_1662);
or U2595 (N_2595,In_984,In_2261);
and U2596 (N_2596,In_232,In_1376);
nand U2597 (N_2597,In_61,In_1898);
and U2598 (N_2598,In_204,In_1623);
xor U2599 (N_2599,In_2102,In_739);
and U2600 (N_2600,In_429,In_697);
or U2601 (N_2601,In_1587,In_1444);
nand U2602 (N_2602,In_1680,In_2106);
and U2603 (N_2603,In_129,In_358);
nor U2604 (N_2604,In_1155,In_1554);
and U2605 (N_2605,In_2118,In_415);
nor U2606 (N_2606,In_1158,In_1056);
and U2607 (N_2607,In_2319,In_1683);
nand U2608 (N_2608,In_432,In_646);
and U2609 (N_2609,In_970,In_678);
xnor U2610 (N_2610,In_2439,In_2090);
nor U2611 (N_2611,In_1970,In_122);
nand U2612 (N_2612,In_2241,In_1987);
and U2613 (N_2613,In_971,In_1438);
or U2614 (N_2614,In_1591,In_1460);
and U2615 (N_2615,In_1010,In_1075);
nor U2616 (N_2616,In_270,In_1306);
and U2617 (N_2617,In_1582,In_910);
nand U2618 (N_2618,In_1892,In_2290);
nand U2619 (N_2619,In_1756,In_2208);
xnor U2620 (N_2620,In_737,In_1102);
nor U2621 (N_2621,In_401,In_566);
nand U2622 (N_2622,In_286,In_2254);
nand U2623 (N_2623,In_1818,In_695);
or U2624 (N_2624,In_1719,In_1826);
nand U2625 (N_2625,In_162,In_294);
xor U2626 (N_2626,In_1515,In_96);
and U2627 (N_2627,In_3,In_1867);
nand U2628 (N_2628,In_1204,In_1560);
nand U2629 (N_2629,In_337,In_1174);
and U2630 (N_2630,In_1304,In_2293);
nand U2631 (N_2631,In_2289,In_1279);
nand U2632 (N_2632,In_1883,In_828);
and U2633 (N_2633,In_2048,In_72);
and U2634 (N_2634,In_1962,In_1465);
or U2635 (N_2635,In_2156,In_1347);
or U2636 (N_2636,In_38,In_417);
nor U2637 (N_2637,In_344,In_362);
nand U2638 (N_2638,In_1804,In_852);
nand U2639 (N_2639,In_413,In_94);
nand U2640 (N_2640,In_1705,In_1479);
or U2641 (N_2641,In_688,In_198);
nor U2642 (N_2642,In_2323,In_837);
nor U2643 (N_2643,In_1947,In_1433);
nand U2644 (N_2644,In_1364,In_1712);
nand U2645 (N_2645,In_990,In_1076);
and U2646 (N_2646,In_900,In_2368);
and U2647 (N_2647,In_1585,In_443);
or U2648 (N_2648,In_805,In_562);
nor U2649 (N_2649,In_2184,In_1227);
or U2650 (N_2650,In_2247,In_2219);
nor U2651 (N_2651,In_351,In_1099);
xnor U2652 (N_2652,In_2382,In_853);
or U2653 (N_2653,In_1843,In_2259);
nand U2654 (N_2654,In_1599,In_1823);
and U2655 (N_2655,In_427,In_2136);
or U2656 (N_2656,In_373,In_724);
and U2657 (N_2657,In_902,In_197);
nor U2658 (N_2658,In_1313,In_669);
nor U2659 (N_2659,In_1775,In_699);
nor U2660 (N_2660,In_1583,In_1445);
nand U2661 (N_2661,In_195,In_1226);
or U2662 (N_2662,In_443,In_882);
or U2663 (N_2663,In_364,In_292);
nor U2664 (N_2664,In_479,In_917);
nor U2665 (N_2665,In_1427,In_1705);
nor U2666 (N_2666,In_1065,In_134);
nor U2667 (N_2667,In_964,In_1535);
and U2668 (N_2668,In_2412,In_20);
nand U2669 (N_2669,In_1155,In_1868);
and U2670 (N_2670,In_2086,In_2059);
or U2671 (N_2671,In_2437,In_2258);
or U2672 (N_2672,In_1596,In_2057);
xor U2673 (N_2673,In_2459,In_664);
nand U2674 (N_2674,In_1990,In_1445);
nand U2675 (N_2675,In_1189,In_1264);
nor U2676 (N_2676,In_1475,In_241);
nor U2677 (N_2677,In_1401,In_2087);
and U2678 (N_2678,In_4,In_2370);
xor U2679 (N_2679,In_1050,In_1400);
and U2680 (N_2680,In_1109,In_1489);
nor U2681 (N_2681,In_266,In_252);
and U2682 (N_2682,In_1495,In_1878);
nor U2683 (N_2683,In_1693,In_1948);
and U2684 (N_2684,In_287,In_1811);
nand U2685 (N_2685,In_766,In_2377);
or U2686 (N_2686,In_1427,In_1464);
nor U2687 (N_2687,In_205,In_1693);
nor U2688 (N_2688,In_369,In_526);
xor U2689 (N_2689,In_1213,In_1796);
nor U2690 (N_2690,In_2252,In_2025);
nor U2691 (N_2691,In_2366,In_2341);
or U2692 (N_2692,In_2421,In_683);
xnor U2693 (N_2693,In_1313,In_1249);
nand U2694 (N_2694,In_976,In_126);
nand U2695 (N_2695,In_2054,In_1646);
and U2696 (N_2696,In_1994,In_1640);
nor U2697 (N_2697,In_1906,In_2265);
and U2698 (N_2698,In_2137,In_1038);
xnor U2699 (N_2699,In_1554,In_2141);
or U2700 (N_2700,In_2285,In_466);
or U2701 (N_2701,In_446,In_907);
and U2702 (N_2702,In_1679,In_471);
nor U2703 (N_2703,In_2447,In_568);
or U2704 (N_2704,In_1742,In_246);
xnor U2705 (N_2705,In_741,In_1797);
xor U2706 (N_2706,In_436,In_1013);
or U2707 (N_2707,In_2038,In_1751);
xnor U2708 (N_2708,In_1161,In_2491);
nor U2709 (N_2709,In_2445,In_1133);
nand U2710 (N_2710,In_2146,In_373);
xnor U2711 (N_2711,In_1010,In_0);
and U2712 (N_2712,In_1166,In_2073);
or U2713 (N_2713,In_543,In_1408);
nor U2714 (N_2714,In_695,In_1766);
nor U2715 (N_2715,In_2091,In_1303);
and U2716 (N_2716,In_2450,In_777);
nand U2717 (N_2717,In_1179,In_1329);
or U2718 (N_2718,In_1993,In_401);
nor U2719 (N_2719,In_1035,In_1263);
and U2720 (N_2720,In_1062,In_2082);
or U2721 (N_2721,In_968,In_1011);
or U2722 (N_2722,In_1270,In_1355);
or U2723 (N_2723,In_1708,In_1509);
and U2724 (N_2724,In_183,In_870);
nand U2725 (N_2725,In_2493,In_1418);
and U2726 (N_2726,In_2186,In_1228);
and U2727 (N_2727,In_2272,In_2091);
or U2728 (N_2728,In_578,In_527);
nor U2729 (N_2729,In_1056,In_1067);
nor U2730 (N_2730,In_787,In_111);
and U2731 (N_2731,In_1562,In_636);
and U2732 (N_2732,In_2164,In_2426);
nand U2733 (N_2733,In_2167,In_39);
nand U2734 (N_2734,In_2403,In_2388);
nand U2735 (N_2735,In_654,In_1442);
or U2736 (N_2736,In_1819,In_275);
nor U2737 (N_2737,In_146,In_2487);
and U2738 (N_2738,In_1787,In_1090);
or U2739 (N_2739,In_1178,In_1370);
or U2740 (N_2740,In_1745,In_1140);
or U2741 (N_2741,In_2079,In_1484);
or U2742 (N_2742,In_1257,In_1674);
nand U2743 (N_2743,In_1873,In_2410);
and U2744 (N_2744,In_1486,In_893);
and U2745 (N_2745,In_1403,In_215);
and U2746 (N_2746,In_1291,In_2401);
nor U2747 (N_2747,In_1057,In_1912);
or U2748 (N_2748,In_302,In_788);
nor U2749 (N_2749,In_1285,In_2372);
or U2750 (N_2750,In_107,In_1464);
or U2751 (N_2751,In_2127,In_71);
nand U2752 (N_2752,In_995,In_325);
nand U2753 (N_2753,In_1029,In_1100);
nor U2754 (N_2754,In_86,In_597);
nand U2755 (N_2755,In_214,In_2076);
or U2756 (N_2756,In_331,In_1275);
and U2757 (N_2757,In_1801,In_95);
and U2758 (N_2758,In_837,In_259);
nor U2759 (N_2759,In_1020,In_1696);
nor U2760 (N_2760,In_1852,In_786);
or U2761 (N_2761,In_522,In_724);
nand U2762 (N_2762,In_316,In_1117);
xnor U2763 (N_2763,In_1336,In_728);
nand U2764 (N_2764,In_1958,In_685);
nor U2765 (N_2765,In_1362,In_2094);
nor U2766 (N_2766,In_1065,In_65);
and U2767 (N_2767,In_981,In_2335);
xnor U2768 (N_2768,In_2313,In_1778);
or U2769 (N_2769,In_1524,In_1443);
xnor U2770 (N_2770,In_2459,In_169);
and U2771 (N_2771,In_247,In_221);
nor U2772 (N_2772,In_204,In_854);
or U2773 (N_2773,In_1449,In_1290);
or U2774 (N_2774,In_2157,In_198);
and U2775 (N_2775,In_255,In_445);
xnor U2776 (N_2776,In_1755,In_2364);
and U2777 (N_2777,In_2281,In_550);
or U2778 (N_2778,In_2418,In_837);
and U2779 (N_2779,In_2315,In_2471);
xor U2780 (N_2780,In_256,In_255);
or U2781 (N_2781,In_145,In_1778);
and U2782 (N_2782,In_309,In_1587);
or U2783 (N_2783,In_1780,In_2484);
or U2784 (N_2784,In_1549,In_2364);
or U2785 (N_2785,In_2372,In_1925);
xor U2786 (N_2786,In_549,In_609);
and U2787 (N_2787,In_1127,In_802);
nand U2788 (N_2788,In_854,In_2451);
nor U2789 (N_2789,In_1275,In_123);
nand U2790 (N_2790,In_1720,In_1619);
nor U2791 (N_2791,In_1218,In_115);
nand U2792 (N_2792,In_1862,In_2477);
or U2793 (N_2793,In_2299,In_1729);
and U2794 (N_2794,In_448,In_1131);
and U2795 (N_2795,In_677,In_2211);
and U2796 (N_2796,In_10,In_1097);
and U2797 (N_2797,In_1622,In_1641);
and U2798 (N_2798,In_1525,In_550);
nor U2799 (N_2799,In_942,In_1259);
or U2800 (N_2800,In_1542,In_64);
or U2801 (N_2801,In_168,In_989);
and U2802 (N_2802,In_1916,In_1470);
nand U2803 (N_2803,In_1122,In_1379);
nor U2804 (N_2804,In_2020,In_908);
nor U2805 (N_2805,In_298,In_926);
or U2806 (N_2806,In_1783,In_627);
nand U2807 (N_2807,In_734,In_179);
nor U2808 (N_2808,In_2001,In_344);
xor U2809 (N_2809,In_2051,In_671);
nor U2810 (N_2810,In_1798,In_1535);
nand U2811 (N_2811,In_381,In_1439);
and U2812 (N_2812,In_1395,In_224);
or U2813 (N_2813,In_545,In_1447);
nor U2814 (N_2814,In_2330,In_1663);
and U2815 (N_2815,In_1459,In_1953);
nand U2816 (N_2816,In_2231,In_793);
and U2817 (N_2817,In_348,In_746);
and U2818 (N_2818,In_348,In_893);
and U2819 (N_2819,In_1854,In_95);
nor U2820 (N_2820,In_2290,In_1035);
xnor U2821 (N_2821,In_1599,In_187);
nand U2822 (N_2822,In_2384,In_2141);
nor U2823 (N_2823,In_746,In_1105);
and U2824 (N_2824,In_693,In_365);
nand U2825 (N_2825,In_1484,In_2037);
nand U2826 (N_2826,In_25,In_507);
nor U2827 (N_2827,In_2252,In_1680);
and U2828 (N_2828,In_866,In_1159);
and U2829 (N_2829,In_1922,In_1007);
or U2830 (N_2830,In_1242,In_1246);
nand U2831 (N_2831,In_758,In_1092);
nor U2832 (N_2832,In_2063,In_2474);
nor U2833 (N_2833,In_999,In_1251);
or U2834 (N_2834,In_2059,In_2178);
xor U2835 (N_2835,In_1381,In_1809);
nand U2836 (N_2836,In_1352,In_1110);
nor U2837 (N_2837,In_435,In_161);
nand U2838 (N_2838,In_2409,In_2273);
or U2839 (N_2839,In_887,In_1590);
nor U2840 (N_2840,In_845,In_1946);
nand U2841 (N_2841,In_781,In_412);
nor U2842 (N_2842,In_2417,In_726);
or U2843 (N_2843,In_2209,In_964);
or U2844 (N_2844,In_913,In_1533);
nand U2845 (N_2845,In_812,In_1765);
nand U2846 (N_2846,In_2362,In_2300);
or U2847 (N_2847,In_450,In_1564);
nand U2848 (N_2848,In_57,In_1041);
nor U2849 (N_2849,In_1355,In_798);
nand U2850 (N_2850,In_327,In_1021);
nand U2851 (N_2851,In_698,In_1030);
or U2852 (N_2852,In_264,In_572);
and U2853 (N_2853,In_2171,In_100);
xor U2854 (N_2854,In_573,In_1152);
nor U2855 (N_2855,In_1791,In_574);
nand U2856 (N_2856,In_1682,In_280);
and U2857 (N_2857,In_310,In_2110);
nor U2858 (N_2858,In_1776,In_2235);
or U2859 (N_2859,In_2196,In_1770);
or U2860 (N_2860,In_1966,In_1677);
nand U2861 (N_2861,In_1839,In_2016);
nor U2862 (N_2862,In_1731,In_1853);
nand U2863 (N_2863,In_980,In_1443);
or U2864 (N_2864,In_284,In_1094);
xor U2865 (N_2865,In_858,In_1917);
or U2866 (N_2866,In_2277,In_1310);
nand U2867 (N_2867,In_1379,In_112);
or U2868 (N_2868,In_2464,In_115);
xor U2869 (N_2869,In_1745,In_317);
nor U2870 (N_2870,In_1056,In_181);
or U2871 (N_2871,In_2324,In_541);
or U2872 (N_2872,In_1688,In_1399);
nor U2873 (N_2873,In_940,In_2338);
and U2874 (N_2874,In_1147,In_1996);
nor U2875 (N_2875,In_286,In_1278);
and U2876 (N_2876,In_2405,In_1747);
nand U2877 (N_2877,In_1484,In_986);
nor U2878 (N_2878,In_1928,In_885);
and U2879 (N_2879,In_816,In_701);
and U2880 (N_2880,In_299,In_280);
nor U2881 (N_2881,In_530,In_461);
nor U2882 (N_2882,In_17,In_1738);
xor U2883 (N_2883,In_1928,In_911);
nor U2884 (N_2884,In_1221,In_678);
nor U2885 (N_2885,In_2256,In_531);
nand U2886 (N_2886,In_304,In_689);
or U2887 (N_2887,In_2332,In_862);
or U2888 (N_2888,In_94,In_1472);
and U2889 (N_2889,In_2150,In_382);
and U2890 (N_2890,In_2125,In_83);
nand U2891 (N_2891,In_294,In_589);
and U2892 (N_2892,In_1070,In_187);
and U2893 (N_2893,In_404,In_2171);
nor U2894 (N_2894,In_1750,In_1063);
or U2895 (N_2895,In_2008,In_1610);
and U2896 (N_2896,In_927,In_1088);
and U2897 (N_2897,In_2077,In_2425);
or U2898 (N_2898,In_1823,In_336);
nor U2899 (N_2899,In_2048,In_417);
or U2900 (N_2900,In_1488,In_1054);
or U2901 (N_2901,In_1431,In_2260);
nor U2902 (N_2902,In_1467,In_683);
or U2903 (N_2903,In_234,In_1700);
nor U2904 (N_2904,In_1024,In_2479);
or U2905 (N_2905,In_800,In_2278);
nand U2906 (N_2906,In_1091,In_1060);
nand U2907 (N_2907,In_2105,In_2375);
xor U2908 (N_2908,In_397,In_2351);
nand U2909 (N_2909,In_226,In_1225);
nor U2910 (N_2910,In_1077,In_1046);
nor U2911 (N_2911,In_142,In_2040);
nand U2912 (N_2912,In_2158,In_1954);
nand U2913 (N_2913,In_1174,In_2122);
nor U2914 (N_2914,In_1010,In_1427);
and U2915 (N_2915,In_397,In_1759);
or U2916 (N_2916,In_287,In_2392);
and U2917 (N_2917,In_887,In_339);
nand U2918 (N_2918,In_1695,In_1503);
nor U2919 (N_2919,In_2072,In_565);
and U2920 (N_2920,In_1984,In_506);
and U2921 (N_2921,In_1962,In_734);
or U2922 (N_2922,In_2482,In_910);
and U2923 (N_2923,In_471,In_981);
and U2924 (N_2924,In_767,In_1603);
and U2925 (N_2925,In_1383,In_770);
nand U2926 (N_2926,In_1685,In_2368);
or U2927 (N_2927,In_515,In_1740);
and U2928 (N_2928,In_134,In_1769);
nor U2929 (N_2929,In_748,In_1574);
or U2930 (N_2930,In_679,In_222);
nor U2931 (N_2931,In_1973,In_2201);
and U2932 (N_2932,In_1147,In_178);
nand U2933 (N_2933,In_2039,In_2112);
nand U2934 (N_2934,In_1730,In_564);
nor U2935 (N_2935,In_2287,In_284);
and U2936 (N_2936,In_1305,In_580);
and U2937 (N_2937,In_2367,In_1206);
and U2938 (N_2938,In_2334,In_929);
or U2939 (N_2939,In_2125,In_74);
or U2940 (N_2940,In_1354,In_785);
and U2941 (N_2941,In_2300,In_815);
and U2942 (N_2942,In_1378,In_416);
xnor U2943 (N_2943,In_2356,In_1337);
or U2944 (N_2944,In_1993,In_926);
xor U2945 (N_2945,In_10,In_1395);
nor U2946 (N_2946,In_1559,In_2386);
nor U2947 (N_2947,In_2235,In_980);
xnor U2948 (N_2948,In_282,In_2239);
or U2949 (N_2949,In_183,In_2199);
or U2950 (N_2950,In_2048,In_2249);
nor U2951 (N_2951,In_2490,In_355);
and U2952 (N_2952,In_1758,In_2317);
or U2953 (N_2953,In_1115,In_278);
nand U2954 (N_2954,In_976,In_189);
nor U2955 (N_2955,In_1859,In_64);
nand U2956 (N_2956,In_1288,In_1717);
nor U2957 (N_2957,In_1381,In_884);
nor U2958 (N_2958,In_1124,In_2132);
or U2959 (N_2959,In_1690,In_910);
nand U2960 (N_2960,In_1950,In_324);
and U2961 (N_2961,In_1663,In_1403);
nand U2962 (N_2962,In_2436,In_249);
and U2963 (N_2963,In_1006,In_2244);
nand U2964 (N_2964,In_1577,In_1705);
and U2965 (N_2965,In_612,In_1356);
and U2966 (N_2966,In_1954,In_1572);
or U2967 (N_2967,In_496,In_180);
nand U2968 (N_2968,In_758,In_1828);
and U2969 (N_2969,In_2499,In_610);
nand U2970 (N_2970,In_1651,In_880);
nand U2971 (N_2971,In_1689,In_196);
nor U2972 (N_2972,In_1385,In_793);
and U2973 (N_2973,In_1924,In_2466);
nand U2974 (N_2974,In_1476,In_2184);
and U2975 (N_2975,In_385,In_2199);
or U2976 (N_2976,In_527,In_271);
nor U2977 (N_2977,In_1749,In_813);
nor U2978 (N_2978,In_964,In_659);
nand U2979 (N_2979,In_549,In_1253);
nor U2980 (N_2980,In_316,In_326);
nand U2981 (N_2981,In_785,In_682);
nand U2982 (N_2982,In_229,In_52);
nor U2983 (N_2983,In_797,In_964);
or U2984 (N_2984,In_760,In_366);
or U2985 (N_2985,In_1698,In_598);
xor U2986 (N_2986,In_59,In_1357);
or U2987 (N_2987,In_2075,In_1360);
xor U2988 (N_2988,In_1931,In_2111);
or U2989 (N_2989,In_34,In_2378);
nand U2990 (N_2990,In_635,In_802);
or U2991 (N_2991,In_1979,In_1086);
and U2992 (N_2992,In_503,In_1167);
nand U2993 (N_2993,In_65,In_2097);
nand U2994 (N_2994,In_1974,In_1555);
nand U2995 (N_2995,In_2284,In_1844);
and U2996 (N_2996,In_201,In_2120);
and U2997 (N_2997,In_475,In_549);
xor U2998 (N_2998,In_602,In_1663);
xnor U2999 (N_2999,In_2369,In_2178);
or U3000 (N_3000,In_2329,In_429);
nand U3001 (N_3001,In_299,In_413);
xnor U3002 (N_3002,In_836,In_1190);
nor U3003 (N_3003,In_1628,In_393);
or U3004 (N_3004,In_615,In_1276);
nand U3005 (N_3005,In_685,In_966);
or U3006 (N_3006,In_169,In_1437);
nor U3007 (N_3007,In_1975,In_202);
xor U3008 (N_3008,In_1866,In_338);
and U3009 (N_3009,In_254,In_1371);
nor U3010 (N_3010,In_1855,In_2007);
and U3011 (N_3011,In_1590,In_715);
nand U3012 (N_3012,In_252,In_1589);
or U3013 (N_3013,In_706,In_1882);
nand U3014 (N_3014,In_1582,In_1094);
or U3015 (N_3015,In_980,In_827);
and U3016 (N_3016,In_2499,In_2204);
and U3017 (N_3017,In_1102,In_610);
and U3018 (N_3018,In_1660,In_871);
nor U3019 (N_3019,In_1696,In_1095);
xor U3020 (N_3020,In_136,In_499);
or U3021 (N_3021,In_2254,In_633);
and U3022 (N_3022,In_444,In_2258);
and U3023 (N_3023,In_789,In_1903);
and U3024 (N_3024,In_1817,In_961);
and U3025 (N_3025,In_879,In_1627);
nor U3026 (N_3026,In_1487,In_2350);
nand U3027 (N_3027,In_1768,In_602);
or U3028 (N_3028,In_1182,In_1811);
or U3029 (N_3029,In_570,In_1679);
and U3030 (N_3030,In_1347,In_2128);
nor U3031 (N_3031,In_837,In_696);
nand U3032 (N_3032,In_842,In_2233);
or U3033 (N_3033,In_1659,In_1742);
and U3034 (N_3034,In_1821,In_1656);
nand U3035 (N_3035,In_2271,In_1193);
xnor U3036 (N_3036,In_1091,In_1429);
nand U3037 (N_3037,In_1659,In_250);
nor U3038 (N_3038,In_1326,In_484);
and U3039 (N_3039,In_2203,In_1235);
nor U3040 (N_3040,In_1522,In_1757);
nor U3041 (N_3041,In_10,In_117);
and U3042 (N_3042,In_682,In_1583);
or U3043 (N_3043,In_1545,In_1804);
nand U3044 (N_3044,In_2085,In_1187);
or U3045 (N_3045,In_260,In_666);
nand U3046 (N_3046,In_509,In_725);
xnor U3047 (N_3047,In_1933,In_373);
nor U3048 (N_3048,In_1946,In_655);
and U3049 (N_3049,In_18,In_896);
nor U3050 (N_3050,In_1405,In_632);
nor U3051 (N_3051,In_397,In_2457);
or U3052 (N_3052,In_172,In_429);
nor U3053 (N_3053,In_1148,In_240);
and U3054 (N_3054,In_1762,In_709);
or U3055 (N_3055,In_1099,In_531);
xnor U3056 (N_3056,In_379,In_1263);
nor U3057 (N_3057,In_154,In_2110);
nor U3058 (N_3058,In_2345,In_514);
or U3059 (N_3059,In_1409,In_61);
or U3060 (N_3060,In_494,In_2323);
xor U3061 (N_3061,In_2483,In_565);
and U3062 (N_3062,In_2441,In_2376);
and U3063 (N_3063,In_1747,In_1796);
and U3064 (N_3064,In_751,In_1423);
nor U3065 (N_3065,In_2424,In_1819);
or U3066 (N_3066,In_2122,In_539);
or U3067 (N_3067,In_368,In_2381);
nor U3068 (N_3068,In_1996,In_964);
xnor U3069 (N_3069,In_900,In_2213);
or U3070 (N_3070,In_514,In_313);
or U3071 (N_3071,In_1384,In_1161);
nand U3072 (N_3072,In_1120,In_1827);
and U3073 (N_3073,In_1248,In_417);
and U3074 (N_3074,In_967,In_907);
and U3075 (N_3075,In_492,In_777);
or U3076 (N_3076,In_2047,In_1121);
and U3077 (N_3077,In_1921,In_1337);
nor U3078 (N_3078,In_916,In_32);
nor U3079 (N_3079,In_1423,In_2289);
and U3080 (N_3080,In_1617,In_268);
nor U3081 (N_3081,In_1661,In_1551);
nor U3082 (N_3082,In_1713,In_990);
and U3083 (N_3083,In_2008,In_2328);
nor U3084 (N_3084,In_1838,In_1924);
xnor U3085 (N_3085,In_713,In_943);
nor U3086 (N_3086,In_509,In_1841);
or U3087 (N_3087,In_1134,In_876);
nand U3088 (N_3088,In_453,In_1352);
and U3089 (N_3089,In_2169,In_2479);
or U3090 (N_3090,In_896,In_2319);
or U3091 (N_3091,In_253,In_829);
and U3092 (N_3092,In_1522,In_711);
nor U3093 (N_3093,In_2147,In_314);
or U3094 (N_3094,In_2409,In_1870);
or U3095 (N_3095,In_1190,In_2495);
or U3096 (N_3096,In_2449,In_460);
nor U3097 (N_3097,In_1117,In_1300);
or U3098 (N_3098,In_1316,In_280);
or U3099 (N_3099,In_1851,In_1460);
nand U3100 (N_3100,In_364,In_150);
nor U3101 (N_3101,In_1682,In_1955);
nand U3102 (N_3102,In_1180,In_708);
nor U3103 (N_3103,In_638,In_1716);
nand U3104 (N_3104,In_1450,In_1518);
nand U3105 (N_3105,In_1777,In_928);
and U3106 (N_3106,In_827,In_2352);
xor U3107 (N_3107,In_1396,In_1625);
nor U3108 (N_3108,In_1474,In_2187);
nand U3109 (N_3109,In_258,In_2344);
xor U3110 (N_3110,In_1776,In_262);
nand U3111 (N_3111,In_531,In_276);
or U3112 (N_3112,In_1565,In_1633);
xnor U3113 (N_3113,In_227,In_1762);
or U3114 (N_3114,In_1213,In_1771);
xnor U3115 (N_3115,In_1567,In_1117);
nor U3116 (N_3116,In_1360,In_1800);
nand U3117 (N_3117,In_1223,In_1367);
nand U3118 (N_3118,In_1700,In_2057);
and U3119 (N_3119,In_471,In_822);
nor U3120 (N_3120,In_463,In_614);
or U3121 (N_3121,In_732,In_1467);
and U3122 (N_3122,In_1329,In_280);
or U3123 (N_3123,In_1222,In_1260);
and U3124 (N_3124,In_773,In_1790);
nand U3125 (N_3125,In_5,In_1345);
or U3126 (N_3126,In_1971,In_1424);
nor U3127 (N_3127,In_1117,In_190);
or U3128 (N_3128,In_2437,In_1401);
or U3129 (N_3129,In_2306,In_425);
and U3130 (N_3130,In_1040,In_1490);
or U3131 (N_3131,In_56,In_2240);
nor U3132 (N_3132,In_1697,In_2426);
xor U3133 (N_3133,In_2008,In_81);
nor U3134 (N_3134,In_1348,In_1421);
nand U3135 (N_3135,In_1624,In_441);
or U3136 (N_3136,In_1602,In_1188);
nand U3137 (N_3137,In_941,In_1871);
nor U3138 (N_3138,In_437,In_1778);
and U3139 (N_3139,In_1111,In_658);
or U3140 (N_3140,In_408,In_1163);
and U3141 (N_3141,In_1837,In_147);
nor U3142 (N_3142,In_2275,In_20);
and U3143 (N_3143,In_1353,In_1649);
nand U3144 (N_3144,In_1662,In_2362);
nor U3145 (N_3145,In_1618,In_108);
xor U3146 (N_3146,In_2118,In_951);
and U3147 (N_3147,In_386,In_1556);
nor U3148 (N_3148,In_2254,In_792);
or U3149 (N_3149,In_2207,In_1297);
or U3150 (N_3150,In_1496,In_1769);
nand U3151 (N_3151,In_2028,In_259);
nand U3152 (N_3152,In_1804,In_1587);
nor U3153 (N_3153,In_833,In_1357);
xnor U3154 (N_3154,In_2014,In_717);
nor U3155 (N_3155,In_2177,In_541);
nor U3156 (N_3156,In_73,In_95);
or U3157 (N_3157,In_51,In_1711);
nand U3158 (N_3158,In_1497,In_1092);
xnor U3159 (N_3159,In_887,In_588);
nand U3160 (N_3160,In_2224,In_1955);
nor U3161 (N_3161,In_2409,In_1306);
and U3162 (N_3162,In_665,In_1493);
and U3163 (N_3163,In_434,In_777);
nor U3164 (N_3164,In_991,In_2478);
nor U3165 (N_3165,In_920,In_1900);
and U3166 (N_3166,In_1383,In_628);
or U3167 (N_3167,In_1716,In_2186);
and U3168 (N_3168,In_5,In_1715);
nand U3169 (N_3169,In_798,In_1950);
and U3170 (N_3170,In_603,In_1027);
nor U3171 (N_3171,In_2219,In_408);
nor U3172 (N_3172,In_1174,In_433);
and U3173 (N_3173,In_2464,In_1724);
and U3174 (N_3174,In_2045,In_2287);
xor U3175 (N_3175,In_1354,In_1445);
or U3176 (N_3176,In_304,In_2489);
nor U3177 (N_3177,In_814,In_425);
or U3178 (N_3178,In_2263,In_1757);
or U3179 (N_3179,In_1641,In_1351);
nand U3180 (N_3180,In_265,In_2479);
and U3181 (N_3181,In_1515,In_1149);
and U3182 (N_3182,In_4,In_2293);
and U3183 (N_3183,In_925,In_1796);
xor U3184 (N_3184,In_265,In_1661);
nand U3185 (N_3185,In_1237,In_2287);
and U3186 (N_3186,In_607,In_468);
or U3187 (N_3187,In_2179,In_2032);
and U3188 (N_3188,In_1449,In_1389);
or U3189 (N_3189,In_298,In_1984);
xor U3190 (N_3190,In_661,In_358);
or U3191 (N_3191,In_2308,In_1635);
or U3192 (N_3192,In_2494,In_703);
nand U3193 (N_3193,In_514,In_1443);
nand U3194 (N_3194,In_1050,In_1977);
nor U3195 (N_3195,In_1733,In_1239);
and U3196 (N_3196,In_2460,In_1922);
nor U3197 (N_3197,In_645,In_1209);
or U3198 (N_3198,In_634,In_1114);
nand U3199 (N_3199,In_354,In_2235);
nand U3200 (N_3200,In_1496,In_140);
nor U3201 (N_3201,In_2210,In_1771);
or U3202 (N_3202,In_727,In_1785);
and U3203 (N_3203,In_1967,In_2006);
nand U3204 (N_3204,In_1397,In_1962);
nand U3205 (N_3205,In_2067,In_2220);
nor U3206 (N_3206,In_454,In_762);
nor U3207 (N_3207,In_399,In_1756);
nand U3208 (N_3208,In_1680,In_1271);
nand U3209 (N_3209,In_2481,In_91);
nor U3210 (N_3210,In_1425,In_1344);
or U3211 (N_3211,In_1171,In_2367);
or U3212 (N_3212,In_2477,In_1612);
xnor U3213 (N_3213,In_1826,In_141);
nand U3214 (N_3214,In_189,In_1129);
xor U3215 (N_3215,In_2410,In_977);
and U3216 (N_3216,In_301,In_1951);
or U3217 (N_3217,In_1428,In_1365);
xor U3218 (N_3218,In_1204,In_1265);
nor U3219 (N_3219,In_2204,In_772);
nand U3220 (N_3220,In_1860,In_1818);
nand U3221 (N_3221,In_753,In_662);
xor U3222 (N_3222,In_1834,In_1647);
and U3223 (N_3223,In_1316,In_1224);
nand U3224 (N_3224,In_2246,In_2361);
nor U3225 (N_3225,In_403,In_134);
or U3226 (N_3226,In_2283,In_1287);
xnor U3227 (N_3227,In_1893,In_770);
or U3228 (N_3228,In_1239,In_1707);
and U3229 (N_3229,In_969,In_1924);
nand U3230 (N_3230,In_2209,In_217);
and U3231 (N_3231,In_1743,In_1478);
or U3232 (N_3232,In_2,In_1709);
nor U3233 (N_3233,In_1624,In_842);
nor U3234 (N_3234,In_2204,In_528);
nor U3235 (N_3235,In_812,In_974);
or U3236 (N_3236,In_1754,In_2377);
nor U3237 (N_3237,In_1696,In_2361);
nor U3238 (N_3238,In_2309,In_2066);
or U3239 (N_3239,In_1418,In_1769);
nor U3240 (N_3240,In_2017,In_2248);
and U3241 (N_3241,In_645,In_2401);
nand U3242 (N_3242,In_1489,In_168);
and U3243 (N_3243,In_678,In_2245);
nand U3244 (N_3244,In_1552,In_2481);
or U3245 (N_3245,In_2374,In_1201);
and U3246 (N_3246,In_731,In_2431);
xnor U3247 (N_3247,In_163,In_1149);
and U3248 (N_3248,In_595,In_944);
or U3249 (N_3249,In_478,In_202);
xor U3250 (N_3250,In_197,In_1103);
nor U3251 (N_3251,In_311,In_718);
nand U3252 (N_3252,In_2091,In_1943);
or U3253 (N_3253,In_656,In_1566);
nor U3254 (N_3254,In_1307,In_1534);
and U3255 (N_3255,In_774,In_2084);
and U3256 (N_3256,In_366,In_1877);
or U3257 (N_3257,In_1420,In_1856);
nor U3258 (N_3258,In_679,In_609);
nand U3259 (N_3259,In_675,In_2127);
and U3260 (N_3260,In_2436,In_1281);
and U3261 (N_3261,In_2028,In_1103);
and U3262 (N_3262,In_1041,In_1921);
and U3263 (N_3263,In_1036,In_1157);
nand U3264 (N_3264,In_2466,In_1);
nor U3265 (N_3265,In_142,In_876);
and U3266 (N_3266,In_1759,In_2301);
and U3267 (N_3267,In_699,In_1047);
nor U3268 (N_3268,In_1271,In_2233);
or U3269 (N_3269,In_284,In_997);
nand U3270 (N_3270,In_2002,In_2263);
or U3271 (N_3271,In_2293,In_60);
nor U3272 (N_3272,In_862,In_629);
nor U3273 (N_3273,In_266,In_304);
nor U3274 (N_3274,In_2215,In_1545);
nor U3275 (N_3275,In_521,In_2222);
or U3276 (N_3276,In_93,In_1157);
nor U3277 (N_3277,In_1989,In_1491);
nor U3278 (N_3278,In_58,In_1959);
nand U3279 (N_3279,In_186,In_1816);
and U3280 (N_3280,In_1124,In_75);
or U3281 (N_3281,In_2171,In_1739);
nand U3282 (N_3282,In_2277,In_2327);
nand U3283 (N_3283,In_147,In_1104);
xor U3284 (N_3284,In_1317,In_835);
and U3285 (N_3285,In_2055,In_133);
nor U3286 (N_3286,In_1137,In_1067);
or U3287 (N_3287,In_651,In_2114);
nand U3288 (N_3288,In_591,In_1598);
or U3289 (N_3289,In_1511,In_1272);
nor U3290 (N_3290,In_2137,In_303);
and U3291 (N_3291,In_1870,In_2205);
or U3292 (N_3292,In_1426,In_2125);
and U3293 (N_3293,In_2319,In_2477);
or U3294 (N_3294,In_1558,In_601);
nand U3295 (N_3295,In_198,In_2472);
or U3296 (N_3296,In_136,In_455);
nor U3297 (N_3297,In_1145,In_945);
and U3298 (N_3298,In_652,In_177);
and U3299 (N_3299,In_1486,In_126);
nand U3300 (N_3300,In_213,In_520);
nor U3301 (N_3301,In_1068,In_256);
nand U3302 (N_3302,In_1276,In_1829);
nand U3303 (N_3303,In_1383,In_2386);
and U3304 (N_3304,In_1500,In_1687);
and U3305 (N_3305,In_665,In_2204);
nor U3306 (N_3306,In_862,In_252);
xnor U3307 (N_3307,In_194,In_242);
nand U3308 (N_3308,In_49,In_2229);
and U3309 (N_3309,In_775,In_758);
and U3310 (N_3310,In_1976,In_1844);
and U3311 (N_3311,In_2032,In_355);
nand U3312 (N_3312,In_979,In_262);
or U3313 (N_3313,In_1847,In_1907);
nand U3314 (N_3314,In_993,In_1252);
nor U3315 (N_3315,In_972,In_1212);
nand U3316 (N_3316,In_1121,In_1217);
or U3317 (N_3317,In_2449,In_996);
nand U3318 (N_3318,In_1063,In_65);
and U3319 (N_3319,In_1633,In_567);
nor U3320 (N_3320,In_613,In_1310);
and U3321 (N_3321,In_1777,In_51);
or U3322 (N_3322,In_757,In_1676);
and U3323 (N_3323,In_782,In_1461);
xnor U3324 (N_3324,In_455,In_1707);
nor U3325 (N_3325,In_510,In_1618);
xnor U3326 (N_3326,In_1127,In_477);
and U3327 (N_3327,In_2446,In_1683);
nand U3328 (N_3328,In_4,In_357);
nand U3329 (N_3329,In_706,In_1625);
nand U3330 (N_3330,In_10,In_478);
xnor U3331 (N_3331,In_2383,In_2419);
or U3332 (N_3332,In_668,In_1407);
nand U3333 (N_3333,In_1980,In_1378);
nor U3334 (N_3334,In_1352,In_1920);
xor U3335 (N_3335,In_2144,In_1102);
nor U3336 (N_3336,In_558,In_1031);
and U3337 (N_3337,In_2245,In_1719);
xnor U3338 (N_3338,In_909,In_917);
or U3339 (N_3339,In_597,In_453);
xnor U3340 (N_3340,In_2277,In_535);
nand U3341 (N_3341,In_906,In_397);
xnor U3342 (N_3342,In_1572,In_531);
nand U3343 (N_3343,In_606,In_1730);
nor U3344 (N_3344,In_1319,In_1014);
and U3345 (N_3345,In_2310,In_1923);
and U3346 (N_3346,In_992,In_1595);
xnor U3347 (N_3347,In_1971,In_1876);
or U3348 (N_3348,In_1169,In_1420);
and U3349 (N_3349,In_1131,In_869);
and U3350 (N_3350,In_343,In_530);
or U3351 (N_3351,In_1251,In_1242);
nor U3352 (N_3352,In_1474,In_378);
or U3353 (N_3353,In_751,In_1333);
and U3354 (N_3354,In_445,In_2161);
and U3355 (N_3355,In_1881,In_293);
nand U3356 (N_3356,In_1695,In_2232);
nor U3357 (N_3357,In_430,In_2413);
and U3358 (N_3358,In_193,In_2397);
nand U3359 (N_3359,In_652,In_2417);
xnor U3360 (N_3360,In_1673,In_1554);
nand U3361 (N_3361,In_563,In_1283);
nor U3362 (N_3362,In_2310,In_874);
nor U3363 (N_3363,In_1823,In_1735);
and U3364 (N_3364,In_857,In_1944);
and U3365 (N_3365,In_1293,In_293);
and U3366 (N_3366,In_733,In_1342);
or U3367 (N_3367,In_2140,In_2157);
or U3368 (N_3368,In_1595,In_1340);
or U3369 (N_3369,In_1479,In_605);
nand U3370 (N_3370,In_308,In_2485);
or U3371 (N_3371,In_1512,In_1894);
nor U3372 (N_3372,In_2412,In_2388);
or U3373 (N_3373,In_524,In_2323);
nand U3374 (N_3374,In_1911,In_540);
and U3375 (N_3375,In_1041,In_496);
nor U3376 (N_3376,In_218,In_185);
and U3377 (N_3377,In_2094,In_2243);
nor U3378 (N_3378,In_733,In_341);
nand U3379 (N_3379,In_2215,In_213);
nor U3380 (N_3380,In_2424,In_1341);
and U3381 (N_3381,In_460,In_2341);
or U3382 (N_3382,In_594,In_1980);
or U3383 (N_3383,In_713,In_2485);
or U3384 (N_3384,In_1142,In_569);
and U3385 (N_3385,In_713,In_2393);
nand U3386 (N_3386,In_1866,In_1375);
xnor U3387 (N_3387,In_1083,In_1983);
and U3388 (N_3388,In_1656,In_1478);
nand U3389 (N_3389,In_1214,In_712);
or U3390 (N_3390,In_303,In_584);
nand U3391 (N_3391,In_1504,In_1289);
nor U3392 (N_3392,In_2219,In_1797);
or U3393 (N_3393,In_2314,In_607);
or U3394 (N_3394,In_859,In_820);
xor U3395 (N_3395,In_269,In_2082);
nor U3396 (N_3396,In_1263,In_217);
nor U3397 (N_3397,In_176,In_920);
or U3398 (N_3398,In_1795,In_1127);
xnor U3399 (N_3399,In_589,In_1931);
nand U3400 (N_3400,In_1949,In_272);
and U3401 (N_3401,In_1499,In_379);
and U3402 (N_3402,In_2086,In_585);
nand U3403 (N_3403,In_175,In_1053);
and U3404 (N_3404,In_1434,In_895);
and U3405 (N_3405,In_71,In_1088);
nand U3406 (N_3406,In_2446,In_2347);
and U3407 (N_3407,In_2005,In_481);
or U3408 (N_3408,In_362,In_1723);
or U3409 (N_3409,In_1701,In_1703);
xnor U3410 (N_3410,In_236,In_2217);
or U3411 (N_3411,In_455,In_194);
xnor U3412 (N_3412,In_1791,In_1247);
nand U3413 (N_3413,In_1648,In_634);
and U3414 (N_3414,In_595,In_2204);
nand U3415 (N_3415,In_1830,In_1319);
and U3416 (N_3416,In_603,In_2224);
or U3417 (N_3417,In_865,In_2428);
nor U3418 (N_3418,In_1843,In_153);
xor U3419 (N_3419,In_1422,In_736);
or U3420 (N_3420,In_1495,In_1167);
and U3421 (N_3421,In_1845,In_2235);
nor U3422 (N_3422,In_968,In_655);
nor U3423 (N_3423,In_260,In_1251);
nand U3424 (N_3424,In_946,In_498);
or U3425 (N_3425,In_534,In_1345);
or U3426 (N_3426,In_1130,In_1800);
xor U3427 (N_3427,In_352,In_1683);
and U3428 (N_3428,In_2073,In_1892);
and U3429 (N_3429,In_1926,In_907);
or U3430 (N_3430,In_1811,In_1144);
nand U3431 (N_3431,In_1424,In_2242);
nand U3432 (N_3432,In_1541,In_299);
nand U3433 (N_3433,In_505,In_1469);
nand U3434 (N_3434,In_698,In_1072);
nand U3435 (N_3435,In_1310,In_1488);
nand U3436 (N_3436,In_470,In_846);
nor U3437 (N_3437,In_1908,In_1102);
nand U3438 (N_3438,In_1042,In_2217);
or U3439 (N_3439,In_520,In_21);
nand U3440 (N_3440,In_1931,In_1268);
nor U3441 (N_3441,In_471,In_2051);
or U3442 (N_3442,In_1008,In_1083);
or U3443 (N_3443,In_308,In_653);
nand U3444 (N_3444,In_1313,In_601);
or U3445 (N_3445,In_1388,In_2268);
and U3446 (N_3446,In_1609,In_37);
and U3447 (N_3447,In_2329,In_2163);
nand U3448 (N_3448,In_2003,In_1821);
nor U3449 (N_3449,In_1405,In_999);
nand U3450 (N_3450,In_714,In_2027);
and U3451 (N_3451,In_1273,In_1932);
and U3452 (N_3452,In_168,In_196);
nand U3453 (N_3453,In_742,In_755);
nor U3454 (N_3454,In_2187,In_627);
or U3455 (N_3455,In_482,In_2430);
nor U3456 (N_3456,In_2235,In_1708);
or U3457 (N_3457,In_138,In_1196);
nor U3458 (N_3458,In_2440,In_458);
nand U3459 (N_3459,In_1289,In_2441);
and U3460 (N_3460,In_2375,In_1651);
or U3461 (N_3461,In_2129,In_1985);
nor U3462 (N_3462,In_471,In_2072);
xor U3463 (N_3463,In_1643,In_2089);
nor U3464 (N_3464,In_452,In_1792);
or U3465 (N_3465,In_1496,In_853);
and U3466 (N_3466,In_1076,In_421);
nand U3467 (N_3467,In_709,In_1178);
nand U3468 (N_3468,In_324,In_2454);
xor U3469 (N_3469,In_2411,In_1893);
nor U3470 (N_3470,In_1973,In_2127);
nand U3471 (N_3471,In_2495,In_1647);
nor U3472 (N_3472,In_1296,In_1726);
nand U3473 (N_3473,In_2372,In_752);
xnor U3474 (N_3474,In_868,In_1585);
nand U3475 (N_3475,In_660,In_2230);
nand U3476 (N_3476,In_810,In_474);
nor U3477 (N_3477,In_33,In_2440);
or U3478 (N_3478,In_2278,In_773);
nor U3479 (N_3479,In_2143,In_883);
or U3480 (N_3480,In_2106,In_2124);
nand U3481 (N_3481,In_1730,In_1835);
nand U3482 (N_3482,In_1129,In_448);
nor U3483 (N_3483,In_1843,In_1044);
and U3484 (N_3484,In_125,In_987);
and U3485 (N_3485,In_1237,In_1369);
xnor U3486 (N_3486,In_1971,In_314);
nor U3487 (N_3487,In_995,In_1726);
xor U3488 (N_3488,In_1492,In_1320);
nor U3489 (N_3489,In_1875,In_1502);
nand U3490 (N_3490,In_612,In_494);
or U3491 (N_3491,In_1078,In_678);
nand U3492 (N_3492,In_1782,In_947);
and U3493 (N_3493,In_1787,In_1671);
and U3494 (N_3494,In_239,In_737);
and U3495 (N_3495,In_1729,In_1955);
nor U3496 (N_3496,In_1018,In_189);
and U3497 (N_3497,In_151,In_807);
nand U3498 (N_3498,In_31,In_268);
nor U3499 (N_3499,In_72,In_558);
or U3500 (N_3500,In_1767,In_2069);
or U3501 (N_3501,In_1327,In_735);
or U3502 (N_3502,In_1277,In_470);
nand U3503 (N_3503,In_486,In_35);
nor U3504 (N_3504,In_1035,In_580);
nand U3505 (N_3505,In_1116,In_674);
nor U3506 (N_3506,In_953,In_212);
xor U3507 (N_3507,In_2029,In_437);
nand U3508 (N_3508,In_534,In_1711);
xor U3509 (N_3509,In_1541,In_305);
nor U3510 (N_3510,In_155,In_2264);
and U3511 (N_3511,In_273,In_2173);
nor U3512 (N_3512,In_2316,In_484);
or U3513 (N_3513,In_2403,In_2472);
nor U3514 (N_3514,In_256,In_2008);
or U3515 (N_3515,In_436,In_1591);
nor U3516 (N_3516,In_1137,In_925);
or U3517 (N_3517,In_2344,In_892);
nand U3518 (N_3518,In_788,In_1786);
nor U3519 (N_3519,In_1465,In_119);
nand U3520 (N_3520,In_2122,In_5);
nor U3521 (N_3521,In_2480,In_2089);
and U3522 (N_3522,In_2093,In_2438);
and U3523 (N_3523,In_1273,In_2370);
and U3524 (N_3524,In_1312,In_352);
nor U3525 (N_3525,In_1505,In_2267);
and U3526 (N_3526,In_2474,In_1805);
nand U3527 (N_3527,In_1694,In_67);
nand U3528 (N_3528,In_483,In_1187);
nor U3529 (N_3529,In_1340,In_1248);
or U3530 (N_3530,In_386,In_771);
nor U3531 (N_3531,In_340,In_972);
xnor U3532 (N_3532,In_2068,In_517);
or U3533 (N_3533,In_1100,In_927);
and U3534 (N_3534,In_272,In_1323);
xnor U3535 (N_3535,In_988,In_1470);
nand U3536 (N_3536,In_1014,In_340);
xnor U3537 (N_3537,In_105,In_1095);
and U3538 (N_3538,In_976,In_365);
nand U3539 (N_3539,In_946,In_22);
nand U3540 (N_3540,In_2265,In_1339);
nor U3541 (N_3541,In_1688,In_1451);
or U3542 (N_3542,In_544,In_2346);
nor U3543 (N_3543,In_1281,In_1499);
or U3544 (N_3544,In_667,In_1360);
nand U3545 (N_3545,In_2114,In_1939);
or U3546 (N_3546,In_1867,In_41);
and U3547 (N_3547,In_2024,In_1994);
nor U3548 (N_3548,In_493,In_1882);
xnor U3549 (N_3549,In_868,In_472);
xnor U3550 (N_3550,In_471,In_1485);
nor U3551 (N_3551,In_1866,In_297);
and U3552 (N_3552,In_595,In_1163);
and U3553 (N_3553,In_950,In_1853);
and U3554 (N_3554,In_2320,In_533);
and U3555 (N_3555,In_2458,In_1826);
or U3556 (N_3556,In_239,In_451);
or U3557 (N_3557,In_2098,In_1040);
and U3558 (N_3558,In_1788,In_934);
xor U3559 (N_3559,In_1646,In_1124);
and U3560 (N_3560,In_1247,In_11);
xnor U3561 (N_3561,In_90,In_2045);
or U3562 (N_3562,In_1653,In_1784);
or U3563 (N_3563,In_948,In_652);
and U3564 (N_3564,In_75,In_595);
nand U3565 (N_3565,In_2416,In_1060);
xor U3566 (N_3566,In_1322,In_1840);
and U3567 (N_3567,In_481,In_390);
xnor U3568 (N_3568,In_1661,In_1856);
nor U3569 (N_3569,In_669,In_955);
nand U3570 (N_3570,In_1585,In_1098);
or U3571 (N_3571,In_1140,In_2108);
xor U3572 (N_3572,In_940,In_1278);
and U3573 (N_3573,In_1181,In_590);
and U3574 (N_3574,In_1678,In_152);
nand U3575 (N_3575,In_2186,In_1424);
nor U3576 (N_3576,In_717,In_526);
nand U3577 (N_3577,In_541,In_2363);
and U3578 (N_3578,In_244,In_1147);
or U3579 (N_3579,In_2252,In_1913);
nand U3580 (N_3580,In_1126,In_518);
xor U3581 (N_3581,In_129,In_771);
nand U3582 (N_3582,In_513,In_287);
nor U3583 (N_3583,In_979,In_1944);
nor U3584 (N_3584,In_369,In_134);
and U3585 (N_3585,In_2101,In_541);
and U3586 (N_3586,In_1016,In_123);
nand U3587 (N_3587,In_463,In_34);
and U3588 (N_3588,In_33,In_834);
nand U3589 (N_3589,In_1680,In_380);
nand U3590 (N_3590,In_2301,In_914);
nand U3591 (N_3591,In_2237,In_221);
and U3592 (N_3592,In_910,In_904);
nor U3593 (N_3593,In_2318,In_2177);
and U3594 (N_3594,In_481,In_549);
or U3595 (N_3595,In_343,In_1097);
xor U3596 (N_3596,In_1321,In_199);
nand U3597 (N_3597,In_914,In_404);
and U3598 (N_3598,In_1483,In_2056);
and U3599 (N_3599,In_755,In_345);
nand U3600 (N_3600,In_1629,In_1925);
nand U3601 (N_3601,In_225,In_871);
xnor U3602 (N_3602,In_1716,In_14);
nand U3603 (N_3603,In_854,In_2098);
nand U3604 (N_3604,In_2337,In_2078);
nand U3605 (N_3605,In_1732,In_199);
or U3606 (N_3606,In_1532,In_2231);
nor U3607 (N_3607,In_1077,In_2099);
and U3608 (N_3608,In_1261,In_592);
nand U3609 (N_3609,In_381,In_2307);
or U3610 (N_3610,In_2312,In_2039);
and U3611 (N_3611,In_1858,In_2062);
and U3612 (N_3612,In_753,In_634);
and U3613 (N_3613,In_1447,In_347);
nand U3614 (N_3614,In_479,In_745);
nand U3615 (N_3615,In_2055,In_1373);
or U3616 (N_3616,In_2023,In_1125);
and U3617 (N_3617,In_939,In_1154);
nor U3618 (N_3618,In_1950,In_1704);
xor U3619 (N_3619,In_2179,In_1585);
nor U3620 (N_3620,In_889,In_1800);
nand U3621 (N_3621,In_878,In_26);
and U3622 (N_3622,In_1085,In_1769);
and U3623 (N_3623,In_605,In_1568);
nor U3624 (N_3624,In_1041,In_2404);
and U3625 (N_3625,In_535,In_223);
nor U3626 (N_3626,In_2496,In_2245);
nor U3627 (N_3627,In_1636,In_184);
nor U3628 (N_3628,In_1312,In_419);
nor U3629 (N_3629,In_2141,In_1526);
nand U3630 (N_3630,In_1663,In_579);
nor U3631 (N_3631,In_2297,In_2337);
nor U3632 (N_3632,In_1511,In_774);
xor U3633 (N_3633,In_726,In_1641);
nor U3634 (N_3634,In_2151,In_1554);
and U3635 (N_3635,In_19,In_2469);
nor U3636 (N_3636,In_1281,In_307);
nor U3637 (N_3637,In_1599,In_1300);
xnor U3638 (N_3638,In_349,In_1557);
or U3639 (N_3639,In_1389,In_2249);
and U3640 (N_3640,In_1299,In_2333);
and U3641 (N_3641,In_279,In_2357);
nand U3642 (N_3642,In_1303,In_99);
or U3643 (N_3643,In_227,In_922);
and U3644 (N_3644,In_2297,In_1910);
or U3645 (N_3645,In_715,In_1132);
or U3646 (N_3646,In_2463,In_348);
nand U3647 (N_3647,In_182,In_1449);
or U3648 (N_3648,In_83,In_238);
nor U3649 (N_3649,In_428,In_1052);
nand U3650 (N_3650,In_1025,In_364);
or U3651 (N_3651,In_510,In_2077);
or U3652 (N_3652,In_292,In_2220);
or U3653 (N_3653,In_2453,In_1689);
and U3654 (N_3654,In_594,In_2009);
nor U3655 (N_3655,In_1769,In_2054);
nand U3656 (N_3656,In_604,In_406);
nand U3657 (N_3657,In_2284,In_213);
or U3658 (N_3658,In_395,In_359);
nand U3659 (N_3659,In_2070,In_1674);
xor U3660 (N_3660,In_1346,In_2127);
nand U3661 (N_3661,In_1130,In_1107);
nand U3662 (N_3662,In_1954,In_954);
or U3663 (N_3663,In_891,In_2090);
and U3664 (N_3664,In_2026,In_2108);
and U3665 (N_3665,In_2368,In_1093);
and U3666 (N_3666,In_455,In_530);
and U3667 (N_3667,In_619,In_2293);
nand U3668 (N_3668,In_67,In_1960);
xor U3669 (N_3669,In_424,In_1442);
nor U3670 (N_3670,In_1332,In_129);
xor U3671 (N_3671,In_837,In_483);
or U3672 (N_3672,In_1955,In_1972);
or U3673 (N_3673,In_2366,In_1864);
nand U3674 (N_3674,In_920,In_1162);
and U3675 (N_3675,In_141,In_604);
nand U3676 (N_3676,In_243,In_2087);
nand U3677 (N_3677,In_1985,In_1063);
and U3678 (N_3678,In_1192,In_1773);
nor U3679 (N_3679,In_244,In_1233);
nand U3680 (N_3680,In_785,In_539);
and U3681 (N_3681,In_242,In_2334);
and U3682 (N_3682,In_1736,In_931);
nor U3683 (N_3683,In_556,In_1437);
nand U3684 (N_3684,In_1522,In_2048);
and U3685 (N_3685,In_1228,In_1575);
or U3686 (N_3686,In_1768,In_1831);
or U3687 (N_3687,In_1893,In_539);
nor U3688 (N_3688,In_2370,In_842);
or U3689 (N_3689,In_1229,In_1060);
nand U3690 (N_3690,In_169,In_1771);
or U3691 (N_3691,In_1607,In_2256);
nand U3692 (N_3692,In_670,In_31);
xor U3693 (N_3693,In_2218,In_122);
nand U3694 (N_3694,In_50,In_1291);
nor U3695 (N_3695,In_1042,In_993);
nand U3696 (N_3696,In_2442,In_1479);
nand U3697 (N_3697,In_462,In_1528);
nor U3698 (N_3698,In_487,In_1696);
nand U3699 (N_3699,In_1080,In_2455);
and U3700 (N_3700,In_687,In_976);
or U3701 (N_3701,In_832,In_1251);
nor U3702 (N_3702,In_2154,In_2227);
nor U3703 (N_3703,In_378,In_1200);
nand U3704 (N_3704,In_795,In_646);
or U3705 (N_3705,In_312,In_141);
or U3706 (N_3706,In_1432,In_373);
nand U3707 (N_3707,In_8,In_1039);
xor U3708 (N_3708,In_1705,In_2024);
or U3709 (N_3709,In_177,In_447);
nor U3710 (N_3710,In_1785,In_1833);
and U3711 (N_3711,In_1030,In_133);
or U3712 (N_3712,In_1665,In_2490);
nand U3713 (N_3713,In_2493,In_1059);
nor U3714 (N_3714,In_1661,In_2040);
and U3715 (N_3715,In_209,In_1859);
nor U3716 (N_3716,In_2221,In_988);
nor U3717 (N_3717,In_59,In_841);
and U3718 (N_3718,In_1684,In_1043);
xor U3719 (N_3719,In_381,In_1494);
or U3720 (N_3720,In_51,In_2051);
and U3721 (N_3721,In_1979,In_374);
and U3722 (N_3722,In_1322,In_899);
or U3723 (N_3723,In_992,In_2490);
nand U3724 (N_3724,In_2202,In_2177);
nand U3725 (N_3725,In_940,In_641);
nand U3726 (N_3726,In_1578,In_1537);
nand U3727 (N_3727,In_234,In_1148);
and U3728 (N_3728,In_835,In_890);
and U3729 (N_3729,In_419,In_567);
and U3730 (N_3730,In_912,In_1786);
and U3731 (N_3731,In_1612,In_120);
nor U3732 (N_3732,In_363,In_2367);
and U3733 (N_3733,In_1741,In_2225);
and U3734 (N_3734,In_480,In_151);
and U3735 (N_3735,In_1151,In_1137);
and U3736 (N_3736,In_2109,In_981);
nor U3737 (N_3737,In_556,In_2394);
nand U3738 (N_3738,In_2430,In_2123);
and U3739 (N_3739,In_391,In_1815);
or U3740 (N_3740,In_1433,In_411);
xor U3741 (N_3741,In_328,In_1807);
and U3742 (N_3742,In_432,In_1622);
nor U3743 (N_3743,In_427,In_2051);
and U3744 (N_3744,In_2427,In_1940);
nand U3745 (N_3745,In_285,In_2332);
nand U3746 (N_3746,In_2106,In_1153);
or U3747 (N_3747,In_2106,In_479);
and U3748 (N_3748,In_1599,In_1738);
nand U3749 (N_3749,In_1795,In_1865);
nand U3750 (N_3750,In_1071,In_2009);
and U3751 (N_3751,In_671,In_1825);
nand U3752 (N_3752,In_2031,In_704);
or U3753 (N_3753,In_2139,In_1517);
xnor U3754 (N_3754,In_2484,In_1993);
nand U3755 (N_3755,In_2172,In_2422);
or U3756 (N_3756,In_1172,In_2377);
and U3757 (N_3757,In_2058,In_2067);
and U3758 (N_3758,In_569,In_873);
and U3759 (N_3759,In_807,In_268);
xnor U3760 (N_3760,In_2168,In_896);
nand U3761 (N_3761,In_1771,In_1024);
or U3762 (N_3762,In_1799,In_1044);
and U3763 (N_3763,In_1453,In_1454);
nand U3764 (N_3764,In_254,In_2129);
and U3765 (N_3765,In_953,In_789);
and U3766 (N_3766,In_2449,In_1869);
and U3767 (N_3767,In_87,In_129);
nand U3768 (N_3768,In_819,In_416);
nand U3769 (N_3769,In_380,In_1741);
nand U3770 (N_3770,In_1823,In_304);
nor U3771 (N_3771,In_1569,In_338);
nor U3772 (N_3772,In_521,In_645);
and U3773 (N_3773,In_2011,In_355);
xnor U3774 (N_3774,In_2147,In_1957);
or U3775 (N_3775,In_139,In_253);
nand U3776 (N_3776,In_2238,In_352);
nor U3777 (N_3777,In_1154,In_1607);
xnor U3778 (N_3778,In_1547,In_799);
nor U3779 (N_3779,In_1418,In_406);
nor U3780 (N_3780,In_417,In_1295);
and U3781 (N_3781,In_1091,In_2415);
nor U3782 (N_3782,In_312,In_2095);
or U3783 (N_3783,In_1058,In_1202);
nand U3784 (N_3784,In_1917,In_1934);
nand U3785 (N_3785,In_1410,In_2308);
and U3786 (N_3786,In_303,In_259);
and U3787 (N_3787,In_1730,In_1474);
nand U3788 (N_3788,In_1844,In_1314);
or U3789 (N_3789,In_649,In_2351);
and U3790 (N_3790,In_1762,In_1311);
or U3791 (N_3791,In_754,In_1272);
nor U3792 (N_3792,In_2493,In_1752);
nor U3793 (N_3793,In_815,In_158);
nand U3794 (N_3794,In_752,In_1160);
nand U3795 (N_3795,In_23,In_15);
or U3796 (N_3796,In_244,In_1029);
nand U3797 (N_3797,In_2301,In_1242);
and U3798 (N_3798,In_394,In_323);
or U3799 (N_3799,In_1578,In_2230);
xnor U3800 (N_3800,In_1162,In_1658);
or U3801 (N_3801,In_1787,In_230);
and U3802 (N_3802,In_2208,In_148);
nor U3803 (N_3803,In_1980,In_2170);
or U3804 (N_3804,In_2353,In_555);
nand U3805 (N_3805,In_2376,In_94);
or U3806 (N_3806,In_1371,In_352);
nor U3807 (N_3807,In_827,In_1011);
nor U3808 (N_3808,In_1315,In_2499);
xnor U3809 (N_3809,In_1433,In_611);
xor U3810 (N_3810,In_1149,In_643);
or U3811 (N_3811,In_1152,In_434);
nor U3812 (N_3812,In_914,In_204);
xnor U3813 (N_3813,In_1713,In_1241);
or U3814 (N_3814,In_1969,In_1054);
nor U3815 (N_3815,In_2270,In_1818);
nor U3816 (N_3816,In_1210,In_786);
nor U3817 (N_3817,In_2400,In_1181);
and U3818 (N_3818,In_166,In_333);
and U3819 (N_3819,In_1310,In_210);
nand U3820 (N_3820,In_1822,In_2368);
or U3821 (N_3821,In_525,In_1826);
nor U3822 (N_3822,In_866,In_1228);
and U3823 (N_3823,In_18,In_2289);
nor U3824 (N_3824,In_2249,In_1630);
nand U3825 (N_3825,In_1047,In_205);
nor U3826 (N_3826,In_154,In_2444);
nor U3827 (N_3827,In_796,In_923);
nor U3828 (N_3828,In_1247,In_1989);
and U3829 (N_3829,In_677,In_1164);
nor U3830 (N_3830,In_1726,In_1282);
xor U3831 (N_3831,In_1983,In_368);
xor U3832 (N_3832,In_1911,In_892);
nor U3833 (N_3833,In_121,In_744);
or U3834 (N_3834,In_1780,In_1216);
nand U3835 (N_3835,In_1269,In_1542);
and U3836 (N_3836,In_1309,In_1534);
nand U3837 (N_3837,In_1375,In_2302);
xnor U3838 (N_3838,In_2103,In_925);
nand U3839 (N_3839,In_2189,In_748);
and U3840 (N_3840,In_1015,In_139);
and U3841 (N_3841,In_1559,In_2163);
nand U3842 (N_3842,In_496,In_1424);
nand U3843 (N_3843,In_1654,In_505);
nor U3844 (N_3844,In_2278,In_1412);
nand U3845 (N_3845,In_1240,In_2422);
and U3846 (N_3846,In_283,In_1544);
or U3847 (N_3847,In_1346,In_2223);
xor U3848 (N_3848,In_1611,In_2240);
nand U3849 (N_3849,In_879,In_868);
or U3850 (N_3850,In_1747,In_931);
nand U3851 (N_3851,In_1716,In_314);
nand U3852 (N_3852,In_2394,In_727);
nor U3853 (N_3853,In_2325,In_2328);
or U3854 (N_3854,In_210,In_1819);
and U3855 (N_3855,In_2152,In_246);
or U3856 (N_3856,In_576,In_265);
xor U3857 (N_3857,In_2046,In_1260);
xor U3858 (N_3858,In_404,In_1694);
or U3859 (N_3859,In_2427,In_1023);
xnor U3860 (N_3860,In_757,In_131);
and U3861 (N_3861,In_1992,In_1499);
nand U3862 (N_3862,In_2490,In_439);
nand U3863 (N_3863,In_1312,In_123);
or U3864 (N_3864,In_1657,In_2175);
and U3865 (N_3865,In_1355,In_1252);
nand U3866 (N_3866,In_959,In_2101);
nor U3867 (N_3867,In_597,In_1718);
and U3868 (N_3868,In_106,In_317);
and U3869 (N_3869,In_1395,In_1524);
nand U3870 (N_3870,In_2198,In_518);
and U3871 (N_3871,In_259,In_2261);
nor U3872 (N_3872,In_1477,In_191);
or U3873 (N_3873,In_2384,In_2175);
or U3874 (N_3874,In_2020,In_130);
and U3875 (N_3875,In_767,In_2456);
xor U3876 (N_3876,In_478,In_1580);
or U3877 (N_3877,In_2282,In_1449);
xnor U3878 (N_3878,In_1396,In_376);
and U3879 (N_3879,In_929,In_2074);
or U3880 (N_3880,In_112,In_1463);
nand U3881 (N_3881,In_1853,In_916);
nor U3882 (N_3882,In_788,In_2286);
nand U3883 (N_3883,In_1101,In_172);
or U3884 (N_3884,In_1654,In_432);
and U3885 (N_3885,In_1659,In_196);
and U3886 (N_3886,In_441,In_491);
nor U3887 (N_3887,In_2469,In_978);
nand U3888 (N_3888,In_1234,In_2303);
nand U3889 (N_3889,In_121,In_2140);
or U3890 (N_3890,In_312,In_1268);
or U3891 (N_3891,In_964,In_2326);
and U3892 (N_3892,In_415,In_271);
nor U3893 (N_3893,In_643,In_80);
nor U3894 (N_3894,In_2128,In_2203);
xor U3895 (N_3895,In_936,In_1916);
and U3896 (N_3896,In_2394,In_795);
xnor U3897 (N_3897,In_601,In_1732);
xor U3898 (N_3898,In_159,In_237);
or U3899 (N_3899,In_402,In_70);
nand U3900 (N_3900,In_296,In_947);
and U3901 (N_3901,In_2039,In_1443);
nand U3902 (N_3902,In_83,In_278);
nor U3903 (N_3903,In_1909,In_1541);
nand U3904 (N_3904,In_702,In_1898);
xnor U3905 (N_3905,In_638,In_1682);
nand U3906 (N_3906,In_883,In_1126);
or U3907 (N_3907,In_952,In_2022);
nor U3908 (N_3908,In_403,In_513);
nor U3909 (N_3909,In_2428,In_1025);
and U3910 (N_3910,In_568,In_2015);
nor U3911 (N_3911,In_1170,In_1952);
and U3912 (N_3912,In_1440,In_1912);
xnor U3913 (N_3913,In_1514,In_2307);
or U3914 (N_3914,In_1354,In_1991);
xor U3915 (N_3915,In_1670,In_756);
and U3916 (N_3916,In_2252,In_683);
nand U3917 (N_3917,In_1725,In_302);
and U3918 (N_3918,In_948,In_688);
or U3919 (N_3919,In_1542,In_742);
or U3920 (N_3920,In_1933,In_512);
nor U3921 (N_3921,In_1276,In_252);
nand U3922 (N_3922,In_1384,In_59);
and U3923 (N_3923,In_277,In_433);
nand U3924 (N_3924,In_1115,In_1168);
and U3925 (N_3925,In_1191,In_761);
nor U3926 (N_3926,In_1508,In_112);
and U3927 (N_3927,In_1333,In_2084);
and U3928 (N_3928,In_85,In_1049);
nand U3929 (N_3929,In_1897,In_2487);
or U3930 (N_3930,In_810,In_1379);
xor U3931 (N_3931,In_1713,In_35);
or U3932 (N_3932,In_947,In_560);
nor U3933 (N_3933,In_1354,In_1449);
or U3934 (N_3934,In_753,In_1903);
nor U3935 (N_3935,In_96,In_1677);
or U3936 (N_3936,In_1364,In_2078);
nand U3937 (N_3937,In_544,In_840);
nor U3938 (N_3938,In_130,In_2477);
and U3939 (N_3939,In_2296,In_2486);
nand U3940 (N_3940,In_1006,In_1553);
xor U3941 (N_3941,In_607,In_1384);
and U3942 (N_3942,In_402,In_837);
or U3943 (N_3943,In_1989,In_540);
xor U3944 (N_3944,In_1445,In_1199);
nand U3945 (N_3945,In_1116,In_581);
nor U3946 (N_3946,In_1882,In_81);
or U3947 (N_3947,In_172,In_1144);
nand U3948 (N_3948,In_593,In_1007);
nor U3949 (N_3949,In_1944,In_888);
and U3950 (N_3950,In_1491,In_2065);
or U3951 (N_3951,In_92,In_274);
nand U3952 (N_3952,In_584,In_277);
or U3953 (N_3953,In_1632,In_1065);
and U3954 (N_3954,In_635,In_1435);
and U3955 (N_3955,In_1025,In_568);
or U3956 (N_3956,In_1455,In_2428);
nor U3957 (N_3957,In_1550,In_1182);
nor U3958 (N_3958,In_777,In_2432);
or U3959 (N_3959,In_2471,In_391);
nand U3960 (N_3960,In_1337,In_145);
nand U3961 (N_3961,In_592,In_74);
nand U3962 (N_3962,In_2155,In_825);
or U3963 (N_3963,In_1383,In_1224);
nand U3964 (N_3964,In_1051,In_479);
and U3965 (N_3965,In_390,In_2461);
nor U3966 (N_3966,In_623,In_1157);
or U3967 (N_3967,In_14,In_1705);
nor U3968 (N_3968,In_1272,In_1885);
nand U3969 (N_3969,In_2429,In_381);
nor U3970 (N_3970,In_2388,In_1155);
nand U3971 (N_3971,In_2005,In_2349);
or U3972 (N_3972,In_689,In_1046);
xor U3973 (N_3973,In_1839,In_1189);
nor U3974 (N_3974,In_1386,In_907);
xor U3975 (N_3975,In_1664,In_1394);
or U3976 (N_3976,In_347,In_1759);
or U3977 (N_3977,In_587,In_1081);
and U3978 (N_3978,In_2434,In_632);
nor U3979 (N_3979,In_1947,In_2375);
xor U3980 (N_3980,In_289,In_1972);
or U3981 (N_3981,In_266,In_1027);
or U3982 (N_3982,In_85,In_1251);
nand U3983 (N_3983,In_2262,In_366);
or U3984 (N_3984,In_1796,In_216);
xor U3985 (N_3985,In_474,In_538);
nor U3986 (N_3986,In_905,In_147);
and U3987 (N_3987,In_140,In_2317);
and U3988 (N_3988,In_1503,In_220);
xor U3989 (N_3989,In_720,In_180);
nor U3990 (N_3990,In_1280,In_468);
and U3991 (N_3991,In_78,In_1914);
nand U3992 (N_3992,In_1247,In_730);
nor U3993 (N_3993,In_2209,In_1507);
nor U3994 (N_3994,In_704,In_1293);
nand U3995 (N_3995,In_1618,In_887);
nand U3996 (N_3996,In_1034,In_884);
xor U3997 (N_3997,In_2137,In_2488);
and U3998 (N_3998,In_458,In_604);
and U3999 (N_3999,In_740,In_2401);
nor U4000 (N_4000,In_1641,In_1284);
or U4001 (N_4001,In_673,In_2014);
nand U4002 (N_4002,In_1739,In_1848);
or U4003 (N_4003,In_309,In_2452);
nand U4004 (N_4004,In_985,In_1067);
nor U4005 (N_4005,In_458,In_2111);
nand U4006 (N_4006,In_805,In_1498);
xnor U4007 (N_4007,In_1977,In_1831);
and U4008 (N_4008,In_1207,In_824);
nand U4009 (N_4009,In_776,In_1214);
nor U4010 (N_4010,In_699,In_1325);
or U4011 (N_4011,In_2413,In_2176);
nand U4012 (N_4012,In_2249,In_1918);
nor U4013 (N_4013,In_1046,In_1684);
or U4014 (N_4014,In_2137,In_1813);
xor U4015 (N_4015,In_965,In_799);
nor U4016 (N_4016,In_314,In_1915);
nor U4017 (N_4017,In_711,In_1031);
nand U4018 (N_4018,In_1115,In_2103);
or U4019 (N_4019,In_2189,In_1914);
or U4020 (N_4020,In_1412,In_1293);
nor U4021 (N_4021,In_846,In_395);
xor U4022 (N_4022,In_1690,In_790);
nand U4023 (N_4023,In_1347,In_1506);
nor U4024 (N_4024,In_922,In_929);
nand U4025 (N_4025,In_1420,In_212);
nor U4026 (N_4026,In_226,In_385);
and U4027 (N_4027,In_1165,In_1444);
or U4028 (N_4028,In_2495,In_1202);
and U4029 (N_4029,In_269,In_445);
and U4030 (N_4030,In_57,In_728);
nor U4031 (N_4031,In_1852,In_2427);
nor U4032 (N_4032,In_1154,In_1730);
and U4033 (N_4033,In_2173,In_186);
nor U4034 (N_4034,In_313,In_2210);
nand U4035 (N_4035,In_1297,In_1609);
nand U4036 (N_4036,In_600,In_2456);
nand U4037 (N_4037,In_1650,In_887);
nor U4038 (N_4038,In_504,In_1834);
nor U4039 (N_4039,In_130,In_746);
and U4040 (N_4040,In_2270,In_2306);
xnor U4041 (N_4041,In_1118,In_361);
nand U4042 (N_4042,In_872,In_1164);
and U4043 (N_4043,In_2110,In_1175);
and U4044 (N_4044,In_748,In_359);
and U4045 (N_4045,In_1174,In_989);
or U4046 (N_4046,In_1201,In_1122);
and U4047 (N_4047,In_183,In_1043);
or U4048 (N_4048,In_2016,In_2126);
or U4049 (N_4049,In_508,In_512);
or U4050 (N_4050,In_2118,In_189);
nand U4051 (N_4051,In_1925,In_1151);
and U4052 (N_4052,In_62,In_1047);
and U4053 (N_4053,In_2405,In_799);
nand U4054 (N_4054,In_2440,In_1628);
and U4055 (N_4055,In_623,In_2318);
nand U4056 (N_4056,In_798,In_684);
nor U4057 (N_4057,In_1472,In_204);
nand U4058 (N_4058,In_1936,In_1384);
or U4059 (N_4059,In_1605,In_2020);
and U4060 (N_4060,In_1329,In_1270);
nand U4061 (N_4061,In_1828,In_1772);
nand U4062 (N_4062,In_455,In_734);
or U4063 (N_4063,In_480,In_235);
nand U4064 (N_4064,In_41,In_1643);
and U4065 (N_4065,In_537,In_115);
nor U4066 (N_4066,In_254,In_1450);
or U4067 (N_4067,In_764,In_143);
or U4068 (N_4068,In_242,In_835);
or U4069 (N_4069,In_846,In_2311);
and U4070 (N_4070,In_2405,In_341);
or U4071 (N_4071,In_1345,In_1472);
nand U4072 (N_4072,In_2324,In_2483);
nand U4073 (N_4073,In_1168,In_1747);
and U4074 (N_4074,In_1981,In_918);
or U4075 (N_4075,In_1415,In_1645);
nor U4076 (N_4076,In_2320,In_2442);
nor U4077 (N_4077,In_1794,In_83);
or U4078 (N_4078,In_990,In_1752);
or U4079 (N_4079,In_2256,In_2189);
nand U4080 (N_4080,In_2147,In_1781);
or U4081 (N_4081,In_582,In_240);
or U4082 (N_4082,In_2069,In_47);
and U4083 (N_4083,In_682,In_605);
xor U4084 (N_4084,In_364,In_822);
and U4085 (N_4085,In_1931,In_69);
and U4086 (N_4086,In_71,In_1732);
nor U4087 (N_4087,In_803,In_2484);
or U4088 (N_4088,In_1403,In_1769);
or U4089 (N_4089,In_237,In_241);
and U4090 (N_4090,In_212,In_2095);
nor U4091 (N_4091,In_1149,In_1133);
or U4092 (N_4092,In_78,In_1404);
nand U4093 (N_4093,In_1925,In_219);
and U4094 (N_4094,In_294,In_411);
nand U4095 (N_4095,In_1267,In_933);
nor U4096 (N_4096,In_2396,In_1233);
and U4097 (N_4097,In_991,In_1520);
nor U4098 (N_4098,In_1165,In_1699);
and U4099 (N_4099,In_2053,In_255);
and U4100 (N_4100,In_1126,In_956);
or U4101 (N_4101,In_617,In_636);
and U4102 (N_4102,In_370,In_124);
nand U4103 (N_4103,In_709,In_2368);
nand U4104 (N_4104,In_1051,In_1621);
and U4105 (N_4105,In_1323,In_411);
and U4106 (N_4106,In_393,In_1526);
nor U4107 (N_4107,In_929,In_1007);
and U4108 (N_4108,In_583,In_1518);
or U4109 (N_4109,In_2114,In_1576);
and U4110 (N_4110,In_1420,In_2375);
and U4111 (N_4111,In_1955,In_459);
and U4112 (N_4112,In_2242,In_1157);
and U4113 (N_4113,In_2228,In_384);
nand U4114 (N_4114,In_1694,In_974);
nor U4115 (N_4115,In_1301,In_2035);
or U4116 (N_4116,In_1331,In_1261);
and U4117 (N_4117,In_1311,In_1432);
or U4118 (N_4118,In_2418,In_2443);
nand U4119 (N_4119,In_2304,In_161);
or U4120 (N_4120,In_1182,In_1798);
nand U4121 (N_4121,In_868,In_2337);
nor U4122 (N_4122,In_323,In_617);
nor U4123 (N_4123,In_1540,In_2041);
xnor U4124 (N_4124,In_739,In_1564);
or U4125 (N_4125,In_1474,In_2427);
and U4126 (N_4126,In_1534,In_874);
and U4127 (N_4127,In_650,In_1740);
nand U4128 (N_4128,In_2276,In_1907);
nor U4129 (N_4129,In_1088,In_1835);
nand U4130 (N_4130,In_141,In_1557);
or U4131 (N_4131,In_724,In_173);
and U4132 (N_4132,In_534,In_1962);
nor U4133 (N_4133,In_504,In_1779);
nand U4134 (N_4134,In_1698,In_173);
and U4135 (N_4135,In_1975,In_1053);
and U4136 (N_4136,In_2492,In_966);
or U4137 (N_4137,In_2178,In_2125);
and U4138 (N_4138,In_346,In_2255);
xor U4139 (N_4139,In_698,In_815);
nor U4140 (N_4140,In_1396,In_711);
nand U4141 (N_4141,In_1909,In_1561);
nand U4142 (N_4142,In_1922,In_2331);
or U4143 (N_4143,In_885,In_2232);
or U4144 (N_4144,In_2179,In_382);
or U4145 (N_4145,In_1099,In_1137);
nor U4146 (N_4146,In_1098,In_2453);
or U4147 (N_4147,In_878,In_1799);
nor U4148 (N_4148,In_1463,In_2207);
or U4149 (N_4149,In_1611,In_2479);
xnor U4150 (N_4150,In_2201,In_172);
xor U4151 (N_4151,In_308,In_1841);
or U4152 (N_4152,In_1885,In_2161);
and U4153 (N_4153,In_550,In_541);
or U4154 (N_4154,In_581,In_2468);
nand U4155 (N_4155,In_1466,In_1422);
and U4156 (N_4156,In_1917,In_1560);
or U4157 (N_4157,In_1156,In_1378);
nor U4158 (N_4158,In_374,In_1122);
xnor U4159 (N_4159,In_2070,In_1718);
xor U4160 (N_4160,In_1193,In_1236);
nor U4161 (N_4161,In_2458,In_115);
nor U4162 (N_4162,In_1417,In_381);
and U4163 (N_4163,In_734,In_2148);
nor U4164 (N_4164,In_329,In_2180);
nor U4165 (N_4165,In_1575,In_978);
or U4166 (N_4166,In_1452,In_240);
nor U4167 (N_4167,In_1548,In_1400);
and U4168 (N_4168,In_185,In_1271);
xnor U4169 (N_4169,In_796,In_1967);
nand U4170 (N_4170,In_260,In_2046);
nor U4171 (N_4171,In_447,In_63);
nor U4172 (N_4172,In_634,In_649);
nand U4173 (N_4173,In_2396,In_997);
and U4174 (N_4174,In_54,In_1738);
and U4175 (N_4175,In_216,In_623);
and U4176 (N_4176,In_1616,In_152);
or U4177 (N_4177,In_1258,In_801);
nand U4178 (N_4178,In_1600,In_2000);
nor U4179 (N_4179,In_1919,In_1432);
nand U4180 (N_4180,In_1227,In_943);
or U4181 (N_4181,In_1435,In_2014);
or U4182 (N_4182,In_1525,In_2098);
nand U4183 (N_4183,In_1661,In_394);
or U4184 (N_4184,In_859,In_2218);
and U4185 (N_4185,In_2254,In_1451);
and U4186 (N_4186,In_864,In_65);
nand U4187 (N_4187,In_1450,In_1081);
nor U4188 (N_4188,In_1386,In_1756);
or U4189 (N_4189,In_967,In_985);
and U4190 (N_4190,In_649,In_985);
nand U4191 (N_4191,In_15,In_1624);
and U4192 (N_4192,In_1423,In_1090);
and U4193 (N_4193,In_2251,In_2218);
nor U4194 (N_4194,In_403,In_2477);
xor U4195 (N_4195,In_1128,In_843);
nor U4196 (N_4196,In_1424,In_1111);
and U4197 (N_4197,In_2185,In_1211);
xor U4198 (N_4198,In_1586,In_635);
nand U4199 (N_4199,In_1932,In_766);
and U4200 (N_4200,In_1424,In_2072);
and U4201 (N_4201,In_1133,In_1666);
or U4202 (N_4202,In_2231,In_1169);
nand U4203 (N_4203,In_1832,In_113);
nor U4204 (N_4204,In_198,In_2354);
xor U4205 (N_4205,In_2432,In_331);
and U4206 (N_4206,In_286,In_856);
and U4207 (N_4207,In_295,In_959);
nand U4208 (N_4208,In_2024,In_633);
nand U4209 (N_4209,In_382,In_91);
nor U4210 (N_4210,In_1105,In_2129);
nand U4211 (N_4211,In_1456,In_136);
or U4212 (N_4212,In_721,In_619);
and U4213 (N_4213,In_1156,In_1859);
or U4214 (N_4214,In_2452,In_352);
nand U4215 (N_4215,In_1867,In_1274);
nand U4216 (N_4216,In_733,In_154);
or U4217 (N_4217,In_508,In_751);
and U4218 (N_4218,In_1887,In_183);
nand U4219 (N_4219,In_1171,In_2386);
and U4220 (N_4220,In_77,In_456);
nand U4221 (N_4221,In_351,In_1914);
and U4222 (N_4222,In_663,In_904);
xnor U4223 (N_4223,In_1875,In_790);
and U4224 (N_4224,In_1210,In_1670);
nand U4225 (N_4225,In_1451,In_1994);
xor U4226 (N_4226,In_551,In_2491);
and U4227 (N_4227,In_2046,In_743);
nor U4228 (N_4228,In_85,In_1529);
nor U4229 (N_4229,In_195,In_2170);
xor U4230 (N_4230,In_802,In_1425);
nand U4231 (N_4231,In_4,In_481);
and U4232 (N_4232,In_1794,In_1125);
xnor U4233 (N_4233,In_954,In_2381);
nor U4234 (N_4234,In_1946,In_2131);
nand U4235 (N_4235,In_1070,In_630);
and U4236 (N_4236,In_2300,In_1377);
and U4237 (N_4237,In_1562,In_1683);
or U4238 (N_4238,In_629,In_1559);
nand U4239 (N_4239,In_2275,In_191);
nor U4240 (N_4240,In_1220,In_1611);
and U4241 (N_4241,In_1629,In_1775);
nor U4242 (N_4242,In_1662,In_1888);
xnor U4243 (N_4243,In_2251,In_1052);
nor U4244 (N_4244,In_105,In_780);
nor U4245 (N_4245,In_1774,In_474);
and U4246 (N_4246,In_596,In_695);
nand U4247 (N_4247,In_1966,In_940);
xor U4248 (N_4248,In_2172,In_540);
nand U4249 (N_4249,In_1820,In_1411);
nand U4250 (N_4250,In_1138,In_1108);
nand U4251 (N_4251,In_1800,In_280);
or U4252 (N_4252,In_1818,In_499);
or U4253 (N_4253,In_2365,In_221);
nor U4254 (N_4254,In_537,In_1347);
and U4255 (N_4255,In_956,In_764);
nand U4256 (N_4256,In_1983,In_1706);
nor U4257 (N_4257,In_1000,In_736);
nor U4258 (N_4258,In_1518,In_184);
nor U4259 (N_4259,In_514,In_2291);
nand U4260 (N_4260,In_204,In_2390);
and U4261 (N_4261,In_1339,In_146);
nand U4262 (N_4262,In_2158,In_2173);
or U4263 (N_4263,In_1464,In_648);
and U4264 (N_4264,In_108,In_2285);
and U4265 (N_4265,In_1797,In_811);
xor U4266 (N_4266,In_1367,In_2057);
nand U4267 (N_4267,In_95,In_2196);
nand U4268 (N_4268,In_528,In_2303);
or U4269 (N_4269,In_1754,In_1440);
or U4270 (N_4270,In_2129,In_1422);
and U4271 (N_4271,In_1089,In_571);
nand U4272 (N_4272,In_1228,In_1366);
or U4273 (N_4273,In_1620,In_2466);
xnor U4274 (N_4274,In_2358,In_1706);
and U4275 (N_4275,In_1126,In_198);
xnor U4276 (N_4276,In_229,In_1578);
nand U4277 (N_4277,In_181,In_275);
and U4278 (N_4278,In_1236,In_424);
nor U4279 (N_4279,In_2497,In_1427);
nand U4280 (N_4280,In_1949,In_1556);
and U4281 (N_4281,In_959,In_1489);
xnor U4282 (N_4282,In_1656,In_145);
and U4283 (N_4283,In_1846,In_1422);
or U4284 (N_4284,In_285,In_181);
nand U4285 (N_4285,In_1287,In_2322);
xor U4286 (N_4286,In_902,In_1859);
xor U4287 (N_4287,In_1775,In_1659);
nor U4288 (N_4288,In_2325,In_1631);
nor U4289 (N_4289,In_1718,In_447);
or U4290 (N_4290,In_266,In_913);
or U4291 (N_4291,In_1645,In_1949);
and U4292 (N_4292,In_2346,In_438);
nand U4293 (N_4293,In_1514,In_516);
xnor U4294 (N_4294,In_2424,In_1010);
nand U4295 (N_4295,In_460,In_2466);
nor U4296 (N_4296,In_2167,In_428);
and U4297 (N_4297,In_9,In_13);
nand U4298 (N_4298,In_619,In_760);
or U4299 (N_4299,In_1778,In_2360);
or U4300 (N_4300,In_121,In_1496);
nor U4301 (N_4301,In_1774,In_1065);
and U4302 (N_4302,In_85,In_1071);
xor U4303 (N_4303,In_534,In_2226);
and U4304 (N_4304,In_1212,In_1035);
nor U4305 (N_4305,In_1476,In_769);
and U4306 (N_4306,In_1807,In_2109);
nor U4307 (N_4307,In_2236,In_2332);
nor U4308 (N_4308,In_113,In_1342);
or U4309 (N_4309,In_1903,In_52);
nand U4310 (N_4310,In_2341,In_565);
nand U4311 (N_4311,In_2224,In_1728);
xnor U4312 (N_4312,In_1992,In_1469);
nor U4313 (N_4313,In_465,In_209);
nand U4314 (N_4314,In_668,In_1339);
and U4315 (N_4315,In_1708,In_2125);
or U4316 (N_4316,In_675,In_127);
and U4317 (N_4317,In_1175,In_84);
or U4318 (N_4318,In_355,In_515);
and U4319 (N_4319,In_1218,In_184);
and U4320 (N_4320,In_515,In_309);
nand U4321 (N_4321,In_944,In_1325);
or U4322 (N_4322,In_406,In_978);
nor U4323 (N_4323,In_541,In_1045);
or U4324 (N_4324,In_1671,In_1121);
or U4325 (N_4325,In_1284,In_2318);
nor U4326 (N_4326,In_1633,In_2275);
or U4327 (N_4327,In_136,In_847);
or U4328 (N_4328,In_268,In_2293);
nor U4329 (N_4329,In_446,In_568);
and U4330 (N_4330,In_1889,In_346);
and U4331 (N_4331,In_2020,In_1901);
nor U4332 (N_4332,In_768,In_447);
nand U4333 (N_4333,In_2262,In_246);
nand U4334 (N_4334,In_1396,In_539);
or U4335 (N_4335,In_800,In_199);
nand U4336 (N_4336,In_2276,In_1597);
and U4337 (N_4337,In_1838,In_1268);
nor U4338 (N_4338,In_1201,In_922);
and U4339 (N_4339,In_1784,In_1626);
or U4340 (N_4340,In_321,In_680);
nand U4341 (N_4341,In_1032,In_419);
nor U4342 (N_4342,In_1782,In_65);
and U4343 (N_4343,In_267,In_656);
nand U4344 (N_4344,In_1019,In_1002);
nand U4345 (N_4345,In_1200,In_435);
nand U4346 (N_4346,In_367,In_143);
and U4347 (N_4347,In_2467,In_1203);
xnor U4348 (N_4348,In_1885,In_1643);
nand U4349 (N_4349,In_432,In_1961);
nand U4350 (N_4350,In_1009,In_512);
nand U4351 (N_4351,In_1693,In_681);
or U4352 (N_4352,In_193,In_290);
or U4353 (N_4353,In_2079,In_637);
and U4354 (N_4354,In_1100,In_991);
nand U4355 (N_4355,In_1949,In_1371);
nor U4356 (N_4356,In_502,In_1891);
nor U4357 (N_4357,In_318,In_837);
nand U4358 (N_4358,In_1856,In_238);
and U4359 (N_4359,In_1873,In_2300);
and U4360 (N_4360,In_2292,In_846);
nand U4361 (N_4361,In_264,In_647);
or U4362 (N_4362,In_14,In_963);
or U4363 (N_4363,In_2478,In_964);
and U4364 (N_4364,In_2364,In_536);
xor U4365 (N_4365,In_426,In_2474);
or U4366 (N_4366,In_1693,In_2095);
nand U4367 (N_4367,In_2034,In_790);
nor U4368 (N_4368,In_391,In_1151);
and U4369 (N_4369,In_393,In_1874);
and U4370 (N_4370,In_2267,In_1453);
xnor U4371 (N_4371,In_9,In_1210);
and U4372 (N_4372,In_363,In_1160);
and U4373 (N_4373,In_541,In_1239);
nand U4374 (N_4374,In_234,In_279);
nor U4375 (N_4375,In_1631,In_2112);
nand U4376 (N_4376,In_27,In_668);
or U4377 (N_4377,In_2025,In_1933);
nor U4378 (N_4378,In_1903,In_973);
nand U4379 (N_4379,In_704,In_1599);
nor U4380 (N_4380,In_595,In_2364);
or U4381 (N_4381,In_1304,In_2409);
nand U4382 (N_4382,In_2468,In_2001);
and U4383 (N_4383,In_1939,In_1737);
or U4384 (N_4384,In_1896,In_883);
or U4385 (N_4385,In_1103,In_1881);
and U4386 (N_4386,In_705,In_1216);
nor U4387 (N_4387,In_2125,In_1019);
nand U4388 (N_4388,In_1444,In_906);
and U4389 (N_4389,In_1725,In_1510);
xnor U4390 (N_4390,In_1932,In_1437);
and U4391 (N_4391,In_685,In_1994);
or U4392 (N_4392,In_762,In_1506);
xnor U4393 (N_4393,In_767,In_240);
or U4394 (N_4394,In_1431,In_1860);
and U4395 (N_4395,In_1629,In_1813);
xor U4396 (N_4396,In_276,In_833);
or U4397 (N_4397,In_578,In_1413);
xnor U4398 (N_4398,In_767,In_1131);
or U4399 (N_4399,In_1167,In_1689);
and U4400 (N_4400,In_1343,In_2123);
and U4401 (N_4401,In_1492,In_1645);
nand U4402 (N_4402,In_1244,In_539);
nor U4403 (N_4403,In_317,In_1913);
nor U4404 (N_4404,In_1387,In_1750);
and U4405 (N_4405,In_4,In_324);
nand U4406 (N_4406,In_1435,In_1421);
or U4407 (N_4407,In_2110,In_1818);
nor U4408 (N_4408,In_493,In_396);
or U4409 (N_4409,In_1567,In_105);
xor U4410 (N_4410,In_269,In_967);
nand U4411 (N_4411,In_602,In_1652);
xnor U4412 (N_4412,In_1241,In_770);
and U4413 (N_4413,In_1014,In_1884);
nand U4414 (N_4414,In_1801,In_1760);
and U4415 (N_4415,In_1751,In_2397);
nor U4416 (N_4416,In_521,In_634);
and U4417 (N_4417,In_2402,In_2391);
nor U4418 (N_4418,In_2227,In_2348);
or U4419 (N_4419,In_68,In_1795);
xor U4420 (N_4420,In_2065,In_1794);
nand U4421 (N_4421,In_1735,In_501);
nor U4422 (N_4422,In_870,In_822);
nor U4423 (N_4423,In_2131,In_99);
or U4424 (N_4424,In_1744,In_1529);
nor U4425 (N_4425,In_1866,In_132);
nor U4426 (N_4426,In_973,In_1191);
nor U4427 (N_4427,In_1591,In_2013);
nand U4428 (N_4428,In_2002,In_2439);
nand U4429 (N_4429,In_1300,In_1293);
or U4430 (N_4430,In_24,In_1702);
or U4431 (N_4431,In_527,In_357);
and U4432 (N_4432,In_2308,In_2148);
xnor U4433 (N_4433,In_2222,In_2435);
and U4434 (N_4434,In_1344,In_534);
and U4435 (N_4435,In_2306,In_747);
nand U4436 (N_4436,In_131,In_1880);
nor U4437 (N_4437,In_1659,In_1604);
xor U4438 (N_4438,In_2117,In_1111);
nand U4439 (N_4439,In_1935,In_1956);
nand U4440 (N_4440,In_1162,In_1927);
xor U4441 (N_4441,In_247,In_1187);
nand U4442 (N_4442,In_361,In_381);
nand U4443 (N_4443,In_1543,In_460);
and U4444 (N_4444,In_2426,In_2281);
nand U4445 (N_4445,In_1399,In_1031);
and U4446 (N_4446,In_1018,In_413);
nand U4447 (N_4447,In_1430,In_1908);
and U4448 (N_4448,In_92,In_1375);
and U4449 (N_4449,In_1101,In_1779);
or U4450 (N_4450,In_2395,In_1873);
and U4451 (N_4451,In_382,In_699);
and U4452 (N_4452,In_1244,In_416);
and U4453 (N_4453,In_1739,In_185);
or U4454 (N_4454,In_218,In_1366);
nor U4455 (N_4455,In_1195,In_2151);
nor U4456 (N_4456,In_1477,In_1519);
nand U4457 (N_4457,In_568,In_2094);
and U4458 (N_4458,In_854,In_332);
nand U4459 (N_4459,In_918,In_270);
nor U4460 (N_4460,In_1215,In_650);
nand U4461 (N_4461,In_1855,In_627);
or U4462 (N_4462,In_1026,In_1546);
or U4463 (N_4463,In_456,In_1521);
and U4464 (N_4464,In_1151,In_47);
or U4465 (N_4465,In_1985,In_2434);
and U4466 (N_4466,In_2012,In_2306);
xor U4467 (N_4467,In_256,In_1923);
or U4468 (N_4468,In_899,In_733);
and U4469 (N_4469,In_2385,In_238);
and U4470 (N_4470,In_104,In_2130);
and U4471 (N_4471,In_889,In_469);
and U4472 (N_4472,In_831,In_997);
nor U4473 (N_4473,In_159,In_559);
nand U4474 (N_4474,In_17,In_2207);
nand U4475 (N_4475,In_1610,In_1726);
nor U4476 (N_4476,In_1754,In_613);
nand U4477 (N_4477,In_1650,In_601);
and U4478 (N_4478,In_1474,In_1440);
xor U4479 (N_4479,In_897,In_1707);
or U4480 (N_4480,In_822,In_882);
nand U4481 (N_4481,In_1190,In_1197);
and U4482 (N_4482,In_1852,In_613);
nor U4483 (N_4483,In_2032,In_15);
or U4484 (N_4484,In_2160,In_2194);
nor U4485 (N_4485,In_1074,In_1896);
and U4486 (N_4486,In_877,In_1701);
nor U4487 (N_4487,In_1347,In_2335);
and U4488 (N_4488,In_2148,In_1934);
xnor U4489 (N_4489,In_547,In_900);
nand U4490 (N_4490,In_1039,In_464);
and U4491 (N_4491,In_878,In_669);
and U4492 (N_4492,In_1135,In_2029);
xor U4493 (N_4493,In_1576,In_25);
or U4494 (N_4494,In_1795,In_1175);
and U4495 (N_4495,In_1140,In_1858);
nand U4496 (N_4496,In_1315,In_2409);
nand U4497 (N_4497,In_2049,In_1055);
or U4498 (N_4498,In_2121,In_527);
nand U4499 (N_4499,In_2488,In_2097);
nor U4500 (N_4500,In_2271,In_774);
and U4501 (N_4501,In_1117,In_380);
or U4502 (N_4502,In_59,In_1542);
nand U4503 (N_4503,In_436,In_1292);
nor U4504 (N_4504,In_1871,In_2224);
and U4505 (N_4505,In_1524,In_1793);
nand U4506 (N_4506,In_2225,In_1934);
or U4507 (N_4507,In_1298,In_43);
nand U4508 (N_4508,In_461,In_430);
nor U4509 (N_4509,In_17,In_1734);
or U4510 (N_4510,In_1635,In_1723);
nor U4511 (N_4511,In_2428,In_378);
or U4512 (N_4512,In_1282,In_532);
nand U4513 (N_4513,In_1801,In_1006);
or U4514 (N_4514,In_589,In_711);
nand U4515 (N_4515,In_1452,In_191);
nand U4516 (N_4516,In_2299,In_515);
nand U4517 (N_4517,In_1647,In_2019);
xor U4518 (N_4518,In_2142,In_2389);
and U4519 (N_4519,In_1248,In_1752);
xnor U4520 (N_4520,In_376,In_1004);
or U4521 (N_4521,In_568,In_2147);
or U4522 (N_4522,In_34,In_1897);
and U4523 (N_4523,In_2397,In_1438);
nand U4524 (N_4524,In_1676,In_2197);
nor U4525 (N_4525,In_270,In_2055);
nor U4526 (N_4526,In_1162,In_174);
nor U4527 (N_4527,In_764,In_1392);
nor U4528 (N_4528,In_639,In_973);
or U4529 (N_4529,In_693,In_1025);
and U4530 (N_4530,In_2488,In_1900);
nand U4531 (N_4531,In_1485,In_1593);
or U4532 (N_4532,In_1858,In_325);
nor U4533 (N_4533,In_1309,In_1231);
nand U4534 (N_4534,In_888,In_849);
nor U4535 (N_4535,In_576,In_2055);
nor U4536 (N_4536,In_1020,In_1683);
or U4537 (N_4537,In_1134,In_1721);
nand U4538 (N_4538,In_515,In_1295);
or U4539 (N_4539,In_666,In_929);
xor U4540 (N_4540,In_2320,In_1860);
nor U4541 (N_4541,In_2302,In_713);
nor U4542 (N_4542,In_2476,In_713);
nand U4543 (N_4543,In_1209,In_996);
and U4544 (N_4544,In_1683,In_1272);
nor U4545 (N_4545,In_2078,In_1667);
nor U4546 (N_4546,In_57,In_575);
or U4547 (N_4547,In_165,In_693);
nor U4548 (N_4548,In_1949,In_2439);
or U4549 (N_4549,In_1617,In_1963);
or U4550 (N_4550,In_1019,In_1849);
xnor U4551 (N_4551,In_2138,In_2424);
nor U4552 (N_4552,In_1148,In_2278);
nand U4553 (N_4553,In_284,In_1494);
nor U4554 (N_4554,In_45,In_2184);
xor U4555 (N_4555,In_1846,In_1283);
nand U4556 (N_4556,In_53,In_681);
nor U4557 (N_4557,In_2147,In_1289);
or U4558 (N_4558,In_1343,In_1137);
and U4559 (N_4559,In_2240,In_1718);
and U4560 (N_4560,In_889,In_1524);
xor U4561 (N_4561,In_2135,In_505);
and U4562 (N_4562,In_1075,In_1396);
or U4563 (N_4563,In_1701,In_2097);
nor U4564 (N_4564,In_2187,In_1324);
nand U4565 (N_4565,In_1491,In_757);
nand U4566 (N_4566,In_551,In_359);
and U4567 (N_4567,In_45,In_322);
nor U4568 (N_4568,In_1801,In_1641);
nor U4569 (N_4569,In_2242,In_2449);
nand U4570 (N_4570,In_2182,In_851);
xor U4571 (N_4571,In_2156,In_1824);
and U4572 (N_4572,In_1719,In_1965);
or U4573 (N_4573,In_1305,In_2122);
nor U4574 (N_4574,In_899,In_1265);
nand U4575 (N_4575,In_1392,In_733);
or U4576 (N_4576,In_1214,In_1215);
and U4577 (N_4577,In_1570,In_222);
and U4578 (N_4578,In_2146,In_2487);
nor U4579 (N_4579,In_2038,In_1381);
nor U4580 (N_4580,In_2397,In_2137);
nor U4581 (N_4581,In_193,In_441);
nor U4582 (N_4582,In_2079,In_904);
nand U4583 (N_4583,In_2050,In_1048);
and U4584 (N_4584,In_1135,In_299);
nand U4585 (N_4585,In_2012,In_904);
and U4586 (N_4586,In_222,In_1536);
nor U4587 (N_4587,In_529,In_919);
nand U4588 (N_4588,In_1602,In_2267);
nor U4589 (N_4589,In_1662,In_2316);
nand U4590 (N_4590,In_747,In_1423);
nand U4591 (N_4591,In_1299,In_315);
or U4592 (N_4592,In_1417,In_1632);
or U4593 (N_4593,In_1046,In_889);
nand U4594 (N_4594,In_1239,In_1315);
or U4595 (N_4595,In_479,In_272);
nor U4596 (N_4596,In_174,In_1439);
nor U4597 (N_4597,In_1414,In_319);
and U4598 (N_4598,In_1080,In_114);
nand U4599 (N_4599,In_897,In_1395);
nor U4600 (N_4600,In_956,In_1367);
nor U4601 (N_4601,In_828,In_1842);
or U4602 (N_4602,In_1501,In_1981);
and U4603 (N_4603,In_1028,In_1314);
or U4604 (N_4604,In_1709,In_517);
nand U4605 (N_4605,In_2275,In_345);
nor U4606 (N_4606,In_433,In_216);
nand U4607 (N_4607,In_1048,In_912);
nand U4608 (N_4608,In_1735,In_2009);
nor U4609 (N_4609,In_1531,In_343);
and U4610 (N_4610,In_732,In_1948);
or U4611 (N_4611,In_152,In_256);
nand U4612 (N_4612,In_1645,In_293);
xnor U4613 (N_4613,In_2255,In_1786);
and U4614 (N_4614,In_1573,In_462);
nor U4615 (N_4615,In_538,In_40);
or U4616 (N_4616,In_1847,In_1421);
or U4617 (N_4617,In_2016,In_1985);
nand U4618 (N_4618,In_1858,In_2468);
nor U4619 (N_4619,In_1297,In_1819);
and U4620 (N_4620,In_1226,In_335);
nand U4621 (N_4621,In_1376,In_2343);
and U4622 (N_4622,In_2310,In_2087);
or U4623 (N_4623,In_524,In_14);
or U4624 (N_4624,In_291,In_2426);
or U4625 (N_4625,In_858,In_325);
nor U4626 (N_4626,In_1221,In_1688);
nand U4627 (N_4627,In_159,In_651);
or U4628 (N_4628,In_300,In_2008);
nor U4629 (N_4629,In_880,In_1687);
nor U4630 (N_4630,In_2277,In_1773);
xor U4631 (N_4631,In_41,In_1850);
nor U4632 (N_4632,In_2159,In_559);
nand U4633 (N_4633,In_1260,In_805);
nand U4634 (N_4634,In_1074,In_1132);
xnor U4635 (N_4635,In_1239,In_1536);
and U4636 (N_4636,In_1602,In_1749);
and U4637 (N_4637,In_2408,In_1190);
nor U4638 (N_4638,In_514,In_1773);
and U4639 (N_4639,In_1712,In_2492);
nor U4640 (N_4640,In_1583,In_566);
nor U4641 (N_4641,In_1117,In_1564);
or U4642 (N_4642,In_947,In_421);
nand U4643 (N_4643,In_2265,In_2114);
and U4644 (N_4644,In_2026,In_2049);
or U4645 (N_4645,In_39,In_183);
or U4646 (N_4646,In_327,In_2047);
nand U4647 (N_4647,In_1392,In_1043);
nand U4648 (N_4648,In_2418,In_1813);
nor U4649 (N_4649,In_2004,In_776);
or U4650 (N_4650,In_2020,In_1492);
xnor U4651 (N_4651,In_530,In_1205);
and U4652 (N_4652,In_1458,In_1911);
nand U4653 (N_4653,In_1783,In_2424);
or U4654 (N_4654,In_722,In_334);
and U4655 (N_4655,In_1672,In_612);
and U4656 (N_4656,In_2303,In_1637);
nand U4657 (N_4657,In_640,In_1036);
or U4658 (N_4658,In_1151,In_1264);
nor U4659 (N_4659,In_201,In_1496);
nand U4660 (N_4660,In_1042,In_1052);
and U4661 (N_4661,In_268,In_2158);
or U4662 (N_4662,In_1813,In_466);
nor U4663 (N_4663,In_2031,In_1706);
and U4664 (N_4664,In_1720,In_802);
or U4665 (N_4665,In_301,In_442);
nor U4666 (N_4666,In_2318,In_1992);
or U4667 (N_4667,In_1047,In_1483);
and U4668 (N_4668,In_433,In_1875);
or U4669 (N_4669,In_186,In_1292);
nor U4670 (N_4670,In_1153,In_1473);
or U4671 (N_4671,In_1467,In_2207);
nor U4672 (N_4672,In_1263,In_2489);
nor U4673 (N_4673,In_2354,In_108);
nor U4674 (N_4674,In_351,In_1745);
nor U4675 (N_4675,In_1037,In_1943);
or U4676 (N_4676,In_1444,In_1841);
nor U4677 (N_4677,In_2401,In_443);
nand U4678 (N_4678,In_664,In_205);
and U4679 (N_4679,In_108,In_640);
and U4680 (N_4680,In_1677,In_1638);
xor U4681 (N_4681,In_2070,In_1642);
nor U4682 (N_4682,In_1065,In_1613);
or U4683 (N_4683,In_1781,In_623);
and U4684 (N_4684,In_1980,In_481);
nor U4685 (N_4685,In_759,In_575);
nand U4686 (N_4686,In_1668,In_571);
nor U4687 (N_4687,In_1869,In_1745);
xnor U4688 (N_4688,In_572,In_1049);
xor U4689 (N_4689,In_60,In_118);
or U4690 (N_4690,In_2097,In_2125);
nand U4691 (N_4691,In_1802,In_1238);
or U4692 (N_4692,In_2464,In_2189);
nand U4693 (N_4693,In_186,In_659);
nor U4694 (N_4694,In_398,In_1423);
nor U4695 (N_4695,In_426,In_419);
or U4696 (N_4696,In_2215,In_2314);
or U4697 (N_4697,In_804,In_701);
or U4698 (N_4698,In_2253,In_193);
nor U4699 (N_4699,In_1328,In_1066);
xor U4700 (N_4700,In_2404,In_2034);
xnor U4701 (N_4701,In_2448,In_456);
nor U4702 (N_4702,In_10,In_2162);
nand U4703 (N_4703,In_786,In_1736);
nand U4704 (N_4704,In_1682,In_1535);
nor U4705 (N_4705,In_369,In_1003);
and U4706 (N_4706,In_2168,In_1628);
or U4707 (N_4707,In_2254,In_1154);
nand U4708 (N_4708,In_926,In_1686);
nor U4709 (N_4709,In_425,In_1360);
nand U4710 (N_4710,In_1771,In_1730);
or U4711 (N_4711,In_656,In_1334);
or U4712 (N_4712,In_726,In_847);
xor U4713 (N_4713,In_1800,In_2296);
nand U4714 (N_4714,In_2187,In_1670);
or U4715 (N_4715,In_510,In_1770);
nor U4716 (N_4716,In_170,In_605);
nand U4717 (N_4717,In_1233,In_1065);
or U4718 (N_4718,In_99,In_479);
nor U4719 (N_4719,In_171,In_1201);
and U4720 (N_4720,In_1953,In_1279);
nor U4721 (N_4721,In_2422,In_73);
xor U4722 (N_4722,In_228,In_2053);
or U4723 (N_4723,In_2482,In_1085);
nand U4724 (N_4724,In_2338,In_961);
nor U4725 (N_4725,In_2181,In_608);
xor U4726 (N_4726,In_1346,In_201);
and U4727 (N_4727,In_1612,In_737);
and U4728 (N_4728,In_2152,In_1367);
and U4729 (N_4729,In_1098,In_2356);
or U4730 (N_4730,In_1206,In_1527);
nor U4731 (N_4731,In_2322,In_2067);
or U4732 (N_4732,In_547,In_59);
or U4733 (N_4733,In_2333,In_1338);
xor U4734 (N_4734,In_76,In_943);
xor U4735 (N_4735,In_790,In_1560);
xor U4736 (N_4736,In_904,In_620);
nand U4737 (N_4737,In_1765,In_1363);
nor U4738 (N_4738,In_887,In_417);
and U4739 (N_4739,In_362,In_949);
or U4740 (N_4740,In_2483,In_496);
nor U4741 (N_4741,In_1406,In_204);
nor U4742 (N_4742,In_1109,In_1552);
and U4743 (N_4743,In_1005,In_660);
xor U4744 (N_4744,In_2000,In_2034);
xnor U4745 (N_4745,In_1170,In_510);
and U4746 (N_4746,In_1607,In_1664);
or U4747 (N_4747,In_901,In_1649);
xnor U4748 (N_4748,In_853,In_2247);
or U4749 (N_4749,In_1014,In_1365);
nand U4750 (N_4750,In_1235,In_100);
xnor U4751 (N_4751,In_141,In_2470);
nand U4752 (N_4752,In_2379,In_1900);
nor U4753 (N_4753,In_1401,In_1479);
nand U4754 (N_4754,In_2204,In_31);
xor U4755 (N_4755,In_965,In_1006);
and U4756 (N_4756,In_2362,In_103);
nand U4757 (N_4757,In_478,In_786);
nor U4758 (N_4758,In_1482,In_982);
and U4759 (N_4759,In_2262,In_1947);
and U4760 (N_4760,In_1135,In_534);
or U4761 (N_4761,In_1933,In_736);
or U4762 (N_4762,In_12,In_2066);
xnor U4763 (N_4763,In_1142,In_1190);
and U4764 (N_4764,In_263,In_1789);
and U4765 (N_4765,In_2193,In_2274);
or U4766 (N_4766,In_688,In_76);
nand U4767 (N_4767,In_924,In_213);
and U4768 (N_4768,In_1180,In_6);
or U4769 (N_4769,In_2488,In_2285);
nor U4770 (N_4770,In_1974,In_1690);
or U4771 (N_4771,In_185,In_882);
and U4772 (N_4772,In_1948,In_310);
or U4773 (N_4773,In_2038,In_2447);
and U4774 (N_4774,In_2003,In_322);
xor U4775 (N_4775,In_2168,In_2203);
and U4776 (N_4776,In_180,In_589);
and U4777 (N_4777,In_1687,In_1149);
or U4778 (N_4778,In_1616,In_739);
nor U4779 (N_4779,In_1373,In_925);
xor U4780 (N_4780,In_1640,In_196);
and U4781 (N_4781,In_1982,In_6);
or U4782 (N_4782,In_244,In_536);
or U4783 (N_4783,In_1440,In_1622);
nand U4784 (N_4784,In_1387,In_138);
nand U4785 (N_4785,In_2031,In_834);
nand U4786 (N_4786,In_1261,In_2325);
and U4787 (N_4787,In_2242,In_1971);
nor U4788 (N_4788,In_2359,In_879);
or U4789 (N_4789,In_796,In_450);
or U4790 (N_4790,In_1634,In_1659);
xor U4791 (N_4791,In_647,In_1570);
nand U4792 (N_4792,In_2253,In_1362);
and U4793 (N_4793,In_1507,In_790);
nor U4794 (N_4794,In_573,In_2112);
nor U4795 (N_4795,In_1021,In_1776);
or U4796 (N_4796,In_348,In_1740);
or U4797 (N_4797,In_146,In_2053);
nand U4798 (N_4798,In_497,In_546);
or U4799 (N_4799,In_838,In_2274);
and U4800 (N_4800,In_996,In_83);
xor U4801 (N_4801,In_102,In_77);
xnor U4802 (N_4802,In_393,In_91);
xnor U4803 (N_4803,In_918,In_325);
nand U4804 (N_4804,In_1748,In_1689);
and U4805 (N_4805,In_989,In_296);
and U4806 (N_4806,In_2212,In_295);
nand U4807 (N_4807,In_2318,In_609);
nand U4808 (N_4808,In_697,In_223);
nand U4809 (N_4809,In_1513,In_1922);
nand U4810 (N_4810,In_1490,In_419);
xnor U4811 (N_4811,In_1110,In_375);
or U4812 (N_4812,In_421,In_2350);
nor U4813 (N_4813,In_428,In_1737);
nand U4814 (N_4814,In_2206,In_1678);
nand U4815 (N_4815,In_1109,In_1643);
and U4816 (N_4816,In_1121,In_1841);
and U4817 (N_4817,In_888,In_1679);
and U4818 (N_4818,In_521,In_2490);
or U4819 (N_4819,In_2466,In_2332);
or U4820 (N_4820,In_821,In_418);
or U4821 (N_4821,In_33,In_1992);
nor U4822 (N_4822,In_931,In_982);
nand U4823 (N_4823,In_1423,In_1913);
nor U4824 (N_4824,In_2494,In_1038);
nand U4825 (N_4825,In_470,In_201);
or U4826 (N_4826,In_1565,In_1136);
xor U4827 (N_4827,In_1810,In_1149);
and U4828 (N_4828,In_54,In_2182);
xnor U4829 (N_4829,In_1050,In_1184);
nor U4830 (N_4830,In_1079,In_349);
nand U4831 (N_4831,In_427,In_878);
nor U4832 (N_4832,In_13,In_2259);
and U4833 (N_4833,In_2235,In_594);
nand U4834 (N_4834,In_1936,In_664);
nand U4835 (N_4835,In_1442,In_1810);
nor U4836 (N_4836,In_2405,In_1022);
nand U4837 (N_4837,In_1301,In_392);
and U4838 (N_4838,In_464,In_2463);
or U4839 (N_4839,In_1472,In_2438);
and U4840 (N_4840,In_257,In_501);
or U4841 (N_4841,In_1641,In_642);
xor U4842 (N_4842,In_166,In_203);
nor U4843 (N_4843,In_2030,In_755);
or U4844 (N_4844,In_91,In_695);
or U4845 (N_4845,In_1778,In_1327);
nor U4846 (N_4846,In_2435,In_292);
nand U4847 (N_4847,In_2473,In_1783);
nor U4848 (N_4848,In_812,In_1572);
nor U4849 (N_4849,In_2340,In_798);
and U4850 (N_4850,In_1766,In_2228);
nor U4851 (N_4851,In_2384,In_1530);
nor U4852 (N_4852,In_373,In_303);
or U4853 (N_4853,In_1762,In_834);
or U4854 (N_4854,In_1544,In_1484);
or U4855 (N_4855,In_1388,In_1714);
nor U4856 (N_4856,In_1539,In_1196);
or U4857 (N_4857,In_606,In_2494);
nand U4858 (N_4858,In_1204,In_1720);
and U4859 (N_4859,In_663,In_107);
nor U4860 (N_4860,In_164,In_2327);
nand U4861 (N_4861,In_1240,In_1498);
nand U4862 (N_4862,In_1419,In_508);
nand U4863 (N_4863,In_1048,In_1490);
nand U4864 (N_4864,In_1659,In_533);
xor U4865 (N_4865,In_1696,In_2212);
or U4866 (N_4866,In_1634,In_38);
or U4867 (N_4867,In_132,In_1011);
nor U4868 (N_4868,In_984,In_1250);
nand U4869 (N_4869,In_56,In_2039);
nand U4870 (N_4870,In_992,In_291);
xor U4871 (N_4871,In_831,In_593);
nor U4872 (N_4872,In_1453,In_1612);
and U4873 (N_4873,In_574,In_1510);
nor U4874 (N_4874,In_1091,In_1530);
and U4875 (N_4875,In_1362,In_469);
nor U4876 (N_4876,In_442,In_539);
nor U4877 (N_4877,In_2086,In_1912);
or U4878 (N_4878,In_89,In_1440);
nand U4879 (N_4879,In_2499,In_129);
and U4880 (N_4880,In_98,In_1552);
and U4881 (N_4881,In_1409,In_1034);
and U4882 (N_4882,In_772,In_720);
or U4883 (N_4883,In_243,In_787);
nand U4884 (N_4884,In_753,In_468);
and U4885 (N_4885,In_687,In_2437);
nor U4886 (N_4886,In_794,In_871);
xnor U4887 (N_4887,In_2270,In_1345);
and U4888 (N_4888,In_1747,In_1730);
or U4889 (N_4889,In_1030,In_2219);
nor U4890 (N_4890,In_816,In_464);
or U4891 (N_4891,In_111,In_1947);
nand U4892 (N_4892,In_1149,In_856);
nor U4893 (N_4893,In_2235,In_2059);
nor U4894 (N_4894,In_1104,In_1303);
xnor U4895 (N_4895,In_1545,In_766);
nand U4896 (N_4896,In_497,In_1278);
and U4897 (N_4897,In_1949,In_2110);
nand U4898 (N_4898,In_1691,In_1886);
nand U4899 (N_4899,In_435,In_1002);
or U4900 (N_4900,In_1966,In_2220);
and U4901 (N_4901,In_158,In_361);
nand U4902 (N_4902,In_542,In_543);
and U4903 (N_4903,In_2354,In_1228);
and U4904 (N_4904,In_2284,In_811);
and U4905 (N_4905,In_2025,In_292);
and U4906 (N_4906,In_800,In_1896);
nor U4907 (N_4907,In_221,In_218);
nor U4908 (N_4908,In_1908,In_489);
and U4909 (N_4909,In_1328,In_722);
nor U4910 (N_4910,In_1734,In_1972);
nand U4911 (N_4911,In_695,In_2244);
and U4912 (N_4912,In_715,In_1007);
nor U4913 (N_4913,In_357,In_1733);
and U4914 (N_4914,In_624,In_2213);
nor U4915 (N_4915,In_1083,In_1210);
or U4916 (N_4916,In_1635,In_2469);
nand U4917 (N_4917,In_1392,In_561);
nand U4918 (N_4918,In_402,In_1665);
or U4919 (N_4919,In_1444,In_600);
nor U4920 (N_4920,In_1655,In_1519);
xnor U4921 (N_4921,In_1569,In_2438);
and U4922 (N_4922,In_583,In_2329);
and U4923 (N_4923,In_1610,In_589);
nand U4924 (N_4924,In_250,In_1375);
nor U4925 (N_4925,In_868,In_2115);
or U4926 (N_4926,In_1074,In_2318);
xnor U4927 (N_4927,In_1655,In_582);
nand U4928 (N_4928,In_1265,In_575);
or U4929 (N_4929,In_208,In_47);
or U4930 (N_4930,In_1293,In_926);
and U4931 (N_4931,In_1058,In_1741);
nor U4932 (N_4932,In_2257,In_1925);
or U4933 (N_4933,In_563,In_1639);
nand U4934 (N_4934,In_618,In_1424);
xor U4935 (N_4935,In_1855,In_1149);
nand U4936 (N_4936,In_396,In_651);
or U4937 (N_4937,In_654,In_1720);
and U4938 (N_4938,In_2195,In_2049);
nor U4939 (N_4939,In_1957,In_2184);
or U4940 (N_4940,In_2376,In_1875);
nor U4941 (N_4941,In_777,In_1861);
or U4942 (N_4942,In_1822,In_2315);
nand U4943 (N_4943,In_2243,In_1291);
or U4944 (N_4944,In_1361,In_1082);
or U4945 (N_4945,In_2024,In_2458);
nor U4946 (N_4946,In_2332,In_2039);
nand U4947 (N_4947,In_1769,In_1247);
nor U4948 (N_4948,In_630,In_1139);
and U4949 (N_4949,In_812,In_467);
or U4950 (N_4950,In_1509,In_1031);
nor U4951 (N_4951,In_2319,In_906);
or U4952 (N_4952,In_136,In_1327);
nand U4953 (N_4953,In_48,In_177);
or U4954 (N_4954,In_474,In_760);
nand U4955 (N_4955,In_93,In_1153);
nor U4956 (N_4956,In_21,In_2300);
and U4957 (N_4957,In_2223,In_661);
nor U4958 (N_4958,In_2342,In_190);
nor U4959 (N_4959,In_419,In_298);
or U4960 (N_4960,In_2213,In_1310);
nor U4961 (N_4961,In_475,In_700);
nand U4962 (N_4962,In_84,In_429);
and U4963 (N_4963,In_2226,In_1295);
xnor U4964 (N_4964,In_926,In_1065);
or U4965 (N_4965,In_885,In_824);
xor U4966 (N_4966,In_836,In_542);
nor U4967 (N_4967,In_488,In_1476);
xnor U4968 (N_4968,In_1674,In_1366);
nand U4969 (N_4969,In_2173,In_2227);
and U4970 (N_4970,In_1939,In_2467);
or U4971 (N_4971,In_2466,In_261);
nor U4972 (N_4972,In_250,In_224);
nor U4973 (N_4973,In_1416,In_2466);
or U4974 (N_4974,In_64,In_1700);
and U4975 (N_4975,In_2194,In_2207);
nand U4976 (N_4976,In_1339,In_944);
xor U4977 (N_4977,In_1313,In_410);
nand U4978 (N_4978,In_2294,In_932);
and U4979 (N_4979,In_2325,In_957);
nand U4980 (N_4980,In_2386,In_1591);
nor U4981 (N_4981,In_1978,In_2336);
xnor U4982 (N_4982,In_1737,In_1187);
or U4983 (N_4983,In_1314,In_1188);
nor U4984 (N_4984,In_144,In_2498);
xor U4985 (N_4985,In_1170,In_1835);
nor U4986 (N_4986,In_685,In_1740);
nand U4987 (N_4987,In_2402,In_1663);
nor U4988 (N_4988,In_1399,In_1923);
nor U4989 (N_4989,In_318,In_1477);
nor U4990 (N_4990,In_885,In_2226);
or U4991 (N_4991,In_824,In_1586);
or U4992 (N_4992,In_1947,In_210);
and U4993 (N_4993,In_2158,In_1972);
and U4994 (N_4994,In_1881,In_1645);
and U4995 (N_4995,In_1290,In_320);
nor U4996 (N_4996,In_222,In_1853);
xnor U4997 (N_4997,In_2348,In_963);
and U4998 (N_4998,In_140,In_50);
nand U4999 (N_4999,In_790,In_1086);
nand U5000 (N_5000,N_2463,N_4983);
nand U5001 (N_5001,N_4027,N_545);
and U5002 (N_5002,N_412,N_1055);
nor U5003 (N_5003,N_2687,N_28);
and U5004 (N_5004,N_4233,N_3625);
or U5005 (N_5005,N_4948,N_4677);
nor U5006 (N_5006,N_2068,N_3121);
nand U5007 (N_5007,N_4092,N_983);
nand U5008 (N_5008,N_674,N_1782);
or U5009 (N_5009,N_565,N_975);
nor U5010 (N_5010,N_3535,N_3876);
or U5011 (N_5011,N_680,N_3753);
and U5012 (N_5012,N_634,N_1315);
nand U5013 (N_5013,N_209,N_3691);
or U5014 (N_5014,N_2202,N_4123);
and U5015 (N_5015,N_2395,N_588);
nor U5016 (N_5016,N_93,N_225);
nand U5017 (N_5017,N_4426,N_4878);
or U5018 (N_5018,N_2679,N_2843);
nand U5019 (N_5019,N_1385,N_1103);
nor U5020 (N_5020,N_2626,N_4393);
nor U5021 (N_5021,N_4375,N_2330);
nor U5022 (N_5022,N_1423,N_560);
and U5023 (N_5023,N_197,N_3811);
nor U5024 (N_5024,N_2677,N_537);
nand U5025 (N_5025,N_2920,N_534);
and U5026 (N_5026,N_89,N_4235);
xor U5027 (N_5027,N_3032,N_1574);
nand U5028 (N_5028,N_1904,N_2266);
nor U5029 (N_5029,N_558,N_4966);
xnor U5030 (N_5030,N_3157,N_427);
nor U5031 (N_5031,N_3628,N_4111);
or U5032 (N_5032,N_2459,N_1923);
nor U5033 (N_5033,N_4640,N_2834);
nand U5034 (N_5034,N_1117,N_180);
nor U5035 (N_5035,N_1935,N_3366);
or U5036 (N_5036,N_4523,N_4729);
nand U5037 (N_5037,N_1133,N_3825);
or U5038 (N_5038,N_2225,N_2454);
or U5039 (N_5039,N_2832,N_3810);
and U5040 (N_5040,N_3562,N_2170);
or U5041 (N_5041,N_943,N_715);
or U5042 (N_5042,N_358,N_1400);
and U5043 (N_5043,N_2806,N_2224);
nand U5044 (N_5044,N_2026,N_946);
xnor U5045 (N_5045,N_4720,N_4833);
and U5046 (N_5046,N_3997,N_757);
or U5047 (N_5047,N_299,N_3508);
or U5048 (N_5048,N_2830,N_4925);
nand U5049 (N_5049,N_3679,N_440);
and U5050 (N_5050,N_3621,N_1870);
nand U5051 (N_5051,N_86,N_3724);
or U5052 (N_5052,N_2747,N_3203);
and U5053 (N_5053,N_4514,N_4324);
or U5054 (N_5054,N_1359,N_1716);
and U5055 (N_5055,N_4617,N_3960);
xor U5056 (N_5056,N_1341,N_2681);
nor U5057 (N_5057,N_1377,N_579);
nand U5058 (N_5058,N_3256,N_316);
and U5059 (N_5059,N_4278,N_442);
nor U5060 (N_5060,N_2570,N_1473);
xnor U5061 (N_5061,N_319,N_3479);
xor U5062 (N_5062,N_4127,N_2305);
and U5063 (N_5063,N_3227,N_1510);
nand U5064 (N_5064,N_3834,N_262);
and U5065 (N_5065,N_1740,N_1928);
nand U5066 (N_5066,N_3831,N_4088);
nor U5067 (N_5067,N_4089,N_1608);
and U5068 (N_5068,N_3421,N_1369);
nand U5069 (N_5069,N_3505,N_1394);
or U5070 (N_5070,N_327,N_230);
nor U5071 (N_5071,N_3352,N_4919);
nor U5072 (N_5072,N_4209,N_1409);
nor U5073 (N_5073,N_751,N_2627);
or U5074 (N_5074,N_810,N_915);
nor U5075 (N_5075,N_1166,N_3446);
and U5076 (N_5076,N_4409,N_3646);
xor U5077 (N_5077,N_1552,N_1425);
nand U5078 (N_5078,N_4718,N_4072);
or U5079 (N_5079,N_4184,N_1067);
nor U5080 (N_5080,N_1879,N_2198);
nor U5081 (N_5081,N_3852,N_232);
nor U5082 (N_5082,N_3739,N_1687);
and U5083 (N_5083,N_819,N_4544);
and U5084 (N_5084,N_1380,N_2942);
nand U5085 (N_5085,N_415,N_2961);
and U5086 (N_5086,N_4414,N_2604);
nor U5087 (N_5087,N_4230,N_1308);
nor U5088 (N_5088,N_4540,N_1407);
nand U5089 (N_5089,N_4903,N_1938);
or U5090 (N_5090,N_714,N_2204);
nor U5091 (N_5091,N_3558,N_22);
or U5092 (N_5092,N_1021,N_1666);
or U5093 (N_5093,N_4124,N_3436);
nand U5094 (N_5094,N_310,N_1154);
nand U5095 (N_5095,N_45,N_2258);
nor U5096 (N_5096,N_730,N_2800);
or U5097 (N_5097,N_1406,N_4897);
and U5098 (N_5098,N_2976,N_2409);
or U5099 (N_5099,N_581,N_1588);
nor U5100 (N_5100,N_1508,N_4328);
or U5101 (N_5101,N_1057,N_1245);
and U5102 (N_5102,N_1395,N_4570);
nand U5103 (N_5103,N_2999,N_969);
nor U5104 (N_5104,N_131,N_4562);
or U5105 (N_5105,N_864,N_2751);
nand U5106 (N_5106,N_1907,N_726);
nand U5107 (N_5107,N_1556,N_4526);
nor U5108 (N_5108,N_1399,N_2853);
or U5109 (N_5109,N_1097,N_629);
nor U5110 (N_5110,N_4013,N_2344);
nor U5111 (N_5111,N_2913,N_3941);
nand U5112 (N_5112,N_2128,N_4344);
and U5113 (N_5113,N_4338,N_4360);
and U5114 (N_5114,N_3878,N_1683);
nor U5115 (N_5115,N_638,N_2090);
nor U5116 (N_5116,N_1124,N_4527);
or U5117 (N_5117,N_1847,N_2636);
nor U5118 (N_5118,N_3861,N_995);
nand U5119 (N_5119,N_1137,N_4771);
nand U5120 (N_5120,N_3368,N_2289);
or U5121 (N_5121,N_935,N_4709);
nand U5122 (N_5122,N_2526,N_3933);
and U5123 (N_5123,N_2595,N_996);
nand U5124 (N_5124,N_1306,N_1464);
or U5125 (N_5125,N_4474,N_356);
and U5126 (N_5126,N_2172,N_2518);
xnor U5127 (N_5127,N_247,N_4790);
or U5128 (N_5128,N_3935,N_3444);
and U5129 (N_5129,N_413,N_1242);
nor U5130 (N_5130,N_833,N_1735);
and U5131 (N_5131,N_4029,N_402);
xor U5132 (N_5132,N_322,N_1271);
nor U5133 (N_5133,N_3307,N_2115);
nand U5134 (N_5134,N_2809,N_828);
and U5135 (N_5135,N_1638,N_4964);
nand U5136 (N_5136,N_1305,N_3836);
nor U5137 (N_5137,N_620,N_3394);
nand U5138 (N_5138,N_2303,N_152);
and U5139 (N_5139,N_3564,N_3439);
or U5140 (N_5140,N_1643,N_2506);
xnor U5141 (N_5141,N_4618,N_788);
nor U5142 (N_5142,N_4542,N_3419);
and U5143 (N_5143,N_676,N_3607);
and U5144 (N_5144,N_574,N_1146);
nand U5145 (N_5145,N_1728,N_863);
xor U5146 (N_5146,N_1089,N_4700);
or U5147 (N_5147,N_3962,N_4007);
nor U5148 (N_5148,N_1975,N_682);
nor U5149 (N_5149,N_4464,N_690);
nand U5150 (N_5150,N_613,N_4488);
nor U5151 (N_5151,N_792,N_1581);
nor U5152 (N_5152,N_1739,N_2150);
nor U5153 (N_5153,N_1202,N_1342);
and U5154 (N_5154,N_4877,N_1796);
xor U5155 (N_5155,N_4810,N_3703);
nor U5156 (N_5156,N_4776,N_1163);
nor U5157 (N_5157,N_4405,N_2745);
nor U5158 (N_5158,N_2455,N_4200);
xor U5159 (N_5159,N_3877,N_4057);
nand U5160 (N_5160,N_3499,N_2233);
and U5161 (N_5161,N_1621,N_2860);
or U5162 (N_5162,N_544,N_3246);
nor U5163 (N_5163,N_3039,N_771);
xor U5164 (N_5164,N_3905,N_4596);
and U5165 (N_5165,N_927,N_4736);
nor U5166 (N_5166,N_1881,N_4675);
or U5167 (N_5167,N_1696,N_4892);
xnor U5168 (N_5168,N_3815,N_4756);
nor U5169 (N_5169,N_1279,N_4453);
nand U5170 (N_5170,N_4524,N_1491);
and U5171 (N_5171,N_92,N_584);
and U5172 (N_5172,N_736,N_1007);
nor U5173 (N_5173,N_2356,N_3349);
and U5174 (N_5174,N_4493,N_3700);
nor U5175 (N_5175,N_752,N_3221);
nand U5176 (N_5176,N_1814,N_2543);
and U5177 (N_5177,N_1397,N_2001);
and U5178 (N_5178,N_2938,N_3822);
xor U5179 (N_5179,N_374,N_4369);
and U5180 (N_5180,N_1127,N_2147);
nor U5181 (N_5181,N_4686,N_1226);
nand U5182 (N_5182,N_888,N_1474);
or U5183 (N_5183,N_653,N_3378);
and U5184 (N_5184,N_128,N_1772);
and U5185 (N_5185,N_4166,N_40);
xor U5186 (N_5186,N_3002,N_699);
or U5187 (N_5187,N_2144,N_2840);
nor U5188 (N_5188,N_3816,N_3609);
nand U5189 (N_5189,N_2673,N_1198);
nor U5190 (N_5190,N_2736,N_2338);
or U5191 (N_5191,N_3552,N_4253);
nand U5192 (N_5192,N_1487,N_1283);
xnor U5193 (N_5193,N_3296,N_3572);
nand U5194 (N_5194,N_1545,N_339);
nand U5195 (N_5195,N_4978,N_3563);
or U5196 (N_5196,N_4711,N_1897);
nand U5197 (N_5197,N_480,N_3687);
or U5198 (N_5198,N_3443,N_535);
nor U5199 (N_5199,N_4448,N_4249);
or U5200 (N_5200,N_330,N_4434);
nor U5201 (N_5201,N_389,N_4186);
nand U5202 (N_5202,N_3914,N_1138);
and U5203 (N_5203,N_473,N_153);
xor U5204 (N_5204,N_4391,N_217);
or U5205 (N_5205,N_4560,N_4248);
or U5206 (N_5206,N_4436,N_1603);
and U5207 (N_5207,N_2336,N_4);
nand U5208 (N_5208,N_1373,N_2028);
nand U5209 (N_5209,N_3202,N_4922);
nor U5210 (N_5210,N_3713,N_2590);
nand U5211 (N_5211,N_3277,N_4268);
nor U5212 (N_5212,N_2583,N_2024);
nand U5213 (N_5213,N_2060,N_3606);
nor U5214 (N_5214,N_4638,N_2359);
and U5215 (N_5215,N_4108,N_429);
nor U5216 (N_5216,N_1627,N_4457);
and U5217 (N_5217,N_1050,N_79);
and U5218 (N_5218,N_3315,N_721);
and U5219 (N_5219,N_461,N_392);
xnor U5220 (N_5220,N_3383,N_1149);
or U5221 (N_5221,N_4207,N_3017);
nor U5222 (N_5222,N_2278,N_4071);
nor U5223 (N_5223,N_769,N_2235);
xnor U5224 (N_5224,N_3775,N_4460);
nor U5225 (N_5225,N_1410,N_4232);
nor U5226 (N_5226,N_4441,N_2408);
nor U5227 (N_5227,N_1027,N_1516);
and U5228 (N_5228,N_3796,N_2689);
and U5229 (N_5229,N_774,N_1557);
nand U5230 (N_5230,N_1818,N_1428);
and U5231 (N_5231,N_4354,N_3071);
xnor U5232 (N_5232,N_658,N_4908);
nor U5233 (N_5233,N_3425,N_2858);
and U5234 (N_5234,N_848,N_3610);
nand U5235 (N_5235,N_4837,N_3080);
nor U5236 (N_5236,N_4969,N_4087);
nor U5237 (N_5237,N_4194,N_3727);
and U5238 (N_5238,N_277,N_939);
and U5239 (N_5239,N_1193,N_3138);
or U5240 (N_5240,N_3243,N_4321);
and U5241 (N_5241,N_524,N_4959);
and U5242 (N_5242,N_4043,N_3653);
nor U5243 (N_5243,N_2520,N_2093);
or U5244 (N_5244,N_117,N_4313);
nor U5245 (N_5245,N_3463,N_2255);
and U5246 (N_5246,N_817,N_1170);
and U5247 (N_5247,N_4886,N_657);
and U5248 (N_5248,N_4952,N_2960);
nor U5249 (N_5249,N_228,N_4423);
xnor U5250 (N_5250,N_1401,N_4094);
nor U5251 (N_5251,N_4707,N_4285);
nand U5252 (N_5252,N_3733,N_3382);
xnor U5253 (N_5253,N_1886,N_268);
nand U5254 (N_5254,N_2536,N_1471);
and U5255 (N_5255,N_3867,N_539);
and U5256 (N_5256,N_921,N_1575);
or U5257 (N_5257,N_137,N_4742);
nor U5258 (N_5258,N_2311,N_1372);
or U5259 (N_5259,N_1789,N_323);
xor U5260 (N_5260,N_3131,N_1921);
and U5261 (N_5261,N_4276,N_778);
nand U5262 (N_5262,N_4951,N_2984);
or U5263 (N_5263,N_3303,N_3532);
or U5264 (N_5264,N_2143,N_1606);
or U5265 (N_5265,N_1172,N_132);
xor U5266 (N_5266,N_2814,N_2782);
or U5267 (N_5267,N_3139,N_3069);
nand U5268 (N_5268,N_3611,N_4734);
or U5269 (N_5269,N_2269,N_4219);
xor U5270 (N_5270,N_149,N_3956);
or U5271 (N_5271,N_4407,N_2398);
nand U5272 (N_5272,N_4340,N_485);
nand U5273 (N_5273,N_1113,N_2181);
nor U5274 (N_5274,N_2394,N_1580);
or U5275 (N_5275,N_4466,N_2433);
and U5276 (N_5276,N_671,N_1667);
and U5277 (N_5277,N_820,N_4511);
nand U5278 (N_5278,N_2867,N_1820);
nor U5279 (N_5279,N_2690,N_3051);
nand U5280 (N_5280,N_836,N_3976);
or U5281 (N_5281,N_1834,N_2314);
or U5282 (N_5282,N_4023,N_2183);
or U5283 (N_5283,N_1629,N_1256);
nor U5284 (N_5284,N_4724,N_639);
nor U5285 (N_5285,N_3824,N_434);
nand U5286 (N_5286,N_550,N_2401);
or U5287 (N_5287,N_4789,N_23);
and U5288 (N_5288,N_3907,N_3591);
nor U5289 (N_5289,N_3838,N_222);
and U5290 (N_5290,N_4961,N_4463);
or U5291 (N_5291,N_3092,N_3327);
or U5292 (N_5292,N_1130,N_3000);
and U5293 (N_5293,N_1004,N_3117);
xor U5294 (N_5294,N_3476,N_42);
or U5295 (N_5295,N_50,N_1060);
nor U5296 (N_5296,N_2199,N_1494);
and U5297 (N_5297,N_525,N_3265);
and U5298 (N_5298,N_3095,N_4368);
nand U5299 (N_5299,N_4678,N_3283);
or U5300 (N_5300,N_1247,N_1720);
and U5301 (N_5301,N_2376,N_3748);
nand U5302 (N_5302,N_2646,N_1432);
nor U5303 (N_5303,N_207,N_551);
xnor U5304 (N_5304,N_1059,N_1176);
or U5305 (N_5305,N_1925,N_2617);
or U5306 (N_5306,N_3006,N_2479);
nor U5307 (N_5307,N_4074,N_3667);
and U5308 (N_5308,N_3862,N_3966);
nor U5309 (N_5309,N_775,N_869);
or U5310 (N_5310,N_1917,N_3214);
xor U5311 (N_5311,N_2633,N_4758);
nand U5312 (N_5312,N_2726,N_3830);
xnor U5313 (N_5313,N_4694,N_3478);
xor U5314 (N_5314,N_4717,N_2);
or U5315 (N_5315,N_1932,N_2080);
nand U5316 (N_5316,N_1609,N_2797);
nor U5317 (N_5317,N_432,N_468);
nor U5318 (N_5318,N_3114,N_2654);
or U5319 (N_5319,N_3016,N_590);
nor U5320 (N_5320,N_2008,N_2811);
or U5321 (N_5321,N_4095,N_1893);
nor U5322 (N_5322,N_2297,N_97);
nor U5323 (N_5323,N_4370,N_3105);
nand U5324 (N_5324,N_3473,N_2772);
and U5325 (N_5325,N_407,N_4716);
or U5326 (N_5326,N_2837,N_3176);
nand U5327 (N_5327,N_3579,N_1761);
or U5328 (N_5328,N_64,N_4665);
nand U5329 (N_5329,N_3964,N_4999);
and U5330 (N_5330,N_1534,N_2606);
nor U5331 (N_5331,N_4843,N_3629);
nor U5332 (N_5332,N_1620,N_276);
nand U5333 (N_5333,N_4159,N_3594);
nand U5334 (N_5334,N_4110,N_2003);
and U5335 (N_5335,N_4054,N_3033);
and U5336 (N_5336,N_3666,N_4894);
and U5337 (N_5337,N_1475,N_2485);
xor U5338 (N_5338,N_3538,N_3374);
nor U5339 (N_5339,N_4195,N_4595);
nand U5340 (N_5340,N_4791,N_3675);
and U5341 (N_5341,N_1776,N_1685);
or U5342 (N_5342,N_4714,N_1604);
or U5343 (N_5343,N_3268,N_2663);
and U5344 (N_5344,N_394,N_2388);
nor U5345 (N_5345,N_595,N_4269);
nor U5346 (N_5346,N_2910,N_1361);
and U5347 (N_5347,N_4705,N_4376);
nand U5348 (N_5348,N_2515,N_852);
or U5349 (N_5349,N_2943,N_1420);
nor U5350 (N_5350,N_4083,N_4084);
xor U5351 (N_5351,N_684,N_2699);
nor U5352 (N_5352,N_4220,N_4044);
and U5353 (N_5353,N_3674,N_4068);
nor U5354 (N_5354,N_129,N_4988);
or U5355 (N_5355,N_3369,N_1595);
nand U5356 (N_5356,N_1,N_3359);
nand U5357 (N_5357,N_1650,N_1773);
and U5358 (N_5358,N_3066,N_133);
nand U5359 (N_5359,N_4004,N_2608);
or U5360 (N_5360,N_4450,N_4612);
xor U5361 (N_5361,N_4051,N_1239);
nand U5362 (N_5362,N_2589,N_4279);
and U5363 (N_5363,N_3042,N_212);
nand U5364 (N_5364,N_1297,N_3123);
and U5365 (N_5365,N_3325,N_842);
nor U5366 (N_5366,N_1184,N_2538);
nor U5367 (N_5367,N_3337,N_2778);
nor U5368 (N_5368,N_3275,N_188);
or U5369 (N_5369,N_897,N_4191);
nand U5370 (N_5370,N_1848,N_2697);
xor U5371 (N_5371,N_169,N_3454);
nand U5372 (N_5372,N_4305,N_2599);
nand U5373 (N_5373,N_1267,N_2936);
xor U5374 (N_5374,N_4041,N_185);
nor U5375 (N_5375,N_248,N_2824);
or U5376 (N_5376,N_3641,N_4385);
nor U5377 (N_5377,N_994,N_1768);
nand U5378 (N_5378,N_4257,N_4876);
nor U5379 (N_5379,N_1223,N_3310);
nand U5380 (N_5380,N_3521,N_4374);
and U5381 (N_5381,N_2541,N_3133);
nor U5382 (N_5382,N_2585,N_635);
or U5383 (N_5383,N_3112,N_371);
nand U5384 (N_5384,N_2352,N_4920);
nand U5385 (N_5385,N_4852,N_1641);
nand U5386 (N_5386,N_2324,N_2117);
or U5387 (N_5387,N_2290,N_3288);
xor U5388 (N_5388,N_2613,N_1482);
or U5389 (N_5389,N_4216,N_3193);
nand U5390 (N_5390,N_2156,N_3686);
xnor U5391 (N_5391,N_2018,N_1398);
or U5392 (N_5392,N_834,N_2270);
xor U5393 (N_5393,N_3736,N_4251);
nand U5394 (N_5394,N_2516,N_1479);
or U5395 (N_5395,N_3682,N_2073);
xor U5396 (N_5396,N_3090,N_2211);
nor U5397 (N_5397,N_772,N_3423);
nand U5398 (N_5398,N_204,N_351);
or U5399 (N_5399,N_4066,N_2568);
and U5400 (N_5400,N_4266,N_3339);
or U5401 (N_5401,N_1757,N_4635);
nor U5402 (N_5402,N_119,N_3531);
and U5403 (N_5403,N_2229,N_166);
or U5404 (N_5404,N_3633,N_3854);
xnor U5405 (N_5405,N_4242,N_919);
or U5406 (N_5406,N_3172,N_2812);
or U5407 (N_5407,N_4745,N_3711);
nand U5408 (N_5408,N_4008,N_3021);
nor U5409 (N_5409,N_705,N_2645);
and U5410 (N_5410,N_4744,N_3965);
nor U5411 (N_5411,N_2505,N_652);
nor U5412 (N_5412,N_4685,N_4916);
and U5413 (N_5413,N_700,N_3460);
and U5414 (N_5414,N_4750,N_3657);
xnor U5415 (N_5415,N_3323,N_3141);
xor U5416 (N_5416,N_1750,N_2969);
or U5417 (N_5417,N_4367,N_3586);
xnor U5418 (N_5418,N_1635,N_1013);
and U5419 (N_5419,N_2801,N_4845);
and U5420 (N_5420,N_3044,N_961);
nor U5421 (N_5421,N_3635,N_90);
or U5422 (N_5422,N_2566,N_4033);
nor U5423 (N_5423,N_3735,N_3088);
or U5424 (N_5424,N_4082,N_594);
nor U5425 (N_5425,N_47,N_1493);
and U5426 (N_5426,N_2142,N_1237);
nor U5427 (N_5427,N_734,N_3714);
nand U5428 (N_5428,N_195,N_987);
nor U5429 (N_5429,N_2901,N_1864);
nand U5430 (N_5430,N_2500,N_4755);
and U5431 (N_5431,N_1514,N_1144);
or U5432 (N_5432,N_2406,N_3546);
nor U5433 (N_5433,N_4769,N_2638);
or U5434 (N_5434,N_1550,N_3177);
nor U5435 (N_5435,N_4848,N_3668);
nand U5436 (N_5436,N_823,N_4055);
nand U5437 (N_5437,N_200,N_1930);
nand U5438 (N_5438,N_3900,N_2898);
nand U5439 (N_5439,N_1519,N_2332);
or U5440 (N_5440,N_2214,N_2524);
nand U5441 (N_5441,N_4401,N_1896);
nor U5442 (N_5442,N_2842,N_2387);
xor U5443 (N_5443,N_4550,N_1501);
or U5444 (N_5444,N_62,N_1995);
and U5445 (N_5445,N_233,N_293);
or U5446 (N_5446,N_1586,N_1019);
and U5447 (N_5447,N_3134,N_1994);
nor U5448 (N_5448,N_1723,N_3401);
and U5449 (N_5449,N_3608,N_240);
nand U5450 (N_5450,N_2537,N_3504);
and U5451 (N_5451,N_3261,N_4264);
and U5452 (N_5452,N_542,N_811);
xnor U5453 (N_5453,N_1663,N_85);
xor U5454 (N_5454,N_164,N_4347);
or U5455 (N_5455,N_1800,N_1709);
nand U5456 (N_5456,N_3472,N_300);
and U5457 (N_5457,N_724,N_399);
nand U5458 (N_5458,N_4246,N_881);
nor U5459 (N_5459,N_4953,N_4732);
nand U5460 (N_5460,N_4483,N_1066);
or U5461 (N_5461,N_2866,N_420);
and U5462 (N_5462,N_4165,N_2383);
nor U5463 (N_5463,N_3052,N_2373);
and U5464 (N_5464,N_1584,N_2740);
xor U5465 (N_5465,N_1568,N_1110);
and U5466 (N_5466,N_124,N_1940);
and U5467 (N_5467,N_3651,N_421);
or U5468 (N_5468,N_3677,N_105);
or U5469 (N_5469,N_1429,N_4781);
and U5470 (N_5470,N_1012,N_2275);
or U5471 (N_5471,N_3364,N_2571);
or U5472 (N_5472,N_3162,N_4960);
xor U5473 (N_5473,N_325,N_1526);
and U5474 (N_5474,N_3974,N_4821);
nand U5475 (N_5475,N_4737,N_2271);
nand U5476 (N_5476,N_3897,N_2862);
or U5477 (N_5477,N_2221,N_1704);
xor U5478 (N_5478,N_3183,N_4019);
and U5479 (N_5479,N_4641,N_4040);
or U5480 (N_5480,N_2413,N_4782);
and U5481 (N_5481,N_4499,N_2733);
and U5482 (N_5482,N_851,N_2277);
xnor U5483 (N_5483,N_1210,N_1924);
xnor U5484 (N_5484,N_4995,N_569);
nor U5485 (N_5485,N_3111,N_1809);
nand U5486 (N_5486,N_444,N_879);
or U5487 (N_5487,N_4203,N_2742);
xor U5488 (N_5488,N_30,N_507);
and U5489 (N_5489,N_4490,N_314);
nand U5490 (N_5490,N_2468,N_3883);
xnor U5491 (N_5491,N_4206,N_688);
nor U5492 (N_5492,N_3395,N_19);
xor U5493 (N_5493,N_1762,N_1591);
or U5494 (N_5494,N_2055,N_732);
nand U5495 (N_5495,N_2574,N_2099);
or U5496 (N_5496,N_3448,N_712);
or U5497 (N_5497,N_3365,N_1644);
nor U5498 (N_5498,N_3818,N_666);
or U5499 (N_5499,N_4162,N_2040);
and U5500 (N_5500,N_859,N_4558);
or U5501 (N_5501,N_3913,N_15);
nor U5502 (N_5502,N_1084,N_2241);
and U5503 (N_5503,N_24,N_794);
nor U5504 (N_5504,N_4343,N_3545);
nand U5505 (N_5505,N_1845,N_4993);
or U5506 (N_5506,N_3293,N_4006);
and U5507 (N_5507,N_4757,N_342);
and U5508 (N_5508,N_2431,N_3240);
and U5509 (N_5509,N_3279,N_2013);
xor U5510 (N_5510,N_3520,N_3318);
nor U5511 (N_5511,N_130,N_2602);
nor U5512 (N_5512,N_2517,N_1408);
nand U5513 (N_5513,N_720,N_4743);
nor U5514 (N_5514,N_556,N_4238);
or U5515 (N_5515,N_4419,N_3084);
nand U5516 (N_5516,N_148,N_646);
xor U5517 (N_5517,N_2790,N_3120);
and U5518 (N_5518,N_1962,N_1551);
or U5519 (N_5519,N_2173,N_2035);
and U5520 (N_5520,N_1295,N_4459);
nor U5521 (N_5521,N_58,N_4888);
or U5522 (N_5522,N_2763,N_1274);
xnor U5523 (N_5523,N_1823,N_3839);
or U5524 (N_5524,N_2787,N_3348);
or U5525 (N_5525,N_4037,N_4890);
and U5526 (N_5526,N_4634,N_4334);
or U5527 (N_5527,N_3789,N_1950);
nand U5528 (N_5528,N_636,N_1148);
nand U5529 (N_5529,N_3160,N_932);
and U5530 (N_5530,N_1703,N_1978);
nor U5531 (N_5531,N_953,N_94);
or U5532 (N_5532,N_2743,N_4901);
nor U5533 (N_5533,N_4864,N_1232);
nor U5534 (N_5534,N_1031,N_144);
xor U5535 (N_5535,N_503,N_2360);
or U5536 (N_5536,N_612,N_4759);
and U5537 (N_5537,N_4433,N_4069);
xor U5538 (N_5538,N_309,N_2161);
and U5539 (N_5539,N_2307,N_1811);
or U5540 (N_5540,N_681,N_1868);
nor U5541 (N_5541,N_655,N_3922);
nand U5542 (N_5542,N_2601,N_4456);
and U5543 (N_5543,N_4224,N_4327);
or U5544 (N_5544,N_1590,N_740);
or U5545 (N_5545,N_3452,N_3484);
and U5546 (N_5546,N_4766,N_3074);
nand U5547 (N_5547,N_4820,N_1500);
or U5548 (N_5548,N_487,N_1119);
or U5549 (N_5549,N_2118,N_2883);
or U5550 (N_5550,N_4614,N_65);
nand U5551 (N_5551,N_4301,N_4898);
and U5552 (N_5552,N_1053,N_3205);
and U5553 (N_5553,N_4802,N_2048);
and U5554 (N_5554,N_2368,N_4721);
nor U5555 (N_5555,N_3731,N_770);
nand U5556 (N_5556,N_3846,N_1688);
or U5557 (N_5557,N_48,N_3187);
and U5558 (N_5558,N_1344,N_2534);
nand U5559 (N_5559,N_1261,N_2662);
nand U5560 (N_5560,N_1662,N_3871);
or U5561 (N_5561,N_650,N_4594);
xnor U5562 (N_5562,N_4606,N_812);
and U5563 (N_5563,N_4818,N_1040);
and U5564 (N_5564,N_2333,N_3281);
nand U5565 (N_5565,N_2921,N_3694);
and U5566 (N_5566,N_713,N_3576);
or U5567 (N_5567,N_1080,N_3420);
xor U5568 (N_5568,N_4261,N_2146);
nor U5569 (N_5569,N_3661,N_1484);
and U5570 (N_5570,N_2159,N_773);
or U5571 (N_5571,N_1513,N_1548);
and U5572 (N_5572,N_3618,N_896);
nor U5573 (N_5573,N_4406,N_98);
nor U5574 (N_5574,N_3587,N_435);
or U5575 (N_5575,N_516,N_1707);
and U5576 (N_5576,N_4860,N_789);
nor U5577 (N_5577,N_3998,N_1876);
nor U5578 (N_5578,N_2973,N_380);
or U5579 (N_5579,N_4786,N_4832);
xnor U5580 (N_5580,N_2464,N_235);
and U5581 (N_5581,N_1542,N_3232);
nand U5582 (N_5582,N_3723,N_522);
nor U5583 (N_5583,N_1499,N_1208);
or U5584 (N_5584,N_4565,N_515);
xor U5585 (N_5585,N_3953,N_2559);
nand U5586 (N_5586,N_962,N_2712);
or U5587 (N_5587,N_3076,N_3720);
nand U5588 (N_5588,N_2109,N_1633);
nor U5589 (N_5589,N_1065,N_4189);
xor U5590 (N_5590,N_1498,N_4016);
and U5591 (N_5591,N_1567,N_3695);
nand U5592 (N_5592,N_4767,N_4987);
or U5593 (N_5593,N_2337,N_4350);
and U5594 (N_5594,N_4795,N_4674);
nor U5595 (N_5595,N_4323,N_2926);
nor U5596 (N_5596,N_1777,N_2991);
nor U5597 (N_5597,N_1098,N_4497);
nor U5598 (N_5598,N_1298,N_3523);
or U5599 (N_5599,N_1675,N_1802);
xnor U5600 (N_5600,N_1072,N_1284);
nand U5601 (N_5601,N_1760,N_805);
and U5602 (N_5602,N_2793,N_1043);
or U5603 (N_5603,N_418,N_1640);
nor U5604 (N_5604,N_728,N_3980);
or U5605 (N_5605,N_3541,N_63);
and U5606 (N_5606,N_1353,N_1830);
nand U5607 (N_5607,N_3742,N_2411);
and U5608 (N_5608,N_3698,N_4143);
and U5609 (N_5609,N_4079,N_1810);
nor U5610 (N_5610,N_3559,N_785);
nand U5611 (N_5611,N_3453,N_1280);
nor U5612 (N_5612,N_2587,N_2249);
nor U5613 (N_5613,N_2966,N_1240);
nor U5614 (N_5614,N_4335,N_510);
nand U5615 (N_5615,N_4101,N_2577);
and U5616 (N_5616,N_2104,N_4982);
nand U5617 (N_5617,N_3892,N_68);
nand U5618 (N_5618,N_4866,N_192);
nor U5619 (N_5619,N_2031,N_2900);
or U5620 (N_5620,N_1960,N_4977);
or U5621 (N_5621,N_4496,N_1502);
nor U5622 (N_5622,N_2049,N_4576);
xnor U5623 (N_5623,N_1585,N_2887);
and U5624 (N_5624,N_803,N_1356);
xor U5625 (N_5625,N_1025,N_675);
or U5626 (N_5626,N_831,N_3367);
and U5627 (N_5627,N_1272,N_4529);
or U5628 (N_5628,N_1527,N_4539);
nand U5629 (N_5629,N_4628,N_3036);
and U5630 (N_5630,N_4868,N_2075);
nand U5631 (N_5631,N_737,N_999);
nor U5632 (N_5632,N_4780,N_6);
nand U5633 (N_5633,N_3253,N_3411);
or U5634 (N_5634,N_2875,N_2492);
nor U5635 (N_5635,N_1669,N_176);
xor U5636 (N_5636,N_4963,N_4749);
nor U5637 (N_5637,N_4476,N_2209);
and U5638 (N_5638,N_1661,N_2917);
xor U5639 (N_5639,N_4250,N_3008);
or U5640 (N_5640,N_3329,N_4454);
nor U5641 (N_5641,N_2392,N_1486);
and U5642 (N_5642,N_3732,N_186);
nor U5643 (N_5643,N_3010,N_317);
or U5644 (N_5644,N_1630,N_3430);
nor U5645 (N_5645,N_3362,N_32);
nand U5646 (N_5646,N_4400,N_3848);
and U5647 (N_5647,N_4164,N_146);
xor U5648 (N_5648,N_3498,N_1140);
and U5649 (N_5649,N_4934,N_66);
nand U5650 (N_5650,N_922,N_4217);
and U5651 (N_5651,N_1509,N_2054);
nor U5652 (N_5652,N_2282,N_3740);
and U5653 (N_5653,N_3996,N_1422);
and U5654 (N_5654,N_2546,N_707);
and U5655 (N_5655,N_4314,N_1216);
xnor U5656 (N_5656,N_1164,N_4531);
nand U5657 (N_5657,N_1922,N_914);
and U5658 (N_5658,N_1674,N_1351);
and U5659 (N_5659,N_1958,N_2243);
or U5660 (N_5660,N_1121,N_2928);
and U5661 (N_5661,N_3230,N_449);
and U5662 (N_5662,N_3124,N_2167);
or U5663 (N_5663,N_286,N_2386);
and U5664 (N_5664,N_4107,N_1861);
and U5665 (N_5665,N_2461,N_743);
and U5666 (N_5666,N_2487,N_3981);
nand U5667 (N_5667,N_289,N_1854);
and U5668 (N_5668,N_3539,N_3393);
nand U5669 (N_5669,N_1825,N_3975);
or U5670 (N_5670,N_2113,N_3774);
or U5671 (N_5671,N_1577,N_189);
nor U5672 (N_5672,N_3343,N_2947);
nand U5673 (N_5673,N_2427,N_627);
xor U5674 (N_5674,N_928,N_4031);
xor U5675 (N_5675,N_1331,N_3969);
xor U5676 (N_5676,N_1889,N_3185);
nand U5677 (N_5677,N_3869,N_2605);
nand U5678 (N_5678,N_108,N_321);
or U5679 (N_5679,N_2539,N_2007);
xnor U5680 (N_5680,N_3652,N_1323);
nand U5681 (N_5681,N_1461,N_2919);
nand U5682 (N_5682,N_1002,N_2807);
or U5683 (N_5683,N_926,N_3650);
nor U5684 (N_5684,N_2667,N_1158);
nand U5685 (N_5685,N_87,N_3402);
or U5686 (N_5686,N_886,N_2770);
and U5687 (N_5687,N_4443,N_1042);
nor U5688 (N_5688,N_1652,N_3483);
nand U5689 (N_5689,N_2705,N_2264);
and U5690 (N_5690,N_3338,N_3083);
nand U5691 (N_5691,N_122,N_271);
nor U5692 (N_5692,N_4779,N_618);
and U5693 (N_5693,N_753,N_1842);
nor U5694 (N_5694,N_183,N_1966);
or U5695 (N_5695,N_4687,N_4398);
nor U5696 (N_5696,N_1679,N_748);
or U5697 (N_5697,N_3450,N_1375);
or U5698 (N_5698,N_2416,N_2456);
and U5699 (N_5699,N_4056,N_4929);
nor U5700 (N_5700,N_4693,N_4410);
nand U5701 (N_5701,N_2625,N_438);
nand U5702 (N_5702,N_1419,N_2734);
or U5703 (N_5703,N_677,N_4399);
and U5704 (N_5704,N_425,N_1206);
or U5705 (N_5705,N_3837,N_4937);
xor U5706 (N_5706,N_988,N_2097);
and U5707 (N_5707,N_4383,N_1672);
nor U5708 (N_5708,N_1983,N_270);
nor U5709 (N_5709,N_1001,N_4684);
nor U5710 (N_5710,N_3688,N_2397);
or U5711 (N_5711,N_1390,N_4653);
or U5712 (N_5712,N_959,N_1217);
or U5713 (N_5713,N_2009,N_4256);
and U5714 (N_5714,N_2544,N_3173);
and U5715 (N_5715,N_4384,N_4332);
and U5716 (N_5716,N_4223,N_1798);
or U5717 (N_5717,N_1795,N_2828);
and U5718 (N_5718,N_4938,N_1979);
nand U5719 (N_5719,N_1637,N_315);
nand U5720 (N_5720,N_1282,N_3518);
nand U5721 (N_5721,N_1028,N_2977);
or U5722 (N_5722,N_4522,N_2119);
nand U5723 (N_5723,N_456,N_211);
nand U5724 (N_5724,N_1951,N_1187);
nor U5725 (N_5725,N_3057,N_3860);
or U5726 (N_5726,N_4117,N_4994);
and U5727 (N_5727,N_1178,N_1221);
nor U5728 (N_5728,N_615,N_302);
nand U5729 (N_5729,N_2562,N_4296);
or U5730 (N_5730,N_3492,N_1128);
xnor U5731 (N_5731,N_4028,N_4656);
and U5732 (N_5732,N_4386,N_2989);
and U5733 (N_5733,N_825,N_443);
or U5734 (N_5734,N_2478,N_3690);
or U5735 (N_5735,N_1944,N_3751);
xnor U5736 (N_5736,N_4715,N_1156);
nor U5737 (N_5737,N_964,N_3407);
nor U5738 (N_5738,N_3923,N_764);
nand U5739 (N_5739,N_1008,N_3597);
and U5740 (N_5740,N_3491,N_3428);
nor U5741 (N_5741,N_1537,N_2959);
nand U5742 (N_5742,N_2871,N_406);
and U5743 (N_5743,N_2789,N_1518);
nand U5744 (N_5744,N_3258,N_1191);
nand U5745 (N_5745,N_2886,N_1753);
nor U5746 (N_5746,N_2390,N_1003);
nor U5747 (N_5747,N_3019,N_4676);
or U5748 (N_5748,N_1909,N_1413);
xnor U5749 (N_5749,N_1598,N_3188);
nand U5750 (N_5750,N_1213,N_4664);
nand U5751 (N_5751,N_4255,N_1708);
and U5752 (N_5752,N_1507,N_4785);
nor U5753 (N_5753,N_1624,N_2177);
nand U5754 (N_5754,N_364,N_27);
and U5755 (N_5755,N_3566,N_1808);
and U5756 (N_5756,N_1976,N_1289);
nor U5757 (N_5757,N_2245,N_2958);
and U5758 (N_5758,N_78,N_4907);
and U5759 (N_5759,N_2780,N_905);
nor U5760 (N_5760,N_243,N_617);
nand U5761 (N_5761,N_2551,N_2683);
or U5762 (N_5762,N_1199,N_1895);
nor U5763 (N_5763,N_3644,N_241);
and U5764 (N_5764,N_2765,N_2967);
nor U5765 (N_5765,N_1578,N_4026);
and U5766 (N_5766,N_735,N_411);
nand U5767 (N_5767,N_891,N_4078);
and U5768 (N_5768,N_4102,N_1087);
nand U5769 (N_5769,N_1522,N_3841);
nor U5770 (N_5770,N_2238,N_3274);
or U5771 (N_5771,N_345,N_4730);
nor U5772 (N_5772,N_1270,N_1715);
or U5773 (N_5773,N_944,N_4566);
nand U5774 (N_5774,N_597,N_1926);
or U5775 (N_5775,N_793,N_4326);
or U5776 (N_5776,N_193,N_1081);
and U5777 (N_5777,N_4131,N_585);
xor U5778 (N_5778,N_306,N_4763);
and U5779 (N_5779,N_455,N_916);
nor U5780 (N_5780,N_2116,N_1388);
or U5781 (N_5781,N_3102,N_4494);
nand U5782 (N_5782,N_4998,N_3344);
and U5783 (N_5783,N_913,N_313);
and U5784 (N_5784,N_2890,N_2162);
or U5785 (N_5785,N_1576,N_4226);
nand U5786 (N_5786,N_1180,N_1301);
and U5787 (N_5787,N_2729,N_1054);
or U5788 (N_5788,N_3631,N_3890);
or U5789 (N_5789,N_3678,N_4752);
or U5790 (N_5790,N_2825,N_3783);
nor U5791 (N_5791,N_4122,N_4169);
xnor U5792 (N_5792,N_2894,N_2678);
xor U5793 (N_5793,N_3286,N_2042);
nand U5794 (N_5794,N_4475,N_3477);
nor U5795 (N_5795,N_4284,N_4010);
nor U5796 (N_5796,N_1105,N_3182);
or U5797 (N_5797,N_2682,N_4294);
xor U5798 (N_5798,N_1936,N_2294);
nand U5799 (N_5799,N_2757,N_1833);
or U5800 (N_5800,N_4912,N_4699);
nand U5801 (N_5801,N_2467,N_4175);
and U5802 (N_5802,N_4298,N_1472);
and U5803 (N_5803,N_739,N_3406);
nor U5804 (N_5804,N_1968,N_2841);
and U5805 (N_5805,N_3779,N_4600);
and U5806 (N_5806,N_4014,N_2512);
and U5807 (N_5807,N_1855,N_3790);
and U5808 (N_5808,N_1073,N_4991);
and U5809 (N_5809,N_2985,N_4955);
nand U5810 (N_5810,N_4104,N_1389);
nand U5811 (N_5811,N_583,N_2598);
xor U5812 (N_5812,N_2727,N_159);
or U5813 (N_5813,N_1564,N_224);
nor U5814 (N_5814,N_1296,N_2558);
and U5815 (N_5815,N_155,N_2384);
nor U5816 (N_5816,N_954,N_156);
nand U5817 (N_5817,N_4746,N_2378);
and U5818 (N_5818,N_4646,N_3561);
and U5819 (N_5819,N_2854,N_8);
and U5820 (N_5820,N_1411,N_4879);
xor U5821 (N_5821,N_941,N_3213);
or U5822 (N_5822,N_3,N_555);
nor U5823 (N_5823,N_529,N_2239);
nor U5824 (N_5824,N_3299,N_1816);
and U5825 (N_5825,N_1931,N_2805);
or U5826 (N_5826,N_4501,N_587);
nor U5827 (N_5827,N_335,N_2429);
and U5828 (N_5828,N_1227,N_3379);
xnor U5829 (N_5829,N_2721,N_4804);
nand U5830 (N_5830,N_1565,N_756);
nor U5831 (N_5831,N_2369,N_279);
xnor U5832 (N_5832,N_386,N_4417);
or U5833 (N_5833,N_1362,N_3785);
or U5834 (N_5834,N_13,N_4733);
nor U5835 (N_5835,N_1139,N_3991);
or U5836 (N_5836,N_3178,N_1214);
or U5837 (N_5837,N_2785,N_482);
nor U5838 (N_5838,N_2694,N_2298);
nor U5839 (N_5839,N_1741,N_1536);
nor U5840 (N_5840,N_1248,N_1579);
and U5841 (N_5841,N_3100,N_2724);
and U5842 (N_5842,N_1263,N_3306);
nand U5843 (N_5843,N_254,N_465);
xnor U5844 (N_5844,N_3543,N_611);
nand U5845 (N_5845,N_2584,N_3280);
nor U5846 (N_5846,N_489,N_172);
nand U5847 (N_5847,N_2346,N_4765);
xnor U5848 (N_5848,N_2322,N_3879);
or U5849 (N_5849,N_3868,N_1327);
xor U5850 (N_5850,N_1183,N_716);
xor U5851 (N_5851,N_575,N_3726);
or U5852 (N_5852,N_3319,N_2857);
nor U5853 (N_5853,N_4225,N_2375);
nand U5854 (N_5854,N_4647,N_4887);
nor U5855 (N_5855,N_263,N_2644);
or U5856 (N_5856,N_2941,N_4857);
xnor U5857 (N_5857,N_982,N_2831);
nor U5858 (N_5858,N_3259,N_3053);
or U5859 (N_5859,N_135,N_4679);
xor U5860 (N_5860,N_990,N_1791);
and U5861 (N_5861,N_4103,N_4346);
nand U5862 (N_5862,N_1812,N_326);
nand U5863 (N_5863,N_3408,N_1980);
nor U5864 (N_5864,N_3903,N_554);
or U5865 (N_5865,N_219,N_861);
or U5866 (N_5866,N_2205,N_1838);
xnor U5867 (N_5867,N_1424,N_1168);
or U5868 (N_5868,N_2185,N_1278);
and U5869 (N_5869,N_4451,N_4352);
nand U5870 (N_5870,N_1262,N_4727);
or U5871 (N_5871,N_4918,N_1076);
nor U5872 (N_5872,N_2335,N_3569);
nand U5873 (N_5873,N_3206,N_4292);
nor U5874 (N_5874,N_3255,N_4624);
nor U5875 (N_5875,N_459,N_4621);
nor U5876 (N_5876,N_1449,N_2676);
nor U5877 (N_5877,N_1505,N_2169);
or U5878 (N_5878,N_4883,N_3381);
xnor U5879 (N_5879,N_4893,N_4632);
nor U5880 (N_5880,N_4545,N_1333);
nand U5881 (N_5881,N_2123,N_2557);
and U5882 (N_5882,N_4981,N_1748);
and U5883 (N_5883,N_3445,N_669);
and U5884 (N_5884,N_904,N_2869);
nor U5885 (N_5885,N_3266,N_3242);
nor U5886 (N_5886,N_2471,N_3375);
nor U5887 (N_5887,N_3026,N_1541);
nand U5888 (N_5888,N_1544,N_2622);
nor U5889 (N_5889,N_1392,N_2777);
nand U5890 (N_5890,N_659,N_2833);
nor U5891 (N_5891,N_3864,N_4826);
or U5892 (N_5892,N_3438,N_301);
or U5893 (N_5893,N_1338,N_521);
and U5894 (N_5894,N_4620,N_1159);
xor U5895 (N_5895,N_4642,N_801);
nand U5896 (N_5896,N_2665,N_2918);
nor U5897 (N_5897,N_3896,N_1211);
or U5898 (N_5898,N_1655,N_2674);
or U5899 (N_5899,N_1758,N_4623);
or U5900 (N_5900,N_1197,N_179);
nand U5901 (N_5901,N_4905,N_493);
or U5902 (N_5902,N_3142,N_4442);
or U5903 (N_5903,N_3647,N_901);
nor U5904 (N_5904,N_3159,N_2469);
and U5905 (N_5905,N_540,N_178);
and U5906 (N_5906,N_4793,N_1885);
nor U5907 (N_5907,N_4357,N_4921);
xnor U5908 (N_5908,N_3118,N_3654);
or U5909 (N_5909,N_4610,N_3548);
nand U5910 (N_5910,N_1786,N_2422);
nand U5911 (N_5911,N_1919,N_1657);
nor U5912 (N_5912,N_2194,N_3065);
and U5913 (N_5913,N_798,N_3449);
xnor U5914 (N_5914,N_4609,N_1167);
and U5915 (N_5915,N_4091,N_3764);
nand U5916 (N_5916,N_1954,N_347);
nand U5917 (N_5917,N_3169,N_622);
and U5918 (N_5918,N_2435,N_3391);
or U5919 (N_5919,N_1450,N_4156);
nor U5920 (N_5920,N_154,N_2507);
nor U5921 (N_5921,N_1063,N_557);
or U5922 (N_5922,N_2127,N_1244);
or U5923 (N_5923,N_3289,N_2481);
or U5924 (N_5924,N_2139,N_3979);
and U5925 (N_5925,N_214,N_393);
nand U5926 (N_5926,N_4467,N_2006);
or U5927 (N_5927,N_336,N_2641);
nor U5928 (N_5928,N_4927,N_1787);
or U5929 (N_5929,N_673,N_2513);
nand U5930 (N_5930,N_1612,N_4824);
or U5931 (N_5931,N_4518,N_4064);
xnor U5932 (N_5932,N_1682,N_4914);
and U5933 (N_5933,N_4437,N_2045);
and U5934 (N_5934,N_4009,N_4613);
or U5935 (N_5935,N_3517,N_4022);
nand U5936 (N_5936,N_2784,N_2767);
xnor U5937 (N_5937,N_4773,N_780);
or U5938 (N_5938,N_1052,N_4137);
nand U5939 (N_5939,N_1319,N_822);
xnor U5940 (N_5940,N_4895,N_965);
nor U5941 (N_5941,N_3904,N_2460);
nand U5942 (N_5942,N_3292,N_1602);
nand U5943 (N_5943,N_1091,N_3475);
nand U5944 (N_5944,N_54,N_2761);
nand U5945 (N_5945,N_4058,N_2069);
nor U5946 (N_5946,N_3595,N_3994);
nand U5947 (N_5947,N_4422,N_4380);
xnor U5948 (N_5948,N_4362,N_3482);
nand U5949 (N_5949,N_727,N_1143);
nand U5950 (N_5950,N_1142,N_1803);
and U5951 (N_5951,N_2323,N_3486);
nand U5952 (N_5952,N_3440,N_1901);
or U5953 (N_5953,N_462,N_2428);
xnor U5954 (N_5954,N_708,N_4306);
or U5955 (N_5955,N_1725,N_685);
and U5956 (N_5956,N_4651,N_1955);
nor U5957 (N_5957,N_4182,N_2201);
or U5958 (N_5958,N_352,N_4517);
nor U5959 (N_5959,N_1102,N_1572);
nand U5960 (N_5960,N_4090,N_2339);
nand U5961 (N_5961,N_4992,N_2061);
and U5962 (N_5962,N_198,N_4065);
or U5963 (N_5963,N_3685,N_1884);
and U5964 (N_5964,N_4541,N_363);
nand U5965 (N_5965,N_4097,N_4295);
or U5966 (N_5966,N_1347,N_1618);
nand U5967 (N_5967,N_1862,N_3305);
nor U5968 (N_5968,N_1532,N_1116);
or U5969 (N_5969,N_4316,N_3585);
or U5970 (N_5970,N_3888,N_2951);
nor U5971 (N_5971,N_1229,N_768);
or U5972 (N_5972,N_453,N_1869);
or U5973 (N_5973,N_3805,N_719);
nor U5974 (N_5974,N_4093,N_1056);
or U5975 (N_5975,N_4871,N_91);
nand U5976 (N_5976,N_3161,N_3497);
xor U5977 (N_5977,N_1872,N_4954);
and U5978 (N_5978,N_1382,N_1804);
and U5979 (N_5979,N_985,N_2775);
nor U5980 (N_5980,N_2094,N_110);
nor U5981 (N_5981,N_1443,N_4829);
nor U5982 (N_5982,N_4355,N_4880);
or U5983 (N_5983,N_4320,N_2027);
nand U5984 (N_5984,N_4472,N_4972);
nor U5985 (N_5985,N_3075,N_626);
and U5986 (N_5986,N_4318,N_2070);
and U5987 (N_5987,N_4412,N_692);
and U5988 (N_5988,N_4590,N_3898);
nand U5989 (N_5989,N_2643,N_4050);
nor U5990 (N_5990,N_275,N_4611);
nand U5991 (N_5991,N_1610,N_4599);
or U5992 (N_5992,N_1483,N_4125);
xor U5993 (N_5993,N_4670,N_236);
nand U5994 (N_5994,N_1778,N_3920);
nor U5995 (N_5995,N_4447,N_796);
or U5996 (N_5996,N_3054,N_2879);
or U5997 (N_5997,N_3547,N_3334);
or U5998 (N_5998,N_3777,N_2304);
and U5999 (N_5999,N_3422,N_4411);
nor U6000 (N_6000,N_2066,N_3063);
nand U6001 (N_6001,N_2994,N_2810);
or U6002 (N_6002,N_4462,N_3495);
xnor U6003 (N_6003,N_2796,N_4525);
or U6004 (N_6004,N_205,N_490);
nor U6005 (N_6005,N_83,N_1417);
nand U6006 (N_6006,N_2446,N_4650);
nor U6007 (N_6007,N_2962,N_3909);
or U6008 (N_6008,N_951,N_171);
nand U6009 (N_6009,N_1846,N_2680);
or U6010 (N_6010,N_3939,N_460);
xnor U6011 (N_6011,N_830,N_3209);
nor U6012 (N_6012,N_643,N_3077);
and U6013 (N_6013,N_3760,N_2219);
or U6014 (N_6014,N_1705,N_1533);
and U6015 (N_6015,N_649,N_4263);
or U6016 (N_6016,N_2095,N_1972);
xor U6017 (N_6017,N_1678,N_2892);
nand U6018 (N_6018,N_2648,N_672);
or U6019 (N_6019,N_782,N_4508);
xor U6020 (N_6020,N_1996,N_948);
nor U6021 (N_6021,N_1111,N_2612);
nor U6022 (N_6022,N_3409,N_1736);
xnor U6023 (N_6023,N_2744,N_2038);
and U6024 (N_6024,N_3925,N_2437);
nor U6025 (N_6025,N_362,N_2501);
and U6026 (N_6026,N_4176,N_4221);
nand U6027 (N_6027,N_4547,N_4427);
nor U6028 (N_6028,N_3786,N_4036);
and U6029 (N_6029,N_4197,N_2573);
nor U6030 (N_6030,N_3208,N_4244);
and U6031 (N_6031,N_2058,N_1254);
or U6032 (N_6032,N_942,N_2135);
nor U6033 (N_6033,N_409,N_3983);
nor U6034 (N_6034,N_4777,N_4741);
and U6035 (N_6035,N_4958,N_3776);
or U6036 (N_6036,N_2870,N_1415);
or U6037 (N_6037,N_3345,N_346);
and U6038 (N_6038,N_3540,N_4163);
or U6039 (N_6039,N_1326,N_4899);
nand U6040 (N_6040,N_3982,N_3302);
or U6041 (N_6041,N_1850,N_1459);
nand U6042 (N_6042,N_779,N_1546);
nand U6043 (N_6043,N_4926,N_1134);
nand U6044 (N_6044,N_1859,N_4096);
xor U6045 (N_6045,N_3676,N_1749);
nand U6046 (N_6046,N_4669,N_1360);
and U6047 (N_6047,N_1045,N_3224);
xnor U6048 (N_6048,N_4484,N_4689);
or U6049 (N_6049,N_4415,N_2813);
or U6050 (N_6050,N_4358,N_2603);
or U6051 (N_6051,N_1370,N_3236);
nor U6052 (N_6052,N_4196,N_2473);
nand U6053 (N_6053,N_1874,N_2286);
and U6054 (N_6054,N_4080,N_376);
nand U6055 (N_6055,N_3536,N_3353);
or U6056 (N_6056,N_4910,N_4739);
and U6057 (N_6057,N_2272,N_1497);
xnor U6058 (N_6058,N_3271,N_2698);
and U6059 (N_6059,N_3360,N_2341);
or U6060 (N_6060,N_1694,N_368);
nand U6061 (N_6061,N_895,N_3328);
xor U6062 (N_6062,N_4809,N_3252);
nor U6063 (N_6063,N_2640,N_4485);
or U6064 (N_6064,N_21,N_1699);
and U6065 (N_6065,N_4477,N_4713);
or U6066 (N_6066,N_1614,N_127);
or U6067 (N_6067,N_2263,N_3503);
nor U6068 (N_6068,N_3604,N_2575);
xnor U6069 (N_6069,N_3554,N_3763);
or U6070 (N_6070,N_2056,N_4940);
or U6071 (N_6071,N_2762,N_261);
nor U6072 (N_6072,N_582,N_4601);
or U6073 (N_6073,N_3801,N_4153);
nor U6074 (N_6074,N_3502,N_3219);
nor U6075 (N_6075,N_4770,N_2382);
and U6076 (N_6076,N_9,N_2441);
xnor U6077 (N_6077,N_2102,N_1835);
or U6078 (N_6078,N_1122,N_4764);
xor U6079 (N_6079,N_931,N_1911);
and U6080 (N_6080,N_1448,N_3684);
nor U6081 (N_6081,N_3106,N_4389);
xor U6082 (N_6082,N_963,N_1673);
nor U6083 (N_6083,N_2020,N_3709);
nor U6084 (N_6084,N_2691,N_4478);
nand U6085 (N_6085,N_3908,N_1330);
xnor U6086 (N_6086,N_2044,N_4487);
or U6087 (N_6087,N_591,N_331);
nand U6088 (N_6088,N_1147,N_1405);
nor U6089 (N_6089,N_2050,N_1676);
nand U6090 (N_6090,N_2017,N_3707);
nor U6091 (N_6091,N_3312,N_4976);
and U6092 (N_6092,N_1228,N_218);
and U6093 (N_6093,N_1300,N_1255);
and U6094 (N_6094,N_383,N_3512);
or U6095 (N_6095,N_4862,N_4471);
and U6096 (N_6096,N_4924,N_3863);
nor U6097 (N_6097,N_559,N_2291);
nand U6098 (N_6098,N_1014,N_2074);
xnor U6099 (N_6099,N_4309,N_3078);
nor U6100 (N_6100,N_1622,N_856);
and U6101 (N_6101,N_2827,N_766);
nand U6102 (N_6102,N_2108,N_3496);
and U6103 (N_6103,N_3916,N_872);
and U6104 (N_6104,N_2130,N_4947);
nand U6105 (N_6105,N_2906,N_1252);
or U6106 (N_6106,N_989,N_2223);
nand U6107 (N_6107,N_1840,N_2896);
nand U6108 (N_6108,N_1123,N_3331);
nor U6109 (N_6109,N_260,N_1477);
xnor U6110 (N_6110,N_287,N_1355);
nor U6111 (N_6111,N_1731,N_4402);
xor U6112 (N_6112,N_1540,N_857);
and U6113 (N_6113,N_661,N_4470);
and U6114 (N_6114,N_3899,N_4896);
or U6115 (N_6115,N_2057,N_3469);
nor U6116 (N_6116,N_4731,N_1596);
and U6117 (N_6117,N_2912,N_2280);
nor U6118 (N_6118,N_2328,N_548);
and U6119 (N_6119,N_610,N_1189);
nor U6120 (N_6120,N_2350,N_142);
and U6121 (N_6121,N_3056,N_4722);
nor U6122 (N_6122,N_741,N_747);
nor U6123 (N_6123,N_763,N_2032);
nand U6124 (N_6124,N_1754,N_1233);
or U6125 (N_6125,N_2025,N_704);
nand U6126 (N_6126,N_3035,N_3455);
or U6127 (N_6127,N_536,N_4260);
xor U6128 (N_6128,N_123,N_2372);
and U6129 (N_6129,N_2675,N_3704);
or U6130 (N_6130,N_945,N_3534);
and U6131 (N_6131,N_161,N_3144);
nand U6132 (N_6132,N_2686,N_923);
xnor U6133 (N_6133,N_3553,N_4160);
or U6134 (N_6134,N_1313,N_3372);
and U6135 (N_6135,N_1431,N_255);
nand U6136 (N_6136,N_39,N_2934);
and U6137 (N_6137,N_2609,N_1525);
and U6138 (N_6138,N_2445,N_696);
nor U6139 (N_6139,N_3060,N_2244);
nand U6140 (N_6140,N_2340,N_3392);
or U6141 (N_6141,N_3340,N_4204);
nand U6142 (N_6142,N_2217,N_1064);
or U6143 (N_6143,N_1717,N_2114);
or U6144 (N_6144,N_4138,N_2450);
nor U6145 (N_6145,N_2347,N_3013);
nor U6146 (N_6146,N_3832,N_2193);
nor U6147 (N_6147,N_295,N_2548);
and U6148 (N_6148,N_1320,N_3316);
or U6149 (N_6149,N_4807,N_2749);
xnor U6150 (N_6150,N_3415,N_2508);
and U6151 (N_6151,N_3692,N_2086);
and U6152 (N_6152,N_1350,N_874);
and U6153 (N_6153,N_3673,N_4128);
nand U6154 (N_6154,N_608,N_3954);
or U6155 (N_6155,N_1416,N_4425);
nand U6156 (N_6156,N_4671,N_2836);
nor U6157 (N_6157,N_2308,N_5);
nor U6158 (N_6158,N_3865,N_1430);
and U6159 (N_6159,N_3333,N_496);
and U6160 (N_6160,N_3845,N_1999);
or U6161 (N_6161,N_3082,N_660);
or U6162 (N_6162,N_4816,N_2616);
and U6163 (N_6163,N_3434,N_397);
nor U6164 (N_6164,N_3137,N_4673);
nor U6165 (N_6165,N_4870,N_4970);
or U6166 (N_6166,N_4666,N_3895);
and U6167 (N_6167,N_1560,N_1281);
nand U6168 (N_6168,N_3873,N_527);
and U6169 (N_6169,N_3741,N_2284);
xnor U6170 (N_6170,N_2972,N_2227);
nor U6171 (N_6171,N_1086,N_3840);
nand U6172 (N_6172,N_1462,N_4812);
or U6173 (N_6173,N_1460,N_2092);
nor U6174 (N_6174,N_3151,N_4702);
nand U6175 (N_6175,N_2476,N_2715);
xor U6176 (N_6176,N_2493,N_3041);
nor U6177 (N_6177,N_1539,N_273);
nor U6178 (N_6178,N_625,N_4480);
nor U6179 (N_6179,N_4046,N_3429);
or U6180 (N_6180,N_3808,N_139);
nand U6181 (N_6181,N_1403,N_1934);
nor U6182 (N_6182,N_2816,N_1058);
nor U6183 (N_6183,N_257,N_3693);
or U6184 (N_6184,N_76,N_1264);
nor U6185 (N_6185,N_414,N_357);
nand U6186 (N_6186,N_3218,N_2996);
nand U6187 (N_6187,N_457,N_4170);
nor U6188 (N_6188,N_4806,N_1783);
and U6189 (N_6189,N_4873,N_3921);
or U6190 (N_6190,N_3179,N_4615);
and U6191 (N_6191,N_3417,N_4388);
and U6192 (N_6192,N_3788,N_34);
or U6193 (N_6193,N_1691,N_3821);
or U6194 (N_6194,N_3196,N_4648);
and U6195 (N_6195,N_1656,N_1075);
nand U6196 (N_6196,N_2774,N_1852);
nand U6197 (N_6197,N_4808,N_1763);
xnor U6198 (N_6198,N_973,N_2292);
or U6199 (N_6199,N_952,N_2421);
nand U6200 (N_6200,N_1503,N_2358);
or U6201 (N_6201,N_3191,N_3522);
or U6202 (N_6202,N_1468,N_4593);
and U6203 (N_6203,N_4690,N_483);
nor U6204 (N_6204,N_410,N_2792);
nand U6205 (N_6205,N_979,N_3474);
nand U6206 (N_6206,N_3881,N_341);
and U6207 (N_6207,N_2226,N_4077);
nand U6208 (N_6208,N_3070,N_3519);
and U6209 (N_6209,N_2746,N_2256);
nor U6210 (N_6210,N_2374,N_2904);
nor U6211 (N_6211,N_3513,N_2527);
nand U6212 (N_6212,N_2660,N_354);
nor U6213 (N_6213,N_1806,N_4578);
nor U6214 (N_6214,N_4073,N_3291);
nor U6215 (N_6215,N_4867,N_2529);
and U6216 (N_6216,N_1292,N_2158);
nand U6217 (N_6217,N_4630,N_3061);
nand U6218 (N_6218,N_1157,N_1162);
xor U6219 (N_6219,N_3910,N_2076);
nand U6220 (N_6220,N_4863,N_799);
and U6221 (N_6221,N_868,N_829);
xnor U6222 (N_6222,N_2719,N_3262);
nand U6223 (N_6223,N_632,N_3043);
nor U6224 (N_6224,N_3186,N_786);
nor U6225 (N_6225,N_2488,N_2895);
nor U6226 (N_6226,N_1445,N_388);
nand U6227 (N_6227,N_2563,N_181);
nor U6228 (N_6228,N_4652,N_2396);
nor U6229 (N_6229,N_4202,N_145);
nand U6230 (N_6230,N_1945,N_2029);
or U6231 (N_6231,N_1101,N_375);
nor U6232 (N_6232,N_1841,N_1726);
xor U6233 (N_6233,N_7,N_508);
xor U6234 (N_6234,N_338,N_502);
nand U6235 (N_6235,N_4420,N_821);
or U6236 (N_6236,N_745,N_2661);
nand U6237 (N_6237,N_4063,N_4192);
xor U6238 (N_6238,N_4842,N_2863);
and U6239 (N_6239,N_2412,N_1769);
or U6240 (N_6240,N_2899,N_571);
nor U6241 (N_6241,N_3079,N_4439);
nor U6242 (N_6242,N_4579,N_3758);
and U6243 (N_6243,N_4608,N_2062);
or U6244 (N_6244,N_2864,N_600);
nand U6245 (N_6245,N_606,N_1182);
nand U6246 (N_6246,N_337,N_2165);
nor U6247 (N_6247,N_3180,N_2195);
nor U6248 (N_6248,N_1088,N_4047);
nor U6249 (N_6249,N_3110,N_2615);
xor U6250 (N_6250,N_3843,N_787);
and U6251 (N_6251,N_4825,N_2310);
nor U6252 (N_6252,N_3347,N_3894);
nor U6253 (N_6253,N_252,N_2876);
or U6254 (N_6254,N_2914,N_2514);
xor U6255 (N_6255,N_3926,N_494);
xor U6256 (N_6256,N_738,N_1780);
xnor U6257 (N_6257,N_1908,N_1929);
nand U6258 (N_6258,N_1660,N_2182);
nor U6259 (N_6259,N_3031,N_3828);
nand U6260 (N_6260,N_3530,N_3931);
nand U6261 (N_6261,N_3147,N_100);
and U6262 (N_6262,N_272,N_274);
nand U6263 (N_6263,N_4854,N_3426);
nor U6264 (N_6264,N_2927,N_203);
and U6265 (N_6265,N_4772,N_486);
nand U6266 (N_6266,N_2861,N_2672);
nand U6267 (N_6267,N_2593,N_1132);
nand U6268 (N_6268,N_408,N_1414);
and U6269 (N_6269,N_2036,N_1774);
or U6270 (N_6270,N_4288,N_549);
nand U6271 (N_6271,N_2216,N_1466);
or U6272 (N_6272,N_2215,N_1435);
or U6273 (N_6273,N_4339,N_2240);
and U6274 (N_6274,N_3109,N_3220);
xnor U6275 (N_6275,N_14,N_3592);
or U6276 (N_6276,N_4302,N_2872);
and U6277 (N_6277,N_2480,N_3320);
or U6278 (N_6278,N_1837,N_2693);
nor U6279 (N_6279,N_2316,N_3250);
nand U6280 (N_6280,N_2279,N_2141);
or U6281 (N_6281,N_1153,N_3619);
nor U6282 (N_6282,N_3326,N_1192);
nand U6283 (N_6283,N_4555,N_2963);
nand U6284 (N_6284,N_3973,N_4917);
nor U6285 (N_6285,N_4218,N_3639);
nor U6286 (N_6286,N_900,N_1902);
xor U6287 (N_6287,N_2377,N_2417);
xor U6288 (N_6288,N_2823,N_1528);
and U6289 (N_6289,N_3578,N_1562);
nand U6290 (N_6290,N_2206,N_4173);
xor U6291 (N_6291,N_1587,N_1093);
and U6292 (N_6292,N_3386,N_433);
nor U6293 (N_6293,N_3582,N_3468);
nor U6294 (N_6294,N_2320,N_4663);
nor U6295 (N_6295,N_458,N_1225);
or U6296 (N_6296,N_423,N_3171);
nand U6297 (N_6297,N_4086,N_2576);
nor U6298 (N_6298,N_1457,N_593);
and U6299 (N_6299,N_3985,N_3632);
and U6300 (N_6300,N_3680,N_3164);
nor U6301 (N_6301,N_165,N_2126);
and U6302 (N_6302,N_2522,N_802);
nand U6303 (N_6303,N_1444,N_246);
nor U6304 (N_6304,N_4017,N_1547);
nor U6305 (N_6305,N_1421,N_2197);
or U6306 (N_6306,N_2893,N_693);
nor U6307 (N_6307,N_4145,N_1670);
and U6308 (N_6308,N_2504,N_2530);
and U6309 (N_6309,N_3853,N_1030);
and U6310 (N_6310,N_2652,N_2634);
nand U6311 (N_6311,N_2874,N_3803);
and U6312 (N_6312,N_416,N_2078);
and U6313 (N_6313,N_4061,N_903);
nor U6314 (N_6314,N_2771,N_3663);
and U6315 (N_6315,N_220,N_776);
and U6316 (N_6316,N_10,N_3986);
and U6317 (N_6317,N_809,N_3081);
nor U6318 (N_6318,N_2220,N_572);
or U6319 (N_6319,N_3978,N_2451);
nor U6320 (N_6320,N_2287,N_1092);
xnor U6321 (N_6321,N_3542,N_3104);
or U6322 (N_6322,N_3665,N_3809);
nand U6323 (N_6323,N_450,N_2367);
and U6324 (N_6324,N_4049,N_1317);
or U6325 (N_6325,N_3424,N_1386);
nor U6326 (N_6326,N_1458,N_4179);
and U6327 (N_6327,N_3304,N_2788);
and U6328 (N_6328,N_202,N_3771);
nand U6329 (N_6329,N_3516,N_4404);
xor U6330 (N_6330,N_4382,N_4038);
nand U6331 (N_6331,N_163,N_1946);
or U6332 (N_6332,N_1062,N_4965);
nand U6333 (N_6333,N_1759,N_870);
and U6334 (N_6334,N_4333,N_644);
and U6335 (N_6335,N_3363,N_2440);
or U6336 (N_6336,N_2768,N_4556);
nand U6337 (N_6337,N_3433,N_1619);
nor U6338 (N_6338,N_2402,N_1589);
nand U6339 (N_6339,N_4397,N_3949);
nor U6340 (N_6340,N_1558,N_294);
nor U6341 (N_6341,N_3557,N_1729);
nand U6342 (N_6342,N_2776,N_3018);
xor U6343 (N_6343,N_3004,N_81);
nor U6344 (N_6344,N_4849,N_43);
or U6345 (N_6345,N_2791,N_2246);
or U6346 (N_6346,N_3526,N_2414);
nor U6347 (N_6347,N_1894,N_1991);
and U6348 (N_6348,N_3489,N_992);
nand U6349 (N_6349,N_3506,N_2357);
nand U6350 (N_6350,N_1623,N_428);
or U6351 (N_6351,N_2592,N_1337);
and U6352 (N_6352,N_1427,N_2203);
nand U6353 (N_6353,N_3995,N_194);
or U6354 (N_6354,N_4838,N_3413);
nor U6355 (N_6355,N_239,N_4931);
nor U6356 (N_6356,N_4535,N_4289);
or U6357 (N_6357,N_4657,N_3556);
nand U6358 (N_6358,N_4452,N_4853);
and U6359 (N_6359,N_99,N_3037);
xnor U6360 (N_6360,N_4174,N_4803);
and U6361 (N_6361,N_4911,N_3400);
or U6362 (N_6362,N_1265,N_2799);
nor U6363 (N_6363,N_1693,N_1569);
nor U6364 (N_6364,N_3241,N_4906);
and U6365 (N_6365,N_2946,N_3893);
nor U6366 (N_6366,N_474,N_1817);
nor U6367 (N_6367,N_3719,N_980);
nor U6368 (N_6368,N_4932,N_115);
or U6369 (N_6369,N_1982,N_447);
or U6370 (N_6370,N_1943,N_4957);
and U6371 (N_6371,N_940,N_4939);
nor U6372 (N_6372,N_518,N_3355);
and U6373 (N_6373,N_2909,N_1336);
nor U6374 (N_6374,N_283,N_4557);
nor U6375 (N_6375,N_4348,N_422);
nand U6376 (N_6376,N_4831,N_1530);
nand U6377 (N_6377,N_974,N_3358);
xor U6378 (N_6378,N_517,N_2565);
nand U6379 (N_6379,N_4797,N_993);
nor U6380 (N_6380,N_3705,N_4489);
nor U6381 (N_6381,N_3943,N_1970);
nor U6382 (N_6382,N_3023,N_1506);
xnor U6383 (N_6383,N_4364,N_3555);
nor U6384 (N_6384,N_1617,N_2370);
or U6385 (N_6385,N_4126,N_2877);
and U6386 (N_6386,N_2952,N_4902);
and U6387 (N_6387,N_4856,N_2781);
or U6388 (N_6388,N_4293,N_80);
nor U6389 (N_6389,N_955,N_20);
xor U6390 (N_6390,N_884,N_2735);
or U6391 (N_6391,N_3085,N_11);
or U6392 (N_6392,N_4161,N_3005);
xnor U6393 (N_6393,N_2728,N_1898);
or U6394 (N_6394,N_3244,N_1383);
nor U6395 (N_6395,N_3593,N_808);
nor U6396 (N_6396,N_564,N_531);
or U6397 (N_6397,N_3581,N_1329);
nand U6398 (N_6398,N_3313,N_1358);
and U6399 (N_6399,N_2847,N_4889);
nand U6400 (N_6400,N_1700,N_1863);
nand U6401 (N_6401,N_4262,N_4030);
nor U6402 (N_6402,N_1335,N_4949);
xor U6403 (N_6403,N_3130,N_2703);
nand U6404 (N_6404,N_2438,N_3769);
nand U6405 (N_6405,N_1135,N_4850);
and U6406 (N_6406,N_1174,N_2400);
and U6407 (N_6407,N_2821,N_1085);
nand U6408 (N_6408,N_2956,N_2494);
nor U6409 (N_6409,N_1343,N_1531);
or U6410 (N_6410,N_2808,N_334);
nor U6411 (N_6411,N_4605,N_3929);
and U6412 (N_6412,N_2572,N_4473);
and U6413 (N_6413,N_4950,N_3958);
nand U6414 (N_6414,N_1665,N_3458);
or U6415 (N_6415,N_3902,N_3387);
nand U6416 (N_6416,N_3007,N_4141);
nor U6417 (N_6417,N_2180,N_4701);
nor U6418 (N_6418,N_2089,N_878);
and U6419 (N_6419,N_452,N_838);
nand U6420 (N_6420,N_2647,N_1829);
or U6421 (N_6421,N_1260,N_391);
or U6422 (N_6422,N_1989,N_4444);
and U6423 (N_6423,N_2783,N_1805);
nor U6424 (N_6424,N_4881,N_2846);
nor U6425 (N_6425,N_33,N_855);
nand U6426 (N_6426,N_3648,N_3336);
or U6427 (N_6427,N_4811,N_187);
xor U6428 (N_6428,N_1985,N_1611);
or U6429 (N_6429,N_305,N_4536);
nor U6430 (N_6430,N_1664,N_2164);
nor U6431 (N_6431,N_4835,N_3936);
nand U6432 (N_6432,N_2365,N_2318);
xor U6433 (N_6433,N_1851,N_296);
or U6434 (N_6434,N_3470,N_3917);
or U6435 (N_6435,N_2642,N_1727);
nor U6436 (N_6436,N_4639,N_2545);
and U6437 (N_6437,N_253,N_138);
xnor U6438 (N_6438,N_2923,N_4076);
or U6439 (N_6439,N_2656,N_1517);
nand U6440 (N_6440,N_2309,N_2998);
nand U6441 (N_6441,N_3135,N_1765);
and U6442 (N_6442,N_466,N_543);
nor U6443 (N_6443,N_1478,N_1706);
or U6444 (N_6444,N_1438,N_1857);
nand U6445 (N_6445,N_2403,N_4291);
nand U6446 (N_6446,N_4098,N_3749);
nand U6447 (N_6447,N_816,N_2610);
and U6448 (N_6448,N_1332,N_4265);
or U6449 (N_6449,N_1948,N_3612);
nor U6450 (N_6450,N_883,N_4834);
nand U6451 (N_6451,N_3584,N_755);
nand U6452 (N_6452,N_284,N_4681);
xnor U6453 (N_6453,N_1529,N_3817);
nand U6454 (N_6454,N_2903,N_3163);
and U6455 (N_6455,N_1891,N_4822);
and U6456 (N_6456,N_4762,N_3645);
or U6457 (N_6457,N_3599,N_3658);
and U6458 (N_6458,N_911,N_2353);
and U6459 (N_6459,N_4719,N_3752);
xnor U6460 (N_6460,N_1456,N_845);
nand U6461 (N_6461,N_4273,N_1692);
nor U6462 (N_6462,N_2418,N_2222);
nand U6463 (N_6463,N_4855,N_1328);
nand U6464 (N_6464,N_566,N_1900);
or U6465 (N_6465,N_4445,N_4528);
xnor U6466 (N_6466,N_4325,N_446);
nand U6467 (N_6467,N_2591,N_2528);
xor U6468 (N_6468,N_4568,N_4312);
and U6469 (N_6469,N_2268,N_2490);
nor U6470 (N_6470,N_4181,N_1078);
nand U6471 (N_6471,N_3544,N_1141);
or U6472 (N_6472,N_4000,N_807);
and U6473 (N_6473,N_2188,N_3738);
or U6474 (N_6474,N_4637,N_1273);
nand U6475 (N_6475,N_4597,N_1888);
and U6476 (N_6476,N_56,N_3802);
nand U6477 (N_6477,N_431,N_4516);
nor U6478 (N_6478,N_2425,N_1346);
xor U6479 (N_6479,N_498,N_1639);
nand U6480 (N_6480,N_2882,N_633);
nand U6481 (N_6481,N_2131,N_2407);
or U6482 (N_6482,N_3835,N_3524);
nor U6483 (N_6483,N_1022,N_967);
xnor U6484 (N_6484,N_3637,N_4183);
and U6485 (N_6485,N_1387,N_1969);
and U6486 (N_6486,N_4941,N_2071);
or U6487 (N_6487,N_520,N_1277);
nor U6488 (N_6488,N_3113,N_589);
nand U6489 (N_6489,N_467,N_3431);
nand U6490 (N_6490,N_3961,N_840);
or U6491 (N_6491,N_1788,N_1559);
nor U6492 (N_6492,N_4239,N_3934);
xnor U6493 (N_6493,N_3977,N_3967);
and U6494 (N_6494,N_2795,N_1878);
nand U6495 (N_6495,N_111,N_1583);
nor U6496 (N_6496,N_4120,N_1402);
nor U6497 (N_6497,N_4012,N_4974);
or U6498 (N_6498,N_1883,N_2868);
and U6499 (N_6499,N_3174,N_3001);
xor U6500 (N_6500,N_4180,N_3718);
and U6501 (N_6501,N_4936,N_519);
or U6502 (N_6502,N_4549,N_281);
or U6503 (N_6503,N_1393,N_4455);
nor U6504 (N_6504,N_865,N_4543);
nand U6505 (N_6505,N_1160,N_4378);
nor U6506 (N_6506,N_3875,N_3254);
xor U6507 (N_6507,N_3850,N_2106);
and U6508 (N_6508,N_3048,N_2580);
nand U6509 (N_6509,N_3301,N_934);
xnor U6510 (N_6510,N_4187,N_750);
nand U6511 (N_6511,N_104,N_2935);
and U6512 (N_6512,N_282,N_1836);
nand U6513 (N_6513,N_3015,N_2915);
nand U6514 (N_6514,N_882,N_2134);
nand U6515 (N_6515,N_1698,N_4157);
nand U6516 (N_6516,N_1751,N_1646);
nand U6517 (N_6517,N_2979,N_2670);
xor U6518 (N_6518,N_2212,N_3403);
and U6519 (N_6519,N_3715,N_1302);
and U6520 (N_6520,N_3217,N_360);
or U6521 (N_6521,N_2248,N_1379);
xor U6522 (N_6522,N_3918,N_1238);
nor U6523 (N_6523,N_711,N_3757);
nor U6524 (N_6524,N_966,N_3490);
and U6525 (N_6525,N_614,N_4844);
or U6526 (N_6526,N_2569,N_4449);
nand U6527 (N_6527,N_2039,N_1801);
nor U6528 (N_6528,N_3672,N_4708);
or U6529 (N_6529,N_2171,N_4980);
xor U6530 (N_6530,N_162,N_2653);
nand U6531 (N_6531,N_4002,N_1026);
nor U6532 (N_6532,N_1196,N_2453);
or U6533 (N_6533,N_790,N_1695);
nand U6534 (N_6534,N_2995,N_4418);
and U6535 (N_6535,N_1807,N_2560);
xor U6536 (N_6536,N_2756,N_3842);
nand U6537 (N_6537,N_3766,N_385);
or U6538 (N_6538,N_280,N_3500);
nor U6539 (N_6539,N_2458,N_725);
and U6540 (N_6540,N_4828,N_4424);
and U6541 (N_6541,N_4564,N_350);
nor U6542 (N_6542,N_328,N_256);
nand U6543 (N_6543,N_2065,N_2829);
or U6544 (N_6544,N_1913,N_3410);
and U6545 (N_6545,N_837,N_2444);
or U6546 (N_6546,N_4290,N_4052);
nor U6547 (N_6547,N_686,N_1871);
and U6548 (N_6548,N_2965,N_3781);
nand U6549 (N_6549,N_3108,N_4167);
nor U6550 (N_6550,N_731,N_1899);
or U6551 (N_6551,N_1756,N_761);
nand U6552 (N_6552,N_4519,N_2704);
nand U6553 (N_6553,N_2363,N_991);
and U6554 (N_6554,N_1467,N_3226);
xnor U6555 (N_6555,N_4946,N_3390);
nand U6556 (N_6556,N_3655,N_3488);
or U6557 (N_6557,N_1219,N_3706);
nor U6558 (N_6558,N_4552,N_3225);
nand U6559 (N_6559,N_238,N_470);
nand U6560 (N_6560,N_624,N_1068);
and U6561 (N_6561,N_2716,N_4345);
or U6562 (N_6562,N_2582,N_609);
nor U6563 (N_6563,N_1543,N_1104);
xnor U6564 (N_6564,N_4787,N_1971);
and U6565 (N_6565,N_1933,N_3759);
nand U6566 (N_6566,N_365,N_77);
or U6567 (N_6567,N_1492,N_1555);
and U6568 (N_6568,N_2327,N_703);
nor U6569 (N_6569,N_1905,N_1083);
nand U6570 (N_6570,N_4660,N_1571);
xor U6571 (N_6571,N_3955,N_4283);
nand U6572 (N_6572,N_1433,N_3216);
nand U6573 (N_6573,N_4506,N_2051);
nor U6574 (N_6574,N_546,N_706);
nand U6575 (N_6575,N_1593,N_1549);
and U6576 (N_6576,N_877,N_4479);
or U6577 (N_6577,N_3636,N_75);
nor U6578 (N_6578,N_2865,N_4553);
or U6579 (N_6579,N_3761,N_4644);
nor U6580 (N_6580,N_3029,N_2100);
and U6581 (N_6581,N_4747,N_3125);
or U6582 (N_6582,N_1957,N_3145);
nand U6583 (N_6583,N_2561,N_4201);
nor U6584 (N_6584,N_2064,N_2632);
nor U6585 (N_6585,N_605,N_601);
and U6586 (N_6586,N_2404,N_1109);
xnor U6587 (N_6587,N_4247,N_1212);
nand U6588 (N_6588,N_3510,N_1231);
or U6589 (N_6589,N_26,N_2651);
and U6590 (N_6590,N_998,N_1436);
nand U6591 (N_6591,N_4431,N_3856);
xnor U6592 (N_6592,N_170,N_3772);
or U6593 (N_6593,N_3014,N_4585);
or U6594 (N_6594,N_1108,N_1179);
or U6595 (N_6595,N_596,N_3389);
and U6596 (N_6596,N_307,N_52);
nand U6597 (N_6597,N_2659,N_184);
and U6598 (N_6598,N_1311,N_3529);
nand U6599 (N_6599,N_2381,N_4968);
and U6600 (N_6600,N_1304,N_949);
nand U6601 (N_6601,N_264,N_701);
or U6602 (N_6602,N_3992,N_2447);
nand U6603 (N_6603,N_2849,N_767);
nor U6604 (N_6604,N_2664,N_3064);
and U6605 (N_6605,N_4133,N_664);
nand U6606 (N_6606,N_4303,N_377);
and U6607 (N_6607,N_2511,N_3930);
or U6608 (N_6608,N_1481,N_683);
or U6609 (N_6609,N_2325,N_2567);
and U6610 (N_6610,N_401,N_3233);
xnor U6611 (N_6611,N_1046,N_4692);
or U6612 (N_6612,N_3560,N_1251);
xor U6613 (N_6613,N_114,N_1734);
nand U6614 (N_6614,N_4581,N_3229);
nand U6615 (N_6615,N_3097,N_4214);
and U6616 (N_6616,N_3799,N_4847);
nor U6617 (N_6617,N_3210,N_3768);
nor U6618 (N_6618,N_269,N_981);
xnor U6619 (N_6619,N_2499,N_2773);
xor U6620 (N_6620,N_2908,N_4574);
or U6621 (N_6621,N_2082,N_744);
xnor U6622 (N_6622,N_3571,N_3200);
or U6623 (N_6623,N_2838,N_4228);
or U6624 (N_6624,N_2990,N_3152);
and U6625 (N_6625,N_2252,N_1490);
xnor U6626 (N_6626,N_3129,N_4119);
or U6627 (N_6627,N_3747,N_3025);
and U6628 (N_6628,N_1964,N_1914);
nand U6629 (N_6629,N_3664,N_1636);
or U6630 (N_6630,N_765,N_1470);
nand U6631 (N_6631,N_4237,N_2011);
nand U6632 (N_6632,N_1831,N_3128);
or U6633 (N_6633,N_477,N_1535);
nand U6634 (N_6634,N_3993,N_2851);
nor U6635 (N_6635,N_2552,N_1161);
and U6636 (N_6636,N_3940,N_1115);
nand U6637 (N_6637,N_3659,N_1321);
nand U6638 (N_6638,N_2929,N_2415);
nor U6639 (N_6639,N_2897,N_2798);
nand U6640 (N_6640,N_2208,N_3617);
and U6641 (N_6641,N_3237,N_4502);
and U6642 (N_6642,N_4928,N_2978);
nor U6643 (N_6643,N_3282,N_1439);
nand U6644 (N_6644,N_3525,N_1345);
xnor U6645 (N_6645,N_866,N_3819);
and U6646 (N_6646,N_3798,N_4532);
or U6647 (N_6647,N_3377,N_2932);
or U6648 (N_6648,N_1718,N_1299);
or U6649 (N_6649,N_4271,N_1582);
and U6650 (N_6650,N_3388,N_4213);
and U6651 (N_6651,N_101,N_2157);
or U6652 (N_6652,N_2163,N_70);
and U6653 (N_6653,N_4571,N_2361);
nand U6654 (N_6654,N_216,N_1194);
or U6655 (N_6655,N_4841,N_175);
xor U6656 (N_6656,N_3493,N_3729);
and U6657 (N_6657,N_3957,N_2922);
or U6658 (N_6658,N_3273,N_4538);
nor U6659 (N_6659,N_3778,N_2380);
or U6660 (N_6660,N_729,N_3485);
and U6661 (N_6661,N_4563,N_182);
and U6662 (N_6662,N_950,N_960);
and U6663 (N_6663,N_1489,N_488);
nand U6664 (N_6664,N_1203,N_1784);
nand U6665 (N_6665,N_3972,N_2355);
nor U6666 (N_6666,N_4446,N_1993);
xor U6667 (N_6667,N_3642,N_511);
nor U6668 (N_6668,N_2482,N_2491);
and U6669 (N_6669,N_3351,N_2975);
xnor U6670 (N_6670,N_804,N_167);
and U6671 (N_6671,N_758,N_4468);
or U6672 (N_6672,N_3146,N_1005);
and U6673 (N_6673,N_3046,N_1710);
xnor U6674 (N_6674,N_1090,N_3812);
nor U6675 (N_6675,N_3622,N_370);
xnor U6676 (N_6676,N_3487,N_4337);
and U6677 (N_6677,N_2738,N_3626);
xnor U6678 (N_6678,N_3928,N_292);
and U6679 (N_6679,N_2046,N_2145);
and U6680 (N_6680,N_885,N_497);
xor U6681 (N_6681,N_49,N_2430);
nand U6682 (N_6682,N_4680,N_4070);
nor U6683 (N_6683,N_29,N_1036);
or U6684 (N_6684,N_3086,N_3385);
nand U6685 (N_6685,N_1849,N_4740);
or U6686 (N_6686,N_3847,N_2329);
or U6687 (N_6687,N_4282,N_2819);
or U6688 (N_6688,N_2426,N_844);
nor U6689 (N_6689,N_3946,N_3263);
nand U6690 (N_6690,N_2650,N_4704);
or U6691 (N_6691,N_1746,N_3087);
nand U6692 (N_6692,N_3912,N_2758);
or U6693 (N_6693,N_3746,N_3712);
nor U6694 (N_6694,N_2474,N_4152);
nor U6695 (N_6695,N_1266,N_3938);
nand U6696 (N_6696,N_4823,N_1512);
and U6697 (N_6697,N_1452,N_4075);
and U6698 (N_6698,N_2120,N_1177);
and U6699 (N_6699,N_173,N_2184);
and U6700 (N_6700,N_4045,N_2253);
nor U6701 (N_6701,N_2880,N_4554);
xnor U6702 (N_6702,N_1918,N_3350);
nand U6703 (N_6703,N_3091,N_2588);
and U6704 (N_6704,N_4515,N_1973);
xnor U6705 (N_6705,N_4379,N_437);
and U6706 (N_6706,N_340,N_3184);
nor U6707 (N_6707,N_4859,N_2174);
nor U6708 (N_6708,N_464,N_4231);
nand U6709 (N_6709,N_3287,N_2549);
and U6710 (N_6710,N_3570,N_924);
and U6711 (N_6711,N_2953,N_3373);
or U6712 (N_6712,N_2345,N_4588);
and U6713 (N_6713,N_3073,N_2317);
nor U6714 (N_6714,N_2754,N_2556);
and U6715 (N_6715,N_298,N_1442);
nor U6716 (N_6716,N_1205,N_2257);
nand U6717 (N_6717,N_500,N_2334);
or U6718 (N_6718,N_3950,N_3223);
xnor U6719 (N_6719,N_1600,N_3399);
nand U6720 (N_6720,N_2804,N_4584);
nor U6721 (N_6721,N_3356,N_4706);
nor U6722 (N_6722,N_3397,N_2472);
or U6723 (N_6723,N_3583,N_4654);
or U6724 (N_6724,N_4481,N_628);
xnor U6725 (N_6725,N_2072,N_3055);
nand U6726 (N_6726,N_2084,N_599);
nand U6727 (N_6727,N_4967,N_1987);
nand U6728 (N_6728,N_1440,N_199);
or U6729 (N_6729,N_908,N_1785);
and U6730 (N_6730,N_4575,N_1561);
nor U6731 (N_6731,N_3404,N_4760);
nand U6732 (N_6732,N_4956,N_2822);
and U6733 (N_6733,N_1915,N_2262);
and U6734 (N_6734,N_4551,N_3882);
or U6735 (N_6735,N_3195,N_451);
nand U6736 (N_6736,N_1563,N_1866);
nand U6737 (N_6737,N_3927,N_3620);
or U6738 (N_6738,N_3858,N_3245);
nand U6739 (N_6739,N_2937,N_3649);
or U6740 (N_6740,N_2154,N_2247);
nor U6741 (N_6741,N_2760,N_4286);
and U6742 (N_6742,N_3154,N_403);
nor U6743 (N_6743,N_971,N_4034);
nor U6744 (N_6744,N_4151,N_4085);
nand U6745 (N_6745,N_718,N_2295);
nand U6746 (N_6746,N_3058,N_2510);
nand U6747 (N_6747,N_61,N_1992);
nor U6748 (N_6748,N_2242,N_4872);
or U6749 (N_6749,N_3844,N_35);
nor U6750 (N_6750,N_1324,N_936);
nor U6751 (N_6751,N_1628,N_2281);
nor U6752 (N_6752,N_783,N_509);
nor U6753 (N_6753,N_3849,N_4788);
nor U6754 (N_6754,N_69,N_4482);
xor U6755 (N_6755,N_4500,N_472);
nor U6756 (N_6756,N_2166,N_530);
nand U6757 (N_6757,N_2564,N_2982);
nand U6758 (N_6758,N_1916,N_512);
nand U6759 (N_6759,N_1681,N_41);
or U6760 (N_6760,N_3924,N_2399);
or U6761 (N_6761,N_3038,N_3968);
nor U6762 (N_6762,N_1129,N_353);
nor U6763 (N_6763,N_3308,N_3565);
nor U6764 (N_6764,N_120,N_1291);
nand U6765 (N_6765,N_2016,N_604);
and U6766 (N_6766,N_1794,N_3189);
or U6767 (N_6767,N_4236,N_3412);
nand U6768 (N_6768,N_2815,N_2700);
or U6769 (N_6769,N_88,N_2019);
and U6770 (N_6770,N_4507,N_3807);
nand U6771 (N_6771,N_3945,N_1626);
and U6772 (N_6772,N_3201,N_4287);
nand U6773 (N_6773,N_4975,N_4698);
or U6774 (N_6774,N_4042,N_2475);
or U6775 (N_6775,N_2443,N_2179);
nand U6776 (N_6776,N_2331,N_3870);
nor U6777 (N_6777,N_4258,N_3603);
nor U6778 (N_6778,N_4135,N_4503);
nor U6779 (N_6779,N_3116,N_3990);
or U6780 (N_6780,N_3989,N_430);
nor U6781 (N_6781,N_4943,N_4891);
nor U6782 (N_6782,N_1819,N_4018);
nor U6783 (N_6783,N_4438,N_2748);
nand U6784 (N_6784,N_95,N_1152);
and U6785 (N_6785,N_1034,N_667);
nor U6786 (N_6786,N_976,N_2844);
nand U6787 (N_6787,N_2657,N_1988);
and U6788 (N_6788,N_4774,N_3780);
nor U6789 (N_6789,N_3730,N_858);
and U6790 (N_6790,N_3947,N_603);
xnor U6791 (N_6791,N_4582,N_1303);
or U6792 (N_6792,N_2129,N_4067);
nand U6793 (N_6793,N_4874,N_2755);
nand U6794 (N_6794,N_3122,N_1391);
xnor U6795 (N_6795,N_1956,N_404);
or U6796 (N_6796,N_1118,N_1286);
and U6797 (N_6797,N_3630,N_177);
or U6798 (N_6798,N_4561,N_4798);
and U6799 (N_6799,N_191,N_938);
or U6800 (N_6800,N_1832,N_1023);
nor U6801 (N_6801,N_2554,N_475);
or U6802 (N_6802,N_3770,N_1151);
xnor U6803 (N_6803,N_1069,N_2160);
nor U6804 (N_6804,N_3970,N_379);
nand U6805 (N_6805,N_1367,N_439);
or U6806 (N_6806,N_1990,N_4935);
nor U6807 (N_6807,N_2041,N_141);
nor U6808 (N_6808,N_4062,N_875);
or U6809 (N_6809,N_3398,N_2273);
nand U6810 (N_6810,N_2236,N_1453);
nand U6811 (N_6811,N_2725,N_4198);
and U6812 (N_6812,N_1259,N_4985);
and U6813 (N_6813,N_1828,N_2695);
or U6814 (N_6814,N_2315,N_3743);
nor U6815 (N_6815,N_1209,N_3285);
nand U6816 (N_6816,N_1312,N_3321);
xnor U6817 (N_6817,N_2581,N_4377);
and U6818 (N_6818,N_1952,N_102);
nand U6819 (N_6819,N_4659,N_698);
and U6820 (N_6820,N_2692,N_2121);
nor U6821 (N_6821,N_3024,N_3527);
or U6822 (N_6822,N_567,N_0);
or U6823 (N_6823,N_36,N_2753);
nand U6824 (N_6824,N_1865,N_832);
and U6825 (N_6825,N_266,N_1875);
xor U6826 (N_6826,N_1942,N_749);
nand U6827 (N_6827,N_3999,N_1446);
nor U6828 (N_6828,N_174,N_3418);
nor U6829 (N_6829,N_3192,N_3247);
nand U6830 (N_6830,N_1220,N_3297);
or U6831 (N_6831,N_578,N_1041);
nor U6832 (N_6832,N_4591,N_1998);
and U6833 (N_6833,N_4586,N_717);
and U6834 (N_6834,N_3481,N_2319);
nand U6835 (N_6835,N_2496,N_1981);
and U6836 (N_6836,N_2122,N_1071);
and U6837 (N_6837,N_448,N_3963);
nor U6838 (N_6838,N_1815,N_1594);
nor U6839 (N_6839,N_1947,N_887);
xor U6840 (N_6840,N_1307,N_621);
and U6841 (N_6841,N_1269,N_1175);
nor U6842 (N_6842,N_3804,N_2540);
and U6843 (N_6843,N_3396,N_2385);
and U6844 (N_6844,N_2010,N_1523);
or U6845 (N_6845,N_2312,N_4996);
or U6846 (N_6846,N_3919,N_1077);
xnor U6847 (N_6847,N_4619,N_4703);
and U6848 (N_6848,N_1937,N_958);
xnor U6849 (N_6849,N_972,N_1755);
nor U6850 (N_6850,N_226,N_710);
nor U6851 (N_6851,N_538,N_4020);
or U6852 (N_6852,N_1314,N_1939);
and U6853 (N_6853,N_4604,N_3901);
or U6854 (N_6854,N_997,N_3701);
and U6855 (N_6855,N_1722,N_349);
nor U6856 (N_6856,N_2873,N_532);
or U6857 (N_6857,N_2442,N_576);
or U6858 (N_6858,N_4168,N_478);
nand U6859 (N_6859,N_2349,N_2628);
nor U6860 (N_6860,N_2707,N_2477);
and U6861 (N_6861,N_2213,N_3119);
nand U6862 (N_6862,N_501,N_1268);
nor U6863 (N_6863,N_4146,N_1651);
and U6864 (N_6864,N_2178,N_395);
nand U6865 (N_6865,N_722,N_1079);
nand U6866 (N_6866,N_2750,N_4005);
or U6867 (N_6867,N_2136,N_31);
nand U6868 (N_6868,N_2351,N_471);
nor U6869 (N_6869,N_4365,N_4885);
and U6870 (N_6870,N_3270,N_2285);
and U6871 (N_6871,N_3003,N_1844);
nor U6872 (N_6872,N_2190,N_4712);
or U6873 (N_6873,N_577,N_2207);
xnor U6874 (N_6874,N_4130,N_3613);
and U6875 (N_6875,N_3380,N_3012);
nand U6876 (N_6876,N_4814,N_3725);
or U6877 (N_6877,N_398,N_3197);
nor U6878 (N_6878,N_2047,N_2302);
and U6879 (N_6879,N_2993,N_3456);
and U6880 (N_6880,N_1465,N_3480);
nor U6881 (N_6881,N_1017,N_2489);
and U6882 (N_6882,N_2596,N_984);
and U6883 (N_6883,N_1339,N_1677);
or U6884 (N_6884,N_3257,N_4280);
nor U6885 (N_6885,N_2096,N_2014);
nor U6886 (N_6886,N_4113,N_4697);
xor U6887 (N_6887,N_918,N_2974);
and U6888 (N_6888,N_2232,N_387);
nor U6889 (N_6889,N_2519,N_4035);
xor U6890 (N_6890,N_2600,N_1000);
nand U6891 (N_6891,N_630,N_3165);
nor U6892 (N_6892,N_3215,N_71);
or U6893 (N_6893,N_1625,N_3459);
or U6894 (N_6894,N_1653,N_3872);
nor U6895 (N_6895,N_4322,N_3660);
xnor U6896 (N_6896,N_1243,N_2631);
nor U6897 (N_6897,N_3096,N_1325);
or U6898 (N_6898,N_2059,N_1290);
nand U6899 (N_6899,N_4109,N_3212);
and U6900 (N_6900,N_2260,N_4003);
or U6901 (N_6901,N_4025,N_237);
and U6902 (N_6902,N_4801,N_2970);
nand U6903 (N_6903,N_67,N_2405);
nand U6904 (N_6904,N_849,N_1632);
or U6905 (N_6905,N_2553,N_4945);
and U6906 (N_6906,N_977,N_4748);
nand U6907 (N_6907,N_843,N_3464);
nor U6908 (N_6908,N_3067,N_2533);
xnor U6909 (N_6909,N_3671,N_2448);
nor U6910 (N_6910,N_3507,N_359);
or U6911 (N_6911,N_3697,N_2826);
xnor U6912 (N_6912,N_1404,N_1051);
or U6913 (N_6913,N_4252,N_3634);
nor U6914 (N_6914,N_2688,N_3670);
or U6915 (N_6915,N_1171,N_3744);
or U6916 (N_6916,N_2081,N_3322);
nor U6917 (N_6917,N_3773,N_4319);
or U6918 (N_6918,N_1363,N_1797);
or U6919 (N_6919,N_4440,N_1236);
nor U6920 (N_6920,N_2112,N_3098);
or U6921 (N_6921,N_3643,N_3072);
nor U6922 (N_6922,N_2769,N_553);
or U6923 (N_6923,N_3745,N_759);
or U6924 (N_6924,N_3211,N_1887);
nor U6925 (N_6925,N_3027,N_244);
or U6926 (N_6926,N_1634,N_1649);
nor U6927 (N_6927,N_4139,N_3238);
or U6928 (N_6928,N_3806,N_2957);
and U6929 (N_6929,N_1599,N_4100);
xor U6930 (N_6930,N_3050,N_3199);
nor U6931 (N_6931,N_3332,N_2306);
and U6932 (N_6932,N_504,N_1496);
and U6933 (N_6933,N_3335,N_4815);
nand U6934 (N_6934,N_2439,N_3115);
nand U6935 (N_6935,N_4308,N_1334);
or U6936 (N_6936,N_678,N_12);
or U6937 (N_6937,N_1125,N_245);
nor U6938 (N_6938,N_1322,N_1039);
xnor U6939 (N_6939,N_631,N_4738);
and U6940 (N_6940,N_3249,N_2891);
and U6941 (N_6941,N_1965,N_4304);
and U6942 (N_6942,N_1732,N_3792);
or U6943 (N_6943,N_4775,N_60);
or U6944 (N_6944,N_1827,N_1654);
nand U6945 (N_6945,N_957,N_3708);
or U6946 (N_6946,N_3317,N_4682);
nor U6947 (N_6947,N_2251,N_2579);
and U6948 (N_6948,N_3820,N_1047);
nor U6949 (N_6949,N_4154,N_1112);
nor U6950 (N_6950,N_1570,N_3754);
or U6951 (N_6951,N_3342,N_4381);
nand U6952 (N_6952,N_2030,N_3136);
nand U6953 (N_6953,N_947,N_1684);
or U6954 (N_6954,N_3784,N_2731);
or U6955 (N_6955,N_2945,N_4408);
or U6956 (N_6956,N_4032,N_4212);
nand U6957 (N_6957,N_3793,N_3944);
xnor U6958 (N_6958,N_4858,N_3465);
and U6959 (N_6959,N_4315,N_2234);
nand U6960 (N_6960,N_4254,N_4118);
and U6961 (N_6961,N_2419,N_373);
or U6962 (N_6962,N_1011,N_2621);
nor U6963 (N_6963,N_3357,N_4688);
or U6964 (N_6964,N_1037,N_4349);
and U6965 (N_6965,N_1813,N_814);
and U6966 (N_6966,N_2732,N_4240);
and U6967 (N_6967,N_2708,N_2364);
nand U6968 (N_6968,N_1276,N_697);
nand U6969 (N_6969,N_4534,N_3683);
or U6970 (N_6970,N_4177,N_4336);
nand U6971 (N_6971,N_3028,N_1920);
nand U6972 (N_6972,N_1250,N_4116);
nand U6973 (N_6973,N_1048,N_4817);
and U6974 (N_6974,N_2607,N_4281);
or U6975 (N_6975,N_4839,N_3222);
nor U6976 (N_6976,N_2525,N_1070);
xor U6977 (N_6977,N_4495,N_1752);
and U6978 (N_6978,N_3767,N_1451);
nor U6979 (N_6979,N_754,N_2124);
xor U6980 (N_6980,N_4915,N_892);
and U6981 (N_6981,N_3959,N_2764);
or U6982 (N_6982,N_4923,N_259);
xor U6983 (N_6983,N_1711,N_116);
nand U6984 (N_6984,N_250,N_3354);
and U6985 (N_6985,N_1257,N_4819);
and U6986 (N_6986,N_4840,N_580);
nor U6987 (N_6987,N_813,N_1120);
nand U6988 (N_6988,N_1201,N_1853);
nor U6989 (N_6989,N_2000,N_2925);
or U6990 (N_6990,N_3550,N_3656);
and U6991 (N_6991,N_1215,N_1418);
nand U6992 (N_6992,N_3175,N_1702);
or U6993 (N_6993,N_3987,N_3148);
and U6994 (N_6994,N_4869,N_2779);
or U6995 (N_6995,N_4142,N_1767);
or U6996 (N_6996,N_1038,N_4513);
or U6997 (N_6997,N_1348,N_3573);
nor U6998 (N_6998,N_2436,N_4185);
and U6999 (N_6999,N_1867,N_384);
and U7000 (N_7000,N_3370,N_1074);
nand U7001 (N_7001,N_344,N_2931);
or U7002 (N_7002,N_4695,N_1686);
and U7003 (N_7003,N_1605,N_670);
nand U7004 (N_7004,N_3800,N_2907);
nand U7005 (N_7005,N_2300,N_3158);
and U7006 (N_7006,N_3702,N_72);
and U7007 (N_7007,N_2635,N_44);
and U7008 (N_7008,N_3627,N_3089);
and U7009 (N_7009,N_3829,N_3551);
xor U7010 (N_7010,N_1371,N_1642);
nor U7011 (N_7011,N_4245,N_3580);
nand U7012 (N_7012,N_4900,N_818);
or U7013 (N_7013,N_2555,N_2110);
nor U7014 (N_7014,N_1032,N_4577);
xor U7015 (N_7015,N_3062,N_3623);
and U7016 (N_7016,N_3932,N_2140);
nand U7017 (N_7017,N_4430,N_96);
xnor U7018 (N_7018,N_4799,N_4048);
nor U7019 (N_7019,N_3194,N_3034);
xnor U7020 (N_7020,N_3099,N_937);
or U7021 (N_7021,N_1566,N_1099);
and U7022 (N_7022,N_4944,N_2210);
or U7023 (N_7023,N_513,N_647);
and U7024 (N_7024,N_1524,N_4307);
nand U7025 (N_7025,N_2547,N_2717);
or U7026 (N_7026,N_4394,N_4171);
and U7027 (N_7027,N_806,N_1082);
or U7028 (N_7028,N_4691,N_1294);
nand U7029 (N_7029,N_733,N_2630);
nand U7030 (N_7030,N_930,N_1515);
nand U7031 (N_7031,N_3887,N_3494);
or U7032 (N_7032,N_4435,N_4372);
nand U7033 (N_7033,N_839,N_4205);
nor U7034 (N_7034,N_3602,N_2714);
nand U7035 (N_7035,N_1963,N_479);
nor U7036 (N_7036,N_4234,N_3717);
and U7037 (N_7037,N_3855,N_4129);
nand U7038 (N_7038,N_107,N_2366);
nor U7039 (N_7039,N_906,N_215);
nand U7040 (N_7040,N_4655,N_978);
nor U7041 (N_7041,N_367,N_3598);
nor U7042 (N_7042,N_1441,N_4667);
nand U7043 (N_7043,N_390,N_2535);
nor U7044 (N_7044,N_1374,N_2971);
nand U7045 (N_7045,N_3511,N_4726);
and U7046 (N_7046,N_1892,N_3794);
nor U7047 (N_7047,N_2410,N_2669);
or U7048 (N_7048,N_3640,N_3791);
and U7049 (N_7049,N_3371,N_2766);
nand U7050 (N_7050,N_4696,N_1253);
nand U7051 (N_7051,N_2261,N_1480);
nand U7052 (N_7052,N_1224,N_4059);
and U7053 (N_7053,N_1554,N_1340);
or U7054 (N_7054,N_4188,N_623);
nand U7055 (N_7055,N_291,N_3951);
nor U7056 (N_7056,N_1822,N_2293);
nand U7057 (N_7057,N_2107,N_134);
and U7058 (N_7058,N_4356,N_668);
or U7059 (N_7059,N_2902,N_3416);
or U7060 (N_7060,N_3874,N_1455);
nor U7061 (N_7061,N_3574,N_3906);
nand U7062 (N_7062,N_419,N_3971);
nor U7063 (N_7063,N_850,N_2033);
nor U7064 (N_7064,N_4211,N_645);
or U7065 (N_7065,N_3376,N_4341);
or U7066 (N_7066,N_3795,N_4602);
nand U7067 (N_7067,N_4371,N_3094);
xor U7068 (N_7068,N_651,N_1793);
nor U7069 (N_7069,N_4754,N_854);
nor U7070 (N_7070,N_3143,N_3942);
or U7071 (N_7071,N_2741,N_3020);
and U7072 (N_7072,N_1488,N_2649);
nand U7073 (N_7073,N_3181,N_2254);
xnor U7074 (N_7074,N_3988,N_3461);
or U7075 (N_7075,N_2614,N_4015);
and U7076 (N_7076,N_2393,N_3284);
xor U7077 (N_7077,N_1877,N_1712);
or U7078 (N_7078,N_16,N_150);
or U7079 (N_7079,N_2888,N_4583);
xor U7080 (N_7080,N_2138,N_2265);
xor U7081 (N_7081,N_4275,N_4387);
nand U7082 (N_7082,N_208,N_2671);
nand U7083 (N_7083,N_2684,N_2542);
nand U7084 (N_7084,N_1738,N_3857);
and U7085 (N_7085,N_1714,N_552);
and U7086 (N_7086,N_3589,N_3047);
nor U7087 (N_7087,N_4661,N_907);
and U7088 (N_7088,N_1318,N_3168);
and U7089 (N_7089,N_902,N_2532);
xor U7090 (N_7090,N_2052,N_3466);
xnor U7091 (N_7091,N_1730,N_3814);
xnor U7092 (N_7092,N_1204,N_1839);
and U7093 (N_7093,N_1106,N_469);
nor U7094 (N_7094,N_4134,N_4115);
nor U7095 (N_7095,N_4629,N_484);
nand U7096 (N_7096,N_1858,N_2722);
and U7097 (N_7097,N_2379,N_4573);
or U7098 (N_7098,N_3528,N_533);
nor U7099 (N_7099,N_3533,N_2924);
xor U7100 (N_7100,N_514,N_3615);
nand U7101 (N_7101,N_1984,N_1737);
or U7102 (N_7102,N_1974,N_2083);
nand U7103 (N_7103,N_797,N_909);
and U7104 (N_7104,N_3568,N_2111);
and U7105 (N_7105,N_1381,N_3272);
xnor U7106 (N_7106,N_640,N_476);
xnor U7107 (N_7107,N_2950,N_2005);
or U7108 (N_7108,N_2088,N_2283);
or U7109 (N_7109,N_1977,N_742);
nand U7110 (N_7110,N_1775,N_4395);
xor U7111 (N_7111,N_3833,N_3204);
and U7112 (N_7112,N_1376,N_3295);
nor U7113 (N_7113,N_51,N_4649);
and U7114 (N_7114,N_4053,N_2817);
and U7115 (N_7115,N_1724,N_1553);
nand U7116 (N_7116,N_2701,N_2191);
and U7117 (N_7117,N_3797,N_1016);
nand U7118 (N_7118,N_4432,N_4792);
and U7119 (N_7119,N_210,N_3537);
nor U7120 (N_7120,N_4830,N_687);
nor U7121 (N_7121,N_1437,N_143);
or U7122 (N_7122,N_956,N_3601);
nor U7123 (N_7123,N_3689,N_846);
nand U7124 (N_7124,N_196,N_3859);
xor U7125 (N_7125,N_2878,N_2502);
nand U7126 (N_7126,N_4274,N_3309);
and U7127 (N_7127,N_2148,N_4509);
nor U7128 (N_7128,N_1349,N_709);
xnor U7129 (N_7129,N_506,N_791);
nor U7130 (N_7130,N_2859,N_2713);
nor U7131 (N_7131,N_1790,N_691);
and U7132 (N_7132,N_343,N_3885);
or U7133 (N_7133,N_396,N_1504);
or U7134 (N_7134,N_1020,N_400);
xnor U7135 (N_7135,N_2988,N_656);
nor U7136 (N_7136,N_1592,N_800);
nor U7137 (N_7137,N_3324,N_4243);
or U7138 (N_7138,N_318,N_2155);
nand U7139 (N_7139,N_2509,N_4645);
or U7140 (N_7140,N_1049,N_2624);
or U7141 (N_7141,N_17,N_1434);
and U7142 (N_7142,N_2288,N_4559);
nand U7143 (N_7143,N_4140,N_4933);
nor U7144 (N_7144,N_547,N_4277);
nor U7145 (N_7145,N_2420,N_2484);
and U7146 (N_7146,N_84,N_2237);
or U7147 (N_7147,N_4099,N_4725);
or U7148 (N_7148,N_665,N_2658);
nor U7149 (N_7149,N_1959,N_4299);
nand U7150 (N_7150,N_1241,N_3040);
xnor U7151 (N_7151,N_4794,N_3765);
and U7152 (N_7152,N_4672,N_1766);
nand U7153 (N_7153,N_505,N_2023);
or U7154 (N_7154,N_2980,N_304);
nand U7155 (N_7155,N_2710,N_4930);
nand U7156 (N_7156,N_3361,N_2685);
nand U7157 (N_7157,N_495,N_1770);
nor U7158 (N_7158,N_1873,N_3314);
nand U7159 (N_7159,N_234,N_4662);
nand U7160 (N_7160,N_303,N_1689);
xor U7161 (N_7161,N_3984,N_3294);
or U7162 (N_7162,N_1095,N_4222);
nand U7163 (N_7163,N_2149,N_3501);
xor U7164 (N_7164,N_1094,N_4942);
nor U7165 (N_7165,N_4486,N_1912);
nor U7166 (N_7166,N_1246,N_4155);
nand U7167 (N_7167,N_3127,N_876);
or U7168 (N_7168,N_4510,N_2343);
nand U7169 (N_7169,N_2578,N_2637);
nand U7170 (N_7170,N_2802,N_607);
nor U7171 (N_7171,N_2354,N_2852);
and U7172 (N_7172,N_3435,N_436);
nor U7173 (N_7173,N_2063,N_4728);
nand U7174 (N_7174,N_586,N_1354);
or U7175 (N_7175,N_3755,N_2424);
and U7176 (N_7176,N_2085,N_541);
and U7177 (N_7177,N_190,N_3149);
or U7178 (N_7178,N_1173,N_311);
xnor U7179 (N_7179,N_2053,N_4603);
nand U7180 (N_7180,N_3756,N_2457);
nor U7181 (N_7181,N_3624,N_4592);
nor U7182 (N_7182,N_2668,N_481);
or U7183 (N_7183,N_267,N_18);
or U7184 (N_7184,N_1100,N_4607);
or U7185 (N_7185,N_4504,N_4330);
or U7186 (N_7186,N_168,N_2192);
xor U7187 (N_7187,N_3948,N_454);
and U7188 (N_7188,N_777,N_4979);
or U7189 (N_7189,N_3441,N_528);
and U7190 (N_7190,N_890,N_382);
nand U7191 (N_7191,N_4001,N_3150);
nand U7192 (N_7192,N_1910,N_4761);
and U7193 (N_7193,N_2189,N_4172);
xnor U7194 (N_7194,N_4199,N_4783);
xor U7195 (N_7195,N_1880,N_1771);
nor U7196 (N_7196,N_1235,N_3330);
and U7197 (N_7197,N_694,N_25);
and U7198 (N_7198,N_2594,N_2043);
or U7199 (N_7199,N_2739,N_2002);
and U7200 (N_7200,N_231,N_2021);
xnor U7201 (N_7201,N_4580,N_4060);
xor U7202 (N_7202,N_2992,N_3575);
nand U7203 (N_7203,N_1024,N_4132);
or U7204 (N_7204,N_4904,N_4884);
nor U7205 (N_7205,N_2015,N_4997);
and U7206 (N_7206,N_2230,N_1107);
or U7207 (N_7207,N_3588,N_2389);
nor U7208 (N_7208,N_570,N_1365);
nand U7209 (N_7209,N_265,N_4106);
or U7210 (N_7210,N_4492,N_695);
nor U7211 (N_7211,N_4039,N_2983);
nor U7212 (N_7212,N_1293,N_3405);
nand U7213 (N_7213,N_968,N_3107);
nand U7214 (N_7214,N_4210,N_1890);
xnor U7215 (N_7215,N_1764,N_2175);
or U7216 (N_7216,N_4984,N_2881);
or U7217 (N_7217,N_2274,N_4633);
nor U7218 (N_7218,N_2794,N_4112);
nand U7219 (N_7219,N_1615,N_121);
nand U7220 (N_7220,N_3170,N_4317);
and U7221 (N_7221,N_2497,N_112);
nor U7222 (N_7222,N_1949,N_125);
nor U7223 (N_7223,N_4587,N_329);
and U7224 (N_7224,N_1613,N_2151);
nor U7225 (N_7225,N_2342,N_1747);
nand U7226 (N_7226,N_2452,N_2955);
nand U7227 (N_7227,N_297,N_3614);
nand U7228 (N_7228,N_2371,N_637);
nor U7229 (N_7229,N_4300,N_642);
xnor U7230 (N_7230,N_2944,N_3126);
or U7231 (N_7231,N_3153,N_2153);
nand U7232 (N_7232,N_288,N_563);
and U7233 (N_7233,N_3030,N_3248);
nand U7234 (N_7234,N_2850,N_2949);
nand U7235 (N_7235,N_912,N_2132);
or U7236 (N_7236,N_862,N_426);
nor U7237 (N_7237,N_1230,N_4796);
and U7238 (N_7238,N_4784,N_4683);
nor U7239 (N_7239,N_3662,N_3269);
or U7240 (N_7240,N_3155,N_4865);
or U7241 (N_7241,N_2619,N_1195);
or U7242 (N_7242,N_4751,N_2885);
nand U7243 (N_7243,N_1601,N_1647);
nand U7244 (N_7244,N_1742,N_2889);
and U7245 (N_7245,N_2997,N_2597);
nand U7246 (N_7246,N_3590,N_140);
or U7247 (N_7247,N_893,N_3826);
nor U7248 (N_7248,N_1035,N_46);
nand U7249 (N_7249,N_4416,N_227);
and U7250 (N_7250,N_1145,N_3049);
or U7251 (N_7251,N_3101,N_2152);
or U7252 (N_7252,N_4846,N_2655);
or U7253 (N_7253,N_2067,N_3616);
nor U7254 (N_7254,N_1986,N_2326);
nor U7255 (N_7255,N_1843,N_1967);
nand U7256 (N_7256,N_424,N_2848);
nor U7257 (N_7257,N_160,N_1659);
xnor U7258 (N_7258,N_126,N_3737);
xor U7259 (N_7259,N_106,N_4403);
or U7260 (N_7260,N_57,N_74);
nand U7261 (N_7261,N_4567,N_1150);
nand U7262 (N_7262,N_4465,N_320);
nor U7263 (N_7263,N_3471,N_4178);
or U7264 (N_7264,N_206,N_2845);
nand U7265 (N_7265,N_815,N_4572);
nor U7266 (N_7266,N_4753,N_4616);
nand U7267 (N_7267,N_1495,N_4626);
and U7268 (N_7268,N_157,N_648);
nor U7269 (N_7269,N_1287,N_2759);
nand U7270 (N_7270,N_2004,N_746);
nand U7271 (N_7271,N_355,N_1188);
or U7272 (N_7272,N_898,N_1426);
or U7273 (N_7273,N_1538,N_2818);
and U7274 (N_7274,N_3156,N_4631);
or U7275 (N_7275,N_366,N_3346);
or U7276 (N_7276,N_663,N_2629);
nor U7277 (N_7277,N_3235,N_880);
nand U7278 (N_7278,N_312,N_221);
and U7279 (N_7279,N_242,N_3251);
nand U7280 (N_7280,N_2267,N_1222);
nand U7281 (N_7281,N_3851,N_2839);
nor U7282 (N_7282,N_1285,N_662);
nor U7283 (N_7283,N_894,N_201);
and U7284 (N_7284,N_616,N_4158);
or U7285 (N_7285,N_3728,N_147);
nor U7286 (N_7286,N_784,N_113);
or U7287 (N_7287,N_4491,N_2620);
nand U7288 (N_7288,N_2752,N_2730);
nand U7289 (N_7289,N_3011,N_2034);
nand U7290 (N_7290,N_762,N_1447);
nand U7291 (N_7291,N_3710,N_3734);
nand U7292 (N_7292,N_4215,N_1009);
nor U7293 (N_7293,N_1010,N_3437);
xnor U7294 (N_7294,N_2905,N_3451);
and U7295 (N_7295,N_405,N_2434);
nand U7296 (N_7296,N_2133,N_3234);
or U7297 (N_7297,N_381,N_4710);
nand U7298 (N_7298,N_2250,N_1469);
and U7299 (N_7299,N_491,N_2313);
and U7300 (N_7300,N_2470,N_1781);
xnor U7301 (N_7301,N_308,N_2187);
nor U7302 (N_7302,N_3549,N_1719);
nor U7303 (N_7303,N_871,N_4011);
nor U7304 (N_7304,N_136,N_853);
or U7305 (N_7305,N_37,N_2012);
nand U7306 (N_7306,N_2855,N_4361);
nand U7307 (N_7307,N_1275,N_3009);
nand U7308 (N_7308,N_4136,N_3298);
or U7309 (N_7309,N_925,N_4021);
and U7310 (N_7310,N_2301,N_860);
nor U7311 (N_7311,N_1366,N_4589);
or U7312 (N_7312,N_986,N_2720);
or U7313 (N_7313,N_1378,N_2495);
and U7314 (N_7314,N_3716,N_4498);
nor U7315 (N_7315,N_3103,N_1114);
and U7316 (N_7316,N_2639,N_562);
nor U7317 (N_7317,N_1131,N_4413);
nand U7318 (N_7318,N_867,N_2523);
or U7319 (N_7319,N_2079,N_3231);
and U7320 (N_7320,N_4768,N_781);
nand U7321 (N_7321,N_4373,N_3891);
xor U7322 (N_7322,N_3384,N_2586);
or U7323 (N_7323,N_3823,N_2462);
nor U7324 (N_7324,N_348,N_103);
or U7325 (N_7325,N_249,N_4366);
xor U7326 (N_7326,N_1463,N_213);
or U7327 (N_7327,N_1906,N_1745);
nor U7328 (N_7328,N_3207,N_3462);
xor U7329 (N_7329,N_2276,N_1631);
nand U7330 (N_7330,N_4813,N_568);
nor U7331 (N_7331,N_4636,N_2623);
and U7332 (N_7332,N_1165,N_4114);
or U7333 (N_7333,N_4973,N_3911);
and U7334 (N_7334,N_2087,N_899);
nor U7335 (N_7335,N_499,N_970);
nor U7336 (N_7336,N_1044,N_2483);
nor U7337 (N_7337,N_4342,N_4882);
or U7338 (N_7338,N_4546,N_1680);
xnor U7339 (N_7339,N_4836,N_598);
or U7340 (N_7340,N_2718,N_2091);
nor U7341 (N_7341,N_59,N_1792);
nand U7342 (N_7342,N_2981,N_3750);
nand U7343 (N_7343,N_3515,N_1671);
or U7344 (N_7344,N_4208,N_3267);
nand U7345 (N_7345,N_2321,N_1856);
xnor U7346 (N_7346,N_4351,N_4622);
nand U7347 (N_7347,N_55,N_361);
and U7348 (N_7348,N_920,N_4149);
nand U7349 (N_7349,N_3696,N_1018);
or U7350 (N_7350,N_3427,N_1396);
and U7351 (N_7351,N_1357,N_2723);
nand U7352 (N_7352,N_2709,N_1384);
nand U7353 (N_7353,N_4962,N_1824);
or U7354 (N_7354,N_4521,N_2101);
nor U7355 (N_7355,N_1779,N_1668);
nand U7356 (N_7356,N_1015,N_2933);
nand U7357 (N_7357,N_3068,N_4990);
and U7358 (N_7358,N_4805,N_4241);
and U7359 (N_7359,N_1511,N_2103);
or U7360 (N_7360,N_118,N_827);
nor U7361 (N_7361,N_1364,N_2218);
nor U7362 (N_7362,N_463,N_3952);
and U7363 (N_7363,N_3915,N_929);
and U7364 (N_7364,N_278,N_372);
nor U7365 (N_7365,N_1821,N_1701);
nand U7366 (N_7366,N_4520,N_723);
nand U7367 (N_7367,N_3787,N_4428);
xor U7368 (N_7368,N_2105,N_2964);
nor U7369 (N_7369,N_492,N_38);
nor U7370 (N_7370,N_561,N_4392);
or U7371 (N_7371,N_1249,N_1520);
or U7372 (N_7372,N_4310,N_2259);
and U7373 (N_7373,N_417,N_2618);
nand U7374 (N_7374,N_4827,N_4331);
nor U7375 (N_7375,N_1181,N_2186);
or U7376 (N_7376,N_3600,N_3722);
or U7377 (N_7377,N_4735,N_2299);
nand U7378 (N_7378,N_3447,N_689);
nor U7379 (N_7379,N_2702,N_3228);
or U7380 (N_7380,N_2948,N_1096);
or U7381 (N_7381,N_3045,N_2391);
nor U7382 (N_7382,N_2987,N_3889);
xnor U7383 (N_7383,N_4533,N_1927);
nand U7384 (N_7384,N_3762,N_2498);
nand U7385 (N_7385,N_4512,N_2503);
and U7386 (N_7386,N_4311,N_4353);
or U7387 (N_7387,N_4458,N_4469);
nor U7388 (N_7388,N_3022,N_2521);
or U7389 (N_7389,N_1061,N_2884);
or U7390 (N_7390,N_4569,N_258);
nor U7391 (N_7391,N_3567,N_917);
nor U7392 (N_7392,N_1597,N_573);
or U7393 (N_7393,N_2200,N_158);
and U7394 (N_7394,N_441,N_1258);
nor U7395 (N_7395,N_3278,N_4359);
or U7396 (N_7396,N_2911,N_4598);
nand U7397 (N_7397,N_2465,N_4800);
nor U7398 (N_7398,N_3190,N_2968);
nand U7399 (N_7399,N_3264,N_1721);
and U7400 (N_7400,N_526,N_3886);
nand U7401 (N_7401,N_3414,N_2196);
and U7402 (N_7402,N_4190,N_2531);
nor U7403 (N_7403,N_4778,N_4267);
nor U7404 (N_7404,N_1309,N_824);
and U7405 (N_7405,N_2611,N_4227);
xnor U7406 (N_7406,N_53,N_2022);
nand U7407 (N_7407,N_3239,N_1616);
and U7408 (N_7408,N_4024,N_1136);
xor U7409 (N_7409,N_1218,N_1288);
xnor U7410 (N_7410,N_1658,N_873);
nor U7411 (N_7411,N_1743,N_2231);
xor U7412 (N_7412,N_1006,N_4989);
and U7413 (N_7413,N_1697,N_1033);
and U7414 (N_7414,N_1169,N_4505);
nand U7415 (N_7415,N_3605,N_4081);
and U7416 (N_7416,N_4971,N_3596);
and U7417 (N_7417,N_285,N_2423);
and U7418 (N_7418,N_4668,N_1234);
xor U7419 (N_7419,N_4658,N_2077);
nand U7420 (N_7420,N_3721,N_847);
nand U7421 (N_7421,N_2296,N_702);
nor U7422 (N_7422,N_795,N_251);
nor U7423 (N_7423,N_4421,N_3093);
or U7424 (N_7424,N_223,N_1799);
xor U7425 (N_7425,N_4148,N_4297);
nor U7426 (N_7426,N_889,N_3059);
nand U7427 (N_7427,N_841,N_2176);
or U7428 (N_7428,N_1368,N_229);
nand U7429 (N_7429,N_4861,N_2711);
nor U7430 (N_7430,N_2432,N_592);
and U7431 (N_7431,N_2803,N_760);
and U7432 (N_7432,N_4627,N_2037);
nor U7433 (N_7433,N_4390,N_1155);
nor U7434 (N_7434,N_1521,N_378);
and U7435 (N_7435,N_1860,N_2820);
nand U7436 (N_7436,N_2449,N_4396);
or U7437 (N_7437,N_4537,N_2666);
and U7438 (N_7438,N_4913,N_2168);
nand U7439 (N_7439,N_1190,N_4625);
nor U7440 (N_7440,N_445,N_2466);
nor U7441 (N_7441,N_1200,N_3457);
or U7442 (N_7442,N_3140,N_4363);
and U7443 (N_7443,N_1645,N_4270);
or U7444 (N_7444,N_4193,N_3290);
and U7445 (N_7445,N_1903,N_2486);
or U7446 (N_7446,N_4272,N_4461);
or U7447 (N_7447,N_835,N_3198);
nor U7448 (N_7448,N_151,N_4429);
or U7449 (N_7449,N_3638,N_4259);
and U7450 (N_7450,N_3300,N_2835);
or U7451 (N_7451,N_3880,N_3514);
nand U7452 (N_7452,N_332,N_369);
nand U7453 (N_7453,N_2737,N_3467);
nand U7454 (N_7454,N_1733,N_82);
nand U7455 (N_7455,N_3681,N_4144);
or U7456 (N_7456,N_3166,N_2916);
and U7457 (N_7457,N_679,N_602);
nor U7458 (N_7458,N_4229,N_826);
and U7459 (N_7459,N_1185,N_1882);
nand U7460 (N_7460,N_324,N_2706);
or U7461 (N_7461,N_1310,N_2348);
nor U7462 (N_7462,N_333,N_2228);
nor U7463 (N_7463,N_4329,N_1961);
nor U7464 (N_7464,N_2940,N_2098);
xnor U7465 (N_7465,N_3132,N_4643);
nor U7466 (N_7466,N_2986,N_2362);
nor U7467 (N_7467,N_4851,N_619);
nor U7468 (N_7468,N_3167,N_1941);
nand U7469 (N_7469,N_4875,N_3699);
or U7470 (N_7470,N_4105,N_2786);
and U7471 (N_7471,N_1713,N_3937);
nand U7472 (N_7472,N_1316,N_641);
or U7473 (N_7473,N_1953,N_654);
and U7474 (N_7474,N_1744,N_1186);
nand U7475 (N_7475,N_3577,N_1454);
nand U7476 (N_7476,N_523,N_2125);
nand U7477 (N_7477,N_1648,N_1476);
nor U7478 (N_7478,N_3341,N_2954);
or U7479 (N_7479,N_3432,N_2930);
nor U7480 (N_7480,N_3669,N_1826);
or U7481 (N_7481,N_3866,N_2550);
or U7482 (N_7482,N_4150,N_4121);
nand U7483 (N_7483,N_1412,N_3260);
nand U7484 (N_7484,N_290,N_1352);
nand U7485 (N_7485,N_3827,N_2939);
and U7486 (N_7486,N_109,N_1207);
nor U7487 (N_7487,N_3884,N_4723);
and U7488 (N_7488,N_2696,N_1997);
nor U7489 (N_7489,N_3813,N_3782);
nand U7490 (N_7490,N_1029,N_3442);
nand U7491 (N_7491,N_4147,N_3311);
and U7492 (N_7492,N_4530,N_1573);
and U7493 (N_7493,N_1607,N_3276);
or U7494 (N_7494,N_73,N_3509);
nor U7495 (N_7495,N_933,N_4909);
nand U7496 (N_7496,N_1690,N_4986);
nor U7497 (N_7497,N_2137,N_4548);
nor U7498 (N_7498,N_1126,N_910);
xor U7499 (N_7499,N_2856,N_1485);
or U7500 (N_7500,N_1077,N_1181);
nor U7501 (N_7501,N_2092,N_1943);
nand U7502 (N_7502,N_783,N_4034);
nor U7503 (N_7503,N_1086,N_2201);
xnor U7504 (N_7504,N_429,N_1010);
and U7505 (N_7505,N_4187,N_745);
nand U7506 (N_7506,N_3265,N_544);
or U7507 (N_7507,N_4476,N_1563);
nor U7508 (N_7508,N_1675,N_2940);
nor U7509 (N_7509,N_2615,N_3345);
or U7510 (N_7510,N_168,N_4772);
nand U7511 (N_7511,N_3512,N_3879);
nor U7512 (N_7512,N_2492,N_3226);
nor U7513 (N_7513,N_3110,N_714);
nand U7514 (N_7514,N_132,N_1118);
or U7515 (N_7515,N_1471,N_3217);
or U7516 (N_7516,N_3389,N_893);
nor U7517 (N_7517,N_237,N_3399);
and U7518 (N_7518,N_3760,N_4080);
nor U7519 (N_7519,N_1265,N_2472);
and U7520 (N_7520,N_2491,N_4255);
nor U7521 (N_7521,N_4294,N_3182);
nor U7522 (N_7522,N_1904,N_3816);
nor U7523 (N_7523,N_3407,N_3930);
nand U7524 (N_7524,N_2036,N_1518);
xor U7525 (N_7525,N_923,N_1822);
nand U7526 (N_7526,N_930,N_3306);
and U7527 (N_7527,N_2798,N_703);
and U7528 (N_7528,N_2968,N_1616);
nand U7529 (N_7529,N_3184,N_69);
or U7530 (N_7530,N_4396,N_4393);
or U7531 (N_7531,N_698,N_4243);
nor U7532 (N_7532,N_1095,N_749);
or U7533 (N_7533,N_431,N_4919);
nand U7534 (N_7534,N_2744,N_4140);
or U7535 (N_7535,N_655,N_3400);
and U7536 (N_7536,N_4185,N_3797);
or U7537 (N_7537,N_802,N_4005);
xnor U7538 (N_7538,N_4983,N_4133);
or U7539 (N_7539,N_1456,N_4872);
nor U7540 (N_7540,N_2881,N_1175);
nor U7541 (N_7541,N_4102,N_4200);
nand U7542 (N_7542,N_3471,N_1860);
nand U7543 (N_7543,N_4029,N_4738);
and U7544 (N_7544,N_3178,N_667);
or U7545 (N_7545,N_17,N_1179);
and U7546 (N_7546,N_2690,N_1721);
nand U7547 (N_7547,N_3984,N_4341);
and U7548 (N_7548,N_3470,N_4639);
or U7549 (N_7549,N_4577,N_301);
or U7550 (N_7550,N_2500,N_3306);
and U7551 (N_7551,N_4868,N_2793);
nand U7552 (N_7552,N_1229,N_136);
nor U7553 (N_7553,N_4643,N_2431);
and U7554 (N_7554,N_17,N_4885);
nand U7555 (N_7555,N_4648,N_2214);
nand U7556 (N_7556,N_3792,N_3119);
or U7557 (N_7557,N_3147,N_2737);
nor U7558 (N_7558,N_1989,N_1568);
or U7559 (N_7559,N_508,N_2777);
or U7560 (N_7560,N_247,N_782);
and U7561 (N_7561,N_1328,N_1289);
and U7562 (N_7562,N_2700,N_2714);
and U7563 (N_7563,N_3563,N_1531);
and U7564 (N_7564,N_2911,N_3903);
nor U7565 (N_7565,N_4502,N_4515);
and U7566 (N_7566,N_2931,N_1333);
nand U7567 (N_7567,N_221,N_4257);
and U7568 (N_7568,N_4724,N_1985);
or U7569 (N_7569,N_1774,N_2662);
nor U7570 (N_7570,N_1835,N_4572);
or U7571 (N_7571,N_3233,N_2668);
xor U7572 (N_7572,N_2414,N_3617);
or U7573 (N_7573,N_1763,N_212);
nand U7574 (N_7574,N_2613,N_1068);
nor U7575 (N_7575,N_345,N_2590);
and U7576 (N_7576,N_860,N_1160);
or U7577 (N_7577,N_1770,N_144);
and U7578 (N_7578,N_1609,N_4155);
nand U7579 (N_7579,N_600,N_136);
or U7580 (N_7580,N_1324,N_4566);
nor U7581 (N_7581,N_1058,N_3933);
or U7582 (N_7582,N_315,N_2052);
or U7583 (N_7583,N_3714,N_3140);
and U7584 (N_7584,N_1357,N_3208);
nor U7585 (N_7585,N_4546,N_3146);
or U7586 (N_7586,N_3506,N_914);
or U7587 (N_7587,N_2050,N_2504);
and U7588 (N_7588,N_834,N_4588);
or U7589 (N_7589,N_30,N_3885);
or U7590 (N_7590,N_3392,N_3825);
nand U7591 (N_7591,N_1128,N_2844);
nor U7592 (N_7592,N_2857,N_2685);
or U7593 (N_7593,N_117,N_44);
nand U7594 (N_7594,N_1809,N_1895);
nor U7595 (N_7595,N_3820,N_3574);
nor U7596 (N_7596,N_4603,N_2516);
nand U7597 (N_7597,N_1574,N_1781);
nor U7598 (N_7598,N_108,N_891);
or U7599 (N_7599,N_2051,N_3733);
and U7600 (N_7600,N_973,N_209);
nor U7601 (N_7601,N_1088,N_2006);
xor U7602 (N_7602,N_2457,N_4870);
nand U7603 (N_7603,N_4617,N_3380);
nor U7604 (N_7604,N_3388,N_4700);
and U7605 (N_7605,N_4520,N_4312);
nor U7606 (N_7606,N_2076,N_402);
nor U7607 (N_7607,N_4206,N_2618);
nor U7608 (N_7608,N_220,N_819);
and U7609 (N_7609,N_4644,N_3311);
xor U7610 (N_7610,N_1679,N_1803);
nor U7611 (N_7611,N_2448,N_3187);
xnor U7612 (N_7612,N_4417,N_75);
or U7613 (N_7613,N_4164,N_2548);
nor U7614 (N_7614,N_3406,N_4535);
nand U7615 (N_7615,N_3940,N_4418);
and U7616 (N_7616,N_2967,N_1254);
nand U7617 (N_7617,N_1848,N_2279);
nor U7618 (N_7618,N_2705,N_2587);
nor U7619 (N_7619,N_3313,N_1452);
nand U7620 (N_7620,N_362,N_1812);
nand U7621 (N_7621,N_575,N_3372);
nand U7622 (N_7622,N_4235,N_4082);
nand U7623 (N_7623,N_4155,N_1558);
or U7624 (N_7624,N_2447,N_342);
nor U7625 (N_7625,N_3070,N_554);
nor U7626 (N_7626,N_3318,N_4095);
nor U7627 (N_7627,N_2013,N_3054);
or U7628 (N_7628,N_2509,N_4080);
nor U7629 (N_7629,N_1216,N_3305);
nand U7630 (N_7630,N_2966,N_3057);
or U7631 (N_7631,N_1613,N_4362);
and U7632 (N_7632,N_2084,N_2088);
nand U7633 (N_7633,N_3296,N_1614);
or U7634 (N_7634,N_3153,N_4878);
xnor U7635 (N_7635,N_854,N_2942);
nand U7636 (N_7636,N_4902,N_2426);
and U7637 (N_7637,N_1066,N_4513);
xor U7638 (N_7638,N_4909,N_1295);
nand U7639 (N_7639,N_4146,N_1405);
nand U7640 (N_7640,N_134,N_921);
and U7641 (N_7641,N_1913,N_4628);
or U7642 (N_7642,N_4394,N_3332);
and U7643 (N_7643,N_3084,N_1293);
or U7644 (N_7644,N_2225,N_1706);
or U7645 (N_7645,N_679,N_1863);
or U7646 (N_7646,N_3769,N_3273);
nand U7647 (N_7647,N_2141,N_1807);
or U7648 (N_7648,N_4082,N_435);
nand U7649 (N_7649,N_2997,N_3258);
or U7650 (N_7650,N_2925,N_1179);
nand U7651 (N_7651,N_32,N_3905);
and U7652 (N_7652,N_4584,N_4776);
nand U7653 (N_7653,N_18,N_4213);
nand U7654 (N_7654,N_1846,N_2116);
or U7655 (N_7655,N_1780,N_1691);
and U7656 (N_7656,N_618,N_2672);
xor U7657 (N_7657,N_2741,N_1861);
nor U7658 (N_7658,N_909,N_1147);
nor U7659 (N_7659,N_2993,N_407);
or U7660 (N_7660,N_2730,N_4432);
nor U7661 (N_7661,N_1392,N_3967);
nor U7662 (N_7662,N_4358,N_1046);
or U7663 (N_7663,N_3713,N_3082);
and U7664 (N_7664,N_4859,N_2292);
nor U7665 (N_7665,N_1032,N_3091);
or U7666 (N_7666,N_2584,N_1544);
xnor U7667 (N_7667,N_204,N_3959);
or U7668 (N_7668,N_766,N_4396);
nand U7669 (N_7669,N_2004,N_3856);
or U7670 (N_7670,N_3884,N_1593);
xor U7671 (N_7671,N_2208,N_2282);
or U7672 (N_7672,N_4984,N_3906);
nand U7673 (N_7673,N_4778,N_1790);
and U7674 (N_7674,N_2875,N_3763);
xnor U7675 (N_7675,N_1714,N_84);
and U7676 (N_7676,N_1956,N_268);
nor U7677 (N_7677,N_4071,N_2407);
nand U7678 (N_7678,N_2423,N_4724);
and U7679 (N_7679,N_1284,N_1225);
nand U7680 (N_7680,N_1567,N_1109);
or U7681 (N_7681,N_681,N_2213);
or U7682 (N_7682,N_2875,N_1643);
or U7683 (N_7683,N_647,N_1459);
nand U7684 (N_7684,N_2093,N_1376);
and U7685 (N_7685,N_2690,N_2512);
or U7686 (N_7686,N_892,N_460);
and U7687 (N_7687,N_1872,N_995);
and U7688 (N_7688,N_772,N_3301);
and U7689 (N_7689,N_4387,N_4564);
and U7690 (N_7690,N_588,N_2783);
or U7691 (N_7691,N_3171,N_844);
or U7692 (N_7692,N_2195,N_2788);
xnor U7693 (N_7693,N_3695,N_4273);
and U7694 (N_7694,N_1578,N_1759);
and U7695 (N_7695,N_1582,N_3121);
and U7696 (N_7696,N_1512,N_2085);
or U7697 (N_7697,N_4531,N_478);
or U7698 (N_7698,N_2141,N_2827);
nor U7699 (N_7699,N_2268,N_85);
and U7700 (N_7700,N_2516,N_1139);
and U7701 (N_7701,N_118,N_2566);
nor U7702 (N_7702,N_2460,N_3327);
nor U7703 (N_7703,N_2584,N_3375);
and U7704 (N_7704,N_2893,N_2342);
xnor U7705 (N_7705,N_1789,N_1211);
nand U7706 (N_7706,N_1272,N_1353);
or U7707 (N_7707,N_3404,N_1856);
or U7708 (N_7708,N_3050,N_1441);
or U7709 (N_7709,N_3008,N_4878);
nor U7710 (N_7710,N_4195,N_4003);
nand U7711 (N_7711,N_1785,N_2841);
nand U7712 (N_7712,N_2192,N_3303);
nor U7713 (N_7713,N_3411,N_2730);
and U7714 (N_7714,N_1363,N_4711);
nand U7715 (N_7715,N_3251,N_3240);
or U7716 (N_7716,N_4991,N_4655);
or U7717 (N_7717,N_4994,N_3984);
nor U7718 (N_7718,N_4548,N_3047);
nor U7719 (N_7719,N_982,N_3500);
xor U7720 (N_7720,N_4645,N_860);
nand U7721 (N_7721,N_1189,N_3315);
nor U7722 (N_7722,N_2059,N_271);
xnor U7723 (N_7723,N_436,N_484);
and U7724 (N_7724,N_3604,N_1722);
nand U7725 (N_7725,N_811,N_3102);
and U7726 (N_7726,N_996,N_4378);
nor U7727 (N_7727,N_641,N_4210);
nor U7728 (N_7728,N_4790,N_343);
or U7729 (N_7729,N_3011,N_4242);
or U7730 (N_7730,N_1093,N_3152);
nand U7731 (N_7731,N_4431,N_3120);
nor U7732 (N_7732,N_263,N_869);
and U7733 (N_7733,N_816,N_2950);
or U7734 (N_7734,N_1848,N_1703);
or U7735 (N_7735,N_357,N_1660);
and U7736 (N_7736,N_2993,N_4062);
nand U7737 (N_7737,N_1542,N_1269);
nor U7738 (N_7738,N_3335,N_4852);
nor U7739 (N_7739,N_1162,N_1901);
and U7740 (N_7740,N_3591,N_18);
nor U7741 (N_7741,N_4514,N_1158);
and U7742 (N_7742,N_1563,N_647);
nor U7743 (N_7743,N_1966,N_2293);
nand U7744 (N_7744,N_1684,N_3968);
nand U7745 (N_7745,N_517,N_4447);
or U7746 (N_7746,N_4912,N_4252);
or U7747 (N_7747,N_1590,N_2830);
nand U7748 (N_7748,N_3578,N_496);
and U7749 (N_7749,N_4122,N_1813);
nand U7750 (N_7750,N_4161,N_2473);
or U7751 (N_7751,N_3597,N_4421);
nor U7752 (N_7752,N_4555,N_4191);
and U7753 (N_7753,N_108,N_4492);
or U7754 (N_7754,N_2371,N_2269);
xor U7755 (N_7755,N_2967,N_3351);
nand U7756 (N_7756,N_861,N_3993);
or U7757 (N_7757,N_4356,N_4847);
nor U7758 (N_7758,N_608,N_1106);
or U7759 (N_7759,N_4117,N_4311);
and U7760 (N_7760,N_4965,N_4407);
nor U7761 (N_7761,N_81,N_3345);
nor U7762 (N_7762,N_2933,N_107);
nor U7763 (N_7763,N_2182,N_4683);
and U7764 (N_7764,N_347,N_1029);
or U7765 (N_7765,N_4340,N_2637);
nand U7766 (N_7766,N_1732,N_2831);
nor U7767 (N_7767,N_4033,N_4986);
and U7768 (N_7768,N_2260,N_1250);
or U7769 (N_7769,N_2653,N_3495);
or U7770 (N_7770,N_1311,N_1372);
or U7771 (N_7771,N_740,N_648);
nand U7772 (N_7772,N_3094,N_383);
and U7773 (N_7773,N_3915,N_4710);
nand U7774 (N_7774,N_3602,N_2528);
and U7775 (N_7775,N_4140,N_2357);
or U7776 (N_7776,N_4179,N_1336);
nor U7777 (N_7777,N_1484,N_3472);
nor U7778 (N_7778,N_3242,N_1255);
or U7779 (N_7779,N_1336,N_3488);
xnor U7780 (N_7780,N_3842,N_3266);
nor U7781 (N_7781,N_3086,N_3133);
nor U7782 (N_7782,N_1952,N_761);
and U7783 (N_7783,N_1477,N_488);
and U7784 (N_7784,N_614,N_481);
and U7785 (N_7785,N_2680,N_571);
and U7786 (N_7786,N_1557,N_899);
or U7787 (N_7787,N_239,N_402);
and U7788 (N_7788,N_3779,N_3055);
or U7789 (N_7789,N_3161,N_1953);
nand U7790 (N_7790,N_2552,N_1924);
nand U7791 (N_7791,N_4057,N_2117);
nand U7792 (N_7792,N_3004,N_3496);
and U7793 (N_7793,N_1159,N_1998);
and U7794 (N_7794,N_4747,N_4822);
xor U7795 (N_7795,N_936,N_842);
or U7796 (N_7796,N_2160,N_1778);
nor U7797 (N_7797,N_3616,N_700);
and U7798 (N_7798,N_982,N_2494);
nor U7799 (N_7799,N_2542,N_3313);
xnor U7800 (N_7800,N_3482,N_469);
or U7801 (N_7801,N_2403,N_4156);
nand U7802 (N_7802,N_4851,N_1076);
nor U7803 (N_7803,N_652,N_1287);
nor U7804 (N_7804,N_4673,N_4985);
nor U7805 (N_7805,N_3705,N_2368);
and U7806 (N_7806,N_3096,N_1296);
or U7807 (N_7807,N_1304,N_1747);
xnor U7808 (N_7808,N_4169,N_3392);
nand U7809 (N_7809,N_2367,N_2138);
nand U7810 (N_7810,N_1650,N_3624);
nand U7811 (N_7811,N_3912,N_3785);
and U7812 (N_7812,N_4571,N_3866);
nor U7813 (N_7813,N_3440,N_4540);
or U7814 (N_7814,N_4827,N_3383);
nor U7815 (N_7815,N_3234,N_3944);
and U7816 (N_7816,N_2734,N_4660);
nor U7817 (N_7817,N_1241,N_183);
and U7818 (N_7818,N_4936,N_4342);
and U7819 (N_7819,N_4866,N_2779);
nand U7820 (N_7820,N_1001,N_382);
nand U7821 (N_7821,N_1363,N_4959);
and U7822 (N_7822,N_2262,N_4807);
or U7823 (N_7823,N_3619,N_3978);
nor U7824 (N_7824,N_1631,N_4076);
or U7825 (N_7825,N_3697,N_758);
and U7826 (N_7826,N_4549,N_1379);
nor U7827 (N_7827,N_645,N_4911);
nor U7828 (N_7828,N_3213,N_1795);
nand U7829 (N_7829,N_2746,N_4456);
nor U7830 (N_7830,N_926,N_2591);
or U7831 (N_7831,N_1217,N_2177);
and U7832 (N_7832,N_4560,N_595);
nand U7833 (N_7833,N_427,N_1861);
or U7834 (N_7834,N_1191,N_2254);
nor U7835 (N_7835,N_2950,N_3503);
nor U7836 (N_7836,N_3842,N_4970);
or U7837 (N_7837,N_2215,N_2881);
nor U7838 (N_7838,N_3991,N_4685);
and U7839 (N_7839,N_3229,N_563);
xor U7840 (N_7840,N_1278,N_851);
xor U7841 (N_7841,N_4239,N_4326);
xor U7842 (N_7842,N_2160,N_3904);
or U7843 (N_7843,N_2780,N_527);
nand U7844 (N_7844,N_2211,N_1085);
nand U7845 (N_7845,N_4942,N_4911);
or U7846 (N_7846,N_4006,N_11);
nor U7847 (N_7847,N_1193,N_1642);
xor U7848 (N_7848,N_901,N_2747);
nor U7849 (N_7849,N_800,N_1394);
or U7850 (N_7850,N_2866,N_662);
and U7851 (N_7851,N_1820,N_1487);
xnor U7852 (N_7852,N_3895,N_2328);
and U7853 (N_7853,N_2988,N_2624);
nor U7854 (N_7854,N_4131,N_4874);
or U7855 (N_7855,N_3791,N_3863);
nand U7856 (N_7856,N_4201,N_733);
nor U7857 (N_7857,N_2798,N_1975);
nand U7858 (N_7858,N_3940,N_3193);
or U7859 (N_7859,N_2303,N_1510);
nor U7860 (N_7860,N_4370,N_4359);
nor U7861 (N_7861,N_1599,N_3808);
nand U7862 (N_7862,N_1481,N_441);
and U7863 (N_7863,N_2760,N_1921);
or U7864 (N_7864,N_4379,N_4327);
xnor U7865 (N_7865,N_1212,N_947);
or U7866 (N_7866,N_4567,N_1354);
nor U7867 (N_7867,N_1237,N_343);
nand U7868 (N_7868,N_1510,N_4417);
or U7869 (N_7869,N_4419,N_3956);
or U7870 (N_7870,N_777,N_2323);
xor U7871 (N_7871,N_2213,N_363);
or U7872 (N_7872,N_3584,N_4881);
or U7873 (N_7873,N_1662,N_1828);
xor U7874 (N_7874,N_3671,N_3730);
and U7875 (N_7875,N_1652,N_3169);
and U7876 (N_7876,N_4893,N_239);
nor U7877 (N_7877,N_2770,N_3338);
nor U7878 (N_7878,N_1967,N_1963);
and U7879 (N_7879,N_4085,N_3160);
or U7880 (N_7880,N_3304,N_2618);
nor U7881 (N_7881,N_2078,N_92);
nor U7882 (N_7882,N_3563,N_4208);
and U7883 (N_7883,N_1046,N_3406);
or U7884 (N_7884,N_3217,N_2698);
or U7885 (N_7885,N_432,N_3513);
nand U7886 (N_7886,N_434,N_3496);
nand U7887 (N_7887,N_4537,N_3348);
and U7888 (N_7888,N_1826,N_388);
nor U7889 (N_7889,N_3506,N_3571);
or U7890 (N_7890,N_4403,N_3399);
nor U7891 (N_7891,N_4839,N_2796);
xnor U7892 (N_7892,N_840,N_4961);
nand U7893 (N_7893,N_1940,N_3874);
or U7894 (N_7894,N_4489,N_4780);
and U7895 (N_7895,N_4291,N_564);
nor U7896 (N_7896,N_1739,N_2728);
and U7897 (N_7897,N_3290,N_2353);
xnor U7898 (N_7898,N_1275,N_4055);
or U7899 (N_7899,N_3789,N_90);
or U7900 (N_7900,N_1567,N_1108);
nand U7901 (N_7901,N_1320,N_1223);
xnor U7902 (N_7902,N_944,N_1500);
xnor U7903 (N_7903,N_4831,N_2173);
or U7904 (N_7904,N_58,N_2260);
and U7905 (N_7905,N_350,N_661);
nor U7906 (N_7906,N_4815,N_222);
and U7907 (N_7907,N_4211,N_3465);
nand U7908 (N_7908,N_2717,N_612);
nor U7909 (N_7909,N_422,N_3244);
and U7910 (N_7910,N_4917,N_2187);
nor U7911 (N_7911,N_404,N_2798);
nor U7912 (N_7912,N_273,N_3221);
xnor U7913 (N_7913,N_4564,N_3337);
and U7914 (N_7914,N_2111,N_4628);
or U7915 (N_7915,N_235,N_3061);
nor U7916 (N_7916,N_3785,N_2506);
nand U7917 (N_7917,N_2029,N_769);
or U7918 (N_7918,N_4143,N_1717);
or U7919 (N_7919,N_249,N_3669);
nand U7920 (N_7920,N_4814,N_256);
or U7921 (N_7921,N_2267,N_3681);
and U7922 (N_7922,N_2709,N_1507);
and U7923 (N_7923,N_3640,N_4155);
and U7924 (N_7924,N_1552,N_727);
nor U7925 (N_7925,N_2411,N_546);
or U7926 (N_7926,N_4941,N_3329);
and U7927 (N_7927,N_4966,N_3540);
and U7928 (N_7928,N_3718,N_4917);
nor U7929 (N_7929,N_1608,N_4213);
or U7930 (N_7930,N_132,N_2337);
nand U7931 (N_7931,N_2502,N_4525);
and U7932 (N_7932,N_2745,N_2900);
nor U7933 (N_7933,N_3377,N_4211);
and U7934 (N_7934,N_2550,N_1827);
nor U7935 (N_7935,N_1210,N_2678);
or U7936 (N_7936,N_2335,N_4895);
nor U7937 (N_7937,N_381,N_928);
and U7938 (N_7938,N_2708,N_3997);
and U7939 (N_7939,N_3047,N_478);
or U7940 (N_7940,N_2963,N_2485);
and U7941 (N_7941,N_3546,N_1239);
or U7942 (N_7942,N_1796,N_4115);
and U7943 (N_7943,N_2300,N_257);
nor U7944 (N_7944,N_2715,N_4181);
and U7945 (N_7945,N_3913,N_2042);
xor U7946 (N_7946,N_3722,N_583);
xor U7947 (N_7947,N_21,N_3054);
or U7948 (N_7948,N_2749,N_1790);
nor U7949 (N_7949,N_218,N_1086);
nor U7950 (N_7950,N_4493,N_3712);
nor U7951 (N_7951,N_3959,N_4525);
nor U7952 (N_7952,N_2397,N_4608);
nor U7953 (N_7953,N_2858,N_3915);
and U7954 (N_7954,N_2383,N_1101);
and U7955 (N_7955,N_4236,N_436);
nor U7956 (N_7956,N_909,N_3587);
or U7957 (N_7957,N_3595,N_1303);
nand U7958 (N_7958,N_3186,N_463);
nand U7959 (N_7959,N_1295,N_2088);
nand U7960 (N_7960,N_726,N_3368);
nor U7961 (N_7961,N_4773,N_1201);
and U7962 (N_7962,N_115,N_2785);
nor U7963 (N_7963,N_1464,N_1671);
nor U7964 (N_7964,N_3609,N_56);
or U7965 (N_7965,N_2831,N_3997);
or U7966 (N_7966,N_2596,N_1051);
nand U7967 (N_7967,N_4206,N_2962);
nand U7968 (N_7968,N_2045,N_596);
and U7969 (N_7969,N_473,N_2460);
nand U7970 (N_7970,N_4552,N_1061);
nor U7971 (N_7971,N_2847,N_3331);
xor U7972 (N_7972,N_272,N_2387);
and U7973 (N_7973,N_2990,N_3645);
and U7974 (N_7974,N_4753,N_1029);
and U7975 (N_7975,N_3207,N_4935);
and U7976 (N_7976,N_154,N_4321);
nand U7977 (N_7977,N_2667,N_300);
nor U7978 (N_7978,N_4550,N_653);
or U7979 (N_7979,N_610,N_104);
nor U7980 (N_7980,N_2755,N_3741);
xnor U7981 (N_7981,N_4459,N_4463);
nor U7982 (N_7982,N_4352,N_889);
or U7983 (N_7983,N_3290,N_4971);
or U7984 (N_7984,N_4071,N_2912);
nand U7985 (N_7985,N_3326,N_4552);
xor U7986 (N_7986,N_1891,N_997);
nand U7987 (N_7987,N_2987,N_847);
nand U7988 (N_7988,N_3197,N_4389);
or U7989 (N_7989,N_4670,N_1375);
xnor U7990 (N_7990,N_1739,N_204);
or U7991 (N_7991,N_1428,N_3023);
nand U7992 (N_7992,N_4567,N_2808);
and U7993 (N_7993,N_3474,N_2959);
nand U7994 (N_7994,N_869,N_1254);
and U7995 (N_7995,N_4218,N_1572);
or U7996 (N_7996,N_3704,N_29);
nor U7997 (N_7997,N_781,N_2559);
and U7998 (N_7998,N_4021,N_870);
nor U7999 (N_7999,N_2831,N_3460);
or U8000 (N_8000,N_319,N_3488);
or U8001 (N_8001,N_1728,N_2362);
nand U8002 (N_8002,N_4209,N_72);
nand U8003 (N_8003,N_1043,N_4610);
nor U8004 (N_8004,N_3168,N_654);
or U8005 (N_8005,N_1919,N_1841);
or U8006 (N_8006,N_4775,N_1794);
or U8007 (N_8007,N_3540,N_1114);
nor U8008 (N_8008,N_4919,N_4055);
nand U8009 (N_8009,N_4593,N_4493);
and U8010 (N_8010,N_1648,N_4500);
xnor U8011 (N_8011,N_1278,N_785);
and U8012 (N_8012,N_972,N_4359);
and U8013 (N_8013,N_1392,N_1947);
or U8014 (N_8014,N_2289,N_820);
xor U8015 (N_8015,N_4586,N_2056);
xnor U8016 (N_8016,N_3618,N_4761);
nor U8017 (N_8017,N_2997,N_3520);
xnor U8018 (N_8018,N_218,N_2430);
nand U8019 (N_8019,N_1149,N_1492);
or U8020 (N_8020,N_586,N_2656);
xor U8021 (N_8021,N_3738,N_3082);
and U8022 (N_8022,N_3904,N_4238);
xnor U8023 (N_8023,N_46,N_4712);
nand U8024 (N_8024,N_2213,N_269);
or U8025 (N_8025,N_3963,N_882);
or U8026 (N_8026,N_2349,N_1996);
nor U8027 (N_8027,N_3647,N_2034);
or U8028 (N_8028,N_1140,N_4425);
and U8029 (N_8029,N_4625,N_1856);
nor U8030 (N_8030,N_1984,N_3200);
and U8031 (N_8031,N_1627,N_1131);
and U8032 (N_8032,N_4219,N_2728);
nor U8033 (N_8033,N_4382,N_3318);
or U8034 (N_8034,N_4823,N_3139);
nand U8035 (N_8035,N_608,N_2981);
and U8036 (N_8036,N_2360,N_243);
or U8037 (N_8037,N_2339,N_2173);
nor U8038 (N_8038,N_3372,N_4164);
or U8039 (N_8039,N_2766,N_2486);
nand U8040 (N_8040,N_79,N_3650);
nand U8041 (N_8041,N_3917,N_3425);
xor U8042 (N_8042,N_3895,N_512);
or U8043 (N_8043,N_4019,N_2297);
xor U8044 (N_8044,N_4178,N_805);
nand U8045 (N_8045,N_3403,N_2268);
xnor U8046 (N_8046,N_4326,N_2873);
and U8047 (N_8047,N_752,N_3176);
nor U8048 (N_8048,N_212,N_2711);
and U8049 (N_8049,N_720,N_168);
or U8050 (N_8050,N_2699,N_778);
nand U8051 (N_8051,N_19,N_1068);
nor U8052 (N_8052,N_2414,N_860);
or U8053 (N_8053,N_1724,N_3977);
or U8054 (N_8054,N_397,N_4315);
and U8055 (N_8055,N_921,N_568);
or U8056 (N_8056,N_665,N_3218);
xnor U8057 (N_8057,N_3098,N_4569);
nand U8058 (N_8058,N_3318,N_2787);
xnor U8059 (N_8059,N_3058,N_3273);
and U8060 (N_8060,N_4345,N_2869);
or U8061 (N_8061,N_4570,N_4856);
nor U8062 (N_8062,N_1861,N_2323);
xor U8063 (N_8063,N_3728,N_4888);
nor U8064 (N_8064,N_1500,N_1311);
nand U8065 (N_8065,N_2214,N_1615);
xor U8066 (N_8066,N_1624,N_4830);
nand U8067 (N_8067,N_145,N_1728);
and U8068 (N_8068,N_3672,N_1945);
and U8069 (N_8069,N_3407,N_2077);
nand U8070 (N_8070,N_401,N_4202);
xor U8071 (N_8071,N_2598,N_3982);
xor U8072 (N_8072,N_2184,N_674);
nor U8073 (N_8073,N_3348,N_1435);
nand U8074 (N_8074,N_480,N_4830);
and U8075 (N_8075,N_4388,N_4963);
nand U8076 (N_8076,N_4172,N_345);
nand U8077 (N_8077,N_4009,N_2538);
and U8078 (N_8078,N_1561,N_3281);
nand U8079 (N_8079,N_1602,N_499);
or U8080 (N_8080,N_1223,N_4428);
nand U8081 (N_8081,N_3320,N_2585);
nor U8082 (N_8082,N_3103,N_3688);
and U8083 (N_8083,N_2604,N_3265);
nor U8084 (N_8084,N_943,N_3712);
or U8085 (N_8085,N_4358,N_592);
and U8086 (N_8086,N_3199,N_3897);
nor U8087 (N_8087,N_1435,N_1901);
nand U8088 (N_8088,N_1898,N_363);
nor U8089 (N_8089,N_509,N_3091);
and U8090 (N_8090,N_448,N_885);
and U8091 (N_8091,N_3162,N_3436);
and U8092 (N_8092,N_3169,N_4699);
nor U8093 (N_8093,N_708,N_2861);
nor U8094 (N_8094,N_2723,N_2316);
nor U8095 (N_8095,N_2510,N_27);
nand U8096 (N_8096,N_3183,N_1730);
or U8097 (N_8097,N_1331,N_1349);
nor U8098 (N_8098,N_3761,N_4459);
or U8099 (N_8099,N_1427,N_1421);
xor U8100 (N_8100,N_4271,N_2785);
or U8101 (N_8101,N_4407,N_855);
or U8102 (N_8102,N_1410,N_1191);
nor U8103 (N_8103,N_196,N_4812);
nand U8104 (N_8104,N_2919,N_4040);
nand U8105 (N_8105,N_4505,N_2000);
and U8106 (N_8106,N_4257,N_3982);
nor U8107 (N_8107,N_3566,N_3378);
nor U8108 (N_8108,N_30,N_4921);
and U8109 (N_8109,N_3050,N_549);
nand U8110 (N_8110,N_4432,N_3006);
nand U8111 (N_8111,N_2621,N_263);
and U8112 (N_8112,N_3595,N_2198);
or U8113 (N_8113,N_3433,N_3470);
nand U8114 (N_8114,N_2517,N_4775);
nand U8115 (N_8115,N_651,N_2011);
and U8116 (N_8116,N_2982,N_2678);
nand U8117 (N_8117,N_3133,N_2335);
nor U8118 (N_8118,N_1041,N_4025);
nor U8119 (N_8119,N_245,N_3625);
xnor U8120 (N_8120,N_2450,N_1750);
nor U8121 (N_8121,N_2315,N_3795);
xor U8122 (N_8122,N_1700,N_397);
and U8123 (N_8123,N_2083,N_2526);
and U8124 (N_8124,N_3573,N_3093);
nor U8125 (N_8125,N_1700,N_104);
nor U8126 (N_8126,N_365,N_4423);
and U8127 (N_8127,N_33,N_123);
or U8128 (N_8128,N_4412,N_513);
nand U8129 (N_8129,N_4122,N_243);
or U8130 (N_8130,N_3194,N_1186);
xor U8131 (N_8131,N_4254,N_4731);
nand U8132 (N_8132,N_1475,N_3896);
xor U8133 (N_8133,N_78,N_3043);
nand U8134 (N_8134,N_2479,N_464);
nand U8135 (N_8135,N_4317,N_4480);
nand U8136 (N_8136,N_3462,N_2443);
nor U8137 (N_8137,N_4045,N_3980);
xor U8138 (N_8138,N_435,N_674);
or U8139 (N_8139,N_3066,N_4430);
nand U8140 (N_8140,N_2926,N_1922);
nand U8141 (N_8141,N_788,N_590);
and U8142 (N_8142,N_581,N_203);
and U8143 (N_8143,N_1630,N_4822);
nand U8144 (N_8144,N_294,N_370);
and U8145 (N_8145,N_3538,N_4180);
nor U8146 (N_8146,N_775,N_75);
nor U8147 (N_8147,N_56,N_2836);
nor U8148 (N_8148,N_3547,N_2841);
xnor U8149 (N_8149,N_60,N_4263);
or U8150 (N_8150,N_501,N_2702);
or U8151 (N_8151,N_1814,N_1275);
or U8152 (N_8152,N_394,N_3484);
nand U8153 (N_8153,N_104,N_2107);
nor U8154 (N_8154,N_4154,N_4259);
and U8155 (N_8155,N_914,N_606);
nand U8156 (N_8156,N_2580,N_1130);
nand U8157 (N_8157,N_1904,N_1605);
or U8158 (N_8158,N_3823,N_701);
or U8159 (N_8159,N_337,N_4851);
nand U8160 (N_8160,N_3926,N_948);
nor U8161 (N_8161,N_2722,N_4833);
and U8162 (N_8162,N_4988,N_206);
nor U8163 (N_8163,N_1783,N_2358);
nand U8164 (N_8164,N_1963,N_755);
or U8165 (N_8165,N_129,N_3027);
nor U8166 (N_8166,N_1332,N_566);
nor U8167 (N_8167,N_1971,N_3854);
and U8168 (N_8168,N_4413,N_2851);
or U8169 (N_8169,N_3154,N_1616);
nor U8170 (N_8170,N_3352,N_740);
or U8171 (N_8171,N_4335,N_1686);
xor U8172 (N_8172,N_1181,N_342);
or U8173 (N_8173,N_1102,N_3104);
and U8174 (N_8174,N_2679,N_662);
and U8175 (N_8175,N_1856,N_2760);
nand U8176 (N_8176,N_55,N_2104);
nor U8177 (N_8177,N_2475,N_2365);
or U8178 (N_8178,N_2651,N_3922);
and U8179 (N_8179,N_488,N_276);
nand U8180 (N_8180,N_2723,N_3565);
nand U8181 (N_8181,N_4889,N_359);
and U8182 (N_8182,N_2984,N_4064);
and U8183 (N_8183,N_1616,N_1332);
nor U8184 (N_8184,N_2832,N_2763);
or U8185 (N_8185,N_3623,N_4327);
and U8186 (N_8186,N_3893,N_85);
nand U8187 (N_8187,N_1592,N_4372);
nor U8188 (N_8188,N_1511,N_2544);
nor U8189 (N_8189,N_1696,N_76);
and U8190 (N_8190,N_1468,N_3081);
or U8191 (N_8191,N_2154,N_4767);
and U8192 (N_8192,N_1293,N_4295);
nor U8193 (N_8193,N_2745,N_629);
nor U8194 (N_8194,N_2016,N_976);
nor U8195 (N_8195,N_4133,N_1249);
xnor U8196 (N_8196,N_1764,N_2884);
or U8197 (N_8197,N_2446,N_1746);
xor U8198 (N_8198,N_3655,N_2849);
and U8199 (N_8199,N_2664,N_837);
nand U8200 (N_8200,N_2992,N_3681);
and U8201 (N_8201,N_4271,N_880);
or U8202 (N_8202,N_3438,N_2636);
xnor U8203 (N_8203,N_469,N_900);
nand U8204 (N_8204,N_1741,N_4056);
nor U8205 (N_8205,N_3921,N_850);
nand U8206 (N_8206,N_3793,N_437);
nand U8207 (N_8207,N_1236,N_389);
nor U8208 (N_8208,N_2655,N_532);
xor U8209 (N_8209,N_2245,N_4926);
and U8210 (N_8210,N_4472,N_724);
nor U8211 (N_8211,N_3849,N_2720);
nor U8212 (N_8212,N_3666,N_4684);
and U8213 (N_8213,N_4697,N_1611);
nand U8214 (N_8214,N_6,N_1977);
nor U8215 (N_8215,N_208,N_1410);
and U8216 (N_8216,N_4557,N_2630);
nor U8217 (N_8217,N_1403,N_3847);
nor U8218 (N_8218,N_1436,N_2932);
nand U8219 (N_8219,N_3116,N_2256);
and U8220 (N_8220,N_168,N_3754);
and U8221 (N_8221,N_4907,N_4580);
xor U8222 (N_8222,N_1740,N_4376);
nor U8223 (N_8223,N_3884,N_1643);
and U8224 (N_8224,N_541,N_3383);
nor U8225 (N_8225,N_2921,N_4546);
nand U8226 (N_8226,N_4607,N_3856);
or U8227 (N_8227,N_440,N_4606);
nor U8228 (N_8228,N_1163,N_1248);
and U8229 (N_8229,N_2603,N_3727);
and U8230 (N_8230,N_3800,N_1596);
nor U8231 (N_8231,N_3513,N_3887);
and U8232 (N_8232,N_4906,N_1246);
xor U8233 (N_8233,N_4242,N_2273);
nor U8234 (N_8234,N_2461,N_3815);
nor U8235 (N_8235,N_3217,N_2812);
and U8236 (N_8236,N_4259,N_1494);
nor U8237 (N_8237,N_2089,N_875);
nor U8238 (N_8238,N_3099,N_2496);
and U8239 (N_8239,N_3399,N_1102);
or U8240 (N_8240,N_4836,N_3866);
nand U8241 (N_8241,N_161,N_2418);
nor U8242 (N_8242,N_2746,N_2939);
and U8243 (N_8243,N_2310,N_456);
nor U8244 (N_8244,N_4381,N_1138);
nor U8245 (N_8245,N_2716,N_158);
and U8246 (N_8246,N_2991,N_371);
or U8247 (N_8247,N_3097,N_4331);
or U8248 (N_8248,N_1940,N_4205);
or U8249 (N_8249,N_1131,N_4156);
nand U8250 (N_8250,N_4231,N_2129);
nor U8251 (N_8251,N_2542,N_604);
nor U8252 (N_8252,N_1943,N_4318);
nor U8253 (N_8253,N_3196,N_331);
xor U8254 (N_8254,N_1830,N_1408);
or U8255 (N_8255,N_1899,N_2397);
nor U8256 (N_8256,N_2242,N_218);
or U8257 (N_8257,N_3716,N_1472);
or U8258 (N_8258,N_711,N_4945);
and U8259 (N_8259,N_1328,N_4014);
nor U8260 (N_8260,N_3259,N_4788);
xor U8261 (N_8261,N_4709,N_2851);
or U8262 (N_8262,N_3224,N_96);
nand U8263 (N_8263,N_4352,N_3688);
xnor U8264 (N_8264,N_3597,N_3106);
or U8265 (N_8265,N_1094,N_2046);
nand U8266 (N_8266,N_879,N_2078);
nor U8267 (N_8267,N_373,N_824);
and U8268 (N_8268,N_3551,N_2642);
nand U8269 (N_8269,N_918,N_2044);
or U8270 (N_8270,N_1432,N_1601);
nor U8271 (N_8271,N_2145,N_1729);
or U8272 (N_8272,N_4780,N_4345);
or U8273 (N_8273,N_3984,N_218);
and U8274 (N_8274,N_2824,N_314);
nand U8275 (N_8275,N_4701,N_2475);
nor U8276 (N_8276,N_2630,N_3239);
nor U8277 (N_8277,N_2852,N_994);
nand U8278 (N_8278,N_3854,N_4768);
nand U8279 (N_8279,N_4823,N_4388);
nor U8280 (N_8280,N_4101,N_2409);
nand U8281 (N_8281,N_1572,N_4626);
nand U8282 (N_8282,N_4362,N_3273);
nor U8283 (N_8283,N_4206,N_234);
and U8284 (N_8284,N_3594,N_197);
or U8285 (N_8285,N_3247,N_581);
or U8286 (N_8286,N_4472,N_4817);
nor U8287 (N_8287,N_4444,N_4898);
or U8288 (N_8288,N_2528,N_3211);
xnor U8289 (N_8289,N_4436,N_3489);
and U8290 (N_8290,N_4310,N_2886);
nand U8291 (N_8291,N_156,N_2690);
nand U8292 (N_8292,N_3301,N_2283);
nor U8293 (N_8293,N_3790,N_2966);
nand U8294 (N_8294,N_4614,N_4006);
and U8295 (N_8295,N_3089,N_3954);
nor U8296 (N_8296,N_733,N_1199);
and U8297 (N_8297,N_1730,N_4831);
and U8298 (N_8298,N_4677,N_4045);
xor U8299 (N_8299,N_4765,N_4207);
xor U8300 (N_8300,N_3345,N_429);
nor U8301 (N_8301,N_389,N_4810);
nor U8302 (N_8302,N_4217,N_4531);
xnor U8303 (N_8303,N_420,N_3376);
nor U8304 (N_8304,N_2786,N_3817);
and U8305 (N_8305,N_4459,N_2787);
nand U8306 (N_8306,N_980,N_4642);
and U8307 (N_8307,N_4055,N_974);
nand U8308 (N_8308,N_3010,N_955);
nand U8309 (N_8309,N_4681,N_4837);
or U8310 (N_8310,N_1453,N_2553);
xor U8311 (N_8311,N_848,N_899);
or U8312 (N_8312,N_3062,N_4909);
or U8313 (N_8313,N_4787,N_721);
nor U8314 (N_8314,N_3487,N_4753);
nor U8315 (N_8315,N_4597,N_2602);
nor U8316 (N_8316,N_4190,N_3364);
or U8317 (N_8317,N_4916,N_2295);
nand U8318 (N_8318,N_2338,N_2645);
nor U8319 (N_8319,N_4919,N_602);
or U8320 (N_8320,N_1333,N_2322);
nor U8321 (N_8321,N_4891,N_1334);
and U8322 (N_8322,N_3908,N_3563);
and U8323 (N_8323,N_2702,N_4183);
and U8324 (N_8324,N_3742,N_3891);
nor U8325 (N_8325,N_265,N_670);
xnor U8326 (N_8326,N_3286,N_1925);
nor U8327 (N_8327,N_152,N_1227);
nor U8328 (N_8328,N_3971,N_320);
and U8329 (N_8329,N_1778,N_2375);
and U8330 (N_8330,N_1956,N_3407);
nor U8331 (N_8331,N_381,N_1377);
nor U8332 (N_8332,N_2546,N_3724);
xnor U8333 (N_8333,N_2035,N_1278);
or U8334 (N_8334,N_4842,N_2277);
nand U8335 (N_8335,N_4724,N_4960);
or U8336 (N_8336,N_117,N_3197);
nor U8337 (N_8337,N_438,N_3507);
and U8338 (N_8338,N_1755,N_117);
or U8339 (N_8339,N_902,N_2929);
nand U8340 (N_8340,N_330,N_1745);
nand U8341 (N_8341,N_2691,N_4439);
or U8342 (N_8342,N_3548,N_2735);
or U8343 (N_8343,N_2160,N_2039);
nand U8344 (N_8344,N_2434,N_171);
xor U8345 (N_8345,N_259,N_2982);
nand U8346 (N_8346,N_646,N_3774);
and U8347 (N_8347,N_3133,N_2093);
and U8348 (N_8348,N_3281,N_614);
and U8349 (N_8349,N_3229,N_948);
or U8350 (N_8350,N_2167,N_1381);
nand U8351 (N_8351,N_3091,N_451);
and U8352 (N_8352,N_2013,N_1984);
and U8353 (N_8353,N_1172,N_4807);
and U8354 (N_8354,N_1035,N_2104);
and U8355 (N_8355,N_695,N_3705);
nand U8356 (N_8356,N_4340,N_3885);
nand U8357 (N_8357,N_2683,N_1192);
and U8358 (N_8358,N_2950,N_1765);
and U8359 (N_8359,N_869,N_4695);
xor U8360 (N_8360,N_2671,N_2582);
and U8361 (N_8361,N_3141,N_3815);
nor U8362 (N_8362,N_4309,N_3658);
and U8363 (N_8363,N_4534,N_4446);
or U8364 (N_8364,N_543,N_2384);
nor U8365 (N_8365,N_2416,N_571);
nor U8366 (N_8366,N_3567,N_2340);
and U8367 (N_8367,N_506,N_1106);
xor U8368 (N_8368,N_3226,N_2137);
nor U8369 (N_8369,N_2162,N_3797);
xor U8370 (N_8370,N_1236,N_3347);
nand U8371 (N_8371,N_1743,N_4998);
or U8372 (N_8372,N_2758,N_3166);
nand U8373 (N_8373,N_1484,N_1253);
nand U8374 (N_8374,N_4370,N_1446);
nand U8375 (N_8375,N_673,N_4759);
nand U8376 (N_8376,N_4511,N_65);
or U8377 (N_8377,N_450,N_2605);
xor U8378 (N_8378,N_110,N_3270);
and U8379 (N_8379,N_4573,N_3966);
nand U8380 (N_8380,N_2677,N_2050);
nor U8381 (N_8381,N_743,N_4730);
or U8382 (N_8382,N_693,N_830);
or U8383 (N_8383,N_2379,N_1167);
nand U8384 (N_8384,N_2450,N_3284);
nor U8385 (N_8385,N_1996,N_1373);
nand U8386 (N_8386,N_4022,N_2423);
xnor U8387 (N_8387,N_2468,N_2058);
nor U8388 (N_8388,N_2461,N_188);
xor U8389 (N_8389,N_2707,N_396);
and U8390 (N_8390,N_4074,N_2302);
nor U8391 (N_8391,N_730,N_3767);
nand U8392 (N_8392,N_1271,N_824);
nor U8393 (N_8393,N_3004,N_3088);
nand U8394 (N_8394,N_3060,N_957);
and U8395 (N_8395,N_4600,N_3544);
or U8396 (N_8396,N_1527,N_1554);
nand U8397 (N_8397,N_1103,N_4945);
or U8398 (N_8398,N_2770,N_617);
and U8399 (N_8399,N_0,N_3902);
or U8400 (N_8400,N_4960,N_2964);
nor U8401 (N_8401,N_2626,N_298);
nand U8402 (N_8402,N_3952,N_52);
or U8403 (N_8403,N_2464,N_217);
nand U8404 (N_8404,N_196,N_1060);
and U8405 (N_8405,N_2445,N_3916);
and U8406 (N_8406,N_2349,N_1173);
nand U8407 (N_8407,N_3054,N_2352);
xnor U8408 (N_8408,N_763,N_116);
xor U8409 (N_8409,N_1995,N_2821);
or U8410 (N_8410,N_4923,N_922);
nor U8411 (N_8411,N_922,N_209);
nand U8412 (N_8412,N_4501,N_2464);
nand U8413 (N_8413,N_3078,N_1103);
xor U8414 (N_8414,N_4783,N_2824);
nor U8415 (N_8415,N_927,N_3995);
nand U8416 (N_8416,N_1049,N_3490);
or U8417 (N_8417,N_1176,N_2429);
and U8418 (N_8418,N_1283,N_2797);
nand U8419 (N_8419,N_3423,N_198);
xnor U8420 (N_8420,N_2637,N_2045);
nand U8421 (N_8421,N_2487,N_2194);
or U8422 (N_8422,N_4100,N_3649);
nor U8423 (N_8423,N_3496,N_4551);
xor U8424 (N_8424,N_209,N_3623);
nand U8425 (N_8425,N_3343,N_2701);
or U8426 (N_8426,N_1099,N_731);
or U8427 (N_8427,N_733,N_3403);
nand U8428 (N_8428,N_1448,N_3415);
and U8429 (N_8429,N_3237,N_4272);
xor U8430 (N_8430,N_2682,N_1808);
and U8431 (N_8431,N_2991,N_1430);
or U8432 (N_8432,N_735,N_1995);
nand U8433 (N_8433,N_829,N_241);
nor U8434 (N_8434,N_4693,N_4995);
and U8435 (N_8435,N_4218,N_2931);
nand U8436 (N_8436,N_474,N_1348);
nor U8437 (N_8437,N_4988,N_3251);
xor U8438 (N_8438,N_1779,N_3762);
nor U8439 (N_8439,N_2779,N_1520);
nand U8440 (N_8440,N_1138,N_3850);
nand U8441 (N_8441,N_3265,N_4341);
or U8442 (N_8442,N_798,N_3015);
nor U8443 (N_8443,N_2488,N_2513);
nor U8444 (N_8444,N_3427,N_4898);
xnor U8445 (N_8445,N_3336,N_879);
or U8446 (N_8446,N_1420,N_4160);
xor U8447 (N_8447,N_3198,N_2519);
and U8448 (N_8448,N_2939,N_875);
and U8449 (N_8449,N_337,N_4427);
nand U8450 (N_8450,N_1727,N_269);
nand U8451 (N_8451,N_37,N_4854);
or U8452 (N_8452,N_4258,N_4838);
nor U8453 (N_8453,N_3459,N_560);
nand U8454 (N_8454,N_3186,N_696);
nand U8455 (N_8455,N_2524,N_1382);
or U8456 (N_8456,N_275,N_3222);
and U8457 (N_8457,N_1331,N_354);
xor U8458 (N_8458,N_4796,N_1591);
nand U8459 (N_8459,N_4725,N_2972);
nand U8460 (N_8460,N_1080,N_3117);
nor U8461 (N_8461,N_4497,N_4830);
or U8462 (N_8462,N_4365,N_1684);
nand U8463 (N_8463,N_2427,N_3491);
nand U8464 (N_8464,N_1737,N_4947);
or U8465 (N_8465,N_4550,N_460);
or U8466 (N_8466,N_316,N_1084);
and U8467 (N_8467,N_3910,N_2991);
nand U8468 (N_8468,N_4899,N_3882);
or U8469 (N_8469,N_1983,N_1422);
and U8470 (N_8470,N_2961,N_2826);
or U8471 (N_8471,N_354,N_621);
and U8472 (N_8472,N_4959,N_1398);
or U8473 (N_8473,N_3505,N_2825);
nor U8474 (N_8474,N_3984,N_1177);
and U8475 (N_8475,N_1727,N_4470);
xor U8476 (N_8476,N_3898,N_4905);
nor U8477 (N_8477,N_2251,N_1330);
nand U8478 (N_8478,N_2762,N_4885);
nand U8479 (N_8479,N_2805,N_3926);
xnor U8480 (N_8480,N_4803,N_3317);
or U8481 (N_8481,N_4776,N_478);
nand U8482 (N_8482,N_1140,N_3147);
nor U8483 (N_8483,N_2084,N_2959);
or U8484 (N_8484,N_2390,N_3404);
or U8485 (N_8485,N_3222,N_4764);
and U8486 (N_8486,N_95,N_1340);
nor U8487 (N_8487,N_1054,N_4123);
or U8488 (N_8488,N_3250,N_2793);
nand U8489 (N_8489,N_351,N_540);
nor U8490 (N_8490,N_1203,N_312);
xnor U8491 (N_8491,N_1800,N_4352);
or U8492 (N_8492,N_2900,N_4850);
nand U8493 (N_8493,N_1570,N_759);
and U8494 (N_8494,N_3445,N_2890);
nand U8495 (N_8495,N_1795,N_2746);
nor U8496 (N_8496,N_1664,N_2452);
and U8497 (N_8497,N_4203,N_2317);
or U8498 (N_8498,N_4876,N_2427);
and U8499 (N_8499,N_2335,N_822);
nand U8500 (N_8500,N_3683,N_1267);
or U8501 (N_8501,N_3936,N_610);
and U8502 (N_8502,N_4275,N_205);
and U8503 (N_8503,N_4661,N_2263);
and U8504 (N_8504,N_2812,N_4175);
nor U8505 (N_8505,N_1710,N_4726);
nand U8506 (N_8506,N_2034,N_2391);
or U8507 (N_8507,N_996,N_4894);
nand U8508 (N_8508,N_1636,N_4616);
nor U8509 (N_8509,N_1650,N_4902);
or U8510 (N_8510,N_4913,N_992);
or U8511 (N_8511,N_4844,N_4453);
nor U8512 (N_8512,N_4137,N_4743);
nor U8513 (N_8513,N_4651,N_3972);
and U8514 (N_8514,N_1444,N_2897);
nand U8515 (N_8515,N_3264,N_559);
nand U8516 (N_8516,N_591,N_379);
nor U8517 (N_8517,N_404,N_1252);
and U8518 (N_8518,N_3882,N_3948);
and U8519 (N_8519,N_3088,N_3955);
and U8520 (N_8520,N_802,N_1504);
or U8521 (N_8521,N_3820,N_1001);
xor U8522 (N_8522,N_4328,N_3089);
or U8523 (N_8523,N_1586,N_2473);
or U8524 (N_8524,N_2640,N_2705);
and U8525 (N_8525,N_3215,N_3490);
and U8526 (N_8526,N_2457,N_4324);
xor U8527 (N_8527,N_4929,N_1077);
nand U8528 (N_8528,N_1506,N_1929);
nand U8529 (N_8529,N_1486,N_4902);
and U8530 (N_8530,N_4284,N_1345);
nand U8531 (N_8531,N_1656,N_2156);
xor U8532 (N_8532,N_622,N_1185);
nor U8533 (N_8533,N_3598,N_4741);
nor U8534 (N_8534,N_3991,N_141);
nand U8535 (N_8535,N_4848,N_1666);
and U8536 (N_8536,N_2545,N_4722);
nand U8537 (N_8537,N_1097,N_1681);
and U8538 (N_8538,N_2858,N_2042);
and U8539 (N_8539,N_3282,N_4533);
or U8540 (N_8540,N_3581,N_874);
and U8541 (N_8541,N_3164,N_4105);
nor U8542 (N_8542,N_4015,N_1094);
xor U8543 (N_8543,N_4164,N_3522);
nand U8544 (N_8544,N_3168,N_2073);
nor U8545 (N_8545,N_203,N_4863);
xor U8546 (N_8546,N_4565,N_217);
xor U8547 (N_8547,N_32,N_669);
or U8548 (N_8548,N_1125,N_4035);
nor U8549 (N_8549,N_1440,N_1719);
nand U8550 (N_8550,N_1153,N_3998);
nor U8551 (N_8551,N_1412,N_3369);
nor U8552 (N_8552,N_3213,N_79);
or U8553 (N_8553,N_4133,N_2986);
and U8554 (N_8554,N_3923,N_3306);
nand U8555 (N_8555,N_2351,N_4485);
nand U8556 (N_8556,N_1779,N_318);
and U8557 (N_8557,N_4206,N_989);
or U8558 (N_8558,N_3826,N_4817);
nand U8559 (N_8559,N_3480,N_634);
nor U8560 (N_8560,N_2167,N_3451);
xnor U8561 (N_8561,N_1348,N_2125);
nor U8562 (N_8562,N_1872,N_71);
or U8563 (N_8563,N_4254,N_1116);
or U8564 (N_8564,N_3007,N_1401);
nor U8565 (N_8565,N_4496,N_3766);
and U8566 (N_8566,N_4312,N_2526);
and U8567 (N_8567,N_3857,N_1387);
xnor U8568 (N_8568,N_2354,N_2596);
or U8569 (N_8569,N_4899,N_129);
nand U8570 (N_8570,N_1749,N_3748);
xnor U8571 (N_8571,N_4889,N_4156);
or U8572 (N_8572,N_2325,N_2689);
xor U8573 (N_8573,N_2974,N_4476);
and U8574 (N_8574,N_2500,N_3488);
xor U8575 (N_8575,N_1348,N_3064);
nand U8576 (N_8576,N_627,N_769);
nor U8577 (N_8577,N_11,N_3920);
or U8578 (N_8578,N_1493,N_2777);
nand U8579 (N_8579,N_2212,N_4504);
nor U8580 (N_8580,N_4845,N_3266);
and U8581 (N_8581,N_3407,N_986);
or U8582 (N_8582,N_240,N_820);
or U8583 (N_8583,N_1965,N_2811);
nor U8584 (N_8584,N_4050,N_4822);
and U8585 (N_8585,N_958,N_211);
or U8586 (N_8586,N_4474,N_805);
nor U8587 (N_8587,N_1385,N_1541);
nand U8588 (N_8588,N_1181,N_3092);
nand U8589 (N_8589,N_2318,N_2490);
nor U8590 (N_8590,N_4768,N_2063);
nor U8591 (N_8591,N_921,N_4299);
xnor U8592 (N_8592,N_152,N_3490);
xnor U8593 (N_8593,N_2342,N_26);
xnor U8594 (N_8594,N_2909,N_4382);
nor U8595 (N_8595,N_1219,N_2625);
nand U8596 (N_8596,N_1454,N_3918);
or U8597 (N_8597,N_470,N_1635);
and U8598 (N_8598,N_1860,N_68);
and U8599 (N_8599,N_4428,N_71);
nand U8600 (N_8600,N_2337,N_2252);
or U8601 (N_8601,N_88,N_405);
and U8602 (N_8602,N_1081,N_671);
and U8603 (N_8603,N_2170,N_2782);
or U8604 (N_8604,N_4944,N_720);
nand U8605 (N_8605,N_282,N_4391);
nand U8606 (N_8606,N_3922,N_312);
nand U8607 (N_8607,N_1272,N_3428);
nor U8608 (N_8608,N_1604,N_4263);
or U8609 (N_8609,N_2449,N_4519);
nand U8610 (N_8610,N_705,N_1781);
and U8611 (N_8611,N_2283,N_217);
and U8612 (N_8612,N_4121,N_714);
or U8613 (N_8613,N_1807,N_248);
nor U8614 (N_8614,N_2712,N_4302);
and U8615 (N_8615,N_2248,N_3333);
nand U8616 (N_8616,N_3900,N_3348);
xor U8617 (N_8617,N_4882,N_1563);
nor U8618 (N_8618,N_4260,N_4123);
nor U8619 (N_8619,N_4108,N_534);
nor U8620 (N_8620,N_672,N_724);
and U8621 (N_8621,N_715,N_974);
nor U8622 (N_8622,N_2513,N_4143);
nand U8623 (N_8623,N_2256,N_1196);
xor U8624 (N_8624,N_1336,N_3683);
or U8625 (N_8625,N_3276,N_2087);
and U8626 (N_8626,N_4316,N_4593);
or U8627 (N_8627,N_2597,N_942);
xnor U8628 (N_8628,N_3169,N_1270);
xnor U8629 (N_8629,N_4266,N_4800);
and U8630 (N_8630,N_2788,N_1716);
and U8631 (N_8631,N_2725,N_595);
or U8632 (N_8632,N_1193,N_1013);
xor U8633 (N_8633,N_2904,N_2598);
and U8634 (N_8634,N_4974,N_3922);
nor U8635 (N_8635,N_1341,N_3686);
or U8636 (N_8636,N_885,N_663);
nor U8637 (N_8637,N_2307,N_2096);
or U8638 (N_8638,N_1212,N_3073);
and U8639 (N_8639,N_2350,N_2702);
nand U8640 (N_8640,N_1844,N_1303);
or U8641 (N_8641,N_2346,N_251);
nor U8642 (N_8642,N_3842,N_2702);
nor U8643 (N_8643,N_2018,N_1477);
nand U8644 (N_8644,N_4131,N_4393);
nor U8645 (N_8645,N_2768,N_2112);
and U8646 (N_8646,N_4329,N_2568);
nand U8647 (N_8647,N_1671,N_4203);
or U8648 (N_8648,N_2931,N_4282);
xnor U8649 (N_8649,N_2400,N_1344);
xnor U8650 (N_8650,N_202,N_2228);
nand U8651 (N_8651,N_4742,N_3212);
or U8652 (N_8652,N_3437,N_4864);
and U8653 (N_8653,N_510,N_768);
xnor U8654 (N_8654,N_4987,N_3096);
nor U8655 (N_8655,N_3920,N_803);
or U8656 (N_8656,N_3394,N_3953);
and U8657 (N_8657,N_4076,N_36);
or U8658 (N_8658,N_4636,N_832);
xnor U8659 (N_8659,N_162,N_2251);
or U8660 (N_8660,N_301,N_3494);
nor U8661 (N_8661,N_2359,N_2463);
nor U8662 (N_8662,N_1631,N_3287);
or U8663 (N_8663,N_4864,N_1960);
and U8664 (N_8664,N_3391,N_943);
or U8665 (N_8665,N_1856,N_1284);
nor U8666 (N_8666,N_570,N_1683);
nor U8667 (N_8667,N_1687,N_3339);
or U8668 (N_8668,N_4927,N_1269);
xnor U8669 (N_8669,N_1986,N_4427);
nand U8670 (N_8670,N_1984,N_903);
and U8671 (N_8671,N_818,N_1522);
or U8672 (N_8672,N_4342,N_1500);
xnor U8673 (N_8673,N_3195,N_3757);
xnor U8674 (N_8674,N_551,N_2656);
and U8675 (N_8675,N_399,N_4843);
and U8676 (N_8676,N_1068,N_1940);
or U8677 (N_8677,N_1192,N_2394);
or U8678 (N_8678,N_3834,N_3079);
nand U8679 (N_8679,N_2687,N_3600);
nand U8680 (N_8680,N_3264,N_3780);
and U8681 (N_8681,N_255,N_409);
and U8682 (N_8682,N_3314,N_1120);
nor U8683 (N_8683,N_32,N_1964);
or U8684 (N_8684,N_590,N_1076);
nor U8685 (N_8685,N_1110,N_4168);
or U8686 (N_8686,N_4809,N_1550);
nand U8687 (N_8687,N_4022,N_2875);
nand U8688 (N_8688,N_1115,N_4155);
or U8689 (N_8689,N_828,N_510);
nand U8690 (N_8690,N_2599,N_1997);
nor U8691 (N_8691,N_3598,N_2822);
xnor U8692 (N_8692,N_2351,N_3530);
and U8693 (N_8693,N_841,N_70);
xor U8694 (N_8694,N_1700,N_1280);
and U8695 (N_8695,N_1996,N_1650);
nor U8696 (N_8696,N_1650,N_2609);
and U8697 (N_8697,N_342,N_3935);
and U8698 (N_8698,N_2695,N_1314);
nor U8699 (N_8699,N_528,N_3402);
nor U8700 (N_8700,N_9,N_2276);
xnor U8701 (N_8701,N_1115,N_470);
and U8702 (N_8702,N_478,N_2486);
and U8703 (N_8703,N_4870,N_4869);
or U8704 (N_8704,N_4084,N_3052);
or U8705 (N_8705,N_4802,N_4690);
xnor U8706 (N_8706,N_4305,N_3330);
and U8707 (N_8707,N_2369,N_3032);
nand U8708 (N_8708,N_3536,N_1489);
nor U8709 (N_8709,N_3565,N_3974);
nor U8710 (N_8710,N_3754,N_1035);
nand U8711 (N_8711,N_3382,N_1304);
nand U8712 (N_8712,N_1060,N_1696);
nand U8713 (N_8713,N_1803,N_451);
or U8714 (N_8714,N_3348,N_2798);
and U8715 (N_8715,N_2480,N_1642);
nand U8716 (N_8716,N_2196,N_3757);
xor U8717 (N_8717,N_940,N_3450);
nand U8718 (N_8718,N_1435,N_3607);
nor U8719 (N_8719,N_2224,N_3357);
xnor U8720 (N_8720,N_1342,N_3361);
nand U8721 (N_8721,N_1458,N_4973);
and U8722 (N_8722,N_1394,N_129);
and U8723 (N_8723,N_3772,N_4625);
and U8724 (N_8724,N_4311,N_1813);
nand U8725 (N_8725,N_465,N_2450);
and U8726 (N_8726,N_4708,N_2111);
nand U8727 (N_8727,N_2624,N_4601);
or U8728 (N_8728,N_3903,N_794);
nor U8729 (N_8729,N_4559,N_744);
and U8730 (N_8730,N_1454,N_544);
or U8731 (N_8731,N_2698,N_2680);
nand U8732 (N_8732,N_2317,N_3502);
and U8733 (N_8733,N_68,N_862);
nand U8734 (N_8734,N_4269,N_1201);
and U8735 (N_8735,N_4893,N_1027);
or U8736 (N_8736,N_2596,N_605);
nand U8737 (N_8737,N_1685,N_4861);
nand U8738 (N_8738,N_4539,N_3051);
or U8739 (N_8739,N_3025,N_996);
nor U8740 (N_8740,N_2265,N_467);
xor U8741 (N_8741,N_4364,N_4763);
and U8742 (N_8742,N_1329,N_2679);
and U8743 (N_8743,N_2987,N_3719);
nand U8744 (N_8744,N_2892,N_2635);
nand U8745 (N_8745,N_856,N_414);
and U8746 (N_8746,N_1125,N_3414);
nor U8747 (N_8747,N_3005,N_787);
and U8748 (N_8748,N_4130,N_4194);
xor U8749 (N_8749,N_457,N_2743);
or U8750 (N_8750,N_2666,N_972);
or U8751 (N_8751,N_145,N_4588);
xor U8752 (N_8752,N_4667,N_2218);
nand U8753 (N_8753,N_2256,N_4003);
and U8754 (N_8754,N_3905,N_1724);
nor U8755 (N_8755,N_1217,N_1372);
nand U8756 (N_8756,N_4813,N_4185);
nand U8757 (N_8757,N_3380,N_3072);
xnor U8758 (N_8758,N_4194,N_671);
nand U8759 (N_8759,N_183,N_2041);
nor U8760 (N_8760,N_2947,N_961);
xor U8761 (N_8761,N_967,N_2265);
or U8762 (N_8762,N_329,N_898);
and U8763 (N_8763,N_2264,N_4330);
xnor U8764 (N_8764,N_3317,N_1108);
xor U8765 (N_8765,N_2783,N_4155);
nor U8766 (N_8766,N_1286,N_4461);
and U8767 (N_8767,N_4871,N_3662);
and U8768 (N_8768,N_332,N_2133);
or U8769 (N_8769,N_2432,N_2721);
nor U8770 (N_8770,N_4089,N_4288);
and U8771 (N_8771,N_241,N_4805);
nand U8772 (N_8772,N_3789,N_2459);
or U8773 (N_8773,N_2543,N_4343);
or U8774 (N_8774,N_4588,N_2169);
or U8775 (N_8775,N_78,N_363);
nand U8776 (N_8776,N_687,N_2070);
and U8777 (N_8777,N_1777,N_4411);
and U8778 (N_8778,N_434,N_3884);
or U8779 (N_8779,N_1928,N_1388);
xor U8780 (N_8780,N_3002,N_2533);
nand U8781 (N_8781,N_2351,N_559);
nand U8782 (N_8782,N_1954,N_2122);
or U8783 (N_8783,N_2947,N_3653);
nor U8784 (N_8784,N_4736,N_2746);
nor U8785 (N_8785,N_4273,N_2743);
nor U8786 (N_8786,N_2798,N_2703);
or U8787 (N_8787,N_838,N_711);
or U8788 (N_8788,N_821,N_1126);
or U8789 (N_8789,N_468,N_4720);
and U8790 (N_8790,N_4408,N_2429);
or U8791 (N_8791,N_2918,N_956);
nand U8792 (N_8792,N_897,N_4278);
and U8793 (N_8793,N_2753,N_2094);
or U8794 (N_8794,N_2543,N_4947);
and U8795 (N_8795,N_4260,N_4690);
nor U8796 (N_8796,N_353,N_2695);
or U8797 (N_8797,N_4637,N_519);
nand U8798 (N_8798,N_4240,N_2651);
and U8799 (N_8799,N_1864,N_1302);
nand U8800 (N_8800,N_4568,N_2866);
and U8801 (N_8801,N_4941,N_1700);
nor U8802 (N_8802,N_368,N_2944);
and U8803 (N_8803,N_4728,N_4791);
nand U8804 (N_8804,N_921,N_419);
nand U8805 (N_8805,N_4022,N_1745);
or U8806 (N_8806,N_89,N_3525);
nand U8807 (N_8807,N_4518,N_774);
and U8808 (N_8808,N_1368,N_50);
nand U8809 (N_8809,N_4299,N_3494);
nand U8810 (N_8810,N_1769,N_2250);
or U8811 (N_8811,N_1742,N_3705);
nand U8812 (N_8812,N_2925,N_808);
xor U8813 (N_8813,N_1381,N_4006);
and U8814 (N_8814,N_3079,N_2811);
nand U8815 (N_8815,N_1853,N_33);
and U8816 (N_8816,N_1267,N_3584);
or U8817 (N_8817,N_1483,N_3192);
nand U8818 (N_8818,N_275,N_4154);
nor U8819 (N_8819,N_2555,N_837);
nand U8820 (N_8820,N_630,N_2607);
and U8821 (N_8821,N_3981,N_1259);
or U8822 (N_8822,N_990,N_4052);
nor U8823 (N_8823,N_458,N_4351);
or U8824 (N_8824,N_4754,N_1999);
and U8825 (N_8825,N_3956,N_341);
nor U8826 (N_8826,N_3086,N_3470);
nand U8827 (N_8827,N_4971,N_1266);
nor U8828 (N_8828,N_2023,N_3164);
or U8829 (N_8829,N_1610,N_4415);
nor U8830 (N_8830,N_2760,N_4327);
xor U8831 (N_8831,N_1873,N_3952);
nor U8832 (N_8832,N_4953,N_93);
and U8833 (N_8833,N_2410,N_740);
nor U8834 (N_8834,N_4350,N_3461);
and U8835 (N_8835,N_579,N_2886);
and U8836 (N_8836,N_1282,N_2633);
and U8837 (N_8837,N_2481,N_2763);
or U8838 (N_8838,N_2714,N_793);
xnor U8839 (N_8839,N_4582,N_1464);
or U8840 (N_8840,N_3534,N_3998);
xor U8841 (N_8841,N_804,N_4062);
nand U8842 (N_8842,N_1787,N_2251);
and U8843 (N_8843,N_4305,N_4635);
nor U8844 (N_8844,N_3536,N_4862);
nand U8845 (N_8845,N_3346,N_2273);
nor U8846 (N_8846,N_900,N_1426);
or U8847 (N_8847,N_1913,N_610);
nand U8848 (N_8848,N_1295,N_553);
or U8849 (N_8849,N_2227,N_3353);
and U8850 (N_8850,N_2843,N_3056);
and U8851 (N_8851,N_2646,N_904);
and U8852 (N_8852,N_906,N_1762);
or U8853 (N_8853,N_2491,N_1509);
and U8854 (N_8854,N_946,N_3215);
or U8855 (N_8855,N_3756,N_1732);
or U8856 (N_8856,N_1755,N_3697);
nor U8857 (N_8857,N_4021,N_3285);
and U8858 (N_8858,N_422,N_2043);
or U8859 (N_8859,N_2368,N_3828);
and U8860 (N_8860,N_213,N_2852);
and U8861 (N_8861,N_3369,N_3493);
and U8862 (N_8862,N_3182,N_3353);
nor U8863 (N_8863,N_4290,N_2387);
nand U8864 (N_8864,N_134,N_3395);
xor U8865 (N_8865,N_2754,N_3016);
nand U8866 (N_8866,N_2360,N_3738);
xor U8867 (N_8867,N_3458,N_3190);
and U8868 (N_8868,N_1447,N_4057);
or U8869 (N_8869,N_3928,N_3219);
and U8870 (N_8870,N_258,N_4031);
xnor U8871 (N_8871,N_3581,N_539);
or U8872 (N_8872,N_143,N_2611);
or U8873 (N_8873,N_4257,N_497);
nor U8874 (N_8874,N_1113,N_4136);
nand U8875 (N_8875,N_1773,N_2403);
nor U8876 (N_8876,N_3764,N_4241);
and U8877 (N_8877,N_1454,N_3307);
nor U8878 (N_8878,N_1781,N_1363);
or U8879 (N_8879,N_4462,N_4209);
nand U8880 (N_8880,N_162,N_2169);
nor U8881 (N_8881,N_1726,N_2901);
or U8882 (N_8882,N_3449,N_3589);
xnor U8883 (N_8883,N_1120,N_1774);
and U8884 (N_8884,N_1148,N_1239);
and U8885 (N_8885,N_3623,N_2297);
or U8886 (N_8886,N_332,N_4910);
nand U8887 (N_8887,N_3243,N_3516);
or U8888 (N_8888,N_498,N_4186);
xnor U8889 (N_8889,N_1985,N_3863);
nor U8890 (N_8890,N_2990,N_3141);
or U8891 (N_8891,N_2569,N_89);
and U8892 (N_8892,N_1622,N_2236);
or U8893 (N_8893,N_2552,N_3840);
nand U8894 (N_8894,N_4959,N_1907);
xnor U8895 (N_8895,N_2233,N_1308);
nand U8896 (N_8896,N_821,N_2493);
nand U8897 (N_8897,N_853,N_189);
or U8898 (N_8898,N_3541,N_3538);
or U8899 (N_8899,N_2320,N_3736);
nand U8900 (N_8900,N_4556,N_95);
xnor U8901 (N_8901,N_4304,N_4805);
xor U8902 (N_8902,N_1758,N_1333);
nor U8903 (N_8903,N_4237,N_2523);
nand U8904 (N_8904,N_4490,N_1937);
nand U8905 (N_8905,N_200,N_889);
nand U8906 (N_8906,N_120,N_634);
and U8907 (N_8907,N_47,N_3682);
and U8908 (N_8908,N_2478,N_229);
nor U8909 (N_8909,N_2603,N_1597);
and U8910 (N_8910,N_1187,N_11);
nand U8911 (N_8911,N_531,N_1635);
or U8912 (N_8912,N_2457,N_2627);
or U8913 (N_8913,N_3972,N_2782);
nand U8914 (N_8914,N_4631,N_2954);
nand U8915 (N_8915,N_2163,N_1726);
or U8916 (N_8916,N_1016,N_2597);
nand U8917 (N_8917,N_3715,N_1571);
xor U8918 (N_8918,N_16,N_4182);
nand U8919 (N_8919,N_3389,N_4804);
or U8920 (N_8920,N_877,N_430);
and U8921 (N_8921,N_2538,N_3018);
nand U8922 (N_8922,N_116,N_561);
nand U8923 (N_8923,N_355,N_4953);
nand U8924 (N_8924,N_118,N_1601);
nand U8925 (N_8925,N_4065,N_1980);
or U8926 (N_8926,N_2941,N_3315);
and U8927 (N_8927,N_191,N_2388);
nor U8928 (N_8928,N_3660,N_2755);
nand U8929 (N_8929,N_564,N_2270);
and U8930 (N_8930,N_1486,N_4195);
and U8931 (N_8931,N_3883,N_2788);
nand U8932 (N_8932,N_3769,N_4264);
or U8933 (N_8933,N_3692,N_105);
nor U8934 (N_8934,N_447,N_1865);
and U8935 (N_8935,N_4384,N_3165);
and U8936 (N_8936,N_1511,N_2096);
nand U8937 (N_8937,N_2935,N_3118);
nand U8938 (N_8938,N_2586,N_1812);
or U8939 (N_8939,N_314,N_2017);
and U8940 (N_8940,N_748,N_4856);
xor U8941 (N_8941,N_1234,N_4983);
and U8942 (N_8942,N_1343,N_552);
nand U8943 (N_8943,N_1679,N_4619);
and U8944 (N_8944,N_368,N_4623);
or U8945 (N_8945,N_3075,N_471);
or U8946 (N_8946,N_875,N_854);
and U8947 (N_8947,N_1419,N_4077);
and U8948 (N_8948,N_2571,N_715);
nand U8949 (N_8949,N_2824,N_4098);
xnor U8950 (N_8950,N_1789,N_3164);
nand U8951 (N_8951,N_3572,N_3930);
nor U8952 (N_8952,N_635,N_1458);
or U8953 (N_8953,N_2061,N_2176);
nand U8954 (N_8954,N_1175,N_3779);
nor U8955 (N_8955,N_3046,N_2185);
nand U8956 (N_8956,N_2282,N_2782);
or U8957 (N_8957,N_4843,N_4334);
or U8958 (N_8958,N_191,N_4013);
or U8959 (N_8959,N_2809,N_3937);
nand U8960 (N_8960,N_2003,N_2174);
or U8961 (N_8961,N_2401,N_1096);
nand U8962 (N_8962,N_1650,N_4115);
nand U8963 (N_8963,N_3565,N_4566);
or U8964 (N_8964,N_3058,N_2829);
and U8965 (N_8965,N_995,N_4933);
nor U8966 (N_8966,N_264,N_1900);
or U8967 (N_8967,N_2150,N_342);
and U8968 (N_8968,N_737,N_1624);
or U8969 (N_8969,N_81,N_4911);
nor U8970 (N_8970,N_499,N_4614);
nor U8971 (N_8971,N_3931,N_2756);
and U8972 (N_8972,N_4555,N_3190);
nor U8973 (N_8973,N_3069,N_3650);
nor U8974 (N_8974,N_1315,N_648);
nand U8975 (N_8975,N_396,N_2431);
nor U8976 (N_8976,N_4014,N_4339);
nand U8977 (N_8977,N_4687,N_52);
nand U8978 (N_8978,N_1859,N_842);
nand U8979 (N_8979,N_4900,N_638);
and U8980 (N_8980,N_3798,N_1869);
nor U8981 (N_8981,N_2273,N_3385);
or U8982 (N_8982,N_2061,N_3250);
nand U8983 (N_8983,N_1138,N_2603);
nor U8984 (N_8984,N_2986,N_868);
nand U8985 (N_8985,N_3021,N_1499);
and U8986 (N_8986,N_4110,N_2540);
nand U8987 (N_8987,N_1516,N_1975);
and U8988 (N_8988,N_2502,N_1400);
nor U8989 (N_8989,N_2072,N_3940);
nand U8990 (N_8990,N_4089,N_1680);
and U8991 (N_8991,N_2214,N_474);
and U8992 (N_8992,N_2956,N_3909);
or U8993 (N_8993,N_1912,N_3187);
or U8994 (N_8994,N_2208,N_1654);
nor U8995 (N_8995,N_1893,N_1443);
or U8996 (N_8996,N_4272,N_3743);
or U8997 (N_8997,N_2910,N_4515);
and U8998 (N_8998,N_342,N_3754);
and U8999 (N_8999,N_3801,N_426);
nand U9000 (N_9000,N_4990,N_4214);
nor U9001 (N_9001,N_1584,N_2204);
nand U9002 (N_9002,N_3760,N_2720);
nor U9003 (N_9003,N_2601,N_455);
and U9004 (N_9004,N_3574,N_3444);
and U9005 (N_9005,N_2008,N_3766);
and U9006 (N_9006,N_422,N_1984);
xor U9007 (N_9007,N_3214,N_1737);
or U9008 (N_9008,N_3930,N_157);
or U9009 (N_9009,N_1315,N_278);
and U9010 (N_9010,N_1233,N_74);
nor U9011 (N_9011,N_2043,N_3168);
nor U9012 (N_9012,N_1571,N_1204);
nand U9013 (N_9013,N_3966,N_566);
nand U9014 (N_9014,N_3281,N_2780);
xor U9015 (N_9015,N_3881,N_2182);
nand U9016 (N_9016,N_1453,N_3341);
and U9017 (N_9017,N_3538,N_1722);
and U9018 (N_9018,N_154,N_3089);
nand U9019 (N_9019,N_4167,N_1287);
or U9020 (N_9020,N_1979,N_936);
and U9021 (N_9021,N_633,N_2466);
and U9022 (N_9022,N_4507,N_4400);
and U9023 (N_9023,N_1598,N_3540);
nor U9024 (N_9024,N_4913,N_226);
xor U9025 (N_9025,N_201,N_1400);
and U9026 (N_9026,N_3285,N_940);
xnor U9027 (N_9027,N_3581,N_1537);
or U9028 (N_9028,N_3233,N_2927);
nand U9029 (N_9029,N_3661,N_3848);
or U9030 (N_9030,N_73,N_3630);
nand U9031 (N_9031,N_2045,N_2442);
or U9032 (N_9032,N_841,N_2811);
nor U9033 (N_9033,N_812,N_612);
xor U9034 (N_9034,N_2482,N_2230);
nand U9035 (N_9035,N_932,N_737);
or U9036 (N_9036,N_3328,N_223);
and U9037 (N_9037,N_3834,N_3519);
nand U9038 (N_9038,N_476,N_550);
xor U9039 (N_9039,N_2160,N_68);
and U9040 (N_9040,N_706,N_960);
nor U9041 (N_9041,N_2377,N_1007);
nand U9042 (N_9042,N_1872,N_3349);
nor U9043 (N_9043,N_3820,N_1745);
nor U9044 (N_9044,N_1939,N_1894);
nand U9045 (N_9045,N_1264,N_4628);
nand U9046 (N_9046,N_3158,N_2181);
and U9047 (N_9047,N_1106,N_3963);
xnor U9048 (N_9048,N_803,N_2194);
nand U9049 (N_9049,N_3552,N_2542);
xnor U9050 (N_9050,N_3976,N_2822);
xnor U9051 (N_9051,N_2280,N_1981);
or U9052 (N_9052,N_711,N_3890);
xor U9053 (N_9053,N_172,N_3490);
nand U9054 (N_9054,N_1400,N_4473);
or U9055 (N_9055,N_389,N_701);
nand U9056 (N_9056,N_2763,N_1488);
or U9057 (N_9057,N_4255,N_3133);
or U9058 (N_9058,N_3920,N_1643);
nand U9059 (N_9059,N_937,N_3516);
nor U9060 (N_9060,N_2508,N_11);
and U9061 (N_9061,N_4381,N_1959);
or U9062 (N_9062,N_3562,N_401);
nor U9063 (N_9063,N_3657,N_2970);
or U9064 (N_9064,N_2191,N_1136);
xor U9065 (N_9065,N_3053,N_2121);
xnor U9066 (N_9066,N_1023,N_3395);
nand U9067 (N_9067,N_4319,N_4122);
nand U9068 (N_9068,N_4375,N_3195);
or U9069 (N_9069,N_791,N_1712);
and U9070 (N_9070,N_2264,N_1305);
nand U9071 (N_9071,N_2495,N_955);
nand U9072 (N_9072,N_38,N_4434);
and U9073 (N_9073,N_87,N_436);
nand U9074 (N_9074,N_4969,N_4028);
and U9075 (N_9075,N_620,N_1837);
nor U9076 (N_9076,N_61,N_900);
or U9077 (N_9077,N_4334,N_1256);
nor U9078 (N_9078,N_1298,N_120);
and U9079 (N_9079,N_506,N_24);
or U9080 (N_9080,N_3266,N_1327);
nand U9081 (N_9081,N_1176,N_2445);
xnor U9082 (N_9082,N_1475,N_3752);
nor U9083 (N_9083,N_848,N_4198);
and U9084 (N_9084,N_2513,N_601);
or U9085 (N_9085,N_439,N_1135);
and U9086 (N_9086,N_1897,N_3817);
or U9087 (N_9087,N_4634,N_602);
nand U9088 (N_9088,N_2787,N_3586);
nand U9089 (N_9089,N_3568,N_1908);
nor U9090 (N_9090,N_1339,N_2778);
and U9091 (N_9091,N_410,N_4063);
and U9092 (N_9092,N_1276,N_3186);
nand U9093 (N_9093,N_1111,N_2106);
nand U9094 (N_9094,N_3430,N_4204);
or U9095 (N_9095,N_4449,N_2055);
or U9096 (N_9096,N_180,N_2592);
nand U9097 (N_9097,N_1103,N_4102);
nor U9098 (N_9098,N_3799,N_525);
nor U9099 (N_9099,N_3285,N_750);
xor U9100 (N_9100,N_2400,N_2038);
and U9101 (N_9101,N_2773,N_566);
nand U9102 (N_9102,N_3724,N_4591);
nor U9103 (N_9103,N_4030,N_483);
nand U9104 (N_9104,N_4535,N_111);
or U9105 (N_9105,N_614,N_4590);
or U9106 (N_9106,N_1542,N_377);
or U9107 (N_9107,N_167,N_2806);
nand U9108 (N_9108,N_1964,N_3767);
nand U9109 (N_9109,N_4676,N_751);
and U9110 (N_9110,N_4794,N_37);
nand U9111 (N_9111,N_1927,N_3093);
nand U9112 (N_9112,N_3141,N_1332);
nor U9113 (N_9113,N_3111,N_3098);
nand U9114 (N_9114,N_3629,N_2203);
and U9115 (N_9115,N_1894,N_308);
and U9116 (N_9116,N_4406,N_4469);
nand U9117 (N_9117,N_4324,N_2188);
nor U9118 (N_9118,N_4512,N_2171);
nor U9119 (N_9119,N_1142,N_2369);
or U9120 (N_9120,N_2614,N_2472);
nand U9121 (N_9121,N_1115,N_2021);
nand U9122 (N_9122,N_836,N_2601);
or U9123 (N_9123,N_1143,N_3730);
and U9124 (N_9124,N_626,N_4663);
nand U9125 (N_9125,N_1833,N_4160);
or U9126 (N_9126,N_830,N_1651);
nand U9127 (N_9127,N_2136,N_2703);
nor U9128 (N_9128,N_1916,N_1154);
and U9129 (N_9129,N_440,N_2407);
and U9130 (N_9130,N_757,N_470);
nand U9131 (N_9131,N_2196,N_305);
or U9132 (N_9132,N_2618,N_3698);
nand U9133 (N_9133,N_753,N_4938);
nor U9134 (N_9134,N_4594,N_697);
xor U9135 (N_9135,N_1836,N_3293);
or U9136 (N_9136,N_1832,N_1802);
and U9137 (N_9137,N_2016,N_1715);
nor U9138 (N_9138,N_4253,N_3899);
xnor U9139 (N_9139,N_3893,N_4198);
or U9140 (N_9140,N_2952,N_3791);
nand U9141 (N_9141,N_2710,N_4786);
nor U9142 (N_9142,N_3823,N_2512);
or U9143 (N_9143,N_4763,N_3861);
and U9144 (N_9144,N_2521,N_3282);
xnor U9145 (N_9145,N_1210,N_3760);
and U9146 (N_9146,N_1141,N_2819);
and U9147 (N_9147,N_4197,N_8);
and U9148 (N_9148,N_4740,N_4626);
or U9149 (N_9149,N_239,N_2951);
nand U9150 (N_9150,N_1680,N_4807);
or U9151 (N_9151,N_3391,N_3023);
nor U9152 (N_9152,N_4942,N_3572);
nor U9153 (N_9153,N_3807,N_2987);
and U9154 (N_9154,N_1837,N_3651);
nor U9155 (N_9155,N_277,N_1280);
nor U9156 (N_9156,N_241,N_975);
nand U9157 (N_9157,N_996,N_1945);
and U9158 (N_9158,N_3067,N_4372);
nand U9159 (N_9159,N_3085,N_4186);
nand U9160 (N_9160,N_1975,N_3266);
nand U9161 (N_9161,N_2385,N_2722);
xnor U9162 (N_9162,N_1678,N_4047);
or U9163 (N_9163,N_3552,N_2897);
or U9164 (N_9164,N_3779,N_4708);
nor U9165 (N_9165,N_4107,N_4001);
nor U9166 (N_9166,N_1481,N_1694);
xor U9167 (N_9167,N_3113,N_2358);
xor U9168 (N_9168,N_1210,N_2447);
nand U9169 (N_9169,N_610,N_850);
and U9170 (N_9170,N_4544,N_2062);
nand U9171 (N_9171,N_1786,N_3601);
xnor U9172 (N_9172,N_1333,N_3916);
nor U9173 (N_9173,N_4043,N_3919);
nand U9174 (N_9174,N_977,N_1126);
nor U9175 (N_9175,N_4821,N_4705);
xor U9176 (N_9176,N_4204,N_4127);
nor U9177 (N_9177,N_4539,N_2433);
nor U9178 (N_9178,N_1328,N_3703);
and U9179 (N_9179,N_4844,N_4471);
or U9180 (N_9180,N_1392,N_751);
and U9181 (N_9181,N_1648,N_4664);
xnor U9182 (N_9182,N_1865,N_2745);
nor U9183 (N_9183,N_4091,N_2516);
nand U9184 (N_9184,N_3800,N_2023);
or U9185 (N_9185,N_217,N_2374);
nor U9186 (N_9186,N_1009,N_3263);
nand U9187 (N_9187,N_4512,N_133);
xnor U9188 (N_9188,N_3028,N_3217);
and U9189 (N_9189,N_2956,N_1262);
xnor U9190 (N_9190,N_2608,N_420);
or U9191 (N_9191,N_2477,N_506);
nor U9192 (N_9192,N_2347,N_2841);
or U9193 (N_9193,N_1985,N_4231);
or U9194 (N_9194,N_4446,N_3715);
nand U9195 (N_9195,N_2467,N_4954);
or U9196 (N_9196,N_2508,N_1820);
or U9197 (N_9197,N_4809,N_1242);
xor U9198 (N_9198,N_3084,N_494);
nor U9199 (N_9199,N_2606,N_241);
nand U9200 (N_9200,N_4292,N_4640);
and U9201 (N_9201,N_708,N_127);
nand U9202 (N_9202,N_4327,N_4705);
nand U9203 (N_9203,N_4888,N_4548);
xor U9204 (N_9204,N_3282,N_2126);
nand U9205 (N_9205,N_3567,N_2634);
or U9206 (N_9206,N_3369,N_1648);
nor U9207 (N_9207,N_1971,N_4380);
nand U9208 (N_9208,N_2582,N_3454);
or U9209 (N_9209,N_3990,N_4627);
nand U9210 (N_9210,N_3058,N_2047);
nand U9211 (N_9211,N_2961,N_3320);
or U9212 (N_9212,N_1821,N_3417);
or U9213 (N_9213,N_956,N_350);
nand U9214 (N_9214,N_4193,N_1599);
nor U9215 (N_9215,N_2354,N_136);
and U9216 (N_9216,N_4528,N_2128);
nand U9217 (N_9217,N_1433,N_676);
xnor U9218 (N_9218,N_3334,N_2205);
nor U9219 (N_9219,N_684,N_2678);
nand U9220 (N_9220,N_1818,N_1948);
xor U9221 (N_9221,N_4045,N_1907);
and U9222 (N_9222,N_2431,N_316);
or U9223 (N_9223,N_3483,N_354);
nor U9224 (N_9224,N_3946,N_990);
xor U9225 (N_9225,N_485,N_1587);
nor U9226 (N_9226,N_1591,N_4712);
xnor U9227 (N_9227,N_3059,N_808);
and U9228 (N_9228,N_297,N_2192);
nand U9229 (N_9229,N_2582,N_2001);
and U9230 (N_9230,N_3154,N_1142);
or U9231 (N_9231,N_48,N_2287);
nor U9232 (N_9232,N_4909,N_2433);
or U9233 (N_9233,N_1357,N_596);
nand U9234 (N_9234,N_179,N_2725);
nor U9235 (N_9235,N_2318,N_4299);
and U9236 (N_9236,N_1447,N_872);
nand U9237 (N_9237,N_4853,N_298);
and U9238 (N_9238,N_4505,N_4696);
or U9239 (N_9239,N_2871,N_1692);
and U9240 (N_9240,N_2654,N_2703);
nor U9241 (N_9241,N_785,N_1138);
and U9242 (N_9242,N_1568,N_4999);
or U9243 (N_9243,N_2302,N_1385);
and U9244 (N_9244,N_1192,N_2494);
and U9245 (N_9245,N_4580,N_4889);
or U9246 (N_9246,N_2145,N_1387);
or U9247 (N_9247,N_2203,N_1585);
nor U9248 (N_9248,N_3078,N_1640);
nand U9249 (N_9249,N_3241,N_2510);
nand U9250 (N_9250,N_379,N_2065);
nand U9251 (N_9251,N_4029,N_4575);
nand U9252 (N_9252,N_21,N_4798);
or U9253 (N_9253,N_4117,N_2199);
or U9254 (N_9254,N_4850,N_1942);
nand U9255 (N_9255,N_3091,N_408);
and U9256 (N_9256,N_399,N_4235);
nand U9257 (N_9257,N_3602,N_2583);
nor U9258 (N_9258,N_309,N_1757);
or U9259 (N_9259,N_4036,N_3142);
or U9260 (N_9260,N_325,N_432);
and U9261 (N_9261,N_400,N_38);
nand U9262 (N_9262,N_4549,N_1715);
nor U9263 (N_9263,N_2185,N_2589);
or U9264 (N_9264,N_1842,N_3242);
or U9265 (N_9265,N_1484,N_252);
nor U9266 (N_9266,N_3828,N_2097);
nor U9267 (N_9267,N_3293,N_3760);
nor U9268 (N_9268,N_3555,N_2928);
nor U9269 (N_9269,N_1866,N_2945);
or U9270 (N_9270,N_518,N_1653);
nor U9271 (N_9271,N_1187,N_1100);
or U9272 (N_9272,N_3481,N_4361);
or U9273 (N_9273,N_1392,N_1166);
nand U9274 (N_9274,N_238,N_2590);
or U9275 (N_9275,N_2057,N_445);
nand U9276 (N_9276,N_4879,N_2518);
nor U9277 (N_9277,N_2021,N_3292);
nor U9278 (N_9278,N_3419,N_3448);
or U9279 (N_9279,N_4043,N_2183);
or U9280 (N_9280,N_1209,N_3468);
nand U9281 (N_9281,N_4507,N_1868);
or U9282 (N_9282,N_150,N_1755);
or U9283 (N_9283,N_2874,N_1246);
and U9284 (N_9284,N_3055,N_2081);
xnor U9285 (N_9285,N_433,N_4892);
nor U9286 (N_9286,N_1445,N_198);
or U9287 (N_9287,N_1871,N_4812);
nand U9288 (N_9288,N_4981,N_4298);
and U9289 (N_9289,N_2043,N_3400);
or U9290 (N_9290,N_2960,N_1753);
and U9291 (N_9291,N_4462,N_3520);
and U9292 (N_9292,N_4300,N_4845);
nor U9293 (N_9293,N_3633,N_692);
nor U9294 (N_9294,N_2893,N_3991);
nor U9295 (N_9295,N_410,N_2791);
nand U9296 (N_9296,N_1074,N_3042);
or U9297 (N_9297,N_1863,N_4179);
or U9298 (N_9298,N_1657,N_870);
and U9299 (N_9299,N_1421,N_4019);
nor U9300 (N_9300,N_1509,N_4028);
nand U9301 (N_9301,N_1467,N_687);
xnor U9302 (N_9302,N_4358,N_2961);
xnor U9303 (N_9303,N_2525,N_2268);
nand U9304 (N_9304,N_925,N_733);
and U9305 (N_9305,N_3321,N_999);
and U9306 (N_9306,N_3633,N_3207);
nor U9307 (N_9307,N_921,N_88);
or U9308 (N_9308,N_1869,N_4195);
nor U9309 (N_9309,N_2036,N_4878);
or U9310 (N_9310,N_2219,N_4826);
or U9311 (N_9311,N_1960,N_4265);
nand U9312 (N_9312,N_4779,N_2058);
or U9313 (N_9313,N_2453,N_1566);
nand U9314 (N_9314,N_379,N_601);
xor U9315 (N_9315,N_1582,N_4193);
nand U9316 (N_9316,N_2300,N_3657);
or U9317 (N_9317,N_2933,N_282);
nand U9318 (N_9318,N_1460,N_319);
or U9319 (N_9319,N_1728,N_990);
and U9320 (N_9320,N_949,N_2610);
nand U9321 (N_9321,N_4714,N_464);
nand U9322 (N_9322,N_1015,N_4565);
and U9323 (N_9323,N_3619,N_3819);
xnor U9324 (N_9324,N_2471,N_3635);
and U9325 (N_9325,N_4432,N_1451);
or U9326 (N_9326,N_3094,N_3825);
nor U9327 (N_9327,N_61,N_2545);
nand U9328 (N_9328,N_1643,N_3219);
nor U9329 (N_9329,N_446,N_506);
or U9330 (N_9330,N_4069,N_3065);
and U9331 (N_9331,N_312,N_1511);
nor U9332 (N_9332,N_1037,N_3231);
or U9333 (N_9333,N_142,N_4828);
nor U9334 (N_9334,N_2041,N_3914);
nor U9335 (N_9335,N_2155,N_4776);
nor U9336 (N_9336,N_4314,N_1883);
nor U9337 (N_9337,N_642,N_3746);
and U9338 (N_9338,N_1866,N_3206);
nor U9339 (N_9339,N_1767,N_1028);
nand U9340 (N_9340,N_4756,N_3341);
xor U9341 (N_9341,N_3970,N_3305);
nor U9342 (N_9342,N_4715,N_2317);
or U9343 (N_9343,N_2815,N_320);
and U9344 (N_9344,N_226,N_834);
nand U9345 (N_9345,N_340,N_3234);
xor U9346 (N_9346,N_4221,N_4559);
nand U9347 (N_9347,N_4829,N_3091);
and U9348 (N_9348,N_4191,N_47);
or U9349 (N_9349,N_4854,N_3680);
or U9350 (N_9350,N_931,N_3360);
or U9351 (N_9351,N_2914,N_240);
nor U9352 (N_9352,N_4510,N_2426);
nand U9353 (N_9353,N_4219,N_3200);
nor U9354 (N_9354,N_1997,N_4739);
or U9355 (N_9355,N_1795,N_1620);
nand U9356 (N_9356,N_2896,N_2775);
xor U9357 (N_9357,N_4103,N_424);
nand U9358 (N_9358,N_3271,N_3445);
and U9359 (N_9359,N_4911,N_2392);
and U9360 (N_9360,N_3611,N_1362);
nand U9361 (N_9361,N_1030,N_1744);
or U9362 (N_9362,N_3933,N_1224);
nand U9363 (N_9363,N_38,N_2813);
and U9364 (N_9364,N_4690,N_2055);
nor U9365 (N_9365,N_2989,N_1886);
nand U9366 (N_9366,N_1841,N_4684);
nor U9367 (N_9367,N_1451,N_4152);
nand U9368 (N_9368,N_505,N_4071);
nor U9369 (N_9369,N_1339,N_3485);
nor U9370 (N_9370,N_2962,N_482);
nand U9371 (N_9371,N_327,N_1471);
nor U9372 (N_9372,N_1559,N_341);
nor U9373 (N_9373,N_724,N_4717);
and U9374 (N_9374,N_2881,N_4686);
or U9375 (N_9375,N_3783,N_2831);
and U9376 (N_9376,N_114,N_3745);
xnor U9377 (N_9377,N_4952,N_2511);
and U9378 (N_9378,N_1942,N_4922);
nand U9379 (N_9379,N_854,N_3476);
or U9380 (N_9380,N_190,N_4190);
nor U9381 (N_9381,N_1497,N_4285);
xor U9382 (N_9382,N_2727,N_152);
nand U9383 (N_9383,N_4193,N_3724);
nor U9384 (N_9384,N_3139,N_72);
and U9385 (N_9385,N_3358,N_307);
xnor U9386 (N_9386,N_591,N_4542);
nand U9387 (N_9387,N_4695,N_792);
nor U9388 (N_9388,N_3309,N_2499);
nand U9389 (N_9389,N_407,N_37);
nor U9390 (N_9390,N_657,N_3572);
nand U9391 (N_9391,N_3198,N_4435);
xnor U9392 (N_9392,N_4930,N_3569);
nor U9393 (N_9393,N_189,N_1971);
or U9394 (N_9394,N_2456,N_3837);
or U9395 (N_9395,N_183,N_3697);
and U9396 (N_9396,N_4167,N_3958);
xor U9397 (N_9397,N_4066,N_2403);
nor U9398 (N_9398,N_341,N_3764);
nor U9399 (N_9399,N_4197,N_113);
nor U9400 (N_9400,N_4655,N_3355);
nor U9401 (N_9401,N_3202,N_1196);
nand U9402 (N_9402,N_2677,N_3303);
xnor U9403 (N_9403,N_970,N_3759);
xor U9404 (N_9404,N_207,N_4029);
xor U9405 (N_9405,N_2136,N_3174);
nor U9406 (N_9406,N_3304,N_4209);
nand U9407 (N_9407,N_2261,N_4879);
xor U9408 (N_9408,N_4668,N_2574);
and U9409 (N_9409,N_4073,N_4282);
nand U9410 (N_9410,N_303,N_617);
nor U9411 (N_9411,N_4962,N_3947);
and U9412 (N_9412,N_3719,N_3633);
or U9413 (N_9413,N_4907,N_4305);
nor U9414 (N_9414,N_4267,N_1683);
nand U9415 (N_9415,N_2717,N_3225);
nor U9416 (N_9416,N_2510,N_4965);
nor U9417 (N_9417,N_2388,N_3673);
or U9418 (N_9418,N_605,N_986);
nor U9419 (N_9419,N_4852,N_3683);
or U9420 (N_9420,N_1909,N_3237);
nor U9421 (N_9421,N_3180,N_2031);
nor U9422 (N_9422,N_1260,N_3528);
and U9423 (N_9423,N_1743,N_931);
nor U9424 (N_9424,N_4003,N_3181);
and U9425 (N_9425,N_4973,N_400);
and U9426 (N_9426,N_1220,N_3363);
xnor U9427 (N_9427,N_780,N_3261);
or U9428 (N_9428,N_3081,N_1888);
and U9429 (N_9429,N_2047,N_3578);
or U9430 (N_9430,N_859,N_4246);
and U9431 (N_9431,N_3616,N_1822);
nand U9432 (N_9432,N_2312,N_117);
nor U9433 (N_9433,N_504,N_2112);
xor U9434 (N_9434,N_2394,N_3005);
nor U9435 (N_9435,N_210,N_4528);
or U9436 (N_9436,N_1180,N_3255);
xor U9437 (N_9437,N_359,N_4161);
and U9438 (N_9438,N_322,N_1764);
nor U9439 (N_9439,N_1389,N_4095);
nand U9440 (N_9440,N_912,N_2833);
nand U9441 (N_9441,N_4335,N_810);
nand U9442 (N_9442,N_453,N_2499);
nor U9443 (N_9443,N_1448,N_4382);
nand U9444 (N_9444,N_1054,N_2078);
and U9445 (N_9445,N_3772,N_3105);
and U9446 (N_9446,N_3484,N_4020);
or U9447 (N_9447,N_3210,N_4912);
or U9448 (N_9448,N_35,N_1542);
or U9449 (N_9449,N_2478,N_4006);
nand U9450 (N_9450,N_4654,N_2573);
nor U9451 (N_9451,N_1651,N_924);
nand U9452 (N_9452,N_2804,N_1893);
nor U9453 (N_9453,N_3699,N_2498);
nand U9454 (N_9454,N_4911,N_1114);
and U9455 (N_9455,N_4942,N_3787);
or U9456 (N_9456,N_3763,N_3473);
or U9457 (N_9457,N_4128,N_150);
or U9458 (N_9458,N_1594,N_4523);
or U9459 (N_9459,N_2635,N_4412);
nand U9460 (N_9460,N_4608,N_1208);
nor U9461 (N_9461,N_3571,N_1477);
xor U9462 (N_9462,N_1953,N_957);
and U9463 (N_9463,N_3854,N_1384);
nor U9464 (N_9464,N_173,N_2289);
and U9465 (N_9465,N_2838,N_1299);
and U9466 (N_9466,N_2394,N_1948);
and U9467 (N_9467,N_1355,N_1163);
and U9468 (N_9468,N_1763,N_4114);
nor U9469 (N_9469,N_1699,N_3797);
nand U9470 (N_9470,N_2118,N_126);
and U9471 (N_9471,N_678,N_2064);
and U9472 (N_9472,N_576,N_259);
xor U9473 (N_9473,N_2998,N_1967);
nor U9474 (N_9474,N_291,N_1490);
or U9475 (N_9475,N_2825,N_1566);
nor U9476 (N_9476,N_2100,N_212);
or U9477 (N_9477,N_1139,N_2544);
and U9478 (N_9478,N_1845,N_3785);
nor U9479 (N_9479,N_4635,N_4247);
or U9480 (N_9480,N_3275,N_3053);
or U9481 (N_9481,N_56,N_182);
or U9482 (N_9482,N_1611,N_2962);
xnor U9483 (N_9483,N_1737,N_1527);
nand U9484 (N_9484,N_4781,N_3895);
xnor U9485 (N_9485,N_3450,N_1625);
and U9486 (N_9486,N_243,N_625);
nand U9487 (N_9487,N_506,N_970);
or U9488 (N_9488,N_326,N_2132);
and U9489 (N_9489,N_4034,N_4118);
nand U9490 (N_9490,N_3799,N_2201);
and U9491 (N_9491,N_3605,N_4910);
nand U9492 (N_9492,N_2606,N_4147);
xnor U9493 (N_9493,N_829,N_182);
and U9494 (N_9494,N_1258,N_3174);
nor U9495 (N_9495,N_286,N_140);
nor U9496 (N_9496,N_2650,N_4748);
or U9497 (N_9497,N_2652,N_704);
xor U9498 (N_9498,N_4948,N_4290);
nand U9499 (N_9499,N_189,N_4050);
nor U9500 (N_9500,N_1814,N_12);
and U9501 (N_9501,N_3274,N_901);
nor U9502 (N_9502,N_4884,N_4414);
or U9503 (N_9503,N_2014,N_3529);
nand U9504 (N_9504,N_3617,N_574);
and U9505 (N_9505,N_2405,N_2120);
and U9506 (N_9506,N_3556,N_699);
and U9507 (N_9507,N_4372,N_4942);
nor U9508 (N_9508,N_3568,N_354);
or U9509 (N_9509,N_3400,N_3219);
nor U9510 (N_9510,N_4826,N_4603);
nand U9511 (N_9511,N_1263,N_924);
or U9512 (N_9512,N_2377,N_1584);
or U9513 (N_9513,N_3402,N_2642);
or U9514 (N_9514,N_4795,N_3954);
and U9515 (N_9515,N_1270,N_2844);
or U9516 (N_9516,N_1872,N_4592);
and U9517 (N_9517,N_2351,N_1278);
and U9518 (N_9518,N_4786,N_2119);
or U9519 (N_9519,N_259,N_1191);
and U9520 (N_9520,N_2459,N_2869);
nand U9521 (N_9521,N_1814,N_2347);
xor U9522 (N_9522,N_3114,N_2338);
or U9523 (N_9523,N_3691,N_2011);
nor U9524 (N_9524,N_1472,N_1032);
nor U9525 (N_9525,N_3215,N_2352);
or U9526 (N_9526,N_930,N_1656);
or U9527 (N_9527,N_304,N_451);
or U9528 (N_9528,N_3959,N_2136);
or U9529 (N_9529,N_4410,N_2262);
and U9530 (N_9530,N_134,N_80);
and U9531 (N_9531,N_3181,N_1046);
or U9532 (N_9532,N_2469,N_1964);
xnor U9533 (N_9533,N_1416,N_4967);
xor U9534 (N_9534,N_1132,N_3038);
xor U9535 (N_9535,N_1524,N_342);
xnor U9536 (N_9536,N_3283,N_4686);
nand U9537 (N_9537,N_770,N_1316);
or U9538 (N_9538,N_2604,N_3524);
nand U9539 (N_9539,N_298,N_2438);
nand U9540 (N_9540,N_125,N_4758);
xnor U9541 (N_9541,N_194,N_1103);
and U9542 (N_9542,N_1221,N_3252);
and U9543 (N_9543,N_4405,N_2482);
nand U9544 (N_9544,N_3345,N_610);
nor U9545 (N_9545,N_4166,N_1678);
nor U9546 (N_9546,N_106,N_3788);
and U9547 (N_9547,N_4508,N_3137);
and U9548 (N_9548,N_4707,N_226);
nor U9549 (N_9549,N_3229,N_3076);
or U9550 (N_9550,N_610,N_4035);
nor U9551 (N_9551,N_3387,N_2304);
and U9552 (N_9552,N_1953,N_4585);
nor U9553 (N_9553,N_3043,N_3102);
xor U9554 (N_9554,N_4597,N_4201);
and U9555 (N_9555,N_4531,N_2573);
and U9556 (N_9556,N_3296,N_3417);
or U9557 (N_9557,N_1861,N_4548);
nor U9558 (N_9558,N_2025,N_4256);
xnor U9559 (N_9559,N_389,N_3639);
or U9560 (N_9560,N_1178,N_50);
or U9561 (N_9561,N_3965,N_290);
or U9562 (N_9562,N_2676,N_3885);
xnor U9563 (N_9563,N_940,N_3645);
and U9564 (N_9564,N_3872,N_1962);
nor U9565 (N_9565,N_2599,N_2838);
and U9566 (N_9566,N_4277,N_4267);
and U9567 (N_9567,N_1178,N_858);
nor U9568 (N_9568,N_8,N_698);
and U9569 (N_9569,N_541,N_3062);
and U9570 (N_9570,N_3987,N_4510);
or U9571 (N_9571,N_1200,N_4935);
or U9572 (N_9572,N_3273,N_2700);
nand U9573 (N_9573,N_609,N_3244);
xor U9574 (N_9574,N_4298,N_812);
and U9575 (N_9575,N_1899,N_3183);
and U9576 (N_9576,N_2497,N_4939);
nor U9577 (N_9577,N_4662,N_4369);
or U9578 (N_9578,N_4967,N_379);
or U9579 (N_9579,N_1626,N_3571);
and U9580 (N_9580,N_636,N_450);
nor U9581 (N_9581,N_1265,N_2309);
nor U9582 (N_9582,N_585,N_3490);
and U9583 (N_9583,N_3419,N_980);
nand U9584 (N_9584,N_2444,N_1317);
nand U9585 (N_9585,N_1512,N_3023);
nand U9586 (N_9586,N_1240,N_4407);
nor U9587 (N_9587,N_4971,N_3958);
or U9588 (N_9588,N_1865,N_4179);
and U9589 (N_9589,N_3365,N_2443);
xnor U9590 (N_9590,N_1929,N_3550);
or U9591 (N_9591,N_3463,N_2298);
or U9592 (N_9592,N_420,N_4338);
nand U9593 (N_9593,N_3651,N_3586);
and U9594 (N_9594,N_3238,N_2769);
nor U9595 (N_9595,N_1043,N_2438);
xor U9596 (N_9596,N_284,N_268);
nand U9597 (N_9597,N_3187,N_1222);
nor U9598 (N_9598,N_775,N_3676);
nor U9599 (N_9599,N_4967,N_3165);
nand U9600 (N_9600,N_793,N_4822);
and U9601 (N_9601,N_3626,N_847);
or U9602 (N_9602,N_2869,N_114);
or U9603 (N_9603,N_3550,N_1427);
xnor U9604 (N_9604,N_1248,N_401);
xnor U9605 (N_9605,N_4187,N_2804);
nand U9606 (N_9606,N_355,N_144);
or U9607 (N_9607,N_2768,N_2049);
nor U9608 (N_9608,N_3048,N_441);
and U9609 (N_9609,N_3590,N_2598);
or U9610 (N_9610,N_258,N_3513);
or U9611 (N_9611,N_4182,N_369);
nand U9612 (N_9612,N_4413,N_2233);
nand U9613 (N_9613,N_4256,N_533);
and U9614 (N_9614,N_2035,N_1704);
nand U9615 (N_9615,N_3559,N_3515);
xnor U9616 (N_9616,N_4156,N_55);
and U9617 (N_9617,N_1413,N_4408);
or U9618 (N_9618,N_209,N_1230);
and U9619 (N_9619,N_4408,N_3136);
nand U9620 (N_9620,N_3195,N_4604);
nor U9621 (N_9621,N_2135,N_1665);
xnor U9622 (N_9622,N_995,N_145);
or U9623 (N_9623,N_2328,N_3027);
nand U9624 (N_9624,N_2053,N_2643);
nand U9625 (N_9625,N_4562,N_4424);
nand U9626 (N_9626,N_2382,N_2408);
nand U9627 (N_9627,N_496,N_4837);
nand U9628 (N_9628,N_3640,N_3687);
nor U9629 (N_9629,N_434,N_51);
nor U9630 (N_9630,N_927,N_2558);
and U9631 (N_9631,N_4837,N_220);
nand U9632 (N_9632,N_940,N_1072);
or U9633 (N_9633,N_1265,N_262);
xnor U9634 (N_9634,N_1763,N_1319);
and U9635 (N_9635,N_550,N_3497);
xor U9636 (N_9636,N_2632,N_4138);
and U9637 (N_9637,N_923,N_3537);
nand U9638 (N_9638,N_2129,N_3760);
nor U9639 (N_9639,N_1416,N_3512);
or U9640 (N_9640,N_4646,N_2022);
nand U9641 (N_9641,N_235,N_3024);
or U9642 (N_9642,N_2055,N_3805);
nand U9643 (N_9643,N_3059,N_4695);
nand U9644 (N_9644,N_1851,N_2);
nor U9645 (N_9645,N_3796,N_1042);
and U9646 (N_9646,N_80,N_3804);
or U9647 (N_9647,N_1523,N_4035);
and U9648 (N_9648,N_1509,N_100);
nand U9649 (N_9649,N_3963,N_2582);
nand U9650 (N_9650,N_1762,N_714);
nor U9651 (N_9651,N_2530,N_3862);
nand U9652 (N_9652,N_1633,N_3197);
or U9653 (N_9653,N_1569,N_2940);
nand U9654 (N_9654,N_4480,N_952);
or U9655 (N_9655,N_386,N_3475);
and U9656 (N_9656,N_4917,N_3826);
and U9657 (N_9657,N_2475,N_2880);
or U9658 (N_9658,N_2345,N_1479);
and U9659 (N_9659,N_757,N_1526);
and U9660 (N_9660,N_2335,N_4232);
and U9661 (N_9661,N_385,N_748);
nand U9662 (N_9662,N_133,N_1569);
nand U9663 (N_9663,N_3217,N_3186);
and U9664 (N_9664,N_4927,N_563);
nor U9665 (N_9665,N_316,N_1104);
and U9666 (N_9666,N_1523,N_2734);
and U9667 (N_9667,N_4204,N_4607);
xnor U9668 (N_9668,N_1785,N_1603);
or U9669 (N_9669,N_2871,N_2275);
nand U9670 (N_9670,N_503,N_3786);
nor U9671 (N_9671,N_2135,N_2300);
or U9672 (N_9672,N_101,N_3546);
xnor U9673 (N_9673,N_4550,N_1966);
nor U9674 (N_9674,N_553,N_3477);
nor U9675 (N_9675,N_3195,N_2261);
nand U9676 (N_9676,N_25,N_2797);
or U9677 (N_9677,N_1461,N_4462);
nor U9678 (N_9678,N_4441,N_744);
nand U9679 (N_9679,N_2373,N_1840);
or U9680 (N_9680,N_1371,N_3981);
and U9681 (N_9681,N_4858,N_4886);
and U9682 (N_9682,N_4994,N_829);
nor U9683 (N_9683,N_2895,N_4689);
nor U9684 (N_9684,N_1209,N_1400);
or U9685 (N_9685,N_2923,N_1967);
nand U9686 (N_9686,N_2957,N_1914);
nor U9687 (N_9687,N_1612,N_3595);
and U9688 (N_9688,N_1293,N_1769);
and U9689 (N_9689,N_4790,N_2721);
nor U9690 (N_9690,N_4805,N_1019);
nand U9691 (N_9691,N_3694,N_327);
and U9692 (N_9692,N_3619,N_4034);
nand U9693 (N_9693,N_2314,N_25);
nor U9694 (N_9694,N_2404,N_3193);
and U9695 (N_9695,N_1227,N_534);
or U9696 (N_9696,N_4633,N_2309);
nand U9697 (N_9697,N_3953,N_1172);
nand U9698 (N_9698,N_856,N_3181);
nand U9699 (N_9699,N_4099,N_4321);
nand U9700 (N_9700,N_3677,N_4277);
nand U9701 (N_9701,N_4844,N_3683);
nand U9702 (N_9702,N_58,N_1014);
and U9703 (N_9703,N_3456,N_3449);
nand U9704 (N_9704,N_4341,N_1763);
nand U9705 (N_9705,N_1095,N_1574);
nor U9706 (N_9706,N_2911,N_1072);
and U9707 (N_9707,N_324,N_1415);
or U9708 (N_9708,N_2003,N_2550);
nor U9709 (N_9709,N_51,N_1994);
nand U9710 (N_9710,N_3260,N_3000);
nand U9711 (N_9711,N_4746,N_4497);
nand U9712 (N_9712,N_3861,N_3047);
nand U9713 (N_9713,N_2809,N_2549);
nor U9714 (N_9714,N_2066,N_1464);
nor U9715 (N_9715,N_629,N_1277);
and U9716 (N_9716,N_4365,N_2242);
xnor U9717 (N_9717,N_2785,N_2160);
or U9718 (N_9718,N_4792,N_2746);
or U9719 (N_9719,N_736,N_3890);
and U9720 (N_9720,N_4567,N_2610);
and U9721 (N_9721,N_598,N_997);
and U9722 (N_9722,N_64,N_1164);
nand U9723 (N_9723,N_1499,N_2589);
and U9724 (N_9724,N_2991,N_942);
and U9725 (N_9725,N_1298,N_3569);
nor U9726 (N_9726,N_4643,N_1030);
xor U9727 (N_9727,N_2932,N_1820);
or U9728 (N_9728,N_4897,N_3769);
nand U9729 (N_9729,N_2632,N_1274);
nand U9730 (N_9730,N_664,N_237);
nand U9731 (N_9731,N_3927,N_1893);
and U9732 (N_9732,N_4969,N_325);
nand U9733 (N_9733,N_3060,N_3842);
nand U9734 (N_9734,N_4392,N_2763);
nor U9735 (N_9735,N_4058,N_4661);
or U9736 (N_9736,N_427,N_4393);
nand U9737 (N_9737,N_2951,N_1210);
or U9738 (N_9738,N_4848,N_2791);
nor U9739 (N_9739,N_3488,N_3100);
nor U9740 (N_9740,N_3810,N_1588);
and U9741 (N_9741,N_1095,N_3324);
and U9742 (N_9742,N_298,N_1125);
nor U9743 (N_9743,N_891,N_2683);
xnor U9744 (N_9744,N_784,N_2554);
and U9745 (N_9745,N_2930,N_4607);
and U9746 (N_9746,N_245,N_1213);
nor U9747 (N_9747,N_1908,N_2854);
and U9748 (N_9748,N_4885,N_2076);
nor U9749 (N_9749,N_1254,N_228);
nand U9750 (N_9750,N_3768,N_4772);
or U9751 (N_9751,N_897,N_3055);
and U9752 (N_9752,N_425,N_4478);
and U9753 (N_9753,N_2618,N_3553);
or U9754 (N_9754,N_2861,N_53);
nor U9755 (N_9755,N_4438,N_1534);
xor U9756 (N_9756,N_2663,N_1870);
or U9757 (N_9757,N_2842,N_532);
or U9758 (N_9758,N_4225,N_4620);
or U9759 (N_9759,N_4113,N_3162);
nand U9760 (N_9760,N_1440,N_2295);
and U9761 (N_9761,N_691,N_3215);
nor U9762 (N_9762,N_4817,N_623);
nand U9763 (N_9763,N_2738,N_4734);
nand U9764 (N_9764,N_2523,N_1810);
or U9765 (N_9765,N_1180,N_918);
or U9766 (N_9766,N_4151,N_1742);
xor U9767 (N_9767,N_3443,N_195);
nand U9768 (N_9768,N_2833,N_462);
nand U9769 (N_9769,N_1695,N_1738);
and U9770 (N_9770,N_2483,N_3355);
nand U9771 (N_9771,N_3380,N_1065);
and U9772 (N_9772,N_2368,N_368);
nor U9773 (N_9773,N_4074,N_2246);
or U9774 (N_9774,N_246,N_4505);
xor U9775 (N_9775,N_416,N_4323);
or U9776 (N_9776,N_3198,N_2373);
and U9777 (N_9777,N_2005,N_3464);
nand U9778 (N_9778,N_1475,N_2877);
or U9779 (N_9779,N_3768,N_3789);
xor U9780 (N_9780,N_1270,N_4889);
or U9781 (N_9781,N_3866,N_3436);
nand U9782 (N_9782,N_618,N_1872);
or U9783 (N_9783,N_4413,N_4776);
and U9784 (N_9784,N_4311,N_2308);
nor U9785 (N_9785,N_2230,N_179);
and U9786 (N_9786,N_3911,N_3466);
and U9787 (N_9787,N_4778,N_4132);
or U9788 (N_9788,N_4571,N_660);
nor U9789 (N_9789,N_597,N_2997);
or U9790 (N_9790,N_3179,N_3711);
nor U9791 (N_9791,N_4545,N_1618);
and U9792 (N_9792,N_2351,N_4298);
or U9793 (N_9793,N_4053,N_1676);
nand U9794 (N_9794,N_912,N_4336);
or U9795 (N_9795,N_3105,N_2043);
xor U9796 (N_9796,N_3956,N_4577);
nand U9797 (N_9797,N_601,N_362);
nand U9798 (N_9798,N_3605,N_3149);
nand U9799 (N_9799,N_2065,N_3368);
or U9800 (N_9800,N_2117,N_2813);
or U9801 (N_9801,N_2906,N_2565);
and U9802 (N_9802,N_804,N_3110);
and U9803 (N_9803,N_3101,N_4950);
xnor U9804 (N_9804,N_2279,N_2928);
xor U9805 (N_9805,N_3630,N_3203);
and U9806 (N_9806,N_3093,N_4827);
and U9807 (N_9807,N_1487,N_3841);
or U9808 (N_9808,N_1496,N_3390);
nand U9809 (N_9809,N_3450,N_1963);
or U9810 (N_9810,N_3721,N_3633);
or U9811 (N_9811,N_3418,N_4444);
nor U9812 (N_9812,N_1877,N_2027);
nand U9813 (N_9813,N_3126,N_4424);
nor U9814 (N_9814,N_2317,N_4550);
and U9815 (N_9815,N_2869,N_328);
nor U9816 (N_9816,N_1192,N_208);
nand U9817 (N_9817,N_2687,N_507);
and U9818 (N_9818,N_3569,N_1156);
and U9819 (N_9819,N_776,N_230);
nand U9820 (N_9820,N_2768,N_3822);
nand U9821 (N_9821,N_2070,N_4991);
or U9822 (N_9822,N_3887,N_3294);
nand U9823 (N_9823,N_3635,N_4796);
or U9824 (N_9824,N_2078,N_4343);
nor U9825 (N_9825,N_842,N_2014);
nor U9826 (N_9826,N_1624,N_2195);
or U9827 (N_9827,N_1740,N_3529);
nand U9828 (N_9828,N_564,N_3063);
nor U9829 (N_9829,N_4025,N_1501);
nand U9830 (N_9830,N_3910,N_2208);
nor U9831 (N_9831,N_2458,N_2000);
nand U9832 (N_9832,N_1911,N_3485);
nand U9833 (N_9833,N_4689,N_4945);
nand U9834 (N_9834,N_4356,N_2682);
xnor U9835 (N_9835,N_1652,N_4573);
nor U9836 (N_9836,N_3950,N_3981);
or U9837 (N_9837,N_1628,N_321);
and U9838 (N_9838,N_446,N_1132);
nor U9839 (N_9839,N_164,N_1607);
or U9840 (N_9840,N_4893,N_4498);
or U9841 (N_9841,N_4663,N_702);
and U9842 (N_9842,N_2507,N_2160);
nand U9843 (N_9843,N_876,N_4498);
nor U9844 (N_9844,N_1517,N_3553);
nor U9845 (N_9845,N_3314,N_39);
or U9846 (N_9846,N_3152,N_723);
or U9847 (N_9847,N_4859,N_2729);
or U9848 (N_9848,N_533,N_1397);
or U9849 (N_9849,N_840,N_2881);
nor U9850 (N_9850,N_4201,N_2096);
nand U9851 (N_9851,N_1407,N_1798);
and U9852 (N_9852,N_449,N_3352);
nor U9853 (N_9853,N_543,N_3073);
nand U9854 (N_9854,N_740,N_2368);
nand U9855 (N_9855,N_3176,N_4325);
or U9856 (N_9856,N_1076,N_3018);
nor U9857 (N_9857,N_3579,N_150);
or U9858 (N_9858,N_3128,N_2987);
or U9859 (N_9859,N_2184,N_916);
nor U9860 (N_9860,N_2273,N_1016);
nor U9861 (N_9861,N_4832,N_3660);
nand U9862 (N_9862,N_2633,N_3213);
xnor U9863 (N_9863,N_1563,N_59);
or U9864 (N_9864,N_3095,N_838);
nand U9865 (N_9865,N_3884,N_3185);
nand U9866 (N_9866,N_2648,N_3315);
or U9867 (N_9867,N_3357,N_1695);
xor U9868 (N_9868,N_4240,N_1402);
nor U9869 (N_9869,N_2696,N_2956);
or U9870 (N_9870,N_3459,N_3100);
xor U9871 (N_9871,N_3573,N_4234);
nand U9872 (N_9872,N_4384,N_1630);
nand U9873 (N_9873,N_2672,N_4199);
nand U9874 (N_9874,N_3732,N_4479);
or U9875 (N_9875,N_714,N_1818);
and U9876 (N_9876,N_4952,N_1629);
or U9877 (N_9877,N_3600,N_4985);
nor U9878 (N_9878,N_2116,N_3238);
xor U9879 (N_9879,N_1355,N_3484);
nand U9880 (N_9880,N_4014,N_3033);
nor U9881 (N_9881,N_4441,N_63);
nor U9882 (N_9882,N_55,N_1619);
and U9883 (N_9883,N_1781,N_445);
nor U9884 (N_9884,N_166,N_3591);
or U9885 (N_9885,N_1645,N_4433);
nand U9886 (N_9886,N_4267,N_3785);
or U9887 (N_9887,N_1841,N_1988);
xnor U9888 (N_9888,N_4143,N_220);
nand U9889 (N_9889,N_4746,N_3844);
or U9890 (N_9890,N_4144,N_2011);
nor U9891 (N_9891,N_4905,N_721);
and U9892 (N_9892,N_188,N_2420);
or U9893 (N_9893,N_4064,N_2118);
or U9894 (N_9894,N_2119,N_3330);
and U9895 (N_9895,N_2585,N_3649);
nor U9896 (N_9896,N_2833,N_4186);
or U9897 (N_9897,N_2563,N_1858);
nand U9898 (N_9898,N_2232,N_704);
or U9899 (N_9899,N_2059,N_751);
and U9900 (N_9900,N_3162,N_603);
nor U9901 (N_9901,N_2505,N_3909);
and U9902 (N_9902,N_1935,N_3160);
or U9903 (N_9903,N_268,N_3840);
xor U9904 (N_9904,N_1984,N_3586);
and U9905 (N_9905,N_609,N_1220);
and U9906 (N_9906,N_2821,N_1953);
and U9907 (N_9907,N_4799,N_2613);
xnor U9908 (N_9908,N_1743,N_1785);
xor U9909 (N_9909,N_2239,N_763);
and U9910 (N_9910,N_4238,N_2833);
or U9911 (N_9911,N_3180,N_1245);
nand U9912 (N_9912,N_1132,N_4629);
or U9913 (N_9913,N_4455,N_2443);
nand U9914 (N_9914,N_3110,N_80);
nand U9915 (N_9915,N_4607,N_2615);
nand U9916 (N_9916,N_1130,N_4891);
or U9917 (N_9917,N_2251,N_168);
and U9918 (N_9918,N_3477,N_1373);
nor U9919 (N_9919,N_4033,N_1288);
nand U9920 (N_9920,N_2328,N_4093);
or U9921 (N_9921,N_1314,N_1174);
and U9922 (N_9922,N_1305,N_1241);
nor U9923 (N_9923,N_2505,N_2869);
xnor U9924 (N_9924,N_1782,N_1679);
and U9925 (N_9925,N_1980,N_2700);
nand U9926 (N_9926,N_72,N_630);
or U9927 (N_9927,N_358,N_39);
or U9928 (N_9928,N_120,N_4983);
nor U9929 (N_9929,N_3958,N_152);
and U9930 (N_9930,N_2325,N_675);
and U9931 (N_9931,N_1920,N_1443);
nor U9932 (N_9932,N_4970,N_4099);
and U9933 (N_9933,N_2394,N_200);
or U9934 (N_9934,N_3527,N_1953);
or U9935 (N_9935,N_423,N_1456);
xnor U9936 (N_9936,N_2085,N_3125);
nand U9937 (N_9937,N_1806,N_994);
xnor U9938 (N_9938,N_4242,N_228);
nor U9939 (N_9939,N_4508,N_4378);
and U9940 (N_9940,N_3963,N_2651);
nor U9941 (N_9941,N_913,N_4075);
or U9942 (N_9942,N_309,N_1851);
nor U9943 (N_9943,N_61,N_4789);
nand U9944 (N_9944,N_635,N_3727);
nand U9945 (N_9945,N_4170,N_4329);
nand U9946 (N_9946,N_3086,N_3105);
nor U9947 (N_9947,N_4940,N_2213);
xor U9948 (N_9948,N_1025,N_4060);
xor U9949 (N_9949,N_459,N_4197);
nor U9950 (N_9950,N_3353,N_2979);
or U9951 (N_9951,N_2608,N_3338);
xor U9952 (N_9952,N_3172,N_171);
and U9953 (N_9953,N_815,N_2529);
or U9954 (N_9954,N_799,N_3800);
or U9955 (N_9955,N_425,N_2441);
nor U9956 (N_9956,N_1822,N_706);
nand U9957 (N_9957,N_2496,N_3860);
nor U9958 (N_9958,N_2307,N_4320);
nor U9959 (N_9959,N_2709,N_2403);
nand U9960 (N_9960,N_4693,N_1876);
or U9961 (N_9961,N_4413,N_4885);
and U9962 (N_9962,N_520,N_1733);
or U9963 (N_9963,N_4994,N_4930);
nand U9964 (N_9964,N_2358,N_2368);
nand U9965 (N_9965,N_478,N_2974);
or U9966 (N_9966,N_3508,N_679);
nand U9967 (N_9967,N_1942,N_2933);
nand U9968 (N_9968,N_3379,N_3686);
xor U9969 (N_9969,N_3870,N_1075);
xnor U9970 (N_9970,N_1344,N_998);
and U9971 (N_9971,N_3763,N_1583);
xnor U9972 (N_9972,N_3391,N_4847);
or U9973 (N_9973,N_2108,N_1023);
nand U9974 (N_9974,N_1859,N_2969);
nand U9975 (N_9975,N_3729,N_4367);
nand U9976 (N_9976,N_4339,N_3851);
nor U9977 (N_9977,N_1737,N_1099);
and U9978 (N_9978,N_3336,N_3600);
nand U9979 (N_9979,N_3598,N_171);
nor U9980 (N_9980,N_800,N_3643);
or U9981 (N_9981,N_4561,N_2701);
nand U9982 (N_9982,N_1317,N_4285);
nor U9983 (N_9983,N_4599,N_2073);
nand U9984 (N_9984,N_3905,N_3467);
xor U9985 (N_9985,N_1399,N_2073);
and U9986 (N_9986,N_4082,N_1777);
nand U9987 (N_9987,N_4416,N_3405);
and U9988 (N_9988,N_448,N_1676);
nor U9989 (N_9989,N_1761,N_560);
and U9990 (N_9990,N_3574,N_1930);
nor U9991 (N_9991,N_56,N_2295);
nand U9992 (N_9992,N_1656,N_2584);
nand U9993 (N_9993,N_1630,N_2650);
or U9994 (N_9994,N_2730,N_3162);
nor U9995 (N_9995,N_3122,N_4477);
and U9996 (N_9996,N_3100,N_4853);
or U9997 (N_9997,N_3994,N_1698);
xor U9998 (N_9998,N_1933,N_3747);
and U9999 (N_9999,N_888,N_1033);
nand U10000 (N_10000,N_9816,N_7093);
xnor U10001 (N_10001,N_6100,N_9082);
nand U10002 (N_10002,N_5756,N_5243);
and U10003 (N_10003,N_6932,N_8743);
and U10004 (N_10004,N_7412,N_9076);
nor U10005 (N_10005,N_9103,N_9129);
xnor U10006 (N_10006,N_8929,N_8609);
nand U10007 (N_10007,N_9712,N_9568);
and U10008 (N_10008,N_5069,N_5609);
and U10009 (N_10009,N_5809,N_5789);
nand U10010 (N_10010,N_7354,N_5320);
and U10011 (N_10011,N_9518,N_7702);
xor U10012 (N_10012,N_7459,N_8313);
nor U10013 (N_10013,N_5373,N_7888);
nor U10014 (N_10014,N_8548,N_6589);
nand U10015 (N_10015,N_7554,N_9771);
and U10016 (N_10016,N_5009,N_8871);
or U10017 (N_10017,N_8889,N_8299);
or U10018 (N_10018,N_8979,N_7697);
nor U10019 (N_10019,N_5084,N_8566);
xor U10020 (N_10020,N_8171,N_9349);
and U10021 (N_10021,N_5890,N_8188);
nand U10022 (N_10022,N_7883,N_9921);
nor U10023 (N_10023,N_5829,N_6054);
or U10024 (N_10024,N_7772,N_8553);
nand U10025 (N_10025,N_9448,N_7581);
nand U10026 (N_10026,N_8995,N_7311);
or U10027 (N_10027,N_8174,N_8868);
nand U10028 (N_10028,N_8404,N_5448);
or U10029 (N_10029,N_9096,N_7935);
and U10030 (N_10030,N_7216,N_5112);
and U10031 (N_10031,N_5331,N_9228);
nor U10032 (N_10032,N_6082,N_9376);
and U10033 (N_10033,N_9273,N_5912);
nand U10034 (N_10034,N_8410,N_9538);
and U10035 (N_10035,N_7503,N_8734);
and U10036 (N_10036,N_8739,N_8006);
nor U10037 (N_10037,N_9791,N_8499);
xor U10038 (N_10038,N_8426,N_8133);
or U10039 (N_10039,N_5173,N_6035);
xor U10040 (N_10040,N_8760,N_7083);
or U10041 (N_10041,N_8844,N_5903);
xor U10042 (N_10042,N_6440,N_9268);
xor U10043 (N_10043,N_5405,N_7975);
nand U10044 (N_10044,N_8418,N_7550);
or U10045 (N_10045,N_9969,N_5509);
nand U10046 (N_10046,N_7568,N_6816);
nor U10047 (N_10047,N_9853,N_9405);
or U10048 (N_10048,N_9209,N_7079);
and U10049 (N_10049,N_5910,N_7687);
nor U10050 (N_10050,N_8272,N_9776);
and U10051 (N_10051,N_9549,N_8789);
xor U10052 (N_10052,N_8998,N_8143);
and U10053 (N_10053,N_8906,N_8054);
and U10054 (N_10054,N_7390,N_7191);
xor U10055 (N_10055,N_6957,N_9399);
or U10056 (N_10056,N_5653,N_6750);
nand U10057 (N_10057,N_7853,N_7054);
and U10058 (N_10058,N_7649,N_8668);
nor U10059 (N_10059,N_9580,N_5929);
and U10060 (N_10060,N_8990,N_9711);
or U10061 (N_10061,N_8599,N_5301);
and U10062 (N_10062,N_8819,N_7743);
nand U10063 (N_10063,N_6926,N_9948);
nor U10064 (N_10064,N_9848,N_6254);
or U10065 (N_10065,N_7086,N_9641);
nand U10066 (N_10066,N_7954,N_6064);
nor U10067 (N_10067,N_6187,N_5453);
nor U10068 (N_10068,N_8126,N_9383);
and U10069 (N_10069,N_7184,N_6891);
nand U10070 (N_10070,N_7931,N_6508);
or U10071 (N_10071,N_8015,N_7317);
nor U10072 (N_10072,N_6296,N_8616);
and U10073 (N_10073,N_8170,N_5853);
or U10074 (N_10074,N_6101,N_7969);
nor U10075 (N_10075,N_7933,N_8047);
nor U10076 (N_10076,N_7343,N_6734);
nand U10077 (N_10077,N_7410,N_9663);
nor U10078 (N_10078,N_7472,N_6320);
nand U10079 (N_10079,N_7283,N_9695);
nand U10080 (N_10080,N_8646,N_5242);
and U10081 (N_10081,N_7721,N_8247);
nor U10082 (N_10082,N_9566,N_8385);
or U10083 (N_10083,N_5870,N_5549);
or U10084 (N_10084,N_6940,N_9840);
or U10085 (N_10085,N_9724,N_6553);
xor U10086 (N_10086,N_5234,N_6302);
and U10087 (N_10087,N_9019,N_8241);
nor U10088 (N_10088,N_9424,N_5891);
xor U10089 (N_10089,N_9253,N_8339);
nand U10090 (N_10090,N_8594,N_5134);
nor U10091 (N_10091,N_5877,N_8664);
and U10092 (N_10092,N_5526,N_5698);
and U10093 (N_10093,N_5452,N_5334);
or U10094 (N_10094,N_7557,N_8136);
nand U10095 (N_10095,N_8970,N_9835);
or U10096 (N_10096,N_6546,N_9151);
nor U10097 (N_10097,N_8628,N_5458);
and U10098 (N_10098,N_6601,N_8758);
or U10099 (N_10099,N_9279,N_5149);
nor U10100 (N_10100,N_8084,N_6586);
nor U10101 (N_10101,N_8211,N_5863);
nand U10102 (N_10102,N_7504,N_6293);
or U10103 (N_10103,N_6216,N_9583);
nor U10104 (N_10104,N_6407,N_8693);
nand U10105 (N_10105,N_6909,N_6885);
xor U10106 (N_10106,N_5236,N_8269);
and U10107 (N_10107,N_7715,N_5446);
and U10108 (N_10108,N_7270,N_9084);
and U10109 (N_10109,N_9824,N_6638);
nor U10110 (N_10110,N_9673,N_8828);
nor U10111 (N_10111,N_6418,N_5090);
nor U10112 (N_10112,N_9274,N_6262);
or U10113 (N_10113,N_5239,N_5318);
or U10114 (N_10114,N_9602,N_6146);
or U10115 (N_10115,N_6286,N_8468);
nand U10116 (N_10116,N_7780,N_7261);
xnor U10117 (N_10117,N_6900,N_8737);
and U10118 (N_10118,N_5374,N_5433);
or U10119 (N_10119,N_7259,N_6132);
and U10120 (N_10120,N_6730,N_6720);
or U10121 (N_10121,N_9831,N_6676);
nor U10122 (N_10122,N_5013,N_8331);
and U10123 (N_10123,N_7921,N_5971);
nand U10124 (N_10124,N_6960,N_9302);
nor U10125 (N_10125,N_7910,N_9558);
nor U10126 (N_10126,N_8782,N_5407);
xor U10127 (N_10127,N_7169,N_5203);
or U10128 (N_10128,N_9978,N_9511);
and U10129 (N_10129,N_7861,N_6121);
xor U10130 (N_10130,N_6191,N_9595);
nor U10131 (N_10131,N_9856,N_6614);
and U10132 (N_10132,N_8402,N_8552);
or U10133 (N_10133,N_5425,N_8569);
or U10134 (N_10134,N_6039,N_7531);
and U10135 (N_10135,N_5854,N_5831);
or U10136 (N_10136,N_5582,N_5488);
or U10137 (N_10137,N_5668,N_8109);
or U10138 (N_10138,N_5873,N_8812);
nor U10139 (N_10139,N_6085,N_9254);
and U10140 (N_10140,N_5628,N_8381);
nor U10141 (N_10141,N_5057,N_7811);
xor U10142 (N_10142,N_5985,N_7075);
nand U10143 (N_10143,N_6092,N_7438);
and U10144 (N_10144,N_6069,N_6571);
nand U10145 (N_10145,N_6768,N_7549);
nor U10146 (N_10146,N_9325,N_7344);
nor U10147 (N_10147,N_6313,N_6918);
nor U10148 (N_10148,N_8715,N_9564);
nand U10149 (N_10149,N_9582,N_6860);
and U10150 (N_10150,N_5945,N_9265);
nand U10151 (N_10151,N_8258,N_5720);
and U10152 (N_10152,N_7378,N_5839);
nor U10153 (N_10153,N_5387,N_6065);
nand U10154 (N_10154,N_9839,N_9038);
xnor U10155 (N_10155,N_8546,N_6465);
and U10156 (N_10156,N_7767,N_8625);
and U10157 (N_10157,N_6139,N_6914);
nor U10158 (N_10158,N_6122,N_6236);
nor U10159 (N_10159,N_7355,N_9515);
nor U10160 (N_10160,N_8669,N_7451);
nor U10161 (N_10161,N_9726,N_6127);
or U10162 (N_10162,N_6387,N_8038);
nand U10163 (N_10163,N_7039,N_9161);
nor U10164 (N_10164,N_6003,N_7489);
or U10165 (N_10165,N_7372,N_7116);
and U10166 (N_10166,N_5753,N_7092);
nand U10167 (N_10167,N_9144,N_8924);
and U10168 (N_10168,N_6812,N_5219);
and U10169 (N_10169,N_5798,N_5467);
xnor U10170 (N_10170,N_6801,N_5792);
or U10171 (N_10171,N_9211,N_7685);
xor U10172 (N_10172,N_8318,N_9529);
nand U10173 (N_10173,N_6607,N_6290);
nand U10174 (N_10174,N_6613,N_7959);
nor U10175 (N_10175,N_6698,N_9427);
nand U10176 (N_10176,N_9772,N_7681);
nor U10177 (N_10177,N_6813,N_8017);
xnor U10178 (N_10178,N_6836,N_6389);
and U10179 (N_10179,N_6202,N_5313);
nor U10180 (N_10180,N_9474,N_9657);
nor U10181 (N_10181,N_6541,N_9392);
or U10182 (N_10182,N_7973,N_7467);
and U10183 (N_10183,N_9430,N_8479);
nand U10184 (N_10184,N_6351,N_8961);
or U10185 (N_10185,N_8037,N_7076);
xnor U10186 (N_10186,N_5815,N_8240);
or U10187 (N_10187,N_8667,N_5991);
or U10188 (N_10188,N_8769,N_6565);
xnor U10189 (N_10189,N_9075,N_7582);
or U10190 (N_10190,N_6797,N_7700);
nand U10191 (N_10191,N_7428,N_8721);
nor U10192 (N_10192,N_8985,N_7331);
nor U10193 (N_10193,N_8659,N_7166);
and U10194 (N_10194,N_5658,N_9309);
nor U10195 (N_10195,N_8325,N_5128);
xor U10196 (N_10196,N_7155,N_5516);
or U10197 (N_10197,N_8901,N_5520);
or U10198 (N_10198,N_5168,N_5258);
xnor U10199 (N_10199,N_7541,N_6526);
nand U10200 (N_10200,N_6584,N_8069);
xnor U10201 (N_10201,N_9944,N_7905);
and U10202 (N_10202,N_6946,N_8535);
or U10203 (N_10203,N_8373,N_9227);
and U10204 (N_10204,N_8401,N_5925);
and U10205 (N_10205,N_6442,N_6081);
or U10206 (N_10206,N_7358,N_8231);
nand U10207 (N_10207,N_8872,N_5772);
or U10208 (N_10208,N_6987,N_9607);
xor U10209 (N_10209,N_8053,N_8491);
and U10210 (N_10210,N_7104,N_9551);
nor U10211 (N_10211,N_5607,N_6350);
or U10212 (N_10212,N_8292,N_9562);
nand U10213 (N_10213,N_6412,N_9913);
or U10214 (N_10214,N_9468,N_5136);
or U10215 (N_10215,N_7591,N_8147);
nor U10216 (N_10216,N_6487,N_9823);
nand U10217 (N_10217,N_5814,N_6419);
xor U10218 (N_10218,N_7073,N_6563);
nand U10219 (N_10219,N_6431,N_7127);
xnor U10220 (N_10220,N_8526,N_6045);
and U10221 (N_10221,N_6503,N_8450);
nor U10222 (N_10222,N_5002,N_8248);
xnor U10223 (N_10223,N_7754,N_5486);
and U10224 (N_10224,N_9591,N_5762);
or U10225 (N_10225,N_9956,N_5087);
xnor U10226 (N_10226,N_9085,N_5916);
and U10227 (N_10227,N_5123,N_9787);
xor U10228 (N_10228,N_7015,N_5339);
and U10229 (N_10229,N_5924,N_5946);
nor U10230 (N_10230,N_8748,N_9132);
and U10231 (N_10231,N_5957,N_8504);
nand U10232 (N_10232,N_7096,N_5198);
xnor U10233 (N_10233,N_8026,N_6997);
nor U10234 (N_10234,N_6425,N_5269);
nor U10235 (N_10235,N_5282,N_5748);
nor U10236 (N_10236,N_9499,N_8003);
and U10237 (N_10237,N_5010,N_7555);
or U10238 (N_10238,N_7873,N_6790);
nand U10239 (N_10239,N_8608,N_7001);
nor U10240 (N_10240,N_7458,N_6219);
nand U10241 (N_10241,N_8962,N_6723);
nor U10242 (N_10242,N_5554,N_9188);
and U10243 (N_10243,N_6102,N_9109);
nand U10244 (N_10244,N_6029,N_8821);
nand U10245 (N_10245,N_7235,N_7768);
nand U10246 (N_10246,N_5113,N_5381);
or U10247 (N_10247,N_9644,N_6529);
nor U10248 (N_10248,N_7561,N_5190);
and U10249 (N_10249,N_5790,N_6361);
and U10250 (N_10250,N_9975,N_5708);
and U10251 (N_10251,N_5127,N_7932);
and U10252 (N_10252,N_8018,N_5583);
nand U10253 (N_10253,N_6748,N_8208);
or U10254 (N_10254,N_7643,N_7886);
nand U10255 (N_10255,N_8722,N_6809);
nand U10256 (N_10256,N_5743,N_5498);
xor U10257 (N_10257,N_6301,N_9322);
and U10258 (N_10258,N_7572,N_5182);
and U10259 (N_10259,N_6754,N_8550);
nor U10260 (N_10260,N_5451,N_9925);
or U10261 (N_10261,N_5600,N_7698);
xor U10262 (N_10262,N_5434,N_9395);
and U10263 (N_10263,N_8577,N_5353);
and U10264 (N_10264,N_7055,N_5968);
nand U10265 (N_10265,N_6845,N_5437);
nand U10266 (N_10266,N_6306,N_7341);
and U10267 (N_10267,N_9304,N_8119);
nand U10268 (N_10268,N_7318,N_9217);
nor U10269 (N_10269,N_5077,N_6319);
nor U10270 (N_10270,N_5962,N_7417);
xor U10271 (N_10271,N_5928,N_5521);
nand U10272 (N_10272,N_9862,N_8585);
nor U10273 (N_10273,N_5625,N_8931);
nor U10274 (N_10274,N_5245,N_8690);
nand U10275 (N_10275,N_7290,N_7110);
nor U10276 (N_10276,N_7774,N_9024);
nand U10277 (N_10277,N_7807,N_5580);
nor U10278 (N_10278,N_8319,N_9780);
nand U10279 (N_10279,N_9504,N_8864);
or U10280 (N_10280,N_8355,N_7406);
and U10281 (N_10281,N_8112,N_8266);
nor U10282 (N_10282,N_5895,N_5060);
nand U10283 (N_10283,N_9301,N_9110);
nor U10284 (N_10284,N_5771,N_9992);
and U10285 (N_10285,N_5726,N_6006);
and U10286 (N_10286,N_6327,N_7926);
and U10287 (N_10287,N_5428,N_8437);
nand U10288 (N_10288,N_7032,N_5881);
or U10289 (N_10289,N_8649,N_6760);
and U10290 (N_10290,N_6277,N_8744);
nor U10291 (N_10291,N_5291,N_8235);
nand U10292 (N_10292,N_8371,N_6846);
nor U10293 (N_10293,N_5704,N_5450);
xor U10294 (N_10294,N_7962,N_5055);
or U10295 (N_10295,N_7540,N_9714);
or U10296 (N_10296,N_9241,N_9857);
nor U10297 (N_10297,N_6835,N_6021);
or U10298 (N_10298,N_7564,N_7456);
and U10299 (N_10299,N_9521,N_9166);
nor U10300 (N_10300,N_9895,N_5862);
and U10301 (N_10301,N_9613,N_5931);
and U10302 (N_10302,N_9198,N_9652);
nand U10303 (N_10303,N_5175,N_5312);
and U10304 (N_10304,N_7018,N_6112);
or U10305 (N_10305,N_8536,N_8545);
nand U10306 (N_10306,N_5289,N_7966);
and U10307 (N_10307,N_6018,N_8455);
or U10308 (N_10308,N_9832,N_9370);
and U10309 (N_10309,N_9156,N_6126);
nand U10310 (N_10310,N_6381,N_6583);
nand U10311 (N_10311,N_5637,N_9509);
nor U10312 (N_10312,N_7469,N_7137);
or U10313 (N_10313,N_9017,N_8048);
and U10314 (N_10314,N_6189,N_5247);
and U10315 (N_10315,N_8592,N_5295);
or U10316 (N_10316,N_8799,N_6386);
or U10317 (N_10317,N_8651,N_9495);
and U10318 (N_10318,N_9805,N_6948);
and U10319 (N_10319,N_5052,N_9484);
and U10320 (N_10320,N_5211,N_9421);
xor U10321 (N_10321,N_5227,N_7193);
nor U10322 (N_10322,N_9725,N_6362);
nor U10323 (N_10323,N_8827,N_6086);
and U10324 (N_10324,N_9199,N_8116);
or U10325 (N_10325,N_9252,N_9500);
and U10326 (N_10326,N_6818,N_6604);
nor U10327 (N_10327,N_8670,N_9642);
or U10328 (N_10328,N_8596,N_8473);
and U10329 (N_10329,N_8315,N_8695);
nand U10330 (N_10330,N_5109,N_6096);
or U10331 (N_10331,N_9410,N_6598);
and U10332 (N_10332,N_6303,N_7402);
nor U10333 (N_10333,N_7695,N_5367);
nand U10334 (N_10334,N_9130,N_9362);
nand U10335 (N_10335,N_8014,N_9384);
and U10336 (N_10336,N_7844,N_6444);
nor U10337 (N_10337,N_6580,N_5755);
xor U10338 (N_10338,N_8542,N_6399);
or U10339 (N_10339,N_6806,N_9236);
and U10340 (N_10340,N_9574,N_7571);
or U10341 (N_10341,N_9890,N_9738);
and U10342 (N_10342,N_6706,N_5271);
nor U10343 (N_10343,N_9874,N_6378);
nor U10344 (N_10344,N_6176,N_6002);
nor U10345 (N_10345,N_8911,N_8959);
or U10346 (N_10346,N_9412,N_9194);
nand U10347 (N_10347,N_9232,N_8267);
and U10348 (N_10348,N_6624,N_6426);
or U10349 (N_10349,N_6186,N_7147);
xor U10350 (N_10350,N_8746,N_7426);
nor U10351 (N_10351,N_8790,N_9950);
or U10352 (N_10352,N_7219,N_8989);
nor U10353 (N_10353,N_5630,N_6304);
and U10354 (N_10354,N_6416,N_7822);
or U10355 (N_10355,N_7634,N_5575);
or U10356 (N_10356,N_7930,N_7411);
nand U10357 (N_10357,N_9258,N_7845);
nand U10358 (N_10358,N_9030,N_5076);
or U10359 (N_10359,N_9855,N_5610);
or U10360 (N_10360,N_7800,N_8102);
and U10361 (N_10361,N_9889,N_8368);
and U10362 (N_10362,N_9098,N_6068);
and U10363 (N_10363,N_8100,N_6751);
nor U10364 (N_10364,N_6198,N_6170);
nand U10365 (N_10365,N_9870,N_5368);
xor U10366 (N_10366,N_6849,N_5493);
or U10367 (N_10367,N_9250,N_7730);
and U10368 (N_10368,N_5484,N_9530);
and U10369 (N_10369,N_9207,N_8785);
or U10370 (N_10370,N_9417,N_7724);
or U10371 (N_10371,N_9523,N_5828);
nand U10372 (N_10372,N_7945,N_9702);
nand U10373 (N_10373,N_8277,N_6036);
or U10374 (N_10374,N_8205,N_6214);
or U10375 (N_10375,N_9981,N_6037);
and U10376 (N_10376,N_7128,N_6382);
nor U10377 (N_10377,N_6385,N_6937);
nor U10378 (N_10378,N_9987,N_9419);
nand U10379 (N_10379,N_6736,N_9080);
and U10380 (N_10380,N_7664,N_6903);
nor U10381 (N_10381,N_7090,N_6791);
or U10382 (N_10382,N_8753,N_7827);
and U10383 (N_10383,N_6853,N_8131);
nor U10384 (N_10384,N_7928,N_9897);
and U10385 (N_10385,N_7638,N_8190);
nand U10386 (N_10386,N_8149,N_8354);
nor U10387 (N_10387,N_7666,N_7474);
nor U10388 (N_10388,N_8486,N_5141);
nand U10389 (N_10389,N_6095,N_8696);
xor U10390 (N_10390,N_7713,N_6309);
or U10391 (N_10391,N_7661,N_7388);
or U10392 (N_10392,N_7894,N_8297);
or U10393 (N_10393,N_9037,N_7907);
nor U10394 (N_10394,N_9438,N_8028);
nand U10395 (N_10395,N_9413,N_9342);
and U10396 (N_10396,N_8412,N_7158);
nand U10397 (N_10397,N_7053,N_6994);
nor U10398 (N_10398,N_9270,N_7944);
and U10399 (N_10399,N_7338,N_9761);
and U10400 (N_10400,N_5431,N_9783);
nand U10401 (N_10401,N_5710,N_9542);
or U10402 (N_10402,N_6328,N_7925);
nand U10403 (N_10403,N_5321,N_7965);
xor U10404 (N_10404,N_6890,N_9074);
xnor U10405 (N_10405,N_6211,N_9540);
and U10406 (N_10406,N_7360,N_8791);
nand U10407 (N_10407,N_8859,N_6014);
or U10408 (N_10408,N_5820,N_5569);
or U10409 (N_10409,N_7512,N_9123);
nand U10410 (N_10410,N_7562,N_7627);
nor U10411 (N_10411,N_7632,N_9875);
nand U10412 (N_10412,N_9152,N_6422);
nor U10413 (N_10413,N_5018,N_7397);
xor U10414 (N_10414,N_9872,N_5274);
nor U10415 (N_10415,N_8389,N_6992);
xor U10416 (N_10416,N_7138,N_5517);
and U10417 (N_10417,N_9456,N_8367);
and U10418 (N_10418,N_7161,N_8180);
xnor U10419 (N_10419,N_8074,N_6915);
or U10420 (N_10420,N_8068,N_5465);
and U10421 (N_10421,N_8714,N_5365);
and U10422 (N_10422,N_6664,N_5598);
nand U10423 (N_10423,N_9418,N_7535);
and U10424 (N_10424,N_5307,N_7528);
nand U10425 (N_10425,N_9271,N_7764);
or U10426 (N_10426,N_5153,N_7887);
nor U10427 (N_10427,N_7080,N_8635);
or U10428 (N_10428,N_9356,N_8207);
or U10429 (N_10429,N_5608,N_6134);
or U10430 (N_10430,N_8615,N_9554);
nor U10431 (N_10431,N_6204,N_7301);
nor U10432 (N_10432,N_7674,N_9612);
nor U10433 (N_10433,N_6814,N_5218);
nor U10434 (N_10434,N_9293,N_6998);
nor U10435 (N_10435,N_9189,N_7679);
or U10436 (N_10436,N_5728,N_9192);
or U10437 (N_10437,N_5299,N_6648);
nand U10438 (N_10438,N_8614,N_7361);
nor U10439 (N_10439,N_6117,N_7113);
nor U10440 (N_10440,N_8786,N_6947);
nor U10441 (N_10441,N_8544,N_7992);
and U10442 (N_10442,N_5477,N_7726);
and U10443 (N_10443,N_6220,N_5260);
xor U10444 (N_10444,N_9317,N_8352);
nor U10445 (N_10445,N_9367,N_9905);
or U10446 (N_10446,N_8880,N_6356);
nand U10447 (N_10447,N_9621,N_6839);
nand U10448 (N_10448,N_5705,N_9454);
and U10449 (N_10449,N_8173,N_7289);
and U10450 (N_10450,N_8802,N_6475);
and U10451 (N_10451,N_5562,N_5277);
nand U10452 (N_10452,N_5143,N_9092);
nand U10453 (N_10453,N_9869,N_6898);
nor U10454 (N_10454,N_6344,N_8927);
or U10455 (N_10455,N_8528,N_9388);
and U10456 (N_10456,N_6680,N_8732);
nand U10457 (N_10457,N_6686,N_9296);
xor U10458 (N_10458,N_7985,N_7645);
nor U10459 (N_10459,N_8988,N_9137);
nor U10460 (N_10460,N_5308,N_5869);
xor U10461 (N_10461,N_5729,N_8971);
and U10462 (N_10462,N_6414,N_6902);
nand U10463 (N_10463,N_5588,N_6484);
nor U10464 (N_10464,N_5847,N_5177);
nor U10465 (N_10465,N_8862,N_6307);
and U10466 (N_10466,N_8547,N_5544);
and U10467 (N_10467,N_7002,N_6771);
or U10468 (N_10468,N_7040,N_8081);
xnor U10469 (N_10469,N_9860,N_5252);
and U10470 (N_10470,N_9704,N_5649);
and U10471 (N_10471,N_8953,N_8833);
nand U10472 (N_10472,N_8195,N_6912);
and U10473 (N_10473,N_7490,N_5797);
or U10474 (N_10474,N_7806,N_7563);
nand U10475 (N_10475,N_5116,N_9894);
nor U10476 (N_10476,N_7952,N_7502);
or U10477 (N_10477,N_9533,N_6201);
and U10478 (N_10478,N_6908,N_9105);
nand U10479 (N_10479,N_7971,N_5068);
xor U10480 (N_10480,N_8478,N_9881);
nand U10481 (N_10481,N_9692,N_9572);
nor U10482 (N_10482,N_7991,N_7972);
and U10483 (N_10483,N_6467,N_7956);
or U10484 (N_10484,N_5603,N_6089);
or U10485 (N_10485,N_9999,N_9575);
nand U10486 (N_10486,N_9608,N_7616);
nand U10487 (N_10487,N_9390,N_9269);
or U10488 (N_10488,N_7016,N_5511);
nor U10489 (N_10489,N_6959,N_7029);
nor U10490 (N_10490,N_8311,N_9078);
and U10491 (N_10491,N_5408,N_8870);
or U10492 (N_10492,N_7707,N_6490);
nor U10493 (N_10493,N_6148,N_6641);
nand U10494 (N_10494,N_5806,N_5265);
and U10495 (N_10495,N_5310,N_8808);
or U10496 (N_10496,N_7069,N_5686);
nand U10497 (N_10497,N_7478,N_6434);
and U10498 (N_10498,N_7941,N_7694);
or U10499 (N_10499,N_6007,N_7120);
or U10500 (N_10500,N_7457,N_7091);
or U10501 (N_10501,N_6501,N_7201);
and U10502 (N_10502,N_9041,N_6564);
nor U10503 (N_10503,N_5292,N_8698);
nor U10504 (N_10504,N_9527,N_9359);
nand U10505 (N_10505,N_9295,N_5541);
nand U10506 (N_10506,N_9878,N_9850);
nor U10507 (N_10507,N_8302,N_7651);
nand U10508 (N_10508,N_6973,N_5210);
xnor U10509 (N_10509,N_7683,N_7588);
nor U10510 (N_10510,N_5371,N_8905);
nand U10511 (N_10511,N_9486,N_9077);
nor U10512 (N_10512,N_9892,N_8013);
nor U10513 (N_10513,N_6534,N_9244);
nand U10514 (N_10514,N_5383,N_8836);
nand U10515 (N_10515,N_7794,N_6135);
nand U10516 (N_10516,N_6077,N_7878);
nand U10517 (N_10517,N_9962,N_7579);
nand U10518 (N_10518,N_7391,N_7297);
and U10519 (N_10519,N_5193,N_9808);
or U10520 (N_10520,N_7313,N_6572);
nand U10521 (N_10521,N_8025,N_8887);
or U10522 (N_10522,N_9798,N_5941);
and U10523 (N_10523,N_7984,N_7346);
nor U10524 (N_10524,N_7977,N_9093);
and U10525 (N_10525,N_9849,N_8497);
and U10526 (N_10526,N_6143,N_9010);
nand U10527 (N_10527,N_5398,N_6535);
nand U10528 (N_10528,N_6371,N_7074);
nor U10529 (N_10529,N_8898,N_7497);
nor U10530 (N_10530,N_8071,N_7114);
nor U10531 (N_10531,N_9520,N_6163);
nor U10532 (N_10532,N_8085,N_5978);
nand U10533 (N_10533,N_8096,N_7396);
nand U10534 (N_10534,N_7008,N_9736);
and U10535 (N_10535,N_5167,N_8772);
and U10536 (N_10536,N_8735,N_5871);
nor U10537 (N_10537,N_6376,N_8809);
xor U10538 (N_10538,N_9893,N_7639);
nor U10539 (N_10539,N_8169,N_7153);
nor U10540 (N_10540,N_5270,N_7159);
xor U10541 (N_10541,N_6567,N_8849);
nand U10542 (N_10542,N_8072,N_5952);
nand U10543 (N_10543,N_9147,N_8443);
or U10544 (N_10544,N_8640,N_6566);
xor U10545 (N_10545,N_6941,N_7696);
nand U10546 (N_10546,N_7937,N_7929);
or U10547 (N_10547,N_5413,N_8510);
and U10548 (N_10548,N_8919,N_5067);
nor U10549 (N_10549,N_6113,N_5059);
nand U10550 (N_10550,N_7659,N_9635);
nand U10551 (N_10551,N_8579,N_7842);
nand U10552 (N_10552,N_5352,N_7709);
nor U10553 (N_10553,N_6196,N_5161);
or U10554 (N_10554,N_5072,N_7433);
nor U10555 (N_10555,N_6780,N_6634);
nor U10556 (N_10556,N_5438,N_5640);
nor U10557 (N_10557,N_5326,N_5401);
and U10558 (N_10558,N_8941,N_7057);
or U10559 (N_10559,N_5133,N_6243);
nand U10560 (N_10560,N_7854,N_7386);
nor U10561 (N_10561,N_8604,N_9974);
xnor U10562 (N_10562,N_7779,N_6173);
and U10563 (N_10563,N_9541,N_8610);
nor U10564 (N_10564,N_6549,N_9289);
nand U10565 (N_10565,N_8306,N_5290);
or U10566 (N_10566,N_9623,N_9433);
nor U10567 (N_10567,N_6451,N_6488);
or U10568 (N_10568,N_9939,N_6928);
nand U10569 (N_10569,N_6958,N_5157);
nor U10570 (N_10570,N_8449,N_9158);
nor U10571 (N_10571,N_7961,N_6699);
and U10572 (N_10572,N_5154,N_5422);
and U10573 (N_10573,N_6391,N_9131);
or U10574 (N_10574,N_5444,N_9475);
or U10575 (N_10575,N_9073,N_7211);
and U10576 (N_10576,N_8958,N_6034);
or U10577 (N_10577,N_7792,N_7279);
nand U10578 (N_10578,N_9502,N_6969);
nor U10579 (N_10579,N_9665,N_8408);
nand U10580 (N_10580,N_9748,N_8834);
nor U10581 (N_10581,N_8111,N_5231);
nand U10582 (N_10582,N_8183,N_7742);
nand U10583 (N_10583,N_6636,N_5361);
and U10584 (N_10584,N_7162,N_9432);
nor U10585 (N_10585,N_8429,N_9004);
nand U10586 (N_10586,N_7825,N_6469);
or U10587 (N_10587,N_5694,N_7766);
xor U10588 (N_10588,N_7760,N_7475);
nand U10589 (N_10589,N_6347,N_6830);
or U10590 (N_10590,N_7189,N_8010);
and U10591 (N_10591,N_8107,N_7421);
xnor U10592 (N_10592,N_6160,N_7675);
or U10593 (N_10593,N_8908,N_9216);
and U10594 (N_10594,N_9949,N_8736);
nand U10595 (N_10595,N_8598,N_7552);
or U10596 (N_10596,N_8291,N_5769);
nor U10597 (N_10597,N_6588,N_6482);
nand U10598 (N_10598,N_5884,N_7601);
nand U10599 (N_10599,N_9380,N_6971);
xnor U10600 (N_10600,N_9995,N_6883);
and U10601 (N_10601,N_5605,N_6019);
nand U10602 (N_10602,N_6756,N_9238);
nor U10603 (N_10603,N_7846,N_8073);
or U10604 (N_10604,N_9843,N_7044);
nor U10605 (N_10605,N_9286,N_9032);
and U10606 (N_10606,N_6681,N_7030);
and U10607 (N_10607,N_8127,N_7109);
nor U10608 (N_10608,N_6510,N_9731);
and U10609 (N_10609,N_9054,N_5117);
nor U10610 (N_10610,N_5131,N_7819);
nor U10611 (N_10611,N_8032,N_6594);
nor U10612 (N_10612,N_5412,N_8249);
and U10613 (N_10613,N_6323,N_9007);
or U10614 (N_10614,N_6192,N_7277);
nor U10615 (N_10615,N_6114,N_9124);
and U10616 (N_10616,N_8718,N_9141);
or U10617 (N_10617,N_9510,N_5261);
nor U10618 (N_10618,N_6721,N_9754);
nand U10619 (N_10619,N_6024,N_8444);
nand U10620 (N_10620,N_6140,N_8848);
or U10621 (N_10621,N_5485,N_7367);
and U10622 (N_10622,N_8080,N_8850);
xor U10623 (N_10623,N_5447,N_7287);
xnor U10624 (N_10624,N_7583,N_9243);
nand U10625 (N_10625,N_5171,N_8515);
and U10626 (N_10626,N_5765,N_9072);
nor U10627 (N_10627,N_7547,N_8392);
and U10628 (N_10628,N_7132,N_7233);
nor U10629 (N_10629,N_8795,N_6632);
nor U10630 (N_10630,N_9774,N_5922);
and U10631 (N_10631,N_7847,N_8797);
and U10632 (N_10632,N_6322,N_5392);
and U10633 (N_10633,N_8245,N_6623);
nor U10634 (N_10634,N_7324,N_9128);
nand U10635 (N_10635,N_6931,N_9656);
nor U10636 (N_10636,N_8794,N_5028);
or U10637 (N_10637,N_7818,N_9437);
nor U10638 (N_10638,N_7786,N_5144);
or U10639 (N_10639,N_6506,N_6055);
or U10640 (N_10640,N_9750,N_8888);
nor U10641 (N_10641,N_8406,N_5824);
and U10642 (N_10642,N_8022,N_9833);
or U10643 (N_10643,N_9311,N_5859);
nor U10644 (N_10644,N_6674,N_5150);
xnor U10645 (N_10645,N_8595,N_8946);
or U10646 (N_10646,N_5779,N_9386);
or U10647 (N_10647,N_8529,N_9045);
nand U10648 (N_10648,N_5178,N_8132);
xor U10649 (N_10649,N_5920,N_8543);
nand U10650 (N_10650,N_6402,N_8326);
and U10651 (N_10651,N_7501,N_5561);
or U10652 (N_10652,N_8756,N_9264);
nor U10653 (N_10653,N_8275,N_9044);
and U10654 (N_10654,N_7867,N_9693);
or U10655 (N_10655,N_8083,N_5894);
nor U10656 (N_10656,N_8146,N_5539);
nand U10657 (N_10657,N_9220,N_8253);
nor U10658 (N_10658,N_9466,N_9852);
xnor U10659 (N_10659,N_9288,N_9299);
nand U10660 (N_10660,N_8694,N_9225);
nor U10661 (N_10661,N_8321,N_5897);
xnor U10662 (N_10662,N_8232,N_9361);
nor U10663 (N_10663,N_6504,N_9912);
nor U10664 (N_10664,N_9976,N_8984);
nand U10665 (N_10665,N_5118,N_5905);
nor U10666 (N_10666,N_7263,N_9947);
and U10667 (N_10667,N_9040,N_5146);
nand U10668 (N_10668,N_8021,N_5825);
nand U10669 (N_10669,N_7185,N_5278);
and U10670 (N_10670,N_7112,N_9633);
nand U10671 (N_10671,N_8879,N_9664);
nand U10672 (N_10672,N_7989,N_8035);
and U10673 (N_10673,N_9865,N_8964);
or U10674 (N_10674,N_6543,N_8829);
xnor U10675 (N_10675,N_8108,N_5403);
or U10676 (N_10676,N_7314,N_6866);
nand U10677 (N_10677,N_7187,N_7328);
and U10678 (N_10678,N_5723,N_9501);
nor U10679 (N_10679,N_5727,N_6728);
or U10680 (N_10680,N_6548,N_5702);
xnor U10681 (N_10681,N_9531,N_8697);
xnor U10682 (N_10682,N_6353,N_6716);
xor U10683 (N_10683,N_9119,N_7198);
nand U10684 (N_10684,N_9603,N_7558);
or U10685 (N_10685,N_9723,N_5502);
nand U10686 (N_10686,N_7167,N_7884);
nand U10687 (N_10687,N_5842,N_5455);
nor U10688 (N_10688,N_7123,N_6802);
and U10689 (N_10689,N_9360,N_9891);
and U10690 (N_10690,N_5606,N_6665);
nor U10691 (N_10691,N_7940,N_7711);
or U10692 (N_10692,N_9452,N_8986);
nand U10693 (N_10693,N_8106,N_8134);
and U10694 (N_10694,N_5416,N_5819);
nor U10695 (N_10695,N_5054,N_6683);
nor U10696 (N_10696,N_7269,N_9393);
or U10697 (N_10697,N_8597,N_7204);
nor U10698 (N_10698,N_9548,N_7890);
nand U10699 (N_10699,N_7609,N_8832);
nand U10700 (N_10700,N_6977,N_9300);
and U10701 (N_10701,N_9537,N_8914);
and U10702 (N_10702,N_6661,N_7493);
or U10703 (N_10703,N_6094,N_6174);
xor U10704 (N_10704,N_8145,N_6496);
nand U10705 (N_10705,N_9794,N_6975);
xnor U10706 (N_10706,N_9573,N_5759);
and U10707 (N_10707,N_6483,N_8061);
nand U10708 (N_10708,N_5103,N_9160);
nor U10709 (N_10709,N_6280,N_5943);
nand U10710 (N_10710,N_7785,N_7976);
nor U10711 (N_10711,N_6659,N_5025);
nor U10712 (N_10712,N_7869,N_9866);
nand U10713 (N_10713,N_9928,N_5773);
or U10714 (N_10714,N_6612,N_5314);
nor U10715 (N_10715,N_6349,N_9276);
and U10716 (N_10716,N_8441,N_8920);
nor U10717 (N_10717,N_6840,N_7446);
and U10718 (N_10718,N_9229,N_7843);
nand U10719 (N_10719,N_7070,N_8316);
and U10720 (N_10720,N_5385,N_6822);
nor U10721 (N_10721,N_8967,N_7917);
nand U10722 (N_10722,N_6287,N_8365);
and U10723 (N_10723,N_7140,N_9063);
nor U10724 (N_10724,N_9267,N_5657);
nor U10725 (N_10725,N_9068,N_9560);
nand U10726 (N_10726,N_5518,N_7596);
or U10727 (N_10727,N_6939,N_5639);
or U10728 (N_10728,N_9983,N_7735);
nand U10729 (N_10729,N_7594,N_5851);
or U10730 (N_10730,N_9666,N_6274);
and U10731 (N_10731,N_8161,N_7126);
xnor U10732 (N_10732,N_8843,N_7146);
nor U10733 (N_10733,N_7374,N_9436);
or U10734 (N_10734,N_7061,N_6710);
nand U10735 (N_10735,N_8448,N_9807);
and U10736 (N_10736,N_8439,N_7436);
and U10737 (N_10737,N_5937,N_5017);
nand U10738 (N_10738,N_8066,N_6251);
nor U10739 (N_10739,N_6722,N_8687);
nor U10740 (N_10740,N_9415,N_8166);
nand U10741 (N_10741,N_5276,N_7408);
nor U10742 (N_10742,N_6000,N_6053);
and U10743 (N_10743,N_5556,N_7300);
and U10744 (N_10744,N_9546,N_9451);
nor U10745 (N_10745,N_9698,N_5306);
or U10746 (N_10746,N_9001,N_6314);
nor U10747 (N_10747,N_5811,N_8379);
nand U10748 (N_10748,N_6460,N_8216);
and U10749 (N_10749,N_5800,N_6996);
and U10750 (N_10750,N_8593,N_6310);
or U10751 (N_10751,N_7282,N_6213);
nor U10752 (N_10752,N_9471,N_8830);
nand U10753 (N_10753,N_5725,N_8965);
and U10754 (N_10754,N_8630,N_8228);
and U10755 (N_10755,N_9793,N_6062);
nand U10756 (N_10756,N_8440,N_6887);
and U10757 (N_10757,N_6587,N_8467);
nand U10758 (N_10758,N_6787,N_8770);
and U10759 (N_10759,N_9721,N_9154);
or U10760 (N_10760,N_9021,N_5188);
nor U10761 (N_10761,N_5199,N_7577);
nor U10762 (N_10762,N_7570,N_5601);
nor U10763 (N_10763,N_8237,N_7337);
nor U10764 (N_10764,N_5006,N_7353);
nand U10765 (N_10765,N_5843,N_7848);
nand U10766 (N_10766,N_8673,N_8563);
and U10767 (N_10767,N_6249,N_6436);
nor U10768 (N_10768,N_9973,N_8360);
xor U10769 (N_10769,N_7942,N_9022);
nor U10770 (N_10770,N_6175,N_7516);
nand U10771 (N_10771,N_5885,N_7836);
nor U10772 (N_10772,N_6456,N_8298);
nor U10773 (N_10773,N_6794,N_8167);
xor U10774 (N_10774,N_5372,N_8672);
xor U10775 (N_10775,N_6530,N_9126);
xnor U10776 (N_10776,N_9447,N_5573);
nand U10777 (N_10777,N_9786,N_8817);
nor U10778 (N_10778,N_6983,N_8286);
nor U10779 (N_10779,N_6905,N_8749);
or U10780 (N_10780,N_8932,N_6498);
nor U10781 (N_10781,N_9543,N_6789);
or U10782 (N_10782,N_8088,N_8641);
nor U10783 (N_10783,N_7784,N_5156);
nor U10784 (N_10784,N_5246,N_8181);
xnor U10785 (N_10785,N_8280,N_6744);
nor U10786 (N_10786,N_6515,N_7765);
nand U10787 (N_10787,N_9887,N_5395);
or U10788 (N_10788,N_7407,N_8709);
or U10789 (N_10789,N_7913,N_6919);
nand U10790 (N_10790,N_5183,N_8397);
xnor U10791 (N_10791,N_8993,N_7835);
nand U10792 (N_10792,N_8784,N_7135);
or U10793 (N_10793,N_7859,N_7206);
or U10794 (N_10794,N_7881,N_8027);
xnor U10795 (N_10795,N_8561,N_6767);
nor U10796 (N_10796,N_5106,N_5040);
and U10797 (N_10797,N_8197,N_8556);
or U10798 (N_10798,N_6354,N_9775);
and U10799 (N_10799,N_7242,N_5932);
and U10800 (N_10800,N_8268,N_8689);
nand U10801 (N_10801,N_7855,N_9516);
or U10802 (N_10802,N_6863,N_5701);
nand U10803 (N_10803,N_8764,N_8781);
nand U10804 (N_10804,N_7463,N_8578);
nand U10805 (N_10805,N_5281,N_9218);
nand U10806 (N_10806,N_9819,N_9029);
or U10807 (N_10807,N_6245,N_9284);
nand U10808 (N_10808,N_6231,N_6647);
or U10809 (N_10809,N_9980,N_5241);
or U10810 (N_10810,N_9170,N_5550);
nor U10811 (N_10811,N_8224,N_8101);
nand U10812 (N_10812,N_5914,N_5338);
or U10813 (N_10813,N_8648,N_6011);
or U10814 (N_10814,N_7443,N_5195);
and U10815 (N_10815,N_6049,N_5342);
or U10816 (N_10816,N_5654,N_9937);
or U10817 (N_10817,N_5836,N_8363);
or U10818 (N_10818,N_7173,N_5648);
and U10819 (N_10819,N_6893,N_8179);
nor U10820 (N_10820,N_7626,N_7950);
nor U10821 (N_10821,N_8341,N_7415);
nor U10822 (N_10822,N_6740,N_9919);
nor U10823 (N_10823,N_7605,N_8184);
nand U10824 (N_10824,N_9260,N_8457);
or U10825 (N_10825,N_5351,N_6892);
or U10826 (N_10826,N_7005,N_7631);
or U10827 (N_10827,N_8420,N_7108);
and U10828 (N_10828,N_8692,N_9492);
xnor U10829 (N_10829,N_7693,N_9120);
or U10830 (N_10830,N_5039,N_5092);
nor U10831 (N_10831,N_8761,N_8831);
nor U10832 (N_10832,N_6075,N_6010);
and U10833 (N_10833,N_8928,N_8203);
nor U10834 (N_10834,N_8281,N_8317);
nor U10835 (N_10835,N_9000,N_5224);
nor U10836 (N_10836,N_6284,N_8532);
nand U10837 (N_10837,N_5463,N_7986);
and U10838 (N_10838,N_8686,N_5294);
nand U10839 (N_10839,N_9746,N_6582);
nor U10840 (N_10840,N_6074,N_9245);
or U10841 (N_10841,N_9180,N_5751);
and U10842 (N_10842,N_9836,N_9347);
or U10843 (N_10843,N_9247,N_7364);
nand U10844 (N_10844,N_7600,N_8092);
and U10845 (N_10845,N_5429,N_5022);
and U10846 (N_10846,N_9766,N_8329);
or U10847 (N_10847,N_8337,N_8779);
and U10848 (N_10848,N_7725,N_9321);
and U10849 (N_10849,N_5466,N_8621);
and U10850 (N_10850,N_9810,N_7274);
nand U10851 (N_10851,N_8803,N_8052);
nor U10852 (N_10852,N_9994,N_7419);
or U10853 (N_10853,N_6786,N_5745);
nor U10854 (N_10854,N_8255,N_8688);
and U10855 (N_10855,N_6334,N_9423);
xnor U10856 (N_10856,N_8727,N_9153);
nor U10857 (N_10857,N_5327,N_9348);
nand U10858 (N_10858,N_8157,N_9226);
nand U10859 (N_10859,N_8503,N_5747);
nor U10860 (N_10860,N_5397,N_6807);
nand U10861 (N_10861,N_9570,N_8075);
nor U10862 (N_10862,N_5414,N_5837);
nor U10863 (N_10863,N_7202,N_7276);
or U10864 (N_10864,N_7589,N_7755);
or U10865 (N_10865,N_7298,N_7874);
nand U10866 (N_10866,N_8707,N_5802);
xnor U10867 (N_10867,N_6499,N_6735);
or U10868 (N_10868,N_8343,N_8679);
nand U10869 (N_10869,N_5974,N_7007);
or U10870 (N_10870,N_7635,N_6441);
nand U10871 (N_10871,N_8278,N_9957);
xor U10872 (N_10872,N_7094,N_8422);
nand U10873 (N_10873,N_9749,N_5322);
nor U10874 (N_10874,N_6321,N_6610);
nor U10875 (N_10875,N_8141,N_9645);
nor U10876 (N_10876,N_6852,N_6083);
nand U10877 (N_10877,N_9728,N_5475);
nand U10878 (N_10878,N_5696,N_9363);
nor U10879 (N_10879,N_6554,N_8762);
or U10880 (N_10880,N_6657,N_6240);
nand U10881 (N_10881,N_8222,N_9960);
nor U10882 (N_10882,N_6758,N_6682);
or U10883 (N_10883,N_5459,N_8708);
or U10884 (N_10884,N_8699,N_6518);
nor U10885 (N_10885,N_9052,N_5122);
or U10886 (N_10886,N_8398,N_5990);
xor U10887 (N_10887,N_7088,N_6569);
xnor U10888 (N_10888,N_6662,N_7863);
and U10889 (N_10889,N_6238,N_9034);
nor U10890 (N_10890,N_7980,N_7383);
nand U10891 (N_10891,N_9959,N_7506);
nor U10892 (N_10892,N_6788,N_8533);
nand U10893 (N_10893,N_9394,N_5742);
and U10894 (N_10894,N_5362,N_7963);
nand U10895 (N_10895,N_7895,N_6763);
nor U10896 (N_10896,N_5963,N_6861);
nor U10897 (N_10897,N_7125,N_5615);
nor U10898 (N_10898,N_9478,N_8187);
nor U10899 (N_10899,N_6001,N_6252);
nand U10900 (N_10900,N_7323,N_9691);
nor U10901 (N_10901,N_6635,N_5186);
nand U10902 (N_10902,N_8506,N_9801);
nand U10903 (N_10903,N_6979,N_7427);
and U10904 (N_10904,N_9659,N_6463);
nor U10905 (N_10905,N_9778,N_5525);
xor U10906 (N_10906,N_6646,N_7542);
xor U10907 (N_10907,N_8130,N_7701);
or U10908 (N_10908,N_7936,N_5194);
nand U10909 (N_10909,N_5961,N_6981);
nor U10910 (N_10910,N_8427,N_6232);
and U10911 (N_10911,N_5947,N_5754);
or U10912 (N_10912,N_7011,N_9259);
or U10913 (N_10913,N_6410,N_7342);
nand U10914 (N_10914,N_7831,N_5302);
nand U10915 (N_10915,N_5064,N_7089);
xor U10916 (N_10916,N_9467,N_6087);
xnor U10917 (N_10917,N_5586,N_9669);
nand U10918 (N_10918,N_8947,N_9434);
and U10919 (N_10919,N_6390,N_6687);
or U10920 (N_10920,N_6764,N_8876);
and U10921 (N_10921,N_6491,N_5557);
or U10922 (N_10922,N_6154,N_9382);
nand U10923 (N_10923,N_8117,N_6162);
or U10924 (N_10924,N_9675,N_5827);
and U10925 (N_10925,N_9619,N_5468);
or U10926 (N_10926,N_8822,N_5911);
nor U10927 (N_10927,N_7769,N_9458);
and U10928 (N_10928,N_5402,N_9545);
or U10929 (N_10929,N_8629,N_9614);
or U10930 (N_10930,N_9316,N_7812);
and U10931 (N_10931,N_5441,N_9569);
or U10932 (N_10932,N_8745,N_9428);
or U10933 (N_10933,N_8178,N_7095);
nand U10934 (N_10934,N_9982,N_6241);
or U10935 (N_10935,N_5959,N_6913);
or U10936 (N_10936,N_7394,N_9996);
and U10937 (N_10937,N_8122,N_7841);
nand U10938 (N_10938,N_8223,N_6466);
nor U10939 (N_10939,N_5835,N_6650);
and U10940 (N_10940,N_5689,N_5531);
nor U10941 (N_10941,N_7336,N_9906);
or U10942 (N_10942,N_6408,N_9100);
nor U10943 (N_10943,N_8742,N_5528);
nand U10944 (N_10944,N_7924,N_5202);
xor U10945 (N_10945,N_9713,N_8518);
or U10946 (N_10946,N_5142,N_9353);
and U10947 (N_10947,N_7828,N_7487);
or U10948 (N_10948,N_9884,N_9535);
nand U10949 (N_10949,N_6639,N_5208);
or U10950 (N_10950,N_9674,N_9708);
or U10951 (N_10951,N_8229,N_8854);
nand U10952 (N_10952,N_8818,N_8846);
nor U10953 (N_10953,N_8041,N_9924);
nor U10954 (N_10954,N_7507,N_6370);
and U10955 (N_10955,N_9990,N_6145);
or U10956 (N_10956,N_5647,N_6897);
nor U10957 (N_10957,N_6020,N_7168);
and U10958 (N_10958,N_8378,N_9335);
or U10959 (N_10959,N_7144,N_9902);
nand U10960 (N_10960,N_7293,N_5691);
or U10961 (N_10961,N_5410,N_8530);
and U10962 (N_10962,N_8459,N_7160);
or U10963 (N_10963,N_6184,N_5003);
or U10964 (N_10964,N_8129,N_7536);
and U10965 (N_10965,N_7617,N_7533);
or U10966 (N_10966,N_5089,N_8644);
and U10967 (N_10967,N_7078,N_9277);
nand U10968 (N_10968,N_5591,N_6911);
nand U10969 (N_10969,N_8470,N_5540);
xor U10970 (N_10970,N_6991,N_6709);
and U10971 (N_10971,N_6631,N_7957);
or U10972 (N_10972,N_7889,N_8677);
xor U10973 (N_10973,N_6520,N_5172);
or U10974 (N_10974,N_9820,N_5255);
or U10975 (N_10975,N_5082,N_9941);
or U10976 (N_10976,N_5960,N_6430);
nor U10977 (N_10977,N_5776,N_7901);
and U10978 (N_10978,N_6358,N_8851);
or U10979 (N_10979,N_9159,N_7452);
nand U10980 (N_10980,N_9070,N_5159);
nor U10981 (N_10981,N_8638,N_6581);
nand U10982 (N_10982,N_9067,N_7770);
and U10983 (N_10983,N_7608,N_9697);
nand U10984 (N_10984,N_5676,N_7899);
and U10985 (N_10985,N_7657,N_9306);
or U10986 (N_10986,N_7920,N_5411);
nor U10987 (N_10987,N_7692,N_6921);
nor U10988 (N_10988,N_5101,N_6649);
nor U10989 (N_10989,N_6747,N_7710);
or U10990 (N_10990,N_5114,N_8265);
nand U10991 (N_10991,N_8517,N_6782);
nor U10992 (N_10992,N_9846,N_8816);
nand U10993 (N_10993,N_9681,N_8461);
xor U10994 (N_10994,N_7484,N_9667);
nand U10995 (N_10995,N_6283,N_7442);
or U10996 (N_10996,N_5663,N_5166);
nand U10997 (N_10997,N_6842,N_8218);
and U10998 (N_10998,N_7964,N_9926);
and U10999 (N_10999,N_8274,N_7911);
nor U11000 (N_11000,N_9710,N_6707);
nor U11001 (N_11001,N_5690,N_9167);
or U11002 (N_11002,N_9859,N_6963);
and U11003 (N_11003,N_9235,N_9911);
and U11004 (N_11004,N_5253,N_9028);
and U11005 (N_11005,N_5031,N_6765);
or U11006 (N_11006,N_5021,N_9668);
nor U11007 (N_11007,N_6239,N_5359);
or U11008 (N_11008,N_7480,N_5777);
and U11009 (N_11009,N_5799,N_5860);
nand U11010 (N_11010,N_9658,N_5120);
nand U11011 (N_11011,N_5213,N_5665);
nor U11012 (N_11012,N_9106,N_9525);
or U11013 (N_11013,N_6803,N_7244);
or U11014 (N_11014,N_7389,N_8680);
and U11015 (N_11015,N_5893,N_9768);
xnor U11016 (N_11016,N_7131,N_8903);
or U11017 (N_11017,N_6325,N_8865);
or U11018 (N_11018,N_7133,N_5670);
and U11019 (N_11019,N_7425,N_8271);
and U11020 (N_11020,N_6925,N_6076);
nor U11021 (N_11021,N_9720,N_9903);
nor U11022 (N_11022,N_7035,N_9181);
and U11023 (N_11023,N_9942,N_7066);
or U11024 (N_11024,N_6719,N_5563);
or U11025 (N_11025,N_5983,N_8307);
nand U11026 (N_11026,N_9867,N_6368);
nand U11027 (N_11027,N_7042,N_5718);
and U11028 (N_11028,N_5409,N_5571);
or U11029 (N_11029,N_9481,N_7714);
nand U11030 (N_11030,N_7580,N_6359);
nand U11031 (N_11031,N_6573,N_5987);
nand U11032 (N_11032,N_9047,N_9409);
nand U11033 (N_11033,N_7900,N_9931);
nor U11034 (N_11034,N_8226,N_7295);
nor U11035 (N_11035,N_5162,N_9814);
nor U11036 (N_11036,N_7860,N_6511);
xnor U11037 (N_11037,N_8560,N_8446);
and U11038 (N_11038,N_8650,N_7902);
or U11039 (N_11039,N_8717,N_7129);
nor U11040 (N_11040,N_5761,N_9627);
and U11041 (N_11041,N_9581,N_7130);
and U11042 (N_11042,N_9314,N_5681);
and U11043 (N_11043,N_5812,N_6169);
or U11044 (N_11044,N_6545,N_7320);
and U11045 (N_11045,N_7870,N_6729);
nand U11046 (N_11046,N_5145,N_8554);
or U11047 (N_11047,N_6403,N_5979);
and U11048 (N_11048,N_5669,N_9310);
nand U11049 (N_11049,N_5977,N_5048);
nor U11050 (N_11050,N_8040,N_8531);
and U11051 (N_11051,N_5311,N_9482);
and U11052 (N_11052,N_5305,N_7882);
nor U11053 (N_11053,N_7099,N_9373);
nor U11054 (N_11054,N_7392,N_5840);
and U11055 (N_11055,N_9145,N_6523);
and U11056 (N_11056,N_8949,N_7741);
or U11057 (N_11057,N_8434,N_7904);
or U11058 (N_11058,N_7302,N_6329);
and U11059 (N_11059,N_9490,N_7646);
or U11060 (N_11060,N_7225,N_7719);
or U11061 (N_11061,N_5581,N_5185);
or U11062 (N_11062,N_5578,N_9343);
nand U11063 (N_11063,N_6672,N_9135);
nand U11064 (N_11064,N_7496,N_9534);
xor U11065 (N_11065,N_7172,N_9491);
nand U11066 (N_11066,N_9125,N_7207);
nand U11067 (N_11067,N_5419,N_8777);
nand U11068 (N_11068,N_8907,N_5356);
and U11069 (N_11069,N_6105,N_7329);
and U11070 (N_11070,N_8121,N_9291);
nor U11071 (N_11071,N_8861,N_7934);
or U11072 (N_11072,N_5005,N_5316);
or U11073 (N_11073,N_9522,N_7031);
or U11074 (N_11074,N_8144,N_8007);
nor U11075 (N_11075,N_8873,N_5666);
nor U11076 (N_11076,N_6318,N_5491);
xnor U11077 (N_11077,N_8220,N_8555);
and U11078 (N_11078,N_5093,N_6966);
nor U11079 (N_11079,N_5232,N_8164);
nand U11080 (N_11080,N_9922,N_7737);
or U11081 (N_11081,N_9407,N_7995);
nand U11082 (N_11082,N_6478,N_5357);
and U11083 (N_11083,N_8881,N_8262);
nand U11084 (N_11084,N_7143,N_5248);
nand U11085 (N_11085,N_5073,N_6888);
nor U11086 (N_11086,N_6690,N_6363);
nor U11087 (N_11087,N_9963,N_5744);
nand U11088 (N_11088,N_8344,N_7654);
and U11089 (N_11089,N_8896,N_8647);
nor U11090 (N_11090,N_7602,N_9611);
xnor U11091 (N_11091,N_8125,N_7663);
nand U11092 (N_11092,N_7230,N_8662);
or U11093 (N_11093,N_6865,N_8740);
and U11094 (N_11094,N_7050,N_9606);
nor U11095 (N_11095,N_7179,N_8607);
xor U11096 (N_11096,N_9350,N_5456);
nor U11097 (N_11097,N_5215,N_5791);
and U11098 (N_11098,N_6298,N_7546);
nand U11099 (N_11099,N_5519,N_8838);
or U11100 (N_11100,N_5662,N_6942);
and U11101 (N_11101,N_6281,N_6628);
or U11102 (N_11102,N_5354,N_8574);
and U11103 (N_11103,N_6955,N_5908);
and U11104 (N_11104,N_6144,N_6536);
and U11105 (N_11105,N_7460,N_8845);
or U11106 (N_11106,N_9508,N_8997);
nand U11107 (N_11107,N_5560,N_8055);
and U11108 (N_11108,N_5546,N_8002);
nand U11109 (N_11109,N_7906,N_6429);
xor U11110 (N_11110,N_8921,N_8624);
and U11111 (N_11111,N_8619,N_5051);
or U11112 (N_11112,N_6964,N_8852);
or U11113 (N_11113,N_8089,N_6435);
and U11114 (N_11114,N_6933,N_8332);
or U11115 (N_11115,N_7947,N_5687);
or U11116 (N_11116,N_5333,N_9684);
or U11117 (N_11117,N_5489,N_7923);
nor U11118 (N_11118,N_6949,N_6671);
and U11119 (N_11119,N_6826,N_6660);
or U11120 (N_11120,N_9177,N_8155);
and U11121 (N_11121,N_6922,N_9179);
or U11122 (N_11122,N_6455,N_5079);
nand U11123 (N_11123,N_7509,N_7464);
and U11124 (N_11124,N_5782,N_8897);
or U11125 (N_11125,N_9777,N_5415);
and U11126 (N_11126,N_5505,N_8591);
nand U11127 (N_11127,N_8787,N_9561);
or U11128 (N_11128,N_9023,N_9339);
nand U11129 (N_11129,N_7020,N_7789);
or U11130 (N_11130,N_7208,N_6899);
and U11131 (N_11131,N_7864,N_5369);
xor U11132 (N_11132,N_6073,N_8357);
or U11133 (N_11133,N_6867,N_5872);
nor U11134 (N_11134,N_5345,N_6445);
nand U11135 (N_11135,N_9176,N_5834);
or U11136 (N_11136,N_7578,N_9812);
and U11137 (N_11137,N_5706,N_9909);
nand U11138 (N_11138,N_8939,N_9584);
xor U11139 (N_11139,N_5482,N_6080);
nand U11140 (N_11140,N_8703,N_9061);
nor U11141 (N_11141,N_9532,N_9201);
or U11142 (N_11142,N_6315,N_9112);
nor U11143 (N_11143,N_7599,N_9979);
nor U11144 (N_11144,N_6779,N_7517);
nand U11145 (N_11145,N_5346,N_5179);
or U11146 (N_11146,N_7087,N_8612);
nand U11147 (N_11147,N_8934,N_7850);
nor U11148 (N_11148,N_6259,N_5110);
and U11149 (N_11149,N_7064,N_9221);
xor U11150 (N_11150,N_6023,N_5000);
and U11151 (N_11151,N_7186,N_9958);
and U11152 (N_11152,N_9646,N_9555);
nor U11153 (N_11153,N_7325,N_9524);
or U11154 (N_11154,N_7665,N_8733);
or U11155 (N_11155,N_5918,N_7224);
xnor U11156 (N_11156,N_9686,N_5044);
xnor U11157 (N_11157,N_8290,N_6072);
or U11158 (N_11158,N_6265,N_8869);
nand U11159 (N_11159,N_9758,N_6316);
nand U11160 (N_11160,N_8631,N_8451);
nand U11161 (N_11161,N_7059,N_9512);
xnor U11162 (N_11162,N_7246,N_9307);
or U11163 (N_11163,N_9883,N_7544);
and U11164 (N_11164,N_5786,N_9813);
and U11165 (N_11165,N_6406,N_7647);
or U11166 (N_11166,N_6131,N_7217);
and U11167 (N_11167,N_8023,N_9283);
nor U11168 (N_11168,N_6823,N_5855);
or U11169 (N_11169,N_5443,N_9882);
nor U11170 (N_11170,N_5981,N_9055);
nor U11171 (N_11171,N_9709,N_9118);
nand U11172 (N_11172,N_5939,N_7453);
and U11173 (N_11173,N_6952,N_7538);
nand U11174 (N_11174,N_5651,N_8860);
nand U11175 (N_11175,N_8227,N_6851);
and U11176 (N_11176,N_5650,N_5135);
and U11177 (N_11177,N_6951,N_6551);
nand U11178 (N_11178,N_5442,N_6025);
or U11179 (N_11179,N_8551,N_8336);
nor U11180 (N_11180,N_5358,N_7520);
or U11181 (N_11181,N_7334,N_9031);
and U11182 (N_11182,N_7098,N_8282);
nor U11183 (N_11183,N_5976,N_6880);
or U11184 (N_11184,N_5216,N_7356);
or U11185 (N_11185,N_8700,N_8835);
nor U11186 (N_11186,N_7060,N_5907);
or U11187 (N_11187,N_5818,N_6984);
nand U11188 (N_11188,N_9257,N_6178);
and U11189 (N_11189,N_5364,N_8000);
nor U11190 (N_11190,N_9649,N_6528);
nor U11191 (N_11191,N_9971,N_5151);
and U11192 (N_11192,N_9039,N_8472);
nand U11193 (N_11193,N_5674,N_5348);
and U11194 (N_11194,N_7880,N_8388);
or U11195 (N_11195,N_7560,N_6016);
nor U11196 (N_11196,N_5917,N_8225);
xor U11197 (N_11197,N_8251,N_7327);
or U11198 (N_11198,N_6778,N_8485);
nand U11199 (N_11199,N_5643,N_9879);
nand U11200 (N_11200,N_5741,N_6181);
and U11201 (N_11201,N_5986,N_6770);
and U11202 (N_11202,N_8639,N_5204);
xor U11203 (N_11203,N_7518,N_9923);
or U11204 (N_11204,N_9435,N_8763);
or U11205 (N_11205,N_6048,N_9139);
and U11206 (N_11206,N_7802,N_9477);
and U11207 (N_11207,N_9416,N_9334);
or U11208 (N_11208,N_6828,N_9876);
nand U11209 (N_11209,N_8793,N_6878);
nand U11210 (N_11210,N_7382,N_7262);
nor U11211 (N_11211,N_5764,N_6542);
nand U11212 (N_11212,N_9332,N_7387);
nor U11213 (N_11213,N_6713,N_8951);
nand U11214 (N_11214,N_9345,N_7395);
nor U11215 (N_11215,N_8123,N_7072);
or U11216 (N_11216,N_8882,N_6104);
nor U11217 (N_11217,N_9797,N_8110);
nor U11218 (N_11218,N_6741,N_9058);
nor U11219 (N_11219,N_6856,N_7673);
nand U11220 (N_11220,N_5462,N_7592);
nand U11221 (N_11221,N_9717,N_5671);
and U11222 (N_11222,N_6275,N_5030);
nor U11223 (N_11223,N_7668,N_7773);
or U11224 (N_11224,N_6237,N_5548);
or U11225 (N_11225,N_5086,N_5487);
xnor U11226 (N_11226,N_7220,N_7033);
or U11227 (N_11227,N_8447,N_9965);
nand U11228 (N_11228,N_9800,N_9972);
nor U11229 (N_11229,N_9961,N_6834);
xnor U11230 (N_11230,N_8206,N_9751);
nand U11231 (N_11231,N_5636,N_8741);
and U11232 (N_11232,N_6938,N_9375);
or U11233 (N_11233,N_9060,N_5098);
and U11234 (N_11234,N_8039,N_6453);
nand U11235 (N_11235,N_7351,N_5496);
nor U11236 (N_11236,N_6644,N_7252);
nand U11237 (N_11237,N_8724,N_6047);
nor U11238 (N_11238,N_8657,N_9842);
nor U11239 (N_11239,N_7398,N_5707);
or U11240 (N_11240,N_7272,N_6221);
nand U11241 (N_11241,N_7228,N_6850);
or U11242 (N_11242,N_5139,N_7803);
or U11243 (N_11243,N_9688,N_9796);
and U11244 (N_11244,N_8568,N_7750);
nand U11245 (N_11245,N_6295,N_8636);
xor U11246 (N_11246,N_8948,N_6247);
or U11247 (N_11247,N_7868,N_9494);
nor U11248 (N_11248,N_5542,N_9185);
or U11249 (N_11249,N_8620,N_6258);
nor U11250 (N_11250,N_8348,N_8863);
xor U11251 (N_11251,N_7483,N_8654);
xnor U11252 (N_11252,N_7105,N_5866);
or U11253 (N_11253,N_9169,N_6561);
nor U11254 (N_11254,N_7405,N_7377);
nor U11255 (N_11255,N_8978,N_5424);
and U11256 (N_11256,N_5695,N_7529);
nand U11257 (N_11257,N_9091,N_6538);
nor U11258 (N_11258,N_9703,N_8380);
xnor U11259 (N_11259,N_9464,N_7106);
or U11260 (N_11260,N_6667,N_7148);
nand U11261 (N_11261,N_8390,N_8944);
xnor U11262 (N_11262,N_8796,N_8396);
and U11263 (N_11263,N_5699,N_7151);
and U11264 (N_11264,N_5589,N_9049);
xor U11265 (N_11265,N_7838,N_5476);
xnor U11266 (N_11266,N_8711,N_8042);
nand U11267 (N_11267,N_9255,N_5457);
xor U11268 (N_11268,N_5682,N_6539);
and U11269 (N_11269,N_8172,N_9003);
or U11270 (N_11270,N_7476,N_5909);
nand U11271 (N_11271,N_6844,N_8372);
nand U11272 (N_11272,N_6742,N_5088);
nor U11273 (N_11273,N_6570,N_5969);
nor U11274 (N_11274,N_6896,N_8713);
or U11275 (N_11275,N_8723,N_6364);
or U11276 (N_11276,N_8036,N_8513);
xor U11277 (N_11277,N_5533,N_7197);
nor U11278 (N_11278,N_5263,N_6651);
or U11279 (N_11279,N_7595,N_9308);
and U11280 (N_11280,N_6617,N_6246);
nand U11281 (N_11281,N_9231,N_8904);
or U11282 (N_11282,N_8603,N_5319);
and U11283 (N_11283,N_9155,N_6831);
nand U11284 (N_11284,N_5220,N_6208);
nand U11285 (N_11285,N_6693,N_8011);
nand U11286 (N_11286,N_6819,N_5404);
nor U11287 (N_11287,N_7028,N_7566);
or U11288 (N_11288,N_5100,N_8209);
or U11289 (N_11289,N_8992,N_5506);
or U11290 (N_11290,N_7943,N_7049);
nand U11291 (N_11291,N_9465,N_7423);
xor U11292 (N_11292,N_5066,N_7294);
nor U11293 (N_11293,N_5567,N_9239);
or U11294 (N_11294,N_8466,N_8716);
and U11295 (N_11295,N_5714,N_6696);
or U11296 (N_11296,N_7258,N_6596);
nand U11297 (N_11297,N_7519,N_9752);
and U11298 (N_11298,N_5716,N_8345);
nor U11299 (N_11299,N_7633,N_8488);
or U11300 (N_11300,N_6194,N_6540);
or U11301 (N_11301,N_8320,N_8915);
or U11302 (N_11302,N_8810,N_5228);
nor U11303 (N_11303,N_7678,N_9240);
xnor U11304 (N_11304,N_7121,N_9051);
and U11305 (N_11305,N_6271,N_5304);
and U11306 (N_11306,N_7801,N_6895);
nor U11307 (N_11307,N_8720,N_7303);
and U11308 (N_11308,N_8661,N_8987);
nor U11309 (N_11309,N_7996,N_6480);
and U11310 (N_11310,N_7849,N_8622);
nand U11311 (N_11311,N_7046,N_6704);
nand U11312 (N_11312,N_8413,N_6576);
nand U11313 (N_11313,N_6227,N_7437);
nand U11314 (N_11314,N_8952,N_5864);
and U11315 (N_11315,N_6712,N_6753);
and U11316 (N_11316,N_7157,N_5887);
and U11317 (N_11317,N_9422,N_9099);
nand U11318 (N_11318,N_7250,N_7667);
and U11319 (N_11319,N_8204,N_6606);
nand U11320 (N_11320,N_5196,N_7471);
and U11321 (N_11321,N_8151,N_8200);
or U11322 (N_11322,N_5915,N_5501);
xor U11323 (N_11323,N_7717,N_5984);
nor U11324 (N_11324,N_9138,N_6177);
or U11325 (N_11325,N_9821,N_6305);
nand U11326 (N_11326,N_7234,N_6424);
and U11327 (N_11327,N_9406,N_8600);
xnor U11328 (N_11328,N_8726,N_8643);
or U11329 (N_11329,N_7149,N_9319);
or U11330 (N_11330,N_6873,N_5833);
nand U11331 (N_11331,N_6346,N_8776);
or U11332 (N_11332,N_6057,N_6881);
or U11333 (N_11333,N_7305,N_6522);
and U11334 (N_11334,N_6070,N_6432);
nand U11335 (N_11335,N_8436,N_8606);
nor U11336 (N_11336,N_9351,N_7821);
nand U11337 (N_11337,N_5254,N_9248);
and U11338 (N_11338,N_8847,N_5852);
xor U11339 (N_11339,N_8757,N_6513);
or U11340 (N_11340,N_8415,N_7909);
and U11341 (N_11341,N_8507,N_5958);
xnor U11342 (N_11342,N_6215,N_6167);
nor U11343 (N_11343,N_6592,N_9626);
xnor U11344 (N_11344,N_5324,N_6377);
and U11345 (N_11345,N_8633,N_8405);
nor U11346 (N_11346,N_8481,N_9873);
and U11347 (N_11347,N_5027,N_7052);
and U11348 (N_11348,N_5377,N_7366);
or U11349 (N_11349,N_6059,N_6182);
or U11350 (N_11350,N_7716,N_5875);
nand U11351 (N_11351,N_8162,N_6137);
and U11352 (N_11352,N_6106,N_5240);
nand U11353 (N_11353,N_7539,N_6058);
or U11354 (N_11354,N_8856,N_7381);
and U11355 (N_11355,N_8312,N_8431);
nand U11356 (N_11356,N_6980,N_9204);
or U11357 (N_11357,N_7788,N_5230);
and U11358 (N_11358,N_7545,N_8477);
nand U11359 (N_11359,N_5165,N_5536);
nand U11360 (N_11360,N_6872,N_5315);
and U11361 (N_11361,N_8857,N_7119);
and U11362 (N_11362,N_6820,N_8454);
or U11363 (N_11363,N_9338,N_8701);
and U11364 (N_11364,N_9183,N_8356);
and U11365 (N_11365,N_8009,N_6521);
nor U11366 (N_11366,N_7213,N_7879);
nand U11367 (N_11367,N_7103,N_7629);
and U11368 (N_11368,N_9651,N_6260);
and U11369 (N_11369,N_7640,N_6005);
and U11370 (N_11370,N_5418,N_8465);
and U11371 (N_11371,N_7723,N_8999);
nand U11372 (N_11372,N_6815,N_7281);
or U11373 (N_11373,N_8346,N_9678);
or U11374 (N_11374,N_6642,N_7027);
nand U11375 (N_11375,N_8257,N_5029);
nand U11376 (N_11376,N_8076,N_8168);
nand U11377 (N_11377,N_9844,N_7858);
nor U11378 (N_11378,N_7455,N_6476);
and U11379 (N_11379,N_6603,N_6458);
nor U11380 (N_11380,N_7248,N_7593);
xor U11381 (N_11381,N_7180,N_5296);
nor U11382 (N_11382,N_6868,N_6161);
or U11383 (N_11383,N_6923,N_9400);
xnor U11384 (N_11384,N_9480,N_8020);
and U11385 (N_11385,N_5644,N_6785);
and U11386 (N_11386,N_8471,N_9735);
nor U11387 (N_11387,N_7637,N_8691);
nand U11388 (N_11388,N_6171,N_9212);
and U11389 (N_11389,N_9578,N_9016);
nor U11390 (N_11390,N_7434,N_7951);
and U11391 (N_11391,N_8945,N_7500);
xor U11392 (N_11392,N_9782,N_9932);
nor U11393 (N_11393,N_7450,N_6516);
and U11394 (N_11394,N_8400,N_9331);
or U11395 (N_11395,N_9753,N_9896);
nor U11396 (N_11396,N_7422,N_8500);
or U11397 (N_11397,N_6330,N_8334);
and U11398 (N_11398,N_9470,N_6012);
nor U11399 (N_11399,N_7399,N_5335);
nand U11400 (N_11400,N_5757,N_7062);
nor U11401 (N_11401,N_7038,N_9440);
nand U11402 (N_11402,N_6336,N_9741);
and U11403 (N_11403,N_5641,N_8705);
nor U11404 (N_11404,N_6253,N_9197);
or U11405 (N_11405,N_6643,N_8138);
and U11406 (N_11406,N_6600,N_6821);
nand U11407 (N_11407,N_9460,N_8148);
nor U11408 (N_11408,N_8685,N_6420);
and U11409 (N_11409,N_7763,N_7689);
nand U11410 (N_11410,N_6859,N_9817);
and U11411 (N_11411,N_8564,N_9187);
nand U11412 (N_11412,N_7613,N_5350);
nand U11413 (N_11413,N_6233,N_9706);
nor U11414 (N_11414,N_9066,N_9585);
nand U11415 (N_11415,N_5184,N_8430);
and U11416 (N_11416,N_5036,N_8825);
or U11417 (N_11417,N_8655,N_8034);
nor U11418 (N_11418,N_7212,N_6961);
or U11419 (N_11419,N_6568,N_6333);
nand U11420 (N_11420,N_8994,N_6532);
nand U11421 (N_11421,N_6061,N_9065);
nand U11422 (N_11422,N_9444,N_5355);
and U11423 (N_11423,N_5795,N_8731);
or U11424 (N_11424,N_5972,N_6493);
nand U11425 (N_11425,N_5481,N_6341);
or U11426 (N_11426,N_7823,N_8250);
and U11427 (N_11427,N_5559,N_6292);
and U11428 (N_11428,N_6669,N_9885);
and U11429 (N_11429,N_9898,N_9009);
nor U11430 (N_11430,N_5071,N_5849);
nand U11431 (N_11431,N_7413,N_9609);
nor U11432 (N_11432,N_5124,N_6773);
nand U11433 (N_11433,N_6225,N_5813);
nand U11434 (N_11434,N_8196,N_8840);
and U11435 (N_11435,N_8702,N_7348);
or U11436 (N_11436,N_6737,N_6272);
and U11437 (N_11437,N_7296,N_5830);
or U11438 (N_11438,N_9934,N_5810);
nand U11439 (N_11439,N_7280,N_6471);
or U11440 (N_11440,N_8191,N_6360);
nor U11441 (N_11441,N_9630,N_8712);
nand U11442 (N_11442,N_5711,N_7744);
nor U11443 (N_11443,N_9915,N_9760);
nand U11444 (N_11444,N_9871,N_8301);
and U11445 (N_11445,N_7628,N_8201);
nand U11446 (N_11446,N_9503,N_9705);
nor U11447 (N_11447,N_5111,N_5400);
or U11448 (N_11448,N_9355,N_7124);
xor U11449 (N_11449,N_5440,N_9648);
nand U11450 (N_11450,N_6015,N_8150);
nand U11451 (N_11451,N_6013,N_8567);
or U11452 (N_11452,N_7922,N_8175);
xnor U11453 (N_11453,N_8386,N_9863);
nand U11454 (N_11454,N_8103,N_6746);
nor U11455 (N_11455,N_7652,N_6999);
and U11456 (N_11456,N_7222,N_5235);
nor U11457 (N_11457,N_9222,N_9624);
nor U11458 (N_11458,N_8495,N_8001);
nor U11459 (N_11459,N_6335,N_7247);
nor U11460 (N_11460,N_9242,N_9453);
nand U11461 (N_11461,N_9372,N_6695);
or U11462 (N_11462,N_7486,N_6575);
and U11463 (N_11463,N_9916,N_7171);
or U11464 (N_11464,N_7194,N_6248);
and U11465 (N_11465,N_7898,N_5579);
or U11466 (N_11466,N_6153,N_9401);
and U11467 (N_11467,N_8279,N_9473);
and U11468 (N_11468,N_5940,N_5538);
xor U11469 (N_11469,N_7000,N_7987);
or U11470 (N_11470,N_6591,N_8051);
xor U11471 (N_11471,N_8839,N_8016);
nand U11472 (N_11472,N_7081,N_8238);
nor U11473 (N_11473,N_7335,N_9431);
xnor U11474 (N_11474,N_6879,N_9357);
nor U11475 (N_11475,N_8391,N_8186);
or U11476 (N_11476,N_7432,N_8115);
nand U11477 (N_11477,N_6705,N_6972);
and U11478 (N_11478,N_6110,N_5577);
nor U11479 (N_11479,N_7771,N_6343);
nor U11480 (N_11480,N_9341,N_9165);
or U11481 (N_11481,N_9377,N_9089);
or U11482 (N_11482,N_7232,N_9985);
nand U11483 (N_11483,N_6028,N_9441);
nand U11484 (N_11484,N_6777,N_7877);
and U11485 (N_11485,N_5104,N_6579);
nand U11486 (N_11486,N_5396,N_7776);
nor U11487 (N_11487,N_7775,N_9718);
nor U11488 (N_11488,N_7026,N_6956);
or U11489 (N_11489,N_8502,N_5256);
or U11490 (N_11490,N_9737,N_5966);
nor U11491 (N_11491,N_8086,N_8387);
nor U11492 (N_11492,N_7444,N_5930);
or U11493 (N_11493,N_8432,N_8710);
nor U11494 (N_11494,N_5479,N_7375);
or U11495 (N_11495,N_7876,N_5623);
xor U11496 (N_11496,N_9694,N_5004);
and U11497 (N_11497,N_8637,N_5189);
and U11498 (N_11498,N_6525,N_6031);
or U11499 (N_11499,N_8618,N_5471);
nand U11500 (N_11500,N_5454,N_6982);
nor U11501 (N_11501,N_7164,N_7857);
nand U11502 (N_11502,N_8571,N_6841);
nor U11503 (N_11503,N_5629,N_7286);
and U11504 (N_11504,N_9149,N_8030);
nand U11505 (N_11505,N_5919,N_7210);
nand U11506 (N_11506,N_9287,N_5992);
nand U11507 (N_11507,N_6962,N_8099);
and U11508 (N_11508,N_5121,N_7188);
or U11509 (N_11509,N_5272,N_6663);
or U11510 (N_11510,N_8033,N_5435);
xor U11511 (N_11511,N_6557,N_6091);
nand U11512 (N_11512,N_8349,N_6500);
nand U11513 (N_11513,N_8433,N_9679);
and U11514 (N_11514,N_5740,N_8521);
nand U11515 (N_11515,N_9069,N_6395);
or U11516 (N_11516,N_6776,N_6278);
nor U11517 (N_11517,N_6620,N_9378);
nor U11518 (N_11518,N_5417,N_7056);
and U11519 (N_11519,N_9945,N_8078);
nor U11520 (N_11520,N_8801,N_9142);
nor U11521 (N_11521,N_7439,N_7241);
nor U11522 (N_11522,N_5512,N_5880);
or U11523 (N_11523,N_5192,N_7810);
nor U11524 (N_11524,N_9108,N_6792);
nor U11525 (N_11525,N_6345,N_5624);
nor U11526 (N_11526,N_7482,N_9977);
nor U11527 (N_11527,N_7347,N_6832);
xnor U11528 (N_11528,N_6107,N_6269);
or U11529 (N_11529,N_9539,N_7176);
xor U11530 (N_11530,N_5317,N_8516);
nand U11531 (N_11531,N_8375,N_9577);
or U11532 (N_11532,N_6317,N_8243);
nand U11533 (N_11533,N_5217,N_9888);
nor U11534 (N_11534,N_8913,N_6299);
or U11535 (N_11535,N_7548,N_9292);
nand U11536 (N_11536,N_7150,N_5788);
nand U11537 (N_11537,N_7619,N_8124);
nor U11538 (N_11538,N_7326,N_8285);
and U11539 (N_11539,N_7214,N_5214);
nor U11540 (N_11540,N_7662,N_9616);
and U11541 (N_11541,N_5293,N_7787);
or U11542 (N_11542,N_9699,N_8416);
and U11543 (N_11543,N_8922,N_8811);
and U11544 (N_11544,N_7556,N_8377);
and U11545 (N_11545,N_7047,N_5888);
or U11546 (N_11546,N_6151,N_6857);
or U11547 (N_11547,N_8304,N_6212);
nand U11548 (N_11548,N_7732,N_8342);
or U11549 (N_11549,N_5249,N_8940);
and U11550 (N_11550,N_8475,N_8980);
nor U11551 (N_11551,N_6976,N_9795);
nand U11552 (N_11552,N_9680,N_7218);
nand U11553 (N_11553,N_9804,N_9088);
or U11554 (N_11554,N_7359,N_6357);
and U11555 (N_11555,N_5733,N_7479);
nor U11556 (N_11556,N_6138,N_7435);
and U11557 (N_11557,N_5074,N_8198);
or U11558 (N_11558,N_8572,N_5652);
nor U11559 (N_11559,N_7265,N_7938);
xor U11560 (N_11560,N_6700,N_8193);
nor U11561 (N_11561,N_8219,N_8463);
nor U11562 (N_11562,N_6605,N_6907);
nand U11563 (N_11563,N_7866,N_9557);
and U11564 (N_11564,N_9743,N_6256);
nor U11565 (N_11565,N_6130,N_9763);
nor U11566 (N_11566,N_6640,N_7891);
and U11567 (N_11567,N_9439,N_7623);
nor U11568 (N_11568,N_7481,N_7783);
and U11569 (N_11569,N_9266,N_8549);
or U11570 (N_11570,N_9014,N_6970);
nand U11571 (N_11571,N_9136,N_7494);
nor U11572 (N_11572,N_6383,N_8097);
and U11573 (N_11573,N_7747,N_6485);
or U11574 (N_11574,N_8456,N_5614);
xor U11575 (N_11575,N_8775,N_9087);
nor U11576 (N_11576,N_8049,N_6375);
or U11577 (N_11577,N_5325,N_7994);
or U11578 (N_11578,N_8509,N_5678);
nor U11579 (N_11579,N_6547,N_8837);
and U11580 (N_11580,N_7063,N_6799);
and U11581 (N_11581,N_5035,N_9854);
nor U11582 (N_11582,N_9904,N_9420);
nand U11583 (N_11583,N_8681,N_8773);
nand U11584 (N_11584,N_6825,N_8558);
or U11585 (N_11585,N_7993,N_9397);
or U11586 (N_11586,N_6311,N_7291);
nor U11587 (N_11587,N_5041,N_5212);
and U11588 (N_11588,N_6374,N_9955);
and U11589 (N_11589,N_7264,N_9385);
nand U11590 (N_11590,N_7205,N_6294);
or U11591 (N_11591,N_7368,N_8158);
or U11592 (N_11592,N_6677,N_8557);
or U11593 (N_11593,N_7574,N_8565);
xnor U11594 (N_11594,N_8890,N_6380);
and U11595 (N_11595,N_7523,N_9759);
or U11596 (N_11596,N_7604,N_6128);
xor U11597 (N_11597,N_8202,N_9547);
nand U11598 (N_11598,N_5209,N_5596);
xnor U11599 (N_11599,N_7384,N_9234);
nand U11600 (N_11600,N_6118,N_9770);
nand U11601 (N_11601,N_7671,N_9696);
nand U11602 (N_11602,N_5460,N_5816);
nor U11603 (N_11603,N_8894,N_9479);
and U11604 (N_11604,N_5158,N_8460);
or U11605 (N_11605,N_5700,N_9739);
nor U11606 (N_11606,N_9727,N_9908);
nand U11607 (N_11607,N_6428,N_6889);
nand U11608 (N_11608,N_8512,N_5735);
nor U11609 (N_11609,N_7575,N_7948);
nand U11610 (N_11610,N_6595,N_9815);
or U11611 (N_11611,N_6944,N_6685);
or U11612 (N_11612,N_6266,N_9168);
and U11613 (N_11613,N_5883,N_9806);
xnor U11614 (N_11614,N_9588,N_8252);
nor U11615 (N_11615,N_7004,N_5999);
or U11616 (N_11616,N_6155,N_5784);
or U11617 (N_11617,N_8087,N_7999);
nor U11618 (N_11618,N_7267,N_6953);
nand U11619 (N_11619,N_7461,N_5936);
nand U11620 (N_11620,N_8242,N_7630);
nand U11621 (N_11621,N_5065,N_5719);
and U11622 (N_11622,N_9966,N_6218);
nand U11623 (N_11623,N_8580,N_7350);
and U11624 (N_11624,N_7084,N_8912);
xnor U11625 (N_11625,N_8523,N_6608);
or U11626 (N_11626,N_5964,N_7537);
or U11627 (N_11627,N_5857,N_5545);
or U11628 (N_11628,N_5340,N_7761);
or U11629 (N_11629,N_6078,N_6910);
nor U11630 (N_11630,N_8330,N_8340);
or U11631 (N_11631,N_6715,N_8239);
and U11632 (N_11632,N_6267,N_9989);
nand U11633 (N_11633,N_8729,N_7307);
and U11634 (N_11634,N_5449,N_8765);
and U11635 (N_11635,N_5604,N_5552);
and U11636 (N_11636,N_7111,N_5283);
xor U11637 (N_11637,N_6702,N_6124);
and U11638 (N_11638,N_5478,N_6046);
or U11639 (N_11639,N_8938,N_6342);
xor U11640 (N_11640,N_5848,N_7748);
or U11641 (N_11641,N_5032,N_7236);
and U11642 (N_11642,N_9700,N_7254);
and U11643 (N_11643,N_8780,N_6447);
nand U11644 (N_11644,N_8519,N_8476);
nor U11645 (N_11645,N_8570,N_5749);
nor U11646 (N_11646,N_6203,N_9660);
nand U11647 (N_11647,N_8423,N_6197);
or U11648 (N_11648,N_8050,N_9661);
nor U11649 (N_11649,N_5645,N_8674);
and U11650 (N_11650,N_6738,N_9320);
xnor U11651 (N_11651,N_8393,N_9163);
and U11652 (N_11652,N_5656,N_5758);
and U11653 (N_11653,N_7182,N_9115);
or U11654 (N_11654,N_9358,N_8767);
or U11655 (N_11655,N_7871,N_7908);
nand U11656 (N_11656,N_5879,N_8082);
nor U11657 (N_11657,N_6411,N_8581);
or U11658 (N_11658,N_6653,N_5007);
nor U11659 (N_11659,N_8295,N_7897);
xor U11660 (N_11660,N_8522,N_5523);
or U11661 (N_11661,N_6090,N_8902);
and U11662 (N_11662,N_6988,N_9476);
or U11663 (N_11663,N_6352,N_8642);
or U11664 (N_11664,N_9567,N_6449);
nand U11665 (N_11665,N_9773,N_6099);
nor U11666 (N_11666,N_8137,N_7333);
nor U11667 (N_11667,N_8104,N_5508);
nand U11668 (N_11668,N_5085,N_7708);
and U11669 (N_11669,N_7829,N_7468);
nand U11670 (N_11670,N_9186,N_7946);
or U11671 (N_11671,N_9629,N_5056);
nand U11672 (N_11672,N_9940,N_8611);
nand U11673 (N_11673,N_5619,N_6052);
nor U11674 (N_11674,N_6051,N_8004);
and U11675 (N_11675,N_5207,N_5734);
or U11676 (N_11676,N_7573,N_6968);
xor U11677 (N_11677,N_9625,N_6459);
or U11678 (N_11678,N_5129,N_8254);
or U11679 (N_11679,N_9113,N_9719);
or U11680 (N_11680,N_7851,N_9861);
and U11681 (N_11681,N_7037,N_7403);
xor U11682 (N_11682,N_5584,N_9497);
or U11683 (N_11683,N_7968,N_6800);
or U11684 (N_11684,N_6678,N_9387);
nand U11685 (N_11685,N_5102,N_8012);
and U11686 (N_11686,N_7498,N_7380);
nand U11687 (N_11687,N_9015,N_9827);
nand U11688 (N_11688,N_5590,N_6088);
nor U11689 (N_11689,N_5126,N_5494);
and U11690 (N_11690,N_6625,N_7117);
nor U11691 (N_11691,N_7777,N_9845);
and U11692 (N_11692,N_5037,N_6843);
and U11693 (N_11693,N_9391,N_9830);
or U11694 (N_11694,N_5337,N_9446);
xor U11695 (N_11695,N_6235,N_7508);
nand U11696 (N_11696,N_9071,N_9364);
or U11697 (N_11697,N_5043,N_6164);
nand U11698 (N_11698,N_5780,N_6223);
nor U11699 (N_11699,N_5026,N_9148);
nand U11700 (N_11700,N_5770,N_6097);
nor U11701 (N_11701,N_9687,N_8300);
xnor U11702 (N_11702,N_9485,N_5616);
nor U11703 (N_11703,N_7034,N_5426);
nand U11704 (N_11704,N_9354,N_5585);
nor U11705 (N_11705,N_6009,N_7953);
nor U11706 (N_11706,N_8065,N_7731);
or U11707 (N_11707,N_8589,N_7393);
and U11708 (N_11708,N_7521,N_9514);
nand U11709 (N_11709,N_5233,N_6658);
and U11710 (N_11710,N_8738,N_7746);
or U11711 (N_11711,N_6798,N_5868);
or U11712 (N_11712,N_8407,N_7625);
and U11713 (N_11713,N_9670,N_5692);
and U11714 (N_11714,N_8353,N_9765);
nand U11715 (N_11715,N_5620,N_5951);
nor U11716 (N_11716,N_6512,N_7285);
nand U11717 (N_11717,N_9280,N_6486);
nor U11718 (N_11718,N_7243,N_5634);
or U11719 (N_11719,N_5070,N_9263);
nor U11720 (N_11720,N_5011,N_5685);
nand U11721 (N_11721,N_6438,N_5389);
and U11722 (N_11722,N_9035,N_6291);
nor U11723 (N_11723,N_9936,N_6255);
and U11724 (N_11724,N_6692,N_5934);
nand U11725 (N_11725,N_6622,N_6379);
nor U11726 (N_11726,N_5251,N_9102);
nor U11727 (N_11727,N_9901,N_5822);
nor U11728 (N_11728,N_5896,N_6986);
nor U11729 (N_11729,N_8751,N_6079);
xor U11730 (N_11730,N_6300,N_9967);
or U11731 (N_11731,N_8056,N_7251);
or U11732 (N_11732,N_8395,N_5328);
or U11733 (N_11733,N_7757,N_9064);
nor U11734 (N_11734,N_6609,N_8525);
and U11735 (N_11735,N_8421,N_6261);
and U11736 (N_11736,N_6043,N_7257);
nand U11737 (N_11737,N_5970,N_8351);
xor U11738 (N_11738,N_8663,N_5599);
xnor U11739 (N_11739,N_6505,N_9297);
nor U11740 (N_11740,N_8182,N_5803);
nand U11741 (N_11741,N_8045,N_9369);
and U11742 (N_11742,N_6749,N_9107);
nand U11743 (N_11743,N_7781,N_5612);
or U11744 (N_11744,N_5679,N_7892);
xor U11745 (N_11745,N_8752,N_5259);
nand U11746 (N_11746,N_9498,N_8877);
or U11747 (N_11747,N_7363,N_9172);
and U11748 (N_11748,N_8656,N_8916);
or U11749 (N_11749,N_8160,N_9643);
and U11750 (N_11750,N_8105,N_5975);
and U11751 (N_11751,N_8310,N_5527);
and U11752 (N_11752,N_8314,N_5592);
nand U11753 (N_11753,N_7610,N_9237);
or U11754 (N_11754,N_9472,N_8527);
and U11755 (N_11755,N_7655,N_9396);
and U11756 (N_11756,N_8185,N_5793);
xnor U11757 (N_11757,N_6862,N_7065);
xor U11758 (N_11758,N_9281,N_5226);
and U11759 (N_11759,N_5683,N_5394);
nand U11760 (N_11760,N_8284,N_8955);
xor U11761 (N_11761,N_7196,N_6206);
xor U11762 (N_11762,N_6769,N_5285);
nand U11763 (N_11763,N_9002,N_9127);
or U11764 (N_11764,N_7837,N_8588);
and U11765 (N_11765,N_7997,N_5709);
or U11766 (N_11766,N_9079,N_6217);
and U11767 (N_11767,N_5406,N_5238);
nand U11768 (N_11768,N_5267,N_9598);
nand U11769 (N_11769,N_9056,N_9526);
or U11770 (N_11770,N_9086,N_9425);
and U11771 (N_11771,N_6142,N_8308);
nand U11772 (N_11772,N_7115,N_9210);
nor U11773 (N_11773,N_6156,N_6168);
nor U11774 (N_11774,N_7622,N_9900);
or U11775 (N_11775,N_6228,N_8666);
or U11776 (N_11776,N_7319,N_8682);
nor U11777 (N_11777,N_6666,N_5886);
and U11778 (N_11778,N_6838,N_6324);
xor U11779 (N_11779,N_6597,N_6761);
or U11780 (N_11780,N_9789,N_6180);
xnor U11781 (N_11781,N_5739,N_7400);
xor U11782 (N_11782,N_6388,N_9571);
and U11783 (N_11783,N_9914,N_8623);
or U11784 (N_11784,N_9469,N_5801);
nor U11785 (N_11785,N_6519,N_9715);
or U11786 (N_11786,N_9116,N_7273);
xnor U11787 (N_11787,N_9622,N_7813);
nand U11788 (N_11788,N_5490,N_6626);
or U11789 (N_11789,N_5906,N_8409);
nand U11790 (N_11790,N_6562,N_5942);
nand U11791 (N_11791,N_5020,N_7373);
and U11792 (N_11792,N_7576,N_7178);
xor U11793 (N_11793,N_5850,N_7473);
nor U11794 (N_11794,N_7532,N_8152);
or U11795 (N_11795,N_7636,N_9285);
or U11796 (N_11796,N_5023,N_7404);
nor U11797 (N_11797,N_7896,N_8296);
nor U11798 (N_11798,N_7100,N_5808);
nand U11799 (N_11799,N_9026,N_6489);
or U11800 (N_11800,N_6877,N_7513);
nor U11801 (N_11801,N_7041,N_7815);
xor U11802 (N_11802,N_6165,N_6264);
and U11803 (N_11803,N_8118,N_5386);
and U11804 (N_11804,N_6874,N_8283);
and U11805 (N_11805,N_5721,N_6811);
nand U11806 (N_11806,N_5933,N_5805);
and U11807 (N_11807,N_7071,N_7852);
nor U11808 (N_11808,N_6038,N_7154);
nor U11809 (N_11809,N_7183,N_6679);
or U11810 (N_11810,N_8382,N_5470);
nor U11811 (N_11811,N_5503,N_7200);
nand U11812 (N_11812,N_7644,N_6784);
and U11813 (N_11813,N_9610,N_7238);
nor U11814 (N_11814,N_5138,N_9594);
and U11815 (N_11815,N_7720,N_7912);
nand U11816 (N_11816,N_7758,N_8866);
nand U11817 (N_11817,N_5155,N_6833);
xor U11818 (N_11818,N_5297,N_7979);
nand U11819 (N_11819,N_6166,N_8977);
nor U11820 (N_11820,N_8874,N_7914);
or U11821 (N_11821,N_5119,N_8886);
nand U11822 (N_11822,N_6229,N_7163);
nand U11823 (N_11823,N_9426,N_7102);
or U11824 (N_11824,N_9825,N_8974);
or U11825 (N_11825,N_5555,N_5343);
or U11826 (N_11826,N_5646,N_7749);
nand U11827 (N_11827,N_7321,N_5250);
and U11828 (N_11828,N_7013,N_5594);
and U11829 (N_11829,N_9986,N_8057);
and U11830 (N_11830,N_7077,N_7441);
nor U11831 (N_11831,N_8261,N_5474);
or U11832 (N_11832,N_5766,N_5867);
nand U11833 (N_11833,N_8883,N_6071);
and U11834 (N_11834,N_6967,N_7177);
nand U11835 (N_11835,N_6123,N_6415);
nand U11836 (N_11836,N_6479,N_5558);
nand U11837 (N_11837,N_7590,N_9329);
and U11838 (N_11838,N_9315,N_8778);
nand U11839 (N_11839,N_5703,N_8627);
nand U11840 (N_11840,N_7142,N_7022);
or U11841 (N_11841,N_9677,N_6230);
and U11842 (N_11842,N_7734,N_6365);
nor U11843 (N_11843,N_6109,N_9487);
or U11844 (N_11844,N_8601,N_5176);
nand U11845 (N_11845,N_5507,N_9639);
nand U11846 (N_11846,N_9747,N_9553);
nor U11847 (N_11847,N_6133,N_8537);
nand U11848 (N_11848,N_6312,N_5672);
or U11849 (N_11849,N_9043,N_6745);
nor U11850 (N_11850,N_7699,N_9587);
xnor U11851 (N_11851,N_9628,N_7401);
nand U11852 (N_11852,N_5286,N_8482);
and U11853 (N_11853,N_9756,N_7559);
nand U11854 (N_11854,N_9544,N_5108);
and U11855 (N_11855,N_7790,N_5169);
nand U11856 (N_11856,N_9059,N_9755);
or U11857 (N_11857,N_8113,N_7729);
nor U11858 (N_11858,N_7684,N_9930);
and U11859 (N_11859,N_7485,N_9809);
nand U11860 (N_11860,N_5019,N_8064);
nor U11861 (N_11861,N_5201,N_6796);
nand U11862 (N_11862,N_5115,N_5938);
and U11863 (N_11863,N_6268,N_7960);
or U11864 (N_11864,N_8878,N_8590);
nor U11865 (N_11865,N_7778,N_9653);
nand U11866 (N_11866,N_5288,N_5635);
or U11867 (N_11867,N_5715,N_8233);
nor U11868 (N_11868,N_9272,N_6448);
or U11869 (N_11869,N_5736,N_6725);
nor U11870 (N_11870,N_7915,N_5688);
nor U11871 (N_11871,N_6995,N_6040);
nand U11872 (N_11872,N_6965,N_6507);
nor U11873 (N_11873,N_9671,N_8807);
nand U11874 (N_11874,N_8798,N_9767);
nor U11875 (N_11875,N_6222,N_7624);
or U11876 (N_11876,N_7618,N_8586);
nor U11877 (N_11877,N_7416,N_5075);
nor U11878 (N_11878,N_5953,N_5844);
nor U11879 (N_11879,N_5205,N_6033);
and U11880 (N_11880,N_7981,N_8327);
xnor U11881 (N_11881,N_8925,N_8541);
and U11882 (N_11882,N_7833,N_7970);
nor U11883 (N_11883,N_9647,N_7118);
xor U11884 (N_11884,N_6147,N_9505);
nand U11885 (N_11885,N_7988,N_5980);
nand U11886 (N_11886,N_6810,N_6655);
nand U11887 (N_11887,N_9984,N_8031);
or U11888 (N_11888,N_8652,N_9205);
nor U11889 (N_11889,N_8366,N_9834);
and U11890 (N_11890,N_7330,N_5551);
or U11891 (N_11891,N_8966,N_6209);
or U11892 (N_11892,N_6026,N_5530);
nand U11893 (N_11893,N_7445,N_7983);
and U11894 (N_11894,N_9993,N_9769);
and U11895 (N_11895,N_7745,N_6766);
nand U11896 (N_11896,N_7606,N_8806);
or U11897 (N_11897,N_8943,N_8490);
or U11898 (N_11898,N_8676,N_8956);
nor U11899 (N_11899,N_5655,N_7429);
nand U11900 (N_11900,N_6537,N_7949);
and U11901 (N_11901,N_9536,N_8058);
xnor U11902 (N_11902,N_8747,N_9133);
or U11903 (N_11903,N_9880,N_6585);
nor U11904 (N_11904,N_6452,N_7339);
nor U11905 (N_11905,N_6497,N_7597);
or U11906 (N_11906,N_6207,N_8077);
nand U11907 (N_11907,N_7752,N_7245);
nand U11908 (N_11908,N_7036,N_5344);
and U11909 (N_11909,N_5132,N_5180);
nor U11910 (N_11910,N_9445,N_5796);
xnor U11911 (N_11911,N_8098,N_8059);
or U11912 (N_11912,N_7706,N_6759);
nand U11913 (N_11913,N_6116,N_7017);
or U11914 (N_11914,N_6718,N_7739);
and U11915 (N_11915,N_7927,N_7365);
or U11916 (N_11916,N_8678,N_7499);
nand U11917 (N_11917,N_5534,N_8221);
nor U11918 (N_11918,N_5279,N_7226);
nor U11919 (N_11919,N_9762,N_5622);
nor U11920 (N_11920,N_7865,N_7703);
nand U11921 (N_11921,N_7466,N_5430);
and U11922 (N_11922,N_7260,N_8855);
or U11923 (N_11923,N_6602,N_6854);
nand U11924 (N_11924,N_9200,N_5049);
nor U11925 (N_11925,N_8276,N_7795);
nand U11926 (N_11926,N_6056,N_6637);
nor U11927 (N_11927,N_9596,N_5950);
and U11928 (N_11928,N_8094,N_9563);
xnor U11929 (N_11929,N_9920,N_6936);
xor U11930 (N_11930,N_5948,N_9722);
or U11931 (N_11931,N_5724,N_5197);
nor U11932 (N_11932,N_7308,N_6774);
xnor U11933 (N_11933,N_5097,N_8487);
xnor U11934 (N_11934,N_9637,N_8213);
or U11935 (N_11935,N_6733,N_9403);
nor U11936 (N_11936,N_9450,N_5330);
or U11937 (N_11937,N_5510,N_6652);
or U11938 (N_11938,N_6450,N_7024);
xor U11939 (N_11939,N_9590,N_5631);
nand U11940 (N_11940,N_5768,N_6930);
or U11941 (N_11941,N_7990,N_8562);
nor U11942 (N_11942,N_8322,N_6781);
nor U11943 (N_11943,N_7753,N_9886);
and U11944 (N_11944,N_6555,N_8813);
nor U11945 (N_11945,N_8411,N_9764);
xor U11946 (N_11946,N_8417,N_5680);
nand U11947 (N_11947,N_9011,N_8771);
nand U11948 (N_11948,N_6717,N_6373);
and U11949 (N_11949,N_7826,N_9463);
or U11950 (N_11950,N_8660,N_8442);
nor U11951 (N_11951,N_7058,N_5576);
nand U11952 (N_11952,N_5902,N_8824);
and U11953 (N_11953,N_9991,N_7511);
or U11954 (N_11954,N_8333,N_7174);
and U11955 (N_11955,N_8024,N_5473);
nor U11956 (N_11956,N_5988,N_5627);
and U11957 (N_11957,N_8135,N_6474);
or U11958 (N_11958,N_9929,N_6404);
or U11959 (N_11959,N_9559,N_6950);
or U11960 (N_11960,N_6250,N_5785);
nor U11961 (N_11961,N_7585,N_7611);
xor U11962 (N_11962,N_7738,N_9837);
nor U11963 (N_11963,N_7691,N_9745);
or U11964 (N_11964,N_5379,N_8374);
nand U11965 (N_11965,N_9858,N_6066);
and U11966 (N_11966,N_9095,N_9294);
and U11967 (N_11967,N_5268,N_7136);
or U11968 (N_11968,N_6179,N_6060);
or U11969 (N_11969,N_5378,N_6297);
nand U11970 (N_11970,N_7598,N_6421);
nor U11971 (N_11971,N_7068,N_6615);
and U11972 (N_11972,N_7918,N_8575);
and U11973 (N_11973,N_9732,N_6224);
nand U11974 (N_11974,N_8969,N_9328);
nand U11975 (N_11975,N_8576,N_7656);
or U11976 (N_11976,N_9952,N_5388);
and U11977 (N_11977,N_9312,N_6618);
and U11978 (N_11978,N_5787,N_8259);
nand U11979 (N_11979,N_6517,N_5107);
or U11980 (N_11980,N_5982,N_5675);
xor U11981 (N_11981,N_6050,N_7495);
or U11982 (N_11982,N_9083,N_8399);
or U11983 (N_11983,N_8062,N_6439);
nor U11984 (N_11984,N_9182,N_9618);
nand U11985 (N_11985,N_8675,N_9742);
nand U11986 (N_11986,N_9802,N_5955);
nor U11987 (N_11987,N_9318,N_7534);
nand U11988 (N_11988,N_8626,N_6762);
nand U11989 (N_11989,N_5492,N_5661);
and U11990 (N_11990,N_7240,N_9933);
nand U11991 (N_11991,N_9256,N_9650);
nand U11992 (N_11992,N_8587,N_5495);
or U11993 (N_11993,N_9701,N_5621);
nand U11994 (N_11994,N_8480,N_9202);
nand U11995 (N_11995,N_5572,N_5826);
nor U11996 (N_11996,N_9190,N_6141);
nand U11997 (N_11997,N_9042,N_7448);
nand U11998 (N_11998,N_8520,N_6901);
and U11999 (N_11999,N_8153,N_7839);
and U12000 (N_12000,N_8458,N_5432);
or U12001 (N_12001,N_7315,N_5926);
and U12002 (N_12002,N_7642,N_8524);
xnor U12003 (N_12003,N_9638,N_8469);
and U12004 (N_12004,N_5626,N_8234);
or U12005 (N_12005,N_9344,N_6590);
or U12006 (N_12006,N_7145,N_5360);
nand U12007 (N_12007,N_7470,N_8419);
and U12008 (N_12008,N_8236,N_9094);
nor U12009 (N_12009,N_9918,N_8719);
nor U12010 (N_12010,N_9927,N_5532);
nand U12011 (N_12011,N_7524,N_9781);
and U12012 (N_12012,N_7292,N_5332);
nor U12013 (N_12013,N_6848,N_9462);
nand U12014 (N_12014,N_9326,N_9173);
and U12015 (N_12015,N_8383,N_8309);
or U12016 (N_12016,N_7454,N_8841);
and U12017 (N_12017,N_5163,N_6369);
and U12018 (N_12018,N_9282,N_8192);
or U12019 (N_12019,N_7798,N_8935);
nand U12020 (N_12020,N_7796,N_6752);
and U12021 (N_12021,N_6708,N_6288);
nor U12022 (N_12022,N_9740,N_8159);
xnor U12023 (N_12023,N_6125,N_8842);
nand U12024 (N_12024,N_7510,N_8338);
or U12025 (N_12025,N_9018,N_8347);
nor U12026 (N_12026,N_9101,N_5899);
or U12027 (N_12027,N_5420,N_5817);
nor U12028 (N_12028,N_9449,N_6772);
or U12029 (N_12029,N_6732,N_9838);
or U12030 (N_12030,N_9175,N_9398);
xor U12031 (N_12031,N_5595,N_6473);
xor U12032 (N_12032,N_8653,N_5993);
and U12033 (N_12033,N_8981,N_7872);
or U12034 (N_12034,N_8428,N_7718);
nor U12035 (N_12035,N_7349,N_9178);
nand U12036 (N_12036,N_6630,N_6724);
and U12037 (N_12037,N_6279,N_6645);
nand U12038 (N_12038,N_9374,N_7249);
and U12039 (N_12039,N_5717,N_9195);
and U12040 (N_12040,N_6629,N_9792);
and U12041 (N_12041,N_9046,N_7958);
nor U12042 (N_12042,N_5876,N_8364);
nand U12043 (N_12043,N_9174,N_9493);
nor U12044 (N_12044,N_9368,N_7420);
xor U12045 (N_12045,N_8256,N_6691);
nand U12046 (N_12046,N_6990,N_8114);
and U12047 (N_12047,N_9617,N_5617);
and U12048 (N_12048,N_5376,N_5973);
nand U12049 (N_12049,N_6120,N_8358);
xnor U12050 (N_12050,N_5900,N_5349);
or U12051 (N_12051,N_6755,N_9414);
or U12052 (N_12052,N_5949,N_7003);
and U12053 (N_12053,N_7229,N_5170);
nor U12054 (N_12054,N_6401,N_6916);
nor U12055 (N_12055,N_5464,N_7447);
nor U12056 (N_12056,N_6552,N_9513);
nor U12057 (N_12057,N_6470,N_9601);
nor U12058 (N_12058,N_7156,N_5222);
nor U12059 (N_12059,N_9790,N_5421);
nor U12060 (N_12060,N_9784,N_8930);
nor U12061 (N_12061,N_9162,N_6616);
nand U12062 (N_12062,N_5994,N_8067);
and U12063 (N_12063,N_8210,N_6633);
and U12064 (N_12064,N_5033,N_6871);
nand U12065 (N_12065,N_7875,N_8154);
nand U12066 (N_12066,N_6392,N_6934);
nor U12067 (N_12067,N_7023,N_8452);
nand U12068 (N_12068,N_5497,N_7409);
nor U12069 (N_12069,N_7430,N_7525);
nor U12070 (N_12070,N_5461,N_8120);
or U12071 (N_12071,N_9111,N_8328);
and U12072 (N_12072,N_8244,N_8573);
nand U12073 (N_12073,N_7067,N_8264);
xnor U12074 (N_12074,N_5081,N_6027);
nand U12075 (N_12075,N_9662,N_8414);
nor U12076 (N_12076,N_8559,N_9379);
nand U12077 (N_12077,N_6041,N_6098);
and U12078 (N_12078,N_9191,N_6276);
or U12079 (N_12079,N_9230,N_5483);
and U12080 (N_12080,N_7195,N_5904);
and U12081 (N_12081,N_9013,N_7793);
xnor U12082 (N_12082,N_9062,N_6405);
or U12083 (N_12083,N_9489,N_5778);
nor U12084 (N_12084,N_7722,N_5611);
nor U12085 (N_12085,N_5024,N_6384);
nor U12086 (N_12086,N_5913,N_7215);
nor U12087 (N_12087,N_6954,N_8493);
nor U12088 (N_12088,N_5015,N_5472);
nor U12089 (N_12089,N_9171,N_8774);
and U12090 (N_12090,N_9143,N_8217);
nand U12091 (N_12091,N_6443,N_7543);
nor U12092 (N_12092,N_5684,N_7759);
or U12093 (N_12093,N_6714,N_7893);
nand U12094 (N_12094,N_7165,N_8293);
nand U12095 (N_12095,N_9313,N_9340);
nor U12096 (N_12096,N_9261,N_6409);
nor U12097 (N_12097,N_5927,N_5164);
and U12098 (N_12098,N_8867,N_9213);
nand U12099 (N_12099,N_9053,N_9389);
nor U12100 (N_12100,N_5287,N_8534);
nand U12101 (N_12101,N_9868,N_7134);
or U12102 (N_12102,N_7209,N_8815);
nand U12103 (N_12103,N_8792,N_5861);
or U12104 (N_12104,N_7449,N_8950);
and U12105 (N_12105,N_8492,N_7006);
or U12106 (N_12106,N_8602,N_9150);
or U12107 (N_12107,N_9455,N_8142);
nor U12108 (N_12108,N_7526,N_7312);
nand U12109 (N_12109,N_7809,N_9365);
nor U12110 (N_12110,N_9818,N_6757);
and U12111 (N_12111,N_8043,N_5080);
nand U12112 (N_12112,N_8975,N_6858);
nor U12113 (N_12113,N_9877,N_8900);
nand U12114 (N_12114,N_9048,N_5034);
nor U12115 (N_12115,N_7266,N_7340);
nor U12116 (N_12116,N_5632,N_6234);
or U12117 (N_12117,N_5499,N_7565);
nand U12118 (N_12118,N_6876,N_8823);
or U12119 (N_12119,N_6022,N_6030);
and U12120 (N_12120,N_8199,N_6989);
or U12121 (N_12121,N_6593,N_6226);
or U12122 (N_12122,N_9640,N_8445);
and U12123 (N_12123,N_8435,N_7175);
and U12124 (N_12124,N_7805,N_5439);
or U12125 (N_12125,N_9951,N_5858);
xnor U12126 (N_12126,N_6017,N_8156);
nand U12127 (N_12127,N_7462,N_8937);
nand U12128 (N_12128,N_6158,N_8046);
or U12129 (N_12129,N_8165,N_6199);
or U12130 (N_12130,N_7527,N_6985);
nor U12131 (N_12131,N_6494,N_9586);
nor U12132 (N_12132,N_7653,N_8044);
nand U12133 (N_12133,N_9907,N_9733);
and U12134 (N_12134,N_6457,N_9223);
nand U12135 (N_12135,N_6136,N_6417);
xnor U12136 (N_12136,N_7239,N_9997);
nand U12137 (N_12137,N_5500,N_6886);
xnor U12138 (N_12138,N_7237,N_9081);
and U12139 (N_12139,N_5965,N_9968);
or U12140 (N_12140,N_6697,N_8505);
nand U12141 (N_12141,N_7019,N_7978);
nand U12142 (N_12142,N_5602,N_6270);
or U12143 (N_12143,N_5570,N_7376);
and U12144 (N_12144,N_9953,N_6870);
and U12145 (N_12145,N_8917,N_5375);
xnor U12146 (N_12146,N_8632,N_9785);
and U12147 (N_12147,N_7522,N_9324);
nor U12148 (N_12148,N_7614,N_7505);
and U12149 (N_12149,N_7051,N_8820);
nand U12150 (N_12150,N_9483,N_6974);
nand U12151 (N_12151,N_5095,N_7418);
xnor U12152 (N_12152,N_5152,N_5664);
xor U12153 (N_12153,N_9707,N_8725);
and U12154 (N_12154,N_8424,N_7586);
xor U12155 (N_12155,N_5303,N_9459);
nor U12156 (N_12156,N_5898,N_6550);
nor U12157 (N_12157,N_7488,N_7998);
xnor U12158 (N_12158,N_9104,N_6332);
and U12159 (N_12159,N_9946,N_9090);
and U12160 (N_12160,N_5524,N_9408);
and U12161 (N_12161,N_8960,N_7431);
or U12162 (N_12162,N_5613,N_6668);
or U12163 (N_12163,N_5062,N_7641);
nor U12164 (N_12164,N_5838,N_9631);
or U12165 (N_12165,N_9938,N_5642);
nor U12166 (N_12166,N_5187,N_6627);
nor U12167 (N_12167,N_9757,N_5221);
nand U12168 (N_12168,N_9799,N_6339);
nor U12169 (N_12169,N_9008,N_5856);
nand U12170 (N_12170,N_5384,N_7255);
or U12171 (N_12171,N_9729,N_9233);
or U12172 (N_12172,N_7669,N_8783);
and U12173 (N_12173,N_6129,N_9203);
nand U12174 (N_12174,N_9411,N_7840);
nor U12175 (N_12175,N_6308,N_7530);
xnor U12176 (N_12176,N_6195,N_9683);
xor U12177 (N_12177,N_5565,N_5147);
xor U12178 (N_12178,N_9196,N_7170);
nand U12179 (N_12179,N_8370,N_8895);
nand U12180 (N_12180,N_5923,N_9206);
nand U12181 (N_12181,N_7268,N_6824);
and U12182 (N_12182,N_6527,N_8909);
xor U12183 (N_12183,N_9636,N_6808);
and U12184 (N_12184,N_6711,N_8483);
nor U12185 (N_12185,N_9589,N_8163);
or U12186 (N_12186,N_5347,N_7712);
and U12187 (N_12187,N_5148,N_7587);
or U12188 (N_12188,N_8858,N_7567);
or U12189 (N_12189,N_5712,N_6611);
nor U12190 (N_12190,N_8484,N_8684);
nor U12191 (N_12191,N_7253,N_6917);
xnor U12192 (N_12192,N_6084,N_6413);
xnor U12193 (N_12193,N_7808,N_7304);
or U12194 (N_12194,N_8933,N_6783);
or U12195 (N_12195,N_5995,N_9779);
and U12196 (N_12196,N_9685,N_9246);
nor U12197 (N_12197,N_9371,N_6159);
and U12198 (N_12198,N_7515,N_8804);
or U12199 (N_12199,N_7553,N_6935);
or U12200 (N_12200,N_7816,N_6906);
nor U12201 (N_12201,N_8140,N_7820);
or U12202 (N_12202,N_7939,N_7192);
or U12203 (N_12203,N_5775,N_8394);
xor U12204 (N_12204,N_8070,N_7371);
nor U12205 (N_12205,N_5237,N_7903);
xnor U12206 (N_12206,N_6149,N_7352);
or U12207 (N_12207,N_7916,N_5390);
xnor U12208 (N_12208,N_5821,N_6621);
and U12209 (N_12209,N_5998,N_9140);
or U12210 (N_12210,N_8918,N_5529);
xnor U12211 (N_12211,N_8270,N_5865);
nor U12212 (N_12212,N_8359,N_7299);
xnor U12213 (N_12213,N_5750,N_9117);
nor U12214 (N_12214,N_5638,N_8768);
nand U12215 (N_12215,N_5889,N_9943);
or U12216 (N_12216,N_8323,N_8246);
and U12217 (N_12217,N_8361,N_5137);
nand U12218 (N_12218,N_9429,N_8091);
nand U12219 (N_12219,N_6675,N_8335);
nor U12220 (N_12220,N_5091,N_5845);
nor U12221 (N_12221,N_6739,N_6670);
and U12222 (N_12222,N_6367,N_7221);
nor U12223 (N_12223,N_9556,N_7332);
xnor U12224 (N_12224,N_9970,N_7974);
or U12225 (N_12225,N_9604,N_8273);
or U12226 (N_12226,N_7414,N_7686);
nand U12227 (N_12227,N_5363,N_9676);
nor U12228 (N_12228,N_5050,N_5618);
and U12229 (N_12229,N_5105,N_9788);
nor U12230 (N_12230,N_7043,N_8605);
nor U12231 (N_12231,N_7607,N_6338);
or U12232 (N_12232,N_9122,N_6337);
and U12233 (N_12233,N_6004,N_8214);
nor U12234 (N_12234,N_6775,N_9193);
or U12235 (N_12235,N_5841,N_8658);
xnor U12236 (N_12236,N_7012,N_6396);
and U12237 (N_12237,N_5677,N_8671);
and U12238 (N_12238,N_5014,N_5574);
and U12239 (N_12239,N_8060,N_7477);
or U12240 (N_12240,N_8189,N_7009);
or U12241 (N_12241,N_6282,N_6694);
nor U12242 (N_12242,N_5996,N_5008);
nor U12243 (N_12243,N_8963,N_5099);
nand U12244 (N_12244,N_8976,N_7621);
nand U12245 (N_12245,N_8376,N_5001);
or U12246 (N_12246,N_9597,N_6183);
nand U12247 (N_12247,N_5794,N_5832);
or U12248 (N_12248,N_6556,N_8230);
nor U12249 (N_12249,N_9899,N_6920);
nand U12250 (N_12250,N_6172,N_8730);
and U12251 (N_12251,N_8634,N_6093);
or U12252 (N_12252,N_8645,N_8957);
and U12253 (N_12253,N_5767,N_8194);
and U12254 (N_12254,N_8750,N_7834);
and U12255 (N_12255,N_9012,N_8584);
nor U12256 (N_12256,N_9443,N_7733);
and U12257 (N_12257,N_9305,N_5047);
nor U12258 (N_12258,N_8090,N_6210);
nor U12259 (N_12259,N_8369,N_7465);
nor U12260 (N_12260,N_7309,N_8350);
and U12261 (N_12261,N_9025,N_8508);
or U12262 (N_12262,N_5366,N_6152);
nor U12263 (N_12263,N_5738,N_9005);
and U12264 (N_12264,N_8923,N_9224);
and U12265 (N_12265,N_6577,N_8425);
xor U12266 (N_12266,N_9366,N_9249);
and U12267 (N_12267,N_8942,N_7284);
and U12268 (N_12268,N_7424,N_6847);
or U12269 (N_12269,N_6032,N_8128);
nand U12270 (N_12270,N_8176,N_9457);
or U12271 (N_12271,N_6257,N_6894);
nor U12272 (N_12272,N_5045,N_9298);
nand U12273 (N_12273,N_6477,N_5660);
xor U12274 (N_12274,N_5731,N_7782);
and U12275 (N_12275,N_5693,N_6119);
nor U12276 (N_12276,N_6673,N_5901);
nand U12277 (N_12277,N_8926,N_8853);
and U12278 (N_12278,N_6619,N_8384);
nor U12279 (N_12279,N_6514,N_5264);
and U12280 (N_12280,N_9033,N_6150);
nand U12281 (N_12281,N_5058,N_9442);
xor U12282 (N_12282,N_5921,N_5882);
or U12283 (N_12283,N_6111,N_7122);
nand U12284 (N_12284,N_6559,N_5393);
nor U12285 (N_12285,N_6200,N_8403);
nand U12286 (N_12286,N_8814,N_9550);
nand U12287 (N_12287,N_8800,N_5380);
nand U12288 (N_12288,N_7085,N_8538);
or U12289 (N_12289,N_7967,N_5229);
nand U12290 (N_12290,N_9917,N_8954);
or U12291 (N_12291,N_7799,N_5257);
or U12292 (N_12292,N_5244,N_6481);
and U12293 (N_12293,N_8498,N_9811);
or U12294 (N_12294,N_6242,N_6793);
nand U12295 (N_12295,N_9496,N_5553);
and U12296 (N_12296,N_7492,N_8008);
and U12297 (N_12297,N_7345,N_6837);
nor U12298 (N_12298,N_8996,N_7199);
nand U12299 (N_12299,N_7357,N_7680);
nor U12300 (N_12300,N_8968,N_9333);
nand U12301 (N_12301,N_8885,N_7814);
xor U12302 (N_12302,N_7705,N_9337);
or U12303 (N_12303,N_7551,N_9672);
nor U12304 (N_12304,N_7728,N_9352);
and U12305 (N_12305,N_5096,N_7740);
nor U12306 (N_12306,N_5125,N_5823);
or U12307 (N_12307,N_7045,N_8079);
nand U12308 (N_12308,N_9935,N_8805);
and U12309 (N_12309,N_6372,N_7658);
and U12310 (N_12310,N_6468,N_5874);
nor U12311 (N_12311,N_5807,N_7615);
and U12312 (N_12312,N_8983,N_8464);
and U12313 (N_12313,N_6804,N_8453);
xor U12314 (N_12314,N_6461,N_5336);
nand U12315 (N_12315,N_7107,N_9134);
nand U12316 (N_12316,N_8260,N_8617);
and U12317 (N_12317,N_9689,N_8683);
nand U12318 (N_12318,N_7817,N_5280);
nor U12319 (N_12319,N_8305,N_5341);
and U12320 (N_12320,N_8540,N_9829);
nor U12321 (N_12321,N_8063,N_7648);
and U12322 (N_12322,N_8704,N_5587);
xor U12323 (N_12323,N_9730,N_8494);
nor U12324 (N_12324,N_5300,N_5191);
nor U12325 (N_12325,N_8489,N_5273);
or U12326 (N_12326,N_7181,N_5746);
nor U12327 (N_12327,N_9278,N_6108);
nand U12328 (N_12328,N_5547,N_7223);
nor U12329 (N_12329,N_7306,N_5160);
and U12330 (N_12330,N_6397,N_6393);
nand U12331 (N_12331,N_9565,N_7856);
or U12332 (N_12332,N_6188,N_6157);
nor U12333 (N_12333,N_5730,N_8303);
and U12334 (N_12334,N_7830,N_7677);
xnor U12335 (N_12335,N_6864,N_7612);
xor U12336 (N_12336,N_8583,N_9592);
nand U12337 (N_12337,N_6743,N_8875);
xor U12338 (N_12338,N_8511,N_5722);
nor U12339 (N_12339,N_6103,N_5399);
xnor U12340 (N_12340,N_5774,N_8263);
nor U12341 (N_12341,N_8501,N_9330);
xor U12342 (N_12342,N_6560,N_8289);
nor U12343 (N_12343,N_5469,N_6578);
nor U12344 (N_12344,N_6472,N_9097);
or U12345 (N_12345,N_6558,N_6464);
nand U12346 (N_12346,N_7316,N_6115);
xor U12347 (N_12347,N_7275,N_9519);
nor U12348 (N_12348,N_6884,N_7014);
nand U12349 (N_12349,N_6993,N_5083);
and U12350 (N_12350,N_8287,N_9251);
nand U12351 (N_12351,N_9157,N_9275);
xnor U12352 (N_12352,N_5935,N_9828);
nor U12353 (N_12353,N_9114,N_8759);
nand U12354 (N_12354,N_6684,N_7227);
and U12355 (N_12355,N_9593,N_5667);
or U12356 (N_12356,N_6855,N_5174);
nor U12357 (N_12357,N_5564,N_8362);
or U12358 (N_12358,N_9036,N_6524);
or U12359 (N_12359,N_6454,N_5262);
and U12360 (N_12360,N_7804,N_8005);
or U12361 (N_12361,N_5737,N_9954);
nor U12362 (N_12362,N_9346,N_9507);
xor U12363 (N_12363,N_8462,N_7514);
nor U12364 (N_12364,N_5181,N_7139);
nand U12365 (N_12365,N_9164,N_6366);
nand U12366 (N_12366,N_8514,N_9910);
nor U12367 (N_12367,N_5673,N_5063);
and U12368 (N_12368,N_9632,N_6945);
or U12369 (N_12369,N_5016,N_6689);
and U12370 (N_12370,N_8892,N_6875);
nand U12371 (N_12371,N_6727,N_7620);
and U12372 (N_12372,N_5382,N_6063);
xnor U12373 (N_12373,N_9146,N_5206);
nor U12374 (N_12374,N_6531,N_9528);
and U12375 (N_12375,N_7288,N_7791);
xor U12376 (N_12376,N_5284,N_9964);
nand U12377 (N_12377,N_8019,N_6400);
nand U12378 (N_12378,N_9208,N_8474);
nand U12379 (N_12379,N_6929,N_7021);
xor U12380 (N_12380,N_7310,N_5781);
and U12381 (N_12381,N_6008,N_9716);
xor U12382 (N_12382,N_7101,N_5391);
or U12383 (N_12383,N_5878,N_7231);
and U12384 (N_12384,N_7919,N_6067);
or U12385 (N_12385,N_9262,N_7736);
and U12386 (N_12386,N_7797,N_7141);
or U12387 (N_12387,N_5846,N_5659);
nand U12388 (N_12388,N_8212,N_7048);
or U12389 (N_12389,N_9006,N_6731);
and U12390 (N_12390,N_8936,N_6190);
nor U12391 (N_12391,N_5046,N_5697);
nand U12392 (N_12392,N_5094,N_5480);
nand U12393 (N_12393,N_5713,N_7491);
nand U12394 (N_12394,N_6533,N_7688);
nor U12395 (N_12395,N_8613,N_7650);
or U12396 (N_12396,N_8910,N_7756);
and U12397 (N_12397,N_6943,N_6355);
xor U12398 (N_12398,N_8893,N_6904);
and U12399 (N_12399,N_9057,N_6817);
or U12400 (N_12400,N_9803,N_9600);
or U12401 (N_12401,N_9605,N_5225);
or U12402 (N_12402,N_5535,N_6688);
nor U12403 (N_12403,N_6462,N_8324);
nand U12404 (N_12404,N_8755,N_6398);
or U12405 (N_12405,N_6423,N_5633);
or U12406 (N_12406,N_9327,N_6244);
nand U12407 (N_12407,N_9734,N_5997);
nand U12408 (N_12408,N_8973,N_7584);
or U12409 (N_12409,N_6289,N_7982);
or U12410 (N_12410,N_5275,N_5078);
or U12411 (N_12411,N_6502,N_6394);
nand U12412 (N_12412,N_8496,N_8826);
or U12413 (N_12413,N_8093,N_8991);
nand U12414 (N_12414,N_5804,N_9634);
and U12415 (N_12415,N_8706,N_9020);
nand U12416 (N_12416,N_7569,N_5989);
xnor U12417 (N_12417,N_8029,N_5597);
nand U12418 (N_12418,N_7379,N_7370);
nor U12419 (N_12419,N_7190,N_9655);
nand U12420 (N_12420,N_5370,N_5130);
nor U12421 (N_12421,N_7362,N_9290);
or U12422 (N_12422,N_6924,N_9552);
nand U12423 (N_12423,N_7762,N_8972);
nand U12424 (N_12424,N_9517,N_6446);
nor U12425 (N_12425,N_5329,N_9488);
nand U12426 (N_12426,N_5298,N_5783);
nand U12427 (N_12427,N_8139,N_5504);
or U12428 (N_12428,N_8539,N_6326);
nand U12429 (N_12429,N_7955,N_5200);
nand U12430 (N_12430,N_8728,N_5053);
nor U12431 (N_12431,N_6869,N_7727);
nor U12432 (N_12432,N_6829,N_5568);
and U12433 (N_12433,N_9336,N_6827);
or U12434 (N_12434,N_6495,N_9214);
nand U12435 (N_12435,N_5944,N_9219);
or U12436 (N_12436,N_5954,N_5061);
xnor U12437 (N_12437,N_6882,N_8177);
and U12438 (N_12438,N_7660,N_9826);
and U12439 (N_12439,N_6205,N_8788);
nand U12440 (N_12440,N_9998,N_6331);
and U12441 (N_12441,N_6433,N_7676);
or U12442 (N_12442,N_7152,N_7025);
or U12443 (N_12443,N_9864,N_5537);
and U12444 (N_12444,N_5309,N_6193);
nor U12445 (N_12445,N_5522,N_6509);
nor U12446 (N_12446,N_5038,N_5012);
nand U12447 (N_12447,N_5323,N_9841);
nand U12448 (N_12448,N_6656,N_5223);
xor U12449 (N_12449,N_7672,N_8899);
xor U12450 (N_12450,N_7704,N_9402);
or U12451 (N_12451,N_9381,N_7278);
nand U12452 (N_12452,N_5892,N_7824);
xor U12453 (N_12453,N_7271,N_8665);
and U12454 (N_12454,N_8884,N_9121);
or U12455 (N_12455,N_7010,N_5752);
nand U12456 (N_12456,N_9620,N_9461);
nor U12457 (N_12457,N_5543,N_9215);
or U12458 (N_12458,N_5956,N_9506);
or U12459 (N_12459,N_7690,N_9579);
nor U12460 (N_12460,N_6927,N_7440);
and U12461 (N_12461,N_6340,N_6599);
and U12462 (N_12462,N_5445,N_6978);
and U12463 (N_12463,N_9847,N_5760);
and U12464 (N_12464,N_7682,N_9682);
or U12465 (N_12465,N_5515,N_8438);
nor U12466 (N_12466,N_5763,N_6544);
nor U12467 (N_12467,N_8766,N_6263);
nor U12468 (N_12468,N_5423,N_5266);
nand U12469 (N_12469,N_7322,N_7603);
and U12470 (N_12470,N_6273,N_9027);
or U12471 (N_12471,N_7082,N_5427);
nor U12472 (N_12472,N_7832,N_5566);
nand U12473 (N_12473,N_7670,N_7862);
nor U12474 (N_12474,N_9690,N_7369);
nand U12475 (N_12475,N_9615,N_9323);
nor U12476 (N_12476,N_8982,N_6427);
and U12477 (N_12477,N_5042,N_9851);
and U12478 (N_12478,N_9744,N_5513);
xnor U12479 (N_12479,N_5732,N_8582);
or U12480 (N_12480,N_8294,N_6437);
nand U12481 (N_12481,N_8754,N_7203);
nor U12482 (N_12482,N_9184,N_5967);
nand U12483 (N_12483,N_8095,N_9988);
nand U12484 (N_12484,N_6654,N_9303);
and U12485 (N_12485,N_6805,N_9654);
nor U12486 (N_12486,N_6492,N_9599);
or U12487 (N_12487,N_9822,N_6703);
nor U12488 (N_12488,N_8891,N_9050);
or U12489 (N_12489,N_6701,N_6044);
xor U12490 (N_12490,N_8288,N_9404);
and U12491 (N_12491,N_6726,N_6348);
nand U12492 (N_12492,N_6795,N_7385);
and U12493 (N_12493,N_7256,N_6574);
nand U12494 (N_12494,N_6042,N_7097);
nand U12495 (N_12495,N_9576,N_7885);
and U12496 (N_12496,N_5514,N_7751);
nor U12497 (N_12497,N_6185,N_5436);
and U12498 (N_12498,N_5593,N_5140);
and U12499 (N_12499,N_8215,N_6285);
and U12500 (N_12500,N_8310,N_6842);
or U12501 (N_12501,N_9655,N_6845);
or U12502 (N_12502,N_9597,N_6192);
xnor U12503 (N_12503,N_5006,N_9716);
and U12504 (N_12504,N_5463,N_5481);
and U12505 (N_12505,N_9601,N_8333);
and U12506 (N_12506,N_8769,N_9362);
nor U12507 (N_12507,N_9237,N_7949);
nor U12508 (N_12508,N_5544,N_9891);
nand U12509 (N_12509,N_9141,N_5996);
xor U12510 (N_12510,N_7831,N_9517);
or U12511 (N_12511,N_9901,N_8052);
nand U12512 (N_12512,N_9159,N_7949);
nand U12513 (N_12513,N_5700,N_6544);
nor U12514 (N_12514,N_7157,N_8144);
or U12515 (N_12515,N_8593,N_6410);
nand U12516 (N_12516,N_9712,N_5664);
nor U12517 (N_12517,N_8058,N_7743);
nand U12518 (N_12518,N_9049,N_8860);
xor U12519 (N_12519,N_9540,N_5845);
nand U12520 (N_12520,N_8766,N_6389);
xor U12521 (N_12521,N_8170,N_6221);
or U12522 (N_12522,N_6942,N_9542);
nor U12523 (N_12523,N_6059,N_8119);
xor U12524 (N_12524,N_6524,N_9010);
nor U12525 (N_12525,N_5666,N_5211);
xnor U12526 (N_12526,N_9187,N_8129);
or U12527 (N_12527,N_5015,N_9976);
nand U12528 (N_12528,N_7233,N_9083);
nand U12529 (N_12529,N_9834,N_5569);
and U12530 (N_12530,N_7832,N_8698);
nor U12531 (N_12531,N_9686,N_8938);
nor U12532 (N_12532,N_7071,N_9377);
nor U12533 (N_12533,N_6101,N_7237);
nand U12534 (N_12534,N_9105,N_7895);
nor U12535 (N_12535,N_7755,N_5742);
or U12536 (N_12536,N_6582,N_6411);
and U12537 (N_12537,N_6476,N_8573);
and U12538 (N_12538,N_7237,N_8206);
and U12539 (N_12539,N_9056,N_6944);
or U12540 (N_12540,N_7449,N_7441);
nor U12541 (N_12541,N_7890,N_5449);
xnor U12542 (N_12542,N_8906,N_6389);
and U12543 (N_12543,N_8731,N_5603);
nor U12544 (N_12544,N_6685,N_5053);
and U12545 (N_12545,N_8568,N_6651);
nor U12546 (N_12546,N_7794,N_5134);
nor U12547 (N_12547,N_8112,N_7655);
and U12548 (N_12548,N_5971,N_9546);
nand U12549 (N_12549,N_5748,N_6148);
xor U12550 (N_12550,N_6029,N_5104);
and U12551 (N_12551,N_5906,N_5225);
xor U12552 (N_12552,N_6079,N_9769);
nor U12553 (N_12553,N_8639,N_9935);
nor U12554 (N_12554,N_9612,N_6696);
nand U12555 (N_12555,N_7643,N_9541);
or U12556 (N_12556,N_7319,N_6858);
nand U12557 (N_12557,N_9891,N_8474);
xnor U12558 (N_12558,N_8457,N_6773);
nand U12559 (N_12559,N_9637,N_6260);
nor U12560 (N_12560,N_9812,N_6168);
xor U12561 (N_12561,N_7462,N_9389);
nand U12562 (N_12562,N_6718,N_7206);
nand U12563 (N_12563,N_6452,N_5361);
or U12564 (N_12564,N_8027,N_5195);
or U12565 (N_12565,N_8139,N_8351);
and U12566 (N_12566,N_8414,N_6902);
xnor U12567 (N_12567,N_5097,N_9760);
xnor U12568 (N_12568,N_6788,N_7148);
nor U12569 (N_12569,N_7686,N_9215);
nand U12570 (N_12570,N_6623,N_9695);
nand U12571 (N_12571,N_9777,N_8741);
or U12572 (N_12572,N_7606,N_5999);
nand U12573 (N_12573,N_5343,N_7275);
and U12574 (N_12574,N_6245,N_6500);
nand U12575 (N_12575,N_7664,N_7820);
xnor U12576 (N_12576,N_9241,N_8225);
nand U12577 (N_12577,N_5719,N_7625);
nand U12578 (N_12578,N_5389,N_5860);
and U12579 (N_12579,N_7657,N_7681);
nor U12580 (N_12580,N_9853,N_5508);
xor U12581 (N_12581,N_9454,N_8417);
nand U12582 (N_12582,N_9807,N_7753);
and U12583 (N_12583,N_6142,N_6492);
nand U12584 (N_12584,N_9672,N_7232);
or U12585 (N_12585,N_9487,N_9475);
and U12586 (N_12586,N_6875,N_6127);
nor U12587 (N_12587,N_7127,N_8744);
and U12588 (N_12588,N_7986,N_9555);
nand U12589 (N_12589,N_7724,N_7678);
or U12590 (N_12590,N_8587,N_8425);
nand U12591 (N_12591,N_5567,N_6552);
or U12592 (N_12592,N_6627,N_7494);
or U12593 (N_12593,N_5090,N_8218);
nand U12594 (N_12594,N_5402,N_6764);
nand U12595 (N_12595,N_5626,N_8451);
or U12596 (N_12596,N_9530,N_6020);
nor U12597 (N_12597,N_8726,N_8972);
or U12598 (N_12598,N_5855,N_8795);
xor U12599 (N_12599,N_8422,N_9698);
or U12600 (N_12600,N_9979,N_6714);
or U12601 (N_12601,N_7679,N_5370);
nand U12602 (N_12602,N_7469,N_9425);
or U12603 (N_12603,N_8785,N_5014);
nor U12604 (N_12604,N_8476,N_5032);
nand U12605 (N_12605,N_7774,N_6296);
nor U12606 (N_12606,N_7106,N_7814);
nand U12607 (N_12607,N_6153,N_6630);
nand U12608 (N_12608,N_9649,N_9225);
and U12609 (N_12609,N_6971,N_8604);
nor U12610 (N_12610,N_5127,N_9699);
and U12611 (N_12611,N_9496,N_8379);
xnor U12612 (N_12612,N_9022,N_9675);
xnor U12613 (N_12613,N_9471,N_5721);
xor U12614 (N_12614,N_9610,N_9420);
nor U12615 (N_12615,N_8355,N_6224);
and U12616 (N_12616,N_8743,N_5281);
nor U12617 (N_12617,N_7066,N_5248);
nor U12618 (N_12618,N_6662,N_7466);
or U12619 (N_12619,N_5686,N_5472);
xor U12620 (N_12620,N_9760,N_8977);
nand U12621 (N_12621,N_7957,N_7096);
nand U12622 (N_12622,N_8705,N_8853);
nand U12623 (N_12623,N_9670,N_5363);
xor U12624 (N_12624,N_5577,N_6108);
nand U12625 (N_12625,N_9611,N_5866);
nor U12626 (N_12626,N_8930,N_6947);
or U12627 (N_12627,N_7663,N_5433);
or U12628 (N_12628,N_6792,N_6110);
or U12629 (N_12629,N_9438,N_6366);
and U12630 (N_12630,N_5466,N_5824);
and U12631 (N_12631,N_9236,N_5234);
nand U12632 (N_12632,N_5456,N_6254);
nor U12633 (N_12633,N_8608,N_7394);
and U12634 (N_12634,N_6892,N_7697);
or U12635 (N_12635,N_8523,N_9446);
nor U12636 (N_12636,N_6395,N_5648);
or U12637 (N_12637,N_6062,N_6099);
or U12638 (N_12638,N_8767,N_8209);
nor U12639 (N_12639,N_6835,N_8948);
xor U12640 (N_12640,N_9906,N_8001);
nand U12641 (N_12641,N_8815,N_7024);
nand U12642 (N_12642,N_9121,N_9698);
nand U12643 (N_12643,N_5426,N_5034);
nor U12644 (N_12644,N_6812,N_8276);
and U12645 (N_12645,N_5582,N_6990);
nand U12646 (N_12646,N_6624,N_9483);
or U12647 (N_12647,N_9680,N_6008);
nand U12648 (N_12648,N_9696,N_9738);
nand U12649 (N_12649,N_5648,N_7418);
and U12650 (N_12650,N_6060,N_5064);
and U12651 (N_12651,N_7081,N_8102);
or U12652 (N_12652,N_9122,N_6131);
or U12653 (N_12653,N_9570,N_8460);
nand U12654 (N_12654,N_6982,N_9939);
and U12655 (N_12655,N_9556,N_6607);
nor U12656 (N_12656,N_7621,N_8525);
nand U12657 (N_12657,N_6077,N_7800);
nand U12658 (N_12658,N_6940,N_8038);
and U12659 (N_12659,N_8769,N_6220);
and U12660 (N_12660,N_8345,N_7607);
nor U12661 (N_12661,N_7820,N_8930);
or U12662 (N_12662,N_9394,N_8160);
nand U12663 (N_12663,N_9249,N_6752);
nand U12664 (N_12664,N_6283,N_6034);
nand U12665 (N_12665,N_5290,N_5704);
or U12666 (N_12666,N_8321,N_9291);
xnor U12667 (N_12667,N_8920,N_6331);
nand U12668 (N_12668,N_5236,N_5649);
nor U12669 (N_12669,N_7617,N_7959);
nand U12670 (N_12670,N_7773,N_7139);
and U12671 (N_12671,N_9868,N_5485);
or U12672 (N_12672,N_9152,N_8732);
and U12673 (N_12673,N_8090,N_8945);
and U12674 (N_12674,N_6105,N_9600);
and U12675 (N_12675,N_7249,N_5064);
or U12676 (N_12676,N_8281,N_6602);
nand U12677 (N_12677,N_8556,N_5349);
or U12678 (N_12678,N_6510,N_6069);
nand U12679 (N_12679,N_7229,N_5392);
nand U12680 (N_12680,N_6798,N_9129);
or U12681 (N_12681,N_7081,N_6792);
nand U12682 (N_12682,N_8520,N_8974);
nor U12683 (N_12683,N_9163,N_8932);
and U12684 (N_12684,N_8557,N_9864);
nand U12685 (N_12685,N_8577,N_7502);
nor U12686 (N_12686,N_5557,N_8884);
or U12687 (N_12687,N_9936,N_7093);
and U12688 (N_12688,N_5961,N_6578);
nor U12689 (N_12689,N_5138,N_7926);
nand U12690 (N_12690,N_9119,N_8908);
nand U12691 (N_12691,N_5641,N_5325);
nand U12692 (N_12692,N_7219,N_8953);
and U12693 (N_12693,N_9110,N_7272);
and U12694 (N_12694,N_5046,N_9038);
nor U12695 (N_12695,N_5726,N_8921);
nand U12696 (N_12696,N_8819,N_7332);
or U12697 (N_12697,N_5073,N_6564);
nor U12698 (N_12698,N_8399,N_9281);
nand U12699 (N_12699,N_9009,N_6711);
and U12700 (N_12700,N_6194,N_6018);
or U12701 (N_12701,N_5048,N_5763);
nand U12702 (N_12702,N_8351,N_5571);
nor U12703 (N_12703,N_9231,N_8892);
or U12704 (N_12704,N_8204,N_8363);
nor U12705 (N_12705,N_6373,N_8792);
nor U12706 (N_12706,N_6413,N_5759);
nand U12707 (N_12707,N_5839,N_7592);
nor U12708 (N_12708,N_9469,N_5513);
and U12709 (N_12709,N_9154,N_8826);
nor U12710 (N_12710,N_7517,N_6971);
nor U12711 (N_12711,N_6455,N_7175);
nor U12712 (N_12712,N_7755,N_6146);
and U12713 (N_12713,N_8864,N_6197);
or U12714 (N_12714,N_6587,N_8976);
and U12715 (N_12715,N_7429,N_5314);
and U12716 (N_12716,N_8575,N_6008);
nand U12717 (N_12717,N_6600,N_9552);
nor U12718 (N_12718,N_6758,N_5619);
nand U12719 (N_12719,N_6993,N_5753);
or U12720 (N_12720,N_7353,N_5748);
xor U12721 (N_12721,N_5252,N_7052);
nor U12722 (N_12722,N_5328,N_8946);
or U12723 (N_12723,N_8910,N_5715);
or U12724 (N_12724,N_5324,N_7739);
nor U12725 (N_12725,N_6733,N_8290);
nor U12726 (N_12726,N_5562,N_8058);
nor U12727 (N_12727,N_7847,N_9726);
nand U12728 (N_12728,N_9341,N_8285);
xnor U12729 (N_12729,N_9187,N_9625);
nand U12730 (N_12730,N_9941,N_5387);
or U12731 (N_12731,N_7531,N_8244);
or U12732 (N_12732,N_6971,N_8811);
and U12733 (N_12733,N_7391,N_7421);
or U12734 (N_12734,N_6227,N_7778);
and U12735 (N_12735,N_8673,N_6301);
nor U12736 (N_12736,N_8798,N_9966);
nand U12737 (N_12737,N_8103,N_8772);
xnor U12738 (N_12738,N_5413,N_9753);
or U12739 (N_12739,N_5281,N_5757);
and U12740 (N_12740,N_5782,N_9499);
or U12741 (N_12741,N_7996,N_5194);
and U12742 (N_12742,N_7035,N_6848);
nor U12743 (N_12743,N_7851,N_8709);
or U12744 (N_12744,N_7802,N_8444);
nand U12745 (N_12745,N_8243,N_9101);
xor U12746 (N_12746,N_7825,N_9974);
and U12747 (N_12747,N_8653,N_9678);
nor U12748 (N_12748,N_5044,N_9978);
xor U12749 (N_12749,N_9391,N_6413);
nand U12750 (N_12750,N_5953,N_5808);
or U12751 (N_12751,N_6230,N_5505);
xnor U12752 (N_12752,N_6724,N_6287);
xor U12753 (N_12753,N_5184,N_7175);
nand U12754 (N_12754,N_8910,N_5143);
nor U12755 (N_12755,N_7193,N_7395);
nor U12756 (N_12756,N_7778,N_7264);
and U12757 (N_12757,N_6563,N_5562);
and U12758 (N_12758,N_5683,N_6414);
or U12759 (N_12759,N_7448,N_7135);
or U12760 (N_12760,N_6891,N_9105);
nand U12761 (N_12761,N_5911,N_8775);
and U12762 (N_12762,N_5456,N_7849);
nor U12763 (N_12763,N_9535,N_7258);
xor U12764 (N_12764,N_5182,N_6911);
nand U12765 (N_12765,N_9152,N_5695);
and U12766 (N_12766,N_5406,N_7713);
or U12767 (N_12767,N_5838,N_8272);
and U12768 (N_12768,N_7568,N_9281);
nor U12769 (N_12769,N_8909,N_9861);
or U12770 (N_12770,N_8742,N_7074);
xor U12771 (N_12771,N_7904,N_9450);
and U12772 (N_12772,N_7622,N_9821);
nor U12773 (N_12773,N_6737,N_5365);
nor U12774 (N_12774,N_8431,N_9859);
or U12775 (N_12775,N_9372,N_6574);
or U12776 (N_12776,N_9471,N_6456);
nor U12777 (N_12777,N_8859,N_7588);
nor U12778 (N_12778,N_7814,N_9337);
nor U12779 (N_12779,N_8554,N_9344);
nand U12780 (N_12780,N_5060,N_9678);
nand U12781 (N_12781,N_7681,N_5343);
or U12782 (N_12782,N_9304,N_7815);
xor U12783 (N_12783,N_8375,N_6851);
nand U12784 (N_12784,N_5003,N_5816);
nor U12785 (N_12785,N_9762,N_7058);
nand U12786 (N_12786,N_5403,N_5637);
or U12787 (N_12787,N_6046,N_6580);
or U12788 (N_12788,N_7210,N_9976);
or U12789 (N_12789,N_8992,N_6014);
and U12790 (N_12790,N_8654,N_6385);
nand U12791 (N_12791,N_7233,N_8207);
nor U12792 (N_12792,N_5457,N_6751);
and U12793 (N_12793,N_8693,N_6702);
or U12794 (N_12794,N_9180,N_9386);
or U12795 (N_12795,N_7893,N_6324);
or U12796 (N_12796,N_5531,N_5952);
and U12797 (N_12797,N_5021,N_9774);
nor U12798 (N_12798,N_5527,N_5373);
nor U12799 (N_12799,N_9056,N_6192);
nand U12800 (N_12800,N_7131,N_9771);
or U12801 (N_12801,N_8438,N_8053);
nor U12802 (N_12802,N_7794,N_8234);
nand U12803 (N_12803,N_9796,N_6632);
and U12804 (N_12804,N_5557,N_9174);
and U12805 (N_12805,N_5737,N_5307);
nor U12806 (N_12806,N_6949,N_9600);
nand U12807 (N_12807,N_8902,N_7675);
and U12808 (N_12808,N_8356,N_7798);
xnor U12809 (N_12809,N_8267,N_6831);
nand U12810 (N_12810,N_8835,N_7343);
and U12811 (N_12811,N_9959,N_5400);
and U12812 (N_12812,N_6043,N_5931);
and U12813 (N_12813,N_5470,N_8789);
or U12814 (N_12814,N_6356,N_7306);
xor U12815 (N_12815,N_8228,N_8896);
and U12816 (N_12816,N_8773,N_7778);
nor U12817 (N_12817,N_6078,N_7418);
and U12818 (N_12818,N_6798,N_8714);
nand U12819 (N_12819,N_9609,N_9822);
or U12820 (N_12820,N_6549,N_5664);
and U12821 (N_12821,N_9605,N_8296);
nor U12822 (N_12822,N_7261,N_9019);
or U12823 (N_12823,N_9416,N_9086);
or U12824 (N_12824,N_8710,N_6798);
or U12825 (N_12825,N_9273,N_6366);
xor U12826 (N_12826,N_8457,N_7107);
nor U12827 (N_12827,N_9585,N_6782);
nand U12828 (N_12828,N_5939,N_9757);
and U12829 (N_12829,N_8769,N_5033);
and U12830 (N_12830,N_6265,N_9901);
and U12831 (N_12831,N_5789,N_8691);
nand U12832 (N_12832,N_7546,N_5338);
nor U12833 (N_12833,N_7535,N_9601);
nand U12834 (N_12834,N_8518,N_9531);
nand U12835 (N_12835,N_9138,N_6280);
nand U12836 (N_12836,N_8496,N_7630);
nand U12837 (N_12837,N_8063,N_6197);
or U12838 (N_12838,N_6194,N_7080);
and U12839 (N_12839,N_9164,N_5789);
nand U12840 (N_12840,N_7809,N_7636);
nor U12841 (N_12841,N_9825,N_6632);
and U12842 (N_12842,N_5638,N_6711);
or U12843 (N_12843,N_5733,N_7031);
nor U12844 (N_12844,N_5661,N_6565);
nor U12845 (N_12845,N_7207,N_7226);
nor U12846 (N_12846,N_9042,N_7663);
xor U12847 (N_12847,N_8449,N_5217);
or U12848 (N_12848,N_8686,N_7334);
xnor U12849 (N_12849,N_5181,N_6665);
and U12850 (N_12850,N_8734,N_5926);
nand U12851 (N_12851,N_9838,N_5825);
xor U12852 (N_12852,N_6294,N_5297);
xor U12853 (N_12853,N_6665,N_5319);
and U12854 (N_12854,N_6982,N_6292);
nand U12855 (N_12855,N_6399,N_8787);
xnor U12856 (N_12856,N_9528,N_9324);
nor U12857 (N_12857,N_5016,N_5391);
nor U12858 (N_12858,N_9974,N_6777);
nor U12859 (N_12859,N_8919,N_5169);
or U12860 (N_12860,N_7144,N_8554);
or U12861 (N_12861,N_9824,N_9338);
or U12862 (N_12862,N_5164,N_7071);
and U12863 (N_12863,N_7839,N_9002);
and U12864 (N_12864,N_6439,N_6343);
nor U12865 (N_12865,N_8954,N_9801);
nor U12866 (N_12866,N_5573,N_7526);
nor U12867 (N_12867,N_9603,N_9819);
nor U12868 (N_12868,N_5946,N_8314);
xnor U12869 (N_12869,N_8196,N_6323);
xor U12870 (N_12870,N_6930,N_8778);
or U12871 (N_12871,N_7691,N_8453);
and U12872 (N_12872,N_7162,N_6458);
nor U12873 (N_12873,N_6789,N_7702);
and U12874 (N_12874,N_9732,N_6447);
or U12875 (N_12875,N_8330,N_7840);
nor U12876 (N_12876,N_9333,N_8436);
and U12877 (N_12877,N_9498,N_6811);
and U12878 (N_12878,N_5125,N_6322);
nor U12879 (N_12879,N_7564,N_9557);
or U12880 (N_12880,N_9217,N_7698);
and U12881 (N_12881,N_7099,N_9057);
xnor U12882 (N_12882,N_7912,N_7103);
xor U12883 (N_12883,N_8307,N_8560);
nand U12884 (N_12884,N_7838,N_9355);
nand U12885 (N_12885,N_9618,N_6901);
nand U12886 (N_12886,N_9774,N_9777);
or U12887 (N_12887,N_6290,N_7554);
nor U12888 (N_12888,N_5927,N_9732);
xor U12889 (N_12889,N_5685,N_8624);
and U12890 (N_12890,N_6541,N_5099);
and U12891 (N_12891,N_8128,N_6586);
nand U12892 (N_12892,N_8934,N_8763);
nor U12893 (N_12893,N_9076,N_8714);
or U12894 (N_12894,N_8963,N_8223);
nand U12895 (N_12895,N_6160,N_9790);
and U12896 (N_12896,N_5882,N_8809);
or U12897 (N_12897,N_9106,N_5924);
nand U12898 (N_12898,N_7755,N_9025);
xor U12899 (N_12899,N_9954,N_5752);
nor U12900 (N_12900,N_8532,N_7734);
and U12901 (N_12901,N_6236,N_9140);
nand U12902 (N_12902,N_6459,N_6754);
xor U12903 (N_12903,N_6787,N_9824);
xnor U12904 (N_12904,N_6492,N_7110);
or U12905 (N_12905,N_8954,N_6905);
nand U12906 (N_12906,N_8619,N_5055);
nand U12907 (N_12907,N_6640,N_5639);
or U12908 (N_12908,N_8784,N_8521);
and U12909 (N_12909,N_7644,N_8123);
nor U12910 (N_12910,N_6893,N_5565);
and U12911 (N_12911,N_8295,N_8302);
and U12912 (N_12912,N_5605,N_8802);
nor U12913 (N_12913,N_5985,N_9129);
nor U12914 (N_12914,N_9130,N_6709);
nand U12915 (N_12915,N_9855,N_8814);
and U12916 (N_12916,N_7226,N_5342);
nand U12917 (N_12917,N_8139,N_9000);
or U12918 (N_12918,N_8575,N_9678);
and U12919 (N_12919,N_7731,N_5108);
or U12920 (N_12920,N_5924,N_6414);
nor U12921 (N_12921,N_7296,N_8525);
or U12922 (N_12922,N_5395,N_8581);
and U12923 (N_12923,N_9807,N_5550);
or U12924 (N_12924,N_7893,N_7448);
xor U12925 (N_12925,N_9231,N_6853);
xnor U12926 (N_12926,N_5833,N_5006);
nor U12927 (N_12927,N_9098,N_5849);
or U12928 (N_12928,N_5436,N_6925);
or U12929 (N_12929,N_8855,N_7989);
nand U12930 (N_12930,N_5207,N_6434);
xor U12931 (N_12931,N_5813,N_9866);
nand U12932 (N_12932,N_8194,N_5876);
and U12933 (N_12933,N_9873,N_6563);
nor U12934 (N_12934,N_7000,N_6272);
nor U12935 (N_12935,N_9243,N_6788);
and U12936 (N_12936,N_7831,N_6268);
and U12937 (N_12937,N_7932,N_9944);
nor U12938 (N_12938,N_8379,N_9338);
nor U12939 (N_12939,N_6957,N_6530);
xnor U12940 (N_12940,N_8703,N_8063);
nor U12941 (N_12941,N_7311,N_9057);
nor U12942 (N_12942,N_7445,N_6826);
xor U12943 (N_12943,N_9002,N_8852);
nor U12944 (N_12944,N_7847,N_9335);
and U12945 (N_12945,N_6559,N_8786);
or U12946 (N_12946,N_5803,N_5190);
nand U12947 (N_12947,N_5131,N_5905);
nand U12948 (N_12948,N_9802,N_8890);
or U12949 (N_12949,N_8200,N_9079);
nand U12950 (N_12950,N_8934,N_8474);
nand U12951 (N_12951,N_5360,N_7578);
nor U12952 (N_12952,N_8449,N_6223);
nor U12953 (N_12953,N_8320,N_5871);
nor U12954 (N_12954,N_9559,N_8655);
xnor U12955 (N_12955,N_9971,N_9358);
or U12956 (N_12956,N_7647,N_8816);
nor U12957 (N_12957,N_6990,N_6677);
nor U12958 (N_12958,N_9616,N_8662);
xor U12959 (N_12959,N_8849,N_9759);
and U12960 (N_12960,N_8916,N_5265);
xor U12961 (N_12961,N_7126,N_7955);
nand U12962 (N_12962,N_5715,N_9939);
nand U12963 (N_12963,N_5630,N_5219);
nand U12964 (N_12964,N_6734,N_9717);
nand U12965 (N_12965,N_8644,N_7136);
and U12966 (N_12966,N_6033,N_7774);
xnor U12967 (N_12967,N_5692,N_9807);
nand U12968 (N_12968,N_9744,N_5462);
and U12969 (N_12969,N_5563,N_9886);
and U12970 (N_12970,N_5023,N_5173);
and U12971 (N_12971,N_6886,N_7961);
and U12972 (N_12972,N_5872,N_5483);
nand U12973 (N_12973,N_7122,N_7761);
and U12974 (N_12974,N_7099,N_6825);
nand U12975 (N_12975,N_8128,N_6635);
and U12976 (N_12976,N_9614,N_9775);
nand U12977 (N_12977,N_9240,N_6211);
nor U12978 (N_12978,N_9150,N_8988);
nor U12979 (N_12979,N_6635,N_5100);
nand U12980 (N_12980,N_8341,N_9735);
nand U12981 (N_12981,N_6555,N_6083);
nor U12982 (N_12982,N_7521,N_5338);
or U12983 (N_12983,N_8740,N_5518);
nor U12984 (N_12984,N_9468,N_6358);
nor U12985 (N_12985,N_8588,N_7592);
and U12986 (N_12986,N_6776,N_7317);
nor U12987 (N_12987,N_8608,N_7960);
or U12988 (N_12988,N_7175,N_5666);
or U12989 (N_12989,N_8931,N_9077);
nor U12990 (N_12990,N_8703,N_6736);
nor U12991 (N_12991,N_9716,N_6924);
or U12992 (N_12992,N_7750,N_9389);
nand U12993 (N_12993,N_6783,N_5284);
or U12994 (N_12994,N_7998,N_8094);
and U12995 (N_12995,N_6950,N_5255);
and U12996 (N_12996,N_6019,N_9733);
and U12997 (N_12997,N_9054,N_7068);
and U12998 (N_12998,N_7878,N_6194);
or U12999 (N_12999,N_9005,N_5540);
or U13000 (N_13000,N_6542,N_8310);
nor U13001 (N_13001,N_9945,N_7658);
nor U13002 (N_13002,N_7648,N_7743);
xor U13003 (N_13003,N_7935,N_7144);
xor U13004 (N_13004,N_6763,N_5004);
nand U13005 (N_13005,N_6741,N_9400);
nand U13006 (N_13006,N_5115,N_8879);
or U13007 (N_13007,N_5516,N_9949);
nand U13008 (N_13008,N_7005,N_9914);
nor U13009 (N_13009,N_6203,N_5475);
nor U13010 (N_13010,N_8838,N_5370);
nor U13011 (N_13011,N_5056,N_5233);
nor U13012 (N_13012,N_5753,N_9578);
or U13013 (N_13013,N_9348,N_8199);
and U13014 (N_13014,N_7913,N_7484);
or U13015 (N_13015,N_9900,N_7173);
nor U13016 (N_13016,N_8746,N_9176);
nand U13017 (N_13017,N_8394,N_9464);
or U13018 (N_13018,N_8492,N_5753);
or U13019 (N_13019,N_6627,N_8339);
xor U13020 (N_13020,N_8657,N_6666);
nor U13021 (N_13021,N_6887,N_8259);
and U13022 (N_13022,N_8548,N_8555);
and U13023 (N_13023,N_7387,N_9407);
nand U13024 (N_13024,N_7971,N_6105);
nand U13025 (N_13025,N_7909,N_9307);
xnor U13026 (N_13026,N_7239,N_6336);
or U13027 (N_13027,N_7475,N_5907);
nand U13028 (N_13028,N_6164,N_9618);
or U13029 (N_13029,N_7206,N_5698);
nor U13030 (N_13030,N_9652,N_9325);
or U13031 (N_13031,N_5166,N_6033);
and U13032 (N_13032,N_5689,N_9521);
nor U13033 (N_13033,N_6131,N_8569);
nor U13034 (N_13034,N_5921,N_7659);
nor U13035 (N_13035,N_9619,N_5654);
and U13036 (N_13036,N_7479,N_6570);
xor U13037 (N_13037,N_7862,N_8218);
and U13038 (N_13038,N_5453,N_8273);
nand U13039 (N_13039,N_7118,N_6206);
nand U13040 (N_13040,N_6679,N_6750);
or U13041 (N_13041,N_5295,N_6282);
or U13042 (N_13042,N_5300,N_5877);
nand U13043 (N_13043,N_7689,N_7778);
xor U13044 (N_13044,N_5440,N_7527);
nand U13045 (N_13045,N_9962,N_8765);
or U13046 (N_13046,N_7949,N_8659);
and U13047 (N_13047,N_9233,N_5950);
nand U13048 (N_13048,N_8258,N_6131);
nor U13049 (N_13049,N_8641,N_6637);
nand U13050 (N_13050,N_7866,N_6855);
nor U13051 (N_13051,N_6368,N_6292);
and U13052 (N_13052,N_5859,N_5620);
nand U13053 (N_13053,N_6062,N_9181);
xor U13054 (N_13054,N_6215,N_5465);
nand U13055 (N_13055,N_9468,N_9967);
nand U13056 (N_13056,N_9182,N_5604);
nand U13057 (N_13057,N_5872,N_6215);
nor U13058 (N_13058,N_7702,N_7984);
nor U13059 (N_13059,N_6255,N_6322);
or U13060 (N_13060,N_6704,N_5429);
nor U13061 (N_13061,N_8747,N_8466);
or U13062 (N_13062,N_9306,N_9434);
and U13063 (N_13063,N_8983,N_7457);
or U13064 (N_13064,N_5521,N_5295);
nor U13065 (N_13065,N_6526,N_7008);
and U13066 (N_13066,N_5993,N_5772);
and U13067 (N_13067,N_9767,N_8409);
nand U13068 (N_13068,N_7600,N_9937);
or U13069 (N_13069,N_8326,N_9386);
nand U13070 (N_13070,N_8532,N_8332);
nand U13071 (N_13071,N_9624,N_6117);
nand U13072 (N_13072,N_8521,N_7487);
nand U13073 (N_13073,N_5712,N_9019);
and U13074 (N_13074,N_9792,N_7829);
or U13075 (N_13075,N_5324,N_5750);
or U13076 (N_13076,N_9652,N_9614);
or U13077 (N_13077,N_6581,N_6995);
nand U13078 (N_13078,N_7600,N_7891);
nand U13079 (N_13079,N_6752,N_8080);
nand U13080 (N_13080,N_5816,N_5758);
xnor U13081 (N_13081,N_5639,N_5955);
and U13082 (N_13082,N_5488,N_7219);
nor U13083 (N_13083,N_5626,N_9234);
nor U13084 (N_13084,N_8887,N_7491);
xnor U13085 (N_13085,N_6304,N_5212);
and U13086 (N_13086,N_7731,N_5734);
nand U13087 (N_13087,N_9126,N_5366);
nor U13088 (N_13088,N_8668,N_7793);
and U13089 (N_13089,N_8413,N_5598);
nand U13090 (N_13090,N_5521,N_6286);
nor U13091 (N_13091,N_9132,N_8235);
nor U13092 (N_13092,N_5176,N_8298);
and U13093 (N_13093,N_5457,N_8734);
or U13094 (N_13094,N_9025,N_6105);
nor U13095 (N_13095,N_9256,N_7143);
nand U13096 (N_13096,N_8648,N_8660);
and U13097 (N_13097,N_8887,N_7377);
and U13098 (N_13098,N_6552,N_5602);
nor U13099 (N_13099,N_6526,N_8630);
and U13100 (N_13100,N_5801,N_5719);
nor U13101 (N_13101,N_9565,N_7677);
or U13102 (N_13102,N_6748,N_9256);
and U13103 (N_13103,N_9351,N_6700);
nand U13104 (N_13104,N_8116,N_9692);
xor U13105 (N_13105,N_7450,N_5368);
nand U13106 (N_13106,N_7172,N_5936);
nor U13107 (N_13107,N_8259,N_6298);
xnor U13108 (N_13108,N_6131,N_5500);
nor U13109 (N_13109,N_5242,N_6322);
and U13110 (N_13110,N_9293,N_7252);
and U13111 (N_13111,N_5621,N_7021);
nand U13112 (N_13112,N_5325,N_5190);
nand U13113 (N_13113,N_8709,N_7515);
or U13114 (N_13114,N_6181,N_8292);
or U13115 (N_13115,N_9611,N_8022);
nand U13116 (N_13116,N_6425,N_9045);
nand U13117 (N_13117,N_5741,N_5819);
and U13118 (N_13118,N_7186,N_8381);
nor U13119 (N_13119,N_9500,N_5722);
or U13120 (N_13120,N_5681,N_5409);
nor U13121 (N_13121,N_7468,N_6834);
and U13122 (N_13122,N_8230,N_7137);
nand U13123 (N_13123,N_8981,N_7485);
xor U13124 (N_13124,N_8809,N_5674);
nand U13125 (N_13125,N_8207,N_6918);
or U13126 (N_13126,N_6276,N_8801);
and U13127 (N_13127,N_9824,N_7676);
or U13128 (N_13128,N_5635,N_7989);
nand U13129 (N_13129,N_7428,N_8420);
and U13130 (N_13130,N_7728,N_8680);
nand U13131 (N_13131,N_7249,N_7695);
and U13132 (N_13132,N_6072,N_8328);
nand U13133 (N_13133,N_6271,N_7842);
and U13134 (N_13134,N_9536,N_7022);
xor U13135 (N_13135,N_6680,N_5525);
nand U13136 (N_13136,N_5910,N_9080);
or U13137 (N_13137,N_8358,N_9953);
nand U13138 (N_13138,N_7462,N_7762);
xor U13139 (N_13139,N_9229,N_5422);
and U13140 (N_13140,N_8416,N_6786);
or U13141 (N_13141,N_9054,N_5899);
nor U13142 (N_13142,N_9639,N_8368);
or U13143 (N_13143,N_5489,N_5157);
xor U13144 (N_13144,N_6255,N_7661);
and U13145 (N_13145,N_6254,N_9162);
nand U13146 (N_13146,N_9531,N_5735);
or U13147 (N_13147,N_9471,N_7106);
nand U13148 (N_13148,N_5891,N_8881);
nand U13149 (N_13149,N_9491,N_5586);
nand U13150 (N_13150,N_7754,N_6780);
and U13151 (N_13151,N_6238,N_5271);
nor U13152 (N_13152,N_7073,N_8819);
and U13153 (N_13153,N_5804,N_5956);
nor U13154 (N_13154,N_5953,N_6225);
nor U13155 (N_13155,N_5491,N_9006);
or U13156 (N_13156,N_5594,N_9849);
nor U13157 (N_13157,N_6150,N_8208);
and U13158 (N_13158,N_6914,N_5109);
nand U13159 (N_13159,N_8455,N_7867);
nand U13160 (N_13160,N_8239,N_8992);
nand U13161 (N_13161,N_6880,N_6242);
xor U13162 (N_13162,N_8734,N_8284);
nor U13163 (N_13163,N_6837,N_5066);
and U13164 (N_13164,N_5163,N_8329);
nand U13165 (N_13165,N_7368,N_6058);
nor U13166 (N_13166,N_5958,N_5752);
or U13167 (N_13167,N_5799,N_7698);
nand U13168 (N_13168,N_5673,N_8467);
or U13169 (N_13169,N_5302,N_9386);
nor U13170 (N_13170,N_8831,N_6099);
nor U13171 (N_13171,N_6707,N_6215);
nor U13172 (N_13172,N_8579,N_7391);
and U13173 (N_13173,N_7781,N_8709);
or U13174 (N_13174,N_9813,N_8619);
and U13175 (N_13175,N_5744,N_9619);
or U13176 (N_13176,N_6149,N_7852);
or U13177 (N_13177,N_8013,N_6277);
or U13178 (N_13178,N_5462,N_8503);
nand U13179 (N_13179,N_5384,N_6739);
and U13180 (N_13180,N_7469,N_6643);
and U13181 (N_13181,N_8243,N_6630);
or U13182 (N_13182,N_8640,N_5997);
nand U13183 (N_13183,N_8535,N_7609);
or U13184 (N_13184,N_8871,N_8694);
or U13185 (N_13185,N_5459,N_9642);
xor U13186 (N_13186,N_7522,N_6100);
and U13187 (N_13187,N_6551,N_5664);
nor U13188 (N_13188,N_8049,N_5752);
or U13189 (N_13189,N_9113,N_8094);
nand U13190 (N_13190,N_8605,N_6376);
and U13191 (N_13191,N_7362,N_5788);
nor U13192 (N_13192,N_5985,N_7912);
nor U13193 (N_13193,N_7057,N_9295);
or U13194 (N_13194,N_8262,N_7730);
or U13195 (N_13195,N_8468,N_5604);
nand U13196 (N_13196,N_5517,N_8564);
or U13197 (N_13197,N_5624,N_9656);
and U13198 (N_13198,N_5991,N_9095);
nor U13199 (N_13199,N_7026,N_8226);
nand U13200 (N_13200,N_8809,N_9907);
nor U13201 (N_13201,N_5706,N_5027);
nor U13202 (N_13202,N_5232,N_7549);
or U13203 (N_13203,N_6056,N_6742);
and U13204 (N_13204,N_9879,N_7502);
nor U13205 (N_13205,N_6795,N_6954);
nor U13206 (N_13206,N_7365,N_6425);
nor U13207 (N_13207,N_8706,N_8995);
xor U13208 (N_13208,N_9547,N_5971);
xor U13209 (N_13209,N_6224,N_5344);
nor U13210 (N_13210,N_7338,N_7536);
nor U13211 (N_13211,N_8983,N_5392);
nand U13212 (N_13212,N_7945,N_5364);
nand U13213 (N_13213,N_9427,N_8015);
nand U13214 (N_13214,N_7720,N_8577);
nor U13215 (N_13215,N_5923,N_7475);
xor U13216 (N_13216,N_8771,N_6202);
nand U13217 (N_13217,N_5981,N_9919);
nor U13218 (N_13218,N_7177,N_7935);
or U13219 (N_13219,N_5437,N_9855);
xor U13220 (N_13220,N_5911,N_6724);
or U13221 (N_13221,N_6155,N_5292);
nor U13222 (N_13222,N_9651,N_8877);
nor U13223 (N_13223,N_8155,N_6346);
and U13224 (N_13224,N_7736,N_6681);
nor U13225 (N_13225,N_8029,N_5291);
or U13226 (N_13226,N_6465,N_5790);
and U13227 (N_13227,N_6309,N_9091);
nor U13228 (N_13228,N_8657,N_8069);
xnor U13229 (N_13229,N_6322,N_8807);
or U13230 (N_13230,N_5122,N_8448);
or U13231 (N_13231,N_7021,N_5647);
or U13232 (N_13232,N_5259,N_6987);
and U13233 (N_13233,N_6592,N_6033);
and U13234 (N_13234,N_8114,N_8527);
xor U13235 (N_13235,N_7865,N_8617);
nor U13236 (N_13236,N_7355,N_6065);
nor U13237 (N_13237,N_9600,N_8493);
nand U13238 (N_13238,N_7642,N_9659);
and U13239 (N_13239,N_8422,N_5881);
nand U13240 (N_13240,N_8435,N_9449);
xor U13241 (N_13241,N_5466,N_7057);
nor U13242 (N_13242,N_5926,N_5183);
nor U13243 (N_13243,N_7841,N_7027);
nor U13244 (N_13244,N_8980,N_5372);
nor U13245 (N_13245,N_7547,N_5414);
nand U13246 (N_13246,N_5252,N_6618);
and U13247 (N_13247,N_7057,N_7432);
or U13248 (N_13248,N_6780,N_7820);
nor U13249 (N_13249,N_7035,N_7538);
nor U13250 (N_13250,N_7632,N_8342);
nand U13251 (N_13251,N_5096,N_7285);
nor U13252 (N_13252,N_6382,N_8649);
or U13253 (N_13253,N_8549,N_8383);
nand U13254 (N_13254,N_5996,N_5916);
and U13255 (N_13255,N_7848,N_8708);
and U13256 (N_13256,N_8615,N_7856);
or U13257 (N_13257,N_6120,N_5323);
nor U13258 (N_13258,N_8716,N_8074);
nand U13259 (N_13259,N_5878,N_6413);
nand U13260 (N_13260,N_5762,N_9556);
and U13261 (N_13261,N_8797,N_7419);
and U13262 (N_13262,N_6880,N_8406);
nor U13263 (N_13263,N_6770,N_6602);
and U13264 (N_13264,N_9655,N_8077);
nand U13265 (N_13265,N_5853,N_7401);
and U13266 (N_13266,N_8223,N_7179);
or U13267 (N_13267,N_5365,N_7469);
nand U13268 (N_13268,N_8852,N_5499);
nor U13269 (N_13269,N_5573,N_9936);
and U13270 (N_13270,N_9507,N_6723);
and U13271 (N_13271,N_5234,N_8494);
nor U13272 (N_13272,N_8751,N_7616);
or U13273 (N_13273,N_5918,N_7345);
or U13274 (N_13274,N_8279,N_5552);
nand U13275 (N_13275,N_7726,N_9030);
nand U13276 (N_13276,N_7043,N_5300);
nand U13277 (N_13277,N_7511,N_8740);
or U13278 (N_13278,N_8496,N_7540);
and U13279 (N_13279,N_7145,N_8968);
nand U13280 (N_13280,N_5679,N_9956);
or U13281 (N_13281,N_5272,N_6978);
nand U13282 (N_13282,N_6122,N_7529);
or U13283 (N_13283,N_6817,N_6699);
and U13284 (N_13284,N_9418,N_9828);
and U13285 (N_13285,N_7790,N_7058);
or U13286 (N_13286,N_9239,N_7844);
nand U13287 (N_13287,N_7930,N_7704);
nand U13288 (N_13288,N_8509,N_6954);
nand U13289 (N_13289,N_7902,N_8316);
or U13290 (N_13290,N_7802,N_6982);
and U13291 (N_13291,N_6830,N_5514);
nor U13292 (N_13292,N_5884,N_7061);
nand U13293 (N_13293,N_6525,N_7099);
and U13294 (N_13294,N_7551,N_6896);
and U13295 (N_13295,N_9229,N_8135);
or U13296 (N_13296,N_9144,N_6901);
nand U13297 (N_13297,N_8144,N_5181);
nor U13298 (N_13298,N_9786,N_8413);
nand U13299 (N_13299,N_8787,N_7471);
and U13300 (N_13300,N_6167,N_9048);
and U13301 (N_13301,N_8166,N_9126);
and U13302 (N_13302,N_5420,N_7342);
nand U13303 (N_13303,N_8690,N_9454);
nor U13304 (N_13304,N_7462,N_9508);
nor U13305 (N_13305,N_6222,N_8192);
nor U13306 (N_13306,N_7189,N_8177);
or U13307 (N_13307,N_6920,N_9823);
and U13308 (N_13308,N_8931,N_8332);
nand U13309 (N_13309,N_5798,N_9094);
nand U13310 (N_13310,N_5326,N_7792);
or U13311 (N_13311,N_8621,N_8959);
nor U13312 (N_13312,N_8387,N_5113);
and U13313 (N_13313,N_6979,N_6760);
and U13314 (N_13314,N_6564,N_9757);
nor U13315 (N_13315,N_8906,N_5633);
nor U13316 (N_13316,N_5002,N_5788);
nand U13317 (N_13317,N_6409,N_7186);
xor U13318 (N_13318,N_6460,N_7405);
or U13319 (N_13319,N_5255,N_6583);
nand U13320 (N_13320,N_6077,N_7234);
nand U13321 (N_13321,N_5875,N_6655);
or U13322 (N_13322,N_5634,N_6009);
and U13323 (N_13323,N_5211,N_6181);
and U13324 (N_13324,N_8402,N_8199);
nand U13325 (N_13325,N_6885,N_9052);
nand U13326 (N_13326,N_6945,N_9785);
nand U13327 (N_13327,N_6929,N_7908);
nor U13328 (N_13328,N_6227,N_6122);
or U13329 (N_13329,N_7862,N_6407);
nor U13330 (N_13330,N_9754,N_6719);
nor U13331 (N_13331,N_6041,N_7083);
nor U13332 (N_13332,N_5937,N_8599);
nand U13333 (N_13333,N_5124,N_8227);
and U13334 (N_13334,N_7908,N_7510);
nor U13335 (N_13335,N_9663,N_9656);
and U13336 (N_13336,N_9188,N_6551);
and U13337 (N_13337,N_9651,N_9564);
or U13338 (N_13338,N_5550,N_6450);
nor U13339 (N_13339,N_6664,N_5199);
nor U13340 (N_13340,N_9227,N_6929);
xnor U13341 (N_13341,N_9697,N_9874);
or U13342 (N_13342,N_9422,N_9331);
nor U13343 (N_13343,N_9063,N_6143);
and U13344 (N_13344,N_7551,N_6073);
or U13345 (N_13345,N_8410,N_8718);
nand U13346 (N_13346,N_9629,N_5331);
xnor U13347 (N_13347,N_8480,N_6686);
nand U13348 (N_13348,N_8119,N_9272);
nor U13349 (N_13349,N_7328,N_5534);
and U13350 (N_13350,N_9551,N_6573);
and U13351 (N_13351,N_8834,N_6915);
and U13352 (N_13352,N_5156,N_8233);
nand U13353 (N_13353,N_8770,N_8921);
and U13354 (N_13354,N_6942,N_8597);
nor U13355 (N_13355,N_8853,N_5144);
and U13356 (N_13356,N_7508,N_5470);
and U13357 (N_13357,N_6307,N_7454);
or U13358 (N_13358,N_7982,N_8070);
xor U13359 (N_13359,N_5555,N_9920);
nor U13360 (N_13360,N_6086,N_9961);
nand U13361 (N_13361,N_9191,N_5271);
nand U13362 (N_13362,N_5541,N_7632);
nor U13363 (N_13363,N_7430,N_9476);
or U13364 (N_13364,N_6426,N_5559);
nand U13365 (N_13365,N_5597,N_6726);
and U13366 (N_13366,N_7380,N_5716);
nand U13367 (N_13367,N_5056,N_9446);
xnor U13368 (N_13368,N_5945,N_8245);
or U13369 (N_13369,N_6207,N_5909);
and U13370 (N_13370,N_6858,N_5819);
or U13371 (N_13371,N_9913,N_9764);
nand U13372 (N_13372,N_6108,N_5605);
or U13373 (N_13373,N_6775,N_7339);
nand U13374 (N_13374,N_7947,N_5173);
or U13375 (N_13375,N_9566,N_6540);
or U13376 (N_13376,N_7744,N_5225);
or U13377 (N_13377,N_7570,N_5864);
or U13378 (N_13378,N_8726,N_6381);
and U13379 (N_13379,N_9706,N_5674);
nand U13380 (N_13380,N_7666,N_8858);
and U13381 (N_13381,N_6146,N_7562);
nor U13382 (N_13382,N_5908,N_5311);
or U13383 (N_13383,N_6112,N_8000);
or U13384 (N_13384,N_6507,N_6914);
nand U13385 (N_13385,N_7854,N_9199);
xnor U13386 (N_13386,N_9728,N_8667);
nand U13387 (N_13387,N_9588,N_7501);
nand U13388 (N_13388,N_5241,N_6486);
nand U13389 (N_13389,N_5045,N_8765);
nor U13390 (N_13390,N_5997,N_5035);
nand U13391 (N_13391,N_7330,N_9117);
nand U13392 (N_13392,N_7590,N_9314);
and U13393 (N_13393,N_8108,N_9672);
and U13394 (N_13394,N_6013,N_8611);
xor U13395 (N_13395,N_7468,N_7940);
xor U13396 (N_13396,N_7067,N_6268);
xor U13397 (N_13397,N_7889,N_8088);
and U13398 (N_13398,N_6476,N_7903);
or U13399 (N_13399,N_8313,N_7467);
or U13400 (N_13400,N_9151,N_9776);
nand U13401 (N_13401,N_5022,N_5980);
or U13402 (N_13402,N_9944,N_9878);
xnor U13403 (N_13403,N_6443,N_7186);
nand U13404 (N_13404,N_9143,N_5261);
nand U13405 (N_13405,N_5202,N_5397);
nand U13406 (N_13406,N_9405,N_9498);
xnor U13407 (N_13407,N_6651,N_9265);
nor U13408 (N_13408,N_8210,N_8084);
nor U13409 (N_13409,N_5845,N_5551);
or U13410 (N_13410,N_9203,N_6622);
or U13411 (N_13411,N_8656,N_9465);
and U13412 (N_13412,N_6282,N_8416);
or U13413 (N_13413,N_9120,N_6472);
or U13414 (N_13414,N_5572,N_8799);
nand U13415 (N_13415,N_9690,N_7397);
nand U13416 (N_13416,N_5897,N_7972);
and U13417 (N_13417,N_5575,N_7463);
nand U13418 (N_13418,N_5396,N_6420);
nor U13419 (N_13419,N_6268,N_8254);
and U13420 (N_13420,N_9344,N_9826);
or U13421 (N_13421,N_9617,N_5318);
xor U13422 (N_13422,N_6348,N_8785);
nand U13423 (N_13423,N_9098,N_8773);
or U13424 (N_13424,N_5157,N_9841);
xor U13425 (N_13425,N_8496,N_7312);
nand U13426 (N_13426,N_9342,N_9542);
or U13427 (N_13427,N_7053,N_6196);
xor U13428 (N_13428,N_9135,N_6670);
nand U13429 (N_13429,N_9377,N_6074);
and U13430 (N_13430,N_9848,N_5214);
and U13431 (N_13431,N_5163,N_8368);
nand U13432 (N_13432,N_8374,N_5818);
and U13433 (N_13433,N_7602,N_9431);
xor U13434 (N_13434,N_8456,N_9063);
nand U13435 (N_13435,N_8987,N_9634);
or U13436 (N_13436,N_6933,N_5198);
nand U13437 (N_13437,N_8919,N_6623);
or U13438 (N_13438,N_6434,N_9823);
nor U13439 (N_13439,N_5302,N_9506);
or U13440 (N_13440,N_7222,N_6169);
xor U13441 (N_13441,N_5112,N_7131);
and U13442 (N_13442,N_7063,N_7501);
and U13443 (N_13443,N_9212,N_5399);
nand U13444 (N_13444,N_6178,N_7840);
or U13445 (N_13445,N_7061,N_8113);
nand U13446 (N_13446,N_9565,N_8411);
nand U13447 (N_13447,N_7772,N_5591);
or U13448 (N_13448,N_9955,N_9228);
nor U13449 (N_13449,N_8877,N_5320);
and U13450 (N_13450,N_7019,N_9317);
or U13451 (N_13451,N_6322,N_9465);
or U13452 (N_13452,N_5321,N_8893);
and U13453 (N_13453,N_5576,N_9340);
and U13454 (N_13454,N_9652,N_5260);
or U13455 (N_13455,N_9734,N_6246);
nand U13456 (N_13456,N_9358,N_7697);
nand U13457 (N_13457,N_9147,N_5379);
nor U13458 (N_13458,N_7224,N_6949);
or U13459 (N_13459,N_5544,N_7765);
nand U13460 (N_13460,N_9135,N_8487);
xor U13461 (N_13461,N_7009,N_9697);
and U13462 (N_13462,N_8663,N_6137);
xor U13463 (N_13463,N_8626,N_6215);
xor U13464 (N_13464,N_9049,N_6807);
or U13465 (N_13465,N_9312,N_8217);
nor U13466 (N_13466,N_9963,N_6223);
nor U13467 (N_13467,N_6443,N_5899);
nor U13468 (N_13468,N_8581,N_6197);
or U13469 (N_13469,N_7807,N_9715);
nor U13470 (N_13470,N_7126,N_5443);
xnor U13471 (N_13471,N_8723,N_6245);
and U13472 (N_13472,N_5046,N_5753);
or U13473 (N_13473,N_8044,N_8820);
nand U13474 (N_13474,N_5602,N_6637);
and U13475 (N_13475,N_7919,N_5769);
nor U13476 (N_13476,N_5208,N_5706);
nor U13477 (N_13477,N_7216,N_5125);
nor U13478 (N_13478,N_9412,N_5040);
or U13479 (N_13479,N_7734,N_8168);
nor U13480 (N_13480,N_6393,N_7476);
nor U13481 (N_13481,N_7521,N_7497);
xnor U13482 (N_13482,N_9678,N_7997);
nand U13483 (N_13483,N_6231,N_5355);
and U13484 (N_13484,N_5082,N_8759);
or U13485 (N_13485,N_5742,N_7593);
nor U13486 (N_13486,N_5462,N_8341);
nand U13487 (N_13487,N_6645,N_8264);
xor U13488 (N_13488,N_7972,N_7520);
or U13489 (N_13489,N_6778,N_9747);
nor U13490 (N_13490,N_9672,N_5188);
and U13491 (N_13491,N_6414,N_5280);
nand U13492 (N_13492,N_8389,N_5837);
xor U13493 (N_13493,N_5020,N_6950);
nand U13494 (N_13494,N_7839,N_8337);
nor U13495 (N_13495,N_6632,N_5562);
nor U13496 (N_13496,N_9185,N_5108);
xor U13497 (N_13497,N_8056,N_7187);
and U13498 (N_13498,N_8955,N_8913);
nand U13499 (N_13499,N_7845,N_8766);
nand U13500 (N_13500,N_9155,N_5348);
nor U13501 (N_13501,N_7609,N_8204);
nor U13502 (N_13502,N_8528,N_6744);
or U13503 (N_13503,N_7543,N_7241);
and U13504 (N_13504,N_6064,N_9279);
nand U13505 (N_13505,N_8869,N_7379);
and U13506 (N_13506,N_6810,N_5575);
and U13507 (N_13507,N_5575,N_5437);
or U13508 (N_13508,N_6481,N_7747);
or U13509 (N_13509,N_9831,N_5178);
nand U13510 (N_13510,N_6396,N_8055);
or U13511 (N_13511,N_9875,N_7623);
and U13512 (N_13512,N_9723,N_7760);
nand U13513 (N_13513,N_8899,N_6321);
nor U13514 (N_13514,N_9528,N_8258);
nand U13515 (N_13515,N_7894,N_7862);
and U13516 (N_13516,N_9571,N_7641);
nand U13517 (N_13517,N_8970,N_5616);
nand U13518 (N_13518,N_5217,N_8026);
or U13519 (N_13519,N_9127,N_8137);
nand U13520 (N_13520,N_5989,N_7679);
or U13521 (N_13521,N_5363,N_6776);
nand U13522 (N_13522,N_7592,N_7340);
xor U13523 (N_13523,N_6753,N_9179);
nor U13524 (N_13524,N_9026,N_9563);
nor U13525 (N_13525,N_9055,N_6880);
nor U13526 (N_13526,N_5622,N_6518);
nor U13527 (N_13527,N_8966,N_6516);
nand U13528 (N_13528,N_7245,N_5665);
or U13529 (N_13529,N_8182,N_9351);
and U13530 (N_13530,N_8493,N_8501);
or U13531 (N_13531,N_8065,N_5750);
nor U13532 (N_13532,N_9076,N_8419);
nand U13533 (N_13533,N_6631,N_8569);
and U13534 (N_13534,N_8604,N_8719);
or U13535 (N_13535,N_9236,N_6742);
and U13536 (N_13536,N_9526,N_7444);
and U13537 (N_13537,N_5208,N_8658);
or U13538 (N_13538,N_5710,N_6956);
nor U13539 (N_13539,N_6075,N_9166);
or U13540 (N_13540,N_9972,N_6067);
and U13541 (N_13541,N_9520,N_8357);
and U13542 (N_13542,N_7191,N_6354);
and U13543 (N_13543,N_9860,N_7773);
or U13544 (N_13544,N_6817,N_9159);
xnor U13545 (N_13545,N_6426,N_6192);
nand U13546 (N_13546,N_8722,N_8209);
and U13547 (N_13547,N_9382,N_8181);
nor U13548 (N_13548,N_6786,N_9473);
nor U13549 (N_13549,N_5609,N_7020);
nand U13550 (N_13550,N_7209,N_9946);
or U13551 (N_13551,N_8442,N_7198);
and U13552 (N_13552,N_9240,N_6178);
nor U13553 (N_13553,N_9023,N_6441);
nor U13554 (N_13554,N_5826,N_7845);
and U13555 (N_13555,N_8020,N_9420);
and U13556 (N_13556,N_5281,N_7741);
xor U13557 (N_13557,N_5494,N_5064);
nand U13558 (N_13558,N_5992,N_8169);
and U13559 (N_13559,N_7167,N_5258);
or U13560 (N_13560,N_8074,N_5414);
nand U13561 (N_13561,N_6920,N_7182);
or U13562 (N_13562,N_9138,N_7622);
nor U13563 (N_13563,N_9731,N_5789);
and U13564 (N_13564,N_9352,N_7837);
and U13565 (N_13565,N_8143,N_5907);
and U13566 (N_13566,N_9688,N_9290);
and U13567 (N_13567,N_8834,N_6868);
nand U13568 (N_13568,N_6574,N_6240);
or U13569 (N_13569,N_5431,N_8705);
nand U13570 (N_13570,N_5742,N_9173);
and U13571 (N_13571,N_7240,N_5372);
and U13572 (N_13572,N_9336,N_7399);
nor U13573 (N_13573,N_8851,N_8417);
and U13574 (N_13574,N_9425,N_9843);
and U13575 (N_13575,N_8831,N_8553);
nand U13576 (N_13576,N_8673,N_6245);
or U13577 (N_13577,N_5817,N_9476);
nand U13578 (N_13578,N_8102,N_9489);
nand U13579 (N_13579,N_5963,N_9725);
and U13580 (N_13580,N_5132,N_5327);
and U13581 (N_13581,N_7224,N_9223);
nor U13582 (N_13582,N_9600,N_7518);
nor U13583 (N_13583,N_7305,N_9131);
xor U13584 (N_13584,N_5139,N_8693);
and U13585 (N_13585,N_5817,N_9929);
nand U13586 (N_13586,N_5436,N_8522);
or U13587 (N_13587,N_5640,N_8456);
nand U13588 (N_13588,N_5966,N_7781);
and U13589 (N_13589,N_7810,N_6214);
nand U13590 (N_13590,N_9994,N_7631);
nor U13591 (N_13591,N_9099,N_7924);
nand U13592 (N_13592,N_9260,N_5077);
nand U13593 (N_13593,N_5799,N_7288);
or U13594 (N_13594,N_9060,N_7643);
and U13595 (N_13595,N_7421,N_6730);
nor U13596 (N_13596,N_8096,N_9811);
or U13597 (N_13597,N_7620,N_8827);
or U13598 (N_13598,N_5636,N_8009);
xnor U13599 (N_13599,N_8518,N_7430);
or U13600 (N_13600,N_6133,N_6111);
xnor U13601 (N_13601,N_9509,N_9979);
or U13602 (N_13602,N_6789,N_9571);
and U13603 (N_13603,N_8403,N_6056);
nand U13604 (N_13604,N_6469,N_6094);
nor U13605 (N_13605,N_5605,N_7978);
nor U13606 (N_13606,N_7141,N_9303);
nand U13607 (N_13607,N_7720,N_7034);
and U13608 (N_13608,N_8218,N_6892);
nand U13609 (N_13609,N_9377,N_7169);
and U13610 (N_13610,N_6509,N_5223);
or U13611 (N_13611,N_9716,N_7856);
xor U13612 (N_13612,N_6557,N_9982);
nor U13613 (N_13613,N_5099,N_7072);
or U13614 (N_13614,N_9010,N_7022);
or U13615 (N_13615,N_5098,N_5269);
and U13616 (N_13616,N_5350,N_7367);
nand U13617 (N_13617,N_5474,N_8750);
or U13618 (N_13618,N_5603,N_5401);
and U13619 (N_13619,N_5942,N_5129);
or U13620 (N_13620,N_5936,N_6526);
nor U13621 (N_13621,N_5280,N_9131);
nand U13622 (N_13622,N_5156,N_5885);
or U13623 (N_13623,N_5344,N_9417);
nor U13624 (N_13624,N_5752,N_7388);
nor U13625 (N_13625,N_6399,N_6085);
or U13626 (N_13626,N_8025,N_7012);
nor U13627 (N_13627,N_8847,N_6845);
or U13628 (N_13628,N_9588,N_9590);
nand U13629 (N_13629,N_6712,N_8432);
or U13630 (N_13630,N_7886,N_7393);
nor U13631 (N_13631,N_9874,N_7907);
xor U13632 (N_13632,N_5340,N_9785);
xor U13633 (N_13633,N_8986,N_7400);
and U13634 (N_13634,N_8070,N_7353);
nand U13635 (N_13635,N_9495,N_7170);
xnor U13636 (N_13636,N_9690,N_6936);
and U13637 (N_13637,N_8721,N_8884);
or U13638 (N_13638,N_5347,N_5577);
xor U13639 (N_13639,N_8820,N_9653);
nand U13640 (N_13640,N_7543,N_5868);
nand U13641 (N_13641,N_5003,N_9739);
nand U13642 (N_13642,N_8449,N_7406);
nand U13643 (N_13643,N_7897,N_8970);
nor U13644 (N_13644,N_5450,N_5294);
or U13645 (N_13645,N_5440,N_8447);
and U13646 (N_13646,N_6714,N_6635);
nand U13647 (N_13647,N_6584,N_7381);
nand U13648 (N_13648,N_7497,N_9323);
and U13649 (N_13649,N_5690,N_8101);
or U13650 (N_13650,N_5810,N_9631);
or U13651 (N_13651,N_8813,N_9164);
or U13652 (N_13652,N_6120,N_8178);
or U13653 (N_13653,N_6948,N_7661);
nor U13654 (N_13654,N_9785,N_5419);
and U13655 (N_13655,N_5972,N_7222);
xor U13656 (N_13656,N_6631,N_6778);
nand U13657 (N_13657,N_9920,N_8584);
or U13658 (N_13658,N_8532,N_5684);
xor U13659 (N_13659,N_6923,N_7867);
and U13660 (N_13660,N_6627,N_8433);
or U13661 (N_13661,N_6272,N_7304);
and U13662 (N_13662,N_6382,N_5306);
and U13663 (N_13663,N_5672,N_7920);
or U13664 (N_13664,N_5285,N_7875);
nor U13665 (N_13665,N_6234,N_6245);
nand U13666 (N_13666,N_9285,N_6475);
or U13667 (N_13667,N_8040,N_6361);
and U13668 (N_13668,N_9699,N_9711);
and U13669 (N_13669,N_9643,N_8847);
nand U13670 (N_13670,N_6546,N_7444);
and U13671 (N_13671,N_9489,N_5170);
or U13672 (N_13672,N_5196,N_8487);
nor U13673 (N_13673,N_9079,N_9787);
nor U13674 (N_13674,N_8131,N_6291);
or U13675 (N_13675,N_8012,N_7347);
nand U13676 (N_13676,N_6789,N_9307);
nand U13677 (N_13677,N_5030,N_9806);
xnor U13678 (N_13678,N_6848,N_9093);
or U13679 (N_13679,N_6070,N_7095);
and U13680 (N_13680,N_5996,N_5887);
or U13681 (N_13681,N_9082,N_6075);
and U13682 (N_13682,N_5192,N_9751);
or U13683 (N_13683,N_9733,N_9753);
or U13684 (N_13684,N_9397,N_5685);
nor U13685 (N_13685,N_8545,N_8057);
and U13686 (N_13686,N_5615,N_8359);
or U13687 (N_13687,N_7806,N_5433);
or U13688 (N_13688,N_8239,N_7896);
or U13689 (N_13689,N_5065,N_9927);
or U13690 (N_13690,N_8013,N_9105);
nor U13691 (N_13691,N_6929,N_9882);
nor U13692 (N_13692,N_6160,N_7367);
nor U13693 (N_13693,N_8514,N_9459);
nor U13694 (N_13694,N_5689,N_9084);
nand U13695 (N_13695,N_5094,N_8079);
and U13696 (N_13696,N_8440,N_9445);
and U13697 (N_13697,N_8752,N_5481);
or U13698 (N_13698,N_5653,N_9708);
nor U13699 (N_13699,N_9489,N_8192);
and U13700 (N_13700,N_9740,N_6678);
and U13701 (N_13701,N_9368,N_7812);
nand U13702 (N_13702,N_8766,N_9858);
xnor U13703 (N_13703,N_6301,N_5817);
and U13704 (N_13704,N_8923,N_7890);
or U13705 (N_13705,N_5829,N_8534);
or U13706 (N_13706,N_6389,N_9217);
and U13707 (N_13707,N_5567,N_8041);
xnor U13708 (N_13708,N_9968,N_8442);
nor U13709 (N_13709,N_7802,N_5003);
and U13710 (N_13710,N_9738,N_5359);
or U13711 (N_13711,N_8426,N_6937);
xnor U13712 (N_13712,N_6632,N_9121);
nand U13713 (N_13713,N_5221,N_9061);
nand U13714 (N_13714,N_8995,N_8681);
nor U13715 (N_13715,N_6259,N_9066);
or U13716 (N_13716,N_8061,N_5724);
or U13717 (N_13717,N_5102,N_8123);
and U13718 (N_13718,N_6321,N_9531);
and U13719 (N_13719,N_9983,N_9707);
and U13720 (N_13720,N_5778,N_8666);
nor U13721 (N_13721,N_6499,N_6387);
or U13722 (N_13722,N_7101,N_7433);
and U13723 (N_13723,N_8668,N_9873);
xor U13724 (N_13724,N_5733,N_6211);
and U13725 (N_13725,N_9293,N_6525);
or U13726 (N_13726,N_8730,N_7426);
or U13727 (N_13727,N_9878,N_8086);
and U13728 (N_13728,N_9237,N_7787);
nor U13729 (N_13729,N_5141,N_8442);
nand U13730 (N_13730,N_6605,N_8106);
nand U13731 (N_13731,N_9975,N_6645);
nor U13732 (N_13732,N_6392,N_6828);
and U13733 (N_13733,N_7531,N_7597);
and U13734 (N_13734,N_8866,N_9065);
nor U13735 (N_13735,N_5199,N_6429);
or U13736 (N_13736,N_6526,N_8127);
nor U13737 (N_13737,N_6602,N_5546);
or U13738 (N_13738,N_6791,N_5026);
or U13739 (N_13739,N_9485,N_8298);
nor U13740 (N_13740,N_9604,N_5025);
xor U13741 (N_13741,N_8597,N_5493);
nor U13742 (N_13742,N_7912,N_9060);
or U13743 (N_13743,N_8470,N_5837);
nor U13744 (N_13744,N_6444,N_9813);
or U13745 (N_13745,N_5268,N_9192);
and U13746 (N_13746,N_9274,N_7541);
or U13747 (N_13747,N_6830,N_8751);
or U13748 (N_13748,N_8578,N_5885);
and U13749 (N_13749,N_6786,N_9318);
and U13750 (N_13750,N_5661,N_7049);
xor U13751 (N_13751,N_6591,N_7991);
nand U13752 (N_13752,N_5048,N_6722);
nand U13753 (N_13753,N_7525,N_9042);
xor U13754 (N_13754,N_8884,N_7848);
or U13755 (N_13755,N_6610,N_9996);
and U13756 (N_13756,N_8387,N_8817);
and U13757 (N_13757,N_6606,N_8336);
xnor U13758 (N_13758,N_6426,N_7665);
xnor U13759 (N_13759,N_9897,N_7621);
and U13760 (N_13760,N_7604,N_8006);
nand U13761 (N_13761,N_9154,N_5404);
or U13762 (N_13762,N_7652,N_9582);
nand U13763 (N_13763,N_6670,N_7237);
and U13764 (N_13764,N_8611,N_5057);
or U13765 (N_13765,N_9469,N_9979);
nor U13766 (N_13766,N_5550,N_6745);
xnor U13767 (N_13767,N_5061,N_9773);
nor U13768 (N_13768,N_9398,N_8945);
xnor U13769 (N_13769,N_6276,N_5695);
or U13770 (N_13770,N_8320,N_7939);
or U13771 (N_13771,N_9072,N_5486);
nor U13772 (N_13772,N_6485,N_6869);
and U13773 (N_13773,N_7043,N_9537);
nand U13774 (N_13774,N_7288,N_8648);
xor U13775 (N_13775,N_8255,N_9572);
and U13776 (N_13776,N_7641,N_7932);
or U13777 (N_13777,N_9289,N_7672);
nand U13778 (N_13778,N_9030,N_6542);
and U13779 (N_13779,N_5624,N_7204);
xnor U13780 (N_13780,N_5812,N_6034);
and U13781 (N_13781,N_8383,N_9742);
or U13782 (N_13782,N_8553,N_5845);
and U13783 (N_13783,N_7787,N_8734);
nand U13784 (N_13784,N_5587,N_6248);
or U13785 (N_13785,N_9692,N_9174);
and U13786 (N_13786,N_8971,N_9400);
and U13787 (N_13787,N_9119,N_9263);
nand U13788 (N_13788,N_6484,N_6864);
and U13789 (N_13789,N_8330,N_9006);
or U13790 (N_13790,N_8519,N_8404);
or U13791 (N_13791,N_5345,N_8640);
xnor U13792 (N_13792,N_5833,N_9381);
nor U13793 (N_13793,N_6692,N_5026);
and U13794 (N_13794,N_6086,N_5397);
or U13795 (N_13795,N_6631,N_6939);
or U13796 (N_13796,N_5521,N_9569);
and U13797 (N_13797,N_9538,N_7096);
nor U13798 (N_13798,N_6904,N_5124);
xnor U13799 (N_13799,N_5051,N_6266);
and U13800 (N_13800,N_6869,N_7711);
or U13801 (N_13801,N_8796,N_7779);
or U13802 (N_13802,N_6272,N_5564);
or U13803 (N_13803,N_9631,N_7453);
nor U13804 (N_13804,N_6130,N_9349);
nor U13805 (N_13805,N_5164,N_5121);
xnor U13806 (N_13806,N_6381,N_7565);
and U13807 (N_13807,N_7265,N_6204);
and U13808 (N_13808,N_5094,N_8340);
nand U13809 (N_13809,N_7829,N_5337);
nor U13810 (N_13810,N_6223,N_6939);
or U13811 (N_13811,N_5113,N_6297);
nor U13812 (N_13812,N_5222,N_6903);
and U13813 (N_13813,N_5984,N_6556);
and U13814 (N_13814,N_8757,N_7343);
nand U13815 (N_13815,N_7236,N_8787);
or U13816 (N_13816,N_7937,N_6159);
nor U13817 (N_13817,N_8879,N_7202);
or U13818 (N_13818,N_7065,N_9134);
nor U13819 (N_13819,N_5300,N_6035);
or U13820 (N_13820,N_9779,N_7219);
xnor U13821 (N_13821,N_7404,N_5266);
or U13822 (N_13822,N_9672,N_7779);
and U13823 (N_13823,N_9642,N_8363);
xnor U13824 (N_13824,N_5205,N_7118);
nand U13825 (N_13825,N_8255,N_8885);
or U13826 (N_13826,N_9469,N_5142);
and U13827 (N_13827,N_8425,N_7715);
nor U13828 (N_13828,N_5927,N_7843);
or U13829 (N_13829,N_8289,N_8487);
or U13830 (N_13830,N_9314,N_5301);
or U13831 (N_13831,N_7212,N_9253);
or U13832 (N_13832,N_5036,N_5244);
xnor U13833 (N_13833,N_9790,N_9559);
nor U13834 (N_13834,N_5319,N_5404);
nand U13835 (N_13835,N_7675,N_7714);
and U13836 (N_13836,N_8115,N_5790);
nand U13837 (N_13837,N_8981,N_7087);
nor U13838 (N_13838,N_8151,N_5812);
and U13839 (N_13839,N_7433,N_7183);
nor U13840 (N_13840,N_5850,N_9416);
nor U13841 (N_13841,N_6391,N_9641);
nor U13842 (N_13842,N_5254,N_5723);
or U13843 (N_13843,N_9929,N_7372);
nor U13844 (N_13844,N_7322,N_8960);
and U13845 (N_13845,N_5681,N_5743);
and U13846 (N_13846,N_5600,N_8352);
or U13847 (N_13847,N_9140,N_6154);
nand U13848 (N_13848,N_9743,N_6432);
xnor U13849 (N_13849,N_7026,N_6291);
and U13850 (N_13850,N_5872,N_8932);
and U13851 (N_13851,N_6597,N_9759);
or U13852 (N_13852,N_5960,N_5939);
nor U13853 (N_13853,N_5325,N_6381);
nand U13854 (N_13854,N_9879,N_6386);
nor U13855 (N_13855,N_9420,N_6840);
and U13856 (N_13856,N_6645,N_5534);
nor U13857 (N_13857,N_5183,N_5828);
nand U13858 (N_13858,N_5120,N_7530);
nand U13859 (N_13859,N_9632,N_7224);
nor U13860 (N_13860,N_5335,N_6534);
nor U13861 (N_13861,N_9675,N_7489);
nand U13862 (N_13862,N_5801,N_8251);
nor U13863 (N_13863,N_9608,N_6286);
nor U13864 (N_13864,N_9550,N_9098);
and U13865 (N_13865,N_7758,N_5782);
nor U13866 (N_13866,N_5063,N_7950);
xor U13867 (N_13867,N_5678,N_8419);
xor U13868 (N_13868,N_5919,N_8990);
and U13869 (N_13869,N_9095,N_7892);
nand U13870 (N_13870,N_9979,N_7828);
xor U13871 (N_13871,N_5240,N_9980);
nand U13872 (N_13872,N_5245,N_9375);
nand U13873 (N_13873,N_8417,N_8606);
and U13874 (N_13874,N_8411,N_6338);
nor U13875 (N_13875,N_8739,N_8078);
nor U13876 (N_13876,N_9836,N_5478);
nor U13877 (N_13877,N_7180,N_6600);
or U13878 (N_13878,N_9681,N_9973);
and U13879 (N_13879,N_8899,N_6674);
nand U13880 (N_13880,N_6597,N_7430);
or U13881 (N_13881,N_5857,N_6168);
nand U13882 (N_13882,N_5502,N_7833);
and U13883 (N_13883,N_6630,N_9916);
or U13884 (N_13884,N_9910,N_7377);
and U13885 (N_13885,N_8717,N_6481);
nand U13886 (N_13886,N_5373,N_6831);
or U13887 (N_13887,N_9248,N_5610);
nand U13888 (N_13888,N_8836,N_9129);
nand U13889 (N_13889,N_5348,N_9398);
and U13890 (N_13890,N_6536,N_8033);
nor U13891 (N_13891,N_8737,N_5619);
nand U13892 (N_13892,N_9514,N_7614);
nor U13893 (N_13893,N_5076,N_8374);
nand U13894 (N_13894,N_6581,N_5303);
nor U13895 (N_13895,N_7219,N_7000);
xnor U13896 (N_13896,N_9013,N_6012);
or U13897 (N_13897,N_5157,N_7465);
and U13898 (N_13898,N_6808,N_8093);
nand U13899 (N_13899,N_7133,N_6879);
nand U13900 (N_13900,N_8729,N_7019);
nand U13901 (N_13901,N_8089,N_6520);
and U13902 (N_13902,N_9914,N_9494);
and U13903 (N_13903,N_7639,N_9393);
and U13904 (N_13904,N_8216,N_6792);
or U13905 (N_13905,N_7844,N_5233);
nand U13906 (N_13906,N_8886,N_6981);
and U13907 (N_13907,N_8745,N_9507);
nor U13908 (N_13908,N_9662,N_6072);
and U13909 (N_13909,N_9719,N_9661);
xnor U13910 (N_13910,N_7763,N_6588);
nor U13911 (N_13911,N_8367,N_8936);
nor U13912 (N_13912,N_9848,N_9721);
or U13913 (N_13913,N_5649,N_7259);
and U13914 (N_13914,N_8933,N_9190);
nand U13915 (N_13915,N_5792,N_6314);
and U13916 (N_13916,N_7200,N_6949);
nor U13917 (N_13917,N_7564,N_7055);
and U13918 (N_13918,N_5106,N_5366);
nor U13919 (N_13919,N_6404,N_6452);
or U13920 (N_13920,N_8584,N_7640);
nor U13921 (N_13921,N_9711,N_6557);
nand U13922 (N_13922,N_6431,N_6393);
and U13923 (N_13923,N_6058,N_6228);
nand U13924 (N_13924,N_7318,N_7016);
or U13925 (N_13925,N_6328,N_5247);
nor U13926 (N_13926,N_6314,N_7770);
xor U13927 (N_13927,N_7687,N_6153);
xnor U13928 (N_13928,N_5304,N_8616);
and U13929 (N_13929,N_9022,N_8237);
or U13930 (N_13930,N_6249,N_9116);
or U13931 (N_13931,N_7198,N_8854);
nand U13932 (N_13932,N_9471,N_6586);
nand U13933 (N_13933,N_9192,N_6986);
nor U13934 (N_13934,N_6582,N_6810);
and U13935 (N_13935,N_7682,N_9257);
or U13936 (N_13936,N_6454,N_6511);
nor U13937 (N_13937,N_6209,N_8477);
or U13938 (N_13938,N_5040,N_6366);
nor U13939 (N_13939,N_5224,N_6992);
xor U13940 (N_13940,N_7340,N_7588);
and U13941 (N_13941,N_5936,N_6917);
and U13942 (N_13942,N_6290,N_7756);
and U13943 (N_13943,N_6631,N_5448);
xnor U13944 (N_13944,N_6126,N_5989);
and U13945 (N_13945,N_8624,N_8084);
nor U13946 (N_13946,N_6750,N_5128);
and U13947 (N_13947,N_5430,N_5075);
nand U13948 (N_13948,N_8055,N_6162);
nand U13949 (N_13949,N_8734,N_6453);
xor U13950 (N_13950,N_9107,N_6892);
and U13951 (N_13951,N_6364,N_6792);
nor U13952 (N_13952,N_5936,N_6444);
nor U13953 (N_13953,N_8705,N_7407);
nor U13954 (N_13954,N_7335,N_9321);
or U13955 (N_13955,N_7524,N_6431);
nand U13956 (N_13956,N_5788,N_6968);
xor U13957 (N_13957,N_6240,N_7192);
and U13958 (N_13958,N_9573,N_7491);
and U13959 (N_13959,N_7006,N_8379);
and U13960 (N_13960,N_5444,N_6689);
or U13961 (N_13961,N_8395,N_7838);
nand U13962 (N_13962,N_7227,N_8264);
nand U13963 (N_13963,N_6035,N_5652);
and U13964 (N_13964,N_9698,N_5938);
or U13965 (N_13965,N_7100,N_7756);
nand U13966 (N_13966,N_6160,N_7359);
and U13967 (N_13967,N_7293,N_6636);
or U13968 (N_13968,N_5394,N_7128);
xnor U13969 (N_13969,N_9310,N_5177);
and U13970 (N_13970,N_7661,N_8762);
nor U13971 (N_13971,N_8724,N_6951);
nor U13972 (N_13972,N_9480,N_9544);
nand U13973 (N_13973,N_6484,N_8254);
nand U13974 (N_13974,N_7890,N_8898);
and U13975 (N_13975,N_8176,N_7683);
or U13976 (N_13976,N_7744,N_5725);
nand U13977 (N_13977,N_9335,N_5652);
nor U13978 (N_13978,N_6443,N_8992);
nand U13979 (N_13979,N_7142,N_7657);
nand U13980 (N_13980,N_9716,N_7964);
nor U13981 (N_13981,N_8787,N_7203);
and U13982 (N_13982,N_6083,N_6993);
and U13983 (N_13983,N_6194,N_7133);
nor U13984 (N_13984,N_9525,N_8134);
xnor U13985 (N_13985,N_6069,N_9129);
nor U13986 (N_13986,N_6594,N_7278);
nor U13987 (N_13987,N_6208,N_9537);
and U13988 (N_13988,N_8560,N_6459);
nand U13989 (N_13989,N_6710,N_8322);
and U13990 (N_13990,N_6308,N_8929);
nor U13991 (N_13991,N_9909,N_5396);
and U13992 (N_13992,N_7563,N_5187);
or U13993 (N_13993,N_5771,N_9237);
nor U13994 (N_13994,N_8086,N_9550);
nand U13995 (N_13995,N_7697,N_6882);
or U13996 (N_13996,N_9796,N_5457);
xor U13997 (N_13997,N_9947,N_5779);
and U13998 (N_13998,N_7191,N_9950);
or U13999 (N_13999,N_5976,N_5226);
or U14000 (N_14000,N_9888,N_9799);
nor U14001 (N_14001,N_5007,N_8949);
and U14002 (N_14002,N_5963,N_6306);
or U14003 (N_14003,N_7923,N_5319);
and U14004 (N_14004,N_9132,N_6312);
nand U14005 (N_14005,N_8317,N_9745);
and U14006 (N_14006,N_5859,N_6079);
or U14007 (N_14007,N_6777,N_9766);
nor U14008 (N_14008,N_6324,N_7317);
or U14009 (N_14009,N_8209,N_8690);
xnor U14010 (N_14010,N_8205,N_9705);
nor U14011 (N_14011,N_8665,N_5372);
nand U14012 (N_14012,N_8856,N_7974);
and U14013 (N_14013,N_5456,N_9918);
or U14014 (N_14014,N_5286,N_7135);
and U14015 (N_14015,N_9599,N_7825);
and U14016 (N_14016,N_7196,N_5115);
nand U14017 (N_14017,N_7336,N_6067);
xor U14018 (N_14018,N_5840,N_6852);
nand U14019 (N_14019,N_7416,N_8543);
nor U14020 (N_14020,N_5628,N_8943);
and U14021 (N_14021,N_7179,N_7027);
nor U14022 (N_14022,N_7207,N_5436);
nand U14023 (N_14023,N_9855,N_9850);
nor U14024 (N_14024,N_9003,N_6942);
and U14025 (N_14025,N_9634,N_6012);
nor U14026 (N_14026,N_5461,N_8393);
nor U14027 (N_14027,N_9567,N_5715);
nand U14028 (N_14028,N_6427,N_8643);
nor U14029 (N_14029,N_6837,N_5084);
and U14030 (N_14030,N_5657,N_8718);
or U14031 (N_14031,N_5224,N_8707);
nand U14032 (N_14032,N_9468,N_5014);
nand U14033 (N_14033,N_9448,N_7961);
nand U14034 (N_14034,N_7955,N_5683);
nand U14035 (N_14035,N_7040,N_9056);
and U14036 (N_14036,N_9516,N_7234);
nand U14037 (N_14037,N_6462,N_9940);
or U14038 (N_14038,N_6257,N_7363);
or U14039 (N_14039,N_6337,N_7996);
nor U14040 (N_14040,N_5383,N_8440);
nor U14041 (N_14041,N_8436,N_9190);
and U14042 (N_14042,N_8067,N_6073);
xnor U14043 (N_14043,N_6045,N_9509);
nand U14044 (N_14044,N_8292,N_8384);
nand U14045 (N_14045,N_8067,N_7556);
and U14046 (N_14046,N_7618,N_9400);
nand U14047 (N_14047,N_7121,N_6690);
nand U14048 (N_14048,N_7161,N_7808);
nand U14049 (N_14049,N_8724,N_6418);
nor U14050 (N_14050,N_7927,N_6528);
or U14051 (N_14051,N_8106,N_7886);
nor U14052 (N_14052,N_5141,N_9801);
and U14053 (N_14053,N_5912,N_9343);
nor U14054 (N_14054,N_8183,N_7028);
or U14055 (N_14055,N_6539,N_9656);
nor U14056 (N_14056,N_7613,N_9400);
or U14057 (N_14057,N_7680,N_7854);
or U14058 (N_14058,N_9417,N_7837);
or U14059 (N_14059,N_8551,N_5128);
nor U14060 (N_14060,N_6707,N_7791);
and U14061 (N_14061,N_7554,N_6819);
nor U14062 (N_14062,N_7619,N_9247);
xnor U14063 (N_14063,N_7531,N_6943);
and U14064 (N_14064,N_9763,N_5648);
and U14065 (N_14065,N_7569,N_5111);
and U14066 (N_14066,N_9690,N_9373);
xnor U14067 (N_14067,N_6366,N_8971);
nand U14068 (N_14068,N_7524,N_9915);
xnor U14069 (N_14069,N_9394,N_6490);
and U14070 (N_14070,N_6212,N_7573);
nand U14071 (N_14071,N_7019,N_7618);
and U14072 (N_14072,N_9235,N_6534);
nor U14073 (N_14073,N_6585,N_9672);
nand U14074 (N_14074,N_8919,N_8088);
and U14075 (N_14075,N_7323,N_5076);
or U14076 (N_14076,N_5246,N_7643);
or U14077 (N_14077,N_8313,N_6349);
nor U14078 (N_14078,N_5201,N_7017);
xor U14079 (N_14079,N_5246,N_7155);
or U14080 (N_14080,N_7996,N_6415);
nand U14081 (N_14081,N_5608,N_9032);
and U14082 (N_14082,N_6084,N_7714);
xnor U14083 (N_14083,N_8157,N_8463);
and U14084 (N_14084,N_7255,N_6784);
nor U14085 (N_14085,N_7429,N_8583);
and U14086 (N_14086,N_5635,N_9511);
and U14087 (N_14087,N_7152,N_7977);
xor U14088 (N_14088,N_5672,N_8837);
nor U14089 (N_14089,N_8051,N_6436);
nor U14090 (N_14090,N_6762,N_9352);
or U14091 (N_14091,N_7972,N_5960);
and U14092 (N_14092,N_7610,N_9798);
nor U14093 (N_14093,N_7539,N_6104);
and U14094 (N_14094,N_5948,N_7050);
and U14095 (N_14095,N_5107,N_5561);
and U14096 (N_14096,N_7661,N_9686);
or U14097 (N_14097,N_9628,N_8982);
nor U14098 (N_14098,N_9101,N_9676);
and U14099 (N_14099,N_7215,N_8848);
or U14100 (N_14100,N_5820,N_5804);
or U14101 (N_14101,N_5626,N_7165);
nand U14102 (N_14102,N_7120,N_7072);
and U14103 (N_14103,N_8802,N_9819);
and U14104 (N_14104,N_7182,N_5622);
xnor U14105 (N_14105,N_7030,N_7869);
nand U14106 (N_14106,N_6082,N_6249);
and U14107 (N_14107,N_8731,N_9031);
and U14108 (N_14108,N_6790,N_8347);
nand U14109 (N_14109,N_8717,N_5251);
nand U14110 (N_14110,N_5103,N_6139);
nand U14111 (N_14111,N_9369,N_8008);
and U14112 (N_14112,N_7989,N_5007);
and U14113 (N_14113,N_8336,N_9166);
nand U14114 (N_14114,N_8421,N_6125);
xnor U14115 (N_14115,N_8030,N_5757);
and U14116 (N_14116,N_6244,N_7308);
nand U14117 (N_14117,N_8523,N_8421);
nand U14118 (N_14118,N_9039,N_5757);
or U14119 (N_14119,N_5834,N_9040);
nor U14120 (N_14120,N_9701,N_8642);
and U14121 (N_14121,N_7760,N_7142);
and U14122 (N_14122,N_8298,N_7075);
xnor U14123 (N_14123,N_6751,N_7947);
nand U14124 (N_14124,N_6622,N_5538);
or U14125 (N_14125,N_5891,N_9105);
or U14126 (N_14126,N_6111,N_6955);
nor U14127 (N_14127,N_5160,N_9046);
and U14128 (N_14128,N_9984,N_6772);
nor U14129 (N_14129,N_6220,N_6311);
and U14130 (N_14130,N_8514,N_7581);
nand U14131 (N_14131,N_5188,N_7622);
nand U14132 (N_14132,N_5227,N_5197);
and U14133 (N_14133,N_7665,N_8769);
nand U14134 (N_14134,N_5131,N_9394);
and U14135 (N_14135,N_9655,N_6200);
xnor U14136 (N_14136,N_6857,N_5385);
nor U14137 (N_14137,N_7309,N_7103);
or U14138 (N_14138,N_9878,N_5570);
or U14139 (N_14139,N_7503,N_7228);
nor U14140 (N_14140,N_8176,N_9113);
and U14141 (N_14141,N_8464,N_8404);
nor U14142 (N_14142,N_6942,N_8606);
nand U14143 (N_14143,N_5836,N_6674);
nand U14144 (N_14144,N_7004,N_5654);
nor U14145 (N_14145,N_8422,N_9475);
nor U14146 (N_14146,N_5871,N_7613);
nor U14147 (N_14147,N_8813,N_6649);
xor U14148 (N_14148,N_8658,N_9524);
nand U14149 (N_14149,N_5562,N_8187);
and U14150 (N_14150,N_9743,N_5262);
or U14151 (N_14151,N_9599,N_5373);
nand U14152 (N_14152,N_6503,N_6418);
nand U14153 (N_14153,N_6666,N_9453);
nor U14154 (N_14154,N_6430,N_7548);
xor U14155 (N_14155,N_6305,N_7866);
or U14156 (N_14156,N_9093,N_9966);
xor U14157 (N_14157,N_8376,N_5917);
and U14158 (N_14158,N_5644,N_7108);
nand U14159 (N_14159,N_9924,N_5046);
and U14160 (N_14160,N_6280,N_9207);
and U14161 (N_14161,N_8637,N_5403);
or U14162 (N_14162,N_9293,N_6550);
nor U14163 (N_14163,N_7083,N_9335);
or U14164 (N_14164,N_8756,N_6026);
or U14165 (N_14165,N_7278,N_9001);
xnor U14166 (N_14166,N_5648,N_6192);
nor U14167 (N_14167,N_8248,N_6469);
nand U14168 (N_14168,N_9388,N_8227);
nand U14169 (N_14169,N_6805,N_6690);
nor U14170 (N_14170,N_7517,N_9926);
or U14171 (N_14171,N_5978,N_5173);
xor U14172 (N_14172,N_7188,N_9281);
and U14173 (N_14173,N_9620,N_9854);
or U14174 (N_14174,N_7285,N_8219);
nor U14175 (N_14175,N_5687,N_7095);
and U14176 (N_14176,N_7561,N_8362);
and U14177 (N_14177,N_5271,N_8727);
nor U14178 (N_14178,N_8826,N_7207);
nand U14179 (N_14179,N_5821,N_9725);
nor U14180 (N_14180,N_9367,N_8476);
xnor U14181 (N_14181,N_5519,N_9911);
nor U14182 (N_14182,N_5804,N_7520);
or U14183 (N_14183,N_7078,N_9790);
or U14184 (N_14184,N_7754,N_7730);
nor U14185 (N_14185,N_5253,N_5198);
nand U14186 (N_14186,N_8394,N_5970);
nand U14187 (N_14187,N_7813,N_9318);
nand U14188 (N_14188,N_5873,N_7433);
and U14189 (N_14189,N_8067,N_7262);
nor U14190 (N_14190,N_7145,N_8352);
and U14191 (N_14191,N_6770,N_8000);
nor U14192 (N_14192,N_5766,N_9427);
nand U14193 (N_14193,N_8544,N_5539);
nor U14194 (N_14194,N_6249,N_9648);
nor U14195 (N_14195,N_5840,N_5186);
and U14196 (N_14196,N_6773,N_7363);
nor U14197 (N_14197,N_5574,N_9314);
nand U14198 (N_14198,N_7406,N_5768);
or U14199 (N_14199,N_9193,N_9674);
and U14200 (N_14200,N_8887,N_9409);
nor U14201 (N_14201,N_5090,N_8371);
or U14202 (N_14202,N_9936,N_6144);
and U14203 (N_14203,N_5288,N_6622);
or U14204 (N_14204,N_5605,N_8315);
nand U14205 (N_14205,N_8468,N_9446);
nand U14206 (N_14206,N_9368,N_9625);
nor U14207 (N_14207,N_5869,N_8856);
or U14208 (N_14208,N_6440,N_6439);
nor U14209 (N_14209,N_9537,N_9013);
and U14210 (N_14210,N_8951,N_9859);
and U14211 (N_14211,N_9594,N_5115);
xnor U14212 (N_14212,N_7814,N_6715);
nor U14213 (N_14213,N_8170,N_9910);
and U14214 (N_14214,N_6223,N_9076);
or U14215 (N_14215,N_9952,N_6212);
nor U14216 (N_14216,N_8066,N_5137);
nor U14217 (N_14217,N_8448,N_7360);
and U14218 (N_14218,N_9075,N_5461);
and U14219 (N_14219,N_5098,N_7192);
nand U14220 (N_14220,N_8404,N_8249);
xor U14221 (N_14221,N_7649,N_9631);
and U14222 (N_14222,N_6493,N_8928);
nand U14223 (N_14223,N_6742,N_5826);
nor U14224 (N_14224,N_8997,N_5439);
and U14225 (N_14225,N_7014,N_5582);
nor U14226 (N_14226,N_6052,N_8655);
nand U14227 (N_14227,N_9411,N_5424);
xor U14228 (N_14228,N_7896,N_6237);
nand U14229 (N_14229,N_6108,N_8821);
and U14230 (N_14230,N_8079,N_5947);
nand U14231 (N_14231,N_5228,N_5976);
or U14232 (N_14232,N_7815,N_6823);
or U14233 (N_14233,N_6585,N_8628);
or U14234 (N_14234,N_5456,N_5064);
or U14235 (N_14235,N_9729,N_8768);
and U14236 (N_14236,N_9279,N_6485);
nand U14237 (N_14237,N_6796,N_6385);
nand U14238 (N_14238,N_7152,N_9246);
nand U14239 (N_14239,N_8884,N_9981);
nor U14240 (N_14240,N_9363,N_7719);
nor U14241 (N_14241,N_8867,N_6488);
and U14242 (N_14242,N_5673,N_9079);
xnor U14243 (N_14243,N_7588,N_9086);
or U14244 (N_14244,N_9770,N_9809);
nor U14245 (N_14245,N_8495,N_8008);
or U14246 (N_14246,N_9176,N_8513);
nand U14247 (N_14247,N_7976,N_8249);
or U14248 (N_14248,N_9270,N_5179);
nor U14249 (N_14249,N_8726,N_5639);
nor U14250 (N_14250,N_8769,N_7608);
nand U14251 (N_14251,N_8034,N_8968);
xnor U14252 (N_14252,N_5246,N_5315);
or U14253 (N_14253,N_9148,N_5584);
or U14254 (N_14254,N_6770,N_6414);
nor U14255 (N_14255,N_7657,N_7231);
or U14256 (N_14256,N_7975,N_6717);
or U14257 (N_14257,N_9623,N_8832);
nand U14258 (N_14258,N_9150,N_5490);
xnor U14259 (N_14259,N_7935,N_7854);
nand U14260 (N_14260,N_5031,N_6417);
and U14261 (N_14261,N_9738,N_6486);
nor U14262 (N_14262,N_5018,N_9452);
nor U14263 (N_14263,N_5872,N_6728);
or U14264 (N_14264,N_6375,N_5715);
nor U14265 (N_14265,N_7226,N_8886);
or U14266 (N_14266,N_8364,N_9428);
and U14267 (N_14267,N_6479,N_8228);
and U14268 (N_14268,N_6922,N_6352);
or U14269 (N_14269,N_9014,N_6725);
nor U14270 (N_14270,N_9025,N_6912);
or U14271 (N_14271,N_9558,N_6727);
xor U14272 (N_14272,N_7011,N_8344);
xor U14273 (N_14273,N_6594,N_5633);
xor U14274 (N_14274,N_5522,N_9435);
or U14275 (N_14275,N_5507,N_6419);
nor U14276 (N_14276,N_7251,N_7076);
nand U14277 (N_14277,N_5194,N_8582);
nor U14278 (N_14278,N_7702,N_6918);
or U14279 (N_14279,N_7062,N_9988);
nor U14280 (N_14280,N_8120,N_7087);
nor U14281 (N_14281,N_9085,N_9138);
xor U14282 (N_14282,N_9770,N_9131);
nor U14283 (N_14283,N_8770,N_5433);
or U14284 (N_14284,N_8936,N_5155);
or U14285 (N_14285,N_8497,N_5073);
and U14286 (N_14286,N_6097,N_8204);
or U14287 (N_14287,N_8446,N_9477);
nor U14288 (N_14288,N_7010,N_7720);
xor U14289 (N_14289,N_9079,N_7413);
nand U14290 (N_14290,N_9764,N_6299);
nor U14291 (N_14291,N_7524,N_8583);
or U14292 (N_14292,N_6723,N_6193);
xnor U14293 (N_14293,N_5524,N_9338);
and U14294 (N_14294,N_7357,N_6526);
or U14295 (N_14295,N_9793,N_8307);
or U14296 (N_14296,N_7550,N_6737);
xnor U14297 (N_14297,N_7110,N_6266);
nand U14298 (N_14298,N_9631,N_6184);
nor U14299 (N_14299,N_9795,N_8119);
nor U14300 (N_14300,N_7537,N_5236);
and U14301 (N_14301,N_8731,N_8496);
and U14302 (N_14302,N_9122,N_9869);
nor U14303 (N_14303,N_9730,N_9140);
and U14304 (N_14304,N_6800,N_5165);
xor U14305 (N_14305,N_8763,N_7620);
or U14306 (N_14306,N_9448,N_8704);
nand U14307 (N_14307,N_8447,N_6102);
nor U14308 (N_14308,N_8653,N_7699);
and U14309 (N_14309,N_7704,N_7123);
or U14310 (N_14310,N_6321,N_8656);
or U14311 (N_14311,N_8591,N_6639);
nand U14312 (N_14312,N_8937,N_8023);
xnor U14313 (N_14313,N_7213,N_9353);
and U14314 (N_14314,N_8792,N_9658);
and U14315 (N_14315,N_9044,N_5652);
or U14316 (N_14316,N_5385,N_8071);
or U14317 (N_14317,N_7625,N_5947);
nand U14318 (N_14318,N_7847,N_8906);
and U14319 (N_14319,N_9383,N_9578);
nand U14320 (N_14320,N_5984,N_5992);
nand U14321 (N_14321,N_7670,N_7287);
and U14322 (N_14322,N_9942,N_8370);
or U14323 (N_14323,N_8442,N_6037);
and U14324 (N_14324,N_8817,N_7748);
and U14325 (N_14325,N_8788,N_7779);
nor U14326 (N_14326,N_8701,N_7000);
nand U14327 (N_14327,N_8012,N_7526);
nand U14328 (N_14328,N_9722,N_9376);
xnor U14329 (N_14329,N_8015,N_8798);
or U14330 (N_14330,N_6609,N_9976);
and U14331 (N_14331,N_7906,N_9676);
or U14332 (N_14332,N_6730,N_8396);
nor U14333 (N_14333,N_7883,N_8974);
xor U14334 (N_14334,N_5330,N_7463);
and U14335 (N_14335,N_7268,N_6993);
or U14336 (N_14336,N_8494,N_7243);
and U14337 (N_14337,N_5538,N_8526);
or U14338 (N_14338,N_5771,N_5815);
nand U14339 (N_14339,N_6119,N_8171);
nand U14340 (N_14340,N_7763,N_8719);
nand U14341 (N_14341,N_5664,N_9088);
and U14342 (N_14342,N_5522,N_5786);
or U14343 (N_14343,N_5518,N_9395);
nor U14344 (N_14344,N_6762,N_6102);
or U14345 (N_14345,N_8827,N_8932);
nand U14346 (N_14346,N_9261,N_7525);
and U14347 (N_14347,N_7880,N_6702);
and U14348 (N_14348,N_8315,N_6882);
nor U14349 (N_14349,N_8084,N_5792);
and U14350 (N_14350,N_7489,N_5497);
nand U14351 (N_14351,N_9978,N_9906);
or U14352 (N_14352,N_9887,N_6075);
or U14353 (N_14353,N_5195,N_6548);
nand U14354 (N_14354,N_6642,N_9064);
xor U14355 (N_14355,N_7284,N_5250);
or U14356 (N_14356,N_8536,N_8855);
nor U14357 (N_14357,N_8304,N_5994);
nor U14358 (N_14358,N_6415,N_6210);
and U14359 (N_14359,N_8182,N_5548);
nand U14360 (N_14360,N_6618,N_5804);
nor U14361 (N_14361,N_6654,N_5369);
nand U14362 (N_14362,N_7880,N_5188);
nand U14363 (N_14363,N_6379,N_5013);
and U14364 (N_14364,N_5167,N_5636);
or U14365 (N_14365,N_6701,N_5414);
xnor U14366 (N_14366,N_8224,N_9526);
xor U14367 (N_14367,N_7230,N_8812);
or U14368 (N_14368,N_7269,N_7465);
xor U14369 (N_14369,N_7174,N_5380);
nor U14370 (N_14370,N_7177,N_6373);
nor U14371 (N_14371,N_7453,N_9709);
and U14372 (N_14372,N_6672,N_6589);
and U14373 (N_14373,N_5427,N_5230);
and U14374 (N_14374,N_6517,N_9351);
nand U14375 (N_14375,N_6945,N_7796);
nor U14376 (N_14376,N_9157,N_5370);
and U14377 (N_14377,N_8634,N_5148);
and U14378 (N_14378,N_5466,N_9252);
and U14379 (N_14379,N_9129,N_8151);
or U14380 (N_14380,N_6057,N_8296);
and U14381 (N_14381,N_6139,N_6487);
nand U14382 (N_14382,N_5967,N_9599);
xor U14383 (N_14383,N_7765,N_7408);
and U14384 (N_14384,N_7964,N_5925);
and U14385 (N_14385,N_8325,N_8647);
and U14386 (N_14386,N_7799,N_9627);
or U14387 (N_14387,N_7185,N_7313);
and U14388 (N_14388,N_5892,N_5725);
nand U14389 (N_14389,N_5296,N_5609);
nand U14390 (N_14390,N_5273,N_5982);
nor U14391 (N_14391,N_5842,N_6542);
and U14392 (N_14392,N_8868,N_8065);
nor U14393 (N_14393,N_9782,N_7156);
and U14394 (N_14394,N_6533,N_7543);
nor U14395 (N_14395,N_7818,N_9214);
and U14396 (N_14396,N_5856,N_6718);
xor U14397 (N_14397,N_6440,N_7288);
nand U14398 (N_14398,N_5543,N_8104);
nand U14399 (N_14399,N_9598,N_5843);
nor U14400 (N_14400,N_5869,N_5166);
nand U14401 (N_14401,N_5450,N_9075);
nand U14402 (N_14402,N_8251,N_5029);
or U14403 (N_14403,N_9273,N_5230);
and U14404 (N_14404,N_6860,N_9598);
nand U14405 (N_14405,N_9047,N_5748);
nand U14406 (N_14406,N_8466,N_6031);
or U14407 (N_14407,N_5159,N_8961);
nand U14408 (N_14408,N_7345,N_5890);
or U14409 (N_14409,N_8619,N_7257);
and U14410 (N_14410,N_8733,N_6543);
nand U14411 (N_14411,N_6044,N_7946);
and U14412 (N_14412,N_7932,N_5040);
nand U14413 (N_14413,N_9549,N_5441);
xor U14414 (N_14414,N_6331,N_8810);
xnor U14415 (N_14415,N_6773,N_6548);
or U14416 (N_14416,N_5528,N_8803);
nor U14417 (N_14417,N_7025,N_9153);
nor U14418 (N_14418,N_7381,N_7012);
or U14419 (N_14419,N_9468,N_8804);
and U14420 (N_14420,N_6599,N_8733);
or U14421 (N_14421,N_8967,N_6141);
nor U14422 (N_14422,N_7618,N_8011);
nor U14423 (N_14423,N_8794,N_6404);
nor U14424 (N_14424,N_5339,N_9323);
nand U14425 (N_14425,N_5446,N_8463);
nand U14426 (N_14426,N_8826,N_9104);
and U14427 (N_14427,N_5971,N_6078);
or U14428 (N_14428,N_9158,N_7822);
and U14429 (N_14429,N_9907,N_9799);
xor U14430 (N_14430,N_9612,N_8781);
nand U14431 (N_14431,N_6615,N_8817);
nand U14432 (N_14432,N_5236,N_7669);
or U14433 (N_14433,N_9640,N_5159);
nand U14434 (N_14434,N_5520,N_8097);
nor U14435 (N_14435,N_7339,N_7420);
or U14436 (N_14436,N_5463,N_5385);
xor U14437 (N_14437,N_6825,N_7376);
nor U14438 (N_14438,N_9858,N_7623);
nand U14439 (N_14439,N_6155,N_9786);
and U14440 (N_14440,N_6921,N_5609);
nand U14441 (N_14441,N_5511,N_6210);
nand U14442 (N_14442,N_8318,N_9332);
and U14443 (N_14443,N_5637,N_6202);
nor U14444 (N_14444,N_9791,N_8862);
or U14445 (N_14445,N_7274,N_6041);
nand U14446 (N_14446,N_5161,N_5511);
or U14447 (N_14447,N_8709,N_5677);
and U14448 (N_14448,N_9966,N_6756);
and U14449 (N_14449,N_6238,N_9188);
nand U14450 (N_14450,N_6950,N_8220);
xor U14451 (N_14451,N_9448,N_9956);
and U14452 (N_14452,N_6181,N_6966);
nor U14453 (N_14453,N_9355,N_6433);
or U14454 (N_14454,N_8860,N_6556);
nor U14455 (N_14455,N_5406,N_7201);
nand U14456 (N_14456,N_8974,N_9963);
nor U14457 (N_14457,N_9400,N_9865);
or U14458 (N_14458,N_5551,N_6364);
nand U14459 (N_14459,N_7184,N_5348);
xnor U14460 (N_14460,N_6731,N_6940);
nor U14461 (N_14461,N_7415,N_8728);
nor U14462 (N_14462,N_6188,N_6135);
nand U14463 (N_14463,N_7142,N_8917);
or U14464 (N_14464,N_9797,N_7878);
nor U14465 (N_14465,N_6388,N_9419);
and U14466 (N_14466,N_7248,N_5899);
xor U14467 (N_14467,N_6214,N_5471);
xor U14468 (N_14468,N_5688,N_8528);
or U14469 (N_14469,N_9222,N_5622);
nand U14470 (N_14470,N_8667,N_9214);
nor U14471 (N_14471,N_8763,N_9730);
nand U14472 (N_14472,N_5297,N_8855);
nor U14473 (N_14473,N_5563,N_9087);
or U14474 (N_14474,N_5905,N_8036);
nand U14475 (N_14475,N_5438,N_7298);
nand U14476 (N_14476,N_6631,N_6625);
nand U14477 (N_14477,N_8876,N_5115);
or U14478 (N_14478,N_8388,N_7485);
nand U14479 (N_14479,N_7376,N_9539);
nor U14480 (N_14480,N_7914,N_7961);
xnor U14481 (N_14481,N_8598,N_8454);
nor U14482 (N_14482,N_8153,N_7484);
or U14483 (N_14483,N_6861,N_5890);
nor U14484 (N_14484,N_8687,N_7285);
or U14485 (N_14485,N_6964,N_5559);
and U14486 (N_14486,N_5901,N_7318);
xor U14487 (N_14487,N_9744,N_8598);
xnor U14488 (N_14488,N_6673,N_5930);
or U14489 (N_14489,N_8032,N_6734);
or U14490 (N_14490,N_8624,N_9417);
nor U14491 (N_14491,N_5317,N_7219);
nand U14492 (N_14492,N_8476,N_5460);
nor U14493 (N_14493,N_7202,N_6195);
nor U14494 (N_14494,N_5166,N_7270);
and U14495 (N_14495,N_5313,N_6221);
nand U14496 (N_14496,N_9906,N_7019);
nand U14497 (N_14497,N_6687,N_5429);
or U14498 (N_14498,N_6373,N_8400);
and U14499 (N_14499,N_5759,N_9319);
nand U14500 (N_14500,N_8806,N_8507);
xnor U14501 (N_14501,N_5255,N_7813);
or U14502 (N_14502,N_9772,N_9944);
and U14503 (N_14503,N_7859,N_8808);
nand U14504 (N_14504,N_8759,N_6767);
or U14505 (N_14505,N_9908,N_9738);
nand U14506 (N_14506,N_9689,N_8919);
nand U14507 (N_14507,N_7818,N_5059);
and U14508 (N_14508,N_5324,N_9497);
nand U14509 (N_14509,N_9061,N_7746);
nand U14510 (N_14510,N_8368,N_5117);
nand U14511 (N_14511,N_8200,N_6491);
xor U14512 (N_14512,N_5261,N_8142);
and U14513 (N_14513,N_7037,N_9918);
nand U14514 (N_14514,N_8160,N_8548);
nor U14515 (N_14515,N_6813,N_6967);
and U14516 (N_14516,N_5843,N_6204);
nand U14517 (N_14517,N_6900,N_6873);
nand U14518 (N_14518,N_8258,N_6199);
and U14519 (N_14519,N_5699,N_8603);
nand U14520 (N_14520,N_8910,N_9664);
nor U14521 (N_14521,N_9296,N_6926);
and U14522 (N_14522,N_6821,N_6332);
and U14523 (N_14523,N_7287,N_6465);
nor U14524 (N_14524,N_5155,N_6459);
and U14525 (N_14525,N_8923,N_9961);
xor U14526 (N_14526,N_6629,N_8702);
and U14527 (N_14527,N_6706,N_9155);
nand U14528 (N_14528,N_6523,N_5421);
and U14529 (N_14529,N_9969,N_8200);
and U14530 (N_14530,N_7347,N_8555);
and U14531 (N_14531,N_9854,N_5848);
and U14532 (N_14532,N_7158,N_8762);
nor U14533 (N_14533,N_8052,N_6193);
or U14534 (N_14534,N_5336,N_8106);
or U14535 (N_14535,N_9000,N_6104);
or U14536 (N_14536,N_6791,N_9024);
nor U14537 (N_14537,N_9630,N_7715);
nor U14538 (N_14538,N_9071,N_8488);
or U14539 (N_14539,N_9764,N_5665);
and U14540 (N_14540,N_5318,N_5438);
and U14541 (N_14541,N_7647,N_5398);
nand U14542 (N_14542,N_9064,N_8602);
nand U14543 (N_14543,N_8805,N_8409);
and U14544 (N_14544,N_6497,N_8200);
nand U14545 (N_14545,N_7300,N_5149);
or U14546 (N_14546,N_9541,N_8367);
or U14547 (N_14547,N_8049,N_7138);
nand U14548 (N_14548,N_7450,N_7791);
nand U14549 (N_14549,N_7492,N_9136);
nand U14550 (N_14550,N_8192,N_6873);
or U14551 (N_14551,N_5768,N_9998);
and U14552 (N_14552,N_7446,N_9546);
xnor U14553 (N_14553,N_9556,N_5782);
nor U14554 (N_14554,N_5929,N_5981);
nor U14555 (N_14555,N_6476,N_8036);
or U14556 (N_14556,N_5129,N_6596);
nor U14557 (N_14557,N_5827,N_9205);
nor U14558 (N_14558,N_8400,N_8158);
nor U14559 (N_14559,N_7410,N_8504);
nor U14560 (N_14560,N_7023,N_8034);
nor U14561 (N_14561,N_6214,N_9152);
or U14562 (N_14562,N_7681,N_5080);
and U14563 (N_14563,N_9903,N_9907);
nand U14564 (N_14564,N_9407,N_6691);
nand U14565 (N_14565,N_9683,N_9946);
or U14566 (N_14566,N_6838,N_6521);
and U14567 (N_14567,N_9397,N_9734);
nor U14568 (N_14568,N_8663,N_5398);
nor U14569 (N_14569,N_9895,N_6006);
or U14570 (N_14570,N_8397,N_5298);
or U14571 (N_14571,N_6048,N_8968);
xnor U14572 (N_14572,N_9541,N_6061);
nor U14573 (N_14573,N_8783,N_7734);
nand U14574 (N_14574,N_8467,N_7215);
nor U14575 (N_14575,N_8958,N_6854);
nand U14576 (N_14576,N_9748,N_9469);
or U14577 (N_14577,N_5699,N_5413);
and U14578 (N_14578,N_9516,N_7209);
or U14579 (N_14579,N_8856,N_5878);
nand U14580 (N_14580,N_5968,N_8090);
or U14581 (N_14581,N_5219,N_9111);
xnor U14582 (N_14582,N_5276,N_7246);
nor U14583 (N_14583,N_6580,N_8094);
and U14584 (N_14584,N_8676,N_6146);
or U14585 (N_14585,N_8039,N_5411);
nor U14586 (N_14586,N_7538,N_8749);
or U14587 (N_14587,N_5020,N_9212);
or U14588 (N_14588,N_8805,N_8987);
and U14589 (N_14589,N_6887,N_9896);
and U14590 (N_14590,N_9099,N_9335);
xor U14591 (N_14591,N_8193,N_9652);
nand U14592 (N_14592,N_7193,N_5827);
and U14593 (N_14593,N_7716,N_6546);
nor U14594 (N_14594,N_6708,N_8488);
nor U14595 (N_14595,N_6817,N_9861);
and U14596 (N_14596,N_5240,N_6050);
or U14597 (N_14597,N_7588,N_8901);
nor U14598 (N_14598,N_9900,N_5086);
or U14599 (N_14599,N_8450,N_9247);
nor U14600 (N_14600,N_6312,N_5866);
and U14601 (N_14601,N_8199,N_7495);
nor U14602 (N_14602,N_9260,N_8957);
nor U14603 (N_14603,N_9983,N_6338);
or U14604 (N_14604,N_5962,N_5010);
nor U14605 (N_14605,N_7069,N_6867);
or U14606 (N_14606,N_8835,N_8893);
and U14607 (N_14607,N_6508,N_5865);
or U14608 (N_14608,N_5276,N_5778);
or U14609 (N_14609,N_7556,N_5159);
nand U14610 (N_14610,N_7914,N_5129);
nand U14611 (N_14611,N_8893,N_5539);
and U14612 (N_14612,N_6876,N_5517);
and U14613 (N_14613,N_7662,N_8949);
or U14614 (N_14614,N_5728,N_6906);
and U14615 (N_14615,N_7679,N_6601);
nor U14616 (N_14616,N_9147,N_5817);
or U14617 (N_14617,N_9918,N_6704);
nand U14618 (N_14618,N_7302,N_7592);
nor U14619 (N_14619,N_7712,N_9104);
nand U14620 (N_14620,N_7305,N_9311);
nor U14621 (N_14621,N_7580,N_9414);
xnor U14622 (N_14622,N_5428,N_6094);
or U14623 (N_14623,N_5466,N_5425);
and U14624 (N_14624,N_9570,N_8895);
xnor U14625 (N_14625,N_8297,N_6729);
and U14626 (N_14626,N_5021,N_9655);
nand U14627 (N_14627,N_8033,N_7614);
nor U14628 (N_14628,N_5202,N_9810);
nor U14629 (N_14629,N_7114,N_9607);
nand U14630 (N_14630,N_5841,N_8483);
nand U14631 (N_14631,N_5189,N_7888);
and U14632 (N_14632,N_6599,N_7153);
or U14633 (N_14633,N_5776,N_9648);
nor U14634 (N_14634,N_7929,N_9713);
and U14635 (N_14635,N_5935,N_9683);
or U14636 (N_14636,N_5653,N_7475);
nor U14637 (N_14637,N_6143,N_8440);
nand U14638 (N_14638,N_9398,N_5904);
and U14639 (N_14639,N_8776,N_8784);
nand U14640 (N_14640,N_7060,N_7917);
or U14641 (N_14641,N_7191,N_8052);
nor U14642 (N_14642,N_7710,N_7147);
or U14643 (N_14643,N_8462,N_8806);
xor U14644 (N_14644,N_8150,N_8650);
nand U14645 (N_14645,N_8288,N_8298);
and U14646 (N_14646,N_8286,N_5120);
and U14647 (N_14647,N_6799,N_8968);
or U14648 (N_14648,N_6609,N_7678);
and U14649 (N_14649,N_6389,N_9530);
and U14650 (N_14650,N_6934,N_8131);
or U14651 (N_14651,N_6544,N_5919);
nand U14652 (N_14652,N_5166,N_6806);
nor U14653 (N_14653,N_6709,N_5879);
nand U14654 (N_14654,N_5843,N_8802);
xor U14655 (N_14655,N_5041,N_8660);
and U14656 (N_14656,N_7219,N_8625);
or U14657 (N_14657,N_6691,N_9908);
nand U14658 (N_14658,N_9122,N_8159);
nand U14659 (N_14659,N_9986,N_5477);
nor U14660 (N_14660,N_9333,N_7048);
nand U14661 (N_14661,N_9252,N_5429);
nand U14662 (N_14662,N_9056,N_8858);
or U14663 (N_14663,N_9622,N_5211);
nand U14664 (N_14664,N_7066,N_9273);
or U14665 (N_14665,N_7340,N_9526);
or U14666 (N_14666,N_9053,N_6980);
nand U14667 (N_14667,N_6496,N_5266);
nor U14668 (N_14668,N_6789,N_5606);
or U14669 (N_14669,N_6175,N_6351);
and U14670 (N_14670,N_6071,N_9912);
and U14671 (N_14671,N_9571,N_6134);
or U14672 (N_14672,N_5769,N_8992);
and U14673 (N_14673,N_6247,N_6741);
nor U14674 (N_14674,N_5037,N_8416);
and U14675 (N_14675,N_9494,N_8306);
xnor U14676 (N_14676,N_6518,N_7976);
and U14677 (N_14677,N_7100,N_8263);
nand U14678 (N_14678,N_6583,N_7966);
nand U14679 (N_14679,N_7282,N_9479);
nor U14680 (N_14680,N_7110,N_9319);
nand U14681 (N_14681,N_8661,N_7270);
nor U14682 (N_14682,N_6624,N_9215);
and U14683 (N_14683,N_8340,N_8382);
nor U14684 (N_14684,N_5067,N_7129);
nor U14685 (N_14685,N_6239,N_7705);
or U14686 (N_14686,N_7154,N_5083);
nor U14687 (N_14687,N_8849,N_5703);
or U14688 (N_14688,N_5582,N_9865);
and U14689 (N_14689,N_5003,N_7097);
or U14690 (N_14690,N_5552,N_9281);
and U14691 (N_14691,N_6255,N_7036);
nor U14692 (N_14692,N_7207,N_9547);
and U14693 (N_14693,N_6880,N_6633);
nand U14694 (N_14694,N_8022,N_9236);
and U14695 (N_14695,N_9466,N_7958);
nor U14696 (N_14696,N_5697,N_8756);
or U14697 (N_14697,N_7906,N_5435);
or U14698 (N_14698,N_7348,N_7091);
or U14699 (N_14699,N_7534,N_6641);
and U14700 (N_14700,N_8911,N_8321);
nor U14701 (N_14701,N_6574,N_9061);
and U14702 (N_14702,N_8804,N_5506);
xnor U14703 (N_14703,N_5464,N_9859);
nor U14704 (N_14704,N_7336,N_6808);
or U14705 (N_14705,N_6574,N_5722);
nand U14706 (N_14706,N_7904,N_5221);
and U14707 (N_14707,N_9715,N_6862);
or U14708 (N_14708,N_8776,N_6942);
nor U14709 (N_14709,N_7675,N_7030);
xnor U14710 (N_14710,N_6529,N_8593);
xnor U14711 (N_14711,N_6031,N_9364);
xnor U14712 (N_14712,N_8184,N_9855);
and U14713 (N_14713,N_9726,N_6367);
nor U14714 (N_14714,N_9318,N_8275);
and U14715 (N_14715,N_9728,N_7974);
or U14716 (N_14716,N_7324,N_9526);
nor U14717 (N_14717,N_8834,N_7698);
nor U14718 (N_14718,N_7103,N_8816);
nor U14719 (N_14719,N_9480,N_9550);
nor U14720 (N_14720,N_9609,N_5276);
and U14721 (N_14721,N_7789,N_6053);
nor U14722 (N_14722,N_6625,N_9318);
or U14723 (N_14723,N_7496,N_9319);
xnor U14724 (N_14724,N_8446,N_6311);
and U14725 (N_14725,N_8622,N_9208);
xnor U14726 (N_14726,N_9640,N_9068);
and U14727 (N_14727,N_8218,N_9989);
nand U14728 (N_14728,N_8128,N_5939);
nand U14729 (N_14729,N_6029,N_9123);
nor U14730 (N_14730,N_9314,N_6684);
or U14731 (N_14731,N_6667,N_5545);
or U14732 (N_14732,N_6422,N_6558);
or U14733 (N_14733,N_6256,N_7142);
or U14734 (N_14734,N_6273,N_8351);
nand U14735 (N_14735,N_5579,N_5155);
xnor U14736 (N_14736,N_8168,N_8790);
or U14737 (N_14737,N_7540,N_8393);
or U14738 (N_14738,N_7579,N_9626);
or U14739 (N_14739,N_8170,N_6460);
nand U14740 (N_14740,N_5410,N_8900);
or U14741 (N_14741,N_9711,N_5904);
or U14742 (N_14742,N_7145,N_5385);
and U14743 (N_14743,N_9098,N_5497);
nand U14744 (N_14744,N_7071,N_9194);
and U14745 (N_14745,N_6650,N_7871);
nor U14746 (N_14746,N_7531,N_6799);
nor U14747 (N_14747,N_6709,N_6118);
nor U14748 (N_14748,N_7518,N_9472);
nand U14749 (N_14749,N_8769,N_7467);
nand U14750 (N_14750,N_6672,N_6529);
nand U14751 (N_14751,N_6649,N_5179);
xor U14752 (N_14752,N_5583,N_5291);
and U14753 (N_14753,N_9801,N_7382);
nand U14754 (N_14754,N_8584,N_8051);
nand U14755 (N_14755,N_8528,N_7264);
and U14756 (N_14756,N_9124,N_5530);
or U14757 (N_14757,N_9355,N_9001);
nand U14758 (N_14758,N_6054,N_5860);
xor U14759 (N_14759,N_9463,N_5420);
nand U14760 (N_14760,N_5119,N_7918);
and U14761 (N_14761,N_8617,N_7092);
nor U14762 (N_14762,N_6627,N_9534);
and U14763 (N_14763,N_6226,N_5528);
nand U14764 (N_14764,N_8320,N_7012);
nor U14765 (N_14765,N_6973,N_7351);
nand U14766 (N_14766,N_9056,N_9618);
and U14767 (N_14767,N_8942,N_8789);
and U14768 (N_14768,N_6508,N_8524);
or U14769 (N_14769,N_9930,N_6478);
and U14770 (N_14770,N_6073,N_5644);
nor U14771 (N_14771,N_6804,N_9260);
nor U14772 (N_14772,N_9213,N_7659);
and U14773 (N_14773,N_9784,N_8645);
nor U14774 (N_14774,N_5868,N_6411);
and U14775 (N_14775,N_9437,N_8365);
nor U14776 (N_14776,N_7327,N_7737);
or U14777 (N_14777,N_7594,N_6525);
nor U14778 (N_14778,N_5423,N_7598);
nand U14779 (N_14779,N_9466,N_6645);
nor U14780 (N_14780,N_6344,N_8835);
or U14781 (N_14781,N_6204,N_8453);
or U14782 (N_14782,N_7497,N_8074);
and U14783 (N_14783,N_5153,N_9330);
and U14784 (N_14784,N_6613,N_5980);
and U14785 (N_14785,N_5907,N_7606);
or U14786 (N_14786,N_6543,N_5655);
nand U14787 (N_14787,N_5265,N_8634);
nor U14788 (N_14788,N_8313,N_9127);
nor U14789 (N_14789,N_8136,N_8377);
and U14790 (N_14790,N_8802,N_7915);
nor U14791 (N_14791,N_9369,N_7960);
xor U14792 (N_14792,N_8690,N_6665);
nor U14793 (N_14793,N_6839,N_8731);
and U14794 (N_14794,N_5954,N_9549);
nand U14795 (N_14795,N_6960,N_7519);
or U14796 (N_14796,N_6364,N_8855);
and U14797 (N_14797,N_7828,N_7084);
xnor U14798 (N_14798,N_8272,N_6416);
nand U14799 (N_14799,N_8107,N_8733);
nand U14800 (N_14800,N_6886,N_7136);
nor U14801 (N_14801,N_9162,N_6036);
and U14802 (N_14802,N_6606,N_6055);
nand U14803 (N_14803,N_5313,N_8930);
nor U14804 (N_14804,N_7515,N_7158);
or U14805 (N_14805,N_8242,N_8630);
and U14806 (N_14806,N_7570,N_9704);
or U14807 (N_14807,N_8074,N_8333);
nand U14808 (N_14808,N_9448,N_6106);
or U14809 (N_14809,N_7703,N_8842);
or U14810 (N_14810,N_8837,N_8372);
nand U14811 (N_14811,N_9587,N_9629);
and U14812 (N_14812,N_5899,N_5515);
nand U14813 (N_14813,N_9277,N_5960);
or U14814 (N_14814,N_7099,N_7346);
and U14815 (N_14815,N_5028,N_8124);
nand U14816 (N_14816,N_9066,N_7021);
nand U14817 (N_14817,N_5106,N_8726);
nand U14818 (N_14818,N_9279,N_5877);
and U14819 (N_14819,N_5594,N_5468);
nand U14820 (N_14820,N_8084,N_9369);
nor U14821 (N_14821,N_8378,N_9085);
nor U14822 (N_14822,N_9784,N_7318);
or U14823 (N_14823,N_9046,N_6205);
xnor U14824 (N_14824,N_6168,N_5589);
nor U14825 (N_14825,N_8113,N_7813);
nand U14826 (N_14826,N_6318,N_6200);
nor U14827 (N_14827,N_7132,N_7351);
or U14828 (N_14828,N_6099,N_8760);
nor U14829 (N_14829,N_9726,N_8652);
and U14830 (N_14830,N_8503,N_5412);
or U14831 (N_14831,N_5477,N_8709);
and U14832 (N_14832,N_5031,N_8479);
and U14833 (N_14833,N_6999,N_7842);
nand U14834 (N_14834,N_9527,N_5697);
and U14835 (N_14835,N_5684,N_5699);
nor U14836 (N_14836,N_7963,N_7156);
and U14837 (N_14837,N_5877,N_8947);
nand U14838 (N_14838,N_8328,N_6125);
or U14839 (N_14839,N_8076,N_6089);
or U14840 (N_14840,N_6082,N_6613);
nand U14841 (N_14841,N_9733,N_9364);
or U14842 (N_14842,N_5814,N_8729);
nor U14843 (N_14843,N_6659,N_5609);
nor U14844 (N_14844,N_7911,N_5793);
nor U14845 (N_14845,N_7644,N_6159);
nand U14846 (N_14846,N_5855,N_6984);
nor U14847 (N_14847,N_9992,N_5835);
and U14848 (N_14848,N_5614,N_9195);
nand U14849 (N_14849,N_9076,N_5675);
nor U14850 (N_14850,N_8830,N_6437);
nor U14851 (N_14851,N_5004,N_7024);
or U14852 (N_14852,N_9771,N_8887);
and U14853 (N_14853,N_7434,N_7896);
nand U14854 (N_14854,N_5171,N_9476);
or U14855 (N_14855,N_6430,N_7542);
and U14856 (N_14856,N_9673,N_9839);
nor U14857 (N_14857,N_8228,N_7499);
and U14858 (N_14858,N_9674,N_6178);
nand U14859 (N_14859,N_5212,N_8913);
nor U14860 (N_14860,N_9083,N_9699);
nor U14861 (N_14861,N_9199,N_6743);
or U14862 (N_14862,N_9444,N_5375);
nor U14863 (N_14863,N_5158,N_5759);
nor U14864 (N_14864,N_5559,N_7023);
nor U14865 (N_14865,N_8122,N_9205);
and U14866 (N_14866,N_5184,N_9297);
or U14867 (N_14867,N_6418,N_6239);
nor U14868 (N_14868,N_7808,N_5714);
nor U14869 (N_14869,N_9259,N_8175);
nand U14870 (N_14870,N_8792,N_5212);
nor U14871 (N_14871,N_5428,N_6967);
and U14872 (N_14872,N_7072,N_7749);
or U14873 (N_14873,N_8514,N_8802);
and U14874 (N_14874,N_5625,N_6104);
nor U14875 (N_14875,N_7126,N_7236);
nand U14876 (N_14876,N_8474,N_8435);
nor U14877 (N_14877,N_9812,N_7096);
nor U14878 (N_14878,N_5243,N_8688);
nor U14879 (N_14879,N_8620,N_6063);
or U14880 (N_14880,N_7175,N_7778);
nor U14881 (N_14881,N_7483,N_6819);
and U14882 (N_14882,N_7135,N_8296);
and U14883 (N_14883,N_7047,N_7283);
or U14884 (N_14884,N_9597,N_5845);
and U14885 (N_14885,N_5621,N_8797);
nor U14886 (N_14886,N_6998,N_7870);
or U14887 (N_14887,N_8818,N_9386);
or U14888 (N_14888,N_8487,N_5068);
nand U14889 (N_14889,N_8015,N_6104);
nand U14890 (N_14890,N_6340,N_6797);
nor U14891 (N_14891,N_6231,N_5804);
nor U14892 (N_14892,N_5307,N_7545);
or U14893 (N_14893,N_8100,N_7319);
nor U14894 (N_14894,N_6913,N_8623);
or U14895 (N_14895,N_7668,N_5403);
or U14896 (N_14896,N_7911,N_5151);
and U14897 (N_14897,N_6893,N_7395);
or U14898 (N_14898,N_7177,N_9327);
and U14899 (N_14899,N_8500,N_9864);
and U14900 (N_14900,N_9160,N_6988);
nor U14901 (N_14901,N_9321,N_9379);
nand U14902 (N_14902,N_7791,N_9027);
nand U14903 (N_14903,N_5582,N_8891);
xor U14904 (N_14904,N_7211,N_8670);
nor U14905 (N_14905,N_8929,N_7145);
nor U14906 (N_14906,N_6918,N_8491);
nand U14907 (N_14907,N_7332,N_8904);
and U14908 (N_14908,N_7971,N_5796);
nor U14909 (N_14909,N_9191,N_5998);
and U14910 (N_14910,N_8986,N_6182);
xnor U14911 (N_14911,N_9089,N_5703);
nor U14912 (N_14912,N_6914,N_8758);
nand U14913 (N_14913,N_6483,N_6417);
nand U14914 (N_14914,N_8473,N_8112);
nor U14915 (N_14915,N_5798,N_9439);
nor U14916 (N_14916,N_7910,N_6701);
and U14917 (N_14917,N_9380,N_8162);
nor U14918 (N_14918,N_7849,N_9529);
nand U14919 (N_14919,N_9566,N_9501);
or U14920 (N_14920,N_7843,N_6344);
and U14921 (N_14921,N_7806,N_7409);
nor U14922 (N_14922,N_5395,N_5736);
and U14923 (N_14923,N_5350,N_9412);
xnor U14924 (N_14924,N_8307,N_7941);
nand U14925 (N_14925,N_7240,N_8494);
nand U14926 (N_14926,N_8879,N_7597);
and U14927 (N_14927,N_5590,N_8416);
or U14928 (N_14928,N_7888,N_6399);
xnor U14929 (N_14929,N_5538,N_8815);
nor U14930 (N_14930,N_9457,N_9261);
nand U14931 (N_14931,N_5843,N_7231);
or U14932 (N_14932,N_7994,N_8816);
and U14933 (N_14933,N_5989,N_9881);
or U14934 (N_14934,N_6824,N_6740);
and U14935 (N_14935,N_6469,N_5040);
nand U14936 (N_14936,N_6492,N_7980);
nand U14937 (N_14937,N_9484,N_6926);
nor U14938 (N_14938,N_5428,N_9145);
nand U14939 (N_14939,N_5234,N_9958);
or U14940 (N_14940,N_8444,N_6904);
nand U14941 (N_14941,N_6417,N_7943);
nor U14942 (N_14942,N_8711,N_7153);
nor U14943 (N_14943,N_5495,N_7497);
or U14944 (N_14944,N_8332,N_6807);
nand U14945 (N_14945,N_8186,N_6511);
nor U14946 (N_14946,N_7383,N_6156);
nand U14947 (N_14947,N_7036,N_6506);
xnor U14948 (N_14948,N_7967,N_6888);
or U14949 (N_14949,N_9815,N_8772);
or U14950 (N_14950,N_5846,N_5555);
nor U14951 (N_14951,N_5365,N_8863);
and U14952 (N_14952,N_7611,N_8792);
nor U14953 (N_14953,N_8489,N_6826);
nor U14954 (N_14954,N_6602,N_7054);
and U14955 (N_14955,N_9375,N_8953);
or U14956 (N_14956,N_8413,N_6596);
nand U14957 (N_14957,N_8377,N_8821);
xnor U14958 (N_14958,N_7014,N_6289);
and U14959 (N_14959,N_6281,N_8418);
nand U14960 (N_14960,N_8941,N_8653);
or U14961 (N_14961,N_9739,N_7628);
and U14962 (N_14962,N_9773,N_7461);
or U14963 (N_14963,N_6610,N_9957);
nor U14964 (N_14964,N_6127,N_6019);
nand U14965 (N_14965,N_9908,N_9144);
or U14966 (N_14966,N_5624,N_8684);
and U14967 (N_14967,N_7267,N_8629);
nand U14968 (N_14968,N_9077,N_6247);
nor U14969 (N_14969,N_7991,N_6996);
or U14970 (N_14970,N_6741,N_6014);
and U14971 (N_14971,N_9383,N_7165);
and U14972 (N_14972,N_9030,N_5522);
and U14973 (N_14973,N_7040,N_6051);
and U14974 (N_14974,N_7218,N_7987);
nand U14975 (N_14975,N_8942,N_9530);
nand U14976 (N_14976,N_6076,N_8067);
nor U14977 (N_14977,N_5591,N_9491);
nand U14978 (N_14978,N_8866,N_9263);
and U14979 (N_14979,N_6157,N_9062);
and U14980 (N_14980,N_6271,N_6143);
nor U14981 (N_14981,N_8465,N_7559);
or U14982 (N_14982,N_8455,N_8645);
and U14983 (N_14983,N_8307,N_5999);
or U14984 (N_14984,N_8750,N_8473);
and U14985 (N_14985,N_7775,N_6736);
nand U14986 (N_14986,N_5802,N_9257);
and U14987 (N_14987,N_7223,N_9727);
nor U14988 (N_14988,N_5877,N_5901);
or U14989 (N_14989,N_8458,N_7156);
xnor U14990 (N_14990,N_9626,N_7669);
or U14991 (N_14991,N_6283,N_6150);
and U14992 (N_14992,N_9199,N_7020);
and U14993 (N_14993,N_5487,N_5912);
nor U14994 (N_14994,N_6182,N_5512);
nand U14995 (N_14995,N_5565,N_9330);
and U14996 (N_14996,N_9295,N_7921);
nor U14997 (N_14997,N_7000,N_5940);
and U14998 (N_14998,N_8083,N_9123);
and U14999 (N_14999,N_6588,N_6652);
nand U15000 (N_15000,N_11411,N_12712);
nor U15001 (N_15001,N_10027,N_13689);
and U15002 (N_15002,N_14430,N_13187);
and U15003 (N_15003,N_11238,N_13300);
nand U15004 (N_15004,N_10291,N_11669);
or U15005 (N_15005,N_10545,N_11444);
and U15006 (N_15006,N_13537,N_14926);
nor U15007 (N_15007,N_11553,N_12486);
or U15008 (N_15008,N_12100,N_11775);
or U15009 (N_15009,N_14773,N_10957);
nand U15010 (N_15010,N_12964,N_11485);
or U15011 (N_15011,N_12250,N_10196);
xnor U15012 (N_15012,N_14275,N_11740);
nand U15013 (N_15013,N_12698,N_13185);
and U15014 (N_15014,N_14972,N_10202);
nand U15015 (N_15015,N_11217,N_14477);
or U15016 (N_15016,N_13433,N_11780);
and U15017 (N_15017,N_10643,N_13457);
and U15018 (N_15018,N_13268,N_14429);
and U15019 (N_15019,N_12848,N_13235);
nand U15020 (N_15020,N_14579,N_12907);
or U15021 (N_15021,N_14688,N_14953);
or U15022 (N_15022,N_10433,N_11715);
and U15023 (N_15023,N_14921,N_11713);
nor U15024 (N_15024,N_14223,N_13744);
and U15025 (N_15025,N_10841,N_10096);
and U15026 (N_15026,N_14603,N_11505);
nor U15027 (N_15027,N_14088,N_12642);
nand U15028 (N_15028,N_13984,N_14628);
and U15029 (N_15029,N_12366,N_12609);
or U15030 (N_15030,N_12011,N_14296);
or U15031 (N_15031,N_14336,N_13389);
nor U15032 (N_15032,N_13461,N_11470);
or U15033 (N_15033,N_11144,N_13327);
nand U15034 (N_15034,N_13378,N_12411);
or U15035 (N_15035,N_12394,N_12413);
nor U15036 (N_15036,N_12565,N_14441);
and U15037 (N_15037,N_13473,N_13896);
and U15038 (N_15038,N_12897,N_11201);
and U15039 (N_15039,N_13617,N_14558);
and U15040 (N_15040,N_14857,N_13421);
or U15041 (N_15041,N_12158,N_12781);
and U15042 (N_15042,N_14616,N_11628);
nand U15043 (N_15043,N_10970,N_13898);
nor U15044 (N_15044,N_10154,N_13644);
xnor U15045 (N_15045,N_10214,N_14484);
nor U15046 (N_15046,N_11325,N_11310);
nand U15047 (N_15047,N_13771,N_14847);
nand U15048 (N_15048,N_10902,N_10183);
nand U15049 (N_15049,N_10699,N_11971);
nor U15050 (N_15050,N_12713,N_10247);
xor U15051 (N_15051,N_13529,N_11951);
and U15052 (N_15052,N_13347,N_11253);
nor U15053 (N_15053,N_12311,N_12336);
xnor U15054 (N_15054,N_10439,N_10157);
and U15055 (N_15055,N_14987,N_10672);
nor U15056 (N_15056,N_14594,N_13713);
or U15057 (N_15057,N_12912,N_13386);
nand U15058 (N_15058,N_11825,N_13346);
and U15059 (N_15059,N_13836,N_12150);
xor U15060 (N_15060,N_11763,N_12408);
nor U15061 (N_15061,N_10769,N_13686);
or U15062 (N_15062,N_11586,N_10899);
xnor U15063 (N_15063,N_11524,N_10285);
nand U15064 (N_15064,N_14500,N_10537);
nor U15065 (N_15065,N_12023,N_11578);
xnor U15066 (N_15066,N_11865,N_12281);
nand U15067 (N_15067,N_13994,N_14333);
and U15068 (N_15068,N_11317,N_11909);
and U15069 (N_15069,N_11748,N_14174);
or U15070 (N_15070,N_14421,N_11620);
nand U15071 (N_15071,N_11488,N_10720);
or U15072 (N_15072,N_11937,N_10849);
and U15073 (N_15073,N_12242,N_12002);
or U15074 (N_15074,N_10279,N_11895);
and U15075 (N_15075,N_12485,N_14766);
or U15076 (N_15076,N_13980,N_14329);
nor U15077 (N_15077,N_14298,N_14013);
and U15078 (N_15078,N_11641,N_13930);
or U15079 (N_15079,N_12490,N_10907);
nor U15080 (N_15080,N_14747,N_12299);
xor U15081 (N_15081,N_11782,N_14540);
nand U15082 (N_15082,N_13171,N_12787);
and U15083 (N_15083,N_14597,N_10510);
and U15084 (N_15084,N_14991,N_10332);
nand U15085 (N_15085,N_11176,N_11543);
xor U15086 (N_15086,N_12314,N_10414);
nor U15087 (N_15087,N_13483,N_11428);
or U15088 (N_15088,N_11001,N_13650);
or U15089 (N_15089,N_11806,N_14533);
nand U15090 (N_15090,N_10138,N_12559);
xor U15091 (N_15091,N_11124,N_14576);
or U15092 (N_15092,N_12248,N_13523);
or U15093 (N_15093,N_10233,N_10634);
nand U15094 (N_15094,N_13586,N_11860);
xor U15095 (N_15095,N_14053,N_12544);
nor U15096 (N_15096,N_12159,N_12994);
nor U15097 (N_15097,N_12106,N_14376);
and U15098 (N_15098,N_10225,N_13398);
nor U15099 (N_15099,N_10996,N_10249);
or U15100 (N_15100,N_13520,N_12228);
or U15101 (N_15101,N_14056,N_14514);
xnor U15102 (N_15102,N_11634,N_13753);
and U15103 (N_15103,N_10175,N_11489);
nand U15104 (N_15104,N_10399,N_10761);
and U15105 (N_15105,N_12518,N_10724);
or U15106 (N_15106,N_10756,N_11929);
or U15107 (N_15107,N_10390,N_12447);
nand U15108 (N_15108,N_13897,N_13556);
nor U15109 (N_15109,N_10264,N_10230);
nor U15110 (N_15110,N_14645,N_12017);
nor U15111 (N_15111,N_14983,N_11548);
or U15112 (N_15112,N_11521,N_10254);
or U15113 (N_15113,N_12693,N_13392);
and U15114 (N_15114,N_12013,N_13033);
nor U15115 (N_15115,N_13008,N_12995);
nand U15116 (N_15116,N_10205,N_11894);
nand U15117 (N_15117,N_10095,N_11550);
nor U15118 (N_15118,N_14145,N_12162);
and U15119 (N_15119,N_13851,N_12445);
nor U15120 (N_15120,N_11472,N_12985);
nor U15121 (N_15121,N_10073,N_12245);
and U15122 (N_15122,N_13338,N_13237);
nand U15123 (N_15123,N_12819,N_10598);
nor U15124 (N_15124,N_11527,N_10698);
nor U15125 (N_15125,N_14444,N_10939);
and U15126 (N_15126,N_12603,N_14982);
or U15127 (N_15127,N_10728,N_13855);
and U15128 (N_15128,N_14212,N_11831);
and U15129 (N_15129,N_10586,N_11816);
nand U15130 (N_15130,N_12719,N_10409);
and U15131 (N_15131,N_14319,N_14506);
xor U15132 (N_15132,N_10870,N_14709);
or U15133 (N_15133,N_12771,N_12662);
and U15134 (N_15134,N_14570,N_10029);
xor U15135 (N_15135,N_13286,N_10132);
or U15136 (N_15136,N_14745,N_14961);
nor U15137 (N_15137,N_11299,N_12058);
nor U15138 (N_15138,N_11027,N_11792);
nand U15139 (N_15139,N_10003,N_13364);
nor U15140 (N_15140,N_12667,N_14634);
or U15141 (N_15141,N_14339,N_10402);
xnor U15142 (N_15142,N_13506,N_10393);
and U15143 (N_15143,N_14101,N_12628);
nor U15144 (N_15144,N_10516,N_11965);
and U15145 (N_15145,N_11762,N_10014);
xor U15146 (N_15146,N_14104,N_13647);
or U15147 (N_15147,N_14064,N_13472);
or U15148 (N_15148,N_10497,N_12085);
nor U15149 (N_15149,N_14633,N_12515);
or U15150 (N_15150,N_12836,N_14572);
nand U15151 (N_15151,N_13569,N_14998);
and U15152 (N_15152,N_10199,N_14496);
nand U15153 (N_15153,N_13165,N_13368);
nor U15154 (N_15154,N_10848,N_12786);
nand U15155 (N_15155,N_14789,N_14111);
nand U15156 (N_15156,N_10991,N_12643);
and U15157 (N_15157,N_12071,N_12065);
nand U15158 (N_15158,N_10059,N_11643);
xor U15159 (N_15159,N_11019,N_11439);
and U15160 (N_15160,N_11468,N_11513);
nor U15161 (N_15161,N_14050,N_11417);
nand U15162 (N_15162,N_14940,N_12549);
xnor U15163 (N_15163,N_11519,N_13273);
or U15164 (N_15164,N_13919,N_12292);
xnor U15165 (N_15165,N_12127,N_12444);
nand U15166 (N_15166,N_13222,N_14286);
and U15167 (N_15167,N_10747,N_11555);
and U15168 (N_15168,N_13833,N_11642);
and U15169 (N_15169,N_11572,N_13721);
or U15170 (N_15170,N_14793,N_10740);
xor U15171 (N_15171,N_10385,N_11083);
nand U15172 (N_15172,N_11125,N_10511);
nand U15173 (N_15173,N_12844,N_13720);
and U15174 (N_15174,N_13212,N_12332);
nand U15175 (N_15175,N_10033,N_11646);
nand U15176 (N_15176,N_12420,N_10024);
and U15177 (N_15177,N_10922,N_11229);
or U15178 (N_15178,N_13487,N_11033);
and U15179 (N_15179,N_11153,N_14650);
nand U15180 (N_15180,N_10321,N_14011);
nand U15181 (N_15181,N_10182,N_10198);
or U15182 (N_15182,N_14000,N_10811);
or U15183 (N_15183,N_10415,N_12126);
nand U15184 (N_15184,N_12689,N_13153);
nand U15185 (N_15185,N_12102,N_11370);
nor U15186 (N_15186,N_11645,N_11295);
and U15187 (N_15187,N_11529,N_10804);
or U15188 (N_15188,N_10591,N_11462);
or U15189 (N_15189,N_12913,N_13901);
or U15190 (N_15190,N_12756,N_10464);
or U15191 (N_15191,N_12562,N_11047);
nand U15192 (N_15192,N_12412,N_14031);
and U15193 (N_15193,N_14621,N_11644);
nand U15194 (N_15194,N_13439,N_13615);
and U15195 (N_15195,N_11157,N_11629);
nand U15196 (N_15196,N_11293,N_11461);
or U15197 (N_15197,N_13460,N_13240);
and U15198 (N_15198,N_10831,N_13942);
and U15199 (N_15199,N_10457,N_14677);
nor U15200 (N_15200,N_12234,N_11403);
or U15201 (N_15201,N_13290,N_11191);
nor U15202 (N_15202,N_13757,N_11708);
nand U15203 (N_15203,N_10584,N_12845);
and U15204 (N_15204,N_11577,N_12355);
nor U15205 (N_15205,N_13755,N_10885);
nand U15206 (N_15206,N_12685,N_12574);
and U15207 (N_15207,N_14358,N_12840);
nor U15208 (N_15208,N_12797,N_14055);
and U15209 (N_15209,N_14911,N_12846);
xor U15210 (N_15210,N_12051,N_11236);
nand U15211 (N_15211,N_14612,N_13043);
nor U15212 (N_15212,N_12620,N_10967);
nand U15213 (N_15213,N_13479,N_12144);
nand U15214 (N_15214,N_11009,N_10891);
nor U15215 (N_15215,N_13913,N_14534);
xnor U15216 (N_15216,N_11766,N_10575);
nand U15217 (N_15217,N_12596,N_12961);
nand U15218 (N_15218,N_12962,N_12927);
nand U15219 (N_15219,N_11297,N_12956);
nand U15220 (N_15220,N_11423,N_10734);
nand U15221 (N_15221,N_10370,N_10859);
nand U15222 (N_15222,N_10383,N_10641);
xor U15223 (N_15223,N_10572,N_13694);
nand U15224 (N_15224,N_13707,N_11649);
or U15225 (N_15225,N_14697,N_12225);
nand U15226 (N_15226,N_14837,N_10937);
and U15227 (N_15227,N_10297,N_13160);
and U15228 (N_15228,N_13480,N_11898);
or U15229 (N_15229,N_11023,N_12438);
nor U15230 (N_15230,N_14620,N_12590);
and U15231 (N_15231,N_12572,N_14306);
nor U15232 (N_15232,N_14505,N_11526);
nand U15233 (N_15233,N_12754,N_10451);
nand U15234 (N_15234,N_14277,N_13403);
nor U15235 (N_15235,N_10305,N_13061);
nor U15236 (N_15236,N_11061,N_11610);
nor U15237 (N_15237,N_12465,N_12622);
nand U15238 (N_15238,N_11820,N_10077);
xor U15239 (N_15239,N_14185,N_13292);
or U15240 (N_15240,N_12570,N_10652);
xor U15241 (N_15241,N_13987,N_10887);
nand U15242 (N_15242,N_12732,N_11355);
nor U15243 (N_15243,N_13228,N_10100);
or U15244 (N_15244,N_13265,N_13001);
nor U15245 (N_15245,N_14191,N_14008);
and U15246 (N_15246,N_14573,N_11939);
or U15247 (N_15247,N_13939,N_13229);
nor U15248 (N_15248,N_12874,N_11114);
xor U15249 (N_15249,N_10889,N_13920);
nand U15250 (N_15250,N_14658,N_10422);
nand U15251 (N_15251,N_11041,N_14080);
nor U15252 (N_15252,N_13345,N_13832);
xor U15253 (N_15253,N_12774,N_11565);
and U15254 (N_15254,N_11626,N_11205);
and U15255 (N_15255,N_12676,N_11405);
or U15256 (N_15256,N_12006,N_14734);
xnor U15257 (N_15257,N_13447,N_14869);
or U15258 (N_15258,N_12267,N_10440);
nor U15259 (N_15259,N_10707,N_13779);
nand U15260 (N_15260,N_11387,N_11487);
nand U15261 (N_15261,N_12612,N_10267);
or U15262 (N_15262,N_11364,N_11227);
or U15263 (N_15263,N_12078,N_11060);
and U15264 (N_15264,N_14816,N_10093);
or U15265 (N_15265,N_12864,N_10362);
nor U15266 (N_15266,N_11322,N_13024);
nand U15267 (N_15267,N_13267,N_11950);
nand U15268 (N_15268,N_13734,N_10022);
or U15269 (N_15269,N_10133,N_10955);
nand U15270 (N_15270,N_12377,N_14760);
nor U15271 (N_15271,N_12548,N_14636);
and U15272 (N_15272,N_13010,N_11833);
nand U15273 (N_15273,N_13716,N_13761);
xnor U15274 (N_15274,N_14220,N_12328);
nor U15275 (N_15275,N_13937,N_10431);
nand U15276 (N_15276,N_14227,N_13515);
and U15277 (N_15277,N_10522,N_13969);
and U15278 (N_15278,N_11822,N_14164);
nor U15279 (N_15279,N_13785,N_11595);
and U15280 (N_15280,N_11535,N_11200);
nand U15281 (N_15281,N_11692,N_10592);
xor U15282 (N_15282,N_12826,N_14196);
nor U15283 (N_15283,N_14109,N_12876);
and U15284 (N_15284,N_13170,N_10054);
or U15285 (N_15285,N_14253,N_10412);
nor U15286 (N_15286,N_13105,N_13727);
and U15287 (N_15287,N_10074,N_10106);
xor U15288 (N_15288,N_14976,N_14459);
or U15289 (N_15289,N_14565,N_11085);
xor U15290 (N_15290,N_12316,N_10517);
nor U15291 (N_15291,N_14412,N_14876);
nand U15292 (N_15292,N_13636,N_14189);
or U15293 (N_15293,N_10913,N_12569);
and U15294 (N_15294,N_10169,N_11503);
nand U15295 (N_15295,N_13876,N_14973);
or U15296 (N_15296,N_10847,N_10644);
nand U15297 (N_15297,N_11188,N_12536);
or U15298 (N_15298,N_11148,N_13029);
or U15299 (N_15299,N_11434,N_10384);
or U15300 (N_15300,N_10723,N_12033);
xnor U15301 (N_15301,N_10371,N_13911);
nor U15302 (N_15302,N_10356,N_14165);
or U15303 (N_15303,N_13294,N_12546);
and U15304 (N_15304,N_13053,N_14874);
nor U15305 (N_15305,N_14786,N_10441);
and U15306 (N_15306,N_13302,N_14963);
nor U15307 (N_15307,N_10338,N_10901);
nand U15308 (N_15308,N_14903,N_12340);
nor U15309 (N_15309,N_11953,N_10231);
nor U15310 (N_15310,N_13603,N_14517);
and U15311 (N_15311,N_10705,N_12296);
or U15312 (N_15312,N_12429,N_10752);
or U15313 (N_15313,N_11700,N_12744);
nand U15314 (N_15314,N_14167,N_10969);
nand U15315 (N_15315,N_11309,N_12313);
or U15316 (N_15316,N_12837,N_10349);
and U15317 (N_15317,N_10374,N_11465);
or U15318 (N_15318,N_12246,N_14784);
or U15319 (N_15319,N_13830,N_13655);
nor U15320 (N_15320,N_13084,N_14831);
and U15321 (N_15321,N_12257,N_14575);
nor U15322 (N_15322,N_11680,N_11290);
and U15323 (N_15323,N_13527,N_12926);
nand U15324 (N_15324,N_10259,N_12911);
or U15325 (N_15325,N_13651,N_13807);
nor U15326 (N_15326,N_11324,N_13058);
nand U15327 (N_15327,N_11506,N_12908);
nand U15328 (N_15328,N_10315,N_12860);
and U15329 (N_15329,N_14622,N_11924);
or U15330 (N_15330,N_14807,N_10442);
nor U15331 (N_15331,N_11873,N_13357);
nor U15332 (N_15332,N_13236,N_12859);
or U15333 (N_15333,N_11025,N_11437);
and U15334 (N_15334,N_14966,N_14691);
and U15335 (N_15335,N_10005,N_13320);
or U15336 (N_15336,N_12714,N_14927);
nor U15337 (N_15337,N_12042,N_14885);
nand U15338 (N_15338,N_10051,N_14992);
and U15339 (N_15339,N_12809,N_12831);
xnor U15340 (N_15340,N_14654,N_12309);
nor U15341 (N_15341,N_12858,N_13289);
nand U15342 (N_15342,N_11129,N_13441);
and U15343 (N_15343,N_10987,N_14450);
nand U15344 (N_15344,N_11976,N_13540);
nor U15345 (N_15345,N_14311,N_10917);
or U15346 (N_15346,N_13384,N_11016);
and U15347 (N_15347,N_10799,N_10058);
nor U15348 (N_15348,N_12645,N_13217);
nor U15349 (N_15349,N_10481,N_14610);
nor U15350 (N_15350,N_13477,N_14556);
nand U15351 (N_15351,N_11852,N_11522);
nor U15352 (N_15352,N_10524,N_11562);
and U15353 (N_15353,N_14454,N_12414);
and U15354 (N_15354,N_12386,N_13178);
nand U15355 (N_15355,N_11908,N_11834);
or U15356 (N_15356,N_10118,N_12200);
and U15357 (N_15357,N_12323,N_12482);
or U15358 (N_15358,N_14110,N_13835);
and U15359 (N_15359,N_11093,N_12416);
nor U15360 (N_15360,N_12816,N_12540);
xnor U15361 (N_15361,N_10428,N_12910);
nand U15362 (N_15362,N_12887,N_11265);
nor U15363 (N_15363,N_14646,N_14467);
nand U15364 (N_15364,N_12221,N_10235);
and U15365 (N_15365,N_12532,N_11804);
nor U15366 (N_15366,N_10026,N_11549);
nor U15367 (N_15367,N_10025,N_11720);
or U15368 (N_15368,N_12492,N_11788);
or U15369 (N_15369,N_12675,N_14855);
and U15370 (N_15370,N_11768,N_10373);
and U15371 (N_15371,N_13900,N_11277);
nor U15372 (N_15372,N_10166,N_10762);
nand U15373 (N_15373,N_10709,N_11162);
nor U15374 (N_15374,N_14337,N_10558);
nor U15375 (N_15375,N_10469,N_11547);
and U15376 (N_15376,N_11271,N_14026);
or U15377 (N_15377,N_10978,N_13844);
nand U15378 (N_15378,N_14070,N_13431);
xor U15379 (N_15379,N_14170,N_10623);
nor U15380 (N_15380,N_10858,N_14303);
and U15381 (N_15381,N_14737,N_10306);
nor U15382 (N_15382,N_14407,N_11486);
xor U15383 (N_15383,N_12959,N_13632);
xnor U15384 (N_15384,N_12352,N_13997);
nor U15385 (N_15385,N_11255,N_13348);
nand U15386 (N_15386,N_14977,N_10821);
nor U15387 (N_15387,N_10964,N_11028);
nor U15388 (N_15388,N_13576,N_11589);
nor U15389 (N_15389,N_11518,N_11818);
nand U15390 (N_15390,N_10304,N_14001);
nor U15391 (N_15391,N_11131,N_10430);
nand U15392 (N_15392,N_10452,N_13780);
or U15393 (N_15393,N_12094,N_11326);
nand U15394 (N_15394,N_10678,N_11542);
and U15395 (N_15395,N_10193,N_13372);
or U15396 (N_15396,N_13322,N_13607);
nand U15397 (N_15397,N_14346,N_12695);
nor U15398 (N_15398,N_10561,N_12119);
nand U15399 (N_15399,N_13739,N_14822);
nand U15400 (N_15400,N_12432,N_12004);
nor U15401 (N_15401,N_13206,N_11625);
nor U15402 (N_15402,N_10764,N_11070);
and U15403 (N_15403,N_11099,N_11197);
nor U15404 (N_15404,N_12624,N_14340);
nand U15405 (N_15405,N_12745,N_12101);
nor U15406 (N_15406,N_11911,N_12778);
and U15407 (N_15407,N_10019,N_13138);
nand U15408 (N_15408,N_13099,N_14527);
nand U15409 (N_15409,N_12294,N_13124);
or U15410 (N_15410,N_11225,N_10485);
and U15411 (N_15411,N_11655,N_12066);
and U15412 (N_15412,N_13137,N_14664);
nand U15413 (N_15413,N_12568,N_12358);
nor U15414 (N_15414,N_14873,N_12271);
nor U15415 (N_15415,N_13554,N_14492);
nor U15416 (N_15416,N_12284,N_13552);
and U15417 (N_15417,N_14529,N_10681);
nand U15418 (N_15418,N_14959,N_10039);
nand U15419 (N_15419,N_12625,N_12584);
nand U15420 (N_15420,N_13422,N_14711);
or U15421 (N_15421,N_13250,N_12951);
or U15422 (N_15422,N_12210,N_13979);
nor U15423 (N_15423,N_12027,N_11583);
or U15424 (N_15424,N_11109,N_13856);
or U15425 (N_15425,N_14845,N_10629);
or U15426 (N_15426,N_12026,N_11422);
nand U15427 (N_15427,N_11116,N_11564);
and U15428 (N_15428,N_14330,N_13108);
or U15429 (N_15429,N_14866,N_14268);
or U15430 (N_15430,N_11560,N_13799);
nor U15431 (N_15431,N_14653,N_14510);
xor U15432 (N_15432,N_11632,N_11308);
and U15433 (N_15433,N_10031,N_10851);
or U15434 (N_15434,N_12674,N_14769);
or U15435 (N_15435,N_10703,N_10742);
nand U15436 (N_15436,N_13884,N_12318);
and U15437 (N_15437,N_10161,N_10053);
or U15438 (N_15438,N_12180,N_10296);
nor U15439 (N_15439,N_14962,N_13623);
and U15440 (N_15440,N_10613,N_12141);
nand U15441 (N_15441,N_10237,N_10590);
or U15442 (N_15442,N_14875,N_11545);
nand U15443 (N_15443,N_11686,N_13886);
and U15444 (N_15444,N_10540,N_11160);
nor U15445 (N_15445,N_11685,N_12512);
and U15446 (N_15446,N_12894,N_10737);
nand U15447 (N_15447,N_10513,N_14539);
nor U15448 (N_15448,N_14373,N_10695);
and U15449 (N_15449,N_12702,N_10805);
or U15450 (N_15450,N_10472,N_12049);
or U15451 (N_15451,N_13704,N_11280);
nand U15452 (N_15452,N_14958,N_13974);
nand U15453 (N_15453,N_11404,N_11474);
nand U15454 (N_15454,N_14686,N_12151);
and U15455 (N_15455,N_12178,N_13588);
nand U15456 (N_15456,N_13555,N_12153);
and U15457 (N_15457,N_10097,N_12524);
and U15458 (N_15458,N_13107,N_14393);
nor U15459 (N_15459,N_12588,N_10162);
nor U15460 (N_15460,N_12830,N_14599);
nand U15461 (N_15461,N_13600,N_12325);
or U15462 (N_15462,N_12436,N_11661);
or U15463 (N_15463,N_10671,N_14578);
and U15464 (N_15464,N_12602,N_10413);
nand U15465 (N_15465,N_10768,N_11544);
and U15466 (N_15466,N_14904,N_12715);
xor U15467 (N_15467,N_11668,N_11399);
nor U15468 (N_15468,N_14217,N_12480);
nor U15469 (N_15469,N_12982,N_14954);
or U15470 (N_15470,N_13400,N_14730);
nor U15471 (N_15471,N_12456,N_11314);
nand U15472 (N_15472,N_12883,N_13245);
nor U15473 (N_15473,N_13924,N_11838);
and U15474 (N_15474,N_14133,N_11126);
and U15475 (N_15475,N_13085,N_13109);
xor U15476 (N_15476,N_14928,N_13711);
or U15477 (N_15477,N_11246,N_10176);
nand U15478 (N_15478,N_12788,N_10823);
nand U15479 (N_15479,N_12670,N_11427);
and U15480 (N_15480,N_10525,N_13745);
and U15481 (N_15481,N_14938,N_13630);
nand U15482 (N_15482,N_12160,N_11879);
xnor U15483 (N_15483,N_13567,N_12811);
xnor U15484 (N_15484,N_14061,N_13680);
nand U15485 (N_15485,N_12262,N_13356);
nor U15486 (N_15486,N_14071,N_11738);
nand U15487 (N_15487,N_14649,N_12498);
nand U15488 (N_15488,N_11262,N_12396);
or U15489 (N_15489,N_13113,N_11758);
nand U15490 (N_15490,N_10324,N_10815);
nand U15491 (N_15491,N_12939,N_11863);
nand U15492 (N_15492,N_13111,N_12497);
or U15493 (N_15493,N_11946,N_12882);
or U15494 (N_15494,N_14304,N_14915);
or U15495 (N_15495,N_12946,N_14965);
xor U15496 (N_15496,N_12750,N_11330);
nor U15497 (N_15497,N_12130,N_14968);
nand U15498 (N_15498,N_14399,N_10090);
nand U15499 (N_15499,N_12729,N_11603);
or U15500 (N_15500,N_14537,N_11471);
and U15501 (N_15501,N_10245,N_11793);
nand U15502 (N_15502,N_10796,N_10527);
nand U15503 (N_15503,N_13452,N_12400);
nor U15504 (N_15504,N_13601,N_13216);
and U15505 (N_15505,N_13722,N_10844);
and U15506 (N_15506,N_12466,N_11492);
xor U15507 (N_15507,N_10108,N_11866);
or U15508 (N_15508,N_14432,N_12827);
xnor U15509 (N_15509,N_11789,N_10581);
nand U15510 (N_15510,N_11258,N_14974);
and U15511 (N_15511,N_11659,N_10521);
nor U15512 (N_15512,N_10462,N_12889);
nor U15513 (N_15513,N_13145,N_11004);
nand U15514 (N_15514,N_10350,N_11102);
nand U15515 (N_15515,N_14986,N_10392);
nand U15516 (N_15516,N_10866,N_12261);
and U15517 (N_15517,N_11613,N_10213);
nor U15518 (N_15518,N_12566,N_12555);
nand U15519 (N_15519,N_14595,N_13354);
or U15520 (N_15520,N_14726,N_13343);
nand U15521 (N_15521,N_12092,N_10755);
nor U15522 (N_15522,N_14232,N_12391);
nand U15523 (N_15523,N_14946,N_10347);
nor U15524 (N_15524,N_11958,N_11755);
nor U15525 (N_15525,N_13989,N_13183);
xor U15526 (N_15526,N_13004,N_14809);
nor U15527 (N_15527,N_14435,N_10048);
and U15528 (N_15528,N_13975,N_10710);
nor U15529 (N_15529,N_12746,N_10673);
nand U15530 (N_15530,N_13710,N_13428);
and U15531 (N_15531,N_14468,N_10933);
nand U15532 (N_15532,N_14117,N_10461);
nor U15533 (N_15533,N_12468,N_13661);
nor U15534 (N_15534,N_13618,N_14497);
nand U15535 (N_15535,N_11663,N_11523);
nand U15536 (N_15536,N_12315,N_11960);
nand U15537 (N_15537,N_13864,N_14367);
and U15538 (N_15538,N_11249,N_10329);
nand U15539 (N_15539,N_11491,N_13380);
nor U15540 (N_15540,N_11388,N_12765);
xor U15541 (N_15541,N_10261,N_11968);
and U15542 (N_15542,N_12381,N_10223);
nand U15543 (N_15543,N_13512,N_14345);
xor U15544 (N_15544,N_10078,N_14759);
nand U15545 (N_15545,N_12129,N_12156);
or U15546 (N_15546,N_12843,N_12998);
and U15547 (N_15547,N_11746,N_14062);
or U15548 (N_15548,N_10126,N_13926);
xnor U15549 (N_15549,N_13990,N_12499);
xnor U15550 (N_15550,N_10606,N_13080);
nor U15551 (N_15551,N_13015,N_13594);
or U15552 (N_15552,N_13585,N_13735);
or U15553 (N_15553,N_12025,N_14841);
or U15554 (N_15554,N_10448,N_12691);
nand U15555 (N_15555,N_12716,N_11426);
nand U15556 (N_15556,N_11218,N_10850);
and U15557 (N_15557,N_12365,N_11594);
nor U15558 (N_15558,N_14222,N_14491);
nor U15559 (N_15559,N_13619,N_14416);
nand U15560 (N_15560,N_14201,N_10153);
and U15561 (N_15561,N_12503,N_14828);
and U15562 (N_15562,N_14630,N_10395);
nor U15563 (N_15563,N_12052,N_14864);
and U15564 (N_15564,N_13196,N_12981);
or U15565 (N_15565,N_14072,N_12280);
nor U15566 (N_15566,N_10144,N_14518);
xor U15567 (N_15567,N_13469,N_14318);
and U15568 (N_15568,N_11985,N_11961);
or U15569 (N_15569,N_13792,N_14979);
nor U15570 (N_15570,N_10170,N_10063);
and U15571 (N_15571,N_14755,N_14402);
and U15572 (N_15572,N_10316,N_11261);
nand U15573 (N_15573,N_11182,N_14370);
xnor U15574 (N_15574,N_10824,N_14933);
or U15575 (N_15575,N_10921,N_14900);
and U15576 (N_15576,N_13157,N_14181);
or U15577 (N_15577,N_12247,N_13125);
and U15578 (N_15578,N_11231,N_11409);
nand U15579 (N_15579,N_10042,N_13430);
nand U15580 (N_15580,N_13494,N_11921);
xor U15581 (N_15581,N_14398,N_12270);
nand U15582 (N_15582,N_11637,N_13970);
or U15583 (N_15583,N_11602,N_10295);
or U15584 (N_15584,N_10625,N_14350);
or U15585 (N_15585,N_12880,N_12808);
nor U15586 (N_15586,N_10318,N_11005);
nor U15587 (N_15587,N_12551,N_13978);
and U15588 (N_15588,N_13489,N_13097);
and U15589 (N_15589,N_13867,N_14770);
nand U15590 (N_15590,N_13508,N_12891);
and U15591 (N_15591,N_12655,N_10785);
nor U15592 (N_15592,N_12020,N_11819);
and U15593 (N_15593,N_13243,N_11941);
nor U15594 (N_15594,N_13525,N_10836);
and U15595 (N_15595,N_11274,N_13119);
nand U15596 (N_15596,N_10493,N_14023);
and U15597 (N_15597,N_11432,N_13514);
or U15598 (N_15598,N_14899,N_13503);
and U15599 (N_15599,N_13582,N_10388);
xnor U15600 (N_15600,N_14929,N_13011);
and U15601 (N_15601,N_14571,N_14424);
nor U15602 (N_15602,N_11079,N_14812);
and U15603 (N_15603,N_13742,N_11240);
nand U15604 (N_15604,N_10416,N_10142);
and U15605 (N_15605,N_12426,N_14294);
or U15606 (N_15606,N_11151,N_14713);
xnor U15607 (N_15607,N_12552,N_12509);
nand U15608 (N_15608,N_14907,N_11257);
nor U15609 (N_15609,N_12348,N_11830);
and U15610 (N_15610,N_13663,N_13246);
or U15611 (N_15611,N_13458,N_13915);
nor U15612 (N_15612,N_13281,N_13412);
or U15613 (N_15613,N_12879,N_14551);
nand U15614 (N_15614,N_10786,N_10239);
nand U15615 (N_15615,N_13701,N_10334);
and U15616 (N_15616,N_14752,N_12139);
and U15617 (N_15617,N_12338,N_12265);
or U15618 (N_15618,N_12289,N_10868);
and U15619 (N_15619,N_12133,N_11846);
nor U15620 (N_15620,N_10856,N_11679);
nand U15621 (N_15621,N_14322,N_11055);
nand U15622 (N_15622,N_14820,N_14149);
nor U15623 (N_15623,N_12186,N_13642);
nand U15624 (N_15624,N_13093,N_11069);
and U15625 (N_15625,N_13775,N_14880);
xor U15626 (N_15626,N_12527,N_14910);
nand U15627 (N_15627,N_12967,N_13961);
xor U15628 (N_15628,N_10702,N_13808);
nor U15629 (N_15629,N_12700,N_14984);
or U15630 (N_15630,N_10156,N_12168);
or U15631 (N_15631,N_12339,N_10884);
nand U15632 (N_15632,N_13450,N_10708);
and U15633 (N_15633,N_14853,N_13350);
nand U15634 (N_15634,N_12099,N_13662);
xnor U15635 (N_15635,N_12048,N_11931);
and U15636 (N_15636,N_14944,N_11066);
xor U15637 (N_15637,N_13595,N_10878);
or U15638 (N_15638,N_13922,N_11998);
nand U15639 (N_15639,N_14700,N_10953);
xnor U15640 (N_15640,N_13221,N_14827);
nor U15641 (N_15641,N_14838,N_12505);
and U15642 (N_15642,N_12748,N_12673);
or U15643 (N_15643,N_12330,N_14592);
or U15644 (N_15644,N_14107,N_10911);
nand U15645 (N_15645,N_13883,N_12016);
nor U15646 (N_15646,N_12598,N_10299);
nand U15647 (N_15647,N_10344,N_13065);
or U15648 (N_15648,N_11494,N_14413);
nand U15649 (N_15649,N_12382,N_12560);
and U15650 (N_15650,N_13885,N_13194);
and U15651 (N_15651,N_14439,N_13259);
and U15652 (N_15652,N_12902,N_13823);
nor U15653 (N_15653,N_11704,N_12116);
or U15654 (N_15654,N_13628,N_13003);
nand U15655 (N_15655,N_13055,N_11759);
nor U15656 (N_15656,N_12968,N_12327);
xnor U15657 (N_15657,N_10207,N_13996);
xnor U15658 (N_15658,N_10380,N_14365);
xnor U15659 (N_15659,N_14442,N_10566);
and U15660 (N_15660,N_14160,N_10049);
and U15661 (N_15661,N_13032,N_14282);
nor U15662 (N_15662,N_10136,N_10314);
and U15663 (N_15663,N_11771,N_10131);
nand U15664 (N_15664,N_11809,N_12523);
nor U15665 (N_15665,N_12034,N_14487);
nand U15666 (N_15666,N_13511,N_11973);
nand U15667 (N_15667,N_11848,N_12259);
and U15668 (N_15668,N_10920,N_14623);
nor U15669 (N_15669,N_14131,N_14415);
nor U15670 (N_15670,N_11454,N_10281);
or U15671 (N_15671,N_11180,N_14395);
nand U15672 (N_15672,N_12564,N_11149);
or U15673 (N_15673,N_12415,N_14420);
or U15674 (N_15674,N_11982,N_12718);
or U15675 (N_15675,N_14455,N_14203);
or U15676 (N_15676,N_13714,N_10604);
nor U15677 (N_15677,N_10578,N_11441);
and U15678 (N_15678,N_14276,N_11107);
or U15679 (N_15679,N_11166,N_14130);
and U15680 (N_15680,N_12725,N_11135);
xor U15681 (N_15681,N_10236,N_13377);
nor U15682 (N_15682,N_11688,N_13411);
nor U15683 (N_15683,N_10122,N_11100);
nor U15684 (N_15684,N_12154,N_14051);
xnor U15685 (N_15685,N_11340,N_10532);
or U15686 (N_15686,N_10480,N_14419);
and U15687 (N_15687,N_11396,N_13130);
and U15688 (N_15688,N_13162,N_12901);
and U15689 (N_15689,N_11222,N_10676);
nor U15690 (N_15690,N_11015,N_14660);
nor U15691 (N_15691,N_11199,N_14155);
nor U15692 (N_15692,N_11536,N_10618);
nor U15693 (N_15693,N_12142,N_12735);
nand U15694 (N_15694,N_12072,N_13927);
and U15695 (N_15695,N_10150,N_14914);
or U15696 (N_15696,N_10611,N_11301);
and U15697 (N_15697,N_11394,N_10757);
and U15698 (N_15698,N_12201,N_13841);
or U15699 (N_15699,N_11460,N_14152);
or U15700 (N_15700,N_14166,N_11251);
xnor U15701 (N_15701,N_14768,N_14655);
nor U15702 (N_15702,N_11881,N_11773);
nor U15703 (N_15703,N_14359,N_11721);
nand U15704 (N_15704,N_14069,N_14719);
xnor U15705 (N_15705,N_11062,N_13271);
nor U15706 (N_15706,N_14731,N_13459);
and U15707 (N_15707,N_12188,N_13812);
nand U15708 (N_15708,N_13287,N_10529);
and U15709 (N_15709,N_12363,N_10429);
or U15710 (N_15710,N_14924,N_12790);
nor U15711 (N_15711,N_10986,N_11981);
nand U15712 (N_15712,N_11241,N_12767);
nor U15713 (N_15713,N_13798,N_13829);
and U15714 (N_15714,N_13025,N_14461);
nand U15715 (N_15715,N_13964,N_12886);
xnor U15716 (N_15716,N_12471,N_14426);
xnor U15717 (N_15717,N_11776,N_12354);
or U15718 (N_15718,N_10130,N_14471);
or U15719 (N_15719,N_12076,N_12448);
nor U15720 (N_15720,N_12388,N_10819);
nor U15721 (N_15721,N_11821,N_11321);
or U15722 (N_15722,N_13191,N_11779);
nor U15723 (N_15723,N_14017,N_10307);
xnor U15724 (N_15724,N_13249,N_14247);
and U15725 (N_15725,N_12211,N_14985);
and U15726 (N_15726,N_11612,N_13308);
or U15727 (N_15727,N_10091,N_12255);
and U15728 (N_15728,N_14640,N_11357);
and U15729 (N_15729,N_14392,N_12915);
or U15730 (N_15730,N_10006,N_10064);
nor U15731 (N_15731,N_12195,N_14079);
or U15732 (N_15732,N_10206,N_14006);
nand U15733 (N_15733,N_11743,N_11110);
nor U15734 (N_15734,N_13131,N_14543);
nand U15735 (N_15735,N_13468,N_10992);
and U15736 (N_15736,N_10877,N_12403);
nand U15737 (N_15737,N_14371,N_10379);
and U15738 (N_15738,N_13762,N_13394);
nand U15739 (N_15739,N_10248,N_14805);
nand U15740 (N_15740,N_10034,N_14067);
nand U15741 (N_15741,N_14931,N_11073);
nand U15742 (N_15742,N_14586,N_11215);
nand U15743 (N_15743,N_14761,N_10226);
nor U15744 (N_15744,N_11673,N_12418);
nand U15745 (N_15745,N_13417,N_10677);
nand U15746 (N_15746,N_12312,N_14835);
nand U15747 (N_15747,N_14685,N_13110);
nor U15748 (N_15748,N_11675,N_10682);
nand U15749 (N_15749,N_13009,N_11614);
nor U15750 (N_15750,N_11917,N_13935);
and U15751 (N_15751,N_13144,N_12112);
nor U15752 (N_15752,N_13828,N_11729);
nor U15753 (N_15753,N_13564,N_11447);
nand U15754 (N_15754,N_10779,N_13522);
nand U15755 (N_15755,N_13054,N_12495);
and U15756 (N_15756,N_14183,N_10990);
nor U15757 (N_15757,N_12899,N_14906);
nor U15758 (N_15758,N_10898,N_14321);
and U15759 (N_15759,N_13905,N_13986);
xnor U15760 (N_15760,N_11778,N_14695);
and U15761 (N_15761,N_11987,N_14290);
nor U15762 (N_15762,N_14014,N_13278);
and U15763 (N_15763,N_10265,N_14829);
nand U15764 (N_15764,N_14758,N_11377);
nor U15765 (N_15765,N_13593,N_13207);
and U15766 (N_15766,N_14662,N_11106);
nand U15767 (N_15767,N_14002,N_11091);
and U15768 (N_15768,N_13878,N_13341);
or U15769 (N_15769,N_10269,N_13899);
nor U15770 (N_15770,N_14048,N_11823);
nand U15771 (N_15771,N_10495,N_10112);
or U15772 (N_15772,N_10687,N_10477);
and U15773 (N_15773,N_13000,N_13132);
and U15774 (N_15774,N_11640,N_12164);
xnor U15775 (N_15775,N_10943,N_14867);
xor U15776 (N_15776,N_14886,N_11735);
nand U15777 (N_15777,N_13679,N_13559);
or U15778 (N_15778,N_10716,N_11674);
xnor U15779 (N_15779,N_10960,N_11358);
nor U15780 (N_15780,N_11540,N_14012);
and U15781 (N_15781,N_10119,N_14821);
or U15782 (N_15782,N_10534,N_11359);
or U15783 (N_15783,N_11630,N_13783);
nor U15784 (N_15784,N_12356,N_11760);
or U15785 (N_15785,N_10602,N_14241);
nand U15786 (N_15786,N_12404,N_12935);
nand U15787 (N_15787,N_13270,N_12446);
nand U15788 (N_15788,N_13225,N_14478);
nor U15789 (N_15789,N_12631,N_10931);
or U15790 (N_15790,N_14360,N_13326);
nor U15791 (N_15791,N_11861,N_11619);
nor U15792 (N_15792,N_10211,N_13598);
or U15793 (N_15793,N_14458,N_14956);
and U15794 (N_15794,N_14774,N_12738);
and U15795 (N_15795,N_13827,N_14211);
or U15796 (N_15796,N_13209,N_12184);
and U15797 (N_15797,N_14960,N_12114);
nor U15798 (N_15798,N_14798,N_12080);
or U15799 (N_15799,N_12766,N_10411);
nor U15800 (N_15800,N_10352,N_13284);
and U15801 (N_15801,N_12258,N_13749);
and U15802 (N_15802,N_12683,N_11223);
and U15803 (N_15803,N_13383,N_13786);
nand U15804 (N_15804,N_11412,N_14128);
nor U15805 (N_15805,N_14590,N_11347);
nand U15806 (N_15806,N_11193,N_11140);
xor U15807 (N_15807,N_14783,N_11288);
nand U15808 (N_15808,N_12230,N_14353);
xnor U15809 (N_15809,N_10526,N_10491);
and U15810 (N_15810,N_14937,N_11344);
and U15811 (N_15811,N_13141,N_12224);
xnor U15812 (N_15812,N_12081,N_14897);
nor U15813 (N_15813,N_14881,N_11169);
xnor U15814 (N_15814,N_12233,N_11117);
nor U15815 (N_15815,N_10741,N_14342);
nor U15816 (N_15816,N_10361,N_10980);
xnor U15817 (N_15817,N_10926,N_11178);
nand U15818 (N_15818,N_10055,N_13765);
or U15819 (N_15819,N_10504,N_12779);
and U15820 (N_15820,N_11751,N_11384);
or U15821 (N_15821,N_10387,N_10069);
and U15822 (N_15822,N_14118,N_13950);
and U15823 (N_15823,N_14794,N_12881);
and U15824 (N_15824,N_10549,N_14765);
and U15825 (N_15825,N_10330,N_12306);
nor U15826 (N_15826,N_12202,N_11035);
nand U15827 (N_15827,N_11925,N_10184);
nand U15828 (N_15828,N_10574,N_14908);
and U15829 (N_15829,N_11090,N_13825);
and U15830 (N_15830,N_13821,N_13002);
nand U15831 (N_15831,N_11017,N_14280);
nor U15832 (N_15832,N_10916,N_14638);
nor U15833 (N_15833,N_11071,N_10890);
and U15834 (N_15834,N_11291,N_10989);
or U15835 (N_15835,N_13624,N_11372);
nor U15836 (N_15836,N_12070,N_10056);
or U15837 (N_15837,N_12463,N_13752);
xnor U15838 (N_15838,N_12706,N_14153);
and U15839 (N_15839,N_10173,N_11877);
and U15840 (N_15840,N_10754,N_14357);
or U15841 (N_15841,N_11769,N_12708);
nor U15842 (N_15842,N_13040,N_13776);
and U15843 (N_15843,N_13039,N_10243);
xor U15844 (N_15844,N_13940,N_12571);
xnor U15845 (N_15845,N_13695,N_12256);
or U15846 (N_15846,N_12227,N_14482);
nor U15847 (N_15847,N_11136,N_11380);
nand U15848 (N_15848,N_13328,N_10816);
nor U15849 (N_15849,N_14692,N_12516);
nor U15850 (N_15850,N_12885,N_12374);
nand U15851 (N_15851,N_12617,N_10331);
nor U15852 (N_15852,N_10092,N_10194);
nand U15853 (N_15853,N_13255,N_13682);
nand U15854 (N_15854,N_11835,N_11279);
and U15855 (N_15855,N_10313,N_13768);
nor U15856 (N_15856,N_14611,N_13370);
or U15857 (N_15857,N_12108,N_12758);
nor U15858 (N_15858,N_12573,N_11051);
nor U15859 (N_15859,N_13404,N_10360);
nor U15860 (N_15860,N_12681,N_13973);
nand U15861 (N_15861,N_14870,N_14038);
nor U15862 (N_15862,N_12854,N_10121);
nand U15863 (N_15863,N_11232,N_12704);
nand U15864 (N_15864,N_11121,N_11747);
and U15865 (N_15865,N_13599,N_14862);
or U15866 (N_15866,N_11532,N_10983);
nand U15867 (N_15867,N_10007,N_10417);
or U15868 (N_15868,N_10910,N_14589);
or U15869 (N_15869,N_11798,N_11756);
nor U15870 (N_15870,N_12930,N_11170);
nand U15871 (N_15871,N_10272,N_10874);
nand U15872 (N_15872,N_10568,N_14913);
or U15873 (N_15873,N_12288,N_10600);
and U15874 (N_15874,N_14266,N_12455);
or U15875 (N_15875,N_13910,N_12193);
and U15876 (N_15876,N_13993,N_13658);
and U15877 (N_15877,N_12124,N_14473);
and U15878 (N_15878,N_10979,N_13437);
nand U15879 (N_15879,N_10904,N_14383);
and U15880 (N_15880,N_14113,N_11761);
xor U15881 (N_15881,N_11988,N_14659);
xnor U15882 (N_15882,N_11219,N_12975);
and U15883 (N_15883,N_12389,N_12740);
nor U15884 (N_15884,N_10909,N_12806);
and U15885 (N_15885,N_10881,N_10167);
or U15886 (N_15886,N_10478,N_13189);
nand U15887 (N_15887,N_11682,N_10776);
and U15888 (N_15888,N_11259,N_11590);
nor U15889 (N_15889,N_11021,N_13393);
or U15890 (N_15890,N_12373,N_10148);
nand U15891 (N_15891,N_11345,N_12909);
or U15892 (N_15892,N_11539,N_12847);
and U15893 (N_15893,N_11870,N_13129);
or U15894 (N_15894,N_13159,N_14052);
or U15895 (N_15895,N_13834,N_11420);
nor U15896 (N_15896,N_11057,N_11002);
nand U15897 (N_15897,N_14674,N_14374);
nor U15898 (N_15898,N_13826,N_11670);
nand U15899 (N_15899,N_12093,N_10771);
nand U15900 (N_15900,N_11616,N_13566);
nand U15901 (N_15901,N_11172,N_11373);
and U15902 (N_15902,N_11875,N_11039);
or U15903 (N_15903,N_13838,N_10627);
nand U15904 (N_15904,N_12098,N_14528);
or U15905 (N_15905,N_11533,N_11184);
nor U15906 (N_15906,N_12273,N_10715);
or U15907 (N_15907,N_12064,N_14325);
and U15908 (N_15908,N_13086,N_12282);
nand U15909 (N_15909,N_11631,N_12473);
nor U15910 (N_15910,N_11986,N_10201);
nand U15911 (N_15911,N_11445,N_13492);
nor U15912 (N_15912,N_10959,N_13665);
and U15913 (N_15913,N_12050,N_14729);
and U15914 (N_15914,N_11919,N_13429);
nor U15915 (N_15915,N_10246,N_14577);
xor U15916 (N_15916,N_13558,N_13958);
nand U15917 (N_15917,N_11618,N_13432);
or U15918 (N_15918,N_14494,N_13643);
nand U15919 (N_15919,N_10721,N_12963);
or U15920 (N_15920,N_10486,N_10807);
or U15921 (N_15921,N_12385,N_10284);
or U15922 (N_15922,N_10465,N_11068);
nand U15923 (N_15923,N_10688,N_13312);
and U15924 (N_15924,N_13382,N_10630);
or U15925 (N_15925,N_11451,N_14554);
nor U15926 (N_15926,N_10621,N_12682);
xor U15927 (N_15927,N_12109,N_10854);
nand U15928 (N_15928,N_10666,N_11382);
nor U15929 (N_15929,N_14251,N_12113);
and U15930 (N_15930,N_11795,N_14362);
nor U15931 (N_15931,N_12319,N_11571);
or U15932 (N_15932,N_12919,N_14735);
or U15933 (N_15933,N_13703,N_12977);
and U15934 (N_15934,N_12749,N_13793);
or U15935 (N_15935,N_10514,N_13729);
nor U15936 (N_15936,N_12215,N_11282);
or U15937 (N_15937,N_13375,N_13536);
or U15938 (N_15938,N_11666,N_10725);
and U15939 (N_15939,N_11183,N_13316);
and U15940 (N_15940,N_10453,N_11089);
nor U15941 (N_15941,N_14788,N_10366);
and U15942 (N_15942,N_13934,N_14047);
or U15943 (N_15943,N_10185,N_13068);
or U15944 (N_15944,N_10177,N_13638);
or U15945 (N_15945,N_13946,N_13499);
or U15946 (N_15946,N_10454,N_14317);
xnor U15947 (N_15947,N_13280,N_12007);
nor U15948 (N_15948,N_10500,N_14083);
and U15949 (N_15949,N_14718,N_12929);
nand U15950 (N_15950,N_13923,N_13982);
nor U15951 (N_15951,N_13484,N_14364);
and U15952 (N_15952,N_13142,N_11436);
nor U15953 (N_15953,N_10002,N_14555);
and U15954 (N_15954,N_11504,N_11609);
nand U15955 (N_15955,N_13435,N_13715);
nand U15956 (N_15956,N_14428,N_11805);
and U15957 (N_15957,N_14757,N_13266);
and U15958 (N_15958,N_12606,N_10842);
and U15959 (N_15959,N_14526,N_11955);
and U15960 (N_15960,N_12199,N_14852);
xnor U15961 (N_15961,N_14483,N_10378);
nor U15962 (N_15962,N_10689,N_13758);
nand U15963 (N_15963,N_12852,N_14918);
nand U15964 (N_15964,N_11210,N_14103);
xnor U15965 (N_15965,N_12709,N_10288);
and U15966 (N_15966,N_14262,N_12326);
or U15967 (N_15967,N_10195,N_11638);
nand U15968 (N_15968,N_12906,N_10186);
nand U15969 (N_15969,N_11096,N_12104);
nand U15970 (N_15970,N_10840,N_11667);
and U15971 (N_15971,N_11874,N_10490);
or U15972 (N_15972,N_13967,N_13070);
nor U15973 (N_15973,N_12805,N_13155);
and U15974 (N_15974,N_11407,N_10770);
and U15975 (N_15975,N_12493,N_11113);
xnor U15976 (N_15976,N_10165,N_14813);
and U15977 (N_15977,N_11607,N_11772);
or U15978 (N_15978,N_14803,N_10968);
and U15979 (N_15979,N_14449,N_11896);
and U15980 (N_15980,N_10924,N_14733);
nand U15981 (N_15981,N_11275,N_13501);
or U15982 (N_15982,N_10282,N_13804);
or U15983 (N_15983,N_12223,N_12648);
nor U15984 (N_15984,N_13692,N_13455);
nor U15985 (N_15985,N_13023,N_13810);
nor U15986 (N_15986,N_12898,N_12393);
nand U15987 (N_15987,N_11975,N_10143);
and U15988 (N_15988,N_12001,N_14656);
and U15989 (N_15989,N_13549,N_14172);
nand U15990 (N_15990,N_13999,N_12626);
or U15991 (N_15991,N_14446,N_10655);
or U15992 (N_15992,N_10023,N_11648);
and U15993 (N_15993,N_13705,N_10492);
or U15994 (N_15994,N_11810,N_13763);
or U15995 (N_15995,N_12666,N_14213);
nor U15996 (N_15996,N_13115,N_11690);
or U15997 (N_15997,N_11683,N_14214);
nand U15998 (N_15998,N_13936,N_11580);
nand U15999 (N_15999,N_11263,N_10985);
nand U16000 (N_16000,N_12417,N_13773);
xnor U16001 (N_16001,N_10727,N_10283);
nand U16002 (N_16002,N_13120,N_12760);
or U16003 (N_16003,N_14902,N_14872);
or U16004 (N_16004,N_13396,N_11165);
and U16005 (N_16005,N_10270,N_13890);
or U16006 (N_16006,N_14772,N_10995);
and U16007 (N_16007,N_12861,N_14242);
nor U16008 (N_16008,N_10692,N_13568);
or U16009 (N_16009,N_13861,N_11155);
nand U16010 (N_16010,N_14186,N_13574);
or U16011 (N_16011,N_12637,N_14095);
xor U16012 (N_16012,N_10224,N_14438);
or U16013 (N_16013,N_14942,N_14891);
or U16014 (N_16014,N_12669,N_11731);
nand U16015 (N_16015,N_10571,N_11947);
nor U16016 (N_16016,N_14190,N_13361);
xnor U16017 (N_16017,N_10425,N_13698);
and U16018 (N_16018,N_14843,N_10976);
xnor U16019 (N_16019,N_11158,N_11078);
nor U16020 (N_16020,N_13177,N_10474);
nor U16021 (N_16021,N_11143,N_11579);
nand U16022 (N_16022,N_12832,N_12692);
or U16023 (N_16023,N_13992,N_14627);
or U16024 (N_16024,N_10323,N_10011);
nand U16025 (N_16025,N_12317,N_10982);
or U16026 (N_16026,N_13195,N_13971);
nand U16027 (N_16027,N_14522,N_13198);
or U16028 (N_16028,N_12583,N_10358);
and U16029 (N_16029,N_12937,N_11306);
and U16030 (N_16030,N_11243,N_13331);
nand U16031 (N_16031,N_14259,N_11438);
nor U16032 (N_16032,N_12008,N_12654);
or U16033 (N_16033,N_12107,N_10544);
or U16034 (N_16034,N_13143,N_11557);
nand U16035 (N_16035,N_12694,N_12989);
nand U16036 (N_16036,N_10748,N_12118);
nand U16037 (N_16037,N_12243,N_10191);
nand U16038 (N_16038,N_10228,N_12149);
nand U16039 (N_16039,N_10009,N_13324);
and U16040 (N_16040,N_11500,N_12724);
nand U16041 (N_16041,N_11699,N_13117);
or U16042 (N_16042,N_13815,N_14151);
xnor U16043 (N_16043,N_11899,N_10192);
nor U16044 (N_16044,N_12851,N_11088);
and U16045 (N_16045,N_13641,N_10701);
nand U16046 (N_16046,N_13562,N_11847);
nor U16047 (N_16047,N_12585,N_12269);
nor U16048 (N_16048,N_13444,N_12095);
and U16049 (N_16049,N_12272,N_10348);
nor U16050 (N_16050,N_12741,N_10814);
and U16051 (N_16051,N_11139,N_12301);
and U16052 (N_16052,N_13976,N_13912);
or U16053 (N_16053,N_14283,N_12996);
or U16054 (N_16054,N_13158,N_10210);
nor U16055 (N_16055,N_13699,N_14859);
and U16056 (N_16056,N_12333,N_13090);
nand U16057 (N_16057,N_10180,N_12035);
or U16058 (N_16058,N_13965,N_11658);
and U16059 (N_16059,N_14663,N_13972);
nor U16060 (N_16060,N_14507,N_14297);
nand U16061 (N_16061,N_11101,N_14666);
and U16062 (N_16062,N_13166,N_11783);
xor U16063 (N_16063,N_13579,N_12238);
xor U16064 (N_16064,N_13299,N_13766);
nor U16065 (N_16065,N_12688,N_14272);
or U16066 (N_16066,N_13092,N_12278);
nand U16067 (N_16067,N_13769,N_10830);
nand U16068 (N_16068,N_14018,N_11393);
xnor U16069 (N_16069,N_12764,N_11817);
nand U16070 (N_16070,N_10573,N_12491);
nand U16071 (N_16071,N_11206,N_10838);
or U16072 (N_16072,N_12043,N_14244);
and U16073 (N_16073,N_12856,N_12783);
nor U16074 (N_16074,N_11410,N_12770);
nand U16075 (N_16075,N_11512,N_14378);
or U16076 (N_16076,N_11496,N_12343);
nand U16077 (N_16077,N_14894,N_10585);
or U16078 (N_16078,N_11880,N_11812);
nor U16079 (N_16079,N_12434,N_11239);
nand U16080 (N_16080,N_11901,N_13612);
or U16081 (N_16081,N_10363,N_14239);
or U16082 (N_16082,N_13391,N_11796);
nand U16083 (N_16083,N_10189,N_14724);
nor U16084 (N_16084,N_14545,N_14024);
and U16085 (N_16085,N_12103,N_10949);
nand U16086 (N_16086,N_10164,N_13448);
or U16087 (N_16087,N_11615,N_13952);
or U16088 (N_16088,N_12476,N_10668);
or U16089 (N_16089,N_10437,N_13344);
nand U16090 (N_16090,N_14969,N_13274);
xnor U16091 (N_16091,N_10810,N_11092);
or U16092 (N_16092,N_13868,N_10693);
nor U16093 (N_16093,N_11725,N_11923);
nor U16094 (N_16094,N_10160,N_13253);
xor U16095 (N_16095,N_14687,N_14049);
nor U16096 (N_16096,N_11585,N_10557);
and U16097 (N_16097,N_14122,N_12479);
nand U16098 (N_16098,N_10612,N_13434);
xnor U16099 (N_16099,N_10158,N_13425);
and U16100 (N_16100,N_14332,N_14042);
nor U16101 (N_16101,N_13397,N_11466);
or U16102 (N_16102,N_11224,N_14299);
xor U16103 (N_16103,N_12580,N_12945);
xor U16104 (N_16104,N_14826,N_14140);
and U16105 (N_16105,N_14289,N_12206);
and U16106 (N_16106,N_14366,N_14849);
nor U16107 (N_16107,N_14625,N_14007);
nand U16108 (N_16108,N_13012,N_12623);
or U16109 (N_16109,N_10444,N_12152);
xor U16110 (N_16110,N_14414,N_12056);
nand U16111 (N_16111,N_11130,N_14462);
or U16112 (N_16112,N_13376,N_13261);
and U16113 (N_16113,N_14943,N_14206);
and U16114 (N_16114,N_11211,N_10030);
or U16115 (N_16115,N_12275,N_11750);
and U16116 (N_16116,N_11914,N_10857);
and U16117 (N_16117,N_14898,N_10240);
or U16118 (N_16118,N_11726,N_11723);
or U16119 (N_16119,N_11087,N_10894);
xnor U16120 (N_16120,N_12812,N_11400);
and U16121 (N_16121,N_14252,N_14207);
and U16122 (N_16122,N_12519,N_11351);
nor U16123 (N_16123,N_11122,N_10258);
nand U16124 (N_16124,N_10473,N_10888);
nand U16125 (N_16125,N_11230,N_11456);
nor U16126 (N_16126,N_14955,N_13323);
nand U16127 (N_16127,N_10222,N_13822);
xor U16128 (N_16128,N_11120,N_12310);
nor U16129 (N_16129,N_10082,N_13330);
xnor U16130 (N_16130,N_10216,N_11179);
and U16131 (N_16131,N_13557,N_12069);
or U16132 (N_16132,N_14889,N_12252);
nand U16133 (N_16133,N_11569,N_10311);
nand U16134 (N_16134,N_10589,N_13706);
nor U16135 (N_16135,N_14919,N_10852);
nand U16136 (N_16136,N_14546,N_11933);
or U16137 (N_16137,N_13353,N_13230);
or U16138 (N_16138,N_10426,N_12324);
nand U16139 (N_16139,N_11416,N_14785);
xnor U16140 (N_16140,N_12183,N_14619);
and U16141 (N_16141,N_10381,N_10648);
or U16142 (N_16142,N_12344,N_13204);
and U16143 (N_16143,N_14707,N_11175);
xnor U16144 (N_16144,N_12055,N_12957);
nor U16145 (N_16145,N_10333,N_13660);
or U16146 (N_16146,N_10792,N_11147);
or U16147 (N_16147,N_12367,N_14096);
and U16148 (N_16148,N_12948,N_11298);
nor U16149 (N_16149,N_11719,N_14354);
nand U16150 (N_16150,N_10273,N_10475);
xnor U16151 (N_16151,N_13916,N_10783);
and U16152 (N_16152,N_11940,N_12349);
or U16153 (N_16153,N_12218,N_11855);
and U16154 (N_16154,N_10212,N_10110);
nand U16155 (N_16155,N_14288,N_10308);
or U16156 (N_16156,N_14314,N_14712);
nor U16157 (N_16157,N_11584,N_12135);
or U16158 (N_16158,N_14549,N_12599);
nand U16159 (N_16159,N_13533,N_12190);
nand U16160 (N_16160,N_14307,N_11244);
or U16161 (N_16161,N_12472,N_13602);
and U16162 (N_16162,N_12165,N_14997);
and U16163 (N_16163,N_14178,N_14787);
xor U16164 (N_16164,N_11209,N_12378);
and U16165 (N_16165,N_12800,N_11323);
and U16166 (N_16166,N_10809,N_10394);
nor U16167 (N_16167,N_13806,N_11386);
or U16168 (N_16168,N_14584,N_14091);
nand U16169 (N_16169,N_13426,N_14547);
or U16170 (N_16170,N_12761,N_12171);
nor U16171 (N_16171,N_13427,N_11514);
or U16172 (N_16172,N_13366,N_14639);
nor U16173 (N_16173,N_12407,N_12928);
nor U16174 (N_16174,N_12216,N_11900);
and U16175 (N_16175,N_13211,N_11477);
nor U16176 (N_16176,N_11186,N_14896);
nand U16177 (N_16177,N_12589,N_12329);
nand U16178 (N_16178,N_12431,N_10449);
or U16179 (N_16179,N_11452,N_13684);
nand U16180 (N_16180,N_11753,N_10679);
xor U16181 (N_16181,N_10219,N_10076);
nand U16182 (N_16182,N_14065,N_10489);
nand U16183 (N_16183,N_13486,N_14347);
nand U16184 (N_16184,N_10950,N_10277);
and U16185 (N_16185,N_13385,N_11737);
or U16186 (N_16186,N_10445,N_10372);
and U16187 (N_16187,N_13877,N_13908);
nor U16188 (N_16188,N_12582,N_12504);
nand U16189 (N_16189,N_11350,N_13121);
xor U16190 (N_16190,N_14187,N_14469);
nand U16191 (N_16191,N_12425,N_10653);
and U16192 (N_16192,N_10607,N_10616);
xor U16193 (N_16193,N_10550,N_11843);
nand U16194 (N_16194,N_13677,N_13051);
nor U16195 (N_16195,N_13702,N_12410);
nor U16196 (N_16196,N_10766,N_14352);
and U16197 (N_16197,N_11270,N_13313);
or U16198 (N_16198,N_10320,N_13251);
nor U16199 (N_16199,N_10660,N_10714);
or U16200 (N_16200,N_10879,N_12010);
nand U16201 (N_16201,N_13652,N_14127);
nand U16202 (N_16202,N_10343,N_10232);
and U16203 (N_16203,N_12663,N_13712);
or U16204 (N_16204,N_10802,N_13988);
or U16205 (N_16205,N_14696,N_14422);
and U16206 (N_16206,N_11574,N_11814);
and U16207 (N_16207,N_12707,N_14033);
nand U16208 (N_16208,N_13134,N_11794);
or U16209 (N_16209,N_10067,N_12931);
nand U16210 (N_16210,N_14802,N_14302);
xor U16211 (N_16211,N_13242,N_11945);
and U16212 (N_16212,N_10117,N_13026);
or U16213 (N_16213,N_10661,N_13546);
nand U16214 (N_16214,N_12496,N_12481);
xor U16215 (N_16215,N_12773,N_14801);
nor U16216 (N_16216,N_14335,N_11289);
nand U16217 (N_16217,N_12793,N_11305);
nor U16218 (N_16218,N_10559,N_14879);
nor U16219 (N_16219,N_10929,N_12513);
xnor U16220 (N_16220,N_10459,N_14472);
xor U16221 (N_16221,N_13100,N_12350);
nor U16222 (N_16222,N_14085,N_12634);
or U16223 (N_16223,N_13303,N_13275);
nor U16224 (N_16224,N_10287,N_13103);
nand U16225 (N_16225,N_12167,N_10608);
and U16226 (N_16226,N_14175,N_13778);
xor U16227 (N_16227,N_13234,N_10507);
or U16228 (N_16228,N_11717,N_14408);
xor U16229 (N_16229,N_14704,N_13918);
nor U16230 (N_16230,N_11141,N_14224);
and U16231 (N_16231,N_12406,N_10386);
xnor U16232 (N_16232,N_13095,N_11354);
nand U16233 (N_16233,N_14780,N_10089);
nor U16234 (N_16234,N_10563,N_11864);
nand U16235 (N_16235,N_13395,N_10128);
and U16236 (N_16236,N_13148,N_13081);
or U16237 (N_16237,N_10085,N_10325);
or U16238 (N_16238,N_14020,N_14043);
nor U16239 (N_16239,N_10145,N_11356);
or U16240 (N_16240,N_11433,N_10919);
or U16241 (N_16241,N_14039,N_14563);
nand U16242 (N_16242,N_10436,N_12677);
and U16243 (N_16243,N_10037,N_13604);
nand U16244 (N_16244,N_10788,N_14596);
or U16245 (N_16245,N_12803,N_12146);
nand U16246 (N_16246,N_10704,N_10365);
or U16247 (N_16247,N_14792,N_11469);
nand U16248 (N_16248,N_13847,N_14403);
and U16249 (N_16249,N_11963,N_10319);
or U16250 (N_16250,N_14058,N_14657);
nand U16251 (N_16251,N_11575,N_12231);
nand U16252 (N_16252,N_11711,N_13575);
and U16253 (N_16253,N_14089,N_11757);
and U16254 (N_16254,N_13741,N_12038);
and U16255 (N_16255,N_10928,N_11727);
nand U16256 (N_16256,N_12769,N_10599);
nand U16257 (N_16257,N_13139,N_11990);
nor U16258 (N_16258,N_14479,N_10104);
or U16259 (N_16259,N_12733,N_10865);
nor U16260 (N_16260,N_10622,N_12375);
xnor U16261 (N_16261,N_10460,N_12457);
or U16262 (N_16262,N_12075,N_10438);
and U16263 (N_16263,N_12639,N_10081);
nor U16264 (N_16264,N_10135,N_11786);
xnor U16265 (N_16265,N_10065,N_12369);
nand U16266 (N_16266,N_12237,N_14391);
or U16267 (N_16267,N_12600,N_11007);
nor U16268 (N_16268,N_10355,N_13069);
or U16269 (N_16269,N_11475,N_11097);
and U16270 (N_16270,N_11600,N_12934);
nand U16271 (N_16271,N_13305,N_13685);
nand U16272 (N_16272,N_12277,N_12219);
and U16273 (N_16273,N_14261,N_11582);
nor U16274 (N_16274,N_14267,N_14848);
or U16275 (N_16275,N_13767,N_14308);
or U16276 (N_16276,N_14550,N_10645);
xor U16277 (N_16277,N_12892,N_12954);
nor U16278 (N_16278,N_11076,N_12320);
nor U16279 (N_16279,N_13627,N_13149);
nor U16280 (N_16280,N_10934,N_12392);
and U16281 (N_16281,N_14147,N_13355);
nor U16282 (N_16282,N_11050,N_13482);
nor U16283 (N_16283,N_14443,N_11744);
nor U16284 (N_16284,N_14255,N_14909);
and U16285 (N_16285,N_12614,N_14059);
nand U16286 (N_16286,N_12742,N_11046);
xnor U16287 (N_16287,N_14326,N_10256);
or U16288 (N_16288,N_10470,N_13875);
xor U16289 (N_16289,N_14967,N_12705);
nand U16290 (N_16290,N_11053,N_10553);
and U16291 (N_16291,N_13887,N_11014);
and U16292 (N_16292,N_10789,N_14916);
nor U16293 (N_16293,N_14037,N_14569);
or U16294 (N_16294,N_13671,N_13565);
and U16295 (N_16295,N_13668,N_11994);
nor U16296 (N_16296,N_10828,N_10897);
and U16297 (N_16297,N_12884,N_13363);
nor U16298 (N_16298,N_14949,N_14310);
nor U16299 (N_16299,N_14643,N_14123);
or U16300 (N_16300,N_11189,N_12019);
xor U16301 (N_16301,N_13597,N_11482);
or U16302 (N_16302,N_11075,N_12298);
nand U16303 (N_16303,N_11854,N_13203);
nor U16304 (N_16304,N_13629,N_11954);
xnor U16305 (N_16305,N_11316,N_13571);
xnor U16306 (N_16306,N_12187,N_14868);
or U16307 (N_16307,N_13797,N_10427);
and U16308 (N_16308,N_10057,N_11103);
nand U16309 (N_16309,N_11010,N_12134);
nand U16310 (N_16310,N_11862,N_11749);
nand U16311 (N_16311,N_13296,N_11559);
nand U16312 (N_16312,N_10760,N_13213);
and U16313 (N_16313,N_12917,N_12220);
and U16314 (N_16314,N_14273,N_12529);
and U16315 (N_16315,N_14460,N_13440);
nand U16316 (N_16316,N_14233,N_14753);
or U16317 (N_16317,N_13169,N_12983);
or U16318 (N_16318,N_11702,N_14387);
and U16319 (N_16319,N_14134,N_14519);
or U16320 (N_16320,N_12387,N_14989);
or U16321 (N_16321,N_10041,N_13052);
nand U16322 (N_16322,N_11850,N_11226);
xor U16323 (N_16323,N_10488,N_12300);
or U16324 (N_16324,N_10583,N_12111);
xnor U16325 (N_16325,N_14173,N_12925);
and U16326 (N_16326,N_13870,N_14097);
nand U16327 (N_16327,N_10620,N_10389);
and U16328 (N_16328,N_13060,N_14221);
nor U16329 (N_16329,N_10482,N_13879);
nand U16330 (N_16330,N_14142,N_10617);
or U16331 (N_16331,N_12345,N_14260);
or U16332 (N_16332,N_12117,N_10718);
nor U16333 (N_16333,N_12604,N_13587);
nand U16334 (N_16334,N_13635,N_10531);
and U16335 (N_16335,N_13502,N_14738);
nor U16336 (N_16336,N_13465,N_11672);
and U16337 (N_16337,N_13580,N_10152);
or U16338 (N_16338,N_10947,N_11414);
and U16339 (N_16339,N_11832,N_10494);
xor U16340 (N_16340,N_11827,N_13490);
and U16341 (N_16341,N_11858,N_10083);
nand U16342 (N_16342,N_12451,N_10908);
nand U16343 (N_16343,N_12627,N_10197);
nor U16344 (N_16344,N_11352,N_11059);
nand U16345 (N_16345,N_12511,N_11926);
nand U16346 (N_16346,N_14583,N_10820);
nor U16347 (N_16347,N_10738,N_11803);
and U16348 (N_16348,N_12163,N_11473);
nand U16349 (N_16349,N_10853,N_13963);
and U16350 (N_16350,N_12508,N_10686);
and U16351 (N_16351,N_13795,N_10984);
and U16352 (N_16352,N_11286,N_11168);
or U16353 (N_16353,N_10456,N_14495);
or U16354 (N_16354,N_10605,N_10260);
and U16355 (N_16355,N_11730,N_13463);
nor U16356 (N_16356,N_10759,N_14331);
xnor U16357 (N_16357,N_14197,N_12401);
nand U16358 (N_16358,N_14947,N_14066);
nand U16359 (N_16359,N_13088,N_13214);
xnor U16360 (N_16360,N_14912,N_12942);
or U16361 (N_16361,N_13681,N_13764);
or U16362 (N_16362,N_14210,N_14502);
and U16363 (N_16363,N_14105,N_11142);
and U16364 (N_16364,N_14489,N_10570);
or U16365 (N_16365,N_14381,N_12044);
nor U16366 (N_16366,N_11145,N_11989);
and U16367 (N_16367,N_14744,N_12335);
and U16368 (N_16368,N_11266,N_12978);
or U16369 (N_16369,N_13676,N_13541);
nand U16370 (N_16370,N_10972,N_13904);
nand U16371 (N_16371,N_13016,N_12263);
and U16372 (N_16372,N_10250,N_14810);
and U16373 (N_16373,N_14032,N_11196);
nor U16374 (N_16374,N_13067,N_12091);
and U16375 (N_16375,N_11883,N_13423);
and U16376 (N_16376,N_10736,N_13747);
and U16377 (N_16377,N_11499,N_12660);
xnor U16378 (N_16378,N_14385,N_14530);
or U16379 (N_16379,N_14108,N_13445);
and U16380 (N_16380,N_14850,N_14893);
nand U16381 (N_16381,N_10667,N_12875);
or U16382 (N_16382,N_10088,N_13163);
nor U16383 (N_16383,N_11133,N_11094);
or U16384 (N_16384,N_11934,N_10004);
nor U16385 (N_16385,N_13968,N_13891);
xor U16386 (N_16386,N_12857,N_14762);
or U16387 (N_16387,N_12067,N_10018);
nor U16388 (N_16388,N_10252,N_11718);
and U16389 (N_16389,N_13087,N_11303);
nand U16390 (N_16390,N_13379,N_14717);
or U16391 (N_16391,N_13813,N_10797);
or U16392 (N_16392,N_12969,N_11331);
nand U16393 (N_16393,N_14041,N_14237);
nor U16394 (N_16394,N_14488,N_14112);
nand U16395 (N_16395,N_11654,N_12458);
nor U16396 (N_16396,N_11481,N_13909);
nand U16397 (N_16397,N_11338,N_12422);
or U16398 (N_16398,N_14447,N_13724);
nor U16399 (N_16399,N_13513,N_12169);
nor U16400 (N_16400,N_12334,N_12772);
and U16401 (N_16401,N_12029,N_12145);
and U16402 (N_16402,N_10726,N_10988);
nand U16403 (N_16403,N_13852,N_11694);
and U16404 (N_16404,N_13948,N_12526);
and U16405 (N_16405,N_14790,N_10541);
nor U16406 (N_16406,N_13325,N_10872);
and U16407 (N_16407,N_13315,N_10044);
xor U16408 (N_16408,N_10787,N_13352);
and U16409 (N_16409,N_11430,N_11724);
nor U16410 (N_16410,N_11784,N_13239);
and U16411 (N_16411,N_12636,N_12036);
nor U16412 (N_16412,N_13182,N_14434);
and U16413 (N_16413,N_14218,N_12653);
or U16414 (N_16414,N_13788,N_13737);
nor U16415 (N_16415,N_10864,N_10923);
nor U16416 (N_16416,N_10238,N_12266);
and U16417 (N_16417,N_14264,N_11098);
nand U16418 (N_16418,N_14219,N_14156);
or U16419 (N_16419,N_12916,N_14806);
or U16420 (N_16420,N_11247,N_12304);
and U16421 (N_16421,N_13983,N_10746);
and U16422 (N_16422,N_12775,N_10855);
nor U16423 (N_16423,N_10730,N_11446);
nand U16424 (N_16424,N_11187,N_13817);
nor U16425 (N_16425,N_11698,N_10217);
nor U16426 (N_16426,N_13128,N_14668);
and U16427 (N_16427,N_14779,N_14015);
or U16428 (N_16428,N_13944,N_11972);
xnor U16429 (N_16429,N_14161,N_13760);
nand U16430 (N_16430,N_10918,N_14411);
nor U16431 (N_16431,N_14030,N_13530);
and U16432 (N_16432,N_10502,N_13337);
or U16433 (N_16433,N_10837,N_12728);
nand U16434 (N_16434,N_10941,N_10781);
xor U16435 (N_16435,N_10535,N_13453);
nor U16436 (N_16436,N_13057,N_12933);
nand U16437 (N_16437,N_14775,N_14804);
xnor U16438 (N_16438,N_11484,N_12346);
nor U16439 (N_16439,N_12368,N_12870);
nand U16440 (N_16440,N_10905,N_10915);
and U16441 (N_16441,N_13669,N_13288);
or U16442 (N_16442,N_11815,N_14291);
and U16443 (N_16443,N_11077,N_11935);
and U16444 (N_16444,N_10353,N_13649);
nor U16445 (N_16445,N_11173,N_13321);
nand U16446 (N_16446,N_12520,N_11697);
xor U16447 (N_16447,N_13903,N_14715);
or U16448 (N_16448,N_11790,N_14782);
nor U16449 (N_16449,N_10706,N_12615);
or U16450 (N_16450,N_13505,N_14728);
and U16451 (N_16451,N_12489,N_14832);
and U16452 (N_16452,N_10640,N_13254);
nand U16453 (N_16453,N_12794,N_12041);
and U16454 (N_16454,N_14137,N_10251);
or U16455 (N_16455,N_11665,N_12890);
and U16456 (N_16456,N_10635,N_10519);
or U16457 (N_16457,N_10745,N_14405);
and U16458 (N_16458,N_12321,N_14476);
and U16459 (N_16459,N_10187,N_11853);
nand U16460 (N_16460,N_14270,N_12115);
nand U16461 (N_16461,N_14511,N_13116);
nor U16462 (N_16462,N_10900,N_13791);
and U16463 (N_16463,N_12390,N_10722);
nor U16464 (N_16464,N_14524,N_12283);
nor U16465 (N_16465,N_14934,N_11770);
or U16466 (N_16466,N_14743,N_12817);
nor U16467 (N_16467,N_11546,N_14892);
and U16468 (N_16468,N_13842,N_12592);
nor U16469 (N_16469,N_14425,N_10137);
or U16470 (N_16470,N_12547,N_10188);
xnor U16471 (N_16471,N_10040,N_14243);
or U16472 (N_16472,N_14604,N_13880);
and U16473 (N_16473,N_12421,N_12721);
or U16474 (N_16474,N_14120,N_12784);
or U16475 (N_16475,N_12701,N_11063);
and U16476 (N_16476,N_12424,N_11008);
or U16477 (N_16477,N_11884,N_12577);
and U16478 (N_16478,N_12943,N_13850);
and U16479 (N_16479,N_14171,N_10587);
nand U16480 (N_16480,N_10633,N_10257);
xnor U16481 (N_16481,N_13381,N_14410);
and U16482 (N_16482,N_13645,N_14349);
nand U16483 (N_16483,N_12581,N_14939);
and U16484 (N_16484,N_13030,N_11889);
or U16485 (N_16485,N_14078,N_14199);
xor U16486 (N_16486,N_13545,N_13902);
or U16487 (N_16487,N_14901,N_13544);
nor U16488 (N_16488,N_10114,N_13774);
nor U16489 (N_16489,N_12541,N_14936);
nand U16490 (N_16490,N_13260,N_13524);
and U16491 (N_16491,N_14871,N_14436);
nand U16492 (N_16492,N_11942,N_10674);
nand U16493 (N_16493,N_12656,N_11383);
and U16494 (N_16494,N_14265,N_10337);
and U16495 (N_16495,N_12575,N_11056);
and U16496 (N_16496,N_11440,N_12488);
and U16497 (N_16497,N_13220,N_12992);
nor U16498 (N_16498,N_13591,N_11128);
nand U16499 (N_16499,N_11397,N_12888);
nand U16500 (N_16500,N_11381,N_10326);
nand U16501 (N_16501,N_14452,N_12148);
and U16502 (N_16502,N_10548,N_14045);
xnor U16503 (N_16503,N_10174,N_14708);
or U16504 (N_16504,N_13014,N_14285);
nor U16505 (N_16505,N_11839,N_11977);
xor U16506 (N_16506,N_14184,N_10675);
nor U16507 (N_16507,N_11660,N_13227);
nand U16508 (N_16508,N_12279,N_12196);
or U16509 (N_16509,N_14819,N_14204);
and U16510 (N_16510,N_12679,N_12587);
or U16511 (N_16511,N_10289,N_11479);
xnor U16512 (N_16512,N_11872,N_13951);
nand U16513 (N_16513,N_13631,N_14922);
nand U16514 (N_16514,N_11695,N_13464);
nor U16515 (N_16515,N_10784,N_11052);
and U16516 (N_16516,N_11605,N_11886);
or U16517 (N_16517,N_12383,N_11030);
nor U16518 (N_16518,N_12535,N_12726);
nor U16519 (N_16519,N_14975,N_12991);
and U16520 (N_16520,N_12166,N_12534);
and U16521 (N_16521,N_14515,N_11678);
and U16522 (N_16522,N_10659,N_12872);
and U16523 (N_16523,N_13526,N_14562);
and U16524 (N_16524,N_14705,N_10861);
and U16525 (N_16525,N_11781,N_14559);
and U16526 (N_16526,N_12232,N_12838);
nand U16527 (N_16527,N_13089,N_10954);
nand U16528 (N_16528,N_10483,N_12993);
or U16529 (N_16529,N_14271,N_10651);
or U16530 (N_16530,N_10610,N_11214);
nand U16531 (N_16531,N_14338,N_13553);
nor U16532 (N_16532,N_14003,N_10833);
nor U16533 (N_16533,N_12647,N_14626);
nor U16534 (N_16534,N_12893,N_13866);
or U16535 (N_16535,N_13860,N_13456);
and U16536 (N_16536,N_12140,N_12136);
and U16537 (N_16537,N_12084,N_14970);
or U16538 (N_16538,N_11042,N_13718);
or U16539 (N_16539,N_14846,N_13666);
nand U16540 (N_16540,N_14121,N_12638);
nor U16541 (N_16541,N_12120,N_11036);
nor U16542 (N_16542,N_13700,N_14176);
and U16543 (N_16543,N_10647,N_12287);
xnor U16544 (N_16544,N_12834,N_11897);
xnor U16545 (N_16545,N_10408,N_11664);
nand U16546 (N_16546,N_12024,N_14671);
and U16547 (N_16547,N_10066,N_14068);
and U16548 (N_16548,N_13895,N_13957);
or U16549 (N_16549,N_12561,N_11868);
and U16550 (N_16550,N_12958,N_11392);
nand U16551 (N_16551,N_10367,N_13135);
and U16552 (N_16552,N_13933,N_11435);
xnor U16553 (N_16553,N_10204,N_11807);
and U16554 (N_16554,N_14404,N_13408);
nand U16555 (N_16555,N_11043,N_13190);
nor U16556 (N_16556,N_11797,N_12362);
and U16557 (N_16557,N_11563,N_13730);
or U16558 (N_16558,N_10419,N_12155);
and U16559 (N_16559,N_11651,N_14932);
nor U16560 (N_16560,N_14029,N_14920);
nor U16561 (N_16561,N_11181,N_11606);
nor U16562 (N_16562,N_13098,N_12828);
nand U16563 (N_16563,N_12083,N_10930);
or U16564 (N_16564,N_14764,N_12239);
and U16565 (N_16565,N_11371,N_12936);
nand U16566 (N_16566,N_10471,N_13301);
nand U16567 (N_16567,N_10278,N_14661);
xnor U16568 (N_16568,N_10467,N_13796);
or U16569 (N_16569,N_12824,N_11003);
or U16570 (N_16570,N_13921,N_10060);
nand U16571 (N_16571,N_11709,N_11105);
nor U16572 (N_16572,N_14229,N_14465);
and U16573 (N_16573,N_10793,N_13906);
nand U16574 (N_16574,N_11449,N_12869);
xnor U16575 (N_16575,N_10172,N_13639);
nor U16576 (N_16576,N_10035,N_10476);
nand U16577 (N_16577,N_12605,N_12514);
or U16578 (N_16578,N_13925,N_11458);
or U16579 (N_16579,N_13481,N_13424);
xor U16580 (N_16580,N_13633,N_11622);
nor U16581 (N_16581,N_11134,N_11464);
and U16582 (N_16582,N_11429,N_11952);
or U16583 (N_16583,N_14057,N_12938);
and U16584 (N_16584,N_14106,N_11448);
nand U16585 (N_16585,N_11362,N_13673);
nor U16586 (N_16586,N_14818,N_13621);
nor U16587 (N_16587,N_14736,N_11032);
nor U16588 (N_16588,N_12398,N_11842);
nand U16589 (N_16589,N_13193,N_13082);
or U16590 (N_16590,N_12170,N_13094);
nor U16591 (N_16591,N_10455,N_11777);
nor U16592 (N_16592,N_12822,N_11333);
or U16593 (N_16593,N_11054,N_12941);
nor U16594 (N_16594,N_14231,N_13258);
or U16595 (N_16595,N_14624,N_10938);
and U16596 (N_16596,N_11552,N_12427);
nand U16597 (N_16597,N_13042,N_10998);
nor U16598 (N_16598,N_10871,N_11425);
nor U16599 (N_16599,N_13717,N_13200);
nor U16600 (N_16600,N_14075,N_12351);
or U16601 (N_16601,N_12268,N_14988);
and U16602 (N_16602,N_12731,N_14617);
nor U16603 (N_16603,N_12291,N_14512);
nor U16604 (N_16604,N_12538,N_13050);
or U16605 (N_16605,N_13226,N_13279);
nand U16606 (N_16606,N_14235,N_12053);
xor U16607 (N_16607,N_12727,N_10215);
or U16608 (N_16608,N_13493,N_10582);
nand U16609 (N_16609,N_10075,N_14274);
or U16610 (N_16610,N_12717,N_12079);
nor U16611 (N_16611,N_11995,N_12123);
nor U16612 (N_16612,N_12128,N_12591);
nand U16613 (N_16613,N_10538,N_14721);
xnor U16614 (N_16614,N_11997,N_14740);
nand U16615 (N_16615,N_10375,N_14727);
xnor U16616 (N_16616,N_14513,N_12302);
or U16617 (N_16617,N_14312,N_13415);
nand U16618 (N_16618,N_11022,N_13390);
nand U16619 (N_16619,N_10028,N_12839);
nand U16620 (N_16620,N_10962,N_12459);
or U16621 (N_16621,N_14683,N_13219);
and U16622 (N_16622,N_12086,N_13147);
xnor U16623 (N_16623,N_14076,N_10713);
nand U16624 (N_16624,N_13732,N_14971);
and U16625 (N_16625,N_13678,N_11156);
or U16626 (N_16626,N_13202,N_12825);
nor U16627 (N_16627,N_10339,N_10382);
xnor U16628 (N_16628,N_11920,N_13442);
and U16629 (N_16629,N_11483,N_10927);
and U16630 (N_16630,N_11656,N_12192);
xnor U16631 (N_16631,N_13388,N_12074);
nand U16632 (N_16632,N_10072,N_13310);
nor U16633 (N_16633,N_13609,N_14999);
nand U16634 (N_16634,N_12423,N_10181);
nand U16635 (N_16635,N_14316,N_14523);
xor U16636 (N_16636,N_12285,N_10533);
nand U16637 (N_16637,N_13570,N_12361);
or U16638 (N_16638,N_13112,N_13362);
nor U16639 (N_16639,N_12475,N_11801);
and U16640 (N_16640,N_12804,N_14027);
nand U16641 (N_16641,N_11185,N_13756);
nor U16642 (N_16642,N_14456,N_10601);
nand U16643 (N_16643,N_14509,N_10155);
nand U16644 (N_16644,N_13451,N_14246);
nor U16645 (N_16645,N_10777,N_14799);
nand U16646 (N_16646,N_12796,N_13359);
nor U16647 (N_16647,N_13333,N_11742);
and U16648 (N_16648,N_14582,N_14084);
nor U16649 (N_16649,N_12097,N_13818);
nand U16650 (N_16650,N_11677,N_10134);
nor U16651 (N_16651,N_13995,N_14964);
or U16652 (N_16652,N_10087,N_10543);
and U16653 (N_16653,N_12450,N_10499);
or U16654 (N_16654,N_12506,N_13241);
nand U16655 (N_16655,N_13264,N_10229);
xor U16656 (N_16656,N_10346,N_13581);
nor U16657 (N_16657,N_11967,N_12402);
xor U16658 (N_16658,N_14644,N_11974);
and U16659 (N_16659,N_12789,N_11154);
and U16660 (N_16660,N_14240,N_11044);
nor U16661 (N_16661,N_14675,N_10914);
nand U16662 (N_16662,N_14139,N_13611);
nand U16663 (N_16663,N_11104,N_13648);
nand U16664 (N_16664,N_11119,N_13943);
nor U16665 (N_16665,N_13256,N_11457);
or U16666 (N_16666,N_14144,N_11058);
or U16667 (N_16667,N_10125,N_12305);
and U16668 (N_16668,N_14749,N_14823);
or U16669 (N_16669,N_12174,N_13839);
or U16670 (N_16670,N_12470,N_13859);
and U16671 (N_16671,N_10569,N_10880);
and U16672 (N_16672,N_12862,N_11693);
nor U16673 (N_16673,N_14248,N_11501);
nand U16674 (N_16674,N_11329,N_12785);
nor U16675 (N_16675,N_10463,N_14498);
nor U16676 (N_16676,N_12014,N_14356);
nor U16677 (N_16677,N_11859,N_10835);
or U16678 (N_16678,N_10015,N_13548);
xnor U16679 (N_16679,N_13561,N_11511);
nand U16680 (N_16680,N_11161,N_10401);
and U16681 (N_16681,N_11568,N_11892);
nor U16682 (N_16682,N_10317,N_10646);
xor U16683 (N_16683,N_14754,N_11728);
or U16684 (N_16684,N_14945,N_10241);
xor U16685 (N_16685,N_14150,N_11245);
or U16686 (N_16686,N_14179,N_14635);
and U16687 (N_16687,N_14102,N_12553);
and U16688 (N_16688,N_14192,N_11876);
nand U16689 (N_16689,N_11567,N_14126);
nor U16690 (N_16690,N_11592,N_13106);
nor U16691 (N_16691,N_14648,N_10536);
nand U16692 (N_16692,N_10624,N_10975);
or U16693 (N_16693,N_13232,N_12737);
xnor U16694 (N_16694,N_12295,N_11115);
nand U16695 (N_16695,N_14389,N_12818);
and U16696 (N_16696,N_14763,N_12537);
or U16697 (N_16697,N_10609,N_14665);
or U16698 (N_16698,N_10739,N_13500);
and U16699 (N_16699,N_11623,N_13577);
and U16700 (N_16700,N_11509,N_11349);
and U16701 (N_16701,N_14884,N_13949);
or U16702 (N_16702,N_13317,N_14236);
or U16703 (N_16703,N_10234,N_14119);
nand U16704 (N_16704,N_13304,N_13349);
nand U16705 (N_16705,N_12462,N_11302);
or U16706 (N_16706,N_12494,N_12110);
or U16707 (N_16707,N_13578,N_10670);
or U16708 (N_16708,N_12594,N_10876);
and U16709 (N_16709,N_10253,N_11064);
nand U16710 (N_16710,N_12121,N_11979);
or U16711 (N_16711,N_11319,N_13777);
nor U16712 (N_16712,N_13985,N_12699);
or U16713 (N_16713,N_10683,N_14372);
nand U16714 (N_16714,N_14327,N_13462);
nor U16715 (N_16715,N_12131,N_13174);
nor U16716 (N_16716,N_14602,N_14238);
nor U16717 (N_16717,N_12073,N_10658);
and U16718 (N_16718,N_12918,N_12661);
nor U16719 (N_16719,N_12641,N_13656);
and U16720 (N_16720,N_12235,N_11841);
nand U16721 (N_16721,N_10665,N_11907);
nor U16722 (N_16722,N_10765,N_10290);
nand U16723 (N_16723,N_14230,N_11732);
nor U16724 (N_16724,N_10825,N_14157);
nand U16725 (N_16725,N_14485,N_13238);
nand U16726 (N_16726,N_10547,N_12522);
and U16727 (N_16727,N_10017,N_12920);
nand U16728 (N_16728,N_12059,N_10302);
nor U16729 (N_16729,N_11639,N_10795);
or U16730 (N_16730,N_10639,N_13809);
and U16731 (N_16731,N_14525,N_11467);
nor U16732 (N_16732,N_10649,N_12554);
nand U16733 (N_16733,N_14313,N_13006);
and U16734 (N_16734,N_10580,N_13626);
nor U16735 (N_16735,N_12125,N_12031);
or U16736 (N_16736,N_13306,N_13215);
nor U16737 (N_16737,N_12177,N_14115);
or U16738 (N_16738,N_10443,N_14601);
nand U16739 (N_16739,N_11932,N_14957);
and U16740 (N_16740,N_12430,N_11084);
and U16741 (N_16741,N_11374,N_14390);
or U16742 (N_16742,N_14004,N_13691);
nand U16743 (N_16743,N_10171,N_11878);
and U16744 (N_16744,N_14022,N_11242);
and U16745 (N_16745,N_14544,N_12469);
or U16746 (N_16746,N_13849,N_13865);
xor U16747 (N_16747,N_14508,N_10883);
and U16748 (N_16748,N_11300,N_14423);
or U16749 (N_16749,N_10564,N_12542);
xor U16750 (N_16750,N_14905,N_10882);
xnor U16751 (N_16751,N_11829,N_13247);
nor U16752 (N_16752,N_12940,N_11983);
or U16753 (N_16753,N_10555,N_11040);
nand U16754 (N_16754,N_12900,N_12062);
nor U16755 (N_16755,N_11712,N_10268);
and U16756 (N_16756,N_14344,N_11696);
or U16757 (N_16757,N_13719,N_12046);
and U16758 (N_16758,N_13693,N_14722);
and U16759 (N_16759,N_14287,N_14216);
xnor U16760 (N_16760,N_11453,N_10000);
nor U16761 (N_16761,N_14860,N_11996);
or U16762 (N_16762,N_10750,N_10012);
nor U16763 (N_16763,N_12556,N_11363);
nand U16764 (N_16764,N_10961,N_13858);
nor U16765 (N_16765,N_13474,N_11150);
xnor U16766 (N_16766,N_14521,N_10867);
and U16767 (N_16767,N_11190,N_13127);
nand U16768 (N_16768,N_10530,N_13074);
xor U16769 (N_16769,N_11928,N_12308);
nand U16770 (N_16770,N_11904,N_11541);
nand U16771 (N_16771,N_11871,N_13035);
xor U16772 (N_16772,N_11315,N_10109);
and U16773 (N_16773,N_11905,N_14678);
nor U16774 (N_16774,N_10773,N_12905);
and U16775 (N_16775,N_13405,N_12501);
and U16776 (N_16776,N_14094,N_10407);
xnor U16777 (N_16777,N_12005,N_10046);
and U16778 (N_16778,N_14226,N_14676);
nand U16779 (N_16779,N_10912,N_10994);
nand U16780 (N_16780,N_10973,N_10735);
or U16781 (N_16781,N_12833,N_13616);
nand U16782 (N_16782,N_12640,N_14895);
and U16783 (N_16783,N_12664,N_11902);
nor U16784 (N_16784,N_14815,N_10892);
and U16785 (N_16785,N_14834,N_11581);
nor U16786 (N_16786,N_12018,N_11970);
nor U16787 (N_16787,N_10576,N_13674);
nand U16788 (N_16788,N_12730,N_11508);
or U16789 (N_16789,N_11408,N_13843);
or U16790 (N_16790,N_11207,N_10528);
and U16791 (N_16791,N_11916,N_11733);
nor U16792 (N_16792,N_14950,N_11292);
nor U16793 (N_16793,N_11930,N_10963);
and U16794 (N_16794,N_12028,N_12621);
or U16795 (N_16795,N_13295,N_11256);
and U16796 (N_16796,N_10286,N_13929);
or U16797 (N_16797,N_10860,N_10220);
nand U16798 (N_16798,N_14363,N_13517);
or U16799 (N_16799,N_10084,N_14480);
and U16800 (N_16800,N_10400,N_10539);
nor U16801 (N_16801,N_13504,N_11341);
nor U16802 (N_16802,N_11650,N_13307);
nand U16803 (N_16803,N_11213,N_12802);
nand U16804 (N_16804,N_11936,N_12337);
nor U16805 (N_16805,N_13625,N_12576);
xnor U16806 (N_16806,N_12510,N_13824);
and U16807 (N_16807,N_10965,N_10863);
or U16808 (N_16808,N_12923,N_14808);
or U16809 (N_16809,N_10826,N_12203);
and U16810 (N_16810,N_14706,N_13063);
or U16811 (N_16811,N_14825,N_12157);
nand U16812 (N_16812,N_14948,N_10208);
nor U16813 (N_16813,N_12672,N_14132);
and U16814 (N_16814,N_14682,N_11888);
nand U16815 (N_16815,N_13314,N_14098);
or U16816 (N_16816,N_10263,N_12868);
and U16817 (N_16817,N_10774,N_11067);
xor U16818 (N_16818,N_10662,N_11741);
or U16819 (N_16819,N_14136,N_14797);
or U16820 (N_16820,N_12652,N_10312);
or U16821 (N_16821,N_14750,N_14748);
nor U16822 (N_16822,N_12567,N_10875);
nor U16823 (N_16823,N_12867,N_10116);
or U16824 (N_16824,N_10327,N_11943);
xnor U16825 (N_16825,N_14542,N_11252);
and U16826 (N_16826,N_14215,N_10935);
nor U16827 (N_16827,N_14328,N_13283);
nor U16828 (N_16828,N_11999,N_12579);
and U16829 (N_16829,N_13819,N_13521);
or U16830 (N_16830,N_12138,N_14320);
and U16831 (N_16831,N_14021,N_14923);
nand U16832 (N_16832,N_14516,N_14830);
or U16833 (N_16833,N_11599,N_14269);
or U16834 (N_16834,N_11194,N_13078);
or U16835 (N_16835,N_13653,N_14036);
or U16836 (N_16836,N_14930,N_12753);
or U16837 (N_16837,N_14858,N_13584);
and U16838 (N_16838,N_10139,N_12009);
xor U16839 (N_16839,N_14990,N_14009);
or U16840 (N_16840,N_14844,N_14693);
and U16841 (N_16841,N_10966,N_12478);
nor U16842 (N_16842,N_14250,N_10303);
and U16843 (N_16843,N_10255,N_12185);
or U16844 (N_16844,N_10546,N_14702);
or U16845 (N_16845,N_13062,N_14324);
nand U16846 (N_16846,N_14406,N_10974);
and U16847 (N_16847,N_11250,N_14548);
and U16848 (N_16848,N_11531,N_11192);
and U16849 (N_16849,N_12290,N_13863);
or U16850 (N_16850,N_13046,N_12082);
nand U16851 (N_16851,N_10958,N_10717);
and U16852 (N_16852,N_13977,N_11342);
and U16853 (N_16853,N_12214,N_10832);
nand U16854 (N_16854,N_12384,N_13073);
or U16855 (N_16855,N_11011,N_11450);
nor U16856 (N_16856,N_11311,N_13369);
nand U16857 (N_16857,N_11516,N_14087);
nand U16858 (N_16858,N_12680,N_14355);
nor U16859 (N_16859,N_11913,N_14710);
or U16860 (N_16860,N_12096,N_10001);
and U16861 (N_16861,N_14824,N_13371);
nor U16862 (N_16862,N_11624,N_14878);
or U16863 (N_16863,N_11671,N_12474);
nand U16864 (N_16864,N_10696,N_11813);
or U16865 (N_16865,N_13436,N_12687);
nand U16866 (N_16866,N_13407,N_10808);
and U16867 (N_16867,N_13005,N_12757);
xor U16868 (N_16868,N_14016,N_12207);
and U16869 (N_16869,N_13066,N_10829);
nor U16870 (N_16870,N_14698,N_12703);
or U16871 (N_16871,N_13401,N_12710);
nand U16872 (N_16872,N_12611,N_14499);
nor U16873 (N_16873,N_14652,N_13497);
or U16874 (N_16874,N_11248,N_14535);
and U16875 (N_16875,N_14379,N_12557);
nor U16876 (N_16876,N_11710,N_13059);
and U16877 (N_16877,N_12960,N_12226);
nor U16878 (N_16878,N_14667,N_11296);
and U16879 (N_16879,N_14917,N_14300);
nand U16880 (N_16880,N_13782,N_13683);
nand U16881 (N_16881,N_12595,N_11840);
nor U16882 (N_16882,N_12521,N_14980);
or U16883 (N_16883,N_10946,N_13857);
nand U16884 (N_16884,N_13277,N_12380);
and U16885 (N_16885,N_12173,N_11267);
nor U16886 (N_16886,N_11706,N_14293);
and U16887 (N_16887,N_12483,N_14129);
or U16888 (N_16888,N_10079,N_12814);
nand U16889 (N_16889,N_12799,N_13928);
and U16890 (N_16890,N_13438,N_10818);
and U16891 (N_16891,N_13551,N_11013);
nand U16892 (N_16892,N_11893,N_13955);
xnor U16893 (N_16893,N_13888,N_12040);
nor U16894 (N_16894,N_10479,N_12649);
xor U16895 (N_16895,N_11264,N_10061);
nor U16896 (N_16896,N_10103,N_10932);
xnor U16897 (N_16897,N_14647,N_11365);
nand U16898 (N_16898,N_14125,N_12607);
nand U16899 (N_16899,N_11108,N_11689);
nor U16900 (N_16900,N_11361,N_14795);
and U16901 (N_16901,N_13151,N_12759);
or U16902 (N_16902,N_12711,N_10869);
nand U16903 (N_16903,N_12763,N_13614);
and U16904 (N_16904,N_12433,N_12990);
or U16905 (N_16905,N_12443,N_10743);
and U16906 (N_16906,N_12039,N_14040);
nor U16907 (N_16907,N_11034,N_10062);
or U16908 (N_16908,N_13172,N_10753);
xor U16909 (N_16909,N_10163,N_14082);
nor U16910 (N_16910,N_13446,N_14044);
nor U16911 (N_16911,N_13728,N_14445);
or U16912 (N_16912,N_12037,N_11332);
nor U16913 (N_16913,N_13150,N_10657);
nor U16914 (N_16914,N_11413,N_10310);
and U16915 (N_16915,N_12896,N_11978);
or U16916 (N_16916,N_11787,N_14606);
nor U16917 (N_16917,N_11082,N_11037);
and U16918 (N_16918,N_14180,N_14732);
and U16919 (N_16919,N_13340,N_10364);
or U16920 (N_16920,N_11287,N_12980);
and U16921 (N_16921,N_13740,N_11903);
nand U16922 (N_16922,N_11268,N_14851);
xor U16923 (N_16923,N_12208,N_12331);
and U16924 (N_16924,N_11687,N_14234);
xnor U16925 (N_16925,N_12254,N_10094);
or U16926 (N_16926,N_14833,N_14532);
or U16927 (N_16927,N_10782,N_12175);
and U16928 (N_16928,N_14796,N_10981);
and U16929 (N_16929,N_11074,N_12047);
or U16930 (N_16930,N_13917,N_11234);
xnor U16931 (N_16931,N_11276,N_13252);
nor U16932 (N_16932,N_10952,N_12684);
xnor U16933 (N_16933,N_14581,N_14475);
nor U16934 (N_16934,N_11956,N_11601);
nor U16935 (N_16935,N_13309,N_13998);
or U16936 (N_16936,N_13123,N_12217);
or U16937 (N_16937,N_14440,N_13532);
or U16938 (N_16938,N_11636,N_14778);
or U16939 (N_16939,N_10999,N_13688);
nand U16940 (N_16940,N_11281,N_10680);
nand U16941 (N_16941,N_10149,N_11517);
nor U16942 (N_16942,N_12063,N_13197);
or U16943 (N_16943,N_13547,N_10642);
nand U16944 (N_16944,N_10447,N_14580);
nand U16945 (N_16945,N_10798,N_11966);
xnor U16946 (N_16946,N_14124,N_10020);
nor U16947 (N_16947,N_11785,N_10862);
nand U16948 (N_16948,N_11045,N_10342);
and U16949 (N_16949,N_11406,N_10664);
or U16950 (N_16950,N_11957,N_13962);
or U16951 (N_16951,N_14701,N_13789);
nor U16952 (N_16952,N_10846,N_10631);
nor U16953 (N_16953,N_12953,N_10951);
xnor U16954 (N_16954,N_13787,N_12877);
nor U16955 (N_16955,N_10218,N_12137);
xor U16956 (N_16956,N_13101,N_13488);
nand U16957 (N_16957,N_14504,N_14182);
nand U16958 (N_16958,N_11112,N_14249);
or U16959 (N_16959,N_14228,N_11980);
nand U16960 (N_16960,N_10124,N_12755);
or U16961 (N_16961,N_14063,N_13622);
nand U16962 (N_16962,N_12987,N_12550);
and U16963 (N_16963,N_10775,N_12132);
or U16964 (N_16964,N_14135,N_13224);
xor U16965 (N_16965,N_14334,N_11597);
nor U16966 (N_16966,N_13041,N_14631);
nand U16967 (N_16967,N_10579,N_13038);
nor U16968 (N_16968,N_14305,N_13146);
and U16969 (N_16969,N_13409,N_13784);
nor U16970 (N_16970,N_12307,N_11086);
nor U16971 (N_16971,N_13332,N_10895);
nand U16972 (N_16972,N_13509,N_14481);
nor U16973 (N_16973,N_11515,N_10032);
nand U16974 (N_16974,N_11318,N_11774);
nor U16975 (N_16975,N_14348,N_11284);
xnor U16976 (N_16976,N_12932,N_13518);
or U16977 (N_16977,N_11127,N_13646);
and U16978 (N_16978,N_10322,N_10016);
xnor U16979 (N_16979,N_11395,N_12449);
xor U16980 (N_16980,N_14800,N_12720);
nand U16981 (N_16981,N_11402,N_12853);
nor U16982 (N_16982,N_13007,N_10508);
xor U16983 (N_16983,N_13342,N_10021);
nand U16984 (N_16984,N_12012,N_10038);
and U16985 (N_16985,N_10896,N_10369);
nand U16986 (N_16986,N_13478,N_14292);
nor U16987 (N_16987,N_13180,N_10446);
and U16988 (N_16988,N_11202,N_11431);
or U16989 (N_16989,N_11739,N_13687);
nor U16990 (N_16990,N_10178,N_11502);
nor U16991 (N_16991,N_10099,N_14090);
nor U16992 (N_16992,N_13104,N_13262);
and U16993 (N_16993,N_14741,N_12360);
xor U16994 (N_16994,N_13534,N_10551);
xnor U16995 (N_16995,N_10800,N_12657);
nor U16996 (N_16996,N_11566,N_11415);
nor U16997 (N_16997,N_14100,N_13076);
xnor U16998 (N_16998,N_11621,N_14162);
and U16999 (N_16999,N_11591,N_13790);
nand U17000 (N_17000,N_12452,N_13291);
xnor U17001 (N_17001,N_13733,N_11260);
nor U17002 (N_17002,N_10812,N_14689);
nor U17003 (N_17003,N_10159,N_10827);
nand U17004 (N_17004,N_13114,N_10280);
nor U17005 (N_17005,N_11969,N_12502);
and U17006 (N_17006,N_11385,N_14295);
or U17007 (N_17007,N_10168,N_14092);
and U17008 (N_17008,N_11336,N_10423);
or U17009 (N_17009,N_11604,N_10466);
or U17010 (N_17010,N_12947,N_13056);
and U17011 (N_17011,N_14587,N_14081);
or U17012 (N_17012,N_12736,N_12635);
and U17013 (N_17013,N_11138,N_11551);
and U17014 (N_17014,N_12563,N_13199);
and U17015 (N_17015,N_13947,N_13021);
and U17016 (N_17016,N_11335,N_14716);
nand U17017 (N_17017,N_12531,N_14501);
and U17018 (N_17018,N_13269,N_11254);
and U17019 (N_17019,N_14158,N_11048);
or U17020 (N_17020,N_13956,N_12586);
nand U17021 (N_17021,N_12970,N_11031);
or U17022 (N_17022,N_11800,N_14433);
nor U17023 (N_17023,N_11391,N_12878);
and U17024 (N_17024,N_14060,N_11337);
nor U17025 (N_17025,N_11587,N_14400);
and U17026 (N_17026,N_11764,N_13374);
xor U17027 (N_17027,N_12850,N_13133);
or U17028 (N_17028,N_10780,N_13019);
and U17029 (N_17029,N_14193,N_13399);
or U17030 (N_17030,N_12419,N_13572);
or U17031 (N_17031,N_13726,N_10839);
or U17032 (N_17032,N_14198,N_10697);
nor U17033 (N_17033,N_13853,N_13064);
or U17034 (N_17034,N_12829,N_13746);
nand U17035 (N_17035,N_14854,N_10997);
or U17036 (N_17036,N_13840,N_12437);
nand U17037 (N_17037,N_10948,N_11869);
xnor U17038 (N_17038,N_10772,N_11328);
nor U17039 (N_17039,N_12976,N_13596);
nand U17040 (N_17040,N_11320,N_12213);
and U17041 (N_17041,N_14418,N_11857);
and U17042 (N_17042,N_11198,N_11915);
and U17043 (N_17043,N_11845,N_14981);
or U17044 (N_17044,N_11221,N_10147);
nor U17045 (N_17045,N_12090,N_12021);
nand U17046 (N_17046,N_14720,N_11608);
nand U17047 (N_17047,N_10763,N_11528);
and U17048 (N_17048,N_12841,N_10886);
xnor U17049 (N_17049,N_11220,N_14005);
or U17050 (N_17050,N_10656,N_13816);
nor U17051 (N_17051,N_13175,N_14086);
or U17052 (N_17052,N_11137,N_13475);
nand U17053 (N_17053,N_14996,N_11419);
xor U17054 (N_17054,N_13672,N_10778);
and U17055 (N_17055,N_10615,N_13406);
and U17056 (N_17056,N_11558,N_12768);
xor U17057 (N_17057,N_14742,N_14814);
nor U17058 (N_17058,N_12807,N_10266);
and U17059 (N_17059,N_13873,N_14856);
or U17060 (N_17060,N_12517,N_14278);
and U17061 (N_17061,N_13637,N_14225);
nor U17062 (N_17062,N_11887,N_11734);
nor U17063 (N_17063,N_10790,N_14245);
or U17064 (N_17064,N_13874,N_13449);
xor U17065 (N_17065,N_12370,N_10744);
and U17066 (N_17066,N_13634,N_14154);
or U17067 (N_17067,N_11307,N_12249);
and U17068 (N_17068,N_12395,N_11038);
nor U17069 (N_17069,N_13013,N_12999);
or U17070 (N_17070,N_12191,N_13820);
or U17071 (N_17071,N_10626,N_11072);
or U17072 (N_17072,N_11348,N_10893);
and U17073 (N_17073,N_10509,N_12143);
or U17074 (N_17074,N_11049,N_14099);
and U17075 (N_17075,N_14375,N_11596);
and U17076 (N_17076,N_10113,N_10690);
or U17077 (N_17077,N_11635,N_12813);
nor U17078 (N_17078,N_14351,N_13831);
or U17079 (N_17079,N_10577,N_13179);
or U17080 (N_17080,N_10801,N_11376);
nand U17081 (N_17081,N_11174,N_13696);
or U17082 (N_17082,N_14427,N_12209);
or U17083 (N_17083,N_14177,N_14143);
nand U17084 (N_17084,N_11991,N_12644);
or U17085 (N_17085,N_11378,N_11163);
nor U17086 (N_17086,N_14448,N_13496);
nor U17087 (N_17087,N_10556,N_10123);
nor U17088 (N_17088,N_13282,N_13659);
nor U17089 (N_17089,N_14257,N_13173);
xnor U17090 (N_17090,N_13188,N_14588);
nor U17091 (N_17091,N_10942,N_10669);
nor U17092 (N_17092,N_10817,N_11722);
or U17093 (N_17093,N_10200,N_13938);
xnor U17094 (N_17094,N_14723,N_13027);
or U17095 (N_17095,N_10597,N_10391);
nor U17096 (N_17096,N_12782,N_14811);
or U17097 (N_17097,N_13894,N_10421);
nand U17098 (N_17098,N_11573,N_12251);
or U17099 (N_17099,N_12003,N_14568);
xor U17100 (N_17100,N_14116,N_14368);
and U17101 (N_17101,N_13168,N_11346);
and U17102 (N_17102,N_11767,N_11849);
and U17103 (N_17103,N_11203,N_11510);
nor U17104 (N_17104,N_10105,N_12397);
or U17105 (N_17105,N_14608,N_14836);
or U17106 (N_17106,N_14169,N_11401);
nor U17107 (N_17107,N_14641,N_12646);
or U17108 (N_17108,N_12222,N_13882);
nand U17109 (N_17109,N_13167,N_14925);
nor U17110 (N_17110,N_11856,N_10111);
and U17111 (N_17111,N_10354,N_12686);
or U17112 (N_17112,N_14888,N_12823);
nand U17113 (N_17113,N_14553,N_11152);
and U17114 (N_17114,N_10636,N_13154);
xnor U17115 (N_17115,N_10498,N_14309);
or U17116 (N_17116,N_11204,N_10010);
nand U17117 (N_17117,N_12632,N_10397);
xnor U17118 (N_17118,N_10293,N_13667);
and U17119 (N_17119,N_11132,N_14301);
xnor U17120 (N_17120,N_12276,N_10300);
or U17121 (N_17121,N_10432,N_14951);
nor U17122 (N_17122,N_14538,N_10405);
or U17123 (N_17123,N_10052,N_13248);
nor U17124 (N_17124,N_12665,N_12924);
nand U17125 (N_17125,N_13981,N_13893);
nor U17126 (N_17126,N_13800,N_12359);
xor U17127 (N_17127,N_13931,N_13690);
nand U17128 (N_17128,N_12610,N_12979);
nand U17129 (N_17129,N_11065,N_12922);
or U17130 (N_17130,N_13476,N_11389);
nand U17131 (N_17131,N_13470,N_11826);
nor U17132 (N_17132,N_13507,N_10506);
and U17133 (N_17133,N_10791,N_11705);
nor U17134 (N_17134,N_11177,N_14146);
nor U17135 (N_17135,N_14567,N_12810);
xnor U17136 (N_17136,N_12795,N_13075);
and U17137 (N_17137,N_12791,N_12286);
xor U17138 (N_17138,N_12364,N_12855);
and U17139 (N_17139,N_10822,N_11368);
nor U17140 (N_17140,N_12971,N_13664);
nor U17141 (N_17141,N_13803,N_10036);
nor U17142 (N_17142,N_14382,N_11802);
and U17143 (N_17143,N_10512,N_13801);
xnor U17144 (N_17144,N_11006,N_11611);
nor U17145 (N_17145,N_10803,N_12236);
and U17146 (N_17146,N_13297,N_14615);
nand U17147 (N_17147,N_10242,N_14025);
nor U17148 (N_17148,N_10244,N_13563);
nand U17149 (N_17149,N_13028,N_13466);
nor U17150 (N_17150,N_11493,N_11593);
xor U17151 (N_17151,N_13872,N_11167);
and U17152 (N_17152,N_13608,N_11195);
or U17153 (N_17153,N_12179,N_14672);
nor U17154 (N_17154,N_10729,N_14703);
or U17155 (N_17155,N_12525,N_12460);
or U17156 (N_17156,N_12229,N_10435);
and U17157 (N_17157,N_14503,N_13020);
or U17158 (N_17158,N_10146,N_13205);
nand U17159 (N_17159,N_12341,N_11360);
nor U17160 (N_17160,N_13837,N_12619);
nand U17161 (N_17161,N_14200,N_10271);
or U17162 (N_17162,N_13516,N_13736);
nor U17163 (N_17163,N_13037,N_10190);
nor U17164 (N_17164,N_10368,N_13367);
or U17165 (N_17165,N_12198,N_12454);
xor U17166 (N_17166,N_13276,N_14490);
nand U17167 (N_17167,N_10008,N_14882);
xnor U17168 (N_17168,N_13402,N_13416);
nor U17169 (N_17169,N_12671,N_13531);
nor U17170 (N_17170,N_10080,N_12439);
nand U17171 (N_17171,N_13675,N_10434);
nand U17172 (N_17172,N_10758,N_11421);
xnor U17173 (N_17173,N_14598,N_10404);
nand U17174 (N_17174,N_13491,N_10179);
nor U17175 (N_17175,N_14574,N_10505);
xor U17176 (N_17176,N_10340,N_12849);
nor U17177 (N_17177,N_14817,N_12260);
nand U17178 (N_17178,N_11294,N_11272);
and U17179 (N_17179,N_10936,N_14114);
nor U17180 (N_17180,N_14195,N_13991);
and U17181 (N_17181,N_14384,N_11867);
xnor U17182 (N_17182,N_11353,N_11662);
nor U17183 (N_17183,N_13471,N_14552);
or U17184 (N_17184,N_11379,N_12944);
nand U17185 (N_17185,N_14746,N_14839);
nand U17186 (N_17186,N_10903,N_11313);
or U17187 (N_17187,N_13794,N_12949);
nand U17188 (N_17188,N_11836,N_11478);
nor U17189 (N_17189,N_13750,N_10203);
nor U17190 (N_17190,N_10925,N_14141);
nor U17191 (N_17191,N_13751,N_13589);
nor U17192 (N_17192,N_13071,N_12955);
or U17193 (N_17193,N_13335,N_12264);
nand U17194 (N_17194,N_11561,N_13519);
nand U17195 (N_17195,N_14564,N_13223);
or U17196 (N_17196,N_11851,N_13329);
and U17197 (N_17197,N_14323,N_11490);
nor U17198 (N_17198,N_14437,N_12835);
or U17199 (N_17199,N_13892,N_13709);
or U17200 (N_17200,N_11312,N_14600);
nor U17201 (N_17201,N_11588,N_12342);
nor U17202 (N_17202,N_13743,N_11938);
and U17203 (N_17203,N_14605,N_13231);
nand U17204 (N_17204,N_12668,N_12914);
nor U17205 (N_17205,N_14028,N_14887);
nand U17206 (N_17206,N_13932,N_12842);
nand U17207 (N_17207,N_10694,N_13140);
and U17208 (N_17208,N_12696,N_11334);
nand U17209 (N_17209,N_14034,N_10588);
nor U17210 (N_17210,N_11020,N_13018);
xor U17211 (N_17211,N_14941,N_12578);
or U17212 (N_17212,N_10700,N_11808);
nor U17213 (N_17213,N_10560,N_13772);
or U17214 (N_17214,N_12871,N_10045);
nand U17215 (N_17215,N_13358,N_11910);
nor U17216 (N_17216,N_13186,N_13192);
or U17217 (N_17217,N_13914,N_12405);
and U17218 (N_17218,N_14725,N_13034);
or U17219 (N_17219,N_11736,N_10294);
and U17220 (N_17220,N_14670,N_13210);
or U17221 (N_17221,N_12105,N_11159);
nor U17222 (N_17222,N_12182,N_10450);
nand U17223 (N_17223,N_14279,N_10221);
and U17224 (N_17224,N_14607,N_12353);
or U17225 (N_17225,N_10468,N_14188);
or U17226 (N_17226,N_12895,N_14863);
and U17227 (N_17227,N_13156,N_10552);
nand U17228 (N_17228,N_11228,N_11837);
and U17229 (N_17229,N_11701,N_13738);
or U17230 (N_17230,N_13218,N_14632);
xor U17231 (N_17231,N_10127,N_10107);
xor U17232 (N_17232,N_11273,N_13036);
xor U17233 (N_17233,N_10945,N_13590);
or U17234 (N_17234,N_13079,N_14541);
nor U17235 (N_17235,N_12618,N_14751);
or U17236 (N_17236,N_13959,N_12974);
nand U17237 (N_17237,N_12204,N_13620);
nand U17238 (N_17238,N_13592,N_12650);
and U17239 (N_17239,N_12274,N_10711);
xor U17240 (N_17240,N_14361,N_11676);
or U17241 (N_17241,N_12616,N_11598);
and U17242 (N_17242,N_14388,N_13096);
nor U17243 (N_17243,N_11627,N_12372);
nor U17244 (N_17244,N_14883,N_12921);
or U17245 (N_17245,N_11476,N_12630);
or U17246 (N_17246,N_12633,N_13257);
and U17247 (N_17247,N_13031,N_14046);
nor U17248 (N_17248,N_10043,N_13814);
and U17249 (N_17249,N_14520,N_13373);
or U17250 (N_17250,N_14771,N_12057);
nand U17251 (N_17251,N_12241,N_12593);
nand U17252 (N_17252,N_14168,N_13418);
nand U17253 (N_17253,N_12952,N_12240);
and U17254 (N_17254,N_10813,N_12801);
nand U17255 (N_17255,N_11964,N_10906);
nor U17256 (N_17256,N_10731,N_12815);
or U17257 (N_17257,N_12464,N_12597);
nand U17258 (N_17258,N_13047,N_11633);
and U17259 (N_17259,N_14208,N_10410);
nor U17260 (N_17260,N_14566,N_12032);
nor U17261 (N_17261,N_14093,N_12409);
or U17262 (N_17262,N_11369,N_14159);
nand U17263 (N_17263,N_14536,N_12659);
xnor U17264 (N_17264,N_13083,N_10691);
nand U17265 (N_17265,N_10520,N_12777);
nor U17266 (N_17266,N_11000,N_11745);
xnor U17267 (N_17267,N_14684,N_13759);
nor U17268 (N_17268,N_13201,N_13022);
nand U17269 (N_17269,N_13184,N_12972);
or U17270 (N_17270,N_14978,N_12780);
xor U17271 (N_17271,N_11984,N_11912);
or U17272 (N_17272,N_13176,N_12507);
xor U17273 (N_17273,N_11390,N_11828);
or U17274 (N_17274,N_12530,N_12000);
nor U17275 (N_17275,N_11233,N_13953);
and U17276 (N_17276,N_14486,N_13560);
and U17277 (N_17277,N_11269,N_11171);
or U17278 (N_17278,N_11216,N_10684);
xnor U17279 (N_17279,N_13122,N_11283);
nor U17280 (N_17280,N_11824,N_10357);
nand U17281 (N_17281,N_14690,N_10977);
xor U17282 (N_17282,N_12147,N_14560);
xor U17283 (N_17283,N_11534,N_10276);
nor U17284 (N_17284,N_10050,N_13606);
nand U17285 (N_17285,N_12747,N_11443);
nand U17286 (N_17286,N_11278,N_11235);
or U17287 (N_17287,N_11681,N_10873);
xor U17288 (N_17288,N_13654,N_13542);
or U17289 (N_17289,N_11480,N_13336);
or U17290 (N_17290,N_14417,N_12441);
nor U17291 (N_17291,N_11164,N_12798);
nand U17292 (N_17292,N_10424,N_13318);
nand U17293 (N_17293,N_14394,N_10593);
nand U17294 (N_17294,N_11375,N_14890);
and U17295 (N_17295,N_12088,N_12212);
nor U17296 (N_17296,N_11208,N_13319);
nand U17297 (N_17297,N_11891,N_13528);
nand U17298 (N_17298,N_11647,N_12077);
nor U17299 (N_17299,N_14343,N_14464);
and U17300 (N_17300,N_10650,N_10993);
nand U17301 (N_17301,N_10101,N_10359);
nand U17302 (N_17302,N_11459,N_13657);
nor U17303 (N_17303,N_14074,N_14451);
or U17304 (N_17304,N_11944,N_12030);
nand U17305 (N_17305,N_11537,N_10503);
and U17306 (N_17306,N_14263,N_14054);
and U17307 (N_17307,N_12500,N_13208);
and U17308 (N_17308,N_10377,N_12061);
nor U17309 (N_17309,N_10515,N_11882);
nand U17310 (N_17310,N_10140,N_13945);
and U17311 (N_17311,N_10834,N_12303);
nor U17312 (N_17312,N_13871,N_11922);
or U17313 (N_17313,N_14637,N_12762);
or U17314 (N_17314,N_11081,N_10484);
nand U17315 (N_17315,N_13413,N_11652);
nand U17316 (N_17316,N_12821,N_11657);
or U17317 (N_17317,N_11791,N_13467);
nand U17318 (N_17318,N_10068,N_14284);
and U17319 (N_17319,N_13907,N_13754);
or U17320 (N_17320,N_14993,N_12722);
and U17321 (N_17321,N_11949,N_14341);
nand U17322 (N_17322,N_11366,N_14256);
nor U17323 (N_17323,N_12863,N_13360);
or U17324 (N_17324,N_13351,N_11327);
and U17325 (N_17325,N_14994,N_13334);
and U17326 (N_17326,N_13091,N_10594);
or U17327 (N_17327,N_11576,N_14861);
or U17328 (N_17328,N_10403,N_11556);
or U17329 (N_17329,N_14380,N_13017);
or U17330 (N_17330,N_13495,N_10098);
or U17331 (N_17331,N_13941,N_10712);
nand U17332 (N_17332,N_14739,N_11962);
nand U17333 (N_17333,N_14493,N_12966);
and U17334 (N_17334,N_10732,N_13233);
nor U17335 (N_17335,N_14877,N_12776);
nand U17336 (N_17336,N_11844,N_12022);
nand U17337 (N_17337,N_11304,N_12903);
or U17338 (N_17338,N_13049,N_10292);
or U17339 (N_17339,N_12371,N_12435);
nor U17340 (N_17340,N_12089,N_14397);
nand U17341 (N_17341,N_12988,N_14681);
and U17342 (N_17342,N_11343,N_13862);
nor U17343 (N_17343,N_10070,N_11029);
nor U17344 (N_17344,N_13805,N_13640);
nand U17345 (N_17345,N_11885,N_11918);
or U17346 (N_17346,N_12950,N_13811);
and U17347 (N_17347,N_10336,N_12357);
xnor U17348 (N_17348,N_11497,N_10115);
and U17349 (N_17349,N_10418,N_13152);
and U17350 (N_17350,N_13272,N_14585);
and U17351 (N_17351,N_12820,N_12751);
and U17352 (N_17352,N_12197,N_13854);
xnor U17353 (N_17353,N_12015,N_14148);
nand U17354 (N_17354,N_12045,N_13723);
or U17355 (N_17355,N_13966,N_14561);
or U17356 (N_17356,N_11339,N_12543);
nor U17357 (N_17357,N_13550,N_14163);
xnor U17358 (N_17358,N_14842,N_13845);
nand U17359 (N_17359,N_12054,N_14466);
nand U17360 (N_17360,N_10458,N_14377);
xnor U17361 (N_17361,N_12189,N_10376);
nor U17362 (N_17362,N_12608,N_14613);
nor U17363 (N_17363,N_11754,N_10227);
nor U17364 (N_17364,N_14651,N_14591);
nor U17365 (N_17365,N_11691,N_11653);
nor U17366 (N_17366,N_10565,N_14401);
and U17367 (N_17367,N_13118,N_12205);
and U17368 (N_17368,N_10619,N_10120);
or U17369 (N_17369,N_12477,N_12752);
or U17370 (N_17370,N_10663,N_10209);
or U17371 (N_17371,N_14463,N_14694);
or U17372 (N_17372,N_11018,N_13045);
or U17373 (N_17373,N_11538,N_10141);
nor U17374 (N_17374,N_10956,N_13583);
xnor U17375 (N_17375,N_12293,N_10971);
or U17376 (N_17376,N_10751,N_14386);
nand U17377 (N_17377,N_11024,N_12697);
nand U17378 (N_17378,N_14396,N_12487);
nand U17379 (N_17379,N_13960,N_12997);
xnor U17380 (N_17380,N_13072,N_12172);
and U17381 (N_17381,N_14470,N_13539);
nor U17382 (N_17382,N_12528,N_13420);
nor U17383 (N_17383,N_12087,N_13365);
or U17384 (N_17384,N_11752,N_10567);
nor U17385 (N_17385,N_10595,N_10632);
xnor U17386 (N_17386,N_12161,N_11570);
and U17387 (N_17387,N_13181,N_14776);
or U17388 (N_17388,N_10298,N_11012);
nand U17389 (N_17389,N_13244,N_12545);
or U17390 (N_17390,N_11617,N_13670);
nor U17391 (N_17391,N_14781,N_12253);
and U17392 (N_17392,N_14202,N_14035);
or U17393 (N_17393,N_14281,N_14593);
nand U17394 (N_17394,N_10301,N_10487);
nor U17395 (N_17395,N_13543,N_13414);
nand U17396 (N_17396,N_10542,N_13498);
nand U17397 (N_17397,N_12865,N_13846);
or U17398 (N_17398,N_10794,N_11285);
and U17399 (N_17399,N_14714,N_10496);
nor U17400 (N_17400,N_10518,N_13044);
and U17401 (N_17401,N_10047,N_12743);
nand U17402 (N_17402,N_11212,N_11520);
nand U17403 (N_17403,N_14791,N_14474);
nand U17404 (N_17404,N_12739,N_11455);
xnor U17405 (N_17405,N_11716,N_13387);
nand U17406 (N_17406,N_11799,N_13605);
and U17407 (N_17407,N_13311,N_10071);
and U17408 (N_17408,N_14618,N_10398);
nor U17409 (N_17409,N_10628,N_10638);
and U17410 (N_17410,N_11026,N_12322);
nor U17411 (N_17411,N_13454,N_14073);
or U17412 (N_17412,N_12347,N_14077);
xnor U17413 (N_17413,N_10129,N_11993);
xnor U17414 (N_17414,N_10345,N_12379);
nor U17415 (N_17415,N_11118,N_12866);
and U17416 (N_17416,N_13708,N_10351);
nor U17417 (N_17417,N_14315,N_13077);
nor U17418 (N_17418,N_12122,N_10719);
nor U17419 (N_17419,N_14756,N_10554);
and U17420 (N_17420,N_13298,N_11146);
nand U17421 (N_17421,N_12792,N_14258);
xor U17422 (N_17422,N_13697,N_11123);
nand U17423 (N_17423,N_13136,N_11525);
or U17424 (N_17424,N_10406,N_11442);
and U17425 (N_17425,N_10341,N_13510);
nand U17426 (N_17426,N_14457,N_12873);
xnor U17427 (N_17427,N_12467,N_12734);
nand U17428 (N_17428,N_14699,N_14777);
and U17429 (N_17429,N_14767,N_12904);
or U17430 (N_17430,N_14840,N_14609);
nor U17431 (N_17431,N_12678,N_12244);
nand U17432 (N_17432,N_12601,N_13573);
xor U17433 (N_17433,N_14673,N_11811);
or U17434 (N_17434,N_11765,N_10396);
or U17435 (N_17435,N_12723,N_10420);
or U17436 (N_17436,N_12453,N_10944);
or U17437 (N_17437,N_14010,N_10603);
and U17438 (N_17438,N_13610,N_11684);
nor U17439 (N_17439,N_12973,N_13263);
and U17440 (N_17440,N_14614,N_14679);
nand U17441 (N_17441,N_13048,N_13538);
or U17442 (N_17442,N_12658,N_14669);
nor U17443 (N_17443,N_13419,N_12461);
or U17444 (N_17444,N_12533,N_13613);
or U17445 (N_17445,N_10733,N_10086);
and U17446 (N_17446,N_14254,N_10637);
and U17447 (N_17447,N_10262,N_11424);
and U17448 (N_17448,N_10843,N_12176);
nor U17449 (N_17449,N_12613,N_13781);
nand U17450 (N_17450,N_10685,N_13731);
and U17451 (N_17451,N_12376,N_11095);
nor U17452 (N_17452,N_10328,N_11707);
nand U17453 (N_17453,N_11080,N_11703);
and U17454 (N_17454,N_13126,N_13443);
nor U17455 (N_17455,N_13881,N_12194);
nand U17456 (N_17456,N_11495,N_10501);
and U17457 (N_17457,N_13339,N_10102);
nor U17458 (N_17458,N_11463,N_11948);
nand U17459 (N_17459,N_14995,N_12651);
nand U17460 (N_17460,N_14431,N_11927);
nand U17461 (N_17461,N_13889,N_10749);
or U17462 (N_17462,N_10596,N_13102);
nand U17463 (N_17463,N_11554,N_11398);
nand U17464 (N_17464,N_14369,N_14209);
xor U17465 (N_17465,N_10274,N_14205);
nand U17466 (N_17466,N_12558,N_13770);
nand U17467 (N_17467,N_13954,N_14531);
and U17468 (N_17468,N_12984,N_14952);
nand U17469 (N_17469,N_10614,N_13802);
nand U17470 (N_17470,N_13164,N_11111);
and U17471 (N_17471,N_10654,N_10845);
or U17472 (N_17472,N_13748,N_12440);
and U17473 (N_17473,N_13535,N_14019);
or U17474 (N_17474,N_11714,N_14935);
nor U17475 (N_17475,N_12297,N_11959);
nor U17476 (N_17476,N_11367,N_12965);
nand U17477 (N_17477,N_13869,N_12060);
or U17478 (N_17478,N_11906,N_14409);
nand U17479 (N_17479,N_11418,N_12690);
or U17480 (N_17480,N_13285,N_12068);
or U17481 (N_17481,N_14194,N_10335);
or U17482 (N_17482,N_12428,N_12442);
and U17483 (N_17483,N_10940,N_14138);
or U17484 (N_17484,N_11890,N_12986);
or U17485 (N_17485,N_10013,N_10562);
and U17486 (N_17486,N_13161,N_11507);
and U17487 (N_17487,N_14680,N_12539);
and U17488 (N_17488,N_12484,N_10309);
nand U17489 (N_17489,N_14557,N_13410);
nand U17490 (N_17490,N_13848,N_12399);
and U17491 (N_17491,N_12629,N_10275);
or U17492 (N_17492,N_14629,N_14453);
xor U17493 (N_17493,N_12181,N_13725);
nand U17494 (N_17494,N_11237,N_13485);
or U17495 (N_17495,N_14642,N_10151);
nor U17496 (N_17496,N_11498,N_14865);
or U17497 (N_17497,N_10767,N_10523);
nand U17498 (N_17498,N_10806,N_13293);
nor U17499 (N_17499,N_11530,N_11992);
nor U17500 (N_17500,N_12754,N_10862);
nand U17501 (N_17501,N_14526,N_12302);
and U17502 (N_17502,N_12252,N_13455);
xor U17503 (N_17503,N_14404,N_14928);
nand U17504 (N_17504,N_12382,N_11763);
or U17505 (N_17505,N_11440,N_14571);
or U17506 (N_17506,N_14583,N_11687);
nor U17507 (N_17507,N_10663,N_11517);
nand U17508 (N_17508,N_13318,N_14068);
and U17509 (N_17509,N_12454,N_14208);
and U17510 (N_17510,N_13546,N_12231);
nand U17511 (N_17511,N_11035,N_10188);
or U17512 (N_17512,N_12399,N_13720);
and U17513 (N_17513,N_14274,N_12178);
nor U17514 (N_17514,N_14609,N_12801);
nor U17515 (N_17515,N_14905,N_10695);
or U17516 (N_17516,N_14029,N_10697);
nor U17517 (N_17517,N_14995,N_14290);
nand U17518 (N_17518,N_14539,N_11370);
or U17519 (N_17519,N_12805,N_13025);
xor U17520 (N_17520,N_10714,N_11187);
nor U17521 (N_17521,N_12673,N_14165);
xnor U17522 (N_17522,N_12237,N_10526);
and U17523 (N_17523,N_10295,N_14279);
nor U17524 (N_17524,N_14751,N_12333);
and U17525 (N_17525,N_10950,N_10267);
or U17526 (N_17526,N_13093,N_12570);
nand U17527 (N_17527,N_14853,N_10766);
nor U17528 (N_17528,N_11032,N_10432);
and U17529 (N_17529,N_13147,N_10429);
xnor U17530 (N_17530,N_14212,N_13996);
nor U17531 (N_17531,N_12747,N_10053);
and U17532 (N_17532,N_13313,N_10250);
nor U17533 (N_17533,N_13560,N_12234);
or U17534 (N_17534,N_14097,N_11908);
nand U17535 (N_17535,N_13220,N_10260);
nor U17536 (N_17536,N_14052,N_10832);
nand U17537 (N_17537,N_11973,N_10997);
nand U17538 (N_17538,N_14030,N_14694);
nand U17539 (N_17539,N_11023,N_10798);
nor U17540 (N_17540,N_10330,N_13569);
and U17541 (N_17541,N_10399,N_10271);
nand U17542 (N_17542,N_14997,N_11745);
and U17543 (N_17543,N_13178,N_10524);
nand U17544 (N_17544,N_10155,N_11972);
or U17545 (N_17545,N_14163,N_10482);
nand U17546 (N_17546,N_12517,N_13296);
xnor U17547 (N_17547,N_14209,N_10800);
nand U17548 (N_17548,N_14913,N_12220);
xor U17549 (N_17549,N_11564,N_12630);
or U17550 (N_17550,N_12740,N_10951);
nand U17551 (N_17551,N_14420,N_13509);
nand U17552 (N_17552,N_12813,N_13531);
nand U17553 (N_17553,N_11030,N_14966);
or U17554 (N_17554,N_14882,N_11229);
or U17555 (N_17555,N_11385,N_11232);
or U17556 (N_17556,N_12393,N_10245);
nand U17557 (N_17557,N_14522,N_11016);
xnor U17558 (N_17558,N_14542,N_13918);
and U17559 (N_17559,N_10029,N_12366);
nor U17560 (N_17560,N_10113,N_11619);
or U17561 (N_17561,N_10882,N_14766);
nor U17562 (N_17562,N_13617,N_14465);
nand U17563 (N_17563,N_10167,N_10397);
xor U17564 (N_17564,N_13209,N_14000);
nor U17565 (N_17565,N_11274,N_12732);
and U17566 (N_17566,N_14180,N_14769);
nor U17567 (N_17567,N_10838,N_14881);
and U17568 (N_17568,N_11201,N_12946);
or U17569 (N_17569,N_10812,N_11053);
and U17570 (N_17570,N_14067,N_12914);
and U17571 (N_17571,N_14527,N_10618);
and U17572 (N_17572,N_10555,N_13382);
and U17573 (N_17573,N_12317,N_13713);
xor U17574 (N_17574,N_12383,N_13023);
nand U17575 (N_17575,N_10831,N_11298);
nand U17576 (N_17576,N_12182,N_14750);
or U17577 (N_17577,N_11697,N_14910);
or U17578 (N_17578,N_11778,N_11106);
nor U17579 (N_17579,N_10806,N_13541);
nand U17580 (N_17580,N_14922,N_13638);
nor U17581 (N_17581,N_13305,N_11113);
nand U17582 (N_17582,N_13822,N_12424);
nand U17583 (N_17583,N_11439,N_12452);
nand U17584 (N_17584,N_14722,N_13556);
nand U17585 (N_17585,N_12732,N_10922);
nand U17586 (N_17586,N_10258,N_13623);
xor U17587 (N_17587,N_11608,N_11174);
and U17588 (N_17588,N_13754,N_14712);
nand U17589 (N_17589,N_10214,N_13996);
or U17590 (N_17590,N_10151,N_14114);
xnor U17591 (N_17591,N_13831,N_10669);
nand U17592 (N_17592,N_10925,N_10177);
nand U17593 (N_17593,N_12887,N_11824);
nand U17594 (N_17594,N_12507,N_10442);
xor U17595 (N_17595,N_13327,N_10514);
and U17596 (N_17596,N_14518,N_11946);
or U17597 (N_17597,N_13501,N_12922);
or U17598 (N_17598,N_13738,N_13808);
nor U17599 (N_17599,N_13920,N_10400);
or U17600 (N_17600,N_14059,N_14940);
or U17601 (N_17601,N_10203,N_12255);
and U17602 (N_17602,N_11604,N_12169);
nand U17603 (N_17603,N_14346,N_12064);
and U17604 (N_17604,N_10437,N_13399);
xnor U17605 (N_17605,N_12384,N_13260);
nor U17606 (N_17606,N_10392,N_11446);
nand U17607 (N_17607,N_10222,N_11334);
nor U17608 (N_17608,N_14265,N_12595);
or U17609 (N_17609,N_11664,N_14010);
and U17610 (N_17610,N_10339,N_14350);
or U17611 (N_17611,N_14268,N_10463);
nand U17612 (N_17612,N_11206,N_11647);
or U17613 (N_17613,N_12441,N_12787);
nand U17614 (N_17614,N_10186,N_10323);
or U17615 (N_17615,N_11306,N_14156);
nand U17616 (N_17616,N_14242,N_14396);
xor U17617 (N_17617,N_11231,N_11795);
nand U17618 (N_17618,N_10324,N_10887);
nor U17619 (N_17619,N_10902,N_14687);
nand U17620 (N_17620,N_14373,N_13264);
and U17621 (N_17621,N_13063,N_13644);
or U17622 (N_17622,N_12283,N_14451);
and U17623 (N_17623,N_13373,N_10058);
nor U17624 (N_17624,N_11512,N_10995);
nand U17625 (N_17625,N_13016,N_14569);
or U17626 (N_17626,N_10117,N_11256);
and U17627 (N_17627,N_14756,N_11414);
xor U17628 (N_17628,N_13018,N_11290);
or U17629 (N_17629,N_11488,N_13642);
nor U17630 (N_17630,N_14310,N_14490);
xor U17631 (N_17631,N_10762,N_10528);
xor U17632 (N_17632,N_13192,N_12884);
or U17633 (N_17633,N_14138,N_14950);
nor U17634 (N_17634,N_10568,N_10114);
nor U17635 (N_17635,N_11857,N_10241);
and U17636 (N_17636,N_11654,N_14969);
xnor U17637 (N_17637,N_13116,N_11476);
or U17638 (N_17638,N_10476,N_13554);
nor U17639 (N_17639,N_13544,N_10716);
nand U17640 (N_17640,N_11505,N_10085);
and U17641 (N_17641,N_13712,N_11895);
nor U17642 (N_17642,N_14803,N_14276);
nand U17643 (N_17643,N_13257,N_10319);
and U17644 (N_17644,N_12048,N_14223);
nand U17645 (N_17645,N_12878,N_12018);
nand U17646 (N_17646,N_14759,N_14841);
or U17647 (N_17647,N_10985,N_14885);
nand U17648 (N_17648,N_13628,N_14965);
and U17649 (N_17649,N_12186,N_11605);
xor U17650 (N_17650,N_11319,N_10878);
xor U17651 (N_17651,N_13806,N_10514);
nand U17652 (N_17652,N_14134,N_12721);
nor U17653 (N_17653,N_14368,N_11630);
xor U17654 (N_17654,N_10869,N_10598);
nor U17655 (N_17655,N_13812,N_14156);
nand U17656 (N_17656,N_14629,N_14442);
nand U17657 (N_17657,N_11821,N_12191);
or U17658 (N_17658,N_11961,N_10286);
nand U17659 (N_17659,N_13773,N_11459);
nor U17660 (N_17660,N_11297,N_12125);
nand U17661 (N_17661,N_12330,N_14450);
xor U17662 (N_17662,N_13352,N_12453);
and U17663 (N_17663,N_13009,N_11908);
or U17664 (N_17664,N_14109,N_13118);
nor U17665 (N_17665,N_14279,N_12039);
nor U17666 (N_17666,N_14128,N_14504);
nand U17667 (N_17667,N_10973,N_12259);
and U17668 (N_17668,N_11265,N_10224);
nor U17669 (N_17669,N_12674,N_14779);
nor U17670 (N_17670,N_10354,N_11572);
nand U17671 (N_17671,N_12997,N_10285);
nand U17672 (N_17672,N_14892,N_12690);
and U17673 (N_17673,N_11052,N_13666);
or U17674 (N_17674,N_12752,N_10691);
xor U17675 (N_17675,N_12939,N_13246);
nor U17676 (N_17676,N_12030,N_11922);
or U17677 (N_17677,N_13182,N_10725);
nand U17678 (N_17678,N_12650,N_11068);
nand U17679 (N_17679,N_11509,N_14871);
nand U17680 (N_17680,N_14341,N_13957);
nor U17681 (N_17681,N_12019,N_11928);
xor U17682 (N_17682,N_13627,N_12064);
or U17683 (N_17683,N_12652,N_11756);
nand U17684 (N_17684,N_10007,N_12931);
nor U17685 (N_17685,N_14704,N_12290);
or U17686 (N_17686,N_10554,N_12592);
and U17687 (N_17687,N_13077,N_11105);
nand U17688 (N_17688,N_14188,N_14388);
or U17689 (N_17689,N_13966,N_13321);
nand U17690 (N_17690,N_12601,N_13220);
and U17691 (N_17691,N_10252,N_12079);
nand U17692 (N_17692,N_11026,N_12896);
and U17693 (N_17693,N_14478,N_13157);
and U17694 (N_17694,N_13022,N_12447);
nand U17695 (N_17695,N_13145,N_13230);
nand U17696 (N_17696,N_11254,N_13992);
nand U17697 (N_17697,N_14564,N_11059);
nand U17698 (N_17698,N_11071,N_12242);
or U17699 (N_17699,N_14087,N_10378);
and U17700 (N_17700,N_13932,N_12618);
and U17701 (N_17701,N_14944,N_13841);
and U17702 (N_17702,N_13331,N_14434);
nor U17703 (N_17703,N_14187,N_11186);
nand U17704 (N_17704,N_10660,N_13400);
xnor U17705 (N_17705,N_14091,N_12917);
or U17706 (N_17706,N_10084,N_12164);
or U17707 (N_17707,N_14016,N_12310);
nand U17708 (N_17708,N_13193,N_11156);
nor U17709 (N_17709,N_10150,N_10457);
nor U17710 (N_17710,N_13573,N_14784);
and U17711 (N_17711,N_11921,N_10132);
or U17712 (N_17712,N_10555,N_13542);
or U17713 (N_17713,N_10621,N_11076);
nand U17714 (N_17714,N_12855,N_11812);
nand U17715 (N_17715,N_11453,N_11349);
or U17716 (N_17716,N_14649,N_10344);
and U17717 (N_17717,N_13643,N_12856);
nand U17718 (N_17718,N_13317,N_14842);
xor U17719 (N_17719,N_10922,N_13203);
and U17720 (N_17720,N_10268,N_12584);
nor U17721 (N_17721,N_10351,N_11030);
and U17722 (N_17722,N_12157,N_10740);
xnor U17723 (N_17723,N_13539,N_14122);
nand U17724 (N_17724,N_11988,N_12058);
nand U17725 (N_17725,N_12534,N_10417);
or U17726 (N_17726,N_14901,N_10789);
xnor U17727 (N_17727,N_11594,N_14134);
or U17728 (N_17728,N_11360,N_12837);
or U17729 (N_17729,N_12399,N_14938);
or U17730 (N_17730,N_11805,N_12221);
and U17731 (N_17731,N_10219,N_14074);
nor U17732 (N_17732,N_10779,N_14221);
and U17733 (N_17733,N_12752,N_14054);
nor U17734 (N_17734,N_11648,N_12958);
nand U17735 (N_17735,N_14774,N_11682);
or U17736 (N_17736,N_10599,N_11162);
nor U17737 (N_17737,N_14351,N_11371);
and U17738 (N_17738,N_13162,N_14699);
or U17739 (N_17739,N_13319,N_13527);
or U17740 (N_17740,N_12748,N_13623);
or U17741 (N_17741,N_11588,N_13126);
and U17742 (N_17742,N_14858,N_14597);
nor U17743 (N_17743,N_13684,N_13622);
nand U17744 (N_17744,N_13672,N_10943);
and U17745 (N_17745,N_13122,N_10545);
and U17746 (N_17746,N_11533,N_13766);
or U17747 (N_17747,N_12405,N_14737);
nand U17748 (N_17748,N_13130,N_13932);
nand U17749 (N_17749,N_10139,N_11382);
or U17750 (N_17750,N_11213,N_14031);
or U17751 (N_17751,N_11633,N_13258);
nor U17752 (N_17752,N_13068,N_12137);
nor U17753 (N_17753,N_13350,N_12052);
xnor U17754 (N_17754,N_10504,N_13086);
and U17755 (N_17755,N_12947,N_13201);
nand U17756 (N_17756,N_12320,N_13449);
or U17757 (N_17757,N_10439,N_11298);
nand U17758 (N_17758,N_12200,N_12073);
nand U17759 (N_17759,N_12531,N_13278);
nor U17760 (N_17760,N_13775,N_10239);
nand U17761 (N_17761,N_13321,N_14107);
and U17762 (N_17762,N_14910,N_12789);
nand U17763 (N_17763,N_12862,N_10267);
nand U17764 (N_17764,N_13224,N_10905);
nor U17765 (N_17765,N_14283,N_10935);
or U17766 (N_17766,N_14502,N_13809);
nor U17767 (N_17767,N_14605,N_13059);
and U17768 (N_17768,N_12356,N_14748);
nor U17769 (N_17769,N_12220,N_14480);
xnor U17770 (N_17770,N_13767,N_10537);
or U17771 (N_17771,N_12099,N_14697);
nor U17772 (N_17772,N_14405,N_13647);
nor U17773 (N_17773,N_13526,N_10775);
nor U17774 (N_17774,N_13541,N_10565);
and U17775 (N_17775,N_10550,N_10052);
and U17776 (N_17776,N_13446,N_13555);
or U17777 (N_17777,N_11156,N_12441);
or U17778 (N_17778,N_14289,N_11997);
nand U17779 (N_17779,N_11454,N_10334);
and U17780 (N_17780,N_14791,N_11320);
and U17781 (N_17781,N_13690,N_12053);
and U17782 (N_17782,N_10907,N_11593);
or U17783 (N_17783,N_10836,N_12040);
nand U17784 (N_17784,N_14827,N_14007);
and U17785 (N_17785,N_10458,N_14546);
nand U17786 (N_17786,N_12027,N_10995);
xor U17787 (N_17787,N_11570,N_13045);
nor U17788 (N_17788,N_14617,N_14419);
nor U17789 (N_17789,N_12223,N_12462);
nor U17790 (N_17790,N_11507,N_11591);
and U17791 (N_17791,N_14239,N_13009);
or U17792 (N_17792,N_14906,N_13415);
or U17793 (N_17793,N_13051,N_10860);
or U17794 (N_17794,N_14449,N_14593);
nand U17795 (N_17795,N_13942,N_13805);
and U17796 (N_17796,N_11753,N_12871);
nand U17797 (N_17797,N_14327,N_14208);
or U17798 (N_17798,N_14910,N_12412);
and U17799 (N_17799,N_14678,N_13330);
xnor U17800 (N_17800,N_13763,N_10179);
xor U17801 (N_17801,N_13424,N_11561);
or U17802 (N_17802,N_13966,N_11417);
nor U17803 (N_17803,N_14830,N_10553);
or U17804 (N_17804,N_14635,N_10427);
nand U17805 (N_17805,N_11830,N_12214);
nand U17806 (N_17806,N_11125,N_14181);
nand U17807 (N_17807,N_13706,N_11555);
xnor U17808 (N_17808,N_13645,N_14290);
nand U17809 (N_17809,N_13337,N_11100);
or U17810 (N_17810,N_13699,N_11919);
or U17811 (N_17811,N_13003,N_11455);
nand U17812 (N_17812,N_11541,N_13151);
nand U17813 (N_17813,N_12001,N_10016);
xor U17814 (N_17814,N_13165,N_13983);
and U17815 (N_17815,N_13124,N_10537);
or U17816 (N_17816,N_12765,N_10713);
or U17817 (N_17817,N_14349,N_13938);
or U17818 (N_17818,N_14047,N_10076);
and U17819 (N_17819,N_10258,N_14246);
nand U17820 (N_17820,N_11013,N_12321);
nor U17821 (N_17821,N_14670,N_14323);
and U17822 (N_17822,N_12688,N_11985);
nor U17823 (N_17823,N_13660,N_13637);
or U17824 (N_17824,N_12784,N_13383);
or U17825 (N_17825,N_14201,N_13746);
and U17826 (N_17826,N_10931,N_13702);
and U17827 (N_17827,N_11161,N_12372);
xor U17828 (N_17828,N_13402,N_14938);
nor U17829 (N_17829,N_11233,N_11741);
nor U17830 (N_17830,N_14359,N_11276);
or U17831 (N_17831,N_13934,N_10853);
and U17832 (N_17832,N_13057,N_10981);
or U17833 (N_17833,N_13419,N_10148);
and U17834 (N_17834,N_10405,N_10963);
nor U17835 (N_17835,N_10713,N_13919);
or U17836 (N_17836,N_11107,N_12849);
and U17837 (N_17837,N_14987,N_11917);
nand U17838 (N_17838,N_11073,N_10720);
xor U17839 (N_17839,N_11200,N_11593);
and U17840 (N_17840,N_13091,N_12892);
or U17841 (N_17841,N_14412,N_11562);
and U17842 (N_17842,N_11471,N_11900);
or U17843 (N_17843,N_14965,N_13566);
nand U17844 (N_17844,N_12624,N_10213);
and U17845 (N_17845,N_13765,N_13413);
xor U17846 (N_17846,N_11816,N_13071);
xnor U17847 (N_17847,N_11182,N_12487);
or U17848 (N_17848,N_13159,N_11534);
nand U17849 (N_17849,N_13689,N_12421);
or U17850 (N_17850,N_12559,N_11382);
and U17851 (N_17851,N_14814,N_11597);
and U17852 (N_17852,N_11092,N_13624);
nand U17853 (N_17853,N_14408,N_10316);
nor U17854 (N_17854,N_13804,N_13930);
and U17855 (N_17855,N_11772,N_10702);
nand U17856 (N_17856,N_13166,N_14655);
nand U17857 (N_17857,N_13142,N_13289);
nor U17858 (N_17858,N_11364,N_12217);
and U17859 (N_17859,N_14758,N_10365);
nand U17860 (N_17860,N_14537,N_14041);
xor U17861 (N_17861,N_12728,N_13039);
and U17862 (N_17862,N_12538,N_11989);
xnor U17863 (N_17863,N_12875,N_10096);
nand U17864 (N_17864,N_12082,N_12619);
or U17865 (N_17865,N_10115,N_12758);
xnor U17866 (N_17866,N_13614,N_13361);
and U17867 (N_17867,N_13743,N_14035);
or U17868 (N_17868,N_11933,N_10188);
or U17869 (N_17869,N_14500,N_13506);
or U17870 (N_17870,N_10348,N_12084);
and U17871 (N_17871,N_12699,N_14948);
and U17872 (N_17872,N_14653,N_13181);
nand U17873 (N_17873,N_11838,N_10217);
nand U17874 (N_17874,N_14749,N_10363);
or U17875 (N_17875,N_11040,N_14220);
nor U17876 (N_17876,N_11097,N_14753);
or U17877 (N_17877,N_14051,N_12015);
nand U17878 (N_17878,N_10392,N_14221);
or U17879 (N_17879,N_10123,N_14110);
and U17880 (N_17880,N_12268,N_12113);
and U17881 (N_17881,N_12261,N_12651);
or U17882 (N_17882,N_13617,N_11186);
nor U17883 (N_17883,N_13034,N_14955);
or U17884 (N_17884,N_10557,N_14992);
xnor U17885 (N_17885,N_11165,N_13053);
nor U17886 (N_17886,N_13751,N_10115);
or U17887 (N_17887,N_13520,N_11838);
nor U17888 (N_17888,N_14871,N_12768);
and U17889 (N_17889,N_13835,N_13779);
nor U17890 (N_17890,N_11738,N_14856);
or U17891 (N_17891,N_14609,N_12496);
nor U17892 (N_17892,N_10476,N_14156);
and U17893 (N_17893,N_14876,N_11144);
nand U17894 (N_17894,N_13402,N_12336);
or U17895 (N_17895,N_13517,N_14957);
nand U17896 (N_17896,N_13087,N_12842);
nor U17897 (N_17897,N_13384,N_12716);
and U17898 (N_17898,N_13169,N_14651);
or U17899 (N_17899,N_12192,N_12533);
and U17900 (N_17900,N_11168,N_14462);
nand U17901 (N_17901,N_11797,N_10511);
and U17902 (N_17902,N_14359,N_13692);
nor U17903 (N_17903,N_11092,N_11571);
nor U17904 (N_17904,N_13059,N_13324);
and U17905 (N_17905,N_11653,N_10880);
or U17906 (N_17906,N_12755,N_11317);
nand U17907 (N_17907,N_11756,N_10110);
nor U17908 (N_17908,N_13997,N_12459);
nand U17909 (N_17909,N_12955,N_13285);
xor U17910 (N_17910,N_11463,N_11544);
and U17911 (N_17911,N_12439,N_10988);
nor U17912 (N_17912,N_12258,N_12325);
xnor U17913 (N_17913,N_14594,N_11411);
nor U17914 (N_17914,N_10310,N_13581);
nor U17915 (N_17915,N_14530,N_12525);
nand U17916 (N_17916,N_12900,N_10037);
nand U17917 (N_17917,N_14823,N_13806);
nor U17918 (N_17918,N_11962,N_13661);
nor U17919 (N_17919,N_11200,N_10167);
xnor U17920 (N_17920,N_11999,N_11482);
nor U17921 (N_17921,N_11667,N_11805);
nand U17922 (N_17922,N_10477,N_13585);
and U17923 (N_17923,N_11513,N_11931);
xnor U17924 (N_17924,N_13516,N_11742);
nand U17925 (N_17925,N_13426,N_10310);
or U17926 (N_17926,N_12587,N_11248);
and U17927 (N_17927,N_12281,N_14568);
xor U17928 (N_17928,N_12166,N_12707);
and U17929 (N_17929,N_10968,N_10929);
nor U17930 (N_17930,N_12497,N_10192);
or U17931 (N_17931,N_10272,N_13066);
and U17932 (N_17932,N_13731,N_14094);
nand U17933 (N_17933,N_10651,N_10373);
nand U17934 (N_17934,N_11024,N_10108);
nor U17935 (N_17935,N_13183,N_13417);
nand U17936 (N_17936,N_11305,N_10041);
or U17937 (N_17937,N_10820,N_10531);
xor U17938 (N_17938,N_12229,N_13405);
and U17939 (N_17939,N_12699,N_14999);
and U17940 (N_17940,N_10232,N_13598);
and U17941 (N_17941,N_13909,N_13925);
nand U17942 (N_17942,N_14878,N_14477);
nand U17943 (N_17943,N_13172,N_10089);
nand U17944 (N_17944,N_11133,N_12782);
nor U17945 (N_17945,N_14508,N_14917);
xnor U17946 (N_17946,N_12266,N_13348);
xnor U17947 (N_17947,N_12495,N_13649);
and U17948 (N_17948,N_10317,N_12879);
nand U17949 (N_17949,N_13585,N_12698);
nand U17950 (N_17950,N_11610,N_12004);
xor U17951 (N_17951,N_13541,N_11506);
or U17952 (N_17952,N_10299,N_11933);
nand U17953 (N_17953,N_13065,N_14405);
and U17954 (N_17954,N_10157,N_10095);
nand U17955 (N_17955,N_13201,N_11371);
and U17956 (N_17956,N_11887,N_10413);
or U17957 (N_17957,N_11011,N_12817);
or U17958 (N_17958,N_10041,N_12107);
nor U17959 (N_17959,N_10091,N_10477);
xnor U17960 (N_17960,N_14519,N_12633);
nor U17961 (N_17961,N_11840,N_13719);
nor U17962 (N_17962,N_10604,N_12969);
nand U17963 (N_17963,N_14797,N_11447);
nor U17964 (N_17964,N_12760,N_13109);
and U17965 (N_17965,N_13012,N_14055);
and U17966 (N_17966,N_11627,N_14755);
nor U17967 (N_17967,N_11352,N_12128);
and U17968 (N_17968,N_14703,N_12794);
or U17969 (N_17969,N_12425,N_11395);
nand U17970 (N_17970,N_14398,N_14139);
nor U17971 (N_17971,N_11586,N_10889);
nand U17972 (N_17972,N_10882,N_14747);
nand U17973 (N_17973,N_13119,N_12982);
nor U17974 (N_17974,N_11980,N_11347);
and U17975 (N_17975,N_12968,N_14755);
xor U17976 (N_17976,N_10060,N_14858);
or U17977 (N_17977,N_10182,N_10246);
nand U17978 (N_17978,N_10292,N_12848);
and U17979 (N_17979,N_13201,N_11878);
nand U17980 (N_17980,N_13802,N_10896);
nor U17981 (N_17981,N_10003,N_11162);
xnor U17982 (N_17982,N_14218,N_10601);
or U17983 (N_17983,N_10083,N_13409);
xor U17984 (N_17984,N_11655,N_11637);
nand U17985 (N_17985,N_14988,N_10540);
or U17986 (N_17986,N_13638,N_14201);
nor U17987 (N_17987,N_11156,N_14358);
and U17988 (N_17988,N_14867,N_11327);
or U17989 (N_17989,N_11930,N_10538);
and U17990 (N_17990,N_10118,N_11885);
and U17991 (N_17991,N_14901,N_12531);
nand U17992 (N_17992,N_12909,N_10227);
nor U17993 (N_17993,N_11699,N_12058);
nand U17994 (N_17994,N_14752,N_11845);
and U17995 (N_17995,N_14626,N_11013);
xor U17996 (N_17996,N_13301,N_10158);
and U17997 (N_17997,N_11576,N_11325);
nor U17998 (N_17998,N_10224,N_13656);
nand U17999 (N_17999,N_13967,N_12311);
or U18000 (N_18000,N_14821,N_12281);
nand U18001 (N_18001,N_12174,N_14149);
nor U18002 (N_18002,N_14172,N_12466);
and U18003 (N_18003,N_12099,N_14395);
nor U18004 (N_18004,N_12674,N_14970);
nor U18005 (N_18005,N_12667,N_13141);
nand U18006 (N_18006,N_14536,N_14777);
or U18007 (N_18007,N_12095,N_14421);
and U18008 (N_18008,N_11512,N_11653);
or U18009 (N_18009,N_12768,N_11712);
and U18010 (N_18010,N_11741,N_11460);
or U18011 (N_18011,N_12667,N_14630);
or U18012 (N_18012,N_11661,N_14234);
nand U18013 (N_18013,N_11307,N_11123);
nor U18014 (N_18014,N_13970,N_13151);
and U18015 (N_18015,N_12583,N_12204);
nand U18016 (N_18016,N_10268,N_13978);
and U18017 (N_18017,N_13350,N_11514);
or U18018 (N_18018,N_14668,N_12125);
or U18019 (N_18019,N_10661,N_10721);
xnor U18020 (N_18020,N_11028,N_14048);
xnor U18021 (N_18021,N_13509,N_11097);
nand U18022 (N_18022,N_11658,N_11292);
or U18023 (N_18023,N_10229,N_13755);
nor U18024 (N_18024,N_13594,N_12189);
or U18025 (N_18025,N_13774,N_10117);
nor U18026 (N_18026,N_14723,N_11749);
nand U18027 (N_18027,N_12659,N_14552);
xnor U18028 (N_18028,N_14606,N_11619);
or U18029 (N_18029,N_13368,N_10871);
nand U18030 (N_18030,N_13911,N_10812);
or U18031 (N_18031,N_14205,N_10266);
nor U18032 (N_18032,N_12644,N_13171);
or U18033 (N_18033,N_10685,N_11306);
nor U18034 (N_18034,N_11530,N_13869);
and U18035 (N_18035,N_10786,N_13998);
nor U18036 (N_18036,N_14133,N_10405);
or U18037 (N_18037,N_10142,N_10527);
nor U18038 (N_18038,N_13441,N_11206);
nand U18039 (N_18039,N_14474,N_13193);
xor U18040 (N_18040,N_10166,N_14052);
or U18041 (N_18041,N_14654,N_10739);
or U18042 (N_18042,N_13535,N_11345);
nor U18043 (N_18043,N_11614,N_10071);
and U18044 (N_18044,N_14109,N_11755);
nand U18045 (N_18045,N_10962,N_12640);
or U18046 (N_18046,N_13603,N_11716);
nand U18047 (N_18047,N_10043,N_10789);
nand U18048 (N_18048,N_11263,N_13378);
and U18049 (N_18049,N_14772,N_13240);
nor U18050 (N_18050,N_13994,N_13929);
nor U18051 (N_18051,N_10300,N_14638);
or U18052 (N_18052,N_11689,N_11385);
and U18053 (N_18053,N_13347,N_11200);
and U18054 (N_18054,N_11654,N_11675);
or U18055 (N_18055,N_12557,N_13768);
nand U18056 (N_18056,N_13281,N_12081);
xor U18057 (N_18057,N_11254,N_13251);
or U18058 (N_18058,N_11052,N_13881);
nand U18059 (N_18059,N_14662,N_12702);
xnor U18060 (N_18060,N_10473,N_11096);
and U18061 (N_18061,N_13609,N_11603);
xor U18062 (N_18062,N_13464,N_11391);
nor U18063 (N_18063,N_13673,N_13619);
or U18064 (N_18064,N_12146,N_13830);
nand U18065 (N_18065,N_11047,N_11151);
or U18066 (N_18066,N_10724,N_13469);
or U18067 (N_18067,N_10274,N_10128);
nor U18068 (N_18068,N_10204,N_13673);
nor U18069 (N_18069,N_14447,N_10355);
and U18070 (N_18070,N_14523,N_13803);
nor U18071 (N_18071,N_10664,N_14618);
nor U18072 (N_18072,N_12562,N_14448);
nor U18073 (N_18073,N_12160,N_10979);
and U18074 (N_18074,N_12021,N_11219);
nor U18075 (N_18075,N_13147,N_11007);
nor U18076 (N_18076,N_12101,N_12505);
or U18077 (N_18077,N_10923,N_10360);
nand U18078 (N_18078,N_10697,N_14415);
and U18079 (N_18079,N_14961,N_11541);
nor U18080 (N_18080,N_13002,N_14352);
nor U18081 (N_18081,N_13045,N_14895);
or U18082 (N_18082,N_14598,N_13398);
nand U18083 (N_18083,N_12824,N_13523);
nor U18084 (N_18084,N_10113,N_12334);
xnor U18085 (N_18085,N_11202,N_14364);
and U18086 (N_18086,N_12081,N_13058);
nand U18087 (N_18087,N_13327,N_14794);
or U18088 (N_18088,N_10576,N_14293);
or U18089 (N_18089,N_12169,N_14481);
nor U18090 (N_18090,N_10502,N_14642);
or U18091 (N_18091,N_14007,N_11578);
and U18092 (N_18092,N_11398,N_11283);
and U18093 (N_18093,N_13562,N_11112);
xor U18094 (N_18094,N_10016,N_11082);
or U18095 (N_18095,N_11518,N_13708);
and U18096 (N_18096,N_14949,N_10964);
and U18097 (N_18097,N_14570,N_12201);
nand U18098 (N_18098,N_11178,N_14765);
or U18099 (N_18099,N_11686,N_12300);
nor U18100 (N_18100,N_12916,N_10440);
and U18101 (N_18101,N_13336,N_14119);
nand U18102 (N_18102,N_10777,N_13101);
or U18103 (N_18103,N_11221,N_13651);
nand U18104 (N_18104,N_11913,N_11983);
or U18105 (N_18105,N_13572,N_12608);
and U18106 (N_18106,N_14635,N_10480);
or U18107 (N_18107,N_14543,N_10433);
and U18108 (N_18108,N_11931,N_13736);
nand U18109 (N_18109,N_10427,N_10255);
and U18110 (N_18110,N_11725,N_11670);
nand U18111 (N_18111,N_11156,N_11539);
and U18112 (N_18112,N_12014,N_14809);
xor U18113 (N_18113,N_10827,N_12502);
and U18114 (N_18114,N_14808,N_14779);
nand U18115 (N_18115,N_11007,N_11289);
or U18116 (N_18116,N_14566,N_10938);
nor U18117 (N_18117,N_12090,N_12160);
and U18118 (N_18118,N_13991,N_12072);
and U18119 (N_18119,N_13926,N_11342);
nand U18120 (N_18120,N_14961,N_13060);
or U18121 (N_18121,N_10569,N_13960);
and U18122 (N_18122,N_12999,N_10730);
nand U18123 (N_18123,N_14543,N_11876);
or U18124 (N_18124,N_14310,N_11426);
or U18125 (N_18125,N_10531,N_10080);
and U18126 (N_18126,N_11341,N_11192);
and U18127 (N_18127,N_10864,N_14046);
and U18128 (N_18128,N_10199,N_11330);
nand U18129 (N_18129,N_14447,N_11359);
or U18130 (N_18130,N_14197,N_13253);
and U18131 (N_18131,N_14213,N_10292);
nand U18132 (N_18132,N_14637,N_14969);
and U18133 (N_18133,N_11827,N_13823);
and U18134 (N_18134,N_12569,N_13677);
nand U18135 (N_18135,N_12960,N_11156);
nand U18136 (N_18136,N_11753,N_12300);
nor U18137 (N_18137,N_14634,N_10122);
or U18138 (N_18138,N_11757,N_14963);
xor U18139 (N_18139,N_11248,N_10712);
nand U18140 (N_18140,N_10489,N_10624);
and U18141 (N_18141,N_12288,N_11439);
and U18142 (N_18142,N_13981,N_12128);
or U18143 (N_18143,N_12991,N_13556);
nor U18144 (N_18144,N_12181,N_13952);
and U18145 (N_18145,N_12194,N_12222);
nor U18146 (N_18146,N_10806,N_14920);
and U18147 (N_18147,N_13750,N_14171);
and U18148 (N_18148,N_11870,N_10128);
and U18149 (N_18149,N_12260,N_10188);
or U18150 (N_18150,N_13350,N_10670);
nor U18151 (N_18151,N_14685,N_12481);
and U18152 (N_18152,N_11184,N_14197);
nor U18153 (N_18153,N_10951,N_11819);
xnor U18154 (N_18154,N_10143,N_11012);
and U18155 (N_18155,N_10258,N_10647);
nor U18156 (N_18156,N_11177,N_10073);
nor U18157 (N_18157,N_12574,N_10154);
nor U18158 (N_18158,N_14293,N_13408);
nand U18159 (N_18159,N_14037,N_13376);
or U18160 (N_18160,N_10563,N_14700);
nand U18161 (N_18161,N_12319,N_14922);
nor U18162 (N_18162,N_12024,N_12857);
or U18163 (N_18163,N_13867,N_11170);
nand U18164 (N_18164,N_14908,N_11326);
nand U18165 (N_18165,N_10670,N_14846);
or U18166 (N_18166,N_13732,N_13625);
and U18167 (N_18167,N_13055,N_11912);
nand U18168 (N_18168,N_14435,N_11592);
or U18169 (N_18169,N_14661,N_11440);
nand U18170 (N_18170,N_10056,N_10120);
nand U18171 (N_18171,N_13835,N_10978);
xor U18172 (N_18172,N_11965,N_12020);
or U18173 (N_18173,N_14144,N_10740);
nor U18174 (N_18174,N_10930,N_10410);
or U18175 (N_18175,N_12267,N_13618);
nor U18176 (N_18176,N_14656,N_12584);
xnor U18177 (N_18177,N_12879,N_12578);
xnor U18178 (N_18178,N_14879,N_11522);
or U18179 (N_18179,N_10482,N_12571);
nor U18180 (N_18180,N_10420,N_10311);
or U18181 (N_18181,N_11305,N_11725);
nor U18182 (N_18182,N_11580,N_11681);
nor U18183 (N_18183,N_13157,N_12883);
nand U18184 (N_18184,N_12778,N_14286);
and U18185 (N_18185,N_12524,N_11712);
or U18186 (N_18186,N_14387,N_13116);
or U18187 (N_18187,N_10110,N_14296);
nand U18188 (N_18188,N_12754,N_10784);
or U18189 (N_18189,N_12350,N_10497);
or U18190 (N_18190,N_11192,N_14452);
or U18191 (N_18191,N_12933,N_11724);
nor U18192 (N_18192,N_10994,N_13769);
nor U18193 (N_18193,N_14915,N_11701);
nand U18194 (N_18194,N_10239,N_10520);
nand U18195 (N_18195,N_14576,N_13889);
and U18196 (N_18196,N_11488,N_11967);
nor U18197 (N_18197,N_10785,N_12664);
nand U18198 (N_18198,N_12381,N_12821);
nor U18199 (N_18199,N_13272,N_10295);
and U18200 (N_18200,N_12947,N_10813);
nand U18201 (N_18201,N_12071,N_13258);
and U18202 (N_18202,N_11438,N_13878);
nand U18203 (N_18203,N_11432,N_10478);
nand U18204 (N_18204,N_14327,N_13628);
and U18205 (N_18205,N_14449,N_11779);
or U18206 (N_18206,N_13607,N_14372);
nand U18207 (N_18207,N_12129,N_12085);
or U18208 (N_18208,N_11805,N_11477);
nor U18209 (N_18209,N_12994,N_13990);
nand U18210 (N_18210,N_12974,N_13262);
nand U18211 (N_18211,N_12073,N_11717);
or U18212 (N_18212,N_10997,N_13199);
nand U18213 (N_18213,N_10637,N_10149);
or U18214 (N_18214,N_10829,N_13020);
nand U18215 (N_18215,N_13654,N_14243);
nand U18216 (N_18216,N_10170,N_14148);
or U18217 (N_18217,N_14585,N_12284);
nand U18218 (N_18218,N_12938,N_12455);
and U18219 (N_18219,N_14854,N_12797);
nand U18220 (N_18220,N_14124,N_14019);
or U18221 (N_18221,N_13218,N_10848);
and U18222 (N_18222,N_10511,N_13601);
or U18223 (N_18223,N_13003,N_11008);
nor U18224 (N_18224,N_14021,N_13418);
and U18225 (N_18225,N_13749,N_12273);
and U18226 (N_18226,N_11884,N_12111);
nand U18227 (N_18227,N_14178,N_13173);
or U18228 (N_18228,N_13505,N_11993);
and U18229 (N_18229,N_12779,N_10733);
nand U18230 (N_18230,N_10563,N_10689);
or U18231 (N_18231,N_12469,N_12819);
nor U18232 (N_18232,N_13490,N_12671);
nor U18233 (N_18233,N_14779,N_14678);
xnor U18234 (N_18234,N_11652,N_12540);
or U18235 (N_18235,N_13007,N_10142);
nor U18236 (N_18236,N_12873,N_11546);
or U18237 (N_18237,N_10121,N_10403);
nor U18238 (N_18238,N_11008,N_12250);
nand U18239 (N_18239,N_11805,N_10549);
nand U18240 (N_18240,N_12214,N_14611);
and U18241 (N_18241,N_13124,N_13315);
nor U18242 (N_18242,N_11520,N_10300);
and U18243 (N_18243,N_11439,N_10867);
nor U18244 (N_18244,N_10572,N_11495);
and U18245 (N_18245,N_10386,N_13819);
and U18246 (N_18246,N_10554,N_13688);
nor U18247 (N_18247,N_10626,N_10199);
or U18248 (N_18248,N_14145,N_11474);
xnor U18249 (N_18249,N_10378,N_14223);
and U18250 (N_18250,N_12645,N_12894);
and U18251 (N_18251,N_14565,N_10263);
xnor U18252 (N_18252,N_13417,N_12739);
nand U18253 (N_18253,N_14281,N_14853);
or U18254 (N_18254,N_14828,N_14093);
nand U18255 (N_18255,N_13988,N_10700);
xnor U18256 (N_18256,N_12182,N_11818);
nor U18257 (N_18257,N_11493,N_11607);
and U18258 (N_18258,N_14654,N_14303);
nand U18259 (N_18259,N_11093,N_14381);
xnor U18260 (N_18260,N_12522,N_11116);
or U18261 (N_18261,N_10451,N_10842);
or U18262 (N_18262,N_12437,N_11205);
or U18263 (N_18263,N_13352,N_11073);
nand U18264 (N_18264,N_13602,N_13585);
nand U18265 (N_18265,N_12433,N_12181);
nor U18266 (N_18266,N_13365,N_11221);
and U18267 (N_18267,N_10424,N_12069);
and U18268 (N_18268,N_13030,N_12623);
nor U18269 (N_18269,N_13530,N_14066);
or U18270 (N_18270,N_10120,N_14406);
nand U18271 (N_18271,N_13159,N_14513);
or U18272 (N_18272,N_13800,N_10795);
and U18273 (N_18273,N_10839,N_10108);
and U18274 (N_18274,N_13322,N_13694);
nand U18275 (N_18275,N_12968,N_12060);
nand U18276 (N_18276,N_14029,N_12489);
and U18277 (N_18277,N_12563,N_12456);
nor U18278 (N_18278,N_11022,N_14138);
nand U18279 (N_18279,N_10769,N_14219);
xnor U18280 (N_18280,N_12602,N_14149);
and U18281 (N_18281,N_10134,N_14085);
and U18282 (N_18282,N_12980,N_11332);
and U18283 (N_18283,N_13729,N_12127);
and U18284 (N_18284,N_12965,N_11443);
or U18285 (N_18285,N_13420,N_13045);
nor U18286 (N_18286,N_14237,N_11858);
nand U18287 (N_18287,N_13423,N_10886);
and U18288 (N_18288,N_10235,N_10427);
and U18289 (N_18289,N_12882,N_13800);
and U18290 (N_18290,N_11456,N_10338);
and U18291 (N_18291,N_14597,N_13200);
and U18292 (N_18292,N_13414,N_11203);
nand U18293 (N_18293,N_10225,N_14420);
or U18294 (N_18294,N_13082,N_13475);
nand U18295 (N_18295,N_14612,N_11327);
or U18296 (N_18296,N_13123,N_10513);
xor U18297 (N_18297,N_10694,N_12905);
nor U18298 (N_18298,N_13570,N_10426);
nand U18299 (N_18299,N_10807,N_13391);
or U18300 (N_18300,N_13505,N_14398);
nand U18301 (N_18301,N_12004,N_13475);
nand U18302 (N_18302,N_10254,N_14740);
nor U18303 (N_18303,N_13279,N_14871);
or U18304 (N_18304,N_10988,N_12734);
or U18305 (N_18305,N_14987,N_14142);
or U18306 (N_18306,N_10955,N_12672);
nand U18307 (N_18307,N_13882,N_13112);
nor U18308 (N_18308,N_10085,N_11607);
nor U18309 (N_18309,N_10522,N_12840);
and U18310 (N_18310,N_13484,N_13022);
nand U18311 (N_18311,N_10313,N_13987);
or U18312 (N_18312,N_12128,N_10024);
nor U18313 (N_18313,N_12231,N_12278);
nand U18314 (N_18314,N_13872,N_12452);
nor U18315 (N_18315,N_13205,N_14541);
nor U18316 (N_18316,N_11825,N_13734);
or U18317 (N_18317,N_10106,N_12984);
nand U18318 (N_18318,N_12217,N_13089);
and U18319 (N_18319,N_10690,N_13750);
or U18320 (N_18320,N_10634,N_10347);
nor U18321 (N_18321,N_14718,N_14074);
xor U18322 (N_18322,N_12850,N_13993);
and U18323 (N_18323,N_11441,N_10495);
and U18324 (N_18324,N_14904,N_14835);
nand U18325 (N_18325,N_13548,N_11621);
xnor U18326 (N_18326,N_13398,N_12059);
nand U18327 (N_18327,N_10673,N_11806);
xor U18328 (N_18328,N_14152,N_11536);
nand U18329 (N_18329,N_10706,N_13430);
and U18330 (N_18330,N_12461,N_12758);
nand U18331 (N_18331,N_12920,N_14162);
and U18332 (N_18332,N_13897,N_12264);
nor U18333 (N_18333,N_12183,N_12986);
nor U18334 (N_18334,N_11608,N_10509);
or U18335 (N_18335,N_11872,N_12859);
nand U18336 (N_18336,N_13060,N_14218);
nand U18337 (N_18337,N_14534,N_14121);
or U18338 (N_18338,N_12303,N_12893);
nor U18339 (N_18339,N_14588,N_12443);
or U18340 (N_18340,N_14650,N_11237);
nand U18341 (N_18341,N_14643,N_13256);
nand U18342 (N_18342,N_10222,N_10926);
nand U18343 (N_18343,N_12052,N_10437);
or U18344 (N_18344,N_11889,N_14420);
nor U18345 (N_18345,N_12781,N_12912);
nor U18346 (N_18346,N_12788,N_13867);
nor U18347 (N_18347,N_11259,N_10481);
xor U18348 (N_18348,N_14439,N_11212);
xor U18349 (N_18349,N_12145,N_13573);
and U18350 (N_18350,N_12358,N_10792);
and U18351 (N_18351,N_14595,N_11013);
nand U18352 (N_18352,N_13738,N_11602);
and U18353 (N_18353,N_10418,N_10165);
nor U18354 (N_18354,N_14276,N_11793);
nor U18355 (N_18355,N_12659,N_13649);
xor U18356 (N_18356,N_12697,N_11595);
nand U18357 (N_18357,N_13627,N_11857);
and U18358 (N_18358,N_12513,N_14307);
nand U18359 (N_18359,N_11591,N_13392);
or U18360 (N_18360,N_13888,N_12734);
or U18361 (N_18361,N_11071,N_13391);
or U18362 (N_18362,N_12631,N_13183);
xor U18363 (N_18363,N_13103,N_10375);
or U18364 (N_18364,N_11002,N_14660);
or U18365 (N_18365,N_12333,N_10269);
or U18366 (N_18366,N_10897,N_11597);
or U18367 (N_18367,N_10742,N_10057);
and U18368 (N_18368,N_14229,N_14872);
xor U18369 (N_18369,N_11614,N_10004);
xor U18370 (N_18370,N_13864,N_11118);
xor U18371 (N_18371,N_10948,N_13328);
nand U18372 (N_18372,N_11870,N_12187);
xor U18373 (N_18373,N_12342,N_10975);
and U18374 (N_18374,N_14646,N_14720);
and U18375 (N_18375,N_13995,N_13457);
or U18376 (N_18376,N_12886,N_12465);
and U18377 (N_18377,N_14200,N_11610);
nor U18378 (N_18378,N_11964,N_11837);
or U18379 (N_18379,N_13527,N_12242);
and U18380 (N_18380,N_12906,N_11156);
or U18381 (N_18381,N_12893,N_11333);
nor U18382 (N_18382,N_14241,N_11831);
nor U18383 (N_18383,N_12476,N_11167);
nand U18384 (N_18384,N_14350,N_12272);
and U18385 (N_18385,N_13314,N_12864);
nand U18386 (N_18386,N_13514,N_13229);
or U18387 (N_18387,N_14539,N_11661);
or U18388 (N_18388,N_10303,N_11673);
and U18389 (N_18389,N_14797,N_10043);
and U18390 (N_18390,N_14023,N_13502);
nand U18391 (N_18391,N_14071,N_13566);
nand U18392 (N_18392,N_11088,N_14320);
or U18393 (N_18393,N_11680,N_11038);
nand U18394 (N_18394,N_11457,N_10068);
or U18395 (N_18395,N_11453,N_12854);
nand U18396 (N_18396,N_13240,N_13094);
and U18397 (N_18397,N_11414,N_12072);
nand U18398 (N_18398,N_13374,N_14412);
or U18399 (N_18399,N_11692,N_11401);
or U18400 (N_18400,N_13881,N_14382);
xor U18401 (N_18401,N_10469,N_13952);
and U18402 (N_18402,N_11414,N_14386);
nor U18403 (N_18403,N_11460,N_11050);
or U18404 (N_18404,N_13678,N_12955);
and U18405 (N_18405,N_11975,N_11311);
and U18406 (N_18406,N_11826,N_14231);
xnor U18407 (N_18407,N_11206,N_14677);
nor U18408 (N_18408,N_13467,N_13290);
or U18409 (N_18409,N_11006,N_11015);
nand U18410 (N_18410,N_14407,N_11737);
and U18411 (N_18411,N_13032,N_10207);
nor U18412 (N_18412,N_13345,N_13409);
nor U18413 (N_18413,N_14922,N_11461);
nand U18414 (N_18414,N_13803,N_14902);
xor U18415 (N_18415,N_10185,N_10994);
and U18416 (N_18416,N_12360,N_10232);
or U18417 (N_18417,N_11874,N_13794);
or U18418 (N_18418,N_13680,N_12614);
nor U18419 (N_18419,N_13140,N_14091);
xor U18420 (N_18420,N_14856,N_12554);
nand U18421 (N_18421,N_12976,N_10082);
xnor U18422 (N_18422,N_12214,N_11207);
or U18423 (N_18423,N_10122,N_12907);
and U18424 (N_18424,N_11640,N_11533);
or U18425 (N_18425,N_14071,N_12153);
and U18426 (N_18426,N_12997,N_14753);
xnor U18427 (N_18427,N_13639,N_12452);
or U18428 (N_18428,N_10196,N_13995);
and U18429 (N_18429,N_10584,N_13415);
and U18430 (N_18430,N_11916,N_11101);
nand U18431 (N_18431,N_13413,N_10028);
or U18432 (N_18432,N_10126,N_14234);
nand U18433 (N_18433,N_14131,N_13987);
and U18434 (N_18434,N_12233,N_13709);
or U18435 (N_18435,N_13545,N_10875);
nand U18436 (N_18436,N_13402,N_12453);
xnor U18437 (N_18437,N_11254,N_14014);
xnor U18438 (N_18438,N_14041,N_14501);
and U18439 (N_18439,N_14703,N_11294);
and U18440 (N_18440,N_10255,N_12434);
xnor U18441 (N_18441,N_13815,N_14376);
and U18442 (N_18442,N_13326,N_13941);
or U18443 (N_18443,N_10091,N_13915);
and U18444 (N_18444,N_12124,N_10604);
xor U18445 (N_18445,N_14541,N_11585);
or U18446 (N_18446,N_14492,N_11933);
xor U18447 (N_18447,N_13586,N_10212);
and U18448 (N_18448,N_10926,N_14351);
nand U18449 (N_18449,N_11877,N_13515);
nand U18450 (N_18450,N_12391,N_11422);
or U18451 (N_18451,N_14129,N_14851);
xnor U18452 (N_18452,N_14278,N_14337);
nand U18453 (N_18453,N_10495,N_14582);
and U18454 (N_18454,N_14255,N_12839);
and U18455 (N_18455,N_10954,N_12674);
nor U18456 (N_18456,N_10640,N_13938);
and U18457 (N_18457,N_10024,N_13998);
or U18458 (N_18458,N_12486,N_14875);
and U18459 (N_18459,N_13073,N_11131);
or U18460 (N_18460,N_13259,N_13765);
nor U18461 (N_18461,N_11238,N_10329);
or U18462 (N_18462,N_14992,N_10601);
and U18463 (N_18463,N_11656,N_12512);
nand U18464 (N_18464,N_14070,N_12784);
nor U18465 (N_18465,N_11605,N_11263);
and U18466 (N_18466,N_12060,N_10225);
xor U18467 (N_18467,N_12981,N_14904);
nor U18468 (N_18468,N_10388,N_10334);
xor U18469 (N_18469,N_12105,N_10494);
nand U18470 (N_18470,N_10410,N_11187);
nand U18471 (N_18471,N_11913,N_13470);
or U18472 (N_18472,N_13132,N_10895);
nand U18473 (N_18473,N_12211,N_12049);
and U18474 (N_18474,N_11146,N_11288);
nor U18475 (N_18475,N_12261,N_14447);
and U18476 (N_18476,N_10323,N_14581);
nor U18477 (N_18477,N_11636,N_14831);
nor U18478 (N_18478,N_14895,N_14310);
xnor U18479 (N_18479,N_14326,N_11992);
nor U18480 (N_18480,N_10434,N_10656);
and U18481 (N_18481,N_13285,N_12147);
nand U18482 (N_18482,N_13102,N_13693);
nand U18483 (N_18483,N_12529,N_10067);
and U18484 (N_18484,N_11437,N_11612);
nand U18485 (N_18485,N_13264,N_13875);
nand U18486 (N_18486,N_13080,N_13509);
or U18487 (N_18487,N_13024,N_11250);
nor U18488 (N_18488,N_11257,N_11577);
xnor U18489 (N_18489,N_13058,N_11108);
or U18490 (N_18490,N_12751,N_12355);
nor U18491 (N_18491,N_14905,N_12076);
nor U18492 (N_18492,N_12379,N_10457);
nor U18493 (N_18493,N_14589,N_14456);
nand U18494 (N_18494,N_11742,N_14597);
or U18495 (N_18495,N_12995,N_14381);
and U18496 (N_18496,N_13193,N_13971);
nor U18497 (N_18497,N_14128,N_12800);
nor U18498 (N_18498,N_13253,N_12620);
nor U18499 (N_18499,N_12558,N_14329);
nor U18500 (N_18500,N_11399,N_10967);
nor U18501 (N_18501,N_10473,N_11963);
nand U18502 (N_18502,N_14041,N_12032);
xnor U18503 (N_18503,N_13514,N_10105);
nand U18504 (N_18504,N_14729,N_12178);
or U18505 (N_18505,N_10278,N_14190);
or U18506 (N_18506,N_14636,N_11443);
and U18507 (N_18507,N_14622,N_12924);
nand U18508 (N_18508,N_12172,N_13461);
nand U18509 (N_18509,N_12317,N_13601);
nor U18510 (N_18510,N_11950,N_13150);
nand U18511 (N_18511,N_13050,N_13219);
nand U18512 (N_18512,N_13691,N_10731);
nor U18513 (N_18513,N_10704,N_11637);
or U18514 (N_18514,N_12489,N_12766);
xnor U18515 (N_18515,N_12909,N_14604);
nor U18516 (N_18516,N_14512,N_14707);
xor U18517 (N_18517,N_10344,N_13939);
or U18518 (N_18518,N_13117,N_10490);
or U18519 (N_18519,N_10776,N_13093);
nor U18520 (N_18520,N_13108,N_10554);
nand U18521 (N_18521,N_14784,N_14984);
and U18522 (N_18522,N_11295,N_10887);
or U18523 (N_18523,N_14475,N_14215);
and U18524 (N_18524,N_13977,N_11675);
nand U18525 (N_18525,N_11316,N_14821);
or U18526 (N_18526,N_12442,N_10585);
and U18527 (N_18527,N_11885,N_10843);
nand U18528 (N_18528,N_12250,N_14154);
and U18529 (N_18529,N_10121,N_11324);
or U18530 (N_18530,N_11462,N_14919);
xor U18531 (N_18531,N_10887,N_10295);
and U18532 (N_18532,N_12277,N_14739);
or U18533 (N_18533,N_13533,N_14949);
nor U18534 (N_18534,N_10781,N_10282);
or U18535 (N_18535,N_12805,N_10984);
and U18536 (N_18536,N_12812,N_13516);
and U18537 (N_18537,N_14269,N_12399);
or U18538 (N_18538,N_11404,N_14653);
and U18539 (N_18539,N_13024,N_10288);
nor U18540 (N_18540,N_14843,N_10182);
nor U18541 (N_18541,N_14227,N_14851);
nand U18542 (N_18542,N_13915,N_10316);
or U18543 (N_18543,N_11464,N_14807);
or U18544 (N_18544,N_14509,N_13165);
and U18545 (N_18545,N_14526,N_10854);
nand U18546 (N_18546,N_10300,N_10621);
xnor U18547 (N_18547,N_13820,N_14528);
nand U18548 (N_18548,N_12648,N_10651);
or U18549 (N_18549,N_13795,N_12793);
nor U18550 (N_18550,N_13562,N_11212);
or U18551 (N_18551,N_11368,N_11037);
nor U18552 (N_18552,N_14008,N_11589);
nor U18553 (N_18553,N_14016,N_14766);
and U18554 (N_18554,N_10015,N_14650);
and U18555 (N_18555,N_11880,N_11899);
nand U18556 (N_18556,N_11472,N_12659);
xnor U18557 (N_18557,N_13332,N_12638);
nand U18558 (N_18558,N_12148,N_11110);
nor U18559 (N_18559,N_13309,N_14498);
nor U18560 (N_18560,N_12308,N_12625);
nor U18561 (N_18561,N_10707,N_10298);
nor U18562 (N_18562,N_10168,N_11566);
xnor U18563 (N_18563,N_13996,N_10930);
or U18564 (N_18564,N_12024,N_11765);
xnor U18565 (N_18565,N_14400,N_13483);
nand U18566 (N_18566,N_12023,N_10108);
nand U18567 (N_18567,N_11347,N_14199);
or U18568 (N_18568,N_12753,N_13135);
and U18569 (N_18569,N_12263,N_13077);
nor U18570 (N_18570,N_10830,N_12794);
nand U18571 (N_18571,N_10786,N_12177);
or U18572 (N_18572,N_10253,N_11878);
nor U18573 (N_18573,N_10371,N_13583);
or U18574 (N_18574,N_10476,N_14126);
or U18575 (N_18575,N_12751,N_12180);
nor U18576 (N_18576,N_14618,N_12526);
and U18577 (N_18577,N_10203,N_10310);
and U18578 (N_18578,N_13372,N_12428);
nand U18579 (N_18579,N_11769,N_11376);
and U18580 (N_18580,N_11603,N_14366);
or U18581 (N_18581,N_14014,N_12588);
nor U18582 (N_18582,N_11064,N_14001);
nand U18583 (N_18583,N_10834,N_13467);
and U18584 (N_18584,N_13124,N_12406);
xor U18585 (N_18585,N_14798,N_14675);
and U18586 (N_18586,N_12230,N_14699);
nand U18587 (N_18587,N_12456,N_11993);
nor U18588 (N_18588,N_13043,N_11844);
nand U18589 (N_18589,N_13058,N_11763);
and U18590 (N_18590,N_12930,N_12446);
nand U18591 (N_18591,N_12212,N_10338);
and U18592 (N_18592,N_14675,N_11755);
and U18593 (N_18593,N_14423,N_10120);
nand U18594 (N_18594,N_14319,N_14779);
nand U18595 (N_18595,N_11125,N_11711);
nor U18596 (N_18596,N_10139,N_10830);
or U18597 (N_18597,N_13805,N_10536);
nand U18598 (N_18598,N_12603,N_11351);
nand U18599 (N_18599,N_13847,N_13750);
and U18600 (N_18600,N_12440,N_13750);
nor U18601 (N_18601,N_10622,N_13713);
nor U18602 (N_18602,N_11403,N_14706);
nor U18603 (N_18603,N_13149,N_11863);
nor U18604 (N_18604,N_13571,N_14147);
nand U18605 (N_18605,N_12146,N_12777);
and U18606 (N_18606,N_14187,N_10837);
nor U18607 (N_18607,N_14122,N_12704);
nand U18608 (N_18608,N_10855,N_11317);
nand U18609 (N_18609,N_12732,N_10091);
and U18610 (N_18610,N_10943,N_12871);
xor U18611 (N_18611,N_12182,N_12755);
and U18612 (N_18612,N_14336,N_13421);
and U18613 (N_18613,N_12408,N_12052);
nand U18614 (N_18614,N_13131,N_12813);
and U18615 (N_18615,N_12575,N_14349);
or U18616 (N_18616,N_14994,N_11404);
nor U18617 (N_18617,N_10945,N_11286);
and U18618 (N_18618,N_10374,N_13659);
nand U18619 (N_18619,N_12747,N_12714);
nand U18620 (N_18620,N_13291,N_10656);
nand U18621 (N_18621,N_14985,N_14402);
nor U18622 (N_18622,N_11577,N_11728);
and U18623 (N_18623,N_14883,N_14429);
xnor U18624 (N_18624,N_14657,N_10168);
or U18625 (N_18625,N_14630,N_14465);
nor U18626 (N_18626,N_12194,N_14126);
or U18627 (N_18627,N_14783,N_14885);
or U18628 (N_18628,N_14950,N_14685);
or U18629 (N_18629,N_11306,N_13492);
nor U18630 (N_18630,N_14522,N_12506);
nor U18631 (N_18631,N_13350,N_11218);
nand U18632 (N_18632,N_12193,N_11805);
nand U18633 (N_18633,N_10251,N_13190);
nor U18634 (N_18634,N_14671,N_13003);
nand U18635 (N_18635,N_11115,N_14529);
nand U18636 (N_18636,N_10167,N_13980);
or U18637 (N_18637,N_13982,N_13605);
xor U18638 (N_18638,N_12565,N_11877);
nand U18639 (N_18639,N_10644,N_12501);
nand U18640 (N_18640,N_14748,N_13209);
nand U18641 (N_18641,N_10112,N_14185);
or U18642 (N_18642,N_11942,N_14241);
nor U18643 (N_18643,N_14271,N_13489);
nor U18644 (N_18644,N_13516,N_12383);
xor U18645 (N_18645,N_13958,N_12535);
nor U18646 (N_18646,N_10589,N_13725);
xnor U18647 (N_18647,N_10511,N_14750);
and U18648 (N_18648,N_13065,N_10512);
nand U18649 (N_18649,N_13395,N_13606);
or U18650 (N_18650,N_12717,N_13773);
nand U18651 (N_18651,N_13278,N_11236);
nor U18652 (N_18652,N_13833,N_12003);
xor U18653 (N_18653,N_10839,N_11070);
xnor U18654 (N_18654,N_14531,N_11036);
and U18655 (N_18655,N_13924,N_11213);
nor U18656 (N_18656,N_14741,N_11318);
nand U18657 (N_18657,N_11086,N_10848);
and U18658 (N_18658,N_13455,N_11517);
nand U18659 (N_18659,N_14023,N_10071);
or U18660 (N_18660,N_12831,N_12069);
or U18661 (N_18661,N_13820,N_12793);
nand U18662 (N_18662,N_14275,N_11917);
nor U18663 (N_18663,N_10652,N_11853);
nand U18664 (N_18664,N_11169,N_11304);
nor U18665 (N_18665,N_14620,N_10098);
and U18666 (N_18666,N_14710,N_14326);
nor U18667 (N_18667,N_13967,N_14925);
and U18668 (N_18668,N_10873,N_13424);
nor U18669 (N_18669,N_11547,N_11022);
or U18670 (N_18670,N_13108,N_11372);
nand U18671 (N_18671,N_13233,N_11760);
and U18672 (N_18672,N_10140,N_13178);
nor U18673 (N_18673,N_11142,N_12166);
nor U18674 (N_18674,N_10451,N_14553);
nor U18675 (N_18675,N_11305,N_12232);
nor U18676 (N_18676,N_11183,N_14392);
nand U18677 (N_18677,N_11452,N_10864);
nand U18678 (N_18678,N_14377,N_13984);
and U18679 (N_18679,N_14668,N_14591);
nand U18680 (N_18680,N_14210,N_12736);
nand U18681 (N_18681,N_14965,N_10614);
or U18682 (N_18682,N_10915,N_11866);
nand U18683 (N_18683,N_11648,N_10491);
nor U18684 (N_18684,N_14122,N_12979);
nor U18685 (N_18685,N_14263,N_12973);
xnor U18686 (N_18686,N_13935,N_12174);
and U18687 (N_18687,N_10231,N_12823);
nand U18688 (N_18688,N_13382,N_11521);
nand U18689 (N_18689,N_14626,N_11359);
and U18690 (N_18690,N_13906,N_10965);
nor U18691 (N_18691,N_10622,N_10821);
nor U18692 (N_18692,N_13310,N_14123);
nand U18693 (N_18693,N_11612,N_11792);
xor U18694 (N_18694,N_13209,N_11399);
or U18695 (N_18695,N_13473,N_13459);
nand U18696 (N_18696,N_10519,N_14511);
and U18697 (N_18697,N_12007,N_14907);
and U18698 (N_18698,N_12671,N_11600);
and U18699 (N_18699,N_14964,N_10171);
nor U18700 (N_18700,N_10200,N_10008);
nand U18701 (N_18701,N_11186,N_10632);
nand U18702 (N_18702,N_11605,N_12021);
xor U18703 (N_18703,N_13226,N_13723);
or U18704 (N_18704,N_13898,N_11320);
or U18705 (N_18705,N_12275,N_10749);
or U18706 (N_18706,N_10700,N_11977);
nand U18707 (N_18707,N_11052,N_11653);
or U18708 (N_18708,N_11128,N_12166);
or U18709 (N_18709,N_10062,N_14200);
nand U18710 (N_18710,N_14642,N_13611);
nor U18711 (N_18711,N_12591,N_11410);
and U18712 (N_18712,N_11432,N_13113);
nand U18713 (N_18713,N_11764,N_12915);
nand U18714 (N_18714,N_14624,N_13487);
and U18715 (N_18715,N_14796,N_12966);
nor U18716 (N_18716,N_13458,N_14546);
or U18717 (N_18717,N_10689,N_14091);
or U18718 (N_18718,N_13370,N_10181);
and U18719 (N_18719,N_11866,N_13943);
and U18720 (N_18720,N_14306,N_10526);
or U18721 (N_18721,N_11032,N_13009);
nor U18722 (N_18722,N_10894,N_10611);
or U18723 (N_18723,N_10064,N_10877);
xnor U18724 (N_18724,N_13309,N_14971);
nor U18725 (N_18725,N_12027,N_14271);
nand U18726 (N_18726,N_10543,N_14468);
and U18727 (N_18727,N_12700,N_12229);
and U18728 (N_18728,N_11805,N_13740);
and U18729 (N_18729,N_10410,N_14238);
and U18730 (N_18730,N_11265,N_11418);
or U18731 (N_18731,N_11298,N_11666);
nor U18732 (N_18732,N_14058,N_12603);
or U18733 (N_18733,N_10216,N_11680);
nand U18734 (N_18734,N_10448,N_14171);
or U18735 (N_18735,N_14499,N_12345);
or U18736 (N_18736,N_11854,N_12946);
and U18737 (N_18737,N_13362,N_12033);
nand U18738 (N_18738,N_12125,N_14697);
or U18739 (N_18739,N_13142,N_12513);
nand U18740 (N_18740,N_13257,N_13409);
nor U18741 (N_18741,N_14566,N_11569);
nand U18742 (N_18742,N_11169,N_13924);
nand U18743 (N_18743,N_14714,N_12414);
nor U18744 (N_18744,N_10011,N_12250);
and U18745 (N_18745,N_14749,N_13149);
xnor U18746 (N_18746,N_14644,N_14054);
nand U18747 (N_18747,N_13351,N_14509);
nand U18748 (N_18748,N_13479,N_14077);
nand U18749 (N_18749,N_14965,N_10543);
nand U18750 (N_18750,N_10417,N_10267);
and U18751 (N_18751,N_14126,N_14538);
nand U18752 (N_18752,N_14174,N_14138);
nor U18753 (N_18753,N_10216,N_14932);
or U18754 (N_18754,N_14934,N_12665);
xnor U18755 (N_18755,N_14605,N_11069);
and U18756 (N_18756,N_14229,N_13219);
nor U18757 (N_18757,N_13346,N_10704);
xor U18758 (N_18758,N_14374,N_14493);
or U18759 (N_18759,N_14083,N_13241);
nor U18760 (N_18760,N_12709,N_13508);
nand U18761 (N_18761,N_11874,N_12976);
xnor U18762 (N_18762,N_14830,N_12026);
nand U18763 (N_18763,N_11415,N_14370);
and U18764 (N_18764,N_14466,N_12448);
and U18765 (N_18765,N_13993,N_11057);
nand U18766 (N_18766,N_13847,N_11424);
or U18767 (N_18767,N_14356,N_13654);
nand U18768 (N_18768,N_12181,N_14351);
nor U18769 (N_18769,N_12565,N_13570);
nand U18770 (N_18770,N_14028,N_14191);
nor U18771 (N_18771,N_10163,N_14851);
or U18772 (N_18772,N_11570,N_13828);
and U18773 (N_18773,N_11281,N_13474);
or U18774 (N_18774,N_10509,N_11719);
xor U18775 (N_18775,N_14219,N_12425);
nor U18776 (N_18776,N_10900,N_14131);
nor U18777 (N_18777,N_11226,N_14736);
or U18778 (N_18778,N_14107,N_13741);
nor U18779 (N_18779,N_12051,N_10482);
nor U18780 (N_18780,N_13168,N_14172);
xnor U18781 (N_18781,N_10180,N_11965);
nor U18782 (N_18782,N_13661,N_13409);
or U18783 (N_18783,N_10219,N_11956);
or U18784 (N_18784,N_10306,N_11603);
or U18785 (N_18785,N_12898,N_11261);
xnor U18786 (N_18786,N_13652,N_11869);
nand U18787 (N_18787,N_11368,N_13172);
nand U18788 (N_18788,N_10783,N_14455);
nor U18789 (N_18789,N_12543,N_14653);
xor U18790 (N_18790,N_10755,N_14809);
nor U18791 (N_18791,N_14999,N_12543);
nand U18792 (N_18792,N_11259,N_13399);
nor U18793 (N_18793,N_13367,N_13889);
nor U18794 (N_18794,N_13230,N_11323);
nor U18795 (N_18795,N_10221,N_13459);
or U18796 (N_18796,N_10156,N_12592);
or U18797 (N_18797,N_10714,N_13144);
and U18798 (N_18798,N_11068,N_10467);
and U18799 (N_18799,N_13972,N_13675);
nand U18800 (N_18800,N_13399,N_14538);
nand U18801 (N_18801,N_12917,N_14663);
or U18802 (N_18802,N_11519,N_10300);
or U18803 (N_18803,N_13432,N_10888);
nand U18804 (N_18804,N_12283,N_11499);
nor U18805 (N_18805,N_12615,N_13689);
nor U18806 (N_18806,N_10643,N_10517);
nand U18807 (N_18807,N_10422,N_13127);
or U18808 (N_18808,N_13454,N_10324);
and U18809 (N_18809,N_11880,N_12934);
xnor U18810 (N_18810,N_14742,N_10771);
nor U18811 (N_18811,N_11804,N_10794);
nand U18812 (N_18812,N_11417,N_11984);
or U18813 (N_18813,N_10009,N_14373);
nand U18814 (N_18814,N_13056,N_13076);
and U18815 (N_18815,N_10602,N_12957);
or U18816 (N_18816,N_12298,N_10718);
xnor U18817 (N_18817,N_14294,N_14461);
and U18818 (N_18818,N_12809,N_10423);
and U18819 (N_18819,N_10820,N_13139);
nor U18820 (N_18820,N_10150,N_14980);
nand U18821 (N_18821,N_13766,N_13722);
xor U18822 (N_18822,N_14977,N_11688);
and U18823 (N_18823,N_10538,N_13706);
or U18824 (N_18824,N_10604,N_10310);
or U18825 (N_18825,N_13649,N_10162);
xor U18826 (N_18826,N_14878,N_11084);
nand U18827 (N_18827,N_11261,N_10793);
and U18828 (N_18828,N_12112,N_13170);
nor U18829 (N_18829,N_13640,N_12008);
or U18830 (N_18830,N_14367,N_11328);
or U18831 (N_18831,N_11379,N_12240);
or U18832 (N_18832,N_12475,N_13479);
xnor U18833 (N_18833,N_13877,N_12812);
nand U18834 (N_18834,N_11002,N_11519);
nand U18835 (N_18835,N_13070,N_10959);
nand U18836 (N_18836,N_11775,N_14630);
or U18837 (N_18837,N_14897,N_10947);
or U18838 (N_18838,N_14711,N_10706);
nand U18839 (N_18839,N_10029,N_12759);
nor U18840 (N_18840,N_11927,N_14138);
and U18841 (N_18841,N_10466,N_10963);
and U18842 (N_18842,N_10359,N_10331);
nand U18843 (N_18843,N_12939,N_10593);
nand U18844 (N_18844,N_13634,N_14375);
nand U18845 (N_18845,N_10224,N_11493);
and U18846 (N_18846,N_14687,N_13019);
and U18847 (N_18847,N_13299,N_12894);
nor U18848 (N_18848,N_13332,N_13617);
nor U18849 (N_18849,N_12262,N_12598);
nor U18850 (N_18850,N_12014,N_13607);
and U18851 (N_18851,N_12692,N_12103);
or U18852 (N_18852,N_14371,N_14700);
nand U18853 (N_18853,N_12260,N_12116);
and U18854 (N_18854,N_12612,N_11751);
nand U18855 (N_18855,N_10633,N_13170);
or U18856 (N_18856,N_13349,N_14426);
nand U18857 (N_18857,N_10751,N_14760);
and U18858 (N_18858,N_11403,N_11131);
or U18859 (N_18859,N_12515,N_13893);
nand U18860 (N_18860,N_10434,N_13346);
and U18861 (N_18861,N_13750,N_10463);
and U18862 (N_18862,N_11225,N_10250);
and U18863 (N_18863,N_12356,N_12668);
and U18864 (N_18864,N_12782,N_12428);
nor U18865 (N_18865,N_11498,N_10842);
nand U18866 (N_18866,N_11025,N_12058);
nor U18867 (N_18867,N_12867,N_14115);
nand U18868 (N_18868,N_12583,N_11796);
xor U18869 (N_18869,N_10243,N_10054);
or U18870 (N_18870,N_13011,N_10537);
nor U18871 (N_18871,N_11097,N_14213);
and U18872 (N_18872,N_12043,N_14920);
and U18873 (N_18873,N_12344,N_10793);
and U18874 (N_18874,N_10024,N_14269);
and U18875 (N_18875,N_11102,N_14337);
and U18876 (N_18876,N_13193,N_10968);
xnor U18877 (N_18877,N_11938,N_11662);
xor U18878 (N_18878,N_11223,N_13631);
or U18879 (N_18879,N_10507,N_10345);
and U18880 (N_18880,N_12942,N_12407);
or U18881 (N_18881,N_10694,N_14902);
xor U18882 (N_18882,N_10830,N_11807);
nor U18883 (N_18883,N_14537,N_12826);
nand U18884 (N_18884,N_14784,N_14628);
nor U18885 (N_18885,N_12147,N_14591);
or U18886 (N_18886,N_13902,N_11246);
or U18887 (N_18887,N_13185,N_14009);
nor U18888 (N_18888,N_14646,N_10215);
xor U18889 (N_18889,N_10923,N_10358);
or U18890 (N_18890,N_10394,N_13928);
or U18891 (N_18891,N_11983,N_13112);
or U18892 (N_18892,N_14072,N_14363);
or U18893 (N_18893,N_10071,N_10624);
and U18894 (N_18894,N_11282,N_12604);
or U18895 (N_18895,N_11555,N_12049);
and U18896 (N_18896,N_13407,N_14801);
nor U18897 (N_18897,N_13003,N_13841);
nand U18898 (N_18898,N_14717,N_11718);
or U18899 (N_18899,N_12576,N_11521);
nand U18900 (N_18900,N_14047,N_11144);
nand U18901 (N_18901,N_11802,N_11473);
and U18902 (N_18902,N_12753,N_11956);
or U18903 (N_18903,N_13786,N_10000);
nand U18904 (N_18904,N_13938,N_13608);
or U18905 (N_18905,N_10197,N_14869);
and U18906 (N_18906,N_12998,N_11048);
or U18907 (N_18907,N_11564,N_14427);
or U18908 (N_18908,N_13711,N_14726);
nand U18909 (N_18909,N_12431,N_10401);
nand U18910 (N_18910,N_12030,N_12756);
nor U18911 (N_18911,N_14219,N_11129);
or U18912 (N_18912,N_10057,N_14041);
or U18913 (N_18913,N_12994,N_13504);
nand U18914 (N_18914,N_11015,N_13451);
or U18915 (N_18915,N_11590,N_11850);
nand U18916 (N_18916,N_13308,N_10532);
or U18917 (N_18917,N_12145,N_11255);
or U18918 (N_18918,N_11788,N_13262);
xnor U18919 (N_18919,N_10987,N_11100);
nor U18920 (N_18920,N_12070,N_12190);
nor U18921 (N_18921,N_10741,N_12371);
and U18922 (N_18922,N_11839,N_14639);
and U18923 (N_18923,N_13713,N_12626);
and U18924 (N_18924,N_14155,N_10807);
nand U18925 (N_18925,N_11830,N_10899);
or U18926 (N_18926,N_10349,N_14286);
and U18927 (N_18927,N_13731,N_14040);
nand U18928 (N_18928,N_11485,N_14438);
or U18929 (N_18929,N_12750,N_14379);
nand U18930 (N_18930,N_10552,N_10029);
and U18931 (N_18931,N_11427,N_10973);
and U18932 (N_18932,N_14999,N_12220);
xor U18933 (N_18933,N_11280,N_11140);
nand U18934 (N_18934,N_11969,N_11650);
and U18935 (N_18935,N_13768,N_11608);
and U18936 (N_18936,N_12552,N_13280);
nand U18937 (N_18937,N_12677,N_10840);
nor U18938 (N_18938,N_11681,N_14089);
xnor U18939 (N_18939,N_10134,N_13394);
or U18940 (N_18940,N_12560,N_14011);
or U18941 (N_18941,N_14636,N_14549);
nor U18942 (N_18942,N_14833,N_14355);
nor U18943 (N_18943,N_10367,N_10929);
and U18944 (N_18944,N_12057,N_12905);
nand U18945 (N_18945,N_12928,N_10663);
and U18946 (N_18946,N_12256,N_11231);
nand U18947 (N_18947,N_11209,N_10383);
or U18948 (N_18948,N_13407,N_11069);
nand U18949 (N_18949,N_11978,N_11780);
nor U18950 (N_18950,N_10925,N_10176);
nand U18951 (N_18951,N_10386,N_11104);
and U18952 (N_18952,N_13018,N_12702);
and U18953 (N_18953,N_10305,N_12543);
nor U18954 (N_18954,N_10058,N_13065);
nor U18955 (N_18955,N_13400,N_13024);
or U18956 (N_18956,N_12632,N_11506);
nor U18957 (N_18957,N_12935,N_11728);
nand U18958 (N_18958,N_13195,N_10785);
xnor U18959 (N_18959,N_14499,N_11422);
nand U18960 (N_18960,N_12544,N_10907);
and U18961 (N_18961,N_14987,N_13242);
and U18962 (N_18962,N_13622,N_13055);
or U18963 (N_18963,N_13495,N_11781);
xor U18964 (N_18964,N_10236,N_14508);
nand U18965 (N_18965,N_10836,N_11002);
nand U18966 (N_18966,N_11411,N_11717);
and U18967 (N_18967,N_13219,N_11335);
nor U18968 (N_18968,N_14413,N_13299);
nand U18969 (N_18969,N_12416,N_14487);
nor U18970 (N_18970,N_12214,N_13197);
nor U18971 (N_18971,N_14482,N_12501);
nand U18972 (N_18972,N_13499,N_10823);
or U18973 (N_18973,N_11681,N_13800);
or U18974 (N_18974,N_11829,N_13659);
and U18975 (N_18975,N_14196,N_13913);
nand U18976 (N_18976,N_10393,N_12236);
nor U18977 (N_18977,N_11663,N_10941);
nand U18978 (N_18978,N_14375,N_10187);
nand U18979 (N_18979,N_11307,N_11338);
nor U18980 (N_18980,N_11018,N_14499);
or U18981 (N_18981,N_13850,N_14151);
or U18982 (N_18982,N_13008,N_10516);
nand U18983 (N_18983,N_12748,N_12888);
nor U18984 (N_18984,N_13049,N_14270);
or U18985 (N_18985,N_12460,N_12219);
nand U18986 (N_18986,N_14658,N_10008);
nor U18987 (N_18987,N_14231,N_10217);
or U18988 (N_18988,N_10085,N_13142);
or U18989 (N_18989,N_13648,N_14014);
nand U18990 (N_18990,N_13711,N_14456);
or U18991 (N_18991,N_14932,N_14294);
nand U18992 (N_18992,N_12076,N_10751);
nor U18993 (N_18993,N_11256,N_12890);
nor U18994 (N_18994,N_13973,N_13467);
or U18995 (N_18995,N_12815,N_12434);
xor U18996 (N_18996,N_13454,N_14303);
nand U18997 (N_18997,N_12424,N_11411);
and U18998 (N_18998,N_14554,N_14482);
nand U18999 (N_18999,N_11954,N_12940);
and U19000 (N_19000,N_13196,N_12544);
or U19001 (N_19001,N_10707,N_11783);
xor U19002 (N_19002,N_10909,N_12863);
and U19003 (N_19003,N_12903,N_12770);
nor U19004 (N_19004,N_13805,N_12265);
nand U19005 (N_19005,N_13251,N_12057);
nand U19006 (N_19006,N_14245,N_11655);
xnor U19007 (N_19007,N_13301,N_10865);
and U19008 (N_19008,N_10590,N_11977);
and U19009 (N_19009,N_11473,N_12418);
nor U19010 (N_19010,N_11753,N_10993);
or U19011 (N_19011,N_14613,N_11476);
nor U19012 (N_19012,N_12814,N_14554);
xor U19013 (N_19013,N_11380,N_10329);
and U19014 (N_19014,N_10429,N_12752);
nand U19015 (N_19015,N_11031,N_11003);
nand U19016 (N_19016,N_10360,N_12576);
nand U19017 (N_19017,N_14758,N_11778);
and U19018 (N_19018,N_13016,N_14847);
and U19019 (N_19019,N_11110,N_11619);
and U19020 (N_19020,N_14496,N_12046);
or U19021 (N_19021,N_11165,N_11889);
and U19022 (N_19022,N_10632,N_12875);
and U19023 (N_19023,N_11075,N_10663);
or U19024 (N_19024,N_13026,N_13141);
nor U19025 (N_19025,N_10182,N_14257);
or U19026 (N_19026,N_14372,N_12549);
nor U19027 (N_19027,N_11880,N_10239);
nor U19028 (N_19028,N_10681,N_13453);
nor U19029 (N_19029,N_12196,N_11609);
and U19030 (N_19030,N_13876,N_12964);
or U19031 (N_19031,N_10172,N_11658);
nand U19032 (N_19032,N_14837,N_12856);
nand U19033 (N_19033,N_12932,N_11587);
or U19034 (N_19034,N_12816,N_12969);
and U19035 (N_19035,N_13935,N_10253);
nand U19036 (N_19036,N_10612,N_12147);
nor U19037 (N_19037,N_10620,N_12861);
nand U19038 (N_19038,N_13960,N_10456);
and U19039 (N_19039,N_13552,N_11500);
nand U19040 (N_19040,N_12555,N_12619);
or U19041 (N_19041,N_13426,N_13198);
nand U19042 (N_19042,N_13938,N_10540);
nor U19043 (N_19043,N_13418,N_10048);
nor U19044 (N_19044,N_11064,N_11491);
nand U19045 (N_19045,N_13766,N_13755);
or U19046 (N_19046,N_10040,N_10062);
and U19047 (N_19047,N_13957,N_14386);
and U19048 (N_19048,N_11464,N_12074);
or U19049 (N_19049,N_10873,N_12052);
and U19050 (N_19050,N_11185,N_10498);
nand U19051 (N_19051,N_12193,N_14841);
and U19052 (N_19052,N_13089,N_11240);
nor U19053 (N_19053,N_11592,N_14438);
xnor U19054 (N_19054,N_14166,N_11803);
nand U19055 (N_19055,N_10348,N_11172);
and U19056 (N_19056,N_11659,N_14969);
and U19057 (N_19057,N_10938,N_14277);
nand U19058 (N_19058,N_11645,N_11564);
and U19059 (N_19059,N_11102,N_11241);
xor U19060 (N_19060,N_13977,N_14300);
nand U19061 (N_19061,N_10649,N_13162);
nand U19062 (N_19062,N_10187,N_10900);
nor U19063 (N_19063,N_10132,N_12016);
and U19064 (N_19064,N_10050,N_11752);
nor U19065 (N_19065,N_14356,N_11295);
or U19066 (N_19066,N_10071,N_10713);
nor U19067 (N_19067,N_11309,N_11676);
or U19068 (N_19068,N_10973,N_12852);
or U19069 (N_19069,N_13642,N_12138);
and U19070 (N_19070,N_13226,N_14166);
and U19071 (N_19071,N_14699,N_12909);
nor U19072 (N_19072,N_14391,N_10538);
nand U19073 (N_19073,N_14677,N_12700);
and U19074 (N_19074,N_13940,N_14175);
nand U19075 (N_19075,N_12522,N_10608);
xnor U19076 (N_19076,N_10668,N_12189);
and U19077 (N_19077,N_13160,N_13572);
xor U19078 (N_19078,N_13396,N_13290);
nor U19079 (N_19079,N_12866,N_13651);
or U19080 (N_19080,N_10441,N_14776);
nor U19081 (N_19081,N_14913,N_14969);
nand U19082 (N_19082,N_13864,N_11115);
or U19083 (N_19083,N_13410,N_11086);
or U19084 (N_19084,N_10518,N_13263);
xor U19085 (N_19085,N_11604,N_13799);
and U19086 (N_19086,N_13144,N_12552);
nand U19087 (N_19087,N_12450,N_14553);
nand U19088 (N_19088,N_11686,N_11294);
or U19089 (N_19089,N_13628,N_10393);
nor U19090 (N_19090,N_11290,N_11368);
nor U19091 (N_19091,N_12868,N_14249);
nor U19092 (N_19092,N_12120,N_14985);
or U19093 (N_19093,N_11871,N_13024);
nand U19094 (N_19094,N_11165,N_14168);
nand U19095 (N_19095,N_11424,N_11309);
or U19096 (N_19096,N_10240,N_10942);
or U19097 (N_19097,N_12723,N_13007);
and U19098 (N_19098,N_14523,N_12372);
and U19099 (N_19099,N_11143,N_13304);
and U19100 (N_19100,N_11687,N_10926);
or U19101 (N_19101,N_12915,N_10890);
or U19102 (N_19102,N_13495,N_10487);
nor U19103 (N_19103,N_10742,N_13633);
and U19104 (N_19104,N_13847,N_10624);
or U19105 (N_19105,N_14428,N_10753);
or U19106 (N_19106,N_14420,N_10567);
nand U19107 (N_19107,N_12372,N_13334);
or U19108 (N_19108,N_12179,N_13519);
nor U19109 (N_19109,N_12384,N_10765);
nand U19110 (N_19110,N_12188,N_14383);
nand U19111 (N_19111,N_14941,N_11071);
or U19112 (N_19112,N_14750,N_14957);
nor U19113 (N_19113,N_10782,N_13770);
nor U19114 (N_19114,N_13615,N_11358);
nor U19115 (N_19115,N_12415,N_12222);
and U19116 (N_19116,N_12228,N_11464);
nand U19117 (N_19117,N_14576,N_10429);
nand U19118 (N_19118,N_10400,N_13295);
nand U19119 (N_19119,N_12343,N_10873);
nor U19120 (N_19120,N_13745,N_11535);
xor U19121 (N_19121,N_13341,N_12705);
nor U19122 (N_19122,N_10683,N_11143);
or U19123 (N_19123,N_12189,N_12390);
and U19124 (N_19124,N_11073,N_12615);
nand U19125 (N_19125,N_10483,N_13389);
or U19126 (N_19126,N_10065,N_13562);
nand U19127 (N_19127,N_14347,N_14739);
or U19128 (N_19128,N_11286,N_13863);
or U19129 (N_19129,N_11585,N_10160);
xnor U19130 (N_19130,N_11888,N_14056);
and U19131 (N_19131,N_11061,N_14342);
and U19132 (N_19132,N_10324,N_14822);
xor U19133 (N_19133,N_11434,N_11183);
and U19134 (N_19134,N_11978,N_13434);
xor U19135 (N_19135,N_11891,N_10328);
nand U19136 (N_19136,N_10155,N_12345);
nor U19137 (N_19137,N_12132,N_14579);
or U19138 (N_19138,N_14330,N_10439);
or U19139 (N_19139,N_10518,N_11889);
nor U19140 (N_19140,N_13803,N_13076);
nor U19141 (N_19141,N_10345,N_12372);
and U19142 (N_19142,N_11195,N_11553);
nor U19143 (N_19143,N_14108,N_12652);
nand U19144 (N_19144,N_10951,N_10487);
and U19145 (N_19145,N_12111,N_12603);
nand U19146 (N_19146,N_12002,N_10284);
and U19147 (N_19147,N_14142,N_14114);
nand U19148 (N_19148,N_14345,N_14086);
nor U19149 (N_19149,N_12631,N_14772);
and U19150 (N_19150,N_11891,N_11775);
nand U19151 (N_19151,N_13120,N_10996);
or U19152 (N_19152,N_10953,N_12619);
xor U19153 (N_19153,N_12023,N_14627);
xnor U19154 (N_19154,N_11201,N_12528);
xor U19155 (N_19155,N_11846,N_14441);
nor U19156 (N_19156,N_14651,N_13243);
nand U19157 (N_19157,N_11671,N_10800);
or U19158 (N_19158,N_13191,N_12402);
and U19159 (N_19159,N_12893,N_11096);
xor U19160 (N_19160,N_12283,N_14501);
and U19161 (N_19161,N_11478,N_11584);
and U19162 (N_19162,N_10981,N_13508);
nand U19163 (N_19163,N_11586,N_14305);
nor U19164 (N_19164,N_13140,N_13554);
xnor U19165 (N_19165,N_14482,N_12208);
nor U19166 (N_19166,N_13970,N_14838);
nor U19167 (N_19167,N_14295,N_14117);
nor U19168 (N_19168,N_13719,N_11781);
and U19169 (N_19169,N_10910,N_11201);
nor U19170 (N_19170,N_14266,N_10717);
and U19171 (N_19171,N_11640,N_11054);
xor U19172 (N_19172,N_14242,N_13582);
nand U19173 (N_19173,N_11746,N_12103);
nor U19174 (N_19174,N_13828,N_14992);
nand U19175 (N_19175,N_10485,N_14931);
and U19176 (N_19176,N_14484,N_14601);
xnor U19177 (N_19177,N_14492,N_10118);
nand U19178 (N_19178,N_13207,N_14750);
xor U19179 (N_19179,N_10756,N_12246);
xnor U19180 (N_19180,N_11934,N_11384);
or U19181 (N_19181,N_13886,N_12117);
xnor U19182 (N_19182,N_10556,N_14542);
nor U19183 (N_19183,N_13255,N_12960);
nand U19184 (N_19184,N_11284,N_14184);
xnor U19185 (N_19185,N_12977,N_11191);
nor U19186 (N_19186,N_10988,N_14195);
or U19187 (N_19187,N_10222,N_14761);
and U19188 (N_19188,N_11546,N_12965);
nand U19189 (N_19189,N_11550,N_10523);
nor U19190 (N_19190,N_14444,N_10975);
nand U19191 (N_19191,N_13331,N_11390);
nand U19192 (N_19192,N_10808,N_10299);
nor U19193 (N_19193,N_13083,N_12719);
nor U19194 (N_19194,N_12478,N_12875);
or U19195 (N_19195,N_10254,N_11500);
xor U19196 (N_19196,N_10606,N_12764);
nor U19197 (N_19197,N_10121,N_12583);
nand U19198 (N_19198,N_11633,N_13055);
nand U19199 (N_19199,N_12091,N_12120);
or U19200 (N_19200,N_13638,N_14226);
nand U19201 (N_19201,N_10070,N_11768);
nand U19202 (N_19202,N_10654,N_13804);
or U19203 (N_19203,N_13772,N_11887);
and U19204 (N_19204,N_14057,N_11989);
or U19205 (N_19205,N_10590,N_12699);
xnor U19206 (N_19206,N_13906,N_10075);
and U19207 (N_19207,N_13092,N_14461);
nor U19208 (N_19208,N_10215,N_10828);
and U19209 (N_19209,N_11005,N_14099);
nor U19210 (N_19210,N_10485,N_14284);
nor U19211 (N_19211,N_12553,N_14238);
or U19212 (N_19212,N_13845,N_13249);
or U19213 (N_19213,N_11490,N_14552);
or U19214 (N_19214,N_12625,N_11832);
nand U19215 (N_19215,N_13962,N_12951);
nor U19216 (N_19216,N_11733,N_12154);
nor U19217 (N_19217,N_10784,N_12237);
and U19218 (N_19218,N_10370,N_13808);
or U19219 (N_19219,N_13026,N_11554);
nor U19220 (N_19220,N_14025,N_10702);
nand U19221 (N_19221,N_11180,N_10321);
nor U19222 (N_19222,N_10384,N_10800);
nor U19223 (N_19223,N_10295,N_10285);
xnor U19224 (N_19224,N_12967,N_11658);
or U19225 (N_19225,N_10808,N_12099);
xor U19226 (N_19226,N_14355,N_13477);
nor U19227 (N_19227,N_13867,N_14068);
and U19228 (N_19228,N_11348,N_14467);
or U19229 (N_19229,N_11814,N_11773);
nand U19230 (N_19230,N_14184,N_14146);
nand U19231 (N_19231,N_11379,N_11607);
or U19232 (N_19232,N_11666,N_12644);
and U19233 (N_19233,N_10135,N_14625);
nor U19234 (N_19234,N_13869,N_12471);
and U19235 (N_19235,N_11606,N_13803);
or U19236 (N_19236,N_13584,N_12504);
and U19237 (N_19237,N_10390,N_12284);
or U19238 (N_19238,N_10744,N_10069);
nor U19239 (N_19239,N_11954,N_11603);
and U19240 (N_19240,N_10869,N_14933);
xor U19241 (N_19241,N_12586,N_10082);
nor U19242 (N_19242,N_13263,N_12688);
nor U19243 (N_19243,N_10148,N_12083);
nand U19244 (N_19244,N_13008,N_10079);
xor U19245 (N_19245,N_14738,N_13181);
nor U19246 (N_19246,N_13862,N_10942);
nand U19247 (N_19247,N_11808,N_10288);
or U19248 (N_19248,N_13047,N_11383);
nor U19249 (N_19249,N_12782,N_14833);
and U19250 (N_19250,N_12347,N_14792);
nand U19251 (N_19251,N_12914,N_12591);
and U19252 (N_19252,N_14179,N_14096);
nand U19253 (N_19253,N_14473,N_14372);
nand U19254 (N_19254,N_10852,N_12931);
nor U19255 (N_19255,N_14159,N_11248);
and U19256 (N_19256,N_12514,N_13940);
and U19257 (N_19257,N_14275,N_12554);
nand U19258 (N_19258,N_12004,N_10158);
nor U19259 (N_19259,N_10173,N_12672);
nand U19260 (N_19260,N_12328,N_10078);
xor U19261 (N_19261,N_12372,N_14696);
or U19262 (N_19262,N_13037,N_13153);
nor U19263 (N_19263,N_11798,N_13552);
nor U19264 (N_19264,N_10431,N_12530);
and U19265 (N_19265,N_10638,N_13058);
and U19266 (N_19266,N_11668,N_14148);
or U19267 (N_19267,N_14103,N_11843);
nand U19268 (N_19268,N_12057,N_14258);
and U19269 (N_19269,N_11122,N_10553);
nand U19270 (N_19270,N_11139,N_10127);
nand U19271 (N_19271,N_13174,N_11600);
nor U19272 (N_19272,N_12956,N_10038);
xor U19273 (N_19273,N_14776,N_12559);
and U19274 (N_19274,N_11482,N_14773);
nor U19275 (N_19275,N_11838,N_11312);
nor U19276 (N_19276,N_11766,N_14296);
and U19277 (N_19277,N_11918,N_11656);
or U19278 (N_19278,N_12365,N_10495);
nor U19279 (N_19279,N_11844,N_12045);
and U19280 (N_19280,N_10785,N_11601);
or U19281 (N_19281,N_13568,N_10659);
or U19282 (N_19282,N_10909,N_14846);
and U19283 (N_19283,N_12095,N_12487);
and U19284 (N_19284,N_14928,N_13063);
nand U19285 (N_19285,N_11492,N_13775);
nand U19286 (N_19286,N_12240,N_14120);
or U19287 (N_19287,N_12428,N_12450);
or U19288 (N_19288,N_14425,N_14256);
and U19289 (N_19289,N_11850,N_14997);
nor U19290 (N_19290,N_11248,N_11107);
and U19291 (N_19291,N_12221,N_10907);
and U19292 (N_19292,N_14000,N_11974);
or U19293 (N_19293,N_14144,N_12799);
and U19294 (N_19294,N_14450,N_12378);
xor U19295 (N_19295,N_13857,N_10575);
and U19296 (N_19296,N_13044,N_14956);
nand U19297 (N_19297,N_14400,N_10261);
and U19298 (N_19298,N_10494,N_12025);
and U19299 (N_19299,N_14609,N_10372);
or U19300 (N_19300,N_14565,N_12231);
nor U19301 (N_19301,N_13821,N_12551);
or U19302 (N_19302,N_11498,N_10604);
nand U19303 (N_19303,N_14102,N_11482);
nor U19304 (N_19304,N_11112,N_11874);
nand U19305 (N_19305,N_10089,N_12478);
and U19306 (N_19306,N_13936,N_14538);
nand U19307 (N_19307,N_14234,N_13457);
or U19308 (N_19308,N_12715,N_14720);
nand U19309 (N_19309,N_11524,N_10415);
nand U19310 (N_19310,N_10580,N_14073);
nand U19311 (N_19311,N_10240,N_11308);
xor U19312 (N_19312,N_14400,N_12423);
xor U19313 (N_19313,N_11706,N_11247);
nand U19314 (N_19314,N_14016,N_10342);
nor U19315 (N_19315,N_14910,N_10795);
or U19316 (N_19316,N_10750,N_11731);
or U19317 (N_19317,N_13450,N_12008);
and U19318 (N_19318,N_10171,N_10851);
nand U19319 (N_19319,N_11566,N_14421);
and U19320 (N_19320,N_11933,N_10652);
xnor U19321 (N_19321,N_12015,N_14981);
and U19322 (N_19322,N_14303,N_10201);
nor U19323 (N_19323,N_11179,N_14453);
xnor U19324 (N_19324,N_13079,N_11383);
nor U19325 (N_19325,N_13691,N_12550);
nand U19326 (N_19326,N_10216,N_11573);
nor U19327 (N_19327,N_14506,N_13549);
nand U19328 (N_19328,N_11689,N_14503);
nand U19329 (N_19329,N_11526,N_14922);
or U19330 (N_19330,N_12024,N_12124);
or U19331 (N_19331,N_14613,N_12350);
xor U19332 (N_19332,N_12360,N_11125);
and U19333 (N_19333,N_13918,N_10992);
nand U19334 (N_19334,N_10150,N_10965);
nand U19335 (N_19335,N_14857,N_12808);
nor U19336 (N_19336,N_10693,N_14039);
or U19337 (N_19337,N_10860,N_12525);
or U19338 (N_19338,N_14289,N_13092);
or U19339 (N_19339,N_10421,N_11134);
nand U19340 (N_19340,N_14823,N_14539);
and U19341 (N_19341,N_11230,N_13571);
xor U19342 (N_19342,N_11238,N_10566);
nor U19343 (N_19343,N_11492,N_12905);
xnor U19344 (N_19344,N_11798,N_10574);
nor U19345 (N_19345,N_10995,N_12498);
nor U19346 (N_19346,N_12106,N_14324);
or U19347 (N_19347,N_14801,N_14617);
nor U19348 (N_19348,N_12937,N_10491);
xnor U19349 (N_19349,N_11681,N_13727);
nand U19350 (N_19350,N_10453,N_12164);
and U19351 (N_19351,N_14900,N_13668);
and U19352 (N_19352,N_14381,N_12138);
or U19353 (N_19353,N_14950,N_10147);
nor U19354 (N_19354,N_14965,N_14857);
nor U19355 (N_19355,N_13631,N_13765);
nor U19356 (N_19356,N_11910,N_13420);
nor U19357 (N_19357,N_11686,N_14728);
xnor U19358 (N_19358,N_14854,N_10441);
xnor U19359 (N_19359,N_11704,N_10672);
nor U19360 (N_19360,N_10113,N_14946);
and U19361 (N_19361,N_14490,N_11205);
nand U19362 (N_19362,N_11598,N_14891);
nand U19363 (N_19363,N_10630,N_11095);
and U19364 (N_19364,N_11163,N_10828);
or U19365 (N_19365,N_12255,N_12278);
or U19366 (N_19366,N_10263,N_10487);
and U19367 (N_19367,N_11970,N_13084);
xnor U19368 (N_19368,N_11705,N_10265);
or U19369 (N_19369,N_12459,N_11526);
and U19370 (N_19370,N_12204,N_13530);
or U19371 (N_19371,N_10227,N_14624);
nor U19372 (N_19372,N_11049,N_14623);
or U19373 (N_19373,N_14087,N_14302);
and U19374 (N_19374,N_13328,N_12834);
nand U19375 (N_19375,N_13344,N_14615);
nand U19376 (N_19376,N_13215,N_13002);
nor U19377 (N_19377,N_10334,N_11494);
and U19378 (N_19378,N_11866,N_12142);
and U19379 (N_19379,N_10425,N_11767);
or U19380 (N_19380,N_10912,N_10204);
nand U19381 (N_19381,N_13537,N_10823);
nor U19382 (N_19382,N_11829,N_14193);
or U19383 (N_19383,N_10492,N_10768);
nand U19384 (N_19384,N_10994,N_14386);
or U19385 (N_19385,N_14625,N_12196);
nand U19386 (N_19386,N_13504,N_14424);
nor U19387 (N_19387,N_12746,N_14054);
nor U19388 (N_19388,N_13178,N_13780);
nor U19389 (N_19389,N_11684,N_10905);
nand U19390 (N_19390,N_11388,N_14370);
or U19391 (N_19391,N_12894,N_10445);
or U19392 (N_19392,N_13171,N_14949);
nand U19393 (N_19393,N_14910,N_12726);
or U19394 (N_19394,N_12421,N_13674);
or U19395 (N_19395,N_13160,N_10181);
nand U19396 (N_19396,N_12176,N_11305);
nor U19397 (N_19397,N_13392,N_14373);
nand U19398 (N_19398,N_14978,N_14482);
nor U19399 (N_19399,N_10603,N_12767);
or U19400 (N_19400,N_11000,N_14156);
nand U19401 (N_19401,N_13838,N_12378);
or U19402 (N_19402,N_13397,N_11627);
or U19403 (N_19403,N_10019,N_10616);
nand U19404 (N_19404,N_14074,N_14507);
or U19405 (N_19405,N_13516,N_11337);
nand U19406 (N_19406,N_13906,N_12299);
or U19407 (N_19407,N_11577,N_13928);
and U19408 (N_19408,N_11789,N_12422);
nor U19409 (N_19409,N_11668,N_10002);
nand U19410 (N_19410,N_12632,N_12253);
nor U19411 (N_19411,N_10333,N_13174);
nand U19412 (N_19412,N_13438,N_11111);
and U19413 (N_19413,N_14529,N_10897);
nand U19414 (N_19414,N_14533,N_14858);
xor U19415 (N_19415,N_10499,N_11415);
nor U19416 (N_19416,N_11457,N_13363);
and U19417 (N_19417,N_12493,N_13025);
nand U19418 (N_19418,N_12147,N_13444);
nor U19419 (N_19419,N_14245,N_13327);
nand U19420 (N_19420,N_14131,N_10234);
and U19421 (N_19421,N_13568,N_11949);
and U19422 (N_19422,N_13559,N_13079);
or U19423 (N_19423,N_13399,N_14371);
nand U19424 (N_19424,N_12972,N_12871);
nand U19425 (N_19425,N_11270,N_13695);
and U19426 (N_19426,N_14492,N_10340);
nand U19427 (N_19427,N_14337,N_14070);
and U19428 (N_19428,N_13957,N_12355);
nand U19429 (N_19429,N_14557,N_11955);
nand U19430 (N_19430,N_10154,N_11414);
nor U19431 (N_19431,N_11374,N_12994);
nand U19432 (N_19432,N_12813,N_11462);
or U19433 (N_19433,N_14957,N_12705);
or U19434 (N_19434,N_10251,N_13157);
or U19435 (N_19435,N_14007,N_14958);
and U19436 (N_19436,N_14790,N_11370);
nor U19437 (N_19437,N_14786,N_13524);
and U19438 (N_19438,N_14842,N_11046);
nor U19439 (N_19439,N_13346,N_13787);
nor U19440 (N_19440,N_14563,N_11853);
xor U19441 (N_19441,N_12396,N_10611);
nor U19442 (N_19442,N_10026,N_10590);
and U19443 (N_19443,N_11031,N_11673);
or U19444 (N_19444,N_13520,N_12435);
nor U19445 (N_19445,N_13045,N_11954);
and U19446 (N_19446,N_12315,N_14063);
nor U19447 (N_19447,N_14644,N_14499);
nor U19448 (N_19448,N_11779,N_10338);
nand U19449 (N_19449,N_11352,N_12669);
xnor U19450 (N_19450,N_12494,N_12193);
or U19451 (N_19451,N_12486,N_11070);
and U19452 (N_19452,N_14780,N_10790);
xor U19453 (N_19453,N_14910,N_10517);
nand U19454 (N_19454,N_11933,N_14922);
and U19455 (N_19455,N_13777,N_11424);
nor U19456 (N_19456,N_12724,N_10262);
nand U19457 (N_19457,N_10262,N_10232);
nor U19458 (N_19458,N_12589,N_11219);
xor U19459 (N_19459,N_13066,N_13971);
nand U19460 (N_19460,N_14641,N_11703);
or U19461 (N_19461,N_12154,N_11715);
nand U19462 (N_19462,N_11937,N_12636);
nand U19463 (N_19463,N_12924,N_11672);
nor U19464 (N_19464,N_12552,N_14199);
or U19465 (N_19465,N_13345,N_13489);
nand U19466 (N_19466,N_14001,N_13460);
or U19467 (N_19467,N_12819,N_13282);
nand U19468 (N_19468,N_12601,N_13800);
nand U19469 (N_19469,N_11753,N_13934);
and U19470 (N_19470,N_14113,N_11007);
nand U19471 (N_19471,N_10539,N_10115);
nor U19472 (N_19472,N_13870,N_13681);
nor U19473 (N_19473,N_11062,N_14969);
and U19474 (N_19474,N_12576,N_14615);
nand U19475 (N_19475,N_10887,N_11321);
nand U19476 (N_19476,N_13852,N_10380);
or U19477 (N_19477,N_14462,N_12407);
nand U19478 (N_19478,N_12450,N_14718);
or U19479 (N_19479,N_10866,N_14666);
nand U19480 (N_19480,N_10367,N_10228);
nor U19481 (N_19481,N_10344,N_10335);
nand U19482 (N_19482,N_14522,N_12848);
or U19483 (N_19483,N_12874,N_11024);
nor U19484 (N_19484,N_11354,N_13812);
xnor U19485 (N_19485,N_14022,N_13355);
nor U19486 (N_19486,N_12868,N_14640);
xor U19487 (N_19487,N_12765,N_14719);
nor U19488 (N_19488,N_14312,N_12504);
nor U19489 (N_19489,N_14474,N_13264);
nor U19490 (N_19490,N_13015,N_12382);
and U19491 (N_19491,N_11444,N_11433);
nor U19492 (N_19492,N_14800,N_11016);
nand U19493 (N_19493,N_10812,N_10214);
nand U19494 (N_19494,N_12999,N_14268);
nand U19495 (N_19495,N_11253,N_12810);
nor U19496 (N_19496,N_14294,N_13324);
xor U19497 (N_19497,N_10007,N_12587);
nor U19498 (N_19498,N_13087,N_14857);
or U19499 (N_19499,N_13757,N_13726);
nor U19500 (N_19500,N_14227,N_11579);
nand U19501 (N_19501,N_11229,N_10066);
nor U19502 (N_19502,N_11928,N_12115);
nand U19503 (N_19503,N_11289,N_12053);
nor U19504 (N_19504,N_11106,N_12602);
or U19505 (N_19505,N_14960,N_14864);
nand U19506 (N_19506,N_14617,N_13638);
nor U19507 (N_19507,N_13683,N_10024);
nor U19508 (N_19508,N_10802,N_10653);
nor U19509 (N_19509,N_12043,N_13602);
and U19510 (N_19510,N_14218,N_14175);
xnor U19511 (N_19511,N_13040,N_11352);
and U19512 (N_19512,N_10555,N_12168);
nor U19513 (N_19513,N_12718,N_12295);
nor U19514 (N_19514,N_10503,N_11931);
nand U19515 (N_19515,N_12448,N_13365);
nand U19516 (N_19516,N_14230,N_11500);
or U19517 (N_19517,N_12483,N_12653);
and U19518 (N_19518,N_10922,N_10766);
or U19519 (N_19519,N_13243,N_10293);
nand U19520 (N_19520,N_11049,N_10288);
and U19521 (N_19521,N_11011,N_12423);
nor U19522 (N_19522,N_10555,N_10954);
and U19523 (N_19523,N_11631,N_11757);
or U19524 (N_19524,N_10091,N_10209);
nand U19525 (N_19525,N_12679,N_13010);
and U19526 (N_19526,N_11000,N_13591);
nand U19527 (N_19527,N_10789,N_14647);
nand U19528 (N_19528,N_12494,N_11524);
or U19529 (N_19529,N_13515,N_14664);
and U19530 (N_19530,N_13873,N_10026);
and U19531 (N_19531,N_13101,N_13867);
nand U19532 (N_19532,N_10540,N_14791);
and U19533 (N_19533,N_11971,N_10799);
nand U19534 (N_19534,N_14927,N_10084);
nor U19535 (N_19535,N_13152,N_14531);
nand U19536 (N_19536,N_13176,N_14037);
or U19537 (N_19537,N_14957,N_12791);
nand U19538 (N_19538,N_10397,N_10267);
nor U19539 (N_19539,N_10177,N_12520);
nand U19540 (N_19540,N_14008,N_10876);
or U19541 (N_19541,N_10221,N_10233);
nand U19542 (N_19542,N_13257,N_10582);
or U19543 (N_19543,N_10449,N_13913);
and U19544 (N_19544,N_12865,N_12184);
nand U19545 (N_19545,N_14055,N_14387);
and U19546 (N_19546,N_10493,N_12031);
and U19547 (N_19547,N_13129,N_13430);
or U19548 (N_19548,N_10302,N_11769);
or U19549 (N_19549,N_11837,N_10690);
or U19550 (N_19550,N_13819,N_11067);
and U19551 (N_19551,N_13756,N_13183);
and U19552 (N_19552,N_13774,N_12574);
and U19553 (N_19553,N_10310,N_10180);
xnor U19554 (N_19554,N_14194,N_13577);
nor U19555 (N_19555,N_14793,N_14637);
nand U19556 (N_19556,N_13690,N_10715);
and U19557 (N_19557,N_10768,N_12184);
or U19558 (N_19558,N_12737,N_14386);
nand U19559 (N_19559,N_11578,N_12152);
and U19560 (N_19560,N_12170,N_11271);
xor U19561 (N_19561,N_10945,N_13000);
xnor U19562 (N_19562,N_13346,N_14793);
or U19563 (N_19563,N_14952,N_11384);
or U19564 (N_19564,N_14764,N_12429);
nand U19565 (N_19565,N_10056,N_12953);
and U19566 (N_19566,N_13353,N_11189);
nor U19567 (N_19567,N_10278,N_13519);
or U19568 (N_19568,N_13938,N_12639);
nand U19569 (N_19569,N_13572,N_12200);
and U19570 (N_19570,N_13002,N_13621);
nand U19571 (N_19571,N_13212,N_10595);
and U19572 (N_19572,N_14483,N_10902);
and U19573 (N_19573,N_14965,N_14678);
nand U19574 (N_19574,N_10226,N_10582);
nand U19575 (N_19575,N_12143,N_11817);
and U19576 (N_19576,N_11660,N_13477);
or U19577 (N_19577,N_12391,N_14602);
and U19578 (N_19578,N_10240,N_13706);
or U19579 (N_19579,N_12290,N_12709);
and U19580 (N_19580,N_14933,N_12361);
nand U19581 (N_19581,N_12562,N_10255);
and U19582 (N_19582,N_10126,N_10450);
and U19583 (N_19583,N_11673,N_13422);
nor U19584 (N_19584,N_12550,N_14932);
or U19585 (N_19585,N_14220,N_11328);
or U19586 (N_19586,N_13782,N_11046);
or U19587 (N_19587,N_11947,N_10720);
nor U19588 (N_19588,N_11428,N_13540);
nor U19589 (N_19589,N_12079,N_12023);
nor U19590 (N_19590,N_11423,N_12461);
nand U19591 (N_19591,N_12023,N_10780);
and U19592 (N_19592,N_11458,N_14570);
or U19593 (N_19593,N_12938,N_10333);
or U19594 (N_19594,N_10943,N_10443);
and U19595 (N_19595,N_11910,N_14796);
nand U19596 (N_19596,N_11987,N_12484);
nand U19597 (N_19597,N_11115,N_10905);
or U19598 (N_19598,N_13189,N_13476);
or U19599 (N_19599,N_13114,N_10910);
nor U19600 (N_19600,N_11835,N_10356);
nand U19601 (N_19601,N_13353,N_12756);
nor U19602 (N_19602,N_14709,N_12634);
nor U19603 (N_19603,N_10830,N_12594);
or U19604 (N_19604,N_12017,N_12823);
xor U19605 (N_19605,N_11497,N_10257);
and U19606 (N_19606,N_10203,N_13252);
nor U19607 (N_19607,N_14982,N_10995);
nand U19608 (N_19608,N_11365,N_12127);
nand U19609 (N_19609,N_12986,N_14678);
or U19610 (N_19610,N_12761,N_13582);
xnor U19611 (N_19611,N_10254,N_10543);
and U19612 (N_19612,N_11566,N_13312);
or U19613 (N_19613,N_10488,N_11555);
or U19614 (N_19614,N_11282,N_14441);
nor U19615 (N_19615,N_14850,N_14957);
and U19616 (N_19616,N_13541,N_14482);
nand U19617 (N_19617,N_13672,N_14602);
nand U19618 (N_19618,N_12426,N_12091);
and U19619 (N_19619,N_12191,N_11438);
and U19620 (N_19620,N_13814,N_10194);
nor U19621 (N_19621,N_10444,N_14350);
nand U19622 (N_19622,N_11433,N_13013);
xnor U19623 (N_19623,N_12280,N_13627);
or U19624 (N_19624,N_11886,N_13000);
xnor U19625 (N_19625,N_14315,N_13717);
nor U19626 (N_19626,N_14120,N_12015);
nor U19627 (N_19627,N_12923,N_13897);
and U19628 (N_19628,N_10895,N_12796);
xor U19629 (N_19629,N_13806,N_14560);
and U19630 (N_19630,N_14338,N_13743);
and U19631 (N_19631,N_10621,N_12902);
nor U19632 (N_19632,N_11642,N_11843);
nor U19633 (N_19633,N_14300,N_12718);
nor U19634 (N_19634,N_11942,N_10845);
or U19635 (N_19635,N_13969,N_11106);
nand U19636 (N_19636,N_11440,N_14474);
or U19637 (N_19637,N_14449,N_10252);
and U19638 (N_19638,N_10709,N_13612);
nand U19639 (N_19639,N_14714,N_12497);
and U19640 (N_19640,N_11913,N_14140);
xnor U19641 (N_19641,N_14925,N_12189);
nor U19642 (N_19642,N_14305,N_11033);
nor U19643 (N_19643,N_12083,N_12932);
xor U19644 (N_19644,N_13667,N_13763);
and U19645 (N_19645,N_10001,N_13037);
xor U19646 (N_19646,N_13760,N_14241);
or U19647 (N_19647,N_14409,N_10139);
nand U19648 (N_19648,N_10212,N_13830);
or U19649 (N_19649,N_12511,N_10396);
nand U19650 (N_19650,N_11249,N_12574);
nand U19651 (N_19651,N_10184,N_13348);
and U19652 (N_19652,N_13427,N_12402);
nor U19653 (N_19653,N_10674,N_10451);
nor U19654 (N_19654,N_11598,N_10049);
or U19655 (N_19655,N_10231,N_10152);
nand U19656 (N_19656,N_12271,N_10509);
nor U19657 (N_19657,N_11649,N_11513);
nand U19658 (N_19658,N_11544,N_10996);
nor U19659 (N_19659,N_11143,N_12582);
or U19660 (N_19660,N_11309,N_14528);
nor U19661 (N_19661,N_14561,N_14807);
nor U19662 (N_19662,N_12678,N_12360);
and U19663 (N_19663,N_12491,N_14260);
or U19664 (N_19664,N_13485,N_13685);
or U19665 (N_19665,N_13578,N_10860);
or U19666 (N_19666,N_13599,N_12465);
and U19667 (N_19667,N_10017,N_14283);
or U19668 (N_19668,N_12125,N_13424);
or U19669 (N_19669,N_14686,N_14548);
nor U19670 (N_19670,N_10373,N_10053);
or U19671 (N_19671,N_13606,N_12678);
or U19672 (N_19672,N_11825,N_12721);
nand U19673 (N_19673,N_12158,N_14320);
or U19674 (N_19674,N_12219,N_12344);
nor U19675 (N_19675,N_12024,N_11364);
nand U19676 (N_19676,N_10471,N_11621);
xnor U19677 (N_19677,N_13335,N_11225);
nand U19678 (N_19678,N_14959,N_14106);
or U19679 (N_19679,N_12042,N_12624);
and U19680 (N_19680,N_13721,N_11793);
or U19681 (N_19681,N_12102,N_14448);
or U19682 (N_19682,N_14360,N_12905);
or U19683 (N_19683,N_12051,N_12900);
xnor U19684 (N_19684,N_10427,N_11698);
or U19685 (N_19685,N_13370,N_13734);
nand U19686 (N_19686,N_14274,N_14249);
nor U19687 (N_19687,N_12975,N_13313);
nand U19688 (N_19688,N_13044,N_10130);
or U19689 (N_19689,N_12924,N_11406);
or U19690 (N_19690,N_14858,N_11307);
nand U19691 (N_19691,N_12225,N_11683);
nand U19692 (N_19692,N_12754,N_12986);
or U19693 (N_19693,N_13922,N_14542);
nand U19694 (N_19694,N_10595,N_10987);
nor U19695 (N_19695,N_10688,N_13872);
and U19696 (N_19696,N_14562,N_13647);
nand U19697 (N_19697,N_12631,N_14417);
nor U19698 (N_19698,N_12607,N_10415);
nor U19699 (N_19699,N_13021,N_12001);
and U19700 (N_19700,N_13317,N_14987);
nor U19701 (N_19701,N_12264,N_14875);
xnor U19702 (N_19702,N_11150,N_11420);
and U19703 (N_19703,N_14360,N_13425);
and U19704 (N_19704,N_13208,N_11712);
or U19705 (N_19705,N_14279,N_14892);
xor U19706 (N_19706,N_10514,N_13289);
nand U19707 (N_19707,N_12183,N_14663);
and U19708 (N_19708,N_12795,N_13833);
nand U19709 (N_19709,N_11798,N_10904);
nand U19710 (N_19710,N_13294,N_14534);
or U19711 (N_19711,N_10400,N_14375);
or U19712 (N_19712,N_14058,N_10582);
and U19713 (N_19713,N_13138,N_11368);
and U19714 (N_19714,N_10634,N_13733);
nor U19715 (N_19715,N_10947,N_14601);
xor U19716 (N_19716,N_11438,N_12519);
xnor U19717 (N_19717,N_14031,N_14199);
xor U19718 (N_19718,N_10319,N_14145);
nand U19719 (N_19719,N_13190,N_12735);
nand U19720 (N_19720,N_10603,N_14766);
or U19721 (N_19721,N_12163,N_12517);
nor U19722 (N_19722,N_11433,N_14304);
nand U19723 (N_19723,N_14545,N_11742);
nand U19724 (N_19724,N_11362,N_12970);
and U19725 (N_19725,N_11005,N_12632);
or U19726 (N_19726,N_14363,N_12442);
and U19727 (N_19727,N_10848,N_14827);
nor U19728 (N_19728,N_10084,N_14423);
nand U19729 (N_19729,N_11542,N_13641);
nand U19730 (N_19730,N_13625,N_13635);
xor U19731 (N_19731,N_13475,N_14867);
or U19732 (N_19732,N_10199,N_11326);
nor U19733 (N_19733,N_14707,N_13195);
and U19734 (N_19734,N_14623,N_12496);
or U19735 (N_19735,N_10165,N_11402);
and U19736 (N_19736,N_14653,N_11547);
or U19737 (N_19737,N_14013,N_12049);
nand U19738 (N_19738,N_11047,N_12136);
nand U19739 (N_19739,N_12910,N_10627);
nand U19740 (N_19740,N_11448,N_13799);
and U19741 (N_19741,N_11863,N_12484);
nor U19742 (N_19742,N_14486,N_12381);
or U19743 (N_19743,N_11035,N_13997);
nor U19744 (N_19744,N_14334,N_11007);
nor U19745 (N_19745,N_14963,N_10490);
nor U19746 (N_19746,N_11132,N_12414);
or U19747 (N_19747,N_11694,N_14030);
or U19748 (N_19748,N_12949,N_14149);
nor U19749 (N_19749,N_11751,N_10188);
nor U19750 (N_19750,N_10062,N_11669);
nor U19751 (N_19751,N_12314,N_11550);
xor U19752 (N_19752,N_14730,N_11836);
xnor U19753 (N_19753,N_12586,N_10818);
nor U19754 (N_19754,N_10808,N_14080);
and U19755 (N_19755,N_10201,N_13334);
and U19756 (N_19756,N_12512,N_13514);
nand U19757 (N_19757,N_10467,N_11784);
and U19758 (N_19758,N_11145,N_12605);
nand U19759 (N_19759,N_14930,N_13073);
nor U19760 (N_19760,N_10688,N_13855);
and U19761 (N_19761,N_11927,N_12980);
and U19762 (N_19762,N_11711,N_12342);
nor U19763 (N_19763,N_13508,N_12073);
and U19764 (N_19764,N_13179,N_11388);
nand U19765 (N_19765,N_10282,N_10387);
and U19766 (N_19766,N_14084,N_13189);
nand U19767 (N_19767,N_11257,N_11765);
xnor U19768 (N_19768,N_12571,N_11281);
nor U19769 (N_19769,N_14030,N_10831);
and U19770 (N_19770,N_14866,N_13381);
nand U19771 (N_19771,N_13698,N_11964);
nand U19772 (N_19772,N_14688,N_10405);
and U19773 (N_19773,N_14423,N_12153);
xor U19774 (N_19774,N_13770,N_13515);
or U19775 (N_19775,N_14601,N_14551);
nor U19776 (N_19776,N_13999,N_11113);
nand U19777 (N_19777,N_14090,N_10043);
nor U19778 (N_19778,N_13216,N_12643);
or U19779 (N_19779,N_12413,N_11528);
and U19780 (N_19780,N_12114,N_13350);
or U19781 (N_19781,N_13727,N_13015);
or U19782 (N_19782,N_11243,N_14507);
or U19783 (N_19783,N_12803,N_11301);
nor U19784 (N_19784,N_12290,N_11341);
or U19785 (N_19785,N_11124,N_12987);
and U19786 (N_19786,N_14895,N_11907);
xnor U19787 (N_19787,N_10609,N_14140);
xnor U19788 (N_19788,N_13817,N_10915);
xor U19789 (N_19789,N_14317,N_11684);
nor U19790 (N_19790,N_11772,N_10320);
or U19791 (N_19791,N_11361,N_12884);
and U19792 (N_19792,N_14851,N_14570);
or U19793 (N_19793,N_11341,N_14077);
and U19794 (N_19794,N_14703,N_14733);
nand U19795 (N_19795,N_13689,N_13946);
nand U19796 (N_19796,N_14916,N_14091);
or U19797 (N_19797,N_11897,N_13769);
or U19798 (N_19798,N_12518,N_12541);
or U19799 (N_19799,N_12846,N_14943);
or U19800 (N_19800,N_13247,N_13703);
or U19801 (N_19801,N_10914,N_13375);
nor U19802 (N_19802,N_10781,N_13439);
and U19803 (N_19803,N_14706,N_12048);
or U19804 (N_19804,N_14076,N_11108);
and U19805 (N_19805,N_10746,N_12199);
nor U19806 (N_19806,N_10215,N_10002);
and U19807 (N_19807,N_10866,N_10494);
and U19808 (N_19808,N_10015,N_12701);
and U19809 (N_19809,N_14515,N_14481);
or U19810 (N_19810,N_13126,N_14738);
and U19811 (N_19811,N_12960,N_14017);
nor U19812 (N_19812,N_14615,N_10145);
and U19813 (N_19813,N_10663,N_12085);
nor U19814 (N_19814,N_12590,N_11479);
nor U19815 (N_19815,N_13558,N_10945);
and U19816 (N_19816,N_14012,N_12187);
nor U19817 (N_19817,N_12031,N_12761);
nand U19818 (N_19818,N_12819,N_14852);
and U19819 (N_19819,N_10859,N_11472);
or U19820 (N_19820,N_14510,N_11124);
nor U19821 (N_19821,N_11025,N_10658);
nand U19822 (N_19822,N_10610,N_12954);
xnor U19823 (N_19823,N_13283,N_14206);
or U19824 (N_19824,N_14012,N_12512);
nand U19825 (N_19825,N_13878,N_12906);
nand U19826 (N_19826,N_13606,N_12561);
xnor U19827 (N_19827,N_12854,N_12446);
or U19828 (N_19828,N_10295,N_13074);
or U19829 (N_19829,N_11506,N_10897);
nand U19830 (N_19830,N_12836,N_13123);
nor U19831 (N_19831,N_12245,N_10713);
nand U19832 (N_19832,N_13943,N_11501);
and U19833 (N_19833,N_12350,N_12425);
nor U19834 (N_19834,N_11248,N_13590);
or U19835 (N_19835,N_14914,N_10557);
nor U19836 (N_19836,N_12912,N_10142);
and U19837 (N_19837,N_14415,N_12569);
nand U19838 (N_19838,N_10608,N_10327);
and U19839 (N_19839,N_12558,N_11323);
nor U19840 (N_19840,N_14680,N_12252);
and U19841 (N_19841,N_10825,N_14186);
or U19842 (N_19842,N_13593,N_10172);
and U19843 (N_19843,N_10890,N_12757);
and U19844 (N_19844,N_13605,N_12764);
nand U19845 (N_19845,N_12567,N_10201);
and U19846 (N_19846,N_14204,N_11686);
nor U19847 (N_19847,N_10789,N_12298);
and U19848 (N_19848,N_11137,N_11543);
xor U19849 (N_19849,N_10933,N_13919);
or U19850 (N_19850,N_13235,N_14922);
or U19851 (N_19851,N_13823,N_11973);
nor U19852 (N_19852,N_13215,N_14698);
xor U19853 (N_19853,N_11373,N_11469);
nand U19854 (N_19854,N_13954,N_12524);
or U19855 (N_19855,N_11237,N_10865);
or U19856 (N_19856,N_14783,N_10994);
nor U19857 (N_19857,N_12275,N_11236);
nand U19858 (N_19858,N_12197,N_12396);
and U19859 (N_19859,N_11749,N_12790);
nand U19860 (N_19860,N_12770,N_12706);
nor U19861 (N_19861,N_11969,N_14376);
xor U19862 (N_19862,N_13868,N_14999);
xnor U19863 (N_19863,N_11021,N_12092);
nor U19864 (N_19864,N_13874,N_14187);
or U19865 (N_19865,N_10079,N_10720);
and U19866 (N_19866,N_14697,N_11547);
nor U19867 (N_19867,N_12177,N_11100);
nand U19868 (N_19868,N_10722,N_14003);
and U19869 (N_19869,N_14501,N_10796);
or U19870 (N_19870,N_11772,N_10489);
or U19871 (N_19871,N_13330,N_13879);
nor U19872 (N_19872,N_11336,N_10551);
and U19873 (N_19873,N_13897,N_13516);
xor U19874 (N_19874,N_10070,N_12833);
xor U19875 (N_19875,N_11927,N_12092);
nand U19876 (N_19876,N_13735,N_13198);
or U19877 (N_19877,N_11386,N_12721);
nand U19878 (N_19878,N_11105,N_10679);
nor U19879 (N_19879,N_10034,N_14101);
or U19880 (N_19880,N_13068,N_11077);
and U19881 (N_19881,N_10140,N_12901);
nor U19882 (N_19882,N_12171,N_12003);
nand U19883 (N_19883,N_11660,N_14400);
nand U19884 (N_19884,N_13293,N_13010);
nor U19885 (N_19885,N_14020,N_14800);
and U19886 (N_19886,N_10914,N_14109);
or U19887 (N_19887,N_12879,N_14191);
xnor U19888 (N_19888,N_10388,N_13383);
nand U19889 (N_19889,N_11694,N_14315);
and U19890 (N_19890,N_12445,N_14486);
nand U19891 (N_19891,N_12818,N_12381);
nor U19892 (N_19892,N_13735,N_13230);
or U19893 (N_19893,N_12550,N_10291);
and U19894 (N_19894,N_10449,N_14672);
nor U19895 (N_19895,N_13818,N_14305);
nor U19896 (N_19896,N_11036,N_11555);
nor U19897 (N_19897,N_10743,N_14075);
nand U19898 (N_19898,N_10899,N_14675);
or U19899 (N_19899,N_14757,N_14144);
nand U19900 (N_19900,N_13393,N_12417);
xor U19901 (N_19901,N_13202,N_11004);
nand U19902 (N_19902,N_13474,N_14498);
nand U19903 (N_19903,N_13485,N_12332);
and U19904 (N_19904,N_14408,N_14811);
nor U19905 (N_19905,N_12446,N_14027);
xnor U19906 (N_19906,N_14389,N_10935);
and U19907 (N_19907,N_10316,N_11551);
xor U19908 (N_19908,N_10386,N_13223);
xnor U19909 (N_19909,N_13622,N_12228);
nor U19910 (N_19910,N_13368,N_14671);
nand U19911 (N_19911,N_10461,N_13328);
nor U19912 (N_19912,N_12302,N_14399);
and U19913 (N_19913,N_10766,N_14647);
nand U19914 (N_19914,N_11591,N_10014);
xnor U19915 (N_19915,N_11888,N_14099);
nor U19916 (N_19916,N_13298,N_12194);
or U19917 (N_19917,N_14332,N_11543);
nor U19918 (N_19918,N_11832,N_13462);
and U19919 (N_19919,N_13187,N_12026);
and U19920 (N_19920,N_11043,N_13623);
nor U19921 (N_19921,N_10189,N_13586);
nor U19922 (N_19922,N_10548,N_13913);
nand U19923 (N_19923,N_12053,N_14773);
or U19924 (N_19924,N_11200,N_11346);
nand U19925 (N_19925,N_12499,N_11796);
and U19926 (N_19926,N_11159,N_12017);
and U19927 (N_19927,N_14393,N_14631);
or U19928 (N_19928,N_14909,N_14564);
or U19929 (N_19929,N_10744,N_10449);
and U19930 (N_19930,N_13141,N_10313);
nor U19931 (N_19931,N_10859,N_11020);
and U19932 (N_19932,N_12298,N_10924);
or U19933 (N_19933,N_13856,N_14003);
nand U19934 (N_19934,N_13511,N_10223);
and U19935 (N_19935,N_12989,N_12134);
nand U19936 (N_19936,N_13604,N_11773);
nor U19937 (N_19937,N_12302,N_14875);
nand U19938 (N_19938,N_13820,N_10763);
xor U19939 (N_19939,N_14348,N_11722);
and U19940 (N_19940,N_13862,N_10010);
and U19941 (N_19941,N_14280,N_14169);
nor U19942 (N_19942,N_11921,N_13853);
nor U19943 (N_19943,N_13018,N_12230);
or U19944 (N_19944,N_14385,N_11657);
nor U19945 (N_19945,N_10519,N_10854);
and U19946 (N_19946,N_12653,N_11346);
or U19947 (N_19947,N_13198,N_13590);
nand U19948 (N_19948,N_12190,N_10508);
nor U19949 (N_19949,N_13276,N_14478);
nor U19950 (N_19950,N_10097,N_14631);
nand U19951 (N_19951,N_11075,N_11035);
or U19952 (N_19952,N_12198,N_14128);
or U19953 (N_19953,N_14355,N_10355);
or U19954 (N_19954,N_11010,N_12947);
and U19955 (N_19955,N_11327,N_10732);
nand U19956 (N_19956,N_10524,N_12375);
nor U19957 (N_19957,N_14842,N_12303);
nor U19958 (N_19958,N_11380,N_12256);
and U19959 (N_19959,N_14294,N_10856);
nand U19960 (N_19960,N_10261,N_12844);
and U19961 (N_19961,N_12945,N_12609);
nand U19962 (N_19962,N_10062,N_14830);
and U19963 (N_19963,N_11015,N_13619);
nand U19964 (N_19964,N_12707,N_10484);
nand U19965 (N_19965,N_10977,N_12083);
and U19966 (N_19966,N_13509,N_12426);
and U19967 (N_19967,N_10487,N_14983);
or U19968 (N_19968,N_10150,N_10787);
xor U19969 (N_19969,N_13153,N_12772);
nand U19970 (N_19970,N_13074,N_10099);
and U19971 (N_19971,N_10428,N_12617);
nand U19972 (N_19972,N_11165,N_13404);
xor U19973 (N_19973,N_11952,N_13436);
xnor U19974 (N_19974,N_12250,N_12982);
nor U19975 (N_19975,N_11025,N_13764);
and U19976 (N_19976,N_10729,N_13814);
or U19977 (N_19977,N_13444,N_13903);
nand U19978 (N_19978,N_14617,N_12875);
xor U19979 (N_19979,N_10957,N_14683);
and U19980 (N_19980,N_12507,N_13470);
and U19981 (N_19981,N_12688,N_11906);
and U19982 (N_19982,N_11222,N_10275);
and U19983 (N_19983,N_14275,N_14438);
xor U19984 (N_19984,N_14245,N_11137);
nor U19985 (N_19985,N_11562,N_12134);
or U19986 (N_19986,N_12305,N_12216);
nand U19987 (N_19987,N_10034,N_10555);
and U19988 (N_19988,N_14408,N_10036);
xnor U19989 (N_19989,N_11944,N_13405);
nor U19990 (N_19990,N_10378,N_14807);
or U19991 (N_19991,N_11077,N_12085);
nand U19992 (N_19992,N_11052,N_11698);
or U19993 (N_19993,N_14595,N_10030);
and U19994 (N_19994,N_14596,N_14570);
or U19995 (N_19995,N_14352,N_12559);
and U19996 (N_19996,N_13350,N_10134);
nand U19997 (N_19997,N_13524,N_14138);
nor U19998 (N_19998,N_12948,N_13055);
xnor U19999 (N_19999,N_10235,N_10262);
nor U20000 (N_20000,N_16627,N_15822);
nor U20001 (N_20001,N_15409,N_18640);
nor U20002 (N_20002,N_17073,N_15261);
and U20003 (N_20003,N_19839,N_18158);
nand U20004 (N_20004,N_15877,N_17322);
nand U20005 (N_20005,N_17519,N_19364);
nor U20006 (N_20006,N_18666,N_18388);
or U20007 (N_20007,N_16678,N_17275);
nand U20008 (N_20008,N_16558,N_19181);
or U20009 (N_20009,N_18625,N_15691);
nand U20010 (N_20010,N_16885,N_19956);
and U20011 (N_20011,N_16267,N_17729);
and U20012 (N_20012,N_18759,N_18806);
or U20013 (N_20013,N_16117,N_15953);
and U20014 (N_20014,N_15482,N_15717);
xnor U20015 (N_20015,N_16962,N_19985);
nor U20016 (N_20016,N_15443,N_15630);
and U20017 (N_20017,N_17038,N_17599);
nand U20018 (N_20018,N_17726,N_15972);
nor U20019 (N_20019,N_15869,N_17806);
or U20020 (N_20020,N_18154,N_18300);
nor U20021 (N_20021,N_15228,N_16033);
xnor U20022 (N_20022,N_15641,N_17916);
and U20023 (N_20023,N_16688,N_16724);
and U20024 (N_20024,N_17460,N_19532);
xnor U20025 (N_20025,N_15695,N_18817);
and U20026 (N_20026,N_18447,N_16555);
nor U20027 (N_20027,N_17120,N_16022);
nand U20028 (N_20028,N_18809,N_17461);
and U20029 (N_20029,N_17154,N_16967);
and U20030 (N_20030,N_18246,N_16895);
xnor U20031 (N_20031,N_15974,N_17072);
xnor U20032 (N_20032,N_18705,N_18429);
xnor U20033 (N_20033,N_15701,N_16234);
or U20034 (N_20034,N_16467,N_18050);
nor U20035 (N_20035,N_17888,N_17257);
and U20036 (N_20036,N_18585,N_16254);
nor U20037 (N_20037,N_19790,N_17477);
nand U20038 (N_20038,N_16485,N_19594);
nand U20039 (N_20039,N_16623,N_19322);
nor U20040 (N_20040,N_19198,N_16565);
nor U20041 (N_20041,N_15518,N_17410);
and U20042 (N_20042,N_17426,N_17628);
nor U20043 (N_20043,N_19155,N_17169);
xnor U20044 (N_20044,N_17756,N_17863);
and U20045 (N_20045,N_17899,N_15897);
or U20046 (N_20046,N_18906,N_19085);
xor U20047 (N_20047,N_18427,N_16447);
nand U20048 (N_20048,N_16387,N_16869);
and U20049 (N_20049,N_16443,N_19080);
or U20050 (N_20050,N_16228,N_17552);
and U20051 (N_20051,N_16178,N_15034);
nor U20052 (N_20052,N_19248,N_18897);
and U20053 (N_20053,N_16986,N_15496);
and U20054 (N_20054,N_15320,N_19402);
nor U20055 (N_20055,N_18579,N_19496);
xnor U20056 (N_20056,N_17068,N_19234);
nand U20057 (N_20057,N_16100,N_16344);
and U20058 (N_20058,N_15799,N_18118);
and U20059 (N_20059,N_16996,N_15159);
nand U20060 (N_20060,N_18903,N_16235);
and U20061 (N_20061,N_17697,N_16844);
nor U20062 (N_20062,N_17828,N_18120);
nand U20063 (N_20063,N_15995,N_17436);
nand U20064 (N_20064,N_19320,N_15485);
nand U20065 (N_20065,N_18849,N_19098);
and U20066 (N_20066,N_15986,N_15620);
nand U20067 (N_20067,N_19396,N_18425);
and U20068 (N_20068,N_15138,N_16489);
nor U20069 (N_20069,N_15322,N_17655);
nor U20070 (N_20070,N_18406,N_19136);
nand U20071 (N_20071,N_17700,N_16583);
or U20072 (N_20072,N_18639,N_17307);
xnor U20073 (N_20073,N_19270,N_18674);
nor U20074 (N_20074,N_16067,N_19240);
and U20075 (N_20075,N_17964,N_15164);
nand U20076 (N_20076,N_19370,N_18708);
and U20077 (N_20077,N_17130,N_19946);
nor U20078 (N_20078,N_17595,N_15240);
nor U20079 (N_20079,N_15807,N_17881);
nor U20080 (N_20080,N_17010,N_15395);
or U20081 (N_20081,N_15929,N_16308);
xnor U20082 (N_20082,N_19176,N_17128);
and U20083 (N_20083,N_17761,N_17047);
nor U20084 (N_20084,N_18880,N_15057);
nor U20085 (N_20085,N_19334,N_17055);
nor U20086 (N_20086,N_15090,N_17298);
nor U20087 (N_20087,N_15110,N_15753);
nand U20088 (N_20088,N_15369,N_17397);
and U20089 (N_20089,N_18096,N_16174);
or U20090 (N_20090,N_18930,N_18994);
and U20091 (N_20091,N_16636,N_16373);
nor U20092 (N_20092,N_16914,N_15829);
nand U20093 (N_20093,N_18170,N_18848);
or U20094 (N_20094,N_15183,N_18490);
nand U20095 (N_20095,N_17640,N_17011);
and U20096 (N_20096,N_16160,N_18859);
or U20097 (N_20097,N_15901,N_16073);
nand U20098 (N_20098,N_19523,N_19197);
or U20099 (N_20099,N_16767,N_17554);
nor U20100 (N_20100,N_19685,N_15656);
nor U20101 (N_20101,N_19141,N_16089);
nor U20102 (N_20102,N_17543,N_18622);
nand U20103 (N_20103,N_19409,N_18982);
nor U20104 (N_20104,N_17727,N_18407);
and U20105 (N_20105,N_15291,N_17938);
or U20106 (N_20106,N_19023,N_15664);
nand U20107 (N_20107,N_16310,N_18220);
xor U20108 (N_20108,N_15321,N_16955);
or U20109 (N_20109,N_17458,N_17665);
nand U20110 (N_20110,N_16091,N_18595);
or U20111 (N_20111,N_17897,N_17845);
nor U20112 (N_20112,N_15716,N_15014);
nand U20113 (N_20113,N_17358,N_15178);
and U20114 (N_20114,N_16109,N_17194);
or U20115 (N_20115,N_18749,N_17695);
and U20116 (N_20116,N_16147,N_18190);
and U20117 (N_20117,N_17550,N_18087);
nor U20118 (N_20118,N_16879,N_19306);
and U20119 (N_20119,N_15107,N_17711);
nor U20120 (N_20120,N_17875,N_15771);
nand U20121 (N_20121,N_15823,N_15751);
nor U20122 (N_20122,N_17712,N_19951);
or U20123 (N_20123,N_18829,N_16587);
or U20124 (N_20124,N_15933,N_15673);
and U20125 (N_20125,N_15464,N_18460);
and U20126 (N_20126,N_17807,N_15151);
or U20127 (N_20127,N_19840,N_17372);
nor U20128 (N_20128,N_18611,N_16113);
nor U20129 (N_20129,N_18433,N_17315);
or U20130 (N_20130,N_19324,N_16735);
or U20131 (N_20131,N_17960,N_15997);
and U20132 (N_20132,N_17575,N_18907);
nand U20133 (N_20133,N_19236,N_16013);
nor U20134 (N_20134,N_17998,N_18163);
and U20135 (N_20135,N_15102,N_18931);
and U20136 (N_20136,N_18767,N_18328);
xnor U20137 (N_20137,N_15996,N_17321);
nand U20138 (N_20138,N_19440,N_15697);
and U20139 (N_20139,N_17547,N_17438);
nor U20140 (N_20140,N_15915,N_17687);
or U20141 (N_20141,N_15837,N_16581);
or U20142 (N_20142,N_18237,N_15096);
or U20143 (N_20143,N_16070,N_15130);
nor U20144 (N_20144,N_18276,N_15682);
nor U20145 (N_20145,N_16051,N_18893);
and U20146 (N_20146,N_18701,N_16226);
nor U20147 (N_20147,N_19533,N_17401);
or U20148 (N_20148,N_18808,N_18201);
nor U20149 (N_20149,N_17814,N_17287);
or U20150 (N_20150,N_16468,N_16118);
nor U20151 (N_20151,N_18978,N_15580);
nand U20152 (N_20152,N_18899,N_18777);
or U20153 (N_20153,N_16352,N_15808);
and U20154 (N_20154,N_19480,N_18288);
or U20155 (N_20155,N_17483,N_19012);
xnor U20156 (N_20156,N_19084,N_18092);
nand U20157 (N_20157,N_18905,N_19040);
or U20158 (N_20158,N_19095,N_15191);
nand U20159 (N_20159,N_17862,N_18366);
or U20160 (N_20160,N_18016,N_18187);
nand U20161 (N_20161,N_19125,N_16090);
and U20162 (N_20162,N_15639,N_17915);
or U20163 (N_20163,N_17970,N_15353);
or U20164 (N_20164,N_16081,N_15040);
xor U20165 (N_20165,N_18617,N_17920);
and U20166 (N_20166,N_16602,N_15358);
nand U20167 (N_20167,N_15329,N_16769);
and U20168 (N_20168,N_16593,N_18732);
nand U20169 (N_20169,N_16224,N_18063);
or U20170 (N_20170,N_16074,N_18493);
nor U20171 (N_20171,N_16338,N_18814);
and U20172 (N_20172,N_16770,N_17549);
nand U20173 (N_20173,N_18748,N_19508);
nand U20174 (N_20174,N_19218,N_15039);
or U20175 (N_20175,N_15103,N_15797);
and U20176 (N_20176,N_19071,N_17997);
nand U20177 (N_20177,N_16193,N_17259);
nand U20178 (N_20178,N_19062,N_18272);
and U20179 (N_20179,N_18226,N_18000);
or U20180 (N_20180,N_17627,N_16144);
nor U20181 (N_20181,N_16573,N_18588);
nand U20182 (N_20182,N_17226,N_16177);
nand U20183 (N_20183,N_17873,N_18877);
nand U20184 (N_20184,N_19608,N_18920);
or U20185 (N_20185,N_19201,N_18721);
or U20186 (N_20186,N_15945,N_18959);
or U20187 (N_20187,N_16370,N_17715);
nand U20188 (N_20188,N_17370,N_16764);
and U20189 (N_20189,N_16086,N_18926);
nand U20190 (N_20190,N_17999,N_18383);
nand U20191 (N_20191,N_15503,N_15908);
nor U20192 (N_20192,N_18231,N_19942);
nand U20193 (N_20193,N_15490,N_19999);
or U20194 (N_20194,N_19656,N_17351);
and U20195 (N_20195,N_17696,N_17951);
nor U20196 (N_20196,N_18027,N_18234);
nor U20197 (N_20197,N_19883,N_15012);
nand U20198 (N_20198,N_16004,N_17124);
nand U20199 (N_20199,N_15694,N_18641);
or U20200 (N_20200,N_18737,N_15554);
and U20201 (N_20201,N_15275,N_19271);
or U20202 (N_20202,N_17473,N_18636);
nor U20203 (N_20203,N_16799,N_17464);
and U20204 (N_20204,N_17754,N_19779);
xor U20205 (N_20205,N_18977,N_15667);
nand U20206 (N_20206,N_16825,N_15396);
nand U20207 (N_20207,N_15839,N_19195);
nor U20208 (N_20208,N_15861,N_17724);
or U20209 (N_20209,N_15731,N_19004);
nor U20210 (N_20210,N_17798,N_17293);
nand U20211 (N_20211,N_18562,N_19327);
nor U20212 (N_20212,N_16528,N_15059);
nand U20213 (N_20213,N_18280,N_19315);
or U20214 (N_20214,N_16060,N_18553);
nand U20215 (N_20215,N_15003,N_16634);
nand U20216 (N_20216,N_17255,N_15394);
xnor U20217 (N_20217,N_18197,N_16153);
nand U20218 (N_20218,N_19529,N_19902);
nor U20219 (N_20219,N_16500,N_17883);
or U20220 (N_20220,N_17272,N_18315);
nand U20221 (N_20221,N_17495,N_16794);
xnor U20222 (N_20222,N_19471,N_18564);
and U20223 (N_20223,N_17793,N_17075);
nand U20224 (N_20224,N_15914,N_19497);
nand U20225 (N_20225,N_17809,N_18505);
nand U20226 (N_20226,N_16657,N_16450);
nor U20227 (N_20227,N_17855,N_18191);
nor U20228 (N_20228,N_15209,N_19474);
nand U20229 (N_20229,N_17859,N_16586);
nand U20230 (N_20230,N_19914,N_17071);
nand U20231 (N_20231,N_16451,N_15427);
xor U20232 (N_20232,N_18103,N_18500);
xnor U20233 (N_20233,N_16214,N_18724);
nand U20234 (N_20234,N_18519,N_17443);
xor U20235 (N_20235,N_16532,N_19089);
nor U20236 (N_20236,N_19318,N_15001);
nor U20237 (N_20237,N_19407,N_16208);
xnor U20238 (N_20238,N_18212,N_18240);
nor U20239 (N_20239,N_18360,N_15608);
and U20240 (N_20240,N_17773,N_16148);
or U20241 (N_20241,N_17136,N_17942);
or U20242 (N_20242,N_15515,N_16479);
and U20243 (N_20243,N_16881,N_17266);
nand U20244 (N_20244,N_18812,N_16376);
nor U20245 (N_20245,N_18065,N_16896);
nand U20246 (N_20246,N_17009,N_19938);
or U20247 (N_20247,N_18056,N_16732);
or U20248 (N_20248,N_19602,N_16921);
nand U20249 (N_20249,N_15679,N_16870);
and U20250 (N_20250,N_16154,N_15136);
nor U20251 (N_20251,N_17768,N_19119);
nand U20252 (N_20252,N_16733,N_19193);
nor U20253 (N_20253,N_18881,N_18340);
and U20254 (N_20254,N_16145,N_19029);
or U20255 (N_20255,N_16563,N_15265);
and U20256 (N_20256,N_18789,N_17015);
or U20257 (N_20257,N_16330,N_15836);
or U20258 (N_20258,N_18794,N_19899);
nand U20259 (N_20259,N_16689,N_17572);
and U20260 (N_20260,N_15309,N_19703);
or U20261 (N_20261,N_16142,N_18761);
nor U20262 (N_20262,N_18164,N_17502);
or U20263 (N_20263,N_15709,N_17675);
and U20264 (N_20264,N_16306,N_19960);
and U20265 (N_20265,N_16853,N_15195);
or U20266 (N_20266,N_18432,N_18682);
and U20267 (N_20267,N_16025,N_18752);
or U20268 (N_20268,N_19027,N_18779);
nand U20269 (N_20269,N_19757,N_16475);
xor U20270 (N_20270,N_18357,N_19622);
and U20271 (N_20271,N_15661,N_16557);
nor U20272 (N_20272,N_15032,N_18725);
or U20273 (N_20273,N_15120,N_17018);
or U20274 (N_20274,N_17208,N_16989);
nor U20275 (N_20275,N_18680,N_16316);
and U20276 (N_20276,N_19607,N_19578);
nand U20277 (N_20277,N_19546,N_18798);
and U20278 (N_20278,N_19880,N_18942);
or U20279 (N_20279,N_15169,N_15865);
nor U20280 (N_20280,N_17432,N_17324);
nand U20281 (N_20281,N_15864,N_15405);
and U20282 (N_20282,N_16612,N_17940);
nand U20283 (N_20283,N_18532,N_18059);
nand U20284 (N_20284,N_19720,N_16683);
nand U20285 (N_20285,N_19549,N_16001);
nor U20286 (N_20286,N_18634,N_18451);
nand U20287 (N_20287,N_18536,N_18608);
nor U20288 (N_20288,N_19127,N_16353);
nand U20289 (N_20289,N_15124,N_15348);
and U20290 (N_20290,N_19791,N_19708);
nand U20291 (N_20291,N_19067,N_15672);
or U20292 (N_20292,N_19473,N_18413);
nor U20293 (N_20293,N_17542,N_15422);
nand U20294 (N_20294,N_16917,N_18359);
nor U20295 (N_20295,N_15959,N_17922);
nor U20296 (N_20296,N_19681,N_17823);
nor U20297 (N_20297,N_15968,N_18888);
nor U20298 (N_20298,N_15549,N_15780);
nand U20299 (N_20299,N_15500,N_16650);
xor U20300 (N_20300,N_18377,N_17521);
nand U20301 (N_20301,N_18476,N_15849);
or U20302 (N_20302,N_16730,N_15636);
or U20303 (N_20303,N_19815,N_15977);
or U20304 (N_20304,N_16977,N_17591);
and U20305 (N_20305,N_17725,N_16048);
nor U20306 (N_20306,N_16960,N_18802);
nand U20307 (N_20307,N_16524,N_19196);
nand U20308 (N_20308,N_19674,N_15165);
and U20309 (N_20309,N_16886,N_16930);
nor U20310 (N_20310,N_19600,N_17593);
nand U20311 (N_20311,N_17160,N_15486);
nor U20312 (N_20312,N_16360,N_18346);
nor U20313 (N_20313,N_15884,N_16806);
nand U20314 (N_20314,N_18022,N_17592);
or U20315 (N_20315,N_19061,N_15834);
nor U20316 (N_20316,N_18953,N_18008);
nor U20317 (N_20317,N_19530,N_17805);
nor U20318 (N_20318,N_15867,N_15243);
and U20319 (N_20319,N_16832,N_19063);
nand U20320 (N_20320,N_18316,N_19599);
or U20321 (N_20321,N_19441,N_17042);
or U20322 (N_20322,N_18067,N_17288);
and U20323 (N_20323,N_19679,N_17203);
xnor U20324 (N_20324,N_16855,N_16426);
and U20325 (N_20325,N_18533,N_19545);
nor U20326 (N_20326,N_16395,N_18150);
or U20327 (N_20327,N_19557,N_19709);
or U20328 (N_20328,N_16668,N_17082);
or U20329 (N_20329,N_16206,N_18672);
or U20330 (N_20330,N_15605,N_16820);
or U20331 (N_20331,N_15802,N_17714);
xnor U20332 (N_20332,N_19255,N_16644);
and U20333 (N_20333,N_18303,N_15631);
nand U20334 (N_20334,N_18203,N_17993);
nand U20335 (N_20335,N_18842,N_18157);
and U20336 (N_20336,N_17548,N_18631);
xor U20337 (N_20337,N_16788,N_17174);
xnor U20338 (N_20338,N_19576,N_17868);
nor U20339 (N_20339,N_15654,N_19531);
or U20340 (N_20340,N_17698,N_19639);
nand U20341 (N_20341,N_18323,N_18871);
nor U20342 (N_20342,N_18879,N_16965);
and U20343 (N_20343,N_19618,N_15167);
nor U20344 (N_20344,N_18756,N_19143);
and U20345 (N_20345,N_17356,N_16165);
or U20346 (N_20346,N_18126,N_16062);
or U20347 (N_20347,N_15339,N_15544);
nand U20348 (N_20348,N_16877,N_16946);
or U20349 (N_20349,N_16401,N_15424);
nand U20350 (N_20350,N_17982,N_19073);
and U20351 (N_20351,N_15705,N_19367);
or U20352 (N_20352,N_17935,N_16579);
or U20353 (N_20353,N_15349,N_19418);
and U20354 (N_20354,N_17959,N_19456);
nor U20355 (N_20355,N_15818,N_16594);
and U20356 (N_20356,N_18075,N_19838);
nand U20357 (N_20357,N_19885,N_17149);
or U20358 (N_20358,N_19287,N_17344);
or U20359 (N_20359,N_19352,N_15800);
or U20360 (N_20360,N_18387,N_18109);
and U20361 (N_20361,N_15928,N_18463);
or U20362 (N_20362,N_17218,N_15337);
nand U20363 (N_20363,N_19107,N_19003);
nor U20364 (N_20364,N_18664,N_15474);
and U20365 (N_20365,N_19845,N_19954);
or U20366 (N_20366,N_19891,N_15457);
nor U20367 (N_20367,N_17292,N_15824);
nor U20368 (N_20368,N_18792,N_18449);
nand U20369 (N_20369,N_18440,N_19871);
and U20370 (N_20370,N_19925,N_16252);
xor U20371 (N_20371,N_15097,N_19099);
nor U20372 (N_20372,N_15913,N_18353);
nand U20373 (N_20373,N_15380,N_17784);
or U20374 (N_20374,N_17220,N_19534);
and U20375 (N_20375,N_18382,N_18475);
nand U20376 (N_20376,N_17973,N_15841);
nor U20377 (N_20377,N_16272,N_17820);
or U20378 (N_20378,N_17747,N_19214);
or U20379 (N_20379,N_18380,N_15895);
or U20380 (N_20380,N_17886,N_17650);
nor U20381 (N_20381,N_19285,N_17406);
nand U20382 (N_20382,N_17340,N_16851);
or U20383 (N_20383,N_18668,N_19087);
and U20384 (N_20384,N_17769,N_15402);
nor U20385 (N_20385,N_18511,N_18249);
nor U20386 (N_20386,N_16078,N_17424);
or U20387 (N_20387,N_15434,N_17744);
xnor U20388 (N_20388,N_16543,N_18758);
nor U20389 (N_20389,N_18145,N_18492);
and U20390 (N_20390,N_15028,N_17199);
nand U20391 (N_20391,N_19233,N_19691);
nor U20392 (N_20392,N_19064,N_15568);
nor U20393 (N_20393,N_15969,N_15367);
nor U20394 (N_20394,N_15277,N_17157);
nor U20395 (N_20395,N_19706,N_19918);
nand U20396 (N_20396,N_18730,N_18155);
nor U20397 (N_20397,N_18326,N_19974);
and U20398 (N_20398,N_19704,N_19392);
or U20399 (N_20399,N_18176,N_19332);
or U20400 (N_20400,N_18494,N_17248);
nor U20401 (N_20401,N_18816,N_19978);
or U20402 (N_20402,N_15477,N_18362);
or U20403 (N_20403,N_18914,N_15430);
nor U20404 (N_20404,N_17243,N_17533);
nand U20405 (N_20405,N_17955,N_18116);
and U20406 (N_20406,N_17923,N_16132);
xnor U20407 (N_20407,N_17109,N_15564);
and U20408 (N_20408,N_18023,N_15144);
nand U20409 (N_20409,N_18970,N_17500);
or U20410 (N_20410,N_16175,N_17636);
nand U20411 (N_20411,N_18918,N_17986);
nor U20412 (N_20412,N_19833,N_16439);
or U20413 (N_20413,N_19964,N_17908);
nor U20414 (N_20414,N_16019,N_15690);
or U20415 (N_20415,N_15406,N_16888);
xor U20416 (N_20416,N_16294,N_15479);
nand U20417 (N_20417,N_18523,N_18541);
and U20418 (N_20418,N_16709,N_18597);
xnor U20419 (N_20419,N_15763,N_17234);
nor U20420 (N_20420,N_19350,N_19200);
nand U20421 (N_20421,N_19586,N_18690);
or U20422 (N_20422,N_15011,N_18657);
and U20423 (N_20423,N_15832,N_15941);
or U20424 (N_20424,N_16544,N_16926);
nor U20425 (N_20425,N_15318,N_19953);
nor U20426 (N_20426,N_15250,N_17450);
xor U20427 (N_20427,N_18313,N_15624);
nor U20428 (N_20428,N_16848,N_19958);
and U20429 (N_20429,N_18466,N_19512);
xnor U20430 (N_20430,N_15094,N_16031);
nand U20431 (N_20431,N_15625,N_15814);
xnor U20432 (N_20432,N_16188,N_17237);
nor U20433 (N_20433,N_18497,N_16686);
or U20434 (N_20434,N_17834,N_17380);
and U20435 (N_20435,N_17232,N_18139);
nand U20436 (N_20436,N_16016,N_19314);
or U20437 (N_20437,N_18943,N_17431);
and U20438 (N_20438,N_19228,N_18077);
and U20439 (N_20439,N_19354,N_17910);
nor U20440 (N_20440,N_17223,N_16220);
nand U20441 (N_20441,N_17091,N_19091);
and U20442 (N_20442,N_19267,N_18363);
xnor U20443 (N_20443,N_16061,N_15200);
nand U20444 (N_20444,N_16497,N_15506);
and U20445 (N_20445,N_17880,N_15080);
xor U20446 (N_20446,N_15362,N_18061);
or U20447 (N_20447,N_17800,N_17144);
or U20448 (N_20448,N_18053,N_19075);
nand U20449 (N_20449,N_19305,N_18450);
nand U20450 (N_20450,N_18117,N_19303);
nor U20451 (N_20451,N_18741,N_16158);
nand U20452 (N_20452,N_15777,N_18957);
nand U20453 (N_20453,N_19031,N_15374);
nor U20454 (N_20454,N_19213,N_16204);
nor U20455 (N_20455,N_18148,N_19309);
nand U20456 (N_20456,N_19208,N_16449);
and U20457 (N_20457,N_15230,N_16569);
nand U20458 (N_20458,N_18872,N_15938);
nand U20459 (N_20459,N_16961,N_16905);
and U20460 (N_20460,N_17532,N_16281);
nand U20461 (N_20461,N_16129,N_15399);
nand U20462 (N_20462,N_16839,N_19363);
nand U20463 (N_20463,N_15619,N_19872);
nand U20464 (N_20464,N_15122,N_17586);
or U20465 (N_20465,N_19921,N_19991);
and U20466 (N_20466,N_19773,N_19949);
or U20467 (N_20467,N_18045,N_18411);
xor U20468 (N_20468,N_15702,N_17618);
nand U20469 (N_20469,N_17430,N_16523);
or U20470 (N_20470,N_16758,N_19976);
and U20471 (N_20471,N_15992,N_15086);
xnor U20472 (N_20472,N_16790,N_15598);
xnor U20473 (N_20473,N_16152,N_17471);
and U20474 (N_20474,N_16846,N_17418);
nor U20475 (N_20475,N_18800,N_16975);
nand U20476 (N_20476,N_19387,N_15127);
nor U20477 (N_20477,N_15488,N_15611);
or U20478 (N_20478,N_16264,N_17622);
nor U20479 (N_20479,N_16850,N_16780);
nor U20480 (N_20480,N_17795,N_16725);
or U20481 (N_20481,N_15534,N_16695);
and U20482 (N_20482,N_16606,N_19513);
and U20483 (N_20483,N_18473,N_15319);
xor U20484 (N_20484,N_16741,N_17968);
and U20485 (N_20485,N_16637,N_18861);
nand U20486 (N_20486,N_15617,N_15882);
nor U20487 (N_20487,N_16796,N_18810);
xnor U20488 (N_20488,N_17630,N_16225);
or U20489 (N_20489,N_16312,N_16517);
nor U20490 (N_20490,N_17146,N_17682);
or U20491 (N_20491,N_18431,N_15622);
or U20492 (N_20492,N_16472,N_18489);
nor U20493 (N_20493,N_19486,N_16538);
nor U20494 (N_20494,N_17354,N_19217);
or U20495 (N_20495,N_17029,N_17896);
or U20496 (N_20496,N_17510,N_19670);
or U20497 (N_20497,N_17398,N_16309);
or U20498 (N_20498,N_18331,N_16922);
or U20499 (N_20499,N_16490,N_18589);
nor U20500 (N_20500,N_15821,N_17413);
and U20501 (N_20501,N_15983,N_18696);
xor U20502 (N_20502,N_16321,N_16864);
and U20503 (N_20503,N_16095,N_17286);
or U20504 (N_20504,N_15081,N_16047);
or U20505 (N_20505,N_17135,N_16936);
or U20506 (N_20506,N_15898,N_16482);
xor U20507 (N_20507,N_16276,N_15494);
and U20508 (N_20508,N_18072,N_18515);
xnor U20509 (N_20509,N_15467,N_15514);
nor U20510 (N_20510,N_15385,N_15843);
or U20511 (N_20511,N_18560,N_19292);
and U20512 (N_20512,N_19043,N_17207);
or U20513 (N_20513,N_16167,N_17299);
xor U20514 (N_20514,N_18575,N_18870);
xnor U20515 (N_20515,N_18512,N_15316);
nand U20516 (N_20516,N_15978,N_16580);
and U20517 (N_20517,N_15779,N_19304);
xnor U20518 (N_20518,N_15952,N_18097);
and U20519 (N_20519,N_17083,N_17977);
or U20520 (N_20520,N_19341,N_16017);
or U20521 (N_20521,N_19741,N_15881);
or U20522 (N_20522,N_15070,N_18769);
and U20523 (N_20523,N_18916,N_15017);
and U20524 (N_20524,N_16366,N_19146);
xnor U20525 (N_20525,N_17201,N_19219);
or U20526 (N_20526,N_17080,N_18669);
nor U20527 (N_20527,N_18221,N_16871);
and U20528 (N_20528,N_17050,N_16958);
xor U20529 (N_20529,N_16970,N_19831);
nor U20530 (N_20530,N_16171,N_17832);
or U20531 (N_20531,N_19105,N_15484);
nand U20532 (N_20532,N_18416,N_19766);
or U20533 (N_20533,N_17484,N_15784);
nor U20534 (N_20534,N_15115,N_15547);
or U20535 (N_20535,N_17360,N_19419);
nor U20536 (N_20536,N_17122,N_17336);
nor U20537 (N_20537,N_16209,N_19368);
xnor U20538 (N_20538,N_19417,N_16242);
xnor U20539 (N_20539,N_18275,N_17309);
or U20540 (N_20540,N_16186,N_16085);
nor U20541 (N_20541,N_16125,N_19752);
nor U20542 (N_20542,N_17138,N_15623);
or U20543 (N_20543,N_15890,N_18199);
and U20544 (N_20544,N_16771,N_19426);
nor U20545 (N_20545,N_19395,N_15312);
and U20546 (N_20546,N_15805,N_18643);
xnor U20547 (N_20547,N_18439,N_18238);
and U20548 (N_20548,N_17639,N_17446);
or U20549 (N_20549,N_19265,N_19888);
and U20550 (N_20550,N_19180,N_16624);
or U20551 (N_20551,N_19436,N_15239);
nor U20552 (N_20552,N_15215,N_18909);
and U20553 (N_20553,N_19747,N_19301);
or U20554 (N_20554,N_16676,N_19613);
and U20555 (N_20555,N_18904,N_16584);
or U20556 (N_20556,N_17159,N_17305);
xor U20557 (N_20557,N_16740,N_18282);
nor U20558 (N_20558,N_19081,N_16945);
nand U20559 (N_20559,N_15604,N_17103);
nand U20560 (N_20560,N_19853,N_18660);
nor U20561 (N_20561,N_18678,N_17290);
nand U20562 (N_20562,N_19191,N_18675);
xnor U20563 (N_20563,N_16941,N_15199);
nand U20564 (N_20564,N_18652,N_18950);
xor U20565 (N_20565,N_19011,N_16050);
nand U20566 (N_20566,N_16480,N_15689);
or U20567 (N_20567,N_16671,N_18596);
nor U20568 (N_20568,N_18426,N_16275);
nand U20569 (N_20569,N_19008,N_17362);
nand U20570 (N_20570,N_19727,N_17147);
xor U20571 (N_20571,N_16863,N_16899);
or U20572 (N_20572,N_19068,N_16176);
nand U20573 (N_20573,N_15013,N_18153);
and U20574 (N_20574,N_15051,N_16841);
or U20575 (N_20575,N_19406,N_17027);
nand U20576 (N_20576,N_19886,N_16715);
nand U20577 (N_20577,N_15046,N_17347);
or U20578 (N_20578,N_16987,N_16168);
or U20579 (N_20579,N_19736,N_18385);
nand U20580 (N_20580,N_15047,N_15739);
nor U20581 (N_20581,N_18940,N_17277);
nor U20582 (N_20582,N_19048,N_18723);
nand U20583 (N_20583,N_15359,N_19920);
nor U20584 (N_20584,N_17282,N_19399);
nor U20585 (N_20585,N_19448,N_16382);
xnor U20586 (N_20586,N_19188,N_19078);
and U20587 (N_20587,N_17872,N_18479);
nor U20588 (N_20588,N_18161,N_17262);
and U20589 (N_20589,N_17758,N_16279);
xnor U20590 (N_20590,N_19860,N_19022);
nand U20591 (N_20591,N_19339,N_15341);
nand U20592 (N_20592,N_19129,N_18876);
nand U20593 (N_20593,N_15655,N_16023);
or U20594 (N_20594,N_16541,N_19721);
nand U20595 (N_20595,N_18948,N_19632);
or U20596 (N_20596,N_19992,N_17269);
nor U20597 (N_20597,N_16002,N_18567);
nand U20598 (N_20598,N_15675,N_19686);
nor U20599 (N_20599,N_19552,N_15475);
nand U20600 (N_20600,N_15525,N_18924);
and U20601 (N_20601,N_19492,N_18350);
xor U20602 (N_20602,N_15456,N_15513);
nand U20603 (N_20603,N_16934,N_18421);
nand U20604 (N_20604,N_18110,N_15234);
or U20605 (N_20605,N_16494,N_19571);
nand U20606 (N_20606,N_18322,N_18980);
nor U20607 (N_20607,N_16184,N_16867);
and U20608 (N_20608,N_19635,N_17377);
and U20609 (N_20609,N_18339,N_18419);
or U20610 (N_20610,N_15449,N_17143);
and U20611 (N_20611,N_15785,N_18021);
and U20612 (N_20612,N_15000,N_15671);
nand U20613 (N_20613,N_15101,N_19221);
or U20614 (N_20614,N_19784,N_16694);
or U20615 (N_20615,N_17066,N_18438);
nor U20616 (N_20616,N_19722,N_18799);
or U20617 (N_20617,N_19278,N_15891);
and U20618 (N_20618,N_16277,N_19947);
and U20619 (N_20619,N_15726,N_17647);
or U20620 (N_20620,N_16545,N_19445);
xnor U20621 (N_20621,N_19555,N_18354);
nand U20622 (N_20622,N_18933,N_16649);
nor U20623 (N_20623,N_17390,N_17205);
nor U20624 (N_20624,N_19126,N_19184);
or U20625 (N_20625,N_19957,N_17405);
nor U20626 (N_20626,N_15025,N_16521);
or U20627 (N_20627,N_18688,N_17161);
xor U20628 (N_20628,N_17557,N_16198);
nor U20629 (N_20629,N_16064,N_18698);
and U20630 (N_20630,N_18343,N_16588);
nand U20631 (N_20631,N_17156,N_17551);
nand U20632 (N_20632,N_16319,N_15756);
nor U20633 (N_20633,N_17209,N_18392);
or U20634 (N_20634,N_18782,N_16621);
or U20635 (N_20635,N_18020,N_17815);
and U20636 (N_20636,N_17468,N_16782);
and U20637 (N_20637,N_15879,N_19483);
or U20638 (N_20638,N_19455,N_15114);
and U20639 (N_20639,N_18123,N_19335);
nand U20640 (N_20640,N_17927,N_17155);
or U20641 (N_20641,N_17753,N_19746);
nand U20642 (N_20642,N_15328,N_17089);
or U20643 (N_20643,N_15157,N_18656);
nor U20644 (N_20644,N_16628,N_16943);
and U20645 (N_20645,N_15728,N_18068);
and U20646 (N_20646,N_15712,N_18151);
and U20647 (N_20647,N_15428,N_18964);
nor U20648 (N_20648,N_16477,N_19385);
nand U20649 (N_20649,N_18358,N_16662);
and U20650 (N_20650,N_19472,N_15934);
nor U20651 (N_20651,N_15920,N_15812);
nor U20652 (N_20652,N_18925,N_17534);
and U20653 (N_20653,N_19001,N_15015);
and U20654 (N_20654,N_17301,N_19575);
or U20655 (N_20655,N_15179,N_16665);
nand U20656 (N_20656,N_17041,N_18299);
and U20657 (N_20657,N_17087,N_19677);
nand U20658 (N_20658,N_16690,N_17777);
nand U20659 (N_20659,N_16397,N_18700);
and U20660 (N_20660,N_15295,N_17825);
or U20661 (N_20661,N_19572,N_16959);
nor U20662 (N_20662,N_15921,N_18728);
and U20663 (N_20663,N_17710,N_16810);
and U20664 (N_20664,N_16356,N_15391);
nand U20665 (N_20665,N_18042,N_15918);
or U20666 (N_20666,N_16104,N_18954);
xor U20667 (N_20667,N_17644,N_16181);
or U20668 (N_20668,N_15313,N_19866);
xor U20669 (N_20669,N_19573,N_16292);
nor U20670 (N_20670,N_17020,N_16367);
and U20671 (N_20671,N_19076,N_15109);
nor U20672 (N_20672,N_17204,N_15980);
xor U20673 (N_20673,N_18618,N_15323);
or U20674 (N_20674,N_15609,N_16389);
nand U20675 (N_20675,N_15252,N_16093);
xnor U20676 (N_20676,N_19930,N_17202);
nand U20677 (N_20677,N_16383,N_17722);
nor U20678 (N_20678,N_18538,N_16777);
and U20679 (N_20679,N_16032,N_19052);
and U20680 (N_20680,N_17333,N_15660);
xor U20681 (N_20681,N_15248,N_19277);
nand U20682 (N_20682,N_17110,N_17211);
nor U20683 (N_20683,N_16736,N_16314);
nand U20684 (N_20684,N_18108,N_15766);
nand U20685 (N_20685,N_19501,N_17363);
nand U20686 (N_20686,N_17933,N_16413);
xor U20687 (N_20687,N_18766,N_19452);
nor U20688 (N_20688,N_19162,N_16938);
and U20689 (N_20689,N_16358,N_19802);
nor U20690 (N_20690,N_19150,N_17113);
nor U20691 (N_20691,N_16010,N_15519);
or U20692 (N_20692,N_17371,N_17026);
and U20693 (N_20693,N_18919,N_16464);
or U20694 (N_20694,N_15652,N_15245);
and U20695 (N_20695,N_18629,N_17705);
nor U20696 (N_20696,N_16288,N_17148);
and U20697 (N_20697,N_16691,N_18378);
nor U20698 (N_20698,N_18780,N_19400);
or U20699 (N_20699,N_18296,N_18032);
nor U20700 (N_20700,N_17150,N_18763);
and U20701 (N_20701,N_17568,N_18069);
nor U20702 (N_20702,N_16562,N_16355);
and U20703 (N_20703,N_16271,N_18820);
nand U20704 (N_20704,N_15987,N_16253);
or U20705 (N_20705,N_16219,N_18011);
nor U20706 (N_20706,N_17439,N_18609);
and U20707 (N_20707,N_19769,N_15154);
nor U20708 (N_20708,N_17302,N_19194);
or U20709 (N_20709,N_15111,N_18771);
nor U20710 (N_20710,N_19021,N_17585);
or U20711 (N_20711,N_18673,N_17088);
nand U20712 (N_20712,N_17037,N_18968);
nor U20713 (N_20713,N_19416,N_17402);
nor U20714 (N_20714,N_16603,N_15737);
nor U20715 (N_20715,N_17329,N_15795);
nor U20716 (N_20716,N_16324,N_17316);
xnor U20717 (N_20717,N_15022,N_18658);
and U20718 (N_20718,N_18935,N_16140);
and U20719 (N_20719,N_18841,N_18868);
nand U20720 (N_20720,N_19751,N_18271);
nand U20721 (N_20721,N_16518,N_16030);
or U20722 (N_20722,N_18891,N_19477);
and U20723 (N_20723,N_15883,N_16195);
and U20724 (N_20724,N_17569,N_19225);
nor U20725 (N_20725,N_15736,N_17779);
nand U20726 (N_20726,N_18774,N_15288);
and U20727 (N_20727,N_19625,N_18894);
nor U20728 (N_20728,N_19836,N_18038);
nand U20729 (N_20729,N_16102,N_16372);
nand U20730 (N_20730,N_15692,N_18811);
nor U20731 (N_20731,N_16719,N_18713);
nor U20732 (N_20732,N_17619,N_17992);
or U20733 (N_20733,N_16164,N_17489);
nand U20734 (N_20734,N_17317,N_15910);
and U20735 (N_20735,N_15408,N_16574);
and U20736 (N_20736,N_16937,N_17475);
and U20737 (N_20737,N_18824,N_16616);
nor U20738 (N_20738,N_19079,N_19268);
and U20739 (N_20739,N_16659,N_15658);
nor U20740 (N_20740,N_18443,N_18029);
xnor U20741 (N_20741,N_19877,N_17917);
nor U20742 (N_20742,N_16084,N_15497);
xor U20743 (N_20743,N_18441,N_18482);
or U20744 (N_20744,N_16131,N_16956);
and U20745 (N_20745,N_18398,N_17115);
nor U20746 (N_20746,N_19186,N_15296);
and U20747 (N_20747,N_17263,N_17811);
nor U20748 (N_20748,N_19631,N_19515);
nand U20749 (N_20749,N_17912,N_15140);
or U20750 (N_20750,N_16241,N_15640);
nand U20751 (N_20751,N_18470,N_18537);
and U20752 (N_20752,N_16099,N_16261);
nor U20753 (N_20753,N_18485,N_17576);
xnor U20754 (N_20754,N_17008,N_17078);
nand U20755 (N_20755,N_16465,N_17635);
and U20756 (N_20756,N_16631,N_19178);
nand U20757 (N_20757,N_16827,N_17801);
nand U20758 (N_20758,N_19086,N_16894);
and U20759 (N_20759,N_18591,N_16748);
nand U20760 (N_20760,N_19518,N_16034);
nand U20761 (N_20761,N_18394,N_17214);
and U20762 (N_20762,N_19585,N_17892);
xor U20763 (N_20763,N_19556,N_19652);
or U20764 (N_20764,N_15446,N_18257);
or U20765 (N_20765,N_15233,N_15258);
nor U20766 (N_20766,N_16575,N_17658);
or U20767 (N_20767,N_16290,N_18209);
and U20768 (N_20768,N_17774,N_17171);
or U20769 (N_20769,N_15299,N_18136);
nor U20770 (N_20770,N_17291,N_15653);
or U20771 (N_20771,N_18208,N_15850);
nor U20772 (N_20772,N_16128,N_17794);
and U20773 (N_20773,N_18222,N_18606);
and U20774 (N_20774,N_18294,N_16374);
and U20775 (N_20775,N_18223,N_15062);
or U20776 (N_20776,N_18152,N_16597);
and U20777 (N_20777,N_17581,N_17215);
or U20778 (N_20778,N_18554,N_15842);
nand U20779 (N_20779,N_15720,N_15875);
xnor U20780 (N_20780,N_17422,N_16437);
xor U20781 (N_20781,N_18801,N_19189);
nor U20782 (N_20782,N_18704,N_18974);
nand U20783 (N_20783,N_19156,N_16556);
or U20784 (N_20784,N_15926,N_18361);
and U20785 (N_20785,N_19627,N_16951);
and U20786 (N_20786,N_15286,N_17142);
nand U20787 (N_20787,N_16026,N_15581);
nand U20788 (N_20788,N_17378,N_17074);
or U20789 (N_20789,N_19716,N_15863);
or U20790 (N_20790,N_17667,N_15210);
or U20791 (N_20791,N_18227,N_16106);
nor U20792 (N_20792,N_15633,N_16632);
and U20793 (N_20793,N_15931,N_15985);
nor U20794 (N_20794,N_17476,N_15037);
xnor U20795 (N_20795,N_16840,N_19689);
or U20796 (N_20796,N_19963,N_15029);
and U20797 (N_20797,N_19275,N_16236);
or U20798 (N_20798,N_19495,N_19481);
nand U20799 (N_20799,N_16585,N_15055);
nand U20800 (N_20800,N_17444,N_17104);
nor U20801 (N_20801,N_15249,N_18367);
or U20802 (N_20802,N_15586,N_18912);
nand U20803 (N_20803,N_15356,N_18293);
nor U20804 (N_20804,N_16831,N_15056);
nor U20805 (N_20805,N_19487,N_15727);
nand U20806 (N_20806,N_18644,N_15613);
nand U20807 (N_20807,N_16289,N_15175);
or U20808 (N_20808,N_16826,N_16315);
nand U20809 (N_20809,N_16763,N_17173);
xnor U20810 (N_20810,N_17216,N_19514);
and U20811 (N_20811,N_16150,N_16496);
and U20812 (N_20812,N_18743,N_17374);
and U20813 (N_20813,N_19413,N_19241);
or U20814 (N_20814,N_16337,N_19680);
and U20815 (N_20815,N_19952,N_18464);
and U20816 (N_20816,N_16098,N_15820);
and U20817 (N_20817,N_19777,N_15649);
and U20818 (N_20818,N_18544,N_15835);
or U20819 (N_20819,N_18577,N_17810);
nand U20820 (N_20820,N_15809,N_17731);
or U20821 (N_20821,N_18983,N_19982);
nor U20822 (N_20822,N_19917,N_17610);
xnor U20823 (N_20823,N_18572,N_16318);
nor U20824 (N_20824,N_17976,N_18430);
or U20825 (N_20825,N_16713,N_17186);
or U20826 (N_20826,N_17121,N_16915);
nand U20827 (N_20827,N_19846,N_19139);
nand U20828 (N_20828,N_17004,N_18107);
nor U20829 (N_20829,N_16697,N_15857);
xor U20830 (N_20830,N_16992,N_16182);
nand U20831 (N_20831,N_16749,N_16708);
nor U20832 (N_20832,N_16744,N_17482);
nor U20833 (N_20833,N_18066,N_19768);
or U20834 (N_20834,N_16700,N_19036);
or U20835 (N_20835,N_16082,N_19245);
nand U20836 (N_20836,N_19222,N_16830);
or U20837 (N_20837,N_15668,N_17451);
and U20838 (N_20838,N_19822,N_16018);
xor U20839 (N_20839,N_17330,N_15084);
and U20840 (N_20840,N_17312,N_19797);
or U20841 (N_20841,N_18522,N_16223);
or U20842 (N_20842,N_19042,N_17659);
and U20843 (N_20843,N_17395,N_17949);
nor U20844 (N_20844,N_16873,N_18706);
nand U20845 (N_20845,N_18348,N_16838);
or U20846 (N_20846,N_16942,N_16645);
and U20847 (N_20847,N_17737,N_15508);
and U20848 (N_20848,N_16212,N_16059);
nand U20849 (N_20849,N_16750,N_19393);
and U20850 (N_20850,N_19118,N_19111);
and U20851 (N_20851,N_15874,N_15194);
and U20852 (N_20852,N_18990,N_17713);
xnor U20853 (N_20853,N_18410,N_18375);
and U20854 (N_20854,N_16139,N_17179);
and U20855 (N_20855,N_17594,N_15006);
xnor U20856 (N_20856,N_15026,N_16779);
or U20857 (N_20857,N_19809,N_15994);
and U20858 (N_20858,N_16000,N_17946);
or U20859 (N_20859,N_15572,N_18804);
or U20860 (N_20860,N_17185,N_18101);
and U20861 (N_20861,N_16190,N_16540);
or U20862 (N_20862,N_17849,N_19174);
nor U20863 (N_20863,N_16274,N_17518);
and U20864 (N_20864,N_15788,N_15492);
or U20865 (N_20865,N_15912,N_18580);
and U20866 (N_20866,N_18060,N_17285);
and U20867 (N_20867,N_18778,N_16222);
nor U20868 (N_20868,N_15610,N_17212);
nand U20869 (N_20869,N_15259,N_19617);
xnor U20870 (N_20870,N_18178,N_18175);
nand U20871 (N_20871,N_15150,N_15281);
or U20872 (N_20872,N_16446,N_17918);
and U20873 (N_20873,N_16862,N_18241);
xnor U20874 (N_20874,N_19059,N_17178);
and U20875 (N_20875,N_16599,N_15419);
nor U20876 (N_20876,N_18863,N_18965);
nor U20877 (N_20877,N_17437,N_15336);
or U20878 (N_20878,N_15118,N_17567);
or U20879 (N_20879,N_15597,N_19805);
xor U20880 (N_20880,N_16630,N_19684);
nand U20881 (N_20881,N_18711,N_18244);
xnor U20882 (N_20882,N_18114,N_19290);
xnor U20883 (N_20883,N_16809,N_18507);
or U20884 (N_20884,N_15095,N_19697);
and U20885 (N_20885,N_19882,N_16610);
or U20886 (N_20886,N_18715,N_17869);
xor U20887 (N_20887,N_17325,N_19535);
nor U20888 (N_20888,N_16380,N_18866);
nor U20889 (N_20889,N_16995,N_16038);
nand U20890 (N_20890,N_15507,N_18613);
xor U20891 (N_20891,N_18781,N_15365);
and U20892 (N_20892,N_17877,N_16527);
and U20893 (N_20893,N_18647,N_19185);
or U20894 (N_20894,N_16371,N_17003);
or U20895 (N_20895,N_15351,N_17093);
and U20896 (N_20896,N_18854,N_18783);
nor U20897 (N_20897,N_15290,N_19969);
xnor U20898 (N_20898,N_15089,N_15827);
xnor U20899 (N_20899,N_15108,N_18232);
or U20900 (N_20900,N_16702,N_18633);
or U20901 (N_20901,N_16684,N_19828);
and U20902 (N_20902,N_18054,N_19259);
and U20903 (N_20903,N_17051,N_15811);
and U20904 (N_20904,N_15602,N_19308);
and U20905 (N_20905,N_17099,N_18287);
nand U20906 (N_20906,N_18593,N_17448);
nor U20907 (N_20907,N_19665,N_16065);
nor U20908 (N_20908,N_16410,N_16618);
or U20909 (N_20909,N_19164,N_16280);
and U20910 (N_20910,N_19311,N_15271);
and U20911 (N_20911,N_16364,N_19892);
or U20912 (N_20912,N_15903,N_18689);
nand U20913 (N_20913,N_19609,N_16080);
or U20914 (N_20914,N_19865,N_15724);
and U20915 (N_20915,N_16944,N_17350);
nand U20916 (N_20916,N_15520,N_19242);
nor U20917 (N_20917,N_17228,N_15971);
or U20918 (N_20918,N_19743,N_15204);
nor U20919 (N_20919,N_16629,N_16282);
nand U20920 (N_20920,N_19927,N_19431);
xor U20921 (N_20921,N_18928,N_19307);
nor U20922 (N_20922,N_17742,N_17515);
nor U20923 (N_20923,N_18393,N_18182);
or U20924 (N_20924,N_15767,N_17934);
nand U20925 (N_20925,N_17947,N_19733);
nand U20926 (N_20926,N_15076,N_17005);
nor U20927 (N_20927,N_15223,N_15902);
or U20928 (N_20928,N_15093,N_16753);
and U20929 (N_20929,N_16405,N_18733);
nor U20930 (N_20930,N_17717,N_19693);
and U20931 (N_20931,N_19858,N_17980);
nand U20932 (N_20932,N_18099,N_19738);
and U20933 (N_20933,N_18314,N_19072);
nand U20934 (N_20934,N_19867,N_19101);
nand U20935 (N_20935,N_15455,N_16155);
nor U20936 (N_20936,N_18312,N_16336);
nand U20937 (N_20937,N_18477,N_16243);
or U20938 (N_20938,N_17812,N_17972);
and U20939 (N_20939,N_17492,N_16357);
nand U20940 (N_20940,N_15775,N_18469);
nand U20941 (N_20941,N_16742,N_19796);
or U20942 (N_20942,N_18219,N_16861);
nor U20943 (N_20943,N_18334,N_16409);
or U20944 (N_20944,N_17273,N_18504);
or U20945 (N_20945,N_15160,N_17236);
xnor U20946 (N_20946,N_17787,N_16112);
and U20947 (N_20947,N_15077,N_15806);
nand U20948 (N_20948,N_17822,N_19446);
xnor U20949 (N_20949,N_15893,N_15787);
and U20950 (N_20950,N_18695,N_19908);
nor U20951 (N_20951,N_18604,N_16834);
nor U20952 (N_20952,N_17663,N_17012);
and U20953 (N_20953,N_19390,N_19653);
nand U20954 (N_20954,N_16427,N_19398);
or U20955 (N_20955,N_19066,N_19567);
nor U20956 (N_20956,N_16124,N_19998);
and U20957 (N_20957,N_19971,N_17393);
and U20958 (N_20958,N_17870,N_17996);
or U20959 (N_20959,N_16707,N_19507);
nand U20960 (N_20960,N_18509,N_17824);
xnor U20961 (N_20961,N_17379,N_15862);
nand U20962 (N_20962,N_15030,N_17749);
and U20963 (N_20963,N_17842,N_17654);
nor U20964 (N_20964,N_19696,N_15612);
nor U20965 (N_20965,N_18242,N_17463);
and U20966 (N_20966,N_19905,N_18295);
nor U20967 (N_20967,N_19582,N_19500);
and U20968 (N_20968,N_16774,N_16448);
nor U20969 (N_20969,N_15134,N_16295);
nor U20970 (N_20970,N_17797,N_17913);
and U20971 (N_20971,N_18167,N_18194);
and U20972 (N_20972,N_15036,N_17420);
and U20973 (N_20973,N_15216,N_15774);
and U20974 (N_20974,N_18274,N_18734);
nor U20975 (N_20975,N_17987,N_18621);
and U20976 (N_20976,N_15182,N_16991);
nor U20977 (N_20977,N_17320,N_19331);
or U20978 (N_20978,N_16721,N_17459);
nand U20979 (N_20979,N_16891,N_16530);
nand U20980 (N_20980,N_18927,N_19910);
nor U20981 (N_20981,N_18755,N_18002);
nand U20982 (N_20982,N_19433,N_16436);
nor U20983 (N_20983,N_17718,N_17723);
nand U20984 (N_20984,N_17063,N_17295);
xor U20985 (N_20985,N_17796,N_17493);
or U20986 (N_20986,N_16567,N_19564);
nor U20987 (N_20987,N_16550,N_19187);
xor U20988 (N_20988,N_19391,N_15335);
nand U20989 (N_20989,N_16502,N_18192);
or U20990 (N_20990,N_17835,N_15722);
or U20991 (N_20991,N_15487,N_18351);
nand U20992 (N_20992,N_19730,N_19026);
and U20993 (N_20993,N_19110,N_16775);
nand U20994 (N_20994,N_18006,N_19264);
nor U20995 (N_20995,N_19979,N_19009);
nor U20996 (N_20996,N_15559,N_18217);
nand U20997 (N_20997,N_17661,N_15651);
nand U20998 (N_20998,N_18548,N_18436);
nand U20999 (N_20999,N_17874,N_18626);
nor U21000 (N_21000,N_19516,N_19377);
or U21001 (N_21001,N_19161,N_16130);
nand U21002 (N_21002,N_16045,N_18546);
nor U21003 (N_21003,N_18183,N_18691);
nor U21004 (N_21004,N_19520,N_19205);
nand U21005 (N_21005,N_18514,N_17022);
or U21006 (N_21006,N_15352,N_18598);
and U21007 (N_21007,N_16800,N_19658);
nor U21008 (N_21008,N_17097,N_19254);
nand U21009 (N_21009,N_18009,N_17059);
xor U21010 (N_21010,N_17914,N_16731);
nand U21011 (N_21011,N_15232,N_19919);
nand U21012 (N_21012,N_18403,N_19355);
nand U21013 (N_21013,N_18409,N_19794);
and U21014 (N_21014,N_15792,N_15306);
nand U21015 (N_21015,N_16993,N_18224);
nor U21016 (N_21016,N_15068,N_16087);
nor U21017 (N_21017,N_17400,N_19807);
nor U21018 (N_21018,N_18508,N_17789);
or U21019 (N_21019,N_17530,N_19995);
or U21020 (N_21020,N_16605,N_15742);
nor U21021 (N_21021,N_16507,N_16743);
nand U21022 (N_21022,N_16681,N_17803);
or U21023 (N_21023,N_15342,N_17514);
nand U21024 (N_21024,N_17782,N_16369);
or U21025 (N_21025,N_16056,N_18389);
nor U21026 (N_21026,N_19898,N_17590);
or U21027 (N_21027,N_15939,N_18442);
xnor U21028 (N_21028,N_15871,N_18830);
nand U21029 (N_21029,N_19881,N_15272);
and U21030 (N_21030,N_19294,N_15714);
and U21031 (N_21031,N_17562,N_16611);
or U21032 (N_21032,N_18785,N_16762);
and U21033 (N_21033,N_15024,N_16483);
nor U21034 (N_21034,N_19932,N_17509);
nor U21035 (N_21035,N_18298,N_18662);
nor U21036 (N_21036,N_17704,N_16519);
and U21037 (N_21037,N_15338,N_16561);
nor U21038 (N_21038,N_19169,N_17944);
nor U21039 (N_21039,N_18853,N_17582);
xor U21040 (N_21040,N_16138,N_15590);
nand U21041 (N_21041,N_19939,N_15447);
or U21042 (N_21042,N_15255,N_15909);
and U21043 (N_21043,N_17606,N_16348);
nand U21044 (N_21044,N_16180,N_16643);
nor U21045 (N_21045,N_17191,N_17034);
nor U21046 (N_21046,N_18702,N_16658);
or U21047 (N_21047,N_19432,N_17499);
nand U21048 (N_21048,N_17346,N_16860);
and U21049 (N_21049,N_19710,N_15262);
nand U21050 (N_21050,N_16954,N_19249);
nor U21051 (N_21051,N_17311,N_17804);
and U21052 (N_21052,N_16675,N_15826);
nor U21053 (N_21053,N_15038,N_16710);
nand U21054 (N_21054,N_17494,N_15758);
and U21055 (N_21055,N_16933,N_19827);
nand U21056 (N_21056,N_16897,N_15198);
nor U21057 (N_21057,N_17520,N_15950);
nand U21058 (N_21058,N_18079,N_15764);
xnor U21059 (N_21059,N_18699,N_16607);
and U21060 (N_21060,N_18875,N_18031);
nand U21061 (N_21061,N_15301,N_19170);
nand U21062 (N_21062,N_16526,N_15188);
xnor U21063 (N_21063,N_19538,N_17841);
and U21064 (N_21064,N_15595,N_18740);
and U21065 (N_21065,N_17561,N_15783);
nand U21066 (N_21066,N_15629,N_15606);
nand U21067 (N_21067,N_16287,N_15343);
and U21068 (N_21068,N_17643,N_19204);
or U21069 (N_21069,N_19148,N_17852);
and U21070 (N_21070,N_17677,N_16411);
nor U21071 (N_21071,N_17381,N_19347);
and U21072 (N_21072,N_15493,N_17657);
and U21073 (N_21073,N_18457,N_19889);
nand U21074 (N_21074,N_19296,N_17002);
nand U21075 (N_21075,N_18583,N_16425);
nor U21076 (N_21076,N_19756,N_19302);
or U21077 (N_21077,N_17615,N_16066);
nand U21078 (N_21078,N_15889,N_18825);
nor U21079 (N_21079,N_16878,N_17133);
and U21080 (N_21080,N_16858,N_18277);
xor U21081 (N_21081,N_15848,N_19132);
and U21082 (N_21082,N_18576,N_19397);
xnor U21083 (N_21083,N_18665,N_17407);
nand U21084 (N_21084,N_16952,N_15270);
nor U21085 (N_21085,N_15516,N_16331);
nor U21086 (N_21086,N_17601,N_18753);
and U21087 (N_21087,N_16009,N_15373);
xor U21088 (N_21088,N_18901,N_16548);
nand U21089 (N_21089,N_15235,N_15063);
or U21090 (N_21090,N_16919,N_18496);
nor U21091 (N_21091,N_18149,N_17588);
and U21092 (N_21092,N_17600,N_19786);
or U21093 (N_21093,N_17775,N_16950);
nand U21094 (N_21094,N_18552,N_17819);
nor U21095 (N_21095,N_16913,N_16291);
nor U21096 (N_21096,N_17187,N_18127);
xnor U21097 (N_21097,N_18111,N_15505);
or U21098 (N_21098,N_19374,N_15112);
nor U21099 (N_21099,N_18844,N_18936);
or U21100 (N_21100,N_19521,N_16533);
or U21101 (N_21101,N_19216,N_16077);
nand U21102 (N_21102,N_18654,N_17539);
and U21103 (N_21103,N_18216,N_19046);
nor U21104 (N_21104,N_15708,N_17054);
nand U21105 (N_21105,N_18128,N_16185);
and U21106 (N_21106,N_15010,N_16134);
nor U21107 (N_21107,N_18525,N_19410);
xor U21108 (N_21108,N_19864,N_15700);
xor U21109 (N_21109,N_18335,N_18852);
nand U21110 (N_21110,N_18481,N_18364);
nand U21111 (N_21111,N_18570,N_19152);
or U21112 (N_21112,N_15184,N_17743);
nor U21113 (N_21113,N_16365,N_16875);
and U21114 (N_21114,N_19203,N_19338);
and U21115 (N_21115,N_15535,N_15173);
and U21116 (N_21116,N_15376,N_19475);
and U21117 (N_21117,N_17969,N_19224);
and U21118 (N_21118,N_19461,N_15287);
or U21119 (N_21119,N_15483,N_18952);
and U21120 (N_21120,N_17296,N_19379);
nor U21121 (N_21121,N_17603,N_15279);
nand U21122 (N_21122,N_16974,N_16481);
and U21123 (N_21123,N_17602,N_16551);
nand U21124 (N_21124,N_16595,N_15501);
nand U21125 (N_21125,N_17838,N_15546);
nand U21126 (N_21126,N_19977,N_19775);
or U21127 (N_21127,N_15566,N_15666);
nor U21128 (N_21128,N_15364,N_17958);
nand U21129 (N_21129,N_16906,N_19547);
or U21130 (N_21130,N_18138,N_17452);
nor U21131 (N_21131,N_16642,N_17479);
nand U21132 (N_21132,N_18373,N_16883);
nor U21133 (N_21133,N_18412,N_19358);
or U21134 (N_21134,N_15469,N_18292);
nand U21135 (N_21135,N_16596,N_17219);
nor U21136 (N_21136,N_17261,N_19644);
or U21137 (N_21137,N_17181,N_15333);
and U21138 (N_21138,N_15963,N_16664);
and U21139 (N_21139,N_15621,N_19673);
nand U21140 (N_21140,N_16969,N_19509);
nor U21141 (N_21141,N_15657,N_18135);
nor U21142 (N_21142,N_19171,N_18661);
nor U21143 (N_21143,N_19987,N_15730);
nand U21144 (N_21144,N_18281,N_15680);
xnor U21145 (N_21145,N_19893,N_19749);
xnor U21146 (N_21146,N_17740,N_15735);
nor U21147 (N_21147,N_17516,N_18616);
and U21148 (N_21148,N_15548,N_15244);
or U21149 (N_21149,N_18044,N_15071);
or U21150 (N_21150,N_19799,N_17006);
or U21151 (N_21151,N_15326,N_16305);
nand U21152 (N_21152,N_15079,N_19427);
or U21153 (N_21153,N_15218,N_16592);
or U21154 (N_21154,N_17052,N_16257);
or U21155 (N_21155,N_18423,N_19428);
nand U21156 (N_21156,N_15186,N_15676);
or U21157 (N_21157,N_16283,N_15523);
nand U21158 (N_21158,N_15851,N_17531);
nand U21159 (N_21159,N_19158,N_15499);
and U21160 (N_21160,N_17435,N_18890);
nor U21161 (N_21161,N_17419,N_19961);
nor U21162 (N_21162,N_18624,N_16564);
or U21163 (N_21163,N_19638,N_18956);
and U21164 (N_21164,N_16362,N_15431);
and U21165 (N_21165,N_17545,N_18188);
nor U21166 (N_21166,N_16772,N_19873);
nand U21167 (N_21167,N_18196,N_16419);
nand U21168 (N_21168,N_15794,N_17123);
xor U21169 (N_21169,N_18047,N_19165);
and U21170 (N_21170,N_19563,N_18727);
and U21171 (N_21171,N_17361,N_15747);
nor U21172 (N_21172,N_17445,N_15561);
and U21173 (N_21173,N_19388,N_18963);
xor U21174 (N_21174,N_17365,N_19782);
and U21175 (N_21175,N_15495,N_18453);
and U21176 (N_21176,N_15642,N_17746);
nand U21177 (N_21177,N_19875,N_15207);
nor U21178 (N_21178,N_16795,N_19542);
nor U21179 (N_21179,N_16417,N_17952);
nand U21180 (N_21180,N_16262,N_15009);
nor U21181 (N_21181,N_18166,N_17375);
and U21182 (N_21182,N_15556,N_17720);
nor U21183 (N_21183,N_19745,N_17571);
nor U21184 (N_21184,N_19758,N_16166);
nor U21185 (N_21185,N_17151,N_18284);
xor U21186 (N_21186,N_18306,N_18772);
nand U21187 (N_21187,N_16021,N_18587);
or U21188 (N_21188,N_15888,N_16737);
nand U21189 (N_21189,N_17085,N_19384);
nand U21190 (N_21190,N_18543,N_17118);
xnor U21191 (N_21191,N_16669,N_15370);
nand U21192 (N_21192,N_18620,N_18390);
xnor U21193 (N_21193,N_15361,N_15379);
nor U21194 (N_21194,N_18165,N_19420);
nand U21195 (N_21195,N_19647,N_16981);
or U21196 (N_21196,N_18703,N_16617);
and U21197 (N_21197,N_19645,N_18932);
and U21198 (N_21198,N_19160,N_15278);
and U21199 (N_21199,N_17056,N_17760);
xor U21200 (N_21200,N_15201,N_16386);
nand U21201 (N_21201,N_16396,N_17247);
or U21202 (N_21202,N_18100,N_15947);
or U21203 (N_21203,N_15563,N_16798);
or U21204 (N_21204,N_15786,N_17102);
and U21205 (N_21205,N_17653,N_17357);
or U21206 (N_21206,N_16968,N_15436);
nand U21207 (N_21207,N_17652,N_15119);
or U21208 (N_21208,N_18266,N_15646);
xnor U21209 (N_21209,N_18997,N_17759);
nand U21210 (N_21210,N_17668,N_19702);
xnor U21211 (N_21211,N_15411,N_15574);
or U21212 (N_21212,N_16363,N_18049);
xnor U21213 (N_21213,N_16141,N_19356);
and U21214 (N_21214,N_18684,N_15964);
and U21215 (N_21215,N_16270,N_17183);
nor U21216 (N_21216,N_18073,N_17728);
nor U21217 (N_21217,N_18371,N_17741);
nand U21218 (N_21218,N_15533,N_18228);
xor U21219 (N_21219,N_18793,N_19227);
nor U21220 (N_21220,N_18189,N_15155);
and U21221 (N_21221,N_17745,N_15264);
and U21222 (N_21222,N_18355,N_18822);
nor U21223 (N_21223,N_16304,N_18981);
or U21224 (N_21224,N_15989,N_16670);
nand U21225 (N_21225,N_15135,N_17386);
or U21226 (N_21226,N_16786,N_18215);
nor U21227 (N_21227,N_17847,N_18499);
or U21228 (N_21228,N_19006,N_15283);
or U21229 (N_21229,N_15274,N_16512);
or U21230 (N_21230,N_18184,N_19298);
nor U21231 (N_21231,N_16932,N_15798);
xnor U21232 (N_21232,N_17131,N_15105);
nor U21233 (N_21233,N_16755,N_16620);
or U21234 (N_21234,N_19715,N_19764);
nor U21235 (N_21235,N_16052,N_16412);
and U21236 (N_21236,N_15330,N_19163);
nand U21237 (N_21237,N_16948,N_18518);
and U21238 (N_21238,N_17953,N_19699);
nand U21239 (N_21239,N_15521,N_18855);
nor U21240 (N_21240,N_16349,N_18590);
and U21241 (N_21241,N_16239,N_16971);
nor U21242 (N_21242,N_17686,N_18750);
xnor U21243 (N_21243,N_15064,N_18989);
or U21244 (N_21244,N_15023,N_18655);
or U21245 (N_21245,N_15478,N_17105);
nor U21246 (N_21246,N_19612,N_17879);
nor U21247 (N_21247,N_18486,N_17898);
xor U21248 (N_21248,N_18757,N_19857);
nand U21249 (N_21249,N_15162,N_19092);
and U21250 (N_21250,N_17919,N_18803);
and U21251 (N_21251,N_15965,N_17389);
nor U21252 (N_21252,N_19055,N_17616);
xor U21253 (N_21253,N_16196,N_15993);
nor U21254 (N_21254,N_18566,N_16738);
and U21255 (N_21255,N_16415,N_18527);
and U21256 (N_21256,N_17672,N_18446);
nand U21257 (N_21257,N_15991,N_17827);
nand U21258 (N_21258,N_18356,N_15018);
and U21259 (N_21259,N_15171,N_15378);
and U21260 (N_21260,N_16159,N_15577);
nor U21261 (N_21261,N_18172,N_15951);
nor U21262 (N_21262,N_18376,N_15260);
or U21263 (N_21263,N_19173,N_18889);
nor U21264 (N_21264,N_19755,N_15582);
nor U21265 (N_21265,N_17831,N_15626);
nor U21266 (N_21266,N_16714,N_16903);
or U21267 (N_21267,N_17508,N_16024);
nand U21268 (N_21268,N_19389,N_16404);
nor U21269 (N_21269,N_15340,N_15454);
or U21270 (N_21270,N_19568,N_17689);
nor U21271 (N_21271,N_18081,N_16776);
nor U21272 (N_21272,N_18896,N_15504);
nor U21273 (N_21273,N_19566,N_15227);
or U21274 (N_21274,N_17537,N_19522);
or U21275 (N_21275,N_15242,N_15246);
and U21276 (N_21276,N_15375,N_19159);
or U21277 (N_21277,N_15975,N_16332);
nor U21278 (N_21278,N_18581,N_18408);
nand U21279 (N_21279,N_16335,N_19876);
and U21280 (N_21280,N_15305,N_17670);
or U21281 (N_21281,N_16660,N_19439);
or U21282 (N_21282,N_18856,N_16255);
nand U21283 (N_21283,N_19629,N_17608);
nor U21284 (N_21284,N_19643,N_17096);
nand U21285 (N_21285,N_19199,N_17061);
nor U21286 (N_21286,N_15973,N_15570);
nand U21287 (N_21287,N_16963,N_19465);
nor U21288 (N_21288,N_17270,N_19010);
xor U21289 (N_21289,N_16351,N_16698);
and U21290 (N_21290,N_15562,N_18813);
nor U21291 (N_21291,N_17837,N_16746);
and U21292 (N_21292,N_15966,N_17016);
and U21293 (N_21293,N_16812,N_15942);
or U21294 (N_21294,N_18677,N_18342);
and U21295 (N_21295,N_16068,N_17326);
nor U21296 (N_21296,N_18132,N_18558);
nand U21297 (N_21297,N_19047,N_19280);
xor U21298 (N_21298,N_15555,N_17866);
xor U21299 (N_21299,N_15531,N_18098);
nor U21300 (N_21300,N_18775,N_17433);
nor U21301 (N_21301,N_16760,N_18437);
and U21302 (N_21302,N_16441,N_17384);
xor U21303 (N_21303,N_17486,N_16931);
or U21304 (N_21304,N_16712,N_15550);
nor U21305 (N_21305,N_15960,N_17693);
or U21306 (N_21306,N_17893,N_17145);
nor U21307 (N_21307,N_17111,N_17979);
or U21308 (N_21308,N_18599,N_16329);
or U21309 (N_21309,N_15540,N_16229);
or U21310 (N_21310,N_18882,N_18310);
nor U21311 (N_21311,N_17184,N_19948);
or U21312 (N_21312,N_16622,N_18720);
nand U21313 (N_21313,N_16385,N_15813);
nor U21314 (N_21314,N_15538,N_18516);
nand U21315 (N_21315,N_16040,N_16768);
nor U21316 (N_21316,N_19167,N_16546);
nand U21317 (N_21317,N_18471,N_16547);
nor U21318 (N_21318,N_16909,N_17785);
and U21319 (N_21319,N_19479,N_19179);
or U21320 (N_21320,N_15048,N_19863);
nor U21321 (N_21321,N_18712,N_15662);
nor U21322 (N_21322,N_19476,N_17488);
xnor U21323 (N_21323,N_19502,N_15355);
or U21324 (N_21324,N_19551,N_17079);
nand U21325 (N_21325,N_15510,N_16110);
and U21326 (N_21326,N_18414,N_19451);
xor U21327 (N_21327,N_17867,N_16007);
and U21328 (N_21328,N_19371,N_19053);
and U21329 (N_21329,N_19032,N_16717);
or U21330 (N_21330,N_19646,N_19595);
and U21331 (N_21331,N_16317,N_19690);
nand U21332 (N_21332,N_15066,N_18173);
or U21333 (N_21333,N_17528,N_18887);
xor U21334 (N_21334,N_16301,N_17077);
xnor U21335 (N_21335,N_15886,N_17735);
nand U21336 (N_21336,N_17684,N_17887);
and U21337 (N_21337,N_16036,N_18255);
nor U21338 (N_21338,N_18884,N_19661);
nor U21339 (N_21339,N_18731,N_16947);
and U21340 (N_21340,N_16250,N_18547);
or U21341 (N_21341,N_18174,N_18386);
and U21342 (N_21342,N_15113,N_18985);
nor U21343 (N_21343,N_16293,N_17699);
or U21344 (N_21344,N_17956,N_18004);
and U21345 (N_21345,N_18368,N_15741);
and U21346 (N_21346,N_19437,N_15350);
or U21347 (N_21347,N_17335,N_17662);
or U21348 (N_21348,N_17092,N_19153);
nand U21349 (N_21349,N_18401,N_19559);
and U21350 (N_21350,N_16473,N_19734);
nor U21351 (N_21351,N_16802,N_17748);
xnor U21352 (N_21352,N_18078,N_19666);
or U21353 (N_21353,N_17062,N_17440);
xor U21354 (N_21354,N_17504,N_16625);
nor U21355 (N_21355,N_19470,N_16300);
and U21356 (N_21356,N_17108,N_16542);
and U21357 (N_21357,N_16114,N_16488);
nor U21358 (N_21358,N_17140,N_16704);
and U21359 (N_21359,N_16520,N_18076);
and U21360 (N_21360,N_15468,N_18305);
xor U21361 (N_21361,N_17039,N_17656);
and U21362 (N_21362,N_15970,N_19366);
nand U21363 (N_21363,N_19263,N_16020);
nor U21364 (N_21364,N_19190,N_18458);
xnor U21365 (N_21365,N_17341,N_18969);
nand U21366 (N_21366,N_17587,N_17721);
nand U21367 (N_21367,N_16729,N_19855);
nand U21368 (N_21368,N_16126,N_19257);
or U21369 (N_21369,N_16792,N_15638);
or U21370 (N_21370,N_18834,N_16256);
or U21371 (N_21371,N_15404,N_17491);
or U21372 (N_21372,N_18913,N_15311);
nand U21373 (N_21373,N_18788,N_16910);
nand U21374 (N_21374,N_17904,N_15147);
nor U21375 (N_21375,N_16054,N_17192);
nand U21376 (N_21376,N_19463,N_19462);
xor U21377 (N_21377,N_16121,N_17909);
nand U21378 (N_21378,N_18465,N_18837);
and U21379 (N_21379,N_16887,N_18651);
nand U21380 (N_21380,N_16476,N_15354);
and U21381 (N_21381,N_16876,N_18555);
xnor U21382 (N_21382,N_16071,N_19640);
nor U21383 (N_21383,N_17119,N_19325);
and U21384 (N_21384,N_15117,N_17415);
nand U21385 (N_21385,N_17553,N_17318);
nand U21386 (N_21386,N_18445,N_17098);
and U21387 (N_21387,N_18311,N_19717);
nand U21388 (N_21388,N_15711,N_18966);
or U21389 (N_21389,N_17991,N_15627);
nor U21390 (N_21390,N_17709,N_19211);
and U21391 (N_21391,N_16706,N_18971);
and U21392 (N_21392,N_17523,N_19123);
and U21393 (N_21393,N_15866,N_15892);
nand U21394 (N_21394,N_17289,N_15828);
nor U21395 (N_21395,N_15707,N_16215);
and U21396 (N_21396,N_16504,N_15470);
nand U21397 (N_21397,N_17988,N_18878);
nor U21398 (N_21398,N_19924,N_15461);
and U21399 (N_21399,N_16908,N_19128);
nand U21400 (N_21400,N_18979,N_15087);
and U21401 (N_21401,N_15628,N_18472);
nand U21402 (N_21402,N_18405,N_16092);
and U21403 (N_21403,N_16398,N_18860);
or U21404 (N_21404,N_16900,N_19293);
or U21405 (N_21405,N_16478,N_16049);
nor U21406 (N_21406,N_16075,N_18635);
nand U21407 (N_21407,N_15387,N_16514);
nand U21408 (N_21408,N_17385,N_19700);
and U21409 (N_21409,N_19489,N_16035);
nand U21410 (N_21410,N_15592,N_18259);
nand U21411 (N_21411,N_18102,N_19192);
and U21412 (N_21412,N_18434,N_19346);
or U21413 (N_21413,N_18474,N_17941);
or U21414 (N_21414,N_15042,N_19931);
nand U21415 (N_21415,N_17067,N_19771);
or U21416 (N_21416,N_19772,N_19279);
nor U21417 (N_21417,N_17327,N_18235);
and U21418 (N_21418,N_16246,N_18495);
nand U21419 (N_21419,N_19678,N_16856);
nor U21420 (N_21420,N_16325,N_15755);
and U21421 (N_21421,N_16601,N_15254);
nor U21422 (N_21422,N_19330,N_17818);
or U21423 (N_21423,N_17634,N_15083);
nor U21424 (N_21424,N_15768,N_16674);
nor U21425 (N_21425,N_18627,N_16238);
nand U21426 (N_21426,N_15776,N_15831);
nand U21427 (N_21427,N_19667,N_16801);
and U21428 (N_21428,N_18565,N_19447);
and U21429 (N_21429,N_18055,N_15943);
xor U21430 (N_21430,N_16127,N_15979);
and U21431 (N_21431,N_15744,N_15088);
or U21432 (N_21432,N_19297,N_17770);
or U21433 (N_21433,N_18747,N_15723);
nor U21434 (N_21434,N_19560,N_18309);
nor U21435 (N_21435,N_19981,N_16505);
or U21436 (N_21436,N_18273,N_19975);
nand U21437 (N_21437,N_17057,N_16818);
nor U21438 (N_21438,N_18162,N_18229);
nand U21439 (N_21439,N_16911,N_19028);
nor U21440 (N_21440,N_15725,N_16882);
nand U21441 (N_21441,N_17830,N_19526);
or U21442 (N_21442,N_17153,N_15530);
nand U21443 (N_21443,N_15746,N_17936);
or U21444 (N_21444,N_18716,N_19288);
and U21445 (N_21445,N_18080,N_19425);
and U21446 (N_21446,N_17342,N_16635);
nor U21447 (N_21447,N_19369,N_18283);
nor U21448 (N_21448,N_16268,N_16498);
nor U21449 (N_21449,N_17428,N_19615);
nand U21450 (N_21450,N_19232,N_18204);
or U21451 (N_21451,N_19247,N_17058);
nor U21452 (N_21452,N_18250,N_18502);
nand U21453 (N_21453,N_19362,N_19074);
xor U21454 (N_21454,N_19103,N_18017);
nand U21455 (N_21455,N_17094,N_16455);
nand U21456 (N_21456,N_17238,N_15224);
nand U21457 (N_21457,N_19360,N_16296);
or U21458 (N_21458,N_16227,N_19134);
nand U21459 (N_21459,N_17193,N_18160);
and U21460 (N_21460,N_15315,N_18988);
nor U21461 (N_21461,N_15193,N_18993);
nor U21462 (N_21462,N_19000,N_18013);
and U21463 (N_21463,N_17222,N_18105);
nand U21464 (N_21464,N_15900,N_17100);
nand U21465 (N_21465,N_15954,N_16939);
nand U21466 (N_21466,N_18823,N_15683);
or U21467 (N_21467,N_18033,N_19340);
and U21468 (N_21468,N_16043,N_18526);
nor U21469 (N_21469,N_15416,N_19574);
nor U21470 (N_21470,N_15180,N_17642);
or U21471 (N_21471,N_15091,N_17678);
nand U21472 (N_21472,N_15596,N_16552);
nand U21473 (N_21473,N_16189,N_19965);
nand U21474 (N_21474,N_19903,N_17036);
nor U21475 (N_21475,N_16791,N_18297);
or U21476 (N_21476,N_18895,N_15132);
or U21477 (N_21477,N_16285,N_19959);
and U21478 (N_21478,N_18815,N_17813);
nand U21479 (N_21479,N_17449,N_15377);
nand U21480 (N_21480,N_18395,N_18468);
nor U21481 (N_21481,N_15955,N_18835);
or U21482 (N_21482,N_18869,N_16399);
nand U21483 (N_21483,N_15762,N_15196);
and U21484 (N_21484,N_16457,N_19149);
nand U21485 (N_21485,N_17808,N_17633);
nor U21486 (N_21486,N_19859,N_18632);
or U21487 (N_21487,N_18141,N_18254);
and U21488 (N_21488,N_17035,N_18104);
nand U21489 (N_21489,N_17175,N_15444);
nand U21490 (N_21490,N_17895,N_19117);
and U21491 (N_21491,N_18396,N_17926);
nor U21492 (N_21492,N_16240,N_15719);
nor U21493 (N_21493,N_19252,N_15789);
nand U21494 (N_21494,N_15293,N_17001);
or U21495 (N_21495,N_19916,N_16466);
or U21496 (N_21496,N_18995,N_19083);
or U21497 (N_21497,N_19108,N_19562);
nor U21498 (N_21498,N_19762,N_19569);
nand U21499 (N_21499,N_16654,N_15870);
xnor U21500 (N_21500,N_17792,N_15962);
nand U21501 (N_21501,N_19811,N_17084);
nand U21502 (N_21502,N_17427,N_16656);
and U21503 (N_21503,N_17975,N_18245);
xnor U21504 (N_21504,N_17240,N_15388);
nor U21505 (N_21505,N_19584,N_19817);
nor U21506 (N_21506,N_16231,N_15618);
xor U21507 (N_21507,N_17466,N_16269);
nor U21508 (N_21508,N_15327,N_17152);
nand U21509 (N_21509,N_19672,N_15721);
and U21510 (N_21510,N_18886,N_19239);
or U21511 (N_21511,N_19856,N_19763);
nand U21512 (N_21512,N_16433,N_15324);
and U21513 (N_21513,N_19731,N_16029);
or U21514 (N_21514,N_17703,N_18088);
nor U21515 (N_21515,N_16266,N_19711);
or U21516 (N_21516,N_19778,N_17570);
nor U21517 (N_21517,N_19291,N_19415);
nor U21518 (N_21518,N_15537,N_18517);
nor U21519 (N_21519,N_18372,N_16661);
nand U21520 (N_21520,N_17000,N_16653);
and U21521 (N_21521,N_17172,N_18428);
nor U21522 (N_21522,N_19412,N_19878);
nand U21523 (N_21523,N_15527,N_18955);
nor U21524 (N_21524,N_17429,N_15770);
and U21525 (N_21525,N_16554,N_17751);
nand U21526 (N_21526,N_16444,N_17306);
or U21527 (N_21527,N_17278,N_17225);
or U21528 (N_21528,N_18615,N_18773);
or U21529 (N_21529,N_15121,N_18171);
xnor U21530 (N_21530,N_15166,N_16859);
nand U21531 (N_21531,N_18586,N_19626);
and U21532 (N_21532,N_16784,N_19896);
nand U21533 (N_21533,N_16957,N_17903);
or U21534 (N_21534,N_19262,N_19019);
nand U21535 (N_21535,N_19122,N_19094);
and U21536 (N_21536,N_15045,N_19597);
and U21537 (N_21537,N_19841,N_18137);
and U21538 (N_21538,N_17367,N_19761);
nor U21539 (N_21539,N_19994,N_17339);
nor U21540 (N_21540,N_16044,N_17790);
and U21541 (N_21541,N_19014,N_18177);
or U21542 (N_21542,N_16696,N_17373);
nand U21543 (N_21543,N_18513,N_15859);
and U21544 (N_21544,N_17352,N_19593);
or U21545 (N_21545,N_17332,N_16726);
or U21546 (N_21546,N_17217,N_15021);
or U21547 (N_21547,N_16259,N_17517);
nand U21548 (N_21548,N_17246,N_19550);
nand U21549 (N_21549,N_19403,N_18491);
xnor U21550 (N_21550,N_15442,N_19984);
and U21551 (N_21551,N_15347,N_18764);
and U21552 (N_21552,N_16471,N_18714);
nand U21553 (N_21553,N_17164,N_17279);
or U21554 (N_21554,N_17692,N_15930);
or U21555 (N_21555,N_17680,N_15999);
xor U21556 (N_21556,N_17676,N_17455);
or U21557 (N_21557,N_19121,N_17382);
or U21558 (N_21558,N_15967,N_18843);
or U21559 (N_21559,N_16745,N_18048);
and U21560 (N_21560,N_15450,N_16469);
nand U21561 (N_21561,N_15403,N_18962);
nand U21562 (N_21562,N_16511,N_15919);
nor U21563 (N_21563,N_18858,N_18214);
or U21564 (N_21564,N_16343,N_15292);
xor U21565 (N_21565,N_17408,N_15360);
and U21566 (N_21566,N_15907,N_15453);
and U21567 (N_21567,N_19033,N_19852);
nand U21568 (N_21568,N_17541,N_17764);
or U21569 (N_21569,N_19375,N_19662);
or U21570 (N_21570,N_16201,N_16265);
nand U21571 (N_21571,N_18444,N_16183);
xnor U21572 (N_21572,N_18286,N_19842);
and U21573 (N_21573,N_19444,N_16734);
nor U21574 (N_21574,N_18448,N_19443);
and U21575 (N_21575,N_18207,N_19458);
and U21576 (N_21576,N_16503,N_16789);
or U21577 (N_21577,N_16508,N_15156);
nand U21578 (N_21578,N_18999,N_17525);
nor U21579 (N_21579,N_16388,N_17040);
or U21580 (N_21580,N_16814,N_15715);
nand U21581 (N_21581,N_17752,N_19663);
xor U21582 (N_21582,N_15858,N_18279);
and U21583 (N_21583,N_15578,N_15511);
and U21584 (N_21584,N_18089,N_17954);
and U21585 (N_21585,N_18709,N_17116);
nand U21586 (N_21586,N_19383,N_15123);
nand U21587 (N_21587,N_15222,N_15856);
nor U21588 (N_21588,N_19801,N_19082);
nor U21589 (N_21589,N_16907,N_15750);
or U21590 (N_21590,N_18261,N_16845);
or U21591 (N_21591,N_16342,N_17404);
or U21592 (N_21592,N_18400,N_17106);
and U21593 (N_21593,N_19286,N_19524);
nand U21594 (N_21594,N_16865,N_16005);
nand U21595 (N_21595,N_15229,N_16434);
nand U21596 (N_21596,N_16928,N_17694);
or U21597 (N_21597,N_17598,N_18559);
and U21598 (N_21598,N_15940,N_17707);
nor U21599 (N_21599,N_17540,N_16994);
or U21600 (N_21600,N_15460,N_17505);
xnor U21601 (N_21601,N_18594,N_17860);
or U21602 (N_21602,N_17249,N_17664);
nand U21603 (N_21603,N_17188,N_18736);
nand U21604 (N_21604,N_18571,N_18267);
nor U21605 (N_21605,N_17060,N_18488);
and U21606 (N_21606,N_16590,N_15289);
nor U21607 (N_21607,N_17864,N_16872);
and U21608 (N_21608,N_19273,N_16211);
nor U21609 (N_21609,N_15685,N_15819);
or U21610 (N_21610,N_16506,N_15644);
and U21611 (N_21611,N_15710,N_16161);
nor U21612 (N_21612,N_17462,N_18085);
and U21613 (N_21613,N_17065,N_17399);
nor U21614 (N_21614,N_18910,N_15790);
nor U21615 (N_21615,N_18883,N_16191);
or U21616 (N_21616,N_19824,N_17901);
and U21617 (N_21617,N_18784,N_19874);
nor U21618 (N_21618,N_15545,N_16854);
and U21619 (N_21619,N_17648,N_17730);
xnor U21620 (N_21620,N_17469,N_19281);
and U21621 (N_21621,N_16323,N_19256);
nor U21622 (N_21622,N_19862,N_16375);
and U21623 (N_21623,N_15421,N_19316);
nor U21624 (N_21624,N_15357,N_19289);
nor U21625 (N_21625,N_15462,N_16972);
or U21626 (N_21626,N_19654,N_18649);
xnor U21627 (N_21627,N_19109,N_17771);
nor U21628 (N_21628,N_15384,N_16057);
nand U21629 (N_21629,N_18347,N_18648);
nor U21630 (N_21630,N_19114,N_15684);
nor U21631 (N_21631,N_19243,N_19237);
or U21632 (N_21632,N_18417,N_17580);
or U21633 (N_21633,N_15512,N_16151);
nand U21634 (N_21634,N_18130,N_15368);
or U21635 (N_21635,N_16042,N_16534);
nand U21636 (N_21636,N_17925,N_15743);
nor U21637 (N_21637,N_16641,N_19937);
nand U21638 (N_21638,N_17971,N_15137);
xor U21639 (N_21639,N_15143,N_15524);
or U21640 (N_21640,N_15307,N_18838);
or U21641 (N_21641,N_19373,N_16244);
and U21642 (N_21642,N_19829,N_16893);
and U21643 (N_21643,N_15899,N_17573);
or U21644 (N_21644,N_18007,N_19183);
or U21645 (N_21645,N_19342,N_16889);
or U21646 (N_21646,N_19596,N_19642);
nor U21647 (N_21647,N_15591,N_18892);
and U21648 (N_21648,N_16718,N_18967);
and U21649 (N_21649,N_18846,N_16278);
or U21650 (N_21650,N_15593,N_19676);
and U21651 (N_21651,N_17876,N_15363);
nand U21652 (N_21652,N_16027,N_18818);
nand U21653 (N_21653,N_19424,N_19517);
or U21654 (N_21654,N_15158,N_17196);
and U21655 (N_21655,N_16146,N_16170);
nand U21656 (N_21656,N_18992,N_19637);
and U21657 (N_21657,N_17496,N_19359);
nand U21658 (N_21658,N_17995,N_16999);
and U21659 (N_21659,N_16751,N_16445);
nand U21660 (N_21660,N_17884,N_15853);
nor U21661 (N_21661,N_19494,N_18996);
and U21662 (N_21662,N_19561,N_16394);
nor U21663 (N_21663,N_17485,N_19460);
nand U21664 (N_21664,N_16591,N_15099);
or U21665 (N_21665,N_15452,N_19812);
or U21666 (N_21666,N_17456,N_17708);
nand U21667 (N_21667,N_15303,N_19449);
nand U21668 (N_21668,N_16406,N_16537);
nor U21669 (N_21669,N_16233,N_16416);
or U21670 (N_21670,N_16982,N_18119);
or U21671 (N_21671,N_15131,N_19922);
nand U21672 (N_21672,N_17200,N_18051);
or U21673 (N_21673,N_19659,N_15092);
nand U21674 (N_21674,N_19246,N_16927);
nand U21675 (N_21675,N_15498,N_15389);
and U21676 (N_21676,N_19498,N_15126);
xnor U21677 (N_21677,N_15146,N_17210);
nand U21678 (N_21678,N_19723,N_16137);
and U21679 (N_21679,N_15772,N_18202);
or U21680 (N_21680,N_19154,N_15778);
nor U21681 (N_21681,N_17180,N_17233);
xnor U21682 (N_21682,N_17069,N_18529);
or U21683 (N_21683,N_19973,N_18336);
or U21684 (N_21684,N_18921,N_16613);
nand U21685 (N_21685,N_15310,N_15816);
or U21686 (N_21686,N_17048,N_19789);
and U21687 (N_21687,N_19623,N_19035);
nand U21688 (N_21688,N_19583,N_18270);
and U21689 (N_21689,N_15924,N_16037);
nor U21690 (N_21690,N_16361,N_19819);
nor U21691 (N_21691,N_17023,N_17848);
and U21692 (N_21692,N_15936,N_15346);
or U21693 (N_21693,N_17780,N_15049);
and U21694 (N_21694,N_19140,N_15880);
or U21695 (N_21695,N_18984,N_18374);
or U21696 (N_21696,N_16747,N_17198);
nand U21697 (N_21697,N_18455,N_17574);
xor U21698 (N_21698,N_19050,N_17781);
or U21699 (N_21699,N_18290,N_17158);
nand U21700 (N_21700,N_18540,N_17921);
nor U21701 (N_21701,N_15922,N_16849);
nand U21702 (N_21702,N_17337,N_19469);
nor U21703 (N_21703,N_19015,N_18260);
nor U21704 (N_21704,N_18827,N_19116);
xnor U21705 (N_21705,N_19759,N_19634);
nor U21706 (N_21706,N_18147,N_19950);
and U21707 (N_21707,N_15473,N_16817);
nand U21708 (N_21708,N_18692,N_15133);
or U21709 (N_21709,N_19624,N_17348);
nand U21710 (N_21710,N_15594,N_18028);
nand U21711 (N_21711,N_15885,N_15398);
nor U21712 (N_21712,N_15670,N_19113);
or U21713 (N_21713,N_16874,N_19650);
xor U21714 (N_21714,N_17127,N_15268);
and U21715 (N_21715,N_18026,N_17423);
nor U21716 (N_21716,N_18435,N_17597);
nor U21717 (N_21717,N_16459,N_15681);
nand U21718 (N_21718,N_18186,N_15873);
nand U21719 (N_21719,N_17114,N_16297);
xor U21720 (N_21720,N_16976,N_19851);
nor U21721 (N_21721,N_16340,N_16221);
or U21722 (N_21722,N_19493,N_16553);
nand U21723 (N_21723,N_19215,N_19732);
nand U21724 (N_21724,N_18840,N_19442);
and U21725 (N_21725,N_19740,N_15325);
or U21726 (N_21726,N_17558,N_16094);
nand U21727 (N_21727,N_15400,N_19137);
or U21728 (N_21728,N_15205,N_19655);
or U21729 (N_21729,N_15840,N_15007);
nor U21730 (N_21730,N_17614,N_16116);
nand U21731 (N_21731,N_15247,N_17750);
or U21732 (N_21732,N_17674,N_18057);
nor U21733 (N_21733,N_19065,N_19464);
and U21734 (N_21734,N_17304,N_19808);
or U21735 (N_21735,N_17706,N_16011);
nand U21736 (N_21736,N_18645,N_15614);
nor U21737 (N_21737,N_19361,N_19913);
and U21738 (N_21738,N_15526,N_19906);
nand U21739 (N_21739,N_19548,N_18263);
xnor U21740 (N_21740,N_18751,N_19688);
nand U21741 (N_21741,N_19323,N_16685);
and U21742 (N_21742,N_16341,N_15584);
or U21743 (N_21743,N_19912,N_19097);
or U21744 (N_21744,N_18024,N_17536);
nand U21745 (N_21745,N_19206,N_15044);
and U21746 (N_21746,N_18121,N_17470);
nor U21747 (N_21747,N_19742,N_18325);
and U21748 (N_21748,N_18744,N_16452);
and U21749 (N_21749,N_18200,N_17053);
nor U21750 (N_21750,N_16055,N_19429);
nand U21751 (N_21751,N_16322,N_19124);
nor U21752 (N_21752,N_16028,N_18034);
or U21753 (N_21753,N_17501,N_16535);
or U21754 (N_21754,N_18252,N_17617);
nor U21755 (N_21755,N_16920,N_17045);
nand U21756 (N_21756,N_19825,N_15698);
nor U21757 (N_21757,N_16379,N_19671);
and U21758 (N_21758,N_16249,N_16402);
and U21759 (N_21759,N_19016,N_18584);
or U21760 (N_21760,N_18569,N_18268);
nand U21761 (N_21761,N_18014,N_19002);
nor U21762 (N_21762,N_19210,N_16163);
and U21763 (N_21763,N_17117,N_19692);
and U21764 (N_21764,N_17538,N_16822);
xor U21765 (N_21765,N_19735,N_18998);
or U21766 (N_21766,N_17512,N_15372);
or U21767 (N_21767,N_15073,N_18619);
and U21768 (N_21768,N_17646,N_18568);
nand U21769 (N_21769,N_19616,N_16194);
nand U21770 (N_21770,N_17990,N_15208);
nor U21771 (N_21771,N_17224,N_16432);
and U21772 (N_21772,N_16378,N_15998);
nand U21773 (N_21773,N_17732,N_15331);
xnor U21774 (N_21774,N_18839,N_19151);
or U21775 (N_21775,N_18637,N_17274);
nand U21776 (N_21776,N_17788,N_16119);
xor U21777 (N_21777,N_15019,N_18574);
nor U21778 (N_21778,N_16263,N_19967);
or U21779 (N_21779,N_16039,N_18857);
or U21780 (N_21780,N_17281,N_19705);
nor U21781 (N_21781,N_18663,N_19382);
nor U21782 (N_21782,N_15413,N_15214);
nor U21783 (N_21783,N_15872,N_17242);
nor U21784 (N_21784,N_17513,N_15297);
and U21785 (N_21785,N_17632,N_15445);
nor U21786 (N_21786,N_19405,N_16997);
nor U21787 (N_21787,N_18991,N_16510);
nor U21788 (N_21788,N_18760,N_19238);
nor U21789 (N_21789,N_15532,N_19565);
and U21790 (N_21790,N_16842,N_18404);
nand U21791 (N_21791,N_17331,N_16493);
or U21792 (N_21792,N_15219,N_19834);
nor U21793 (N_21793,N_17284,N_15266);
and U21794 (N_21794,N_19553,N_16813);
or U21795 (N_21795,N_16811,N_19499);
xnor U21796 (N_21796,N_15579,N_17197);
and U21797 (N_21797,N_17252,N_19590);
or U21798 (N_21798,N_15896,N_15435);
and U21799 (N_21799,N_18503,N_15058);
or U21800 (N_21800,N_19687,N_16898);
nor U21801 (N_21801,N_19056,N_16424);
or U21802 (N_21802,N_17660,N_19701);
xnor U21803 (N_21803,N_18225,N_15220);
or U21804 (N_21804,N_18454,N_18951);
nor U21805 (N_21805,N_15269,N_19321);
nor U21806 (N_21806,N_19698,N_17739);
nor U21807 (N_21807,N_16101,N_17334);
nand U21808 (N_21808,N_17467,N_15221);
nand U21809 (N_21809,N_17844,N_15845);
xnor U21810 (N_21810,N_16608,N_16442);
nand U21811 (N_21811,N_18605,N_16307);
xor U21812 (N_21812,N_17560,N_17978);
and U21813 (N_21813,N_15603,N_19621);
nand U21814 (N_21814,N_16218,N_18349);
and U21815 (N_21815,N_15420,N_18253);
nand U21816 (N_21816,N_17937,N_15031);
nand U21817 (N_21817,N_17945,N_19488);
nand U21818 (N_21818,N_18796,N_15713);
and U21819 (N_21819,N_17125,N_17265);
nand U21820 (N_21820,N_15304,N_15517);
or U21821 (N_21821,N_15585,N_18041);
nand U21822 (N_21822,N_15576,N_16403);
or U21823 (N_21823,N_19490,N_16778);
xor U21824 (N_21824,N_15027,N_16647);
and U21825 (N_21825,N_15237,N_17137);
xor U21826 (N_21826,N_15407,N_18338);
or U21827 (N_21827,N_18908,N_17929);
and U21828 (N_21828,N_18090,N_19202);
xnor U21829 (N_21829,N_15185,N_17930);
nand U21830 (N_21830,N_17524,N_19282);
or U21831 (N_21831,N_16699,N_17629);
or U21832 (N_21832,N_15502,N_15587);
or U21833 (N_21833,N_17025,N_15923);
nor U21834 (N_21834,N_18917,N_18185);
nand U21835 (N_21835,N_15145,N_15830);
nand U21836 (N_21836,N_19253,N_19781);
or U21837 (N_21837,N_15463,N_16823);
and U21838 (N_21838,N_19209,N_16985);
nand U21839 (N_21839,N_18019,N_18667);
and U21840 (N_21840,N_17139,N_19739);
nor U21841 (N_21841,N_18318,N_19131);
nand U21842 (N_21842,N_15509,N_19261);
xnor U21843 (N_21843,N_16716,N_17981);
and U21844 (N_21844,N_15583,N_19013);
or U21845 (N_21845,N_15916,N_17028);
nand U21846 (N_21846,N_16536,N_16638);
and U21847 (N_21847,N_16765,N_15203);
xnor U21848 (N_21848,N_15236,N_16438);
nand U21849 (N_21849,N_17487,N_18679);
and U21850 (N_21850,N_17840,N_18557);
and U21851 (N_21851,N_18046,N_16578);
nand U21852 (N_21852,N_15565,N_16549);
or U21853 (N_21853,N_16414,N_19598);
or U21854 (N_21854,N_16728,N_18332);
nand U21855 (N_21855,N_17856,N_19904);
and U21856 (N_21856,N_17170,N_15401);
or U21857 (N_21857,N_15932,N_19633);
nand U21858 (N_21858,N_15177,N_18330);
or U21859 (N_21859,N_19182,N_17343);
and U21860 (N_21860,N_19030,N_16111);
and U21861 (N_21861,N_16815,N_15075);
and U21862 (N_21862,N_16006,N_19348);
or U21863 (N_21863,N_16626,N_16041);
nand U21864 (N_21864,N_17966,N_19923);
xor U21865 (N_21865,N_16754,N_18094);
and U21866 (N_21866,N_18623,N_19558);
or U21867 (N_21867,N_15440,N_18329);
nor U21868 (N_21868,N_16273,N_16456);
or U21869 (N_21869,N_18487,N_19057);
and U21870 (N_21870,N_18535,N_17763);
nand U21871 (N_21871,N_18520,N_17353);
nor U21872 (N_21872,N_17624,N_15217);
nand U21873 (N_21873,N_18670,N_19543);
or U21874 (N_21874,N_15601,N_16247);
and U21875 (N_21875,N_15852,N_18938);
nor U21876 (N_21876,N_19060,N_18864);
and U21877 (N_21877,N_15197,N_17497);
or U21878 (N_21878,N_16251,N_15528);
or U21879 (N_21879,N_19226,N_16408);
nor U21880 (N_21880,N_15284,N_17163);
nor U21881 (N_21881,N_15981,N_15397);
or U21882 (N_21882,N_19619,N_17786);
nor U21883 (N_21883,N_15294,N_15061);
or U21884 (N_21884,N_16531,N_18384);
or U21885 (N_21885,N_16663,N_16890);
and U21886 (N_21886,N_17323,N_16377);
or U21887 (N_21887,N_19336,N_18865);
nor U21888 (N_21888,N_16487,N_18694);
nand U21889 (N_21889,N_19986,N_17239);
nor U21890 (N_21890,N_16929,N_19887);
and U21891 (N_21891,N_15153,N_18193);
and U21892 (N_21892,N_19135,N_15917);
nand U21893 (N_21893,N_18739,N_17885);
nand U21894 (N_21894,N_17556,N_19038);
and U21895 (N_21895,N_19519,N_19980);
nor U21896 (N_21896,N_16582,N_18874);
nor U21897 (N_21897,N_15317,N_18851);
nor U21898 (N_21898,N_15176,N_15393);
nor U21899 (N_21899,N_18230,N_15781);
xor U21900 (N_21900,N_16619,N_19725);
nor U21901 (N_21901,N_19810,N_18391);
or U21902 (N_21902,N_18106,N_19767);
or U21903 (N_21903,N_19018,N_15648);
nor U21904 (N_21904,N_19884,N_16492);
and U21905 (N_21905,N_16230,N_15615);
and U21906 (N_21906,N_19528,N_19748);
nand U21907 (N_21907,N_18612,N_19848);
or U21908 (N_21908,N_19788,N_15459);
and U21909 (N_21909,N_17086,N_15607);
nand U21910 (N_21910,N_15480,N_18352);
and U21911 (N_21911,N_15982,N_16589);
and U21912 (N_21912,N_15543,N_18911);
xnor U21913 (N_21913,N_17851,N_17014);
nor U21914 (N_21914,N_15161,N_16008);
or U21915 (N_21915,N_17765,N_17480);
and U21916 (N_21916,N_18929,N_18582);
nor U21917 (N_21917,N_17733,N_19394);
and U21918 (N_21918,N_17506,N_18484);
nand U21919 (N_21919,N_18898,N_17229);
nor U21920 (N_21920,N_18845,N_18462);
nand U21921 (N_21921,N_16667,N_16105);
or U21922 (N_21922,N_15067,N_19505);
xor U21923 (N_21923,N_17507,N_16752);
or U21924 (N_21924,N_19365,N_16420);
xnor U21925 (N_21925,N_18319,N_19792);
nor U21926 (N_21926,N_16679,N_16216);
and U21927 (N_21927,N_19376,N_16298);
nand U21928 (N_21928,N_18765,N_19603);
and U21929 (N_21929,N_16491,N_15285);
nand U21930 (N_21930,N_15669,N_16384);
nor U21931 (N_21931,N_19177,N_18483);
and U21932 (N_21932,N_18146,N_17701);
nor U21933 (N_21933,N_15632,N_18344);
and U21934 (N_21934,N_16722,N_17626);
nor U21935 (N_21935,N_17783,N_18074);
and U21936 (N_21936,N_17244,N_19968);
or U21937 (N_21937,N_15383,N_18324);
nand U21938 (N_21938,N_15560,N_19349);
nand U21939 (N_21939,N_18269,N_17260);
nor U21940 (N_21940,N_19450,N_15082);
nand U21941 (N_21941,N_19750,N_16677);
nand U21942 (N_21942,N_18058,N_19760);
or U21943 (N_21943,N_19328,N_17858);
and U21944 (N_21944,N_19636,N_17907);
and U21945 (N_21945,N_15104,N_15838);
nand U21946 (N_21946,N_16460,N_18370);
or U21947 (N_21947,N_16474,N_19404);
or U21948 (N_21948,N_15050,N_17107);
nor U21949 (N_21949,N_18001,N_18610);
and U21950 (N_21950,N_17546,N_16525);
nor U21951 (N_21951,N_18415,N_16381);
nor U21952 (N_21952,N_18083,N_18762);
or U21953 (N_21953,N_15441,N_18308);
nand U21954 (N_21954,N_16609,N_17511);
nor U21955 (N_21955,N_19776,N_15659);
and U21956 (N_21956,N_19940,N_19345);
nand U21957 (N_21957,N_15868,N_18521);
or U21958 (N_21958,N_16393,N_16108);
or U21959 (N_21959,N_17294,N_18646);
and U21960 (N_21960,N_18341,N_19601);
or U21961 (N_21961,N_16964,N_17303);
nor U21962 (N_21962,N_18790,N_18717);
nand U21963 (N_21963,N_16773,N_16072);
nand U21964 (N_21964,N_19380,N_16727);
nor U21965 (N_21965,N_17772,N_15106);
nor U21966 (N_21966,N_19849,N_16334);
and U21967 (N_21967,N_17833,N_18143);
nor U21968 (N_21968,N_17865,N_18180);
xor U21969 (N_21969,N_15053,N_16390);
or U21970 (N_21970,N_16797,N_19729);
or U21971 (N_21971,N_18205,N_15065);
nand U21972 (N_21972,N_19020,N_17702);
or U21973 (N_21973,N_19813,N_18302);
nor U21974 (N_21974,N_18561,N_15190);
or U21975 (N_21975,N_17417,N_19614);
nand U21976 (N_21976,N_15192,N_19744);
and U21977 (N_21977,N_16339,N_15804);
nor U21978 (N_21978,N_15571,N_16990);
or U21979 (N_21979,N_18501,N_16916);
nand U21980 (N_21980,N_18506,N_15476);
xnor U21981 (N_21981,N_19381,N_18602);
or U21982 (N_21982,N_17890,N_15472);
nand U21983 (N_21983,N_16847,N_15225);
or U21984 (N_21984,N_17589,N_16866);
nor U21985 (N_21985,N_16615,N_19269);
nor U21986 (N_21986,N_19879,N_18972);
nand U21987 (N_21987,N_17250,N_15371);
nand U21988 (N_21988,N_15732,N_16053);
or U21989 (N_21989,N_15267,N_16303);
or U21990 (N_21990,N_16328,N_15696);
nor U21991 (N_21991,N_19051,N_19037);
and U21992 (N_21992,N_17264,N_15437);
nor U21993 (N_21993,N_19421,N_17836);
or U21994 (N_21994,N_18534,N_18379);
nand U21995 (N_21995,N_16440,N_17231);
or U21996 (N_21996,N_15529,N_15163);
nand U21997 (N_21997,N_17611,N_15904);
nor U21998 (N_21998,N_19695,N_19714);
xnor U21999 (N_21999,N_15754,N_17719);
or U22000 (N_22000,N_19313,N_18140);
xnor U22001 (N_22001,N_18062,N_19070);
and U22002 (N_22002,N_16723,N_17412);
xnor U22003 (N_22003,N_16120,N_19694);
or U22004 (N_22004,N_16302,N_18211);
nand U22005 (N_22005,N_17024,N_19283);
and U22006 (N_22006,N_15273,N_16761);
nand U22007 (N_22007,N_15035,N_15846);
or U22008 (N_22008,N_16953,N_18819);
and U22009 (N_22009,N_19284,N_19511);
nor U22010 (N_22010,N_15944,N_17434);
or U22011 (N_22011,N_19166,N_18776);
nor U22012 (N_22012,N_17490,N_16600);
nand U22013 (N_22013,N_19718,N_17905);
and U22014 (N_22014,N_19592,N_19054);
nor U22015 (N_22015,N_15202,N_18071);
nand U22016 (N_22016,N_16421,N_16217);
nand U22017 (N_22017,N_15677,N_17641);
nor U22018 (N_22018,N_19728,N_16327);
nor U22019 (N_22019,N_15060,N_19034);
nor U22020 (N_22020,N_16299,N_17253);
or U22021 (N_22021,N_18015,N_19408);
or U22022 (N_22022,N_19175,N_17230);
or U22023 (N_22023,N_19231,N_19276);
or U22024 (N_22024,N_18545,N_15569);
and U22025 (N_22025,N_15465,N_19482);
and U22026 (N_22026,N_19719,N_17620);
nor U22027 (N_22027,N_18946,N_17526);
and U22028 (N_22028,N_17308,N_17256);
nand U22029 (N_22029,N_16884,N_18671);
nor U22030 (N_22030,N_17766,N_19832);
nor U22031 (N_22031,N_17447,N_17359);
or U22032 (N_22032,N_19660,N_17857);
and U22033 (N_22033,N_18337,N_16172);
nand U22034 (N_22034,N_19260,N_19897);
nor U22035 (N_22035,N_17267,N_15308);
nor U22036 (N_22036,N_15536,N_19669);
nand U22037 (N_22037,N_19230,N_15729);
xnor U22038 (N_22038,N_15761,N_19936);
or U22039 (N_22039,N_19843,N_18304);
or U22040 (N_22040,N_18614,N_19955);
nor U22041 (N_22041,N_17076,N_19830);
nor U22042 (N_22042,N_17388,N_19795);
and U22043 (N_22043,N_18528,N_18091);
nor U22044 (N_22044,N_16179,N_16570);
and U22045 (N_22045,N_16462,N_16568);
nor U22046 (N_22046,N_19017,N_19102);
or U22047 (N_22047,N_15241,N_19536);
or U22048 (N_22048,N_16966,N_16123);
xnor U22049 (N_22049,N_19935,N_18233);
and U22050 (N_22050,N_16088,N_19570);
nand U22051 (N_22051,N_17168,N_17383);
and U22052 (N_22052,N_18262,N_19142);
or U22053 (N_22053,N_19605,N_18397);
and U22054 (N_22054,N_15643,N_15414);
xor U22055 (N_22055,N_16103,N_17070);
or U22056 (N_22056,N_18134,N_19115);
and U22057 (N_22057,N_16486,N_18653);
or U22058 (N_22058,N_18052,N_18923);
and U22059 (N_22059,N_18125,N_16868);
nor U22060 (N_22060,N_18005,N_16843);
nor U22061 (N_22061,N_15345,N_16122);
xnor U22062 (N_22062,N_17645,N_16857);
nor U22063 (N_22063,N_19130,N_15302);
xnor U22064 (N_22064,N_16248,N_19466);
nand U22065 (N_22065,N_18285,N_16205);
nand U22066 (N_22066,N_19468,N_16980);
and U22067 (N_22067,N_18258,N_15927);
and U22068 (N_22068,N_18251,N_15844);
nor U22069 (N_22069,N_17167,N_15298);
nand U22070 (N_22070,N_17671,N_19814);
and U22071 (N_22071,N_16756,N_19793);
and U22072 (N_22072,N_15280,N_19484);
nor U22073 (N_22073,N_18821,N_15706);
and U22074 (N_22074,N_17555,N_15734);
or U22075 (N_22075,N_15815,N_17376);
and U22076 (N_22076,N_19933,N_15748);
xor U22077 (N_22077,N_15181,N_17442);
xnor U22078 (N_22078,N_16682,N_17165);
nor U22079 (N_22079,N_18542,N_17338);
or U22080 (N_22080,N_17691,N_19682);
nand U22081 (N_22081,N_16703,N_19997);
and U22082 (N_22082,N_19820,N_16237);
nor U22083 (N_22083,N_18112,N_17853);
or U22084 (N_22084,N_17013,N_17716);
and U22085 (N_22085,N_18218,N_19168);
nand U22086 (N_22086,N_16202,N_15935);
nand U22087 (N_22087,N_17638,N_19485);
nand U22088 (N_22088,N_18805,N_17081);
nand U22089 (N_22089,N_16924,N_17843);
nor U22090 (N_22090,N_18960,N_17271);
and U22091 (N_22091,N_19310,N_17943);
and U22092 (N_22092,N_16793,N_17498);
and U22093 (N_22093,N_19804,N_16260);
or U22094 (N_22094,N_18524,N_17221);
nor U22095 (N_22095,N_18043,N_19344);
and U22096 (N_22096,N_17021,N_15213);
nand U22097 (N_22097,N_16640,N_18320);
and U22098 (N_22098,N_16529,N_15020);
nor U22099 (N_22099,N_16720,N_15757);
or U22100 (N_22100,N_17757,N_18461);
nand U22101 (N_22101,N_18915,N_18573);
and U22102 (N_22102,N_16484,N_16311);
xnor U22103 (N_22103,N_16187,N_16173);
xnor U22104 (N_22104,N_15390,N_17276);
nand U22105 (N_22105,N_18131,N_16012);
nand U22106 (N_22106,N_19077,N_19837);
and U22107 (N_22107,N_19581,N_18301);
and U22108 (N_22108,N_16115,N_15810);
nand U22109 (N_22109,N_17134,N_17939);
and U22110 (N_22110,N_16805,N_19713);
nand U22111 (N_22111,N_16598,N_19945);
and U22112 (N_22112,N_18885,N_19941);
nor U22113 (N_22113,N_19787,N_17637);
and U22114 (N_22114,N_15002,N_17612);
or U22115 (N_22115,N_19990,N_17129);
and U22116 (N_22116,N_18726,N_18693);
nor U22117 (N_22117,N_19453,N_17957);
xnor U22118 (N_22118,N_15366,N_19664);
and U22119 (N_22119,N_19478,N_15098);
xor U22120 (N_22120,N_15334,N_19966);
xor U22121 (N_22121,N_19577,N_16107);
nand U22122 (N_22122,N_15069,N_17906);
or U22123 (N_22123,N_17669,N_19934);
and U22124 (N_22124,N_19724,N_19220);
nor U22125 (N_22125,N_17871,N_17478);
xnor U22126 (N_22126,N_17166,N_15567);
nand U22127 (N_22127,N_16345,N_16666);
nor U22128 (N_22128,N_16998,N_19648);
nor U22129 (N_22129,N_17985,N_15876);
nand U22130 (N_22130,N_18239,N_18742);
xnor U22131 (N_22131,N_19683,N_19620);
nand U22132 (N_22132,N_17911,N_15573);
nor U22133 (N_22133,N_19707,N_16435);
and U22134 (N_22134,N_17416,N_18124);
and U22135 (N_22135,N_17030,N_15551);
or U22136 (N_22136,N_16135,N_16143);
and U22137 (N_22137,N_18826,N_18478);
nor U22138 (N_22138,N_17465,N_17126);
nor U22139 (N_22139,N_18236,N_16829);
nor U22140 (N_22140,N_19088,N_17474);
and U22141 (N_22141,N_18786,N_16501);
and U22142 (N_22142,N_17300,N_17882);
nor U22143 (N_22143,N_19326,N_15860);
or U22144 (N_22144,N_16097,N_18676);
nand U22145 (N_22145,N_18369,N_16454);
and U22146 (N_22146,N_15958,N_16513);
nor U22147 (N_22147,N_16925,N_17297);
nand U22148 (N_22148,N_17177,N_15332);
and U22149 (N_22149,N_18333,N_16978);
or U22150 (N_22150,N_15052,N_16046);
or U22151 (N_22151,N_17527,N_18934);
xor U22152 (N_22152,N_17894,N_18941);
or U22153 (N_22153,N_19510,N_18770);
and U22154 (N_22154,N_16918,N_17681);
or U22155 (N_22155,N_18480,N_19504);
or U22156 (N_22156,N_17932,N_19737);
nor U22157 (N_22157,N_17049,N_18010);
nor U22158 (N_22158,N_15575,N_18947);
xor U22159 (N_22159,N_19229,N_15005);
xor U22160 (N_22160,N_17472,N_15174);
or U22161 (N_22161,N_19900,N_17195);
and U22162 (N_22162,N_16326,N_15415);
and U22163 (N_22163,N_16803,N_17564);
or U22164 (N_22164,N_16687,N_15439);
and U22165 (N_22165,N_17961,N_19295);
and U22166 (N_22166,N_18642,N_18181);
or U22167 (N_22167,N_16368,N_19611);
nor U22168 (N_22168,N_17391,N_18807);
nand U22169 (N_22169,N_19337,N_17481);
nand U22170 (N_22170,N_19333,N_15170);
nor U22171 (N_22171,N_16833,N_19058);
xor U22172 (N_22172,N_18030,N_15263);
or U22173 (N_22173,N_15381,N_19835);
and U22174 (N_22174,N_16807,N_16892);
nand U22175 (N_22175,N_16983,N_16429);
or U22176 (N_22176,N_16199,N_17625);
and U22177 (N_22177,N_15425,N_18975);
nor U22178 (N_22178,N_15773,N_16284);
nor U22179 (N_22179,N_18291,N_18198);
nand U22180 (N_22180,N_16313,N_17254);
nor U22181 (N_22181,N_17583,N_16604);
xor U22182 (N_22182,N_16566,N_16333);
or U22183 (N_22183,N_19587,N_18169);
nor U22184 (N_22184,N_19821,N_15817);
nand U22185 (N_22185,N_18424,N_19414);
nand U22186 (N_22186,N_19630,N_15253);
nor U22187 (N_22187,N_16069,N_18710);
nor U22188 (N_22188,N_18531,N_19041);
nor U22189 (N_22189,N_16245,N_18681);
and U22190 (N_22190,N_15168,N_18828);
nand U22191 (N_22191,N_17861,N_18707);
or U22192 (N_22192,N_18142,N_19972);
nand U22193 (N_22193,N_16672,N_15990);
nand U22194 (N_22194,N_19459,N_18144);
or U22195 (N_22195,N_19312,N_15803);
nor U22196 (N_22196,N_16808,N_19503);
or U22197 (N_22197,N_17355,N_18607);
nor U22198 (N_22198,N_17453,N_18156);
xor U22199 (N_22199,N_18601,N_15552);
xnor U22200 (N_22200,N_19138,N_19100);
nor U22201 (N_22201,N_17738,N_15522);
nor U22202 (N_22202,N_15760,N_16949);
nand U22203 (N_22203,N_17649,N_19540);
nor U22204 (N_22204,N_16136,N_15854);
or U22205 (N_22205,N_17101,N_17802);
or U22206 (N_22206,N_17182,N_15733);
and U22207 (N_22207,N_17928,N_19506);
or U22208 (N_22208,N_19783,N_15539);
nand U22209 (N_22209,N_18012,N_18195);
nor U22210 (N_22210,N_16133,N_19527);
and U22211 (N_22211,N_19147,N_16783);
or U22212 (N_22212,N_15072,N_15553);
or U22213 (N_22213,N_15769,N_17673);
nand U22214 (N_22214,N_19606,N_17328);
or U22215 (N_22215,N_16347,N_16213);
xor U22216 (N_22216,N_17392,N_18973);
nand U22217 (N_22217,N_18550,N_17736);
nand U22218 (N_22218,N_19024,N_19823);
nand U22219 (N_22219,N_18797,N_17368);
nor U22220 (N_22220,N_15212,N_18683);
or U22221 (N_22221,N_16572,N_18365);
and U22222 (N_22222,N_16648,N_18768);
or U22223 (N_22223,N_18210,N_15206);
and U22224 (N_22224,N_17690,N_18317);
nand U22225 (N_22225,N_16470,N_19588);
nor U22226 (N_22226,N_17948,N_18873);
nand U22227 (N_22227,N_17414,N_16973);
nand U22228 (N_22228,N_17963,N_15451);
and U22229 (N_22229,N_19928,N_18256);
nand U22230 (N_22230,N_17989,N_16258);
nand U22231 (N_22231,N_15887,N_19454);
nand U22232 (N_22232,N_15637,N_17245);
nor U22233 (N_22233,N_15686,N_19422);
nor U22234 (N_22234,N_17535,N_17227);
nor U22235 (N_22235,N_19580,N_17387);
nand U22236 (N_22236,N_15599,N_18697);
xnor U22237 (N_22237,N_19411,N_17962);
nand U22238 (N_22238,N_18685,N_19025);
nand U22239 (N_22239,N_19926,N_15074);
and U22240 (N_22240,N_18687,N_15100);
nand U22241 (N_22241,N_15878,N_15687);
nand U22242 (N_22242,N_17425,N_18795);
or U22243 (N_22243,N_18402,N_19929);
nor U22244 (N_22244,N_15957,N_17529);
nor U22245 (N_22245,N_19675,N_17816);
nor U22246 (N_22246,N_16354,N_19401);
or U22247 (N_22247,N_19668,N_18600);
and U22248 (N_22248,N_18247,N_19144);
nor U22249 (N_22249,N_17044,N_16828);
nand U22250 (N_22250,N_19157,N_19901);
nor U22251 (N_22251,N_18939,N_18213);
and U22252 (N_22252,N_15432,N_19765);
nand U22253 (N_22253,N_17189,N_17683);
or U22254 (N_22254,N_16495,N_15956);
nand U22255 (N_22255,N_15141,N_17621);
and U22256 (N_22256,N_17283,N_16509);
nand U22257 (N_22257,N_19657,N_15793);
nand U22258 (N_22258,N_19039,N_16418);
or U22259 (N_22259,N_15008,N_15976);
and U22260 (N_22260,N_16083,N_15282);
nand U22261 (N_22261,N_19133,N_15688);
nor U22262 (N_22262,N_19223,N_16757);
nor U22263 (N_22263,N_17577,N_17900);
and U22264 (N_22264,N_17878,N_19712);
nor U22265 (N_22265,N_19911,N_16392);
and U22266 (N_22266,N_17967,N_17579);
nor U22267 (N_22267,N_19386,N_19907);
or U22268 (N_22268,N_17095,N_15129);
nor U22269 (N_22269,N_15438,N_15833);
nand U22270 (N_22270,N_17046,N_18082);
and U22271 (N_22271,N_16559,N_15847);
nand U22272 (N_22272,N_16852,N_17206);
nand U22273 (N_22273,N_17950,N_16463);
or U22274 (N_22274,N_18976,N_16576);
and U22275 (N_22275,N_19430,N_16655);
nor U22276 (N_22276,N_18452,N_18902);
or U22277 (N_22277,N_17666,N_18563);
or U22278 (N_22278,N_16407,N_16816);
nand U22279 (N_22279,N_19423,N_15946);
or U22280 (N_22280,N_17931,N_17821);
nand U22281 (N_22281,N_15825,N_16836);
or U22282 (N_22282,N_17596,N_18862);
nor U22283 (N_22283,N_18735,N_15911);
nor U22284 (N_22284,N_15616,N_16359);
and U22285 (N_22285,N_19774,N_18168);
and U22286 (N_22286,N_17902,N_19909);
nor U22287 (N_22287,N_18738,N_15426);
nand U22288 (N_22288,N_16515,N_15043);
nand U22289 (N_22289,N_17345,N_16923);
nor U22290 (N_22290,N_18718,N_17829);
xnor U22291 (N_22291,N_16692,N_19854);
nand U22292 (N_22292,N_17679,N_17984);
or U22293 (N_22293,N_15782,N_18638);
or U22294 (N_22294,N_19591,N_17019);
nand U22295 (N_22295,N_16350,N_19988);
or U22296 (N_22296,N_15226,N_18345);
and U22297 (N_22297,N_16739,N_16824);
and U22298 (N_22298,N_19806,N_17778);
xor U22299 (N_22299,N_15152,N_18729);
xor U22300 (N_22300,N_18093,N_17688);
and U22301 (N_22301,N_17503,N_17396);
or U22302 (N_22302,N_18381,N_16759);
nand U22303 (N_22303,N_17251,N_17032);
and U22304 (N_22304,N_18945,N_19525);
nor U22305 (N_22305,N_18115,N_19351);
and U22306 (N_22306,N_19850,N_17213);
or U22307 (N_22307,N_15635,N_19457);
or U22308 (N_22308,N_16935,N_16200);
xor U22309 (N_22309,N_16430,N_17965);
or U22310 (N_22310,N_17578,N_15645);
and U22311 (N_22311,N_15738,N_15148);
nor U22312 (N_22312,N_17605,N_15665);
or U22313 (N_22313,N_15796,N_16819);
nand U22314 (N_22314,N_19120,N_16901);
nand U22315 (N_22315,N_16346,N_16014);
nor U22316 (N_22316,N_18206,N_18040);
and U22317 (N_22317,N_15458,N_17313);
and U22318 (N_22318,N_16984,N_18456);
xor U22319 (N_22319,N_15116,N_16423);
and U22320 (N_22320,N_16539,N_19993);
and U22321 (N_22321,N_15704,N_18754);
nor U22322 (N_22322,N_17314,N_19319);
nor U22323 (N_22323,N_18944,N_15855);
nor U22324 (N_22324,N_17364,N_19541);
and U22325 (N_22325,N_19770,N_17817);
and U22326 (N_22326,N_18459,N_17685);
nand U22327 (N_22327,N_18922,N_17017);
and U22328 (N_22328,N_16149,N_17033);
or U22329 (N_22329,N_16673,N_19317);
and U22330 (N_22330,N_16453,N_16192);
and U22331 (N_22331,N_15187,N_16705);
nand U22332 (N_22332,N_19649,N_15448);
or U22333 (N_22333,N_16169,N_17369);
nand U22334 (N_22334,N_18987,N_18122);
and U22335 (N_22335,N_18179,N_15961);
or U22336 (N_22336,N_17850,N_17162);
xnor U22337 (N_22337,N_15906,N_19554);
xor U22338 (N_22338,N_16096,N_18086);
and U22339 (N_22339,N_16499,N_18850);
and U22340 (N_22340,N_18422,N_19434);
xor U22341 (N_22341,N_19069,N_16821);
and U22342 (N_22342,N_15481,N_16079);
and U22343 (N_22343,N_15650,N_18787);
or U22344 (N_22344,N_19329,N_16156);
or U22345 (N_22345,N_17734,N_16428);
xor U22346 (N_22346,N_19300,N_18628);
nor U22347 (N_22347,N_16571,N_17064);
nor U22348 (N_22348,N_17235,N_18265);
nand U22349 (N_22349,N_18264,N_15759);
nor U22350 (N_22350,N_16207,N_16651);
nand U22351 (N_22351,N_19890,N_16197);
or U22352 (N_22352,N_16422,N_15139);
and U22353 (N_22353,N_19785,N_19818);
and U22354 (N_22354,N_17826,N_16912);
or U22355 (N_22355,N_17924,N_15276);
or U22356 (N_22356,N_15433,N_17349);
and U22357 (N_22357,N_15699,N_16979);
and U22358 (N_22358,N_17846,N_17631);
or U22359 (N_22359,N_15491,N_15211);
nor U22360 (N_22360,N_15386,N_15344);
xor U22361 (N_22361,N_16058,N_18418);
nand U22362 (N_22362,N_19803,N_19372);
nor U22363 (N_22363,N_18833,N_19798);
nand U22364 (N_22364,N_15085,N_16785);
nand U22365 (N_22365,N_18003,N_18831);
or U22366 (N_22366,N_19726,N_19816);
nor U22367 (N_22367,N_15231,N_15740);
xnor U22368 (N_22368,N_18847,N_19045);
and U22369 (N_22369,N_18420,N_19258);
nand U22370 (N_22370,N_18836,N_19145);
nand U22371 (N_22371,N_15004,N_18467);
xnor U22372 (N_22372,N_19096,N_19604);
xnor U22373 (N_22373,N_18064,N_18498);
nand U22374 (N_22374,N_18037,N_19894);
nor U22375 (N_22375,N_17280,N_18603);
and U22376 (N_22376,N_17767,N_16400);
nor U22377 (N_22377,N_18289,N_17031);
or U22378 (N_22378,N_18592,N_16210);
xor U22379 (N_22379,N_15542,N_17604);
nor U22380 (N_22380,N_17974,N_19438);
nor U22381 (N_22381,N_18321,N_16461);
and U22382 (N_22382,N_15801,N_17559);
xor U22383 (N_22383,N_16522,N_16680);
and U22384 (N_22384,N_18659,N_16904);
nor U22385 (N_22385,N_18630,N_18867);
or U22386 (N_22386,N_15752,N_18539);
nor U22387 (N_22387,N_18510,N_15558);
or U22388 (N_22388,N_15984,N_15471);
and U22389 (N_22389,N_16639,N_16232);
nor U22390 (N_22390,N_19272,N_15937);
xor U22391 (N_22391,N_19943,N_19435);
nor U22392 (N_22392,N_15382,N_16837);
nand U22393 (N_22393,N_19780,N_19005);
or U22394 (N_22394,N_17090,N_15948);
and U22395 (N_22395,N_15925,N_18129);
nand U22396 (N_22396,N_19090,N_17994);
and U22397 (N_22397,N_18900,N_16693);
nand U22398 (N_22398,N_17565,N_19212);
or U22399 (N_22399,N_19244,N_17889);
nand U22400 (N_22400,N_17983,N_16804);
xor U22401 (N_22401,N_17651,N_17776);
and U22402 (N_22402,N_17891,N_17411);
nand U22403 (N_22403,N_16652,N_17544);
or U22404 (N_22404,N_16766,N_18791);
or U22405 (N_22405,N_17441,N_15016);
or U22406 (N_22406,N_15894,N_19266);
nor U22407 (N_22407,N_19800,N_18949);
xnor U22408 (N_22408,N_16940,N_19251);
nand U22409 (N_22409,N_15588,N_15791);
nor U22410 (N_22410,N_15423,N_15314);
or U22411 (N_22411,N_18549,N_16646);
nor U22412 (N_22412,N_19869,N_18095);
and U22413 (N_22413,N_18036,N_17112);
nor U22414 (N_22414,N_18746,N_17190);
or U22415 (N_22415,N_15589,N_19353);
or U22416 (N_22416,N_15172,N_19895);
or U22417 (N_22417,N_17409,N_18530);
and U22418 (N_22418,N_19753,N_17176);
nor U22419 (N_22419,N_15149,N_17854);
or U22420 (N_22420,N_15988,N_16063);
nor U22421 (N_22421,N_15417,N_19861);
nor U22422 (N_22422,N_19844,N_15392);
nand U22423 (N_22423,N_19544,N_18551);
and U22424 (N_22424,N_18327,N_18243);
nand U22425 (N_22425,N_19754,N_15765);
or U22426 (N_22426,N_18578,N_19983);
or U22427 (N_22427,N_17623,N_16577);
or U22428 (N_22428,N_19628,N_19944);
nor U22429 (N_22429,N_15541,N_19641);
nor U22430 (N_22430,N_15949,N_16157);
or U22431 (N_22431,N_19299,N_18722);
or U22432 (N_22432,N_15634,N_19870);
or U22433 (N_22433,N_16162,N_19250);
and U22434 (N_22434,N_16781,N_19044);
xor U22435 (N_22435,N_16203,N_15125);
nand U22436 (N_22436,N_15557,N_18307);
xnor U22437 (N_22437,N_15142,N_17457);
and U22438 (N_22438,N_16701,N_19357);
nand U22439 (N_22439,N_18719,N_18686);
or U22440 (N_22440,N_15718,N_15745);
nor U22441 (N_22441,N_18159,N_18961);
nand U22442 (N_22442,N_19491,N_15429);
nor U22443 (N_22443,N_17522,N_15410);
nor U22444 (N_22444,N_18084,N_17613);
and U22445 (N_22445,N_17755,N_19112);
or U22446 (N_22446,N_19826,N_17258);
and U22447 (N_22447,N_16614,N_17762);
and U22448 (N_22448,N_17799,N_16458);
nor U22449 (N_22449,N_18937,N_18556);
nand U22450 (N_22450,N_16560,N_19996);
nand U22451 (N_22451,N_18278,N_19093);
xnor U22452 (N_22452,N_17007,N_15033);
nor U22453 (N_22453,N_19172,N_16902);
and U22454 (N_22454,N_17403,N_15041);
or U22455 (N_22455,N_19343,N_19378);
or U22456 (N_22456,N_19651,N_15703);
and U22457 (N_22457,N_17607,N_17584);
xor U22458 (N_22458,N_17394,N_15256);
xor U22459 (N_22459,N_19589,N_19579);
xor U22460 (N_22460,N_18113,N_16787);
or U22461 (N_22461,N_18832,N_19007);
nor U22462 (N_22462,N_16633,N_18650);
nand U22463 (N_22463,N_16988,N_18958);
or U22464 (N_22464,N_18399,N_15905);
nor U22465 (N_22465,N_18018,N_15647);
and U22466 (N_22466,N_19207,N_19539);
nand U22467 (N_22467,N_19537,N_19467);
nand U22468 (N_22468,N_19962,N_17454);
or U22469 (N_22469,N_16286,N_15489);
and U22470 (N_22470,N_15749,N_17268);
nand U22471 (N_22471,N_15054,N_15078);
nand U22472 (N_22472,N_18745,N_15600);
or U22473 (N_22473,N_16320,N_19915);
or U22474 (N_22474,N_16711,N_17566);
xor U22475 (N_22475,N_17310,N_18039);
nand U22476 (N_22476,N_15678,N_19104);
or U22477 (N_22477,N_16015,N_17132);
nor U22478 (N_22478,N_17839,N_18133);
and U22479 (N_22479,N_19847,N_15257);
nand U22480 (N_22480,N_17241,N_18025);
and U22481 (N_22481,N_18070,N_17609);
and U22482 (N_22482,N_15251,N_18986);
and U22483 (N_22483,N_16003,N_17421);
and U22484 (N_22484,N_16076,N_15674);
and U22485 (N_22485,N_16880,N_15418);
and U22486 (N_22486,N_15412,N_19235);
nor U22487 (N_22487,N_16391,N_19868);
nand U22488 (N_22488,N_19989,N_17366);
and U22489 (N_22489,N_15189,N_18035);
nor U22490 (N_22490,N_17791,N_15238);
and U22491 (N_22491,N_15693,N_17563);
and U22492 (N_22492,N_17141,N_17043);
xnor U22493 (N_22493,N_17319,N_15466);
or U22494 (N_22494,N_15663,N_19610);
or U22495 (N_22495,N_18248,N_16516);
nor U22496 (N_22496,N_19970,N_19274);
or U22497 (N_22497,N_15128,N_19106);
nor U22498 (N_22498,N_16431,N_16835);
or U22499 (N_22499,N_19049,N_15300);
nor U22500 (N_22500,N_15894,N_15581);
or U22501 (N_22501,N_17395,N_17876);
nor U22502 (N_22502,N_18042,N_19687);
and U22503 (N_22503,N_18381,N_19575);
nand U22504 (N_22504,N_19234,N_19365);
xnor U22505 (N_22505,N_18110,N_19090);
xor U22506 (N_22506,N_18181,N_19790);
and U22507 (N_22507,N_19348,N_17115);
or U22508 (N_22508,N_18791,N_16205);
xor U22509 (N_22509,N_18154,N_19930);
xor U22510 (N_22510,N_15352,N_18276);
xor U22511 (N_22511,N_15252,N_15787);
or U22512 (N_22512,N_15691,N_19559);
or U22513 (N_22513,N_19416,N_15361);
or U22514 (N_22514,N_19483,N_15318);
xor U22515 (N_22515,N_18186,N_15115);
nor U22516 (N_22516,N_18004,N_17817);
and U22517 (N_22517,N_17783,N_19767);
and U22518 (N_22518,N_15717,N_18690);
nand U22519 (N_22519,N_19138,N_18997);
xnor U22520 (N_22520,N_16917,N_16434);
and U22521 (N_22521,N_15339,N_15181);
nor U22522 (N_22522,N_15041,N_16891);
nor U22523 (N_22523,N_16620,N_19916);
or U22524 (N_22524,N_15758,N_19753);
nand U22525 (N_22525,N_15012,N_16309);
and U22526 (N_22526,N_18862,N_18625);
nand U22527 (N_22527,N_19021,N_15667);
nand U22528 (N_22528,N_19347,N_16314);
and U22529 (N_22529,N_15994,N_15156);
nand U22530 (N_22530,N_15328,N_18161);
nand U22531 (N_22531,N_15251,N_16414);
nand U22532 (N_22532,N_16425,N_17392);
and U22533 (N_22533,N_18416,N_16118);
or U22534 (N_22534,N_19425,N_18159);
nand U22535 (N_22535,N_19134,N_17308);
or U22536 (N_22536,N_19963,N_16885);
nand U22537 (N_22537,N_19099,N_18562);
and U22538 (N_22538,N_19542,N_15849);
and U22539 (N_22539,N_17378,N_17604);
and U22540 (N_22540,N_16186,N_18391);
nand U22541 (N_22541,N_15379,N_17361);
nand U22542 (N_22542,N_15052,N_19898);
nand U22543 (N_22543,N_19434,N_17772);
and U22544 (N_22544,N_17399,N_18198);
nand U22545 (N_22545,N_17876,N_17933);
or U22546 (N_22546,N_19454,N_15082);
and U22547 (N_22547,N_19652,N_15793);
nor U22548 (N_22548,N_17570,N_19180);
nand U22549 (N_22549,N_19372,N_16793);
and U22550 (N_22550,N_15202,N_17689);
or U22551 (N_22551,N_15908,N_16477);
or U22552 (N_22552,N_17793,N_19262);
nor U22553 (N_22553,N_17569,N_16196);
xor U22554 (N_22554,N_15813,N_18844);
or U22555 (N_22555,N_15703,N_19300);
nand U22556 (N_22556,N_18578,N_17304);
or U22557 (N_22557,N_15812,N_19018);
and U22558 (N_22558,N_16184,N_18336);
nand U22559 (N_22559,N_17147,N_16284);
nor U22560 (N_22560,N_17545,N_19614);
and U22561 (N_22561,N_17679,N_18395);
and U22562 (N_22562,N_18664,N_17492);
or U22563 (N_22563,N_18736,N_17155);
and U22564 (N_22564,N_16934,N_16738);
and U22565 (N_22565,N_19626,N_16036);
nor U22566 (N_22566,N_17944,N_18941);
or U22567 (N_22567,N_16602,N_16543);
xor U22568 (N_22568,N_18980,N_19679);
nor U22569 (N_22569,N_18914,N_16967);
or U22570 (N_22570,N_15591,N_15736);
xnor U22571 (N_22571,N_15137,N_17400);
nor U22572 (N_22572,N_16205,N_19290);
and U22573 (N_22573,N_16380,N_19285);
xor U22574 (N_22574,N_19950,N_16793);
nor U22575 (N_22575,N_17062,N_17338);
nor U22576 (N_22576,N_18732,N_16949);
and U22577 (N_22577,N_17268,N_18914);
or U22578 (N_22578,N_19675,N_15205);
or U22579 (N_22579,N_15329,N_19305);
and U22580 (N_22580,N_18533,N_18831);
nand U22581 (N_22581,N_18331,N_15695);
xor U22582 (N_22582,N_19791,N_16001);
nand U22583 (N_22583,N_17345,N_16057);
nor U22584 (N_22584,N_15160,N_15518);
nand U22585 (N_22585,N_19661,N_19585);
nor U22586 (N_22586,N_18111,N_16715);
and U22587 (N_22587,N_18709,N_17142);
xnor U22588 (N_22588,N_16213,N_15968);
nand U22589 (N_22589,N_15886,N_18053);
nor U22590 (N_22590,N_17295,N_19638);
and U22591 (N_22591,N_17745,N_15670);
or U22592 (N_22592,N_17357,N_18673);
xor U22593 (N_22593,N_16799,N_15188);
nand U22594 (N_22594,N_19247,N_16422);
nor U22595 (N_22595,N_17679,N_18071);
and U22596 (N_22596,N_15665,N_19483);
and U22597 (N_22597,N_19565,N_15331);
nor U22598 (N_22598,N_15301,N_15772);
or U22599 (N_22599,N_16776,N_17239);
and U22600 (N_22600,N_19946,N_19797);
nor U22601 (N_22601,N_16154,N_19588);
nor U22602 (N_22602,N_18090,N_18303);
nand U22603 (N_22603,N_15349,N_19948);
nor U22604 (N_22604,N_17396,N_16986);
and U22605 (N_22605,N_16368,N_18593);
nand U22606 (N_22606,N_17526,N_15160);
nand U22607 (N_22607,N_15622,N_19913);
and U22608 (N_22608,N_15293,N_17440);
or U22609 (N_22609,N_18912,N_16069);
or U22610 (N_22610,N_19212,N_19032);
and U22611 (N_22611,N_19141,N_17639);
xnor U22612 (N_22612,N_17802,N_16533);
nand U22613 (N_22613,N_19886,N_18220);
and U22614 (N_22614,N_18091,N_19861);
nor U22615 (N_22615,N_17530,N_15980);
nand U22616 (N_22616,N_17258,N_16783);
and U22617 (N_22617,N_18385,N_18384);
or U22618 (N_22618,N_19159,N_15976);
nand U22619 (N_22619,N_15731,N_15219);
nor U22620 (N_22620,N_16887,N_16112);
xor U22621 (N_22621,N_15247,N_15308);
nor U22622 (N_22622,N_15741,N_16913);
nand U22623 (N_22623,N_18449,N_17648);
or U22624 (N_22624,N_19581,N_18572);
xnor U22625 (N_22625,N_18167,N_18675);
xnor U22626 (N_22626,N_18712,N_18515);
nor U22627 (N_22627,N_18878,N_17539);
nand U22628 (N_22628,N_17846,N_16273);
nand U22629 (N_22629,N_18596,N_19066);
or U22630 (N_22630,N_19221,N_16248);
and U22631 (N_22631,N_15836,N_15145);
and U22632 (N_22632,N_17565,N_16711);
nor U22633 (N_22633,N_16677,N_17860);
or U22634 (N_22634,N_18089,N_16185);
and U22635 (N_22635,N_15546,N_15203);
nand U22636 (N_22636,N_17862,N_17547);
or U22637 (N_22637,N_18855,N_19714);
nand U22638 (N_22638,N_18848,N_17667);
nand U22639 (N_22639,N_19304,N_17581);
nand U22640 (N_22640,N_16059,N_17431);
nor U22641 (N_22641,N_15503,N_15804);
nand U22642 (N_22642,N_16989,N_15755);
nor U22643 (N_22643,N_17527,N_18412);
and U22644 (N_22644,N_17640,N_19841);
and U22645 (N_22645,N_15549,N_17577);
nor U22646 (N_22646,N_16368,N_17770);
nor U22647 (N_22647,N_17631,N_16277);
nor U22648 (N_22648,N_19076,N_19619);
and U22649 (N_22649,N_17003,N_17936);
or U22650 (N_22650,N_19141,N_17553);
xnor U22651 (N_22651,N_19815,N_18799);
nand U22652 (N_22652,N_18273,N_19118);
or U22653 (N_22653,N_19231,N_19030);
nand U22654 (N_22654,N_15641,N_19152);
nand U22655 (N_22655,N_17799,N_15001);
and U22656 (N_22656,N_16224,N_15823);
xnor U22657 (N_22657,N_17043,N_19992);
nor U22658 (N_22658,N_17373,N_15317);
and U22659 (N_22659,N_19850,N_16974);
nand U22660 (N_22660,N_15860,N_18870);
nor U22661 (N_22661,N_17284,N_18946);
and U22662 (N_22662,N_19105,N_17091);
or U22663 (N_22663,N_15478,N_17911);
nand U22664 (N_22664,N_18206,N_16956);
nor U22665 (N_22665,N_16942,N_17799);
nor U22666 (N_22666,N_17589,N_15280);
or U22667 (N_22667,N_16167,N_16730);
and U22668 (N_22668,N_18192,N_16856);
and U22669 (N_22669,N_15391,N_15204);
nor U22670 (N_22670,N_16908,N_17549);
nand U22671 (N_22671,N_18371,N_17709);
nor U22672 (N_22672,N_17897,N_18218);
nor U22673 (N_22673,N_17675,N_15558);
or U22674 (N_22674,N_19884,N_18404);
nor U22675 (N_22675,N_19677,N_17825);
and U22676 (N_22676,N_18815,N_18679);
or U22677 (N_22677,N_17977,N_17488);
and U22678 (N_22678,N_17269,N_15781);
or U22679 (N_22679,N_15118,N_17356);
nor U22680 (N_22680,N_17007,N_17943);
xnor U22681 (N_22681,N_18663,N_15412);
nand U22682 (N_22682,N_16628,N_19240);
or U22683 (N_22683,N_16493,N_18606);
and U22684 (N_22684,N_18367,N_18893);
nor U22685 (N_22685,N_17044,N_16089);
nor U22686 (N_22686,N_15226,N_16016);
nand U22687 (N_22687,N_18779,N_19785);
nor U22688 (N_22688,N_16205,N_17512);
nand U22689 (N_22689,N_17440,N_17942);
and U22690 (N_22690,N_16814,N_17920);
nor U22691 (N_22691,N_18122,N_18595);
nor U22692 (N_22692,N_15421,N_16143);
and U22693 (N_22693,N_15560,N_16176);
nand U22694 (N_22694,N_15128,N_16217);
nand U22695 (N_22695,N_19795,N_15508);
nor U22696 (N_22696,N_18146,N_18114);
nand U22697 (N_22697,N_18962,N_17214);
or U22698 (N_22698,N_16649,N_17445);
and U22699 (N_22699,N_18523,N_16000);
nor U22700 (N_22700,N_16390,N_17500);
nand U22701 (N_22701,N_17924,N_17218);
nor U22702 (N_22702,N_18560,N_19386);
nor U22703 (N_22703,N_19094,N_18433);
nand U22704 (N_22704,N_18090,N_16055);
nor U22705 (N_22705,N_16720,N_19864);
xnor U22706 (N_22706,N_16817,N_18362);
xnor U22707 (N_22707,N_17743,N_15701);
nand U22708 (N_22708,N_18206,N_18052);
nand U22709 (N_22709,N_15020,N_18728);
xnor U22710 (N_22710,N_16435,N_16408);
and U22711 (N_22711,N_18935,N_17157);
nand U22712 (N_22712,N_17003,N_19390);
or U22713 (N_22713,N_17235,N_15342);
nand U22714 (N_22714,N_18255,N_19654);
and U22715 (N_22715,N_16276,N_17336);
nor U22716 (N_22716,N_17483,N_18246);
and U22717 (N_22717,N_15859,N_15219);
nor U22718 (N_22718,N_18351,N_17499);
nor U22719 (N_22719,N_17333,N_17014);
and U22720 (N_22720,N_15500,N_19041);
or U22721 (N_22721,N_15624,N_19581);
xor U22722 (N_22722,N_16175,N_18931);
nand U22723 (N_22723,N_18423,N_15075);
nor U22724 (N_22724,N_17795,N_18857);
nand U22725 (N_22725,N_19728,N_18750);
or U22726 (N_22726,N_17163,N_16315);
xor U22727 (N_22727,N_15580,N_16035);
and U22728 (N_22728,N_17683,N_17195);
nand U22729 (N_22729,N_16923,N_16345);
nor U22730 (N_22730,N_15688,N_16249);
nor U22731 (N_22731,N_18425,N_18031);
nor U22732 (N_22732,N_15395,N_17893);
nor U22733 (N_22733,N_19527,N_19017);
nand U22734 (N_22734,N_19625,N_16003);
or U22735 (N_22735,N_19482,N_16013);
nand U22736 (N_22736,N_18593,N_19800);
or U22737 (N_22737,N_19760,N_17490);
nand U22738 (N_22738,N_19231,N_18172);
nor U22739 (N_22739,N_16884,N_17606);
and U22740 (N_22740,N_15372,N_15163);
or U22741 (N_22741,N_15400,N_18299);
or U22742 (N_22742,N_19534,N_15663);
and U22743 (N_22743,N_15037,N_17357);
or U22744 (N_22744,N_18039,N_15587);
or U22745 (N_22745,N_17967,N_15720);
nand U22746 (N_22746,N_18811,N_16957);
and U22747 (N_22747,N_17591,N_16692);
or U22748 (N_22748,N_16702,N_18600);
or U22749 (N_22749,N_16585,N_17101);
nand U22750 (N_22750,N_19382,N_19490);
nor U22751 (N_22751,N_17516,N_18037);
and U22752 (N_22752,N_16681,N_17484);
and U22753 (N_22753,N_15040,N_17870);
nor U22754 (N_22754,N_16863,N_17467);
or U22755 (N_22755,N_17079,N_15995);
nor U22756 (N_22756,N_19225,N_16790);
nor U22757 (N_22757,N_19137,N_16260);
or U22758 (N_22758,N_16991,N_18231);
or U22759 (N_22759,N_16975,N_17835);
nor U22760 (N_22760,N_19568,N_15471);
nor U22761 (N_22761,N_17573,N_15829);
and U22762 (N_22762,N_19679,N_18547);
nor U22763 (N_22763,N_16776,N_15910);
nor U22764 (N_22764,N_16703,N_19602);
nor U22765 (N_22765,N_17404,N_19162);
and U22766 (N_22766,N_19237,N_19719);
xnor U22767 (N_22767,N_18784,N_17763);
nand U22768 (N_22768,N_17919,N_18236);
nor U22769 (N_22769,N_15619,N_19921);
or U22770 (N_22770,N_19864,N_18752);
nand U22771 (N_22771,N_19185,N_18043);
or U22772 (N_22772,N_18605,N_15881);
xor U22773 (N_22773,N_16083,N_17955);
or U22774 (N_22774,N_19987,N_16031);
nand U22775 (N_22775,N_16510,N_15564);
nor U22776 (N_22776,N_16827,N_18205);
nor U22777 (N_22777,N_18474,N_15748);
nand U22778 (N_22778,N_17780,N_15175);
nand U22779 (N_22779,N_18641,N_19865);
and U22780 (N_22780,N_18350,N_16995);
and U22781 (N_22781,N_17338,N_17158);
nand U22782 (N_22782,N_18102,N_19195);
nor U22783 (N_22783,N_15323,N_18122);
and U22784 (N_22784,N_16555,N_18229);
and U22785 (N_22785,N_15202,N_19540);
nor U22786 (N_22786,N_17330,N_17554);
xnor U22787 (N_22787,N_18749,N_18838);
nor U22788 (N_22788,N_19384,N_19302);
nor U22789 (N_22789,N_15755,N_16938);
or U22790 (N_22790,N_19112,N_18927);
and U22791 (N_22791,N_15328,N_18262);
or U22792 (N_22792,N_15422,N_17487);
and U22793 (N_22793,N_19177,N_17217);
or U22794 (N_22794,N_16922,N_18187);
and U22795 (N_22795,N_17935,N_15336);
or U22796 (N_22796,N_17532,N_19954);
or U22797 (N_22797,N_18321,N_16219);
and U22798 (N_22798,N_16878,N_18896);
nand U22799 (N_22799,N_19268,N_19129);
nand U22800 (N_22800,N_19361,N_19445);
and U22801 (N_22801,N_16386,N_16456);
or U22802 (N_22802,N_19912,N_16946);
nor U22803 (N_22803,N_16917,N_17785);
nor U22804 (N_22804,N_19118,N_19331);
or U22805 (N_22805,N_17210,N_16788);
and U22806 (N_22806,N_15931,N_19271);
nor U22807 (N_22807,N_18275,N_18578);
and U22808 (N_22808,N_15371,N_19128);
or U22809 (N_22809,N_15841,N_15988);
nor U22810 (N_22810,N_16381,N_19494);
xor U22811 (N_22811,N_16622,N_17128);
nor U22812 (N_22812,N_19313,N_15852);
or U22813 (N_22813,N_16666,N_18498);
nand U22814 (N_22814,N_15402,N_19692);
and U22815 (N_22815,N_16384,N_17778);
or U22816 (N_22816,N_15469,N_17608);
or U22817 (N_22817,N_16327,N_18096);
or U22818 (N_22818,N_16113,N_16075);
xor U22819 (N_22819,N_15732,N_16430);
nor U22820 (N_22820,N_16072,N_17286);
or U22821 (N_22821,N_16773,N_19372);
xor U22822 (N_22822,N_15120,N_15517);
nor U22823 (N_22823,N_19072,N_16266);
xnor U22824 (N_22824,N_19463,N_15981);
nor U22825 (N_22825,N_17067,N_15089);
or U22826 (N_22826,N_17691,N_17421);
or U22827 (N_22827,N_15415,N_19683);
nand U22828 (N_22828,N_15216,N_17194);
nor U22829 (N_22829,N_18855,N_18460);
and U22830 (N_22830,N_19429,N_18319);
nand U22831 (N_22831,N_16762,N_18718);
and U22832 (N_22832,N_18327,N_18754);
or U22833 (N_22833,N_19769,N_16199);
nand U22834 (N_22834,N_19460,N_16961);
nand U22835 (N_22835,N_16152,N_16434);
xnor U22836 (N_22836,N_15898,N_17303);
nand U22837 (N_22837,N_18281,N_16974);
or U22838 (N_22838,N_19758,N_18026);
or U22839 (N_22839,N_18359,N_16945);
nor U22840 (N_22840,N_19418,N_15668);
nand U22841 (N_22841,N_15783,N_17946);
or U22842 (N_22842,N_15296,N_15458);
or U22843 (N_22843,N_16972,N_18462);
xor U22844 (N_22844,N_18451,N_15644);
xnor U22845 (N_22845,N_19755,N_18218);
or U22846 (N_22846,N_18307,N_16548);
or U22847 (N_22847,N_17516,N_17948);
or U22848 (N_22848,N_19962,N_15066);
or U22849 (N_22849,N_17537,N_15480);
nand U22850 (N_22850,N_18406,N_16232);
or U22851 (N_22851,N_16554,N_17221);
or U22852 (N_22852,N_17597,N_16588);
and U22853 (N_22853,N_16212,N_16681);
and U22854 (N_22854,N_19909,N_18788);
nor U22855 (N_22855,N_19848,N_19798);
and U22856 (N_22856,N_18012,N_15235);
and U22857 (N_22857,N_17320,N_16812);
xnor U22858 (N_22858,N_16305,N_18078);
nor U22859 (N_22859,N_15896,N_18267);
nand U22860 (N_22860,N_19561,N_15113);
xnor U22861 (N_22861,N_19739,N_16551);
nor U22862 (N_22862,N_15154,N_17375);
nor U22863 (N_22863,N_15415,N_17843);
or U22864 (N_22864,N_16621,N_17550);
and U22865 (N_22865,N_16628,N_19301);
nand U22866 (N_22866,N_19151,N_15422);
nand U22867 (N_22867,N_15499,N_16929);
nand U22868 (N_22868,N_18004,N_19241);
or U22869 (N_22869,N_16583,N_16861);
or U22870 (N_22870,N_15415,N_18910);
or U22871 (N_22871,N_17527,N_19801);
nand U22872 (N_22872,N_15503,N_19950);
and U22873 (N_22873,N_16354,N_16279);
nand U22874 (N_22874,N_19514,N_15636);
nand U22875 (N_22875,N_17036,N_19248);
or U22876 (N_22876,N_15325,N_17803);
xor U22877 (N_22877,N_17978,N_18697);
nor U22878 (N_22878,N_18549,N_17139);
xnor U22879 (N_22879,N_16604,N_15487);
and U22880 (N_22880,N_16887,N_15955);
nand U22881 (N_22881,N_19764,N_16882);
nand U22882 (N_22882,N_16723,N_15088);
and U22883 (N_22883,N_15443,N_19573);
or U22884 (N_22884,N_17441,N_17079);
nor U22885 (N_22885,N_18046,N_18549);
and U22886 (N_22886,N_19947,N_15384);
nor U22887 (N_22887,N_15576,N_18026);
or U22888 (N_22888,N_18115,N_19554);
nand U22889 (N_22889,N_15533,N_16903);
nand U22890 (N_22890,N_18086,N_17749);
nor U22891 (N_22891,N_16882,N_16354);
nand U22892 (N_22892,N_15386,N_19232);
and U22893 (N_22893,N_16448,N_17578);
nor U22894 (N_22894,N_18113,N_19426);
or U22895 (N_22895,N_15531,N_18046);
nand U22896 (N_22896,N_17444,N_19611);
or U22897 (N_22897,N_17082,N_18291);
or U22898 (N_22898,N_17672,N_18202);
nor U22899 (N_22899,N_15392,N_16100);
nor U22900 (N_22900,N_15932,N_17085);
nand U22901 (N_22901,N_19249,N_15270);
and U22902 (N_22902,N_15553,N_19101);
and U22903 (N_22903,N_19134,N_17191);
nor U22904 (N_22904,N_17521,N_19915);
or U22905 (N_22905,N_17792,N_16542);
nor U22906 (N_22906,N_15923,N_17580);
nor U22907 (N_22907,N_17940,N_18106);
nand U22908 (N_22908,N_17382,N_19560);
and U22909 (N_22909,N_19796,N_17017);
and U22910 (N_22910,N_19183,N_15031);
or U22911 (N_22911,N_18203,N_18486);
nand U22912 (N_22912,N_16190,N_18340);
nor U22913 (N_22913,N_16696,N_19755);
or U22914 (N_22914,N_16620,N_17269);
or U22915 (N_22915,N_19790,N_15789);
nor U22916 (N_22916,N_17772,N_17475);
and U22917 (N_22917,N_16145,N_16002);
xnor U22918 (N_22918,N_19639,N_16887);
xnor U22919 (N_22919,N_16905,N_17101);
or U22920 (N_22920,N_16417,N_15033);
and U22921 (N_22921,N_17928,N_19965);
or U22922 (N_22922,N_18054,N_16766);
nor U22923 (N_22923,N_16433,N_18482);
or U22924 (N_22924,N_17439,N_17773);
nand U22925 (N_22925,N_17766,N_15619);
or U22926 (N_22926,N_19793,N_18084);
nand U22927 (N_22927,N_17372,N_18110);
nand U22928 (N_22928,N_17426,N_16753);
nor U22929 (N_22929,N_17546,N_16962);
nor U22930 (N_22930,N_17397,N_18277);
and U22931 (N_22931,N_18061,N_15696);
xor U22932 (N_22932,N_16238,N_17528);
or U22933 (N_22933,N_16607,N_18953);
or U22934 (N_22934,N_17575,N_16931);
or U22935 (N_22935,N_18538,N_15589);
or U22936 (N_22936,N_19626,N_19905);
nor U22937 (N_22937,N_16847,N_18759);
and U22938 (N_22938,N_15421,N_18719);
nand U22939 (N_22939,N_15333,N_15560);
nor U22940 (N_22940,N_16439,N_18327);
nand U22941 (N_22941,N_18350,N_19450);
nand U22942 (N_22942,N_15282,N_15331);
nor U22943 (N_22943,N_18724,N_15455);
and U22944 (N_22944,N_16002,N_17907);
or U22945 (N_22945,N_15033,N_18437);
nand U22946 (N_22946,N_19128,N_16653);
xnor U22947 (N_22947,N_17114,N_18481);
xnor U22948 (N_22948,N_19455,N_19658);
xor U22949 (N_22949,N_15576,N_17680);
nand U22950 (N_22950,N_19976,N_19588);
and U22951 (N_22951,N_17185,N_17965);
and U22952 (N_22952,N_19192,N_15210);
nor U22953 (N_22953,N_15684,N_17329);
nor U22954 (N_22954,N_16944,N_19187);
and U22955 (N_22955,N_16451,N_18805);
xnor U22956 (N_22956,N_17096,N_19133);
nand U22957 (N_22957,N_18552,N_17768);
and U22958 (N_22958,N_18472,N_16922);
and U22959 (N_22959,N_15962,N_19123);
and U22960 (N_22960,N_16755,N_15297);
xor U22961 (N_22961,N_15656,N_16232);
or U22962 (N_22962,N_19029,N_17856);
nand U22963 (N_22963,N_15998,N_19192);
and U22964 (N_22964,N_17224,N_18228);
or U22965 (N_22965,N_15245,N_17397);
nor U22966 (N_22966,N_17197,N_18107);
nor U22967 (N_22967,N_17059,N_17323);
and U22968 (N_22968,N_19298,N_18656);
or U22969 (N_22969,N_15505,N_15486);
nor U22970 (N_22970,N_16498,N_19914);
nand U22971 (N_22971,N_19039,N_19886);
nand U22972 (N_22972,N_17147,N_16643);
nor U22973 (N_22973,N_16672,N_18819);
or U22974 (N_22974,N_15913,N_16412);
or U22975 (N_22975,N_16341,N_15763);
or U22976 (N_22976,N_19692,N_15600);
nand U22977 (N_22977,N_19959,N_15757);
nand U22978 (N_22978,N_16881,N_15491);
or U22979 (N_22979,N_16263,N_18241);
or U22980 (N_22980,N_17430,N_15997);
nand U22981 (N_22981,N_18752,N_19387);
and U22982 (N_22982,N_18190,N_19158);
or U22983 (N_22983,N_15928,N_18732);
or U22984 (N_22984,N_16585,N_18029);
nor U22985 (N_22985,N_17950,N_19791);
xnor U22986 (N_22986,N_17163,N_18685);
nand U22987 (N_22987,N_19225,N_18542);
nor U22988 (N_22988,N_18634,N_17800);
or U22989 (N_22989,N_18803,N_17284);
nor U22990 (N_22990,N_19857,N_17132);
nand U22991 (N_22991,N_15059,N_15105);
xor U22992 (N_22992,N_17841,N_19006);
or U22993 (N_22993,N_17945,N_15282);
or U22994 (N_22994,N_15218,N_17777);
nor U22995 (N_22995,N_18295,N_17845);
and U22996 (N_22996,N_15307,N_19215);
nor U22997 (N_22997,N_17242,N_18519);
nor U22998 (N_22998,N_15477,N_17575);
nand U22999 (N_22999,N_15048,N_16450);
nand U23000 (N_23000,N_15088,N_17801);
and U23001 (N_23001,N_19753,N_16748);
or U23002 (N_23002,N_18898,N_19455);
or U23003 (N_23003,N_15560,N_17651);
or U23004 (N_23004,N_19962,N_19310);
and U23005 (N_23005,N_16648,N_17499);
and U23006 (N_23006,N_18451,N_18775);
nor U23007 (N_23007,N_15999,N_19729);
xnor U23008 (N_23008,N_17045,N_17334);
nand U23009 (N_23009,N_15552,N_17259);
and U23010 (N_23010,N_16300,N_16269);
nor U23011 (N_23011,N_15483,N_17475);
nand U23012 (N_23012,N_17928,N_15047);
and U23013 (N_23013,N_18333,N_15551);
nand U23014 (N_23014,N_15628,N_17003);
nor U23015 (N_23015,N_18940,N_17677);
and U23016 (N_23016,N_16473,N_16658);
and U23017 (N_23017,N_17070,N_15498);
nand U23018 (N_23018,N_18523,N_18717);
and U23019 (N_23019,N_16838,N_18041);
or U23020 (N_23020,N_16247,N_17583);
and U23021 (N_23021,N_19308,N_17369);
and U23022 (N_23022,N_16695,N_18996);
or U23023 (N_23023,N_15109,N_19603);
or U23024 (N_23024,N_19897,N_16843);
and U23025 (N_23025,N_15464,N_17373);
or U23026 (N_23026,N_18870,N_15188);
or U23027 (N_23027,N_18951,N_15093);
nor U23028 (N_23028,N_15323,N_17890);
or U23029 (N_23029,N_18149,N_15051);
and U23030 (N_23030,N_16320,N_17450);
and U23031 (N_23031,N_17542,N_17250);
nand U23032 (N_23032,N_18812,N_19010);
and U23033 (N_23033,N_15743,N_16645);
xor U23034 (N_23034,N_18604,N_15978);
xnor U23035 (N_23035,N_18191,N_18313);
or U23036 (N_23036,N_18332,N_16692);
and U23037 (N_23037,N_16598,N_16554);
nor U23038 (N_23038,N_17111,N_16182);
nand U23039 (N_23039,N_15084,N_18692);
or U23040 (N_23040,N_19527,N_18874);
or U23041 (N_23041,N_18081,N_18638);
nor U23042 (N_23042,N_16246,N_17855);
nand U23043 (N_23043,N_16226,N_15621);
and U23044 (N_23044,N_19138,N_16890);
nor U23045 (N_23045,N_16358,N_15017);
and U23046 (N_23046,N_17519,N_16705);
nand U23047 (N_23047,N_15932,N_18708);
and U23048 (N_23048,N_17948,N_18898);
nand U23049 (N_23049,N_18772,N_15760);
or U23050 (N_23050,N_18700,N_17026);
nor U23051 (N_23051,N_18631,N_16657);
xnor U23052 (N_23052,N_18547,N_17173);
nor U23053 (N_23053,N_15007,N_15358);
nor U23054 (N_23054,N_18193,N_15018);
and U23055 (N_23055,N_19262,N_18702);
nand U23056 (N_23056,N_19000,N_15863);
or U23057 (N_23057,N_18955,N_19870);
or U23058 (N_23058,N_16465,N_17705);
nor U23059 (N_23059,N_15209,N_16026);
or U23060 (N_23060,N_16039,N_16802);
or U23061 (N_23061,N_17862,N_19268);
or U23062 (N_23062,N_17027,N_16017);
or U23063 (N_23063,N_18787,N_15092);
and U23064 (N_23064,N_16154,N_19462);
or U23065 (N_23065,N_17371,N_17908);
xor U23066 (N_23066,N_18744,N_15671);
nor U23067 (N_23067,N_18040,N_18993);
nor U23068 (N_23068,N_19205,N_19063);
and U23069 (N_23069,N_15734,N_18001);
or U23070 (N_23070,N_19710,N_18010);
or U23071 (N_23071,N_16369,N_17284);
nor U23072 (N_23072,N_18248,N_16783);
nand U23073 (N_23073,N_18835,N_16792);
nor U23074 (N_23074,N_17855,N_18517);
xor U23075 (N_23075,N_17266,N_17770);
nand U23076 (N_23076,N_16532,N_19461);
nand U23077 (N_23077,N_18505,N_16156);
or U23078 (N_23078,N_17065,N_18562);
or U23079 (N_23079,N_15831,N_18464);
or U23080 (N_23080,N_18234,N_16196);
nor U23081 (N_23081,N_18775,N_17732);
nand U23082 (N_23082,N_19300,N_17153);
and U23083 (N_23083,N_16378,N_19300);
or U23084 (N_23084,N_15852,N_15549);
and U23085 (N_23085,N_19829,N_15698);
nor U23086 (N_23086,N_17592,N_16880);
nand U23087 (N_23087,N_16628,N_16588);
and U23088 (N_23088,N_15883,N_19248);
nand U23089 (N_23089,N_17241,N_16117);
and U23090 (N_23090,N_15756,N_15957);
nor U23091 (N_23091,N_18756,N_19301);
or U23092 (N_23092,N_15838,N_15198);
or U23093 (N_23093,N_16114,N_15834);
xnor U23094 (N_23094,N_19493,N_17569);
xor U23095 (N_23095,N_17908,N_19858);
xor U23096 (N_23096,N_19752,N_16053);
xnor U23097 (N_23097,N_15656,N_15364);
and U23098 (N_23098,N_18690,N_18979);
nor U23099 (N_23099,N_16786,N_19687);
or U23100 (N_23100,N_16739,N_19353);
and U23101 (N_23101,N_19317,N_19261);
nor U23102 (N_23102,N_18924,N_15200);
or U23103 (N_23103,N_18167,N_19214);
and U23104 (N_23104,N_17806,N_17155);
nand U23105 (N_23105,N_16310,N_16154);
nor U23106 (N_23106,N_15489,N_18295);
nor U23107 (N_23107,N_17384,N_17804);
nor U23108 (N_23108,N_16145,N_15276);
or U23109 (N_23109,N_18543,N_17643);
xor U23110 (N_23110,N_17721,N_17491);
nor U23111 (N_23111,N_16933,N_16221);
or U23112 (N_23112,N_16094,N_19812);
nor U23113 (N_23113,N_16726,N_15523);
or U23114 (N_23114,N_19491,N_17614);
nor U23115 (N_23115,N_16409,N_15714);
or U23116 (N_23116,N_18488,N_16957);
nand U23117 (N_23117,N_18008,N_18086);
and U23118 (N_23118,N_17767,N_17353);
and U23119 (N_23119,N_15700,N_16133);
nand U23120 (N_23120,N_17576,N_18359);
nand U23121 (N_23121,N_19452,N_19991);
nand U23122 (N_23122,N_15375,N_19951);
nor U23123 (N_23123,N_16023,N_19427);
or U23124 (N_23124,N_16310,N_17357);
or U23125 (N_23125,N_15593,N_17498);
and U23126 (N_23126,N_17474,N_19026);
nor U23127 (N_23127,N_19793,N_18410);
and U23128 (N_23128,N_17915,N_19012);
nor U23129 (N_23129,N_19020,N_15450);
or U23130 (N_23130,N_15935,N_17233);
or U23131 (N_23131,N_15237,N_16666);
nand U23132 (N_23132,N_16861,N_18948);
nor U23133 (N_23133,N_15507,N_19247);
xor U23134 (N_23134,N_18879,N_17115);
nand U23135 (N_23135,N_15701,N_19252);
and U23136 (N_23136,N_18714,N_19795);
xor U23137 (N_23137,N_19684,N_15326);
or U23138 (N_23138,N_18257,N_18182);
or U23139 (N_23139,N_19635,N_16493);
xor U23140 (N_23140,N_15512,N_18283);
nand U23141 (N_23141,N_18795,N_19201);
nor U23142 (N_23142,N_15381,N_19655);
or U23143 (N_23143,N_18234,N_19308);
and U23144 (N_23144,N_18094,N_15489);
nor U23145 (N_23145,N_19020,N_16987);
and U23146 (N_23146,N_16676,N_15517);
and U23147 (N_23147,N_15714,N_17605);
and U23148 (N_23148,N_19965,N_19088);
nor U23149 (N_23149,N_16472,N_15377);
or U23150 (N_23150,N_19938,N_17739);
and U23151 (N_23151,N_15520,N_16029);
nand U23152 (N_23152,N_18540,N_17712);
nor U23153 (N_23153,N_17728,N_19084);
or U23154 (N_23154,N_19772,N_19334);
nor U23155 (N_23155,N_18388,N_16199);
nor U23156 (N_23156,N_18993,N_19157);
xnor U23157 (N_23157,N_19992,N_17976);
and U23158 (N_23158,N_18250,N_16353);
nand U23159 (N_23159,N_16279,N_19122);
or U23160 (N_23160,N_19144,N_15617);
nand U23161 (N_23161,N_17906,N_18181);
nor U23162 (N_23162,N_15103,N_19753);
nor U23163 (N_23163,N_18937,N_19792);
xnor U23164 (N_23164,N_17747,N_16308);
and U23165 (N_23165,N_15813,N_18465);
or U23166 (N_23166,N_16099,N_18195);
nor U23167 (N_23167,N_19035,N_15900);
or U23168 (N_23168,N_18863,N_15347);
and U23169 (N_23169,N_17347,N_16831);
nor U23170 (N_23170,N_16414,N_15885);
or U23171 (N_23171,N_15393,N_17743);
nor U23172 (N_23172,N_17662,N_17417);
nor U23173 (N_23173,N_17256,N_18923);
nor U23174 (N_23174,N_17212,N_17877);
and U23175 (N_23175,N_17148,N_18107);
and U23176 (N_23176,N_19033,N_19017);
nand U23177 (N_23177,N_15968,N_16200);
nor U23178 (N_23178,N_18723,N_18354);
or U23179 (N_23179,N_18150,N_16352);
or U23180 (N_23180,N_16135,N_16361);
nor U23181 (N_23181,N_16694,N_15683);
nor U23182 (N_23182,N_15880,N_18335);
nand U23183 (N_23183,N_17668,N_19408);
nand U23184 (N_23184,N_19791,N_19194);
or U23185 (N_23185,N_17723,N_16735);
nand U23186 (N_23186,N_18691,N_17542);
or U23187 (N_23187,N_16814,N_16268);
and U23188 (N_23188,N_15600,N_16285);
and U23189 (N_23189,N_19108,N_16950);
xnor U23190 (N_23190,N_15031,N_15435);
nor U23191 (N_23191,N_17682,N_16473);
and U23192 (N_23192,N_17408,N_15205);
or U23193 (N_23193,N_17901,N_19799);
nor U23194 (N_23194,N_15588,N_15704);
and U23195 (N_23195,N_16478,N_16683);
nor U23196 (N_23196,N_16265,N_16065);
and U23197 (N_23197,N_18802,N_19570);
nand U23198 (N_23198,N_15048,N_16127);
and U23199 (N_23199,N_17320,N_18039);
and U23200 (N_23200,N_19585,N_18662);
nor U23201 (N_23201,N_19286,N_18374);
or U23202 (N_23202,N_15533,N_17798);
xnor U23203 (N_23203,N_16178,N_18163);
nor U23204 (N_23204,N_18799,N_19018);
and U23205 (N_23205,N_16842,N_19783);
or U23206 (N_23206,N_18678,N_17313);
or U23207 (N_23207,N_15207,N_17983);
nand U23208 (N_23208,N_17961,N_18906);
and U23209 (N_23209,N_19515,N_19503);
or U23210 (N_23210,N_19246,N_17141);
nor U23211 (N_23211,N_19418,N_19285);
nor U23212 (N_23212,N_17967,N_15798);
and U23213 (N_23213,N_19189,N_19029);
and U23214 (N_23214,N_17968,N_18182);
nor U23215 (N_23215,N_16551,N_17989);
nand U23216 (N_23216,N_18742,N_15649);
xnor U23217 (N_23217,N_18181,N_18503);
and U23218 (N_23218,N_17401,N_17790);
or U23219 (N_23219,N_16429,N_16400);
and U23220 (N_23220,N_19728,N_18018);
and U23221 (N_23221,N_16300,N_19326);
or U23222 (N_23222,N_16898,N_17129);
and U23223 (N_23223,N_15369,N_18693);
or U23224 (N_23224,N_18593,N_19176);
and U23225 (N_23225,N_17229,N_17629);
or U23226 (N_23226,N_15959,N_15912);
nor U23227 (N_23227,N_16764,N_16744);
or U23228 (N_23228,N_17092,N_18467);
and U23229 (N_23229,N_18070,N_16309);
nor U23230 (N_23230,N_19747,N_15299);
or U23231 (N_23231,N_18676,N_16200);
nand U23232 (N_23232,N_19900,N_16588);
and U23233 (N_23233,N_15924,N_18476);
and U23234 (N_23234,N_15084,N_18256);
nand U23235 (N_23235,N_19931,N_16889);
or U23236 (N_23236,N_18110,N_19145);
and U23237 (N_23237,N_19929,N_18765);
nand U23238 (N_23238,N_15460,N_19177);
and U23239 (N_23239,N_17201,N_18984);
and U23240 (N_23240,N_15820,N_16015);
and U23241 (N_23241,N_18451,N_16005);
xnor U23242 (N_23242,N_18575,N_15466);
and U23243 (N_23243,N_15853,N_19693);
nor U23244 (N_23244,N_17363,N_15981);
nand U23245 (N_23245,N_15481,N_18490);
and U23246 (N_23246,N_16941,N_18195);
and U23247 (N_23247,N_16724,N_19536);
and U23248 (N_23248,N_18406,N_17489);
nor U23249 (N_23249,N_16290,N_17199);
or U23250 (N_23250,N_19903,N_17055);
and U23251 (N_23251,N_16967,N_18310);
nand U23252 (N_23252,N_15069,N_15532);
and U23253 (N_23253,N_19108,N_18044);
xnor U23254 (N_23254,N_19116,N_16985);
or U23255 (N_23255,N_17948,N_17710);
nor U23256 (N_23256,N_17760,N_15787);
nand U23257 (N_23257,N_17995,N_18481);
nor U23258 (N_23258,N_17444,N_15611);
or U23259 (N_23259,N_19852,N_18597);
xor U23260 (N_23260,N_18367,N_16767);
nor U23261 (N_23261,N_19911,N_17545);
nand U23262 (N_23262,N_15175,N_18740);
and U23263 (N_23263,N_15250,N_19244);
and U23264 (N_23264,N_18713,N_19170);
and U23265 (N_23265,N_17585,N_15114);
nor U23266 (N_23266,N_18587,N_17984);
or U23267 (N_23267,N_17546,N_16341);
nand U23268 (N_23268,N_16741,N_19257);
nand U23269 (N_23269,N_17907,N_15331);
xor U23270 (N_23270,N_19081,N_18415);
and U23271 (N_23271,N_17311,N_19148);
nand U23272 (N_23272,N_18652,N_18779);
or U23273 (N_23273,N_16941,N_15855);
nand U23274 (N_23274,N_15073,N_19249);
xor U23275 (N_23275,N_18393,N_16436);
or U23276 (N_23276,N_17388,N_16820);
and U23277 (N_23277,N_19329,N_15996);
or U23278 (N_23278,N_19153,N_18720);
nor U23279 (N_23279,N_18139,N_19081);
nand U23280 (N_23280,N_19643,N_15238);
nor U23281 (N_23281,N_18053,N_18587);
nor U23282 (N_23282,N_15762,N_15686);
nor U23283 (N_23283,N_16239,N_16479);
and U23284 (N_23284,N_15211,N_18915);
nand U23285 (N_23285,N_15190,N_18625);
or U23286 (N_23286,N_19343,N_19352);
and U23287 (N_23287,N_19507,N_16103);
or U23288 (N_23288,N_16945,N_17179);
nand U23289 (N_23289,N_15608,N_17426);
or U23290 (N_23290,N_18012,N_19957);
or U23291 (N_23291,N_15613,N_19429);
or U23292 (N_23292,N_16304,N_15840);
nand U23293 (N_23293,N_16726,N_17804);
xor U23294 (N_23294,N_17860,N_18948);
nand U23295 (N_23295,N_18318,N_17522);
nand U23296 (N_23296,N_16706,N_17435);
or U23297 (N_23297,N_18100,N_17337);
nor U23298 (N_23298,N_17135,N_18593);
and U23299 (N_23299,N_17387,N_18147);
nor U23300 (N_23300,N_18470,N_17048);
nand U23301 (N_23301,N_18395,N_17551);
or U23302 (N_23302,N_18855,N_19336);
nor U23303 (N_23303,N_17710,N_16020);
nand U23304 (N_23304,N_18230,N_17100);
and U23305 (N_23305,N_16862,N_16741);
and U23306 (N_23306,N_17611,N_17788);
and U23307 (N_23307,N_18928,N_15314);
nand U23308 (N_23308,N_15814,N_15787);
and U23309 (N_23309,N_16751,N_18400);
nor U23310 (N_23310,N_15106,N_16171);
nor U23311 (N_23311,N_15807,N_15991);
nand U23312 (N_23312,N_16572,N_18374);
nand U23313 (N_23313,N_19095,N_15491);
xor U23314 (N_23314,N_17145,N_18767);
and U23315 (N_23315,N_19110,N_19574);
nand U23316 (N_23316,N_15523,N_18027);
nor U23317 (N_23317,N_19315,N_19735);
or U23318 (N_23318,N_16406,N_16736);
nand U23319 (N_23319,N_19093,N_15607);
nand U23320 (N_23320,N_18682,N_18044);
nand U23321 (N_23321,N_18308,N_16276);
nor U23322 (N_23322,N_15811,N_15307);
or U23323 (N_23323,N_17530,N_17736);
and U23324 (N_23324,N_16339,N_15168);
or U23325 (N_23325,N_16258,N_15208);
nand U23326 (N_23326,N_15635,N_18944);
nand U23327 (N_23327,N_19315,N_18776);
and U23328 (N_23328,N_18999,N_17634);
and U23329 (N_23329,N_16753,N_18589);
nand U23330 (N_23330,N_17182,N_17575);
xor U23331 (N_23331,N_15503,N_18377);
or U23332 (N_23332,N_18646,N_18765);
nor U23333 (N_23333,N_19662,N_19765);
or U23334 (N_23334,N_17371,N_19683);
or U23335 (N_23335,N_15934,N_18767);
nor U23336 (N_23336,N_15879,N_19862);
or U23337 (N_23337,N_19500,N_15731);
nand U23338 (N_23338,N_18493,N_17193);
nand U23339 (N_23339,N_16177,N_17968);
or U23340 (N_23340,N_16365,N_17669);
nand U23341 (N_23341,N_16853,N_17371);
nand U23342 (N_23342,N_18298,N_16080);
nor U23343 (N_23343,N_16388,N_17706);
nor U23344 (N_23344,N_15083,N_19215);
nand U23345 (N_23345,N_19982,N_15294);
nand U23346 (N_23346,N_18978,N_19103);
xor U23347 (N_23347,N_15629,N_16038);
and U23348 (N_23348,N_16589,N_19334);
and U23349 (N_23349,N_15284,N_19052);
nor U23350 (N_23350,N_17531,N_18313);
nand U23351 (N_23351,N_17884,N_15052);
nor U23352 (N_23352,N_18136,N_16647);
and U23353 (N_23353,N_18722,N_17834);
nand U23354 (N_23354,N_15217,N_15799);
and U23355 (N_23355,N_17235,N_16992);
nand U23356 (N_23356,N_17373,N_18664);
or U23357 (N_23357,N_15932,N_17435);
or U23358 (N_23358,N_19105,N_19405);
nor U23359 (N_23359,N_19183,N_15335);
and U23360 (N_23360,N_16138,N_19842);
or U23361 (N_23361,N_18240,N_16955);
and U23362 (N_23362,N_16937,N_16194);
nor U23363 (N_23363,N_16367,N_16020);
nor U23364 (N_23364,N_15279,N_16016);
nor U23365 (N_23365,N_15972,N_19109);
and U23366 (N_23366,N_16197,N_18069);
or U23367 (N_23367,N_16174,N_16274);
and U23368 (N_23368,N_15584,N_16853);
nand U23369 (N_23369,N_17915,N_17517);
nor U23370 (N_23370,N_16405,N_16719);
xnor U23371 (N_23371,N_17798,N_17038);
and U23372 (N_23372,N_19956,N_16427);
or U23373 (N_23373,N_16454,N_17716);
nand U23374 (N_23374,N_18954,N_16401);
nor U23375 (N_23375,N_19808,N_17613);
nor U23376 (N_23376,N_18454,N_17598);
and U23377 (N_23377,N_15723,N_16965);
or U23378 (N_23378,N_15157,N_15456);
or U23379 (N_23379,N_19012,N_15619);
and U23380 (N_23380,N_16142,N_15970);
and U23381 (N_23381,N_18138,N_18516);
nor U23382 (N_23382,N_16867,N_17356);
or U23383 (N_23383,N_16762,N_15221);
xor U23384 (N_23384,N_16228,N_17180);
and U23385 (N_23385,N_15514,N_16693);
nand U23386 (N_23386,N_17660,N_19444);
or U23387 (N_23387,N_16258,N_18409);
and U23388 (N_23388,N_17001,N_19831);
or U23389 (N_23389,N_16394,N_16546);
and U23390 (N_23390,N_16026,N_17537);
nand U23391 (N_23391,N_18941,N_16598);
or U23392 (N_23392,N_15159,N_19067);
nor U23393 (N_23393,N_17896,N_16016);
xor U23394 (N_23394,N_18924,N_16786);
nor U23395 (N_23395,N_15724,N_18749);
nand U23396 (N_23396,N_17072,N_16584);
nor U23397 (N_23397,N_19277,N_19411);
and U23398 (N_23398,N_17819,N_16230);
nand U23399 (N_23399,N_15214,N_18592);
xor U23400 (N_23400,N_18144,N_18478);
nor U23401 (N_23401,N_15464,N_17702);
or U23402 (N_23402,N_18621,N_16182);
and U23403 (N_23403,N_19720,N_19738);
and U23404 (N_23404,N_15820,N_15115);
or U23405 (N_23405,N_16540,N_16000);
nor U23406 (N_23406,N_16846,N_16719);
nand U23407 (N_23407,N_19718,N_15721);
and U23408 (N_23408,N_16227,N_18300);
or U23409 (N_23409,N_18584,N_16168);
and U23410 (N_23410,N_15812,N_17547);
nand U23411 (N_23411,N_16032,N_17023);
or U23412 (N_23412,N_15471,N_16670);
xor U23413 (N_23413,N_19888,N_17874);
nor U23414 (N_23414,N_19456,N_18157);
or U23415 (N_23415,N_18782,N_19447);
nor U23416 (N_23416,N_15508,N_17389);
nor U23417 (N_23417,N_18294,N_16419);
or U23418 (N_23418,N_17262,N_17367);
or U23419 (N_23419,N_18549,N_18255);
and U23420 (N_23420,N_18083,N_18865);
or U23421 (N_23421,N_16857,N_17262);
nand U23422 (N_23422,N_17633,N_15292);
xor U23423 (N_23423,N_15909,N_15848);
nor U23424 (N_23424,N_19566,N_19811);
nand U23425 (N_23425,N_19196,N_15983);
xor U23426 (N_23426,N_19042,N_19713);
nor U23427 (N_23427,N_19932,N_18468);
and U23428 (N_23428,N_16013,N_15633);
nand U23429 (N_23429,N_15644,N_18341);
or U23430 (N_23430,N_18654,N_18534);
nand U23431 (N_23431,N_18739,N_19105);
or U23432 (N_23432,N_19621,N_18609);
or U23433 (N_23433,N_17679,N_16745);
and U23434 (N_23434,N_16360,N_17506);
nor U23435 (N_23435,N_17153,N_17859);
and U23436 (N_23436,N_17570,N_18574);
xor U23437 (N_23437,N_19633,N_17639);
nand U23438 (N_23438,N_17476,N_19258);
and U23439 (N_23439,N_18674,N_18907);
nor U23440 (N_23440,N_18780,N_18392);
nand U23441 (N_23441,N_15456,N_18261);
or U23442 (N_23442,N_15556,N_17596);
and U23443 (N_23443,N_16761,N_17279);
and U23444 (N_23444,N_17058,N_17405);
nor U23445 (N_23445,N_19169,N_17129);
and U23446 (N_23446,N_17684,N_17915);
nor U23447 (N_23447,N_16766,N_15758);
and U23448 (N_23448,N_16135,N_18302);
nor U23449 (N_23449,N_19285,N_19937);
nor U23450 (N_23450,N_19770,N_15482);
nand U23451 (N_23451,N_16465,N_18350);
nand U23452 (N_23452,N_19748,N_16725);
nand U23453 (N_23453,N_19697,N_18450);
nor U23454 (N_23454,N_18592,N_17769);
and U23455 (N_23455,N_19061,N_16654);
nor U23456 (N_23456,N_17287,N_15120);
xor U23457 (N_23457,N_16414,N_19115);
nand U23458 (N_23458,N_16260,N_19328);
nand U23459 (N_23459,N_18299,N_19685);
nand U23460 (N_23460,N_19121,N_16473);
nor U23461 (N_23461,N_17284,N_15152);
nand U23462 (N_23462,N_17867,N_16392);
and U23463 (N_23463,N_18042,N_18597);
nor U23464 (N_23464,N_15126,N_16166);
nand U23465 (N_23465,N_15028,N_17728);
or U23466 (N_23466,N_18827,N_15981);
or U23467 (N_23467,N_19209,N_16673);
and U23468 (N_23468,N_17162,N_18225);
nand U23469 (N_23469,N_17098,N_17845);
or U23470 (N_23470,N_18263,N_15131);
nand U23471 (N_23471,N_16346,N_19040);
nor U23472 (N_23472,N_17393,N_16159);
and U23473 (N_23473,N_16281,N_16663);
nor U23474 (N_23474,N_16228,N_15645);
and U23475 (N_23475,N_18372,N_18701);
nor U23476 (N_23476,N_19680,N_18966);
nand U23477 (N_23477,N_16899,N_19269);
nor U23478 (N_23478,N_15262,N_19851);
and U23479 (N_23479,N_19904,N_15720);
or U23480 (N_23480,N_17618,N_15879);
nand U23481 (N_23481,N_16471,N_17952);
or U23482 (N_23482,N_18036,N_19673);
nor U23483 (N_23483,N_17121,N_16687);
nor U23484 (N_23484,N_17032,N_19364);
nor U23485 (N_23485,N_17871,N_16025);
or U23486 (N_23486,N_16746,N_16250);
and U23487 (N_23487,N_18193,N_15652);
nand U23488 (N_23488,N_18287,N_19498);
and U23489 (N_23489,N_16536,N_17013);
nor U23490 (N_23490,N_17884,N_15942);
and U23491 (N_23491,N_19335,N_17313);
or U23492 (N_23492,N_15692,N_19319);
nand U23493 (N_23493,N_19015,N_17760);
and U23494 (N_23494,N_17287,N_17772);
nor U23495 (N_23495,N_16633,N_15154);
or U23496 (N_23496,N_16346,N_16277);
nor U23497 (N_23497,N_15643,N_16787);
xor U23498 (N_23498,N_18836,N_17895);
xnor U23499 (N_23499,N_17168,N_18382);
xnor U23500 (N_23500,N_18994,N_19777);
or U23501 (N_23501,N_15850,N_17162);
xnor U23502 (N_23502,N_17665,N_18545);
xnor U23503 (N_23503,N_18531,N_18795);
xor U23504 (N_23504,N_19994,N_17826);
nor U23505 (N_23505,N_17941,N_15559);
and U23506 (N_23506,N_15521,N_17400);
nand U23507 (N_23507,N_15845,N_19443);
and U23508 (N_23508,N_18846,N_18397);
nand U23509 (N_23509,N_19618,N_18893);
or U23510 (N_23510,N_17219,N_17386);
or U23511 (N_23511,N_17447,N_16176);
nor U23512 (N_23512,N_16128,N_15765);
nand U23513 (N_23513,N_18471,N_17831);
or U23514 (N_23514,N_16870,N_19848);
and U23515 (N_23515,N_19241,N_19133);
and U23516 (N_23516,N_19399,N_19077);
and U23517 (N_23517,N_15594,N_19711);
nor U23518 (N_23518,N_19582,N_17969);
or U23519 (N_23519,N_17631,N_15733);
nor U23520 (N_23520,N_16809,N_17096);
xor U23521 (N_23521,N_16839,N_18721);
or U23522 (N_23522,N_19114,N_18300);
nor U23523 (N_23523,N_19379,N_16815);
or U23524 (N_23524,N_17423,N_19837);
nor U23525 (N_23525,N_16921,N_18496);
xnor U23526 (N_23526,N_15590,N_18242);
nand U23527 (N_23527,N_16730,N_17596);
xnor U23528 (N_23528,N_19566,N_17080);
and U23529 (N_23529,N_18613,N_19433);
and U23530 (N_23530,N_16852,N_15499);
nor U23531 (N_23531,N_15759,N_15240);
nor U23532 (N_23532,N_19308,N_17193);
or U23533 (N_23533,N_17838,N_17361);
xnor U23534 (N_23534,N_15899,N_19166);
and U23535 (N_23535,N_19467,N_19094);
or U23536 (N_23536,N_18492,N_16711);
nand U23537 (N_23537,N_19057,N_16736);
xnor U23538 (N_23538,N_15451,N_19354);
or U23539 (N_23539,N_17004,N_19483);
nand U23540 (N_23540,N_19228,N_19545);
or U23541 (N_23541,N_17387,N_17030);
and U23542 (N_23542,N_15958,N_18320);
and U23543 (N_23543,N_15076,N_15449);
xor U23544 (N_23544,N_16038,N_19537);
nor U23545 (N_23545,N_17449,N_16259);
nand U23546 (N_23546,N_19174,N_18207);
and U23547 (N_23547,N_17731,N_15557);
nand U23548 (N_23548,N_15406,N_17521);
nand U23549 (N_23549,N_19029,N_17908);
nand U23550 (N_23550,N_18154,N_19178);
xor U23551 (N_23551,N_19016,N_18341);
and U23552 (N_23552,N_19366,N_18900);
and U23553 (N_23553,N_19354,N_18011);
xnor U23554 (N_23554,N_19765,N_16109);
and U23555 (N_23555,N_19783,N_19378);
nand U23556 (N_23556,N_15323,N_15259);
and U23557 (N_23557,N_15551,N_17173);
and U23558 (N_23558,N_18915,N_18393);
nor U23559 (N_23559,N_15248,N_17327);
or U23560 (N_23560,N_15162,N_18131);
nand U23561 (N_23561,N_16909,N_18706);
nand U23562 (N_23562,N_15172,N_16256);
and U23563 (N_23563,N_18289,N_19600);
nor U23564 (N_23564,N_18933,N_18190);
nor U23565 (N_23565,N_17842,N_19501);
or U23566 (N_23566,N_16871,N_16341);
and U23567 (N_23567,N_16071,N_15305);
nand U23568 (N_23568,N_17106,N_15859);
nand U23569 (N_23569,N_17761,N_15878);
nor U23570 (N_23570,N_17000,N_17035);
xnor U23571 (N_23571,N_16828,N_15350);
and U23572 (N_23572,N_15009,N_18554);
and U23573 (N_23573,N_16914,N_17174);
or U23574 (N_23574,N_15459,N_18910);
nor U23575 (N_23575,N_18209,N_19816);
or U23576 (N_23576,N_16912,N_16904);
and U23577 (N_23577,N_17218,N_17363);
or U23578 (N_23578,N_16697,N_16499);
or U23579 (N_23579,N_15130,N_15481);
and U23580 (N_23580,N_16467,N_18165);
and U23581 (N_23581,N_19922,N_19250);
xor U23582 (N_23582,N_17418,N_17857);
nand U23583 (N_23583,N_15393,N_16626);
and U23584 (N_23584,N_18066,N_16949);
or U23585 (N_23585,N_18321,N_17057);
and U23586 (N_23586,N_18781,N_19884);
or U23587 (N_23587,N_17389,N_15901);
and U23588 (N_23588,N_19522,N_19093);
or U23589 (N_23589,N_19708,N_15046);
or U23590 (N_23590,N_18589,N_17267);
or U23591 (N_23591,N_19040,N_19910);
nor U23592 (N_23592,N_17365,N_15320);
nand U23593 (N_23593,N_15385,N_15581);
nor U23594 (N_23594,N_17902,N_15650);
and U23595 (N_23595,N_16454,N_16704);
nand U23596 (N_23596,N_17135,N_15075);
or U23597 (N_23597,N_16980,N_19752);
and U23598 (N_23598,N_19617,N_16164);
nand U23599 (N_23599,N_15940,N_18191);
nand U23600 (N_23600,N_17441,N_19010);
nor U23601 (N_23601,N_15107,N_16185);
and U23602 (N_23602,N_17883,N_18532);
xnor U23603 (N_23603,N_17154,N_16717);
nand U23604 (N_23604,N_17634,N_15088);
and U23605 (N_23605,N_17346,N_19929);
or U23606 (N_23606,N_16256,N_18634);
or U23607 (N_23607,N_15138,N_16667);
or U23608 (N_23608,N_17201,N_17460);
nand U23609 (N_23609,N_16794,N_18476);
nor U23610 (N_23610,N_15646,N_19958);
nor U23611 (N_23611,N_19585,N_19487);
nand U23612 (N_23612,N_16182,N_15358);
or U23613 (N_23613,N_15992,N_18512);
nand U23614 (N_23614,N_16065,N_19611);
or U23615 (N_23615,N_19730,N_16931);
or U23616 (N_23616,N_18434,N_16971);
nor U23617 (N_23617,N_17095,N_15912);
or U23618 (N_23618,N_16766,N_16158);
and U23619 (N_23619,N_17221,N_19158);
or U23620 (N_23620,N_17372,N_18141);
xnor U23621 (N_23621,N_18577,N_19765);
nor U23622 (N_23622,N_19234,N_16422);
and U23623 (N_23623,N_16239,N_18654);
nor U23624 (N_23624,N_15168,N_15924);
and U23625 (N_23625,N_18651,N_16296);
or U23626 (N_23626,N_16037,N_17560);
and U23627 (N_23627,N_18496,N_16039);
nand U23628 (N_23628,N_19679,N_17016);
nand U23629 (N_23629,N_18870,N_16284);
or U23630 (N_23630,N_17074,N_19714);
nor U23631 (N_23631,N_17911,N_19751);
or U23632 (N_23632,N_19365,N_19216);
nand U23633 (N_23633,N_15224,N_17851);
and U23634 (N_23634,N_17263,N_17114);
and U23635 (N_23635,N_18697,N_16922);
nand U23636 (N_23636,N_16134,N_16523);
nand U23637 (N_23637,N_15662,N_19402);
nor U23638 (N_23638,N_15461,N_15499);
nand U23639 (N_23639,N_16420,N_16180);
or U23640 (N_23640,N_18480,N_17523);
or U23641 (N_23641,N_16027,N_18566);
or U23642 (N_23642,N_15459,N_18649);
nor U23643 (N_23643,N_18942,N_15060);
and U23644 (N_23644,N_16581,N_18290);
or U23645 (N_23645,N_18715,N_18729);
or U23646 (N_23646,N_18614,N_19803);
xnor U23647 (N_23647,N_16368,N_16476);
and U23648 (N_23648,N_17939,N_15694);
nand U23649 (N_23649,N_19088,N_15572);
nand U23650 (N_23650,N_17261,N_19830);
nor U23651 (N_23651,N_15050,N_17434);
xnor U23652 (N_23652,N_19951,N_18030);
nor U23653 (N_23653,N_19885,N_15038);
and U23654 (N_23654,N_18574,N_17020);
xor U23655 (N_23655,N_16942,N_19980);
nor U23656 (N_23656,N_16074,N_19138);
and U23657 (N_23657,N_19064,N_19026);
or U23658 (N_23658,N_19028,N_15450);
nor U23659 (N_23659,N_18765,N_18848);
nand U23660 (N_23660,N_15601,N_15284);
nand U23661 (N_23661,N_15633,N_16337);
or U23662 (N_23662,N_15208,N_18482);
or U23663 (N_23663,N_19259,N_15840);
nand U23664 (N_23664,N_19311,N_15643);
and U23665 (N_23665,N_19196,N_16436);
nand U23666 (N_23666,N_19148,N_18113);
or U23667 (N_23667,N_19532,N_17665);
or U23668 (N_23668,N_18534,N_17629);
or U23669 (N_23669,N_15860,N_18232);
and U23670 (N_23670,N_16088,N_19043);
nand U23671 (N_23671,N_16213,N_16123);
nor U23672 (N_23672,N_17410,N_19403);
and U23673 (N_23673,N_15202,N_19998);
and U23674 (N_23674,N_18730,N_16427);
and U23675 (N_23675,N_18460,N_19719);
or U23676 (N_23676,N_19464,N_15413);
nor U23677 (N_23677,N_19055,N_16589);
and U23678 (N_23678,N_18037,N_15313);
or U23679 (N_23679,N_17643,N_15253);
nor U23680 (N_23680,N_15225,N_17270);
nand U23681 (N_23681,N_18580,N_19606);
nor U23682 (N_23682,N_15189,N_16144);
nand U23683 (N_23683,N_19109,N_16753);
and U23684 (N_23684,N_19347,N_16431);
and U23685 (N_23685,N_16125,N_19187);
and U23686 (N_23686,N_17356,N_16662);
nand U23687 (N_23687,N_18823,N_17144);
nand U23688 (N_23688,N_17872,N_16997);
or U23689 (N_23689,N_18771,N_19827);
or U23690 (N_23690,N_16098,N_16139);
nor U23691 (N_23691,N_18116,N_16093);
nor U23692 (N_23692,N_19301,N_15884);
and U23693 (N_23693,N_17037,N_17613);
or U23694 (N_23694,N_19463,N_19810);
xnor U23695 (N_23695,N_15056,N_18603);
and U23696 (N_23696,N_17669,N_15037);
nor U23697 (N_23697,N_18754,N_18259);
xnor U23698 (N_23698,N_18389,N_18596);
and U23699 (N_23699,N_17400,N_18674);
or U23700 (N_23700,N_17905,N_16281);
and U23701 (N_23701,N_19381,N_18394);
and U23702 (N_23702,N_17860,N_17066);
or U23703 (N_23703,N_17334,N_19183);
nor U23704 (N_23704,N_15930,N_15299);
nor U23705 (N_23705,N_18886,N_15237);
nor U23706 (N_23706,N_15465,N_17602);
nor U23707 (N_23707,N_16396,N_19481);
and U23708 (N_23708,N_16942,N_15817);
or U23709 (N_23709,N_18759,N_18732);
or U23710 (N_23710,N_16605,N_16574);
or U23711 (N_23711,N_15839,N_19907);
nor U23712 (N_23712,N_18748,N_17781);
nand U23713 (N_23713,N_15070,N_19080);
and U23714 (N_23714,N_17255,N_19589);
nor U23715 (N_23715,N_19468,N_19072);
or U23716 (N_23716,N_17477,N_18366);
nor U23717 (N_23717,N_17700,N_18116);
and U23718 (N_23718,N_18735,N_19709);
nor U23719 (N_23719,N_19379,N_17402);
nor U23720 (N_23720,N_19793,N_15473);
xnor U23721 (N_23721,N_15342,N_17273);
nor U23722 (N_23722,N_15110,N_16815);
nor U23723 (N_23723,N_17915,N_15946);
nor U23724 (N_23724,N_19141,N_17075);
and U23725 (N_23725,N_16949,N_15171);
nor U23726 (N_23726,N_18419,N_17161);
xor U23727 (N_23727,N_17377,N_16701);
and U23728 (N_23728,N_18226,N_18760);
nand U23729 (N_23729,N_18566,N_17260);
nor U23730 (N_23730,N_17356,N_18489);
or U23731 (N_23731,N_19105,N_17373);
or U23732 (N_23732,N_16740,N_15081);
and U23733 (N_23733,N_16617,N_16744);
xnor U23734 (N_23734,N_18460,N_15527);
nor U23735 (N_23735,N_19741,N_19918);
or U23736 (N_23736,N_16364,N_17162);
or U23737 (N_23737,N_18323,N_18521);
nand U23738 (N_23738,N_18582,N_18308);
xnor U23739 (N_23739,N_16704,N_16696);
nand U23740 (N_23740,N_18787,N_15582);
nand U23741 (N_23741,N_17357,N_19388);
nand U23742 (N_23742,N_18356,N_17092);
nand U23743 (N_23743,N_15606,N_15400);
xor U23744 (N_23744,N_17819,N_19030);
nor U23745 (N_23745,N_16767,N_16870);
xor U23746 (N_23746,N_17775,N_18138);
or U23747 (N_23747,N_15801,N_17135);
nor U23748 (N_23748,N_16210,N_17571);
or U23749 (N_23749,N_19378,N_15451);
nor U23750 (N_23750,N_18024,N_18665);
nand U23751 (N_23751,N_16110,N_19124);
nor U23752 (N_23752,N_18863,N_15475);
or U23753 (N_23753,N_15629,N_16207);
nand U23754 (N_23754,N_15823,N_16344);
and U23755 (N_23755,N_18356,N_17254);
and U23756 (N_23756,N_18815,N_17461);
or U23757 (N_23757,N_18088,N_16463);
nand U23758 (N_23758,N_17266,N_19427);
nor U23759 (N_23759,N_17467,N_15825);
nor U23760 (N_23760,N_17370,N_18368);
nor U23761 (N_23761,N_19544,N_18108);
xnor U23762 (N_23762,N_16977,N_17119);
or U23763 (N_23763,N_19015,N_17107);
nor U23764 (N_23764,N_17340,N_19196);
nor U23765 (N_23765,N_18779,N_18041);
xor U23766 (N_23766,N_16785,N_16556);
xnor U23767 (N_23767,N_18941,N_18217);
xnor U23768 (N_23768,N_15813,N_15346);
nor U23769 (N_23769,N_17796,N_18897);
nand U23770 (N_23770,N_17902,N_16670);
nor U23771 (N_23771,N_16466,N_17841);
nor U23772 (N_23772,N_18183,N_19589);
and U23773 (N_23773,N_19717,N_18667);
and U23774 (N_23774,N_16570,N_19779);
or U23775 (N_23775,N_18632,N_18015);
nand U23776 (N_23776,N_17484,N_15195);
or U23777 (N_23777,N_19464,N_15486);
nand U23778 (N_23778,N_15158,N_19274);
nor U23779 (N_23779,N_15689,N_17451);
and U23780 (N_23780,N_15925,N_18127);
nand U23781 (N_23781,N_19426,N_16522);
and U23782 (N_23782,N_18506,N_17781);
nand U23783 (N_23783,N_19311,N_17524);
and U23784 (N_23784,N_19216,N_19583);
nand U23785 (N_23785,N_16308,N_18322);
nor U23786 (N_23786,N_19700,N_15198);
nor U23787 (N_23787,N_19121,N_17778);
nor U23788 (N_23788,N_17235,N_15023);
nand U23789 (N_23789,N_17098,N_17223);
nand U23790 (N_23790,N_19456,N_19870);
and U23791 (N_23791,N_15673,N_19043);
nand U23792 (N_23792,N_16915,N_18825);
nor U23793 (N_23793,N_18760,N_15482);
and U23794 (N_23794,N_15354,N_19225);
or U23795 (N_23795,N_18467,N_18933);
nor U23796 (N_23796,N_19089,N_19759);
and U23797 (N_23797,N_15647,N_17959);
xnor U23798 (N_23798,N_17635,N_17197);
nand U23799 (N_23799,N_15367,N_16316);
nand U23800 (N_23800,N_19072,N_18555);
or U23801 (N_23801,N_19526,N_15283);
or U23802 (N_23802,N_17508,N_19372);
nand U23803 (N_23803,N_15126,N_16109);
or U23804 (N_23804,N_16732,N_17494);
nor U23805 (N_23805,N_15158,N_19588);
nand U23806 (N_23806,N_17761,N_18882);
and U23807 (N_23807,N_15773,N_16373);
and U23808 (N_23808,N_18750,N_17594);
nor U23809 (N_23809,N_16524,N_16652);
nor U23810 (N_23810,N_15218,N_19994);
and U23811 (N_23811,N_17659,N_18345);
and U23812 (N_23812,N_15772,N_16867);
nand U23813 (N_23813,N_19360,N_19902);
and U23814 (N_23814,N_19657,N_19603);
nand U23815 (N_23815,N_18237,N_15282);
or U23816 (N_23816,N_17317,N_15196);
or U23817 (N_23817,N_16195,N_18580);
nand U23818 (N_23818,N_17025,N_16639);
nor U23819 (N_23819,N_16859,N_15935);
nor U23820 (N_23820,N_18382,N_16680);
or U23821 (N_23821,N_19961,N_17918);
xor U23822 (N_23822,N_17006,N_18806);
nand U23823 (N_23823,N_17083,N_16849);
nand U23824 (N_23824,N_16932,N_16957);
nand U23825 (N_23825,N_15788,N_19454);
nand U23826 (N_23826,N_19976,N_19704);
and U23827 (N_23827,N_19550,N_19328);
and U23828 (N_23828,N_18720,N_15984);
and U23829 (N_23829,N_18347,N_17432);
nor U23830 (N_23830,N_15909,N_17257);
and U23831 (N_23831,N_16523,N_16285);
or U23832 (N_23832,N_16858,N_18071);
nor U23833 (N_23833,N_19084,N_17276);
and U23834 (N_23834,N_17013,N_18423);
and U23835 (N_23835,N_18090,N_17304);
or U23836 (N_23836,N_17320,N_15279);
and U23837 (N_23837,N_15354,N_17709);
nand U23838 (N_23838,N_18495,N_16448);
nor U23839 (N_23839,N_15205,N_17673);
or U23840 (N_23840,N_17347,N_16738);
nand U23841 (N_23841,N_18502,N_15057);
and U23842 (N_23842,N_19027,N_19088);
xnor U23843 (N_23843,N_18316,N_18726);
nor U23844 (N_23844,N_16860,N_19597);
and U23845 (N_23845,N_16631,N_15489);
or U23846 (N_23846,N_18863,N_15411);
and U23847 (N_23847,N_17569,N_17011);
nor U23848 (N_23848,N_16431,N_17228);
or U23849 (N_23849,N_18653,N_19012);
nor U23850 (N_23850,N_18011,N_16023);
and U23851 (N_23851,N_16536,N_16383);
or U23852 (N_23852,N_15332,N_18689);
nand U23853 (N_23853,N_16032,N_16710);
nor U23854 (N_23854,N_17252,N_17515);
nor U23855 (N_23855,N_16526,N_15823);
and U23856 (N_23856,N_15756,N_16543);
or U23857 (N_23857,N_15423,N_15992);
nor U23858 (N_23858,N_18942,N_18309);
and U23859 (N_23859,N_15323,N_15604);
nor U23860 (N_23860,N_16170,N_16123);
nor U23861 (N_23861,N_15570,N_16492);
nand U23862 (N_23862,N_19822,N_17842);
nand U23863 (N_23863,N_15329,N_19131);
or U23864 (N_23864,N_16465,N_19756);
nand U23865 (N_23865,N_15535,N_18570);
or U23866 (N_23866,N_15412,N_17617);
or U23867 (N_23867,N_15526,N_16564);
xor U23868 (N_23868,N_19218,N_17004);
nor U23869 (N_23869,N_17551,N_15871);
and U23870 (N_23870,N_16042,N_15927);
and U23871 (N_23871,N_16043,N_15040);
and U23872 (N_23872,N_16207,N_16310);
nand U23873 (N_23873,N_18292,N_17468);
nand U23874 (N_23874,N_15346,N_15769);
and U23875 (N_23875,N_15078,N_19650);
and U23876 (N_23876,N_18378,N_16326);
xor U23877 (N_23877,N_19775,N_18556);
nor U23878 (N_23878,N_18777,N_17469);
xnor U23879 (N_23879,N_15086,N_17418);
nand U23880 (N_23880,N_16613,N_16318);
and U23881 (N_23881,N_18598,N_17204);
or U23882 (N_23882,N_16946,N_16807);
and U23883 (N_23883,N_17975,N_17650);
nand U23884 (N_23884,N_15293,N_15872);
nor U23885 (N_23885,N_15601,N_17009);
nor U23886 (N_23886,N_19025,N_16711);
nor U23887 (N_23887,N_15058,N_16212);
nor U23888 (N_23888,N_19362,N_19578);
and U23889 (N_23889,N_15868,N_18058);
and U23890 (N_23890,N_18089,N_18551);
and U23891 (N_23891,N_17159,N_16060);
nand U23892 (N_23892,N_17140,N_19412);
or U23893 (N_23893,N_18886,N_16354);
nor U23894 (N_23894,N_17833,N_16752);
nand U23895 (N_23895,N_15063,N_18962);
nand U23896 (N_23896,N_18157,N_16433);
and U23897 (N_23897,N_15463,N_19630);
or U23898 (N_23898,N_17001,N_16050);
and U23899 (N_23899,N_15939,N_17938);
xnor U23900 (N_23900,N_15360,N_16175);
or U23901 (N_23901,N_16667,N_15956);
nor U23902 (N_23902,N_19610,N_19874);
and U23903 (N_23903,N_18315,N_17679);
nand U23904 (N_23904,N_16604,N_19112);
nor U23905 (N_23905,N_17691,N_19219);
or U23906 (N_23906,N_18450,N_16008);
nand U23907 (N_23907,N_19376,N_17739);
or U23908 (N_23908,N_19395,N_18236);
nor U23909 (N_23909,N_17224,N_18819);
nand U23910 (N_23910,N_15218,N_15864);
and U23911 (N_23911,N_16545,N_16432);
and U23912 (N_23912,N_15238,N_16104);
nor U23913 (N_23913,N_16921,N_17067);
nor U23914 (N_23914,N_16955,N_18551);
or U23915 (N_23915,N_19871,N_15043);
nand U23916 (N_23916,N_19941,N_18036);
and U23917 (N_23917,N_15292,N_19661);
and U23918 (N_23918,N_18281,N_17968);
nor U23919 (N_23919,N_18432,N_17703);
or U23920 (N_23920,N_19565,N_18866);
nand U23921 (N_23921,N_17991,N_16463);
or U23922 (N_23922,N_16268,N_15186);
xor U23923 (N_23923,N_19576,N_19117);
and U23924 (N_23924,N_18046,N_18109);
or U23925 (N_23925,N_15526,N_17710);
xor U23926 (N_23926,N_16616,N_16051);
or U23927 (N_23927,N_18027,N_18236);
xor U23928 (N_23928,N_15488,N_17473);
or U23929 (N_23929,N_18101,N_15302);
and U23930 (N_23930,N_15303,N_18052);
or U23931 (N_23931,N_18243,N_19795);
nor U23932 (N_23932,N_18689,N_15925);
nor U23933 (N_23933,N_17847,N_18660);
nand U23934 (N_23934,N_19135,N_19036);
nand U23935 (N_23935,N_19362,N_19735);
and U23936 (N_23936,N_16535,N_18937);
nand U23937 (N_23937,N_18967,N_15530);
nand U23938 (N_23938,N_19573,N_18595);
nor U23939 (N_23939,N_18673,N_17490);
or U23940 (N_23940,N_19223,N_18912);
nand U23941 (N_23941,N_19180,N_15695);
nor U23942 (N_23942,N_16833,N_16135);
nand U23943 (N_23943,N_15831,N_18075);
and U23944 (N_23944,N_15164,N_16193);
nor U23945 (N_23945,N_15717,N_15334);
nand U23946 (N_23946,N_19499,N_19294);
xor U23947 (N_23947,N_16303,N_16075);
nand U23948 (N_23948,N_17857,N_19747);
or U23949 (N_23949,N_19295,N_16101);
nand U23950 (N_23950,N_18003,N_15389);
nand U23951 (N_23951,N_17343,N_17174);
or U23952 (N_23952,N_19478,N_16498);
nand U23953 (N_23953,N_18834,N_16842);
nor U23954 (N_23954,N_18397,N_17071);
nand U23955 (N_23955,N_15413,N_15184);
nor U23956 (N_23956,N_18813,N_17275);
and U23957 (N_23957,N_16597,N_18253);
nand U23958 (N_23958,N_18545,N_15727);
or U23959 (N_23959,N_17929,N_16921);
nor U23960 (N_23960,N_19944,N_16246);
and U23961 (N_23961,N_15287,N_18632);
or U23962 (N_23962,N_16739,N_19613);
nand U23963 (N_23963,N_19529,N_19895);
or U23964 (N_23964,N_19655,N_18812);
xor U23965 (N_23965,N_17955,N_17981);
xnor U23966 (N_23966,N_15627,N_18351);
nor U23967 (N_23967,N_18547,N_16342);
nor U23968 (N_23968,N_15993,N_19745);
xnor U23969 (N_23969,N_18005,N_18826);
xor U23970 (N_23970,N_15623,N_16066);
and U23971 (N_23971,N_16918,N_15635);
nand U23972 (N_23972,N_16449,N_15209);
nor U23973 (N_23973,N_15954,N_16918);
nor U23974 (N_23974,N_17600,N_16277);
nand U23975 (N_23975,N_18014,N_17962);
and U23976 (N_23976,N_16179,N_18767);
nor U23977 (N_23977,N_16513,N_18693);
nor U23978 (N_23978,N_17024,N_15975);
nand U23979 (N_23979,N_19070,N_16575);
or U23980 (N_23980,N_18297,N_15891);
nand U23981 (N_23981,N_18785,N_19831);
nor U23982 (N_23982,N_16158,N_18069);
and U23983 (N_23983,N_16742,N_19178);
nor U23984 (N_23984,N_17297,N_17105);
nand U23985 (N_23985,N_16802,N_19049);
nand U23986 (N_23986,N_17996,N_17843);
nand U23987 (N_23987,N_19337,N_17449);
nand U23988 (N_23988,N_17701,N_15289);
nand U23989 (N_23989,N_18116,N_15698);
and U23990 (N_23990,N_15883,N_17938);
nand U23991 (N_23991,N_19176,N_15580);
or U23992 (N_23992,N_17234,N_19511);
or U23993 (N_23993,N_17810,N_18026);
and U23994 (N_23994,N_19305,N_19749);
or U23995 (N_23995,N_19924,N_18661);
or U23996 (N_23996,N_16211,N_18641);
nor U23997 (N_23997,N_18802,N_16587);
nand U23998 (N_23998,N_18416,N_15976);
or U23999 (N_23999,N_19429,N_16011);
nor U24000 (N_24000,N_18685,N_18787);
and U24001 (N_24001,N_18117,N_17359);
nor U24002 (N_24002,N_19687,N_16722);
or U24003 (N_24003,N_19410,N_17544);
and U24004 (N_24004,N_16356,N_16946);
nor U24005 (N_24005,N_16239,N_15889);
nand U24006 (N_24006,N_19071,N_16799);
nor U24007 (N_24007,N_18193,N_16985);
xor U24008 (N_24008,N_18747,N_18725);
and U24009 (N_24009,N_19728,N_18305);
nor U24010 (N_24010,N_18262,N_19492);
or U24011 (N_24011,N_17386,N_15240);
nor U24012 (N_24012,N_19839,N_17418);
nor U24013 (N_24013,N_19839,N_16691);
or U24014 (N_24014,N_17832,N_15163);
or U24015 (N_24015,N_15106,N_18535);
or U24016 (N_24016,N_17494,N_18149);
or U24017 (N_24017,N_16062,N_17651);
nand U24018 (N_24018,N_15241,N_16448);
and U24019 (N_24019,N_16813,N_19403);
or U24020 (N_24020,N_17196,N_15972);
xor U24021 (N_24021,N_18255,N_16794);
nor U24022 (N_24022,N_17061,N_19238);
nand U24023 (N_24023,N_16599,N_16624);
or U24024 (N_24024,N_18156,N_19036);
and U24025 (N_24025,N_17923,N_15586);
nand U24026 (N_24026,N_18777,N_19618);
and U24027 (N_24027,N_19880,N_16379);
and U24028 (N_24028,N_17687,N_17866);
nor U24029 (N_24029,N_15819,N_16365);
nor U24030 (N_24030,N_18837,N_17287);
nor U24031 (N_24031,N_16312,N_16835);
and U24032 (N_24032,N_17371,N_19951);
nand U24033 (N_24033,N_17378,N_15760);
or U24034 (N_24034,N_19033,N_18093);
or U24035 (N_24035,N_19234,N_17817);
nor U24036 (N_24036,N_17050,N_17041);
nor U24037 (N_24037,N_15457,N_19433);
nand U24038 (N_24038,N_19084,N_16651);
nand U24039 (N_24039,N_16480,N_18801);
nand U24040 (N_24040,N_19110,N_18198);
or U24041 (N_24041,N_16525,N_19785);
or U24042 (N_24042,N_15940,N_15784);
and U24043 (N_24043,N_16753,N_18984);
or U24044 (N_24044,N_15598,N_15172);
xnor U24045 (N_24045,N_19444,N_15342);
nor U24046 (N_24046,N_16303,N_16090);
or U24047 (N_24047,N_19199,N_16042);
and U24048 (N_24048,N_15416,N_18279);
nor U24049 (N_24049,N_17844,N_16109);
nor U24050 (N_24050,N_18389,N_15892);
or U24051 (N_24051,N_15577,N_18045);
xnor U24052 (N_24052,N_15470,N_17491);
nand U24053 (N_24053,N_16117,N_15053);
and U24054 (N_24054,N_19115,N_15000);
xor U24055 (N_24055,N_19632,N_15874);
and U24056 (N_24056,N_15800,N_17241);
or U24057 (N_24057,N_19493,N_16443);
nand U24058 (N_24058,N_16566,N_16241);
nor U24059 (N_24059,N_16829,N_18879);
or U24060 (N_24060,N_16873,N_17711);
nand U24061 (N_24061,N_15556,N_17422);
or U24062 (N_24062,N_15669,N_15134);
nor U24063 (N_24063,N_19401,N_19561);
and U24064 (N_24064,N_19099,N_18869);
nand U24065 (N_24065,N_15517,N_18459);
nor U24066 (N_24066,N_17377,N_19570);
nand U24067 (N_24067,N_15453,N_15275);
nor U24068 (N_24068,N_19746,N_16111);
xnor U24069 (N_24069,N_17317,N_16460);
and U24070 (N_24070,N_15057,N_16856);
nand U24071 (N_24071,N_17410,N_19328);
nor U24072 (N_24072,N_17036,N_16771);
nor U24073 (N_24073,N_18682,N_16296);
nor U24074 (N_24074,N_17269,N_19808);
and U24075 (N_24075,N_15618,N_19435);
xnor U24076 (N_24076,N_15937,N_16673);
nor U24077 (N_24077,N_17795,N_17576);
or U24078 (N_24078,N_16402,N_19189);
or U24079 (N_24079,N_15645,N_18318);
nor U24080 (N_24080,N_16342,N_17429);
xor U24081 (N_24081,N_18674,N_18954);
nor U24082 (N_24082,N_19910,N_15896);
nand U24083 (N_24083,N_15541,N_16210);
and U24084 (N_24084,N_19318,N_17764);
nor U24085 (N_24085,N_17769,N_15873);
nand U24086 (N_24086,N_18266,N_18236);
nor U24087 (N_24087,N_19668,N_15992);
and U24088 (N_24088,N_17263,N_16411);
nand U24089 (N_24089,N_16404,N_17464);
xor U24090 (N_24090,N_16072,N_15392);
nor U24091 (N_24091,N_19483,N_19452);
or U24092 (N_24092,N_19993,N_15745);
nor U24093 (N_24093,N_17324,N_19818);
or U24094 (N_24094,N_16125,N_19242);
and U24095 (N_24095,N_17089,N_18635);
or U24096 (N_24096,N_15745,N_15197);
or U24097 (N_24097,N_15753,N_17927);
nor U24098 (N_24098,N_19999,N_17635);
or U24099 (N_24099,N_17462,N_16906);
nand U24100 (N_24100,N_17914,N_16884);
nor U24101 (N_24101,N_16750,N_16063);
nor U24102 (N_24102,N_17528,N_16245);
nor U24103 (N_24103,N_16385,N_17971);
and U24104 (N_24104,N_15102,N_18050);
nand U24105 (N_24105,N_18876,N_15942);
or U24106 (N_24106,N_18800,N_18467);
or U24107 (N_24107,N_17794,N_17352);
nand U24108 (N_24108,N_15901,N_19520);
xnor U24109 (N_24109,N_19913,N_19261);
and U24110 (N_24110,N_17721,N_17502);
and U24111 (N_24111,N_15807,N_16406);
xor U24112 (N_24112,N_18051,N_15050);
or U24113 (N_24113,N_17820,N_15667);
xnor U24114 (N_24114,N_15183,N_15834);
or U24115 (N_24115,N_17528,N_19429);
or U24116 (N_24116,N_17272,N_19219);
nor U24117 (N_24117,N_16066,N_16202);
nand U24118 (N_24118,N_17347,N_15976);
and U24119 (N_24119,N_17705,N_15683);
xnor U24120 (N_24120,N_15946,N_17423);
nand U24121 (N_24121,N_19446,N_16909);
nor U24122 (N_24122,N_15387,N_18817);
xor U24123 (N_24123,N_17360,N_16323);
and U24124 (N_24124,N_18838,N_19842);
nor U24125 (N_24125,N_15816,N_19835);
and U24126 (N_24126,N_16639,N_16707);
nor U24127 (N_24127,N_15992,N_19612);
or U24128 (N_24128,N_19671,N_18641);
nand U24129 (N_24129,N_19638,N_16075);
nand U24130 (N_24130,N_17915,N_16338);
nor U24131 (N_24131,N_15505,N_15907);
or U24132 (N_24132,N_15257,N_15737);
nand U24133 (N_24133,N_17560,N_19320);
nand U24134 (N_24134,N_15551,N_18025);
and U24135 (N_24135,N_16684,N_19630);
xnor U24136 (N_24136,N_18838,N_19202);
nor U24137 (N_24137,N_16113,N_19025);
and U24138 (N_24138,N_17574,N_17315);
nor U24139 (N_24139,N_16984,N_19228);
nand U24140 (N_24140,N_18839,N_18913);
nand U24141 (N_24141,N_18355,N_19253);
and U24142 (N_24142,N_15667,N_16209);
and U24143 (N_24143,N_16447,N_15041);
or U24144 (N_24144,N_16180,N_18512);
nand U24145 (N_24145,N_19481,N_18102);
xnor U24146 (N_24146,N_19239,N_15758);
nor U24147 (N_24147,N_15233,N_16401);
nand U24148 (N_24148,N_15006,N_18816);
xnor U24149 (N_24149,N_19609,N_15981);
xnor U24150 (N_24150,N_17824,N_16534);
nor U24151 (N_24151,N_18674,N_19687);
nor U24152 (N_24152,N_17966,N_16522);
nor U24153 (N_24153,N_18754,N_17452);
nand U24154 (N_24154,N_15654,N_19869);
or U24155 (N_24155,N_15865,N_18971);
nor U24156 (N_24156,N_17647,N_15048);
nor U24157 (N_24157,N_18721,N_19080);
and U24158 (N_24158,N_15449,N_18691);
and U24159 (N_24159,N_15060,N_17659);
nor U24160 (N_24160,N_16252,N_19222);
nor U24161 (N_24161,N_16053,N_18883);
nand U24162 (N_24162,N_16974,N_17987);
xnor U24163 (N_24163,N_17502,N_16334);
nor U24164 (N_24164,N_17452,N_16360);
nand U24165 (N_24165,N_16477,N_18809);
and U24166 (N_24166,N_16450,N_15811);
and U24167 (N_24167,N_18516,N_18006);
and U24168 (N_24168,N_15860,N_18167);
nor U24169 (N_24169,N_18200,N_18480);
nor U24170 (N_24170,N_15298,N_16916);
or U24171 (N_24171,N_19533,N_19207);
or U24172 (N_24172,N_19476,N_16111);
nand U24173 (N_24173,N_17558,N_15497);
xnor U24174 (N_24174,N_17627,N_17357);
nor U24175 (N_24175,N_17968,N_17103);
xnor U24176 (N_24176,N_19324,N_19649);
and U24177 (N_24177,N_17695,N_19608);
nor U24178 (N_24178,N_16422,N_17645);
nor U24179 (N_24179,N_18634,N_17487);
nand U24180 (N_24180,N_17244,N_17022);
and U24181 (N_24181,N_15731,N_15761);
nand U24182 (N_24182,N_19235,N_15186);
nor U24183 (N_24183,N_16713,N_18240);
and U24184 (N_24184,N_18766,N_17281);
nand U24185 (N_24185,N_18470,N_18633);
and U24186 (N_24186,N_18790,N_18843);
nand U24187 (N_24187,N_17552,N_17940);
nand U24188 (N_24188,N_18656,N_18119);
nor U24189 (N_24189,N_18238,N_18877);
xor U24190 (N_24190,N_16374,N_17011);
nor U24191 (N_24191,N_15596,N_17842);
nand U24192 (N_24192,N_17950,N_15469);
nor U24193 (N_24193,N_18450,N_18588);
nor U24194 (N_24194,N_16213,N_15248);
and U24195 (N_24195,N_15900,N_18881);
or U24196 (N_24196,N_16587,N_19792);
nor U24197 (N_24197,N_16361,N_19312);
nand U24198 (N_24198,N_19180,N_16099);
nand U24199 (N_24199,N_15727,N_15949);
nor U24200 (N_24200,N_17726,N_18353);
or U24201 (N_24201,N_17070,N_16077);
or U24202 (N_24202,N_18460,N_15911);
nor U24203 (N_24203,N_16535,N_18994);
nor U24204 (N_24204,N_17612,N_16730);
xnor U24205 (N_24205,N_17739,N_15656);
and U24206 (N_24206,N_18379,N_17143);
or U24207 (N_24207,N_17337,N_18363);
nand U24208 (N_24208,N_18877,N_17145);
or U24209 (N_24209,N_17764,N_16274);
nor U24210 (N_24210,N_19208,N_18642);
xnor U24211 (N_24211,N_18828,N_17067);
nand U24212 (N_24212,N_18774,N_17556);
and U24213 (N_24213,N_15756,N_15054);
xnor U24214 (N_24214,N_19483,N_18391);
xnor U24215 (N_24215,N_17538,N_16209);
xnor U24216 (N_24216,N_16283,N_17152);
xor U24217 (N_24217,N_15171,N_16407);
or U24218 (N_24218,N_16577,N_15515);
or U24219 (N_24219,N_19075,N_18520);
and U24220 (N_24220,N_15286,N_15665);
nand U24221 (N_24221,N_19233,N_19658);
xor U24222 (N_24222,N_15809,N_15031);
nor U24223 (N_24223,N_16463,N_16251);
or U24224 (N_24224,N_17150,N_16800);
and U24225 (N_24225,N_17492,N_18976);
nor U24226 (N_24226,N_17207,N_18829);
and U24227 (N_24227,N_18836,N_15225);
nor U24228 (N_24228,N_18525,N_19641);
xor U24229 (N_24229,N_17978,N_15235);
and U24230 (N_24230,N_18984,N_17717);
or U24231 (N_24231,N_18250,N_19868);
xor U24232 (N_24232,N_17733,N_16325);
or U24233 (N_24233,N_17151,N_17476);
or U24234 (N_24234,N_18523,N_15654);
nor U24235 (N_24235,N_15512,N_17063);
nor U24236 (N_24236,N_16930,N_18434);
nand U24237 (N_24237,N_19266,N_16696);
nor U24238 (N_24238,N_17160,N_15211);
or U24239 (N_24239,N_17785,N_16571);
nor U24240 (N_24240,N_16675,N_19191);
or U24241 (N_24241,N_17235,N_19291);
nor U24242 (N_24242,N_16600,N_19076);
or U24243 (N_24243,N_19027,N_19853);
nand U24244 (N_24244,N_19592,N_17597);
xor U24245 (N_24245,N_17940,N_17265);
and U24246 (N_24246,N_16979,N_16339);
nand U24247 (N_24247,N_19353,N_19857);
and U24248 (N_24248,N_17275,N_19284);
nor U24249 (N_24249,N_15876,N_16357);
xor U24250 (N_24250,N_18668,N_19330);
nand U24251 (N_24251,N_17963,N_17546);
and U24252 (N_24252,N_16086,N_18306);
nor U24253 (N_24253,N_19705,N_16981);
or U24254 (N_24254,N_19509,N_19960);
nor U24255 (N_24255,N_16392,N_17890);
nor U24256 (N_24256,N_19965,N_19869);
or U24257 (N_24257,N_15333,N_18431);
nand U24258 (N_24258,N_18757,N_16276);
and U24259 (N_24259,N_16706,N_16464);
and U24260 (N_24260,N_15962,N_17091);
and U24261 (N_24261,N_17778,N_19924);
or U24262 (N_24262,N_17845,N_16431);
or U24263 (N_24263,N_15711,N_18226);
nor U24264 (N_24264,N_19365,N_19499);
or U24265 (N_24265,N_19335,N_19619);
or U24266 (N_24266,N_16814,N_15805);
nor U24267 (N_24267,N_15262,N_16316);
or U24268 (N_24268,N_18765,N_15072);
xnor U24269 (N_24269,N_15419,N_15087);
or U24270 (N_24270,N_17352,N_19233);
or U24271 (N_24271,N_15054,N_19151);
and U24272 (N_24272,N_18123,N_17398);
or U24273 (N_24273,N_16144,N_17559);
nand U24274 (N_24274,N_17376,N_18859);
and U24275 (N_24275,N_19401,N_16370);
nor U24276 (N_24276,N_17748,N_19826);
or U24277 (N_24277,N_17919,N_15041);
nor U24278 (N_24278,N_17821,N_17937);
nand U24279 (N_24279,N_15508,N_16725);
or U24280 (N_24280,N_15001,N_19848);
and U24281 (N_24281,N_19853,N_17564);
and U24282 (N_24282,N_17079,N_18310);
and U24283 (N_24283,N_15681,N_17087);
or U24284 (N_24284,N_18828,N_16018);
nor U24285 (N_24285,N_15775,N_17895);
nor U24286 (N_24286,N_16691,N_18859);
or U24287 (N_24287,N_16796,N_15474);
xnor U24288 (N_24288,N_15267,N_15414);
nor U24289 (N_24289,N_15859,N_17786);
nor U24290 (N_24290,N_18789,N_16183);
nand U24291 (N_24291,N_17369,N_18615);
nor U24292 (N_24292,N_19999,N_15554);
and U24293 (N_24293,N_18517,N_18771);
and U24294 (N_24294,N_19607,N_15439);
xnor U24295 (N_24295,N_17821,N_15397);
xor U24296 (N_24296,N_17527,N_19304);
xor U24297 (N_24297,N_18863,N_19354);
nor U24298 (N_24298,N_19337,N_19266);
and U24299 (N_24299,N_16148,N_19978);
nor U24300 (N_24300,N_19449,N_15155);
and U24301 (N_24301,N_18278,N_15089);
and U24302 (N_24302,N_17350,N_18986);
and U24303 (N_24303,N_15521,N_19834);
and U24304 (N_24304,N_19468,N_15988);
and U24305 (N_24305,N_18477,N_15780);
and U24306 (N_24306,N_17631,N_15365);
nor U24307 (N_24307,N_19225,N_17264);
and U24308 (N_24308,N_19240,N_19374);
xnor U24309 (N_24309,N_17340,N_19926);
nand U24310 (N_24310,N_16017,N_17469);
xnor U24311 (N_24311,N_15205,N_15378);
nor U24312 (N_24312,N_18696,N_17513);
xor U24313 (N_24313,N_15352,N_15109);
or U24314 (N_24314,N_19512,N_19547);
and U24315 (N_24315,N_17775,N_15793);
and U24316 (N_24316,N_15752,N_15751);
or U24317 (N_24317,N_15831,N_19847);
xor U24318 (N_24318,N_15078,N_15981);
xnor U24319 (N_24319,N_18221,N_16263);
nor U24320 (N_24320,N_16416,N_15875);
and U24321 (N_24321,N_16978,N_15974);
xnor U24322 (N_24322,N_18304,N_19899);
nor U24323 (N_24323,N_18953,N_16410);
or U24324 (N_24324,N_17828,N_19521);
or U24325 (N_24325,N_15614,N_16988);
or U24326 (N_24326,N_17525,N_17901);
nand U24327 (N_24327,N_16615,N_18815);
and U24328 (N_24328,N_17229,N_15679);
nand U24329 (N_24329,N_17836,N_17088);
or U24330 (N_24330,N_19182,N_15949);
nand U24331 (N_24331,N_17404,N_19031);
and U24332 (N_24332,N_17408,N_19157);
nor U24333 (N_24333,N_16960,N_18164);
xor U24334 (N_24334,N_17421,N_18981);
nor U24335 (N_24335,N_19491,N_16097);
nand U24336 (N_24336,N_16434,N_17452);
xor U24337 (N_24337,N_18090,N_18392);
nand U24338 (N_24338,N_19662,N_18616);
or U24339 (N_24339,N_16459,N_16674);
nand U24340 (N_24340,N_16315,N_15603);
nand U24341 (N_24341,N_18510,N_16188);
nor U24342 (N_24342,N_18753,N_19577);
nand U24343 (N_24343,N_17212,N_18445);
nand U24344 (N_24344,N_15218,N_16824);
and U24345 (N_24345,N_18046,N_15380);
nor U24346 (N_24346,N_18970,N_19489);
nor U24347 (N_24347,N_16075,N_19668);
or U24348 (N_24348,N_19664,N_19266);
nand U24349 (N_24349,N_15590,N_19602);
nand U24350 (N_24350,N_17997,N_18519);
nor U24351 (N_24351,N_17406,N_16173);
and U24352 (N_24352,N_17696,N_16697);
nand U24353 (N_24353,N_18641,N_18738);
and U24354 (N_24354,N_17576,N_18047);
or U24355 (N_24355,N_15214,N_16227);
nand U24356 (N_24356,N_16130,N_17276);
xor U24357 (N_24357,N_16561,N_19265);
nand U24358 (N_24358,N_18479,N_19132);
and U24359 (N_24359,N_16236,N_18396);
nor U24360 (N_24360,N_18334,N_19475);
nor U24361 (N_24361,N_15153,N_16830);
nand U24362 (N_24362,N_17446,N_15227);
and U24363 (N_24363,N_16751,N_18247);
nor U24364 (N_24364,N_17237,N_19923);
and U24365 (N_24365,N_15230,N_17408);
nand U24366 (N_24366,N_16891,N_18536);
nand U24367 (N_24367,N_17813,N_19198);
nand U24368 (N_24368,N_15338,N_15098);
or U24369 (N_24369,N_15878,N_15482);
nor U24370 (N_24370,N_19227,N_19578);
nor U24371 (N_24371,N_19087,N_16445);
nand U24372 (N_24372,N_17442,N_15106);
nand U24373 (N_24373,N_18965,N_16082);
or U24374 (N_24374,N_15200,N_18472);
and U24375 (N_24375,N_18942,N_16669);
or U24376 (N_24376,N_19064,N_18174);
xor U24377 (N_24377,N_15811,N_15356);
and U24378 (N_24378,N_18218,N_17348);
nand U24379 (N_24379,N_15797,N_17298);
or U24380 (N_24380,N_19961,N_18305);
nand U24381 (N_24381,N_16446,N_18297);
xnor U24382 (N_24382,N_17319,N_18147);
and U24383 (N_24383,N_16403,N_16625);
nor U24384 (N_24384,N_18824,N_15845);
and U24385 (N_24385,N_15616,N_15270);
nor U24386 (N_24386,N_19003,N_16880);
xor U24387 (N_24387,N_17102,N_16930);
and U24388 (N_24388,N_15513,N_17079);
or U24389 (N_24389,N_19460,N_17278);
nor U24390 (N_24390,N_18799,N_19200);
or U24391 (N_24391,N_19893,N_16414);
and U24392 (N_24392,N_18461,N_19965);
and U24393 (N_24393,N_16880,N_19667);
xor U24394 (N_24394,N_16635,N_16247);
nor U24395 (N_24395,N_15503,N_18186);
xnor U24396 (N_24396,N_16452,N_17212);
and U24397 (N_24397,N_17337,N_17315);
and U24398 (N_24398,N_15986,N_16911);
nand U24399 (N_24399,N_17962,N_15945);
nor U24400 (N_24400,N_15793,N_16985);
or U24401 (N_24401,N_16793,N_16870);
or U24402 (N_24402,N_18151,N_16910);
or U24403 (N_24403,N_17967,N_17205);
and U24404 (N_24404,N_19893,N_17741);
nor U24405 (N_24405,N_16117,N_19901);
and U24406 (N_24406,N_18732,N_19669);
or U24407 (N_24407,N_16992,N_15800);
xnor U24408 (N_24408,N_19284,N_19952);
or U24409 (N_24409,N_16518,N_16622);
xnor U24410 (N_24410,N_17968,N_19221);
nand U24411 (N_24411,N_15834,N_18066);
or U24412 (N_24412,N_19842,N_15219);
or U24413 (N_24413,N_17276,N_15609);
xnor U24414 (N_24414,N_17029,N_15434);
nand U24415 (N_24415,N_15820,N_16035);
or U24416 (N_24416,N_18918,N_17357);
nand U24417 (N_24417,N_19779,N_18942);
nor U24418 (N_24418,N_16931,N_19503);
and U24419 (N_24419,N_16875,N_16981);
xor U24420 (N_24420,N_17329,N_17066);
nand U24421 (N_24421,N_15651,N_16187);
nand U24422 (N_24422,N_16786,N_16833);
and U24423 (N_24423,N_19828,N_15778);
nand U24424 (N_24424,N_17559,N_18148);
nor U24425 (N_24425,N_18080,N_16819);
or U24426 (N_24426,N_19001,N_19073);
nand U24427 (N_24427,N_18341,N_17504);
or U24428 (N_24428,N_17600,N_18020);
or U24429 (N_24429,N_15174,N_16991);
xor U24430 (N_24430,N_16396,N_18067);
xor U24431 (N_24431,N_16487,N_15319);
or U24432 (N_24432,N_16746,N_15369);
and U24433 (N_24433,N_15527,N_16475);
and U24434 (N_24434,N_19618,N_16542);
and U24435 (N_24435,N_18931,N_16286);
nor U24436 (N_24436,N_17230,N_18736);
and U24437 (N_24437,N_15029,N_17545);
or U24438 (N_24438,N_16669,N_15980);
and U24439 (N_24439,N_17628,N_15375);
nor U24440 (N_24440,N_19387,N_19657);
and U24441 (N_24441,N_15408,N_17433);
or U24442 (N_24442,N_17382,N_17185);
and U24443 (N_24443,N_17851,N_18877);
or U24444 (N_24444,N_17440,N_18933);
or U24445 (N_24445,N_19849,N_19185);
and U24446 (N_24446,N_16588,N_16919);
nor U24447 (N_24447,N_16734,N_16908);
and U24448 (N_24448,N_18343,N_18070);
or U24449 (N_24449,N_19738,N_19554);
or U24450 (N_24450,N_18899,N_18246);
or U24451 (N_24451,N_16762,N_15097);
and U24452 (N_24452,N_17388,N_17298);
nor U24453 (N_24453,N_15294,N_18622);
nand U24454 (N_24454,N_16712,N_16403);
or U24455 (N_24455,N_19114,N_18454);
and U24456 (N_24456,N_19097,N_15326);
nand U24457 (N_24457,N_18285,N_18610);
and U24458 (N_24458,N_17169,N_19771);
and U24459 (N_24459,N_17107,N_19057);
and U24460 (N_24460,N_19639,N_15507);
or U24461 (N_24461,N_17620,N_15705);
or U24462 (N_24462,N_18654,N_16442);
nor U24463 (N_24463,N_16237,N_19705);
and U24464 (N_24464,N_17509,N_18067);
xor U24465 (N_24465,N_19547,N_16415);
or U24466 (N_24466,N_16044,N_19615);
and U24467 (N_24467,N_17173,N_17413);
nor U24468 (N_24468,N_17085,N_18863);
nand U24469 (N_24469,N_18915,N_17255);
or U24470 (N_24470,N_18547,N_16261);
or U24471 (N_24471,N_17100,N_18811);
nor U24472 (N_24472,N_19289,N_19530);
and U24473 (N_24473,N_18136,N_15230);
nor U24474 (N_24474,N_17197,N_16886);
nor U24475 (N_24475,N_19034,N_18242);
xor U24476 (N_24476,N_19899,N_15501);
xor U24477 (N_24477,N_15545,N_18895);
nand U24478 (N_24478,N_18510,N_16558);
and U24479 (N_24479,N_17287,N_16147);
xor U24480 (N_24480,N_15318,N_18212);
xnor U24481 (N_24481,N_18165,N_19211);
and U24482 (N_24482,N_18335,N_18558);
nand U24483 (N_24483,N_15821,N_17213);
or U24484 (N_24484,N_17123,N_16756);
nand U24485 (N_24485,N_15266,N_15067);
nor U24486 (N_24486,N_17794,N_17829);
nand U24487 (N_24487,N_18447,N_17815);
nor U24488 (N_24488,N_16000,N_15403);
nor U24489 (N_24489,N_17269,N_16041);
nor U24490 (N_24490,N_19604,N_19911);
nor U24491 (N_24491,N_15499,N_15968);
nand U24492 (N_24492,N_18535,N_19944);
and U24493 (N_24493,N_17291,N_19609);
nand U24494 (N_24494,N_18361,N_18690);
and U24495 (N_24495,N_18129,N_18018);
nand U24496 (N_24496,N_16947,N_19441);
nand U24497 (N_24497,N_16665,N_17178);
and U24498 (N_24498,N_18672,N_18798);
xor U24499 (N_24499,N_17098,N_15999);
nor U24500 (N_24500,N_19987,N_15817);
nand U24501 (N_24501,N_17449,N_18875);
nor U24502 (N_24502,N_19539,N_19584);
nor U24503 (N_24503,N_16445,N_18124);
nor U24504 (N_24504,N_19657,N_16786);
nand U24505 (N_24505,N_19063,N_19166);
and U24506 (N_24506,N_19626,N_17904);
nand U24507 (N_24507,N_19684,N_18973);
and U24508 (N_24508,N_19044,N_19379);
or U24509 (N_24509,N_18855,N_17831);
xnor U24510 (N_24510,N_17929,N_16044);
nor U24511 (N_24511,N_15284,N_17400);
or U24512 (N_24512,N_18397,N_15675);
nand U24513 (N_24513,N_19879,N_18469);
and U24514 (N_24514,N_19880,N_16272);
or U24515 (N_24515,N_19737,N_17926);
xnor U24516 (N_24516,N_17054,N_16977);
and U24517 (N_24517,N_19174,N_17935);
nand U24518 (N_24518,N_19301,N_19305);
and U24519 (N_24519,N_19375,N_16978);
and U24520 (N_24520,N_16967,N_19962);
and U24521 (N_24521,N_16205,N_19666);
nor U24522 (N_24522,N_17597,N_15345);
nor U24523 (N_24523,N_17104,N_18315);
nand U24524 (N_24524,N_17562,N_16409);
nand U24525 (N_24525,N_19871,N_19489);
nor U24526 (N_24526,N_19002,N_17307);
or U24527 (N_24527,N_19917,N_17091);
nand U24528 (N_24528,N_15234,N_19226);
and U24529 (N_24529,N_19566,N_18422);
nor U24530 (N_24530,N_16149,N_17206);
or U24531 (N_24531,N_16337,N_18046);
or U24532 (N_24532,N_18192,N_16977);
nor U24533 (N_24533,N_15764,N_17309);
nor U24534 (N_24534,N_19040,N_19275);
and U24535 (N_24535,N_18251,N_15252);
nor U24536 (N_24536,N_15391,N_15137);
or U24537 (N_24537,N_15168,N_16932);
and U24538 (N_24538,N_19479,N_16594);
nor U24539 (N_24539,N_19341,N_19964);
nand U24540 (N_24540,N_15479,N_15523);
and U24541 (N_24541,N_17378,N_18873);
nand U24542 (N_24542,N_15547,N_18164);
nor U24543 (N_24543,N_16341,N_15474);
nand U24544 (N_24544,N_17827,N_17753);
and U24545 (N_24545,N_19512,N_16675);
and U24546 (N_24546,N_18600,N_17595);
nand U24547 (N_24547,N_17205,N_19404);
nor U24548 (N_24548,N_16251,N_18583);
or U24549 (N_24549,N_19410,N_16567);
nand U24550 (N_24550,N_18029,N_16588);
and U24551 (N_24551,N_19225,N_18940);
and U24552 (N_24552,N_17003,N_18061);
or U24553 (N_24553,N_16363,N_18870);
nor U24554 (N_24554,N_17022,N_15325);
or U24555 (N_24555,N_17361,N_19658);
and U24556 (N_24556,N_16696,N_19886);
nand U24557 (N_24557,N_15944,N_18771);
and U24558 (N_24558,N_18620,N_17596);
nor U24559 (N_24559,N_15190,N_16912);
nor U24560 (N_24560,N_19632,N_18189);
xor U24561 (N_24561,N_18032,N_15183);
or U24562 (N_24562,N_16274,N_16988);
or U24563 (N_24563,N_16069,N_16341);
nor U24564 (N_24564,N_18464,N_15064);
nor U24565 (N_24565,N_16544,N_15954);
or U24566 (N_24566,N_18193,N_16926);
and U24567 (N_24567,N_17686,N_19794);
nand U24568 (N_24568,N_18494,N_16338);
or U24569 (N_24569,N_17888,N_15662);
nand U24570 (N_24570,N_17230,N_16394);
or U24571 (N_24571,N_18064,N_15156);
or U24572 (N_24572,N_17648,N_19377);
and U24573 (N_24573,N_19499,N_15358);
nand U24574 (N_24574,N_16515,N_19900);
or U24575 (N_24575,N_19536,N_17651);
nor U24576 (N_24576,N_15945,N_17067);
nor U24577 (N_24577,N_18669,N_16584);
xnor U24578 (N_24578,N_16809,N_15385);
or U24579 (N_24579,N_19296,N_19978);
or U24580 (N_24580,N_16157,N_18161);
and U24581 (N_24581,N_15642,N_16524);
and U24582 (N_24582,N_16588,N_19348);
and U24583 (N_24583,N_19629,N_17207);
and U24584 (N_24584,N_18092,N_19347);
xor U24585 (N_24585,N_17610,N_17322);
xor U24586 (N_24586,N_16984,N_15664);
nor U24587 (N_24587,N_19542,N_16977);
and U24588 (N_24588,N_16192,N_15931);
and U24589 (N_24589,N_16178,N_19434);
nor U24590 (N_24590,N_15850,N_19862);
nor U24591 (N_24591,N_16671,N_19615);
and U24592 (N_24592,N_16771,N_17098);
or U24593 (N_24593,N_17544,N_16337);
nor U24594 (N_24594,N_19606,N_17063);
nand U24595 (N_24595,N_15534,N_16179);
or U24596 (N_24596,N_18334,N_15104);
nor U24597 (N_24597,N_19368,N_19473);
xor U24598 (N_24598,N_19855,N_19090);
and U24599 (N_24599,N_19706,N_15025);
nand U24600 (N_24600,N_17415,N_19201);
or U24601 (N_24601,N_15705,N_15906);
and U24602 (N_24602,N_19786,N_17187);
xor U24603 (N_24603,N_17684,N_15203);
nand U24604 (N_24604,N_17079,N_16208);
nand U24605 (N_24605,N_17867,N_15760);
nor U24606 (N_24606,N_15632,N_18619);
nor U24607 (N_24607,N_19556,N_15325);
or U24608 (N_24608,N_15029,N_19793);
nor U24609 (N_24609,N_15613,N_19219);
or U24610 (N_24610,N_16795,N_17085);
nor U24611 (N_24611,N_19214,N_18675);
nand U24612 (N_24612,N_19060,N_16758);
nor U24613 (N_24613,N_15280,N_18982);
nand U24614 (N_24614,N_15762,N_17435);
nor U24615 (N_24615,N_16122,N_15824);
nand U24616 (N_24616,N_15234,N_19002);
nor U24617 (N_24617,N_18350,N_17292);
nor U24618 (N_24618,N_19057,N_17024);
or U24619 (N_24619,N_15038,N_16355);
nor U24620 (N_24620,N_15213,N_17943);
xnor U24621 (N_24621,N_18021,N_19720);
nor U24622 (N_24622,N_16105,N_16274);
nor U24623 (N_24623,N_15707,N_15907);
nand U24624 (N_24624,N_15763,N_18550);
xor U24625 (N_24625,N_15427,N_18744);
and U24626 (N_24626,N_19787,N_16434);
nor U24627 (N_24627,N_17139,N_16132);
or U24628 (N_24628,N_16182,N_15696);
nand U24629 (N_24629,N_17782,N_18226);
and U24630 (N_24630,N_15143,N_16500);
nor U24631 (N_24631,N_16280,N_17874);
nor U24632 (N_24632,N_16917,N_18149);
nand U24633 (N_24633,N_17073,N_16668);
and U24634 (N_24634,N_16293,N_15616);
nor U24635 (N_24635,N_15382,N_19633);
and U24636 (N_24636,N_17692,N_17469);
or U24637 (N_24637,N_16484,N_18315);
nor U24638 (N_24638,N_15301,N_17997);
or U24639 (N_24639,N_16067,N_17184);
nand U24640 (N_24640,N_15150,N_16802);
xor U24641 (N_24641,N_17250,N_15267);
nand U24642 (N_24642,N_17907,N_19489);
xor U24643 (N_24643,N_16821,N_18861);
and U24644 (N_24644,N_17153,N_17165);
or U24645 (N_24645,N_19256,N_15710);
and U24646 (N_24646,N_17842,N_19409);
nand U24647 (N_24647,N_17329,N_15426);
or U24648 (N_24648,N_15234,N_19394);
nor U24649 (N_24649,N_17019,N_15266);
nand U24650 (N_24650,N_19451,N_18837);
and U24651 (N_24651,N_16116,N_18374);
or U24652 (N_24652,N_17002,N_16934);
xnor U24653 (N_24653,N_17012,N_16078);
nand U24654 (N_24654,N_15417,N_15643);
and U24655 (N_24655,N_18048,N_18965);
and U24656 (N_24656,N_16071,N_15350);
xor U24657 (N_24657,N_16648,N_17021);
or U24658 (N_24658,N_18593,N_15058);
nand U24659 (N_24659,N_15557,N_17618);
nand U24660 (N_24660,N_15675,N_17895);
or U24661 (N_24661,N_15691,N_15533);
xnor U24662 (N_24662,N_19712,N_15656);
nor U24663 (N_24663,N_15641,N_16800);
nor U24664 (N_24664,N_16091,N_19384);
nand U24665 (N_24665,N_17199,N_16739);
or U24666 (N_24666,N_17840,N_19157);
nand U24667 (N_24667,N_17059,N_19825);
nand U24668 (N_24668,N_17831,N_16656);
or U24669 (N_24669,N_18917,N_16564);
and U24670 (N_24670,N_19059,N_16854);
nor U24671 (N_24671,N_15001,N_19549);
nand U24672 (N_24672,N_19778,N_18798);
nor U24673 (N_24673,N_17983,N_18177);
nor U24674 (N_24674,N_19199,N_19881);
nor U24675 (N_24675,N_18591,N_15179);
nor U24676 (N_24676,N_18695,N_18464);
nor U24677 (N_24677,N_19374,N_19746);
nand U24678 (N_24678,N_16508,N_18328);
nand U24679 (N_24679,N_16910,N_16714);
xor U24680 (N_24680,N_16929,N_19720);
nand U24681 (N_24681,N_19886,N_18870);
nor U24682 (N_24682,N_15961,N_16965);
or U24683 (N_24683,N_19715,N_17646);
nand U24684 (N_24684,N_17241,N_17215);
and U24685 (N_24685,N_15637,N_16369);
xnor U24686 (N_24686,N_17994,N_18208);
or U24687 (N_24687,N_16025,N_16297);
nor U24688 (N_24688,N_18271,N_16653);
and U24689 (N_24689,N_16932,N_16276);
xor U24690 (N_24690,N_15153,N_15866);
nand U24691 (N_24691,N_16895,N_17760);
and U24692 (N_24692,N_16500,N_16854);
or U24693 (N_24693,N_16208,N_16892);
xor U24694 (N_24694,N_17651,N_19113);
and U24695 (N_24695,N_16491,N_18751);
nor U24696 (N_24696,N_15198,N_15709);
nor U24697 (N_24697,N_19957,N_17934);
and U24698 (N_24698,N_19376,N_19110);
and U24699 (N_24699,N_16472,N_17558);
and U24700 (N_24700,N_16813,N_17347);
nor U24701 (N_24701,N_15551,N_16754);
nand U24702 (N_24702,N_16188,N_19381);
and U24703 (N_24703,N_17161,N_19252);
and U24704 (N_24704,N_15586,N_16997);
and U24705 (N_24705,N_17190,N_19155);
and U24706 (N_24706,N_16243,N_19003);
or U24707 (N_24707,N_15449,N_17619);
or U24708 (N_24708,N_19311,N_19117);
nor U24709 (N_24709,N_19746,N_16545);
and U24710 (N_24710,N_15226,N_18340);
or U24711 (N_24711,N_18221,N_17011);
or U24712 (N_24712,N_17714,N_15367);
nand U24713 (N_24713,N_16743,N_19417);
and U24714 (N_24714,N_17121,N_18622);
nor U24715 (N_24715,N_16838,N_18290);
nor U24716 (N_24716,N_16786,N_19166);
nand U24717 (N_24717,N_15248,N_17981);
or U24718 (N_24718,N_19379,N_15512);
and U24719 (N_24719,N_17202,N_15953);
or U24720 (N_24720,N_15051,N_17439);
or U24721 (N_24721,N_15994,N_15669);
xor U24722 (N_24722,N_16523,N_16958);
or U24723 (N_24723,N_16034,N_18375);
or U24724 (N_24724,N_16281,N_17684);
nor U24725 (N_24725,N_16500,N_19279);
or U24726 (N_24726,N_18505,N_17652);
and U24727 (N_24727,N_15040,N_16437);
nor U24728 (N_24728,N_19385,N_17456);
and U24729 (N_24729,N_15261,N_17209);
nor U24730 (N_24730,N_18267,N_18560);
nand U24731 (N_24731,N_16879,N_17838);
or U24732 (N_24732,N_16763,N_15890);
and U24733 (N_24733,N_17880,N_17178);
or U24734 (N_24734,N_15021,N_19599);
nor U24735 (N_24735,N_18406,N_19018);
nor U24736 (N_24736,N_16657,N_16020);
nand U24737 (N_24737,N_17566,N_15237);
or U24738 (N_24738,N_18749,N_17438);
and U24739 (N_24739,N_17180,N_18021);
nand U24740 (N_24740,N_17872,N_16019);
or U24741 (N_24741,N_17650,N_15043);
nand U24742 (N_24742,N_15182,N_17283);
and U24743 (N_24743,N_15866,N_19726);
nor U24744 (N_24744,N_16536,N_17000);
nor U24745 (N_24745,N_19734,N_18795);
nand U24746 (N_24746,N_15672,N_15714);
nor U24747 (N_24747,N_15752,N_19388);
nand U24748 (N_24748,N_16930,N_18345);
xor U24749 (N_24749,N_16160,N_16592);
or U24750 (N_24750,N_15227,N_18739);
nor U24751 (N_24751,N_16640,N_15590);
and U24752 (N_24752,N_16398,N_17576);
and U24753 (N_24753,N_18273,N_18297);
and U24754 (N_24754,N_18269,N_19861);
and U24755 (N_24755,N_18378,N_16396);
xor U24756 (N_24756,N_15310,N_16043);
nand U24757 (N_24757,N_18546,N_17936);
nand U24758 (N_24758,N_16551,N_15951);
nor U24759 (N_24759,N_16969,N_15257);
and U24760 (N_24760,N_15047,N_19738);
and U24761 (N_24761,N_16549,N_19901);
or U24762 (N_24762,N_18636,N_19625);
nand U24763 (N_24763,N_16579,N_18497);
or U24764 (N_24764,N_17077,N_19110);
nor U24765 (N_24765,N_17949,N_18714);
nor U24766 (N_24766,N_16663,N_16015);
nor U24767 (N_24767,N_17438,N_17262);
nand U24768 (N_24768,N_19337,N_15279);
or U24769 (N_24769,N_17285,N_17950);
and U24770 (N_24770,N_18389,N_19641);
and U24771 (N_24771,N_15228,N_16323);
and U24772 (N_24772,N_16450,N_16838);
xnor U24773 (N_24773,N_18959,N_17236);
nand U24774 (N_24774,N_15437,N_18477);
xor U24775 (N_24775,N_19572,N_16163);
or U24776 (N_24776,N_18305,N_15292);
and U24777 (N_24777,N_15200,N_17617);
nor U24778 (N_24778,N_19015,N_16435);
nand U24779 (N_24779,N_19487,N_16206);
or U24780 (N_24780,N_16314,N_19098);
xor U24781 (N_24781,N_15376,N_18496);
and U24782 (N_24782,N_16248,N_19330);
nor U24783 (N_24783,N_16321,N_19626);
nor U24784 (N_24784,N_16088,N_15278);
nand U24785 (N_24785,N_19256,N_17958);
nor U24786 (N_24786,N_16559,N_18891);
nand U24787 (N_24787,N_18422,N_19222);
and U24788 (N_24788,N_16276,N_17288);
or U24789 (N_24789,N_15139,N_17531);
nand U24790 (N_24790,N_18752,N_18916);
nand U24791 (N_24791,N_17595,N_16540);
nor U24792 (N_24792,N_18371,N_19846);
and U24793 (N_24793,N_15020,N_16238);
and U24794 (N_24794,N_15146,N_18557);
or U24795 (N_24795,N_18202,N_15223);
nand U24796 (N_24796,N_16559,N_15066);
and U24797 (N_24797,N_15696,N_19509);
or U24798 (N_24798,N_16650,N_15742);
and U24799 (N_24799,N_19484,N_16600);
nor U24800 (N_24800,N_16772,N_18821);
or U24801 (N_24801,N_18842,N_18139);
and U24802 (N_24802,N_19513,N_17802);
xnor U24803 (N_24803,N_15948,N_15018);
nand U24804 (N_24804,N_18497,N_19755);
nor U24805 (N_24805,N_18246,N_15208);
xnor U24806 (N_24806,N_18859,N_16581);
nor U24807 (N_24807,N_17215,N_18129);
and U24808 (N_24808,N_17192,N_17649);
xnor U24809 (N_24809,N_19674,N_19182);
or U24810 (N_24810,N_17752,N_16699);
or U24811 (N_24811,N_19893,N_16011);
nor U24812 (N_24812,N_16120,N_17150);
or U24813 (N_24813,N_15591,N_19915);
nor U24814 (N_24814,N_19873,N_16840);
and U24815 (N_24815,N_18872,N_19600);
nor U24816 (N_24816,N_17408,N_17956);
and U24817 (N_24817,N_18753,N_18380);
nand U24818 (N_24818,N_15992,N_15646);
or U24819 (N_24819,N_18806,N_16886);
and U24820 (N_24820,N_16211,N_19397);
xnor U24821 (N_24821,N_17842,N_15622);
and U24822 (N_24822,N_19643,N_16584);
and U24823 (N_24823,N_18090,N_19359);
and U24824 (N_24824,N_15556,N_17726);
and U24825 (N_24825,N_18147,N_16930);
nand U24826 (N_24826,N_16094,N_18662);
or U24827 (N_24827,N_15514,N_18840);
or U24828 (N_24828,N_15116,N_19369);
nand U24829 (N_24829,N_19652,N_16728);
or U24830 (N_24830,N_16566,N_18507);
nand U24831 (N_24831,N_17847,N_18884);
xnor U24832 (N_24832,N_18189,N_19902);
nand U24833 (N_24833,N_18474,N_18749);
xnor U24834 (N_24834,N_17613,N_16671);
nor U24835 (N_24835,N_19528,N_18708);
or U24836 (N_24836,N_16425,N_17536);
nand U24837 (N_24837,N_16515,N_16797);
nand U24838 (N_24838,N_15270,N_15375);
or U24839 (N_24839,N_17737,N_18227);
nand U24840 (N_24840,N_19575,N_17204);
nand U24841 (N_24841,N_17855,N_15972);
nor U24842 (N_24842,N_18701,N_16761);
and U24843 (N_24843,N_17128,N_18570);
nand U24844 (N_24844,N_16978,N_18787);
or U24845 (N_24845,N_19527,N_17608);
or U24846 (N_24846,N_19276,N_19427);
nand U24847 (N_24847,N_19319,N_18538);
xor U24848 (N_24848,N_19360,N_15164);
nand U24849 (N_24849,N_15556,N_18460);
and U24850 (N_24850,N_18261,N_17542);
nand U24851 (N_24851,N_19582,N_16166);
nand U24852 (N_24852,N_15181,N_15249);
nand U24853 (N_24853,N_16900,N_16934);
nand U24854 (N_24854,N_15478,N_16699);
and U24855 (N_24855,N_15770,N_15957);
or U24856 (N_24856,N_15917,N_16911);
and U24857 (N_24857,N_16576,N_17867);
nand U24858 (N_24858,N_18346,N_17562);
xor U24859 (N_24859,N_18730,N_17955);
nor U24860 (N_24860,N_16028,N_19076);
or U24861 (N_24861,N_18865,N_19395);
or U24862 (N_24862,N_18284,N_15392);
xnor U24863 (N_24863,N_19911,N_19301);
and U24864 (N_24864,N_18886,N_15389);
or U24865 (N_24865,N_17547,N_19921);
nor U24866 (N_24866,N_15785,N_18734);
nor U24867 (N_24867,N_17984,N_19204);
nor U24868 (N_24868,N_18436,N_17340);
or U24869 (N_24869,N_17233,N_19138);
or U24870 (N_24870,N_17046,N_19642);
or U24871 (N_24871,N_15432,N_16067);
nor U24872 (N_24872,N_16549,N_15756);
nor U24873 (N_24873,N_19844,N_17466);
nand U24874 (N_24874,N_15464,N_17971);
and U24875 (N_24875,N_18959,N_16341);
or U24876 (N_24876,N_18515,N_16286);
and U24877 (N_24877,N_18221,N_17628);
or U24878 (N_24878,N_15767,N_16680);
and U24879 (N_24879,N_18251,N_18498);
nand U24880 (N_24880,N_19982,N_17106);
nor U24881 (N_24881,N_18976,N_19189);
nand U24882 (N_24882,N_19458,N_15284);
xor U24883 (N_24883,N_15933,N_15441);
nor U24884 (N_24884,N_17246,N_15535);
or U24885 (N_24885,N_18050,N_15493);
nor U24886 (N_24886,N_15752,N_16908);
xnor U24887 (N_24887,N_16529,N_19745);
or U24888 (N_24888,N_15311,N_18638);
nor U24889 (N_24889,N_18112,N_16568);
or U24890 (N_24890,N_15207,N_17902);
xor U24891 (N_24891,N_16386,N_19246);
and U24892 (N_24892,N_17654,N_19733);
and U24893 (N_24893,N_17466,N_17388);
nand U24894 (N_24894,N_17020,N_16521);
nand U24895 (N_24895,N_16053,N_17572);
and U24896 (N_24896,N_15369,N_18863);
nor U24897 (N_24897,N_18313,N_15219);
or U24898 (N_24898,N_17613,N_17532);
nand U24899 (N_24899,N_19974,N_18008);
nand U24900 (N_24900,N_19489,N_16888);
nand U24901 (N_24901,N_16650,N_18257);
or U24902 (N_24902,N_15517,N_18576);
nor U24903 (N_24903,N_15010,N_17651);
nand U24904 (N_24904,N_15844,N_19084);
or U24905 (N_24905,N_17059,N_17154);
or U24906 (N_24906,N_19104,N_15107);
and U24907 (N_24907,N_15957,N_16247);
and U24908 (N_24908,N_18233,N_17193);
nor U24909 (N_24909,N_17914,N_18326);
xor U24910 (N_24910,N_18857,N_18260);
or U24911 (N_24911,N_16042,N_17962);
nand U24912 (N_24912,N_19794,N_16557);
or U24913 (N_24913,N_16778,N_15961);
nor U24914 (N_24914,N_16785,N_18905);
or U24915 (N_24915,N_18369,N_17182);
and U24916 (N_24916,N_18061,N_16202);
or U24917 (N_24917,N_18214,N_16253);
or U24918 (N_24918,N_17735,N_16695);
nor U24919 (N_24919,N_17027,N_16232);
nor U24920 (N_24920,N_19680,N_17563);
or U24921 (N_24921,N_19156,N_19871);
xor U24922 (N_24922,N_17240,N_16963);
or U24923 (N_24923,N_16283,N_19988);
nor U24924 (N_24924,N_18338,N_18556);
nand U24925 (N_24925,N_16823,N_16005);
and U24926 (N_24926,N_16834,N_17092);
xor U24927 (N_24927,N_16799,N_19362);
nand U24928 (N_24928,N_18979,N_18832);
xor U24929 (N_24929,N_17329,N_15891);
nor U24930 (N_24930,N_15559,N_15629);
nand U24931 (N_24931,N_18491,N_16451);
nand U24932 (N_24932,N_16438,N_19722);
and U24933 (N_24933,N_17505,N_16209);
and U24934 (N_24934,N_15479,N_16198);
nand U24935 (N_24935,N_17998,N_18504);
nand U24936 (N_24936,N_18653,N_18397);
and U24937 (N_24937,N_18287,N_17335);
nor U24938 (N_24938,N_18302,N_18960);
and U24939 (N_24939,N_19756,N_17110);
or U24940 (N_24940,N_17222,N_16589);
nor U24941 (N_24941,N_17885,N_15973);
or U24942 (N_24942,N_17347,N_17716);
nor U24943 (N_24943,N_19717,N_16329);
and U24944 (N_24944,N_17236,N_18881);
or U24945 (N_24945,N_17442,N_17051);
nand U24946 (N_24946,N_16134,N_16463);
or U24947 (N_24947,N_17427,N_19825);
nor U24948 (N_24948,N_17251,N_16265);
nor U24949 (N_24949,N_19045,N_16980);
nand U24950 (N_24950,N_19746,N_18982);
and U24951 (N_24951,N_17416,N_15810);
or U24952 (N_24952,N_18045,N_19022);
nor U24953 (N_24953,N_16453,N_17607);
xor U24954 (N_24954,N_17905,N_17659);
nor U24955 (N_24955,N_15847,N_16093);
or U24956 (N_24956,N_16719,N_17091);
nand U24957 (N_24957,N_16754,N_16546);
and U24958 (N_24958,N_19437,N_19040);
nor U24959 (N_24959,N_15520,N_18959);
nand U24960 (N_24960,N_18696,N_19495);
xor U24961 (N_24961,N_19523,N_15201);
xor U24962 (N_24962,N_19051,N_15767);
nand U24963 (N_24963,N_19781,N_18358);
nand U24964 (N_24964,N_15008,N_17778);
nor U24965 (N_24965,N_18618,N_19354);
and U24966 (N_24966,N_16500,N_19073);
nor U24967 (N_24967,N_19229,N_18633);
or U24968 (N_24968,N_17643,N_15375);
and U24969 (N_24969,N_16708,N_16669);
nand U24970 (N_24970,N_15857,N_18364);
or U24971 (N_24971,N_15984,N_19632);
xnor U24972 (N_24972,N_19587,N_19063);
nor U24973 (N_24973,N_15805,N_17623);
nor U24974 (N_24974,N_16972,N_15040);
and U24975 (N_24975,N_15513,N_16223);
xnor U24976 (N_24976,N_19059,N_19184);
and U24977 (N_24977,N_16341,N_16709);
or U24978 (N_24978,N_17710,N_17173);
or U24979 (N_24979,N_16526,N_17854);
and U24980 (N_24980,N_18806,N_16815);
and U24981 (N_24981,N_17379,N_16921);
or U24982 (N_24982,N_16370,N_17110);
nor U24983 (N_24983,N_16513,N_17489);
nor U24984 (N_24984,N_18913,N_15361);
and U24985 (N_24985,N_15744,N_16059);
or U24986 (N_24986,N_16547,N_19354);
and U24987 (N_24987,N_18362,N_18428);
nand U24988 (N_24988,N_16224,N_15231);
nor U24989 (N_24989,N_19042,N_15061);
or U24990 (N_24990,N_19419,N_17925);
nand U24991 (N_24991,N_15087,N_15966);
nor U24992 (N_24992,N_18374,N_18757);
nand U24993 (N_24993,N_18803,N_16450);
and U24994 (N_24994,N_16817,N_16467);
nor U24995 (N_24995,N_15412,N_17252);
nand U24996 (N_24996,N_16157,N_16292);
nor U24997 (N_24997,N_16615,N_19787);
and U24998 (N_24998,N_16193,N_19052);
nand U24999 (N_24999,N_17071,N_16536);
nand UO_0 (O_0,N_23029,N_22976);
nand UO_1 (O_1,N_20135,N_23910);
xor UO_2 (O_2,N_24498,N_20098);
xor UO_3 (O_3,N_22914,N_21391);
and UO_4 (O_4,N_24573,N_22385);
nand UO_5 (O_5,N_21999,N_23975);
or UO_6 (O_6,N_20353,N_21998);
nor UO_7 (O_7,N_24627,N_23843);
and UO_8 (O_8,N_21670,N_24342);
and UO_9 (O_9,N_21582,N_22598);
and UO_10 (O_10,N_21790,N_24440);
or UO_11 (O_11,N_23328,N_21749);
xor UO_12 (O_12,N_22613,N_24412);
and UO_13 (O_13,N_23579,N_20171);
and UO_14 (O_14,N_21569,N_21930);
and UO_15 (O_15,N_20830,N_20928);
and UO_16 (O_16,N_21285,N_21466);
nand UO_17 (O_17,N_23243,N_20515);
nor UO_18 (O_18,N_22559,N_23139);
and UO_19 (O_19,N_22384,N_20723);
nor UO_20 (O_20,N_20937,N_22907);
nor UO_21 (O_21,N_24591,N_20368);
nor UO_22 (O_22,N_23747,N_20963);
nor UO_23 (O_23,N_22859,N_23428);
and UO_24 (O_24,N_20616,N_20557);
and UO_25 (O_25,N_21113,N_21169);
or UO_26 (O_26,N_24650,N_23124);
nor UO_27 (O_27,N_23069,N_21452);
nor UO_28 (O_28,N_23636,N_20671);
nor UO_29 (O_29,N_20980,N_22338);
nand UO_30 (O_30,N_24017,N_22948);
and UO_31 (O_31,N_22390,N_22647);
or UO_32 (O_32,N_21610,N_22840);
nand UO_33 (O_33,N_24348,N_22224);
xor UO_34 (O_34,N_24629,N_20144);
or UO_35 (O_35,N_23160,N_24835);
or UO_36 (O_36,N_24187,N_23797);
and UO_37 (O_37,N_23840,N_22349);
or UO_38 (O_38,N_20177,N_20179);
or UO_39 (O_39,N_24942,N_20925);
or UO_40 (O_40,N_20014,N_21762);
and UO_41 (O_41,N_24202,N_23759);
nor UO_42 (O_42,N_23202,N_21655);
nand UO_43 (O_43,N_24507,N_23021);
or UO_44 (O_44,N_20800,N_20683);
nor UO_45 (O_45,N_24170,N_20173);
or UO_46 (O_46,N_21812,N_22792);
and UO_47 (O_47,N_22370,N_21995);
or UO_48 (O_48,N_21882,N_24387);
nor UO_49 (O_49,N_23896,N_24977);
xor UO_50 (O_50,N_24588,N_21904);
nor UO_51 (O_51,N_24418,N_23960);
nor UO_52 (O_52,N_20011,N_22697);
nand UO_53 (O_53,N_22211,N_22794);
or UO_54 (O_54,N_23944,N_20664);
nor UO_55 (O_55,N_20362,N_23716);
nand UO_56 (O_56,N_23077,N_24075);
nand UO_57 (O_57,N_23489,N_22098);
nand UO_58 (O_58,N_21606,N_21756);
or UO_59 (O_59,N_21835,N_22767);
nor UO_60 (O_60,N_22626,N_20570);
or UO_61 (O_61,N_23079,N_21000);
nand UO_62 (O_62,N_24105,N_20359);
and UO_63 (O_63,N_22120,N_24385);
or UO_64 (O_64,N_20523,N_21873);
or UO_65 (O_65,N_24667,N_23694);
nand UO_66 (O_66,N_23658,N_21676);
nor UO_67 (O_67,N_21679,N_20086);
nor UO_68 (O_68,N_21609,N_24386);
and UO_69 (O_69,N_21155,N_23946);
and UO_70 (O_70,N_20453,N_23325);
or UO_71 (O_71,N_23281,N_21320);
nor UO_72 (O_72,N_21289,N_23048);
nand UO_73 (O_73,N_24201,N_24943);
or UO_74 (O_74,N_23121,N_23780);
xor UO_75 (O_75,N_20155,N_22869);
nor UO_76 (O_76,N_22268,N_20957);
nor UO_77 (O_77,N_23955,N_22898);
or UO_78 (O_78,N_21953,N_23935);
nand UO_79 (O_79,N_20078,N_22660);
nand UO_80 (O_80,N_20236,N_22395);
and UO_81 (O_81,N_23627,N_23958);
nand UO_82 (O_82,N_24619,N_21312);
or UO_83 (O_83,N_21051,N_20278);
nor UO_84 (O_84,N_21920,N_20959);
or UO_85 (O_85,N_22029,N_20667);
nand UO_86 (O_86,N_20705,N_20844);
or UO_87 (O_87,N_24554,N_20713);
nor UO_88 (O_88,N_23692,N_20355);
nor UO_89 (O_89,N_21740,N_23287);
nand UO_90 (O_90,N_20599,N_20894);
xor UO_91 (O_91,N_20228,N_20465);
or UO_92 (O_92,N_22352,N_23407);
nand UO_93 (O_93,N_22426,N_23740);
or UO_94 (O_94,N_20710,N_23259);
and UO_95 (O_95,N_23689,N_22278);
xor UO_96 (O_96,N_22151,N_21378);
nor UO_97 (O_97,N_20906,N_20855);
and UO_98 (O_98,N_21933,N_23280);
and UO_99 (O_99,N_22146,N_24431);
and UO_100 (O_100,N_22518,N_23999);
or UO_101 (O_101,N_23963,N_24042);
nor UO_102 (O_102,N_23597,N_23679);
nand UO_103 (O_103,N_22602,N_21187);
nor UO_104 (O_104,N_21591,N_24182);
or UO_105 (O_105,N_23702,N_20121);
or UO_106 (O_106,N_21978,N_20506);
or UO_107 (O_107,N_24450,N_20137);
nand UO_108 (O_108,N_21695,N_21766);
and UO_109 (O_109,N_20986,N_20912);
and UO_110 (O_110,N_20130,N_24612);
nor UO_111 (O_111,N_24155,N_23872);
and UO_112 (O_112,N_24358,N_24363);
or UO_113 (O_113,N_20150,N_23777);
or UO_114 (O_114,N_20672,N_22520);
nor UO_115 (O_115,N_20929,N_23286);
nand UO_116 (O_116,N_20433,N_21152);
or UO_117 (O_117,N_20482,N_24928);
and UO_118 (O_118,N_24141,N_21970);
nand UO_119 (O_119,N_23097,N_23841);
and UO_120 (O_120,N_23932,N_24026);
nor UO_121 (O_121,N_20068,N_22297);
xor UO_122 (O_122,N_24258,N_24484);
nor UO_123 (O_123,N_24491,N_22679);
nand UO_124 (O_124,N_24955,N_20307);
and UO_125 (O_125,N_21417,N_23918);
or UO_126 (O_126,N_21759,N_23903);
nand UO_127 (O_127,N_24396,N_24020);
and UO_128 (O_128,N_20352,N_23371);
and UO_129 (O_129,N_24854,N_22072);
and UO_130 (O_130,N_24508,N_20378);
and UO_131 (O_131,N_22593,N_22881);
nor UO_132 (O_132,N_20062,N_20954);
and UO_133 (O_133,N_22551,N_20138);
and UO_134 (O_134,N_22889,N_23421);
and UO_135 (O_135,N_24559,N_22011);
nand UO_136 (O_136,N_21375,N_23793);
and UO_137 (O_137,N_21821,N_24641);
nor UO_138 (O_138,N_22190,N_24297);
nand UO_139 (O_139,N_20707,N_22777);
xor UO_140 (O_140,N_21434,N_21036);
or UO_141 (O_141,N_23762,N_21634);
or UO_142 (O_142,N_20084,N_21657);
nor UO_143 (O_143,N_22635,N_20376);
and UO_144 (O_144,N_24748,N_22568);
nand UO_145 (O_145,N_23902,N_24433);
xnor UO_146 (O_146,N_23183,N_22300);
nand UO_147 (O_147,N_24133,N_24785);
xnor UO_148 (O_148,N_23835,N_20493);
or UO_149 (O_149,N_22282,N_21771);
nand UO_150 (O_150,N_23188,N_23576);
and UO_151 (O_151,N_22644,N_23363);
or UO_152 (O_152,N_23945,N_24540);
or UO_153 (O_153,N_22921,N_20250);
or UO_154 (O_154,N_22958,N_23900);
or UO_155 (O_155,N_23413,N_22639);
nand UO_156 (O_156,N_20087,N_23058);
xor UO_157 (O_157,N_21031,N_20814);
nor UO_158 (O_158,N_21271,N_20106);
or UO_159 (O_159,N_24286,N_22342);
and UO_160 (O_160,N_23211,N_23155);
nand UO_161 (O_161,N_23892,N_21996);
nor UO_162 (O_162,N_20642,N_23558);
and UO_163 (O_163,N_22149,N_21424);
nand UO_164 (O_164,N_21418,N_23603);
and UO_165 (O_165,N_24095,N_22612);
nand UO_166 (O_166,N_22439,N_23172);
and UO_167 (O_167,N_23770,N_21564);
or UO_168 (O_168,N_24671,N_20140);
or UO_169 (O_169,N_20417,N_21142);
nor UO_170 (O_170,N_23100,N_20881);
or UO_171 (O_171,N_20456,N_22562);
or UO_172 (O_172,N_23909,N_24516);
or UO_173 (O_173,N_23232,N_22037);
xor UO_174 (O_174,N_22633,N_24195);
or UO_175 (O_175,N_20735,N_22734);
nand UO_176 (O_176,N_20818,N_23296);
nor UO_177 (O_177,N_23837,N_21573);
nand UO_178 (O_178,N_22521,N_20819);
or UO_179 (O_179,N_21209,N_23541);
nor UO_180 (O_180,N_24562,N_21469);
xor UO_181 (O_181,N_24359,N_21863);
and UO_182 (O_182,N_22817,N_22448);
or UO_183 (O_183,N_20991,N_21060);
and UO_184 (O_184,N_24390,N_22141);
and UO_185 (O_185,N_20466,N_20627);
and UO_186 (O_186,N_23465,N_24626);
nor UO_187 (O_187,N_23344,N_23847);
or UO_188 (O_188,N_24850,N_24913);
or UO_189 (O_189,N_24154,N_21077);
and UO_190 (O_190,N_24683,N_24765);
nor UO_191 (O_191,N_24309,N_20467);
or UO_192 (O_192,N_20170,N_24566);
and UO_193 (O_193,N_24300,N_21718);
or UO_194 (O_194,N_21621,N_24244);
and UO_195 (O_195,N_20758,N_21221);
and UO_196 (O_196,N_24113,N_22990);
nand UO_197 (O_197,N_21144,N_23640);
nor UO_198 (O_198,N_20793,N_22417);
and UO_199 (O_199,N_23518,N_21767);
or UO_200 (O_200,N_23581,N_20679);
and UO_201 (O_201,N_24163,N_20286);
and UO_202 (O_202,N_20785,N_22970);
nor UO_203 (O_203,N_24362,N_22173);
nand UO_204 (O_204,N_23306,N_22706);
and UO_205 (O_205,N_23175,N_21688);
nor UO_206 (O_206,N_22293,N_20879);
nor UO_207 (O_207,N_21846,N_24570);
nand UO_208 (O_208,N_23967,N_20113);
or UO_209 (O_209,N_24245,N_24282);
and UO_210 (O_210,N_20588,N_22761);
nand UO_211 (O_211,N_20477,N_23655);
and UO_212 (O_212,N_21611,N_22319);
xor UO_213 (O_213,N_21504,N_23814);
nand UO_214 (O_214,N_22851,N_20348);
and UO_215 (O_215,N_23113,N_20509);
or UO_216 (O_216,N_23893,N_22466);
or UO_217 (O_217,N_24538,N_21415);
nand UO_218 (O_218,N_23527,N_22205);
nor UO_219 (O_219,N_20973,N_20988);
or UO_220 (O_220,N_22858,N_23057);
nor UO_221 (O_221,N_22063,N_20408);
and UO_222 (O_222,N_21181,N_24689);
and UO_223 (O_223,N_22802,N_23867);
xor UO_224 (O_224,N_23018,N_20784);
nand UO_225 (O_225,N_23566,N_24274);
or UO_226 (O_226,N_20851,N_20909);
or UO_227 (O_227,N_23123,N_22493);
and UO_228 (O_228,N_22513,N_20478);
nand UO_229 (O_229,N_21758,N_21108);
nand UO_230 (O_230,N_21720,N_22453);
xnor UO_231 (O_231,N_24224,N_24164);
and UO_232 (O_232,N_21824,N_24401);
nand UO_233 (O_233,N_21241,N_21827);
nand UO_234 (O_234,N_23300,N_22930);
or UO_235 (O_235,N_21689,N_20694);
and UO_236 (O_236,N_23792,N_20418);
and UO_237 (O_237,N_24524,N_24298);
nand UO_238 (O_238,N_23844,N_23961);
and UO_239 (O_239,N_20184,N_23794);
nor UO_240 (O_240,N_24514,N_20834);
and UO_241 (O_241,N_23972,N_21991);
nand UO_242 (O_242,N_20951,N_20497);
nand UO_243 (O_243,N_22780,N_20526);
nor UO_244 (O_244,N_21521,N_21095);
or UO_245 (O_245,N_24991,N_21176);
xnor UO_246 (O_246,N_21130,N_22507);
nor UO_247 (O_247,N_22285,N_24241);
or UO_248 (O_248,N_23115,N_20805);
xor UO_249 (O_249,N_24435,N_22910);
nand UO_250 (O_250,N_23378,N_24515);
nand UO_251 (O_251,N_24166,N_22575);
or UO_252 (O_252,N_20858,N_23870);
and UO_253 (O_253,N_23218,N_23998);
and UO_254 (O_254,N_23703,N_20282);
nand UO_255 (O_255,N_20558,N_21367);
and UO_256 (O_256,N_22431,N_22523);
and UO_257 (O_257,N_22042,N_21788);
and UO_258 (O_258,N_23912,N_21772);
nor UO_259 (O_259,N_22228,N_24144);
nand UO_260 (O_260,N_21588,N_22103);
nand UO_261 (O_261,N_20652,N_24509);
and UO_262 (O_262,N_24242,N_21224);
and UO_263 (O_263,N_23699,N_22893);
nand UO_264 (O_264,N_24628,N_20208);
nor UO_265 (O_265,N_22045,N_23509);
or UO_266 (O_266,N_21931,N_20993);
nor UO_267 (O_267,N_21279,N_20468);
nand UO_268 (O_268,N_21994,N_23379);
nor UO_269 (O_269,N_21120,N_23979);
nor UO_270 (O_270,N_23153,N_23082);
nand UO_271 (O_271,N_24833,N_24319);
or UO_272 (O_272,N_22630,N_20065);
nor UO_273 (O_273,N_21165,N_20345);
xnor UO_274 (O_274,N_24609,N_23686);
and UO_275 (O_275,N_22100,N_21966);
xor UO_276 (O_276,N_21467,N_24829);
or UO_277 (O_277,N_24781,N_22737);
nand UO_278 (O_278,N_24879,N_22218);
nor UO_279 (O_279,N_24256,N_23411);
xor UO_280 (O_280,N_24279,N_23244);
and UO_281 (O_281,N_21149,N_24295);
xor UO_282 (O_282,N_21058,N_20235);
nor UO_283 (O_283,N_22789,N_20393);
nand UO_284 (O_284,N_22161,N_20238);
nand UO_285 (O_285,N_24198,N_21032);
nor UO_286 (O_286,N_24158,N_24060);
or UO_287 (O_287,N_20053,N_23587);
nor UO_288 (O_288,N_22185,N_20054);
or UO_289 (O_289,N_23158,N_24531);
nor UO_290 (O_290,N_21944,N_24010);
and UO_291 (O_291,N_21210,N_23663);
or UO_292 (O_292,N_21349,N_21485);
nand UO_293 (O_293,N_23273,N_20296);
or UO_294 (O_294,N_20488,N_22208);
nor UO_295 (O_295,N_24473,N_21708);
nand UO_296 (O_296,N_23223,N_21770);
or UO_297 (O_297,N_24252,N_22331);
and UO_298 (O_298,N_23733,N_22363);
nand UO_299 (O_299,N_21997,N_21600);
nand UO_300 (O_300,N_22927,N_20441);
nor UO_301 (O_301,N_24079,N_20504);
nand UO_302 (O_302,N_24383,N_21881);
nand UO_303 (O_303,N_20522,N_24221);
xnor UO_304 (O_304,N_24581,N_21910);
and UO_305 (O_305,N_21735,N_23106);
nand UO_306 (O_306,N_20079,N_21653);
nor UO_307 (O_307,N_22492,N_24409);
and UO_308 (O_308,N_24129,N_20483);
nor UO_309 (O_309,N_22487,N_24486);
or UO_310 (O_310,N_20984,N_22603);
nor UO_311 (O_311,N_21022,N_20326);
and UO_312 (O_312,N_24556,N_23024);
and UO_313 (O_313,N_23933,N_20055);
nand UO_314 (O_314,N_23570,N_21494);
or UO_315 (O_315,N_24594,N_20254);
or UO_316 (O_316,N_20443,N_20424);
nor UO_317 (O_317,N_22839,N_21705);
nand UO_318 (O_318,N_24771,N_23250);
xnor UO_319 (O_319,N_24937,N_20043);
and UO_320 (O_320,N_21184,N_24495);
nor UO_321 (O_321,N_24679,N_22692);
nor UO_322 (O_322,N_23451,N_24767);
or UO_323 (O_323,N_24981,N_20853);
nor UO_324 (O_324,N_23006,N_22757);
and UO_325 (O_325,N_20941,N_23612);
nor UO_326 (O_326,N_23865,N_21331);
nand UO_327 (O_327,N_22280,N_21448);
xor UO_328 (O_328,N_23196,N_20439);
nand UO_329 (O_329,N_21015,N_23238);
nand UO_330 (O_330,N_24862,N_20840);
nand UO_331 (O_331,N_24188,N_23226);
xnor UO_332 (O_332,N_23105,N_23341);
nand UO_333 (O_333,N_22303,N_22801);
nor UO_334 (O_334,N_22102,N_21902);
nand UO_335 (O_335,N_22750,N_24194);
nor UO_336 (O_336,N_23394,N_22629);
nor UO_337 (O_337,N_23635,N_21477);
nand UO_338 (O_338,N_24798,N_22867);
xnor UO_339 (O_339,N_22194,N_23824);
nand UO_340 (O_340,N_22200,N_23441);
nand UO_341 (O_341,N_22749,N_20803);
and UO_342 (O_342,N_20197,N_23142);
and UO_343 (O_343,N_24983,N_23810);
nand UO_344 (O_344,N_20035,N_23878);
nand UO_345 (O_345,N_23071,N_23681);
and UO_346 (O_346,N_21760,N_23129);
nand UO_347 (O_347,N_21337,N_21177);
or UO_348 (O_348,N_21536,N_21831);
and UO_349 (O_349,N_21733,N_23497);
nand UO_350 (O_350,N_24614,N_22250);
or UO_351 (O_351,N_20530,N_23205);
nand UO_352 (O_352,N_24296,N_20028);
and UO_353 (O_353,N_22708,N_21739);
or UO_354 (O_354,N_23102,N_24485);
or UO_355 (O_355,N_24369,N_20081);
xor UO_356 (O_356,N_24929,N_24326);
or UO_357 (O_357,N_21212,N_22275);
nand UO_358 (O_358,N_23633,N_20152);
nor UO_359 (O_359,N_21444,N_20330);
nand UO_360 (O_360,N_24522,N_22118);
or UO_361 (O_361,N_24809,N_23853);
nor UO_362 (O_362,N_22152,N_22261);
xor UO_363 (O_363,N_24544,N_20400);
nor UO_364 (O_364,N_22314,N_23424);
nand UO_365 (O_365,N_22525,N_24014);
xor UO_366 (O_366,N_23305,N_22649);
nor UO_367 (O_367,N_22371,N_20195);
xnor UO_368 (O_368,N_21493,N_21123);
or UO_369 (O_369,N_23073,N_20227);
and UO_370 (O_370,N_20132,N_24230);
or UO_371 (O_371,N_22561,N_23003);
and UO_372 (O_372,N_24247,N_24743);
or UO_373 (O_373,N_24189,N_22712);
nand UO_374 (O_374,N_23751,N_21354);
or UO_375 (O_375,N_22873,N_24052);
or UO_376 (O_376,N_21304,N_23440);
xnor UO_377 (O_377,N_23191,N_21935);
nand UO_378 (O_378,N_20560,N_20787);
or UO_379 (O_379,N_24846,N_20310);
nand UO_380 (O_380,N_21268,N_22396);
and UO_381 (O_381,N_21731,N_21549);
and UO_382 (O_382,N_21678,N_24535);
or UO_383 (O_383,N_20585,N_24847);
and UO_384 (O_384,N_20974,N_23680);
nor UO_385 (O_385,N_20444,N_22591);
and UO_386 (O_386,N_20036,N_22748);
and UO_387 (O_387,N_21801,N_23236);
nor UO_388 (O_388,N_22140,N_20625);
nand UO_389 (O_389,N_21666,N_20623);
nor UO_390 (O_390,N_20968,N_21604);
nand UO_391 (O_391,N_21537,N_21915);
or UO_392 (O_392,N_21937,N_22989);
xor UO_393 (O_393,N_21748,N_20938);
or UO_394 (O_394,N_21656,N_21692);
nor UO_395 (O_395,N_21507,N_22271);
nor UO_396 (O_396,N_23430,N_22286);
nor UO_397 (O_397,N_20712,N_23829);
nand UO_398 (O_398,N_21002,N_20145);
nand UO_399 (O_399,N_23199,N_23053);
or UO_400 (O_400,N_22425,N_21357);
nand UO_401 (O_401,N_21359,N_24789);
nand UO_402 (O_402,N_20711,N_22435);
nand UO_403 (O_403,N_22341,N_22061);
nand UO_404 (O_404,N_21746,N_23608);
or UO_405 (O_405,N_21328,N_21200);
nor UO_406 (O_406,N_22198,N_21018);
xor UO_407 (O_407,N_22189,N_20581);
and UO_408 (O_408,N_24137,N_20017);
or UO_409 (O_409,N_24962,N_23538);
nand UO_410 (O_410,N_20041,N_20922);
and UO_411 (O_411,N_20426,N_20921);
or UO_412 (O_412,N_22415,N_24877);
or UO_413 (O_413,N_20458,N_24897);
xor UO_414 (O_414,N_22419,N_24775);
and UO_415 (O_415,N_22924,N_23542);
and UO_416 (O_416,N_22961,N_23161);
or UO_417 (O_417,N_22862,N_22822);
nand UO_418 (O_418,N_20440,N_24225);
and UO_419 (O_419,N_20841,N_22330);
nor UO_420 (O_420,N_21829,N_22281);
and UO_421 (O_421,N_20660,N_23856);
xnor UO_422 (O_422,N_22292,N_21353);
and UO_423 (O_423,N_23406,N_23215);
nor UO_424 (O_424,N_20969,N_21932);
or UO_425 (O_425,N_20726,N_22219);
nor UO_426 (O_426,N_22014,N_21426);
and UO_427 (O_427,N_20918,N_20047);
or UO_428 (O_428,N_22409,N_22707);
or UO_429 (O_429,N_23613,N_20645);
nor UO_430 (O_430,N_20252,N_21061);
nand UO_431 (O_431,N_24265,N_24994);
or UO_432 (O_432,N_20559,N_22516);
xor UO_433 (O_433,N_20284,N_23045);
and UO_434 (O_434,N_23643,N_20165);
nor UO_435 (O_435,N_23786,N_23745);
nand UO_436 (O_436,N_20018,N_20429);
nand UO_437 (O_437,N_21358,N_24766);
nor UO_438 (O_438,N_22508,N_23255);
or UO_439 (O_439,N_24982,N_23688);
nor UO_440 (O_440,N_23864,N_23649);
nand UO_441 (O_441,N_20024,N_21722);
and UO_442 (O_442,N_23673,N_21104);
and UO_443 (O_443,N_22947,N_20976);
and UO_444 (O_444,N_22312,N_24382);
and UO_445 (O_445,N_21332,N_21986);
and UO_446 (O_446,N_21050,N_22437);
nand UO_447 (O_447,N_20731,N_24577);
nor UO_448 (O_448,N_22870,N_20886);
nand UO_449 (O_449,N_23746,N_20129);
nor UO_450 (O_450,N_22548,N_23295);
nand UO_451 (O_451,N_21121,N_24161);
nand UO_452 (O_452,N_21511,N_20823);
nand UO_453 (O_453,N_20962,N_24726);
nand UO_454 (O_454,N_20849,N_23025);
and UO_455 (O_455,N_21094,N_22528);
nor UO_456 (O_456,N_23517,N_21816);
or UO_457 (O_457,N_22830,N_21398);
nand UO_458 (O_458,N_22696,N_23198);
nor UO_459 (O_459,N_22248,N_22857);
nor UO_460 (O_460,N_22442,N_22532);
nor UO_461 (O_461,N_22236,N_23177);
nor UO_462 (O_462,N_20692,N_21076);
nor UO_463 (O_463,N_20510,N_23513);
or UO_464 (O_464,N_21581,N_21680);
and UO_465 (O_465,N_20438,N_20745);
nor UO_466 (O_466,N_23730,N_21065);
and UO_467 (O_467,N_21566,N_24532);
and UO_468 (O_468,N_23785,N_21178);
or UO_469 (O_469,N_24529,N_22450);
nand UO_470 (O_470,N_24536,N_24739);
or UO_471 (O_471,N_24036,N_21458);
and UO_472 (O_472,N_23988,N_21616);
nand UO_473 (O_473,N_23811,N_22413);
and UO_474 (O_474,N_24223,N_24366);
nor UO_475 (O_475,N_21750,N_20060);
nand UO_476 (O_476,N_20702,N_20397);
or UO_477 (O_477,N_22535,N_23044);
nor UO_478 (O_478,N_24177,N_21470);
and UO_479 (O_479,N_23365,N_21183);
and UO_480 (O_480,N_23194,N_24682);
xor UO_481 (O_481,N_23744,N_20409);
nand UO_482 (O_482,N_21729,N_21895);
nand UO_483 (O_483,N_22628,N_24449);
and UO_484 (O_484,N_21161,N_24453);
or UO_485 (O_485,N_22824,N_23264);
nor UO_486 (O_486,N_23766,N_21407);
and UO_487 (O_487,N_21526,N_21732);
and UO_488 (O_488,N_23398,N_24590);
nor UO_489 (O_489,N_22109,N_23302);
nand UO_490 (O_490,N_24857,N_22595);
nand UO_491 (O_491,N_24299,N_20865);
and UO_492 (O_492,N_24493,N_22445);
or UO_493 (O_493,N_20746,N_23422);
nand UO_494 (O_494,N_20031,N_22375);
nor UO_495 (O_495,N_22847,N_22049);
nor UO_496 (O_496,N_23995,N_20704);
nor UO_497 (O_497,N_24002,N_24009);
nand UO_498 (O_498,N_24192,N_23446);
or UO_499 (O_499,N_20390,N_20529);
nor UO_500 (O_500,N_22615,N_21699);
and UO_501 (O_501,N_24321,N_22793);
nand UO_502 (O_502,N_20817,N_23146);
and UO_503 (O_503,N_24839,N_24914);
nand UO_504 (O_504,N_22852,N_24061);
or UO_505 (O_505,N_23741,N_22322);
nand UO_506 (O_506,N_24757,N_21909);
nor UO_507 (O_507,N_22046,N_21383);
and UO_508 (O_508,N_23089,N_23239);
nor UO_509 (O_509,N_20049,N_24584);
nor UO_510 (O_510,N_20975,N_20926);
xnor UO_511 (O_511,N_24721,N_20224);
and UO_512 (O_512,N_21495,N_23532);
nor UO_513 (O_513,N_22308,N_21940);
and UO_514 (O_514,N_20846,N_22624);
or UO_515 (O_515,N_20248,N_23732);
nand UO_516 (O_516,N_23469,N_21186);
and UO_517 (O_517,N_20421,N_22685);
nor UO_518 (O_518,N_22768,N_23775);
xor UO_519 (O_519,N_24527,N_22320);
and UO_520 (O_520,N_20946,N_24618);
nand UO_521 (O_521,N_23370,N_22007);
nor UO_522 (O_522,N_20042,N_20386);
nand UO_523 (O_523,N_22157,N_24264);
and UO_524 (O_524,N_20162,N_21292);
nor UO_525 (O_525,N_23789,N_20255);
nand UO_526 (O_526,N_21780,N_21921);
or UO_527 (O_527,N_21419,N_20654);
or UO_528 (O_528,N_23323,N_24510);
and UO_529 (O_529,N_20548,N_20044);
nand UO_530 (O_530,N_23374,N_23393);
or UO_531 (O_531,N_22254,N_24080);
and UO_532 (O_532,N_22294,N_24381);
xor UO_533 (O_533,N_24350,N_22485);
xnor UO_534 (O_534,N_21518,N_20476);
and UO_535 (O_535,N_22981,N_23156);
xor UO_536 (O_536,N_20773,N_24499);
nor UO_537 (O_537,N_22469,N_24634);
xnor UO_538 (O_538,N_20251,N_23752);
nor UO_539 (O_539,N_24374,N_24179);
or UO_540 (O_540,N_21968,N_24888);
and UO_541 (O_541,N_21217,N_20939);
nand UO_542 (O_542,N_22489,N_23334);
xnor UO_543 (O_543,N_22549,N_24446);
nor UO_544 (O_544,N_24324,N_24400);
nor UO_545 (O_545,N_20073,N_23180);
and UO_546 (O_546,N_24772,N_23645);
nand UO_547 (O_547,N_22746,N_23200);
and UO_548 (O_548,N_21249,N_20459);
nor UO_549 (O_549,N_24056,N_21936);
nand UO_550 (O_550,N_23476,N_20958);
or UO_551 (O_551,N_20786,N_23482);
and UO_552 (O_552,N_24000,N_21815);
nand UO_553 (O_553,N_21726,N_23041);
xnor UO_554 (O_554,N_21885,N_22166);
or UO_555 (O_555,N_20315,N_23099);
nor UO_556 (O_556,N_21845,N_23863);
nand UO_557 (O_557,N_23167,N_20513);
or UO_558 (O_558,N_22664,N_22674);
nor UO_559 (O_559,N_24368,N_23190);
nand UO_560 (O_560,N_21590,N_22356);
or UO_561 (O_561,N_20464,N_22229);
nand UO_562 (O_562,N_23671,N_20914);
nor UO_563 (O_563,N_20337,N_24999);
nand UO_564 (O_564,N_24470,N_20026);
and UO_565 (O_565,N_23711,N_24367);
xor UO_566 (O_566,N_23969,N_20677);
or UO_567 (O_567,N_20586,N_21035);
or UO_568 (O_568,N_24807,N_20835);
and UO_569 (O_569,N_23085,N_24249);
nand UO_570 (O_570,N_24394,N_23005);
nand UO_571 (O_571,N_20537,N_24153);
or UO_572 (O_572,N_20948,N_20943);
or UO_573 (O_573,N_20617,N_24727);
and UO_574 (O_574,N_22329,N_24959);
nor UO_575 (O_575,N_22259,N_23297);
nor UO_576 (O_576,N_21284,N_23135);
or UO_577 (O_577,N_24115,N_23715);
nor UO_578 (O_578,N_21214,N_24558);
and UO_579 (O_579,N_20698,N_21266);
and UO_580 (O_580,N_21302,N_20864);
or UO_581 (O_581,N_21871,N_24370);
xor UO_582 (O_582,N_22298,N_23667);
or UO_583 (O_583,N_21420,N_23605);
xor UO_584 (O_584,N_20927,N_23956);
or UO_585 (O_585,N_21884,N_20681);
nand UO_586 (O_586,N_22751,N_23298);
or UO_587 (O_587,N_23050,N_24403);
and UO_588 (O_588,N_22172,N_24415);
or UO_589 (O_589,N_21747,N_20333);
nand UO_590 (O_590,N_21006,N_23882);
nand UO_591 (O_591,N_21532,N_20720);
or UO_592 (O_592,N_22875,N_22723);
nand UO_593 (O_593,N_24148,N_20994);
nand UO_594 (O_594,N_22482,N_23049);
xnor UO_595 (O_595,N_20552,N_22998);
or UO_596 (O_596,N_24866,N_22705);
nor UO_597 (O_597,N_23083,N_23973);
xnor UO_598 (O_598,N_23753,N_21842);
or UO_599 (O_599,N_24266,N_20647);
nor UO_600 (O_600,N_23019,N_21451);
nand UO_601 (O_601,N_21361,N_24672);
and UO_602 (O_602,N_23127,N_20420);
xnor UO_603 (O_603,N_21742,N_21390);
nand UO_604 (O_604,N_21201,N_20160);
and UO_605 (O_605,N_23550,N_23385);
nand UO_606 (O_606,N_21833,N_20604);
nor UO_607 (O_607,N_20085,N_22527);
nor UO_608 (O_608,N_24452,N_23914);
or UO_609 (O_609,N_21593,N_23065);
nor UO_610 (O_610,N_23657,N_20191);
nor UO_611 (O_611,N_23262,N_24697);
or UO_612 (O_612,N_24948,N_24867);
and UO_613 (O_613,N_20214,N_22018);
and UO_614 (O_614,N_23543,N_21502);
xnor UO_615 (O_615,N_20633,N_21291);
nand UO_616 (O_616,N_20202,N_20675);
or UO_617 (O_617,N_22931,N_23372);
nor UO_618 (O_618,N_23248,N_24891);
nand UO_619 (O_619,N_20892,N_23676);
or UO_620 (O_620,N_20734,N_21719);
nor UO_621 (O_621,N_21457,N_23496);
nor UO_622 (O_622,N_24734,N_24474);
nor UO_623 (O_623,N_21132,N_22094);
or UO_624 (O_624,N_24797,N_21531);
nand UO_625 (O_625,N_22803,N_22452);
xor UO_626 (O_626,N_22318,N_23981);
or UO_627 (O_627,N_24422,N_21851);
and UO_628 (O_628,N_22531,N_24869);
nand UO_629 (O_629,N_21492,N_20167);
or UO_630 (O_630,N_24755,N_23908);
nand UO_631 (O_631,N_20212,N_24477);
nor UO_632 (O_632,N_23881,N_22288);
and UO_633 (O_633,N_21213,N_24746);
and UO_634 (O_634,N_23529,N_22906);
nand UO_635 (O_635,N_24965,N_24373);
or UO_636 (O_636,N_21207,N_20690);
nor UO_637 (O_637,N_22481,N_20001);
xnor UO_638 (O_638,N_24630,N_20192);
nand UO_639 (O_639,N_24238,N_21482);
xor UO_640 (O_640,N_20587,N_22034);
and UO_641 (O_641,N_23116,N_20809);
or UO_642 (O_642,N_20484,N_22441);
nand UO_643 (O_643,N_24813,N_20843);
or UO_644 (O_644,N_21175,N_24892);
and UO_645 (O_645,N_20635,N_21222);
or UO_646 (O_646,N_20541,N_21117);
and UO_647 (O_647,N_21473,N_22992);
xor UO_648 (O_648,N_23884,N_20995);
or UO_649 (O_649,N_24045,N_24131);
or UO_650 (O_650,N_24699,N_23072);
or UO_651 (O_651,N_21027,N_22719);
nand UO_652 (O_652,N_20543,N_22972);
xnor UO_653 (O_653,N_20431,N_23926);
and UO_654 (O_654,N_22740,N_20945);
or UO_655 (O_655,N_23293,N_22742);
nor UO_656 (O_656,N_22617,N_22731);
and UO_657 (O_657,N_23015,N_20154);
and UO_658 (O_658,N_22062,N_24178);
nor UO_659 (O_659,N_24763,N_24533);
and UO_660 (O_660,N_21674,N_24651);
nor UO_661 (O_661,N_21955,N_24901);
nand UO_662 (O_662,N_22587,N_23567);
or UO_663 (O_663,N_21189,N_21057);
or UO_664 (O_664,N_20309,N_24126);
nand UO_665 (O_665,N_24711,N_22067);
and UO_666 (O_666,N_20760,N_22025);
or UO_667 (O_667,N_24995,N_21350);
nand UO_668 (O_668,N_23522,N_23022);
or UO_669 (O_669,N_24024,N_20689);
or UO_670 (O_670,N_24622,N_23719);
nor UO_671 (O_671,N_23414,N_21298);
or UO_672 (O_672,N_22006,N_24545);
nand UO_673 (O_673,N_20934,N_23787);
nor UO_674 (O_674,N_23848,N_21408);
nor UO_675 (O_675,N_22714,N_22052);
xnor UO_676 (O_676,N_24206,N_21074);
nor UO_677 (O_677,N_22888,N_24130);
or UO_678 (O_678,N_22769,N_22913);
xor UO_679 (O_679,N_22519,N_21886);
xor UO_680 (O_680,N_22468,N_23357);
nor UO_681 (O_681,N_23631,N_20999);
xor UO_682 (O_682,N_23477,N_23825);
nand UO_683 (O_683,N_21776,N_22908);
and UO_684 (O_684,N_21414,N_20189);
nand UO_685 (O_685,N_21592,N_22348);
and UO_686 (O_686,N_20312,N_22252);
and UO_687 (O_687,N_23492,N_24621);
or UO_688 (O_688,N_20485,N_22831);
and UO_689 (O_689,N_20051,N_24871);
or UO_690 (O_690,N_23195,N_23707);
and UO_691 (O_691,N_22943,N_23551);
and UO_692 (O_692,N_24512,N_24259);
nand UO_693 (O_693,N_21980,N_22455);
nand UO_694 (O_694,N_24832,N_23754);
and UO_695 (O_695,N_24478,N_21409);
and UO_696 (O_696,N_21706,N_24044);
nor UO_697 (O_697,N_21958,N_21791);
xnor UO_698 (O_698,N_24722,N_21379);
nand UO_699 (O_699,N_20684,N_20546);
nand UO_700 (O_700,N_22882,N_24310);
nor UO_701 (O_701,N_20966,N_24873);
or UO_702 (O_702,N_24214,N_24361);
and UO_703 (O_703,N_22950,N_24117);
or UO_704 (O_704,N_23120,N_24693);
nor UO_705 (O_705,N_21675,N_23768);
nor UO_706 (O_706,N_20201,N_20606);
nor UO_707 (O_707,N_23526,N_24229);
or UO_708 (O_708,N_22317,N_24924);
and UO_709 (O_709,N_21257,N_22967);
and UO_710 (O_710,N_23845,N_23107);
or UO_711 (O_711,N_20933,N_21033);
nor UO_712 (O_712,N_21946,N_23891);
nor UO_713 (O_713,N_21805,N_21230);
nand UO_714 (O_714,N_21346,N_22573);
or UO_715 (O_715,N_24638,N_22806);
nand UO_716 (O_716,N_24142,N_21836);
or UO_717 (O_717,N_23828,N_22786);
nand UO_718 (O_718,N_20854,N_22267);
or UO_719 (O_719,N_24551,N_20792);
nor UO_720 (O_720,N_20607,N_24207);
nor UO_721 (O_721,N_22191,N_20637);
and UO_722 (O_722,N_23277,N_21404);
xor UO_723 (O_723,N_21270,N_20732);
xnor UO_724 (O_724,N_20204,N_20003);
or UO_725 (O_725,N_24673,N_24413);
nor UO_726 (O_726,N_22982,N_23193);
or UO_727 (O_727,N_24261,N_21671);
nand UO_728 (O_728,N_20520,N_24030);
nor UO_729 (O_729,N_20446,N_22702);
nor UO_730 (O_730,N_22753,N_22365);
or UO_731 (O_731,N_24909,N_24287);
and UO_732 (O_732,N_24425,N_24341);
nand UO_733 (O_733,N_22915,N_22262);
or UO_734 (O_734,N_21195,N_24330);
nor UO_735 (O_735,N_20046,N_21167);
and UO_736 (O_736,N_20622,N_21803);
and UO_737 (O_737,N_24458,N_21669);
or UO_738 (O_738,N_23136,N_20923);
and UO_739 (O_739,N_21309,N_24647);
nand UO_740 (O_740,N_22187,N_22412);
nand UO_741 (O_741,N_21055,N_23928);
nand UO_742 (O_742,N_21710,N_20940);
nand UO_743 (O_743,N_20534,N_23319);
and UO_744 (O_744,N_22808,N_22050);
nand UO_745 (O_745,N_23659,N_20334);
nor UO_746 (O_746,N_22775,N_21602);
or UO_747 (O_747,N_24941,N_24881);
or UO_748 (O_748,N_23122,N_21081);
or UO_749 (O_749,N_21314,N_24934);
nand UO_750 (O_750,N_20264,N_22903);
and UO_751 (O_751,N_23350,N_23096);
nor UO_752 (O_752,N_21193,N_24146);
nand UO_753 (O_753,N_23778,N_24648);
and UO_754 (O_754,N_23462,N_21240);
or UO_755 (O_755,N_22097,N_24407);
nand UO_756 (O_756,N_21598,N_21517);
or UO_757 (O_757,N_23266,N_21109);
or UO_758 (O_758,N_24741,N_21003);
and UO_759 (O_759,N_24354,N_20366);
and UO_760 (O_760,N_22904,N_21550);
and UO_761 (O_761,N_21244,N_21509);
or UO_762 (O_762,N_20952,N_22890);
and UO_763 (O_763,N_22678,N_24794);
and UO_764 (O_764,N_23980,N_24964);
and UO_765 (O_765,N_22952,N_22060);
nor UO_766 (O_766,N_21365,N_23487);
or UO_767 (O_767,N_24110,N_23448);
nand UO_768 (O_768,N_23861,N_21734);
nor UO_769 (O_769,N_20209,N_24517);
xor UO_770 (O_770,N_23304,N_21868);
nor UO_771 (O_771,N_20216,N_21806);
nand UO_772 (O_772,N_24884,N_24692);
or UO_773 (O_773,N_20992,N_21498);
nand UO_774 (O_774,N_22648,N_24625);
or UO_775 (O_775,N_23086,N_23359);
nor UO_776 (O_776,N_23993,N_22032);
or UO_777 (O_777,N_21927,N_21286);
or UO_778 (O_778,N_23506,N_23565);
or UO_779 (O_779,N_20399,N_21131);
or UO_780 (O_780,N_23162,N_21639);
nand UO_781 (O_781,N_22608,N_23763);
or UO_782 (O_782,N_24680,N_21376);
nor UO_783 (O_783,N_24889,N_23399);
nand UO_784 (O_784,N_22815,N_20148);
xor UO_785 (O_785,N_22563,N_20639);
xnor UO_786 (O_786,N_22572,N_23818);
and UO_787 (O_787,N_20826,N_22076);
and UO_788 (O_788,N_22766,N_22073);
or UO_789 (O_789,N_22695,N_20866);
and UO_790 (O_790,N_23820,N_20536);
or UO_791 (O_791,N_20402,N_21456);
nor UO_792 (O_792,N_20316,N_21410);
xor UO_793 (O_793,N_21837,N_21607);
or UO_794 (O_794,N_23391,N_21906);
xor UO_795 (O_795,N_23684,N_21103);
nor UO_796 (O_796,N_22885,N_22689);
nand UO_797 (O_797,N_20023,N_20776);
nand UO_798 (O_798,N_21701,N_22088);
or UO_799 (O_799,N_24702,N_24430);
xor UO_800 (O_800,N_23735,N_23478);
nor UO_801 (O_801,N_22225,N_21883);
or UO_802 (O_802,N_23375,N_24215);
xnor UO_803 (O_803,N_23367,N_22474);
nor UO_804 (O_804,N_23546,N_24378);
xor UO_805 (O_805,N_24885,N_20469);
nor UO_806 (O_806,N_24908,N_20470);
nor UO_807 (O_807,N_22814,N_20790);
or UO_808 (O_808,N_22717,N_23952);
xnor UO_809 (O_809,N_24560,N_22810);
or UO_810 (O_810,N_23545,N_20989);
nor UO_811 (O_811,N_21001,N_23216);
nor UO_812 (O_812,N_23665,N_21079);
or UO_813 (O_813,N_22323,N_22392);
nand UO_814 (O_814,N_23028,N_22180);
nor UO_815 (O_815,N_22763,N_22681);
nand UO_816 (O_816,N_22727,N_22538);
nor UO_817 (O_817,N_23227,N_24066);
xor UO_818 (O_818,N_22897,N_21574);
nor UO_819 (O_819,N_22821,N_24145);
nand UO_820 (O_820,N_24550,N_24204);
nand UO_821 (O_821,N_21192,N_20900);
xnor UO_822 (O_822,N_23382,N_23204);
and UO_823 (O_823,N_24865,N_23459);
nor UO_824 (O_824,N_24831,N_22115);
nand UO_825 (O_825,N_23092,N_24098);
or UO_826 (O_826,N_22502,N_23523);
nor UO_827 (O_827,N_22670,N_21311);
nand UO_828 (O_828,N_23410,N_23395);
nor UO_829 (O_829,N_22257,N_22979);
nand UO_830 (O_830,N_22788,N_23212);
or UO_831 (O_831,N_22953,N_24615);
or UO_832 (O_832,N_21009,N_21500);
and UO_833 (O_833,N_20317,N_22744);
nor UO_834 (O_834,N_23816,N_22984);
and UO_835 (O_835,N_21893,N_23376);
nand UO_836 (O_836,N_22816,N_22934);
nand UO_837 (O_837,N_22651,N_23147);
xor UO_838 (O_838,N_22328,N_24334);
and UO_839 (O_839,N_20859,N_21499);
and UO_840 (O_840,N_24073,N_24481);
or UO_841 (O_841,N_22028,N_20367);
nor UO_842 (O_842,N_20022,N_22020);
nand UO_843 (O_843,N_21580,N_22724);
and UO_844 (O_844,N_22597,N_20602);
nand UO_845 (O_845,N_24424,N_22940);
nor UO_846 (O_846,N_22845,N_20761);
nand UO_847 (O_847,N_21865,N_24159);
or UO_848 (O_848,N_22554,N_20299);
or UO_849 (O_849,N_22326,N_20763);
nand UO_850 (O_850,N_21070,N_22132);
xor UO_851 (O_851,N_20935,N_23493);
and UO_852 (O_852,N_20605,N_24031);
nor UO_853 (O_853,N_22854,N_24631);
and UO_854 (O_854,N_21465,N_22584);
or UO_855 (O_855,N_23027,N_23662);
or UO_856 (O_856,N_22069,N_23392);
nand UO_857 (O_857,N_23638,N_24349);
xor UO_858 (O_858,N_24805,N_24978);
and UO_859 (O_859,N_21557,N_20012);
and UO_860 (O_860,N_23321,N_23589);
or UO_861 (O_861,N_24759,N_22336);
xnor UO_862 (O_862,N_20432,N_21565);
or UO_863 (O_863,N_22008,N_21754);
nor UO_864 (O_864,N_21983,N_22960);
nor UO_865 (O_865,N_24479,N_20562);
nor UO_866 (O_866,N_20532,N_24108);
nand UO_867 (O_867,N_22515,N_20178);
and UO_868 (O_868,N_21368,N_21162);
and UO_869 (O_869,N_22099,N_22969);
and UO_870 (O_870,N_23207,N_24084);
or UO_871 (O_871,N_21533,N_20369);
nor UO_872 (O_872,N_20847,N_20103);
or UO_873 (O_873,N_24655,N_23809);
nand UO_874 (O_874,N_24096,N_21717);
or UO_875 (O_875,N_20153,N_20982);
and UO_876 (O_876,N_21133,N_21947);
nand UO_877 (O_877,N_21394,N_22249);
or UO_878 (O_878,N_21635,N_21231);
xor UO_879 (O_879,N_23203,N_20398);
and UO_880 (O_880,N_21101,N_21396);
nor UO_881 (O_881,N_22027,N_20442);
or UO_882 (O_882,N_24051,N_21489);
or UO_883 (O_883,N_20842,N_23557);
xor UO_884 (O_884,N_20241,N_24325);
or UO_885 (O_885,N_21124,N_24875);
and UO_886 (O_886,N_24542,N_22374);
or UO_887 (O_887,N_22463,N_22460);
xnor UO_888 (O_888,N_23755,N_22760);
nand UO_889 (O_889,N_24567,N_24997);
and UO_890 (O_890,N_21914,N_21808);
or UO_891 (O_891,N_20351,N_22074);
nor UO_892 (O_892,N_21151,N_24973);
nand UO_893 (O_893,N_24088,N_23249);
and UO_894 (O_894,N_22217,N_20266);
and UO_895 (O_895,N_22423,N_20093);
and UO_896 (O_896,N_23159,N_21263);
and UO_897 (O_897,N_23674,N_22688);
or UO_898 (O_898,N_23584,N_22399);
nor UO_899 (O_899,N_22372,N_21684);
nand UO_900 (O_900,N_24007,N_24389);
nand UO_901 (O_901,N_23620,N_24377);
or UO_902 (O_902,N_24289,N_21597);
or UO_903 (O_903,N_24663,N_20944);
nand UO_904 (O_904,N_20924,N_21185);
or UO_905 (O_905,N_24008,N_22242);
nand UO_906 (O_906,N_21505,N_21397);
nand UO_907 (O_907,N_24190,N_22555);
or UO_908 (O_908,N_24267,N_22163);
nor UO_909 (O_909,N_22726,N_22274);
or UO_910 (O_910,N_22059,N_22051);
and UO_911 (O_911,N_23206,N_20739);
nand UO_912 (O_912,N_24372,N_21579);
or UO_913 (O_913,N_22427,N_23533);
and UO_914 (O_914,N_22728,N_21650);
and UO_915 (O_915,N_21911,N_23512);
and UO_916 (O_916,N_24883,N_20298);
or UO_917 (O_917,N_24028,N_24323);
and UO_918 (O_918,N_22735,N_21601);
nand UO_919 (O_919,N_24758,N_21340);
and UO_920 (O_920,N_21682,N_22290);
and UO_921 (O_921,N_23519,N_23225);
nand UO_922 (O_922,N_20318,N_21317);
and UO_923 (O_923,N_24127,N_20496);
and UO_924 (O_924,N_20820,N_23552);
nand UO_925 (O_925,N_24005,N_21262);
nor UO_926 (O_926,N_21487,N_23834);
and UO_927 (O_927,N_22411,N_21483);
and UO_928 (O_928,N_20159,N_20643);
nand UO_929 (O_929,N_20313,N_23850);
or UO_930 (O_930,N_22357,N_24787);
nand UO_931 (O_931,N_21437,N_23426);
nand UO_932 (O_932,N_23626,N_24443);
and UO_933 (O_933,N_24585,N_24255);
nand UO_934 (O_934,N_23968,N_21741);
xnor UO_935 (O_935,N_24804,N_24212);
nor UO_936 (O_936,N_20824,N_22243);
or UO_937 (O_937,N_24753,N_21778);
and UO_938 (O_938,N_21558,N_24777);
or UO_939 (O_939,N_24041,N_22686);
nand UO_940 (O_940,N_23209,N_23361);
and UO_941 (O_941,N_21439,N_24706);
nand UO_942 (O_942,N_23783,N_23883);
and UO_943 (O_943,N_21711,N_24861);
and UO_944 (O_944,N_21313,N_22404);
or UO_945 (O_945,N_20561,N_21852);
or UO_946 (O_946,N_22917,N_24275);
nand UO_947 (O_947,N_22053,N_21260);
nand UO_948 (O_948,N_21907,N_21736);
nand UO_949 (O_949,N_20768,N_20289);
or UO_950 (O_950,N_23355,N_20016);
and UO_951 (O_951,N_21993,N_22868);
xor UO_952 (O_952,N_22133,N_24849);
nor UO_953 (O_953,N_22747,N_24971);
and UO_954 (O_954,N_21715,N_24784);
nor UO_955 (O_955,N_23358,N_21283);
or UO_956 (O_956,N_24863,N_24786);
nor UO_957 (O_957,N_20489,N_22610);
or UO_958 (O_958,N_22933,N_21453);
or UO_959 (O_959,N_23078,N_20525);
or UO_960 (O_960,N_23154,N_22305);
and UO_961 (O_961,N_20281,N_22856);
xor UO_962 (O_962,N_22335,N_22641);
nor UO_963 (O_963,N_20237,N_22337);
xnor UO_964 (O_964,N_20174,N_22203);
and UO_965 (O_965,N_21630,N_20211);
nand UO_966 (O_966,N_23390,N_21080);
or UO_967 (O_967,N_22577,N_24938);
xor UO_968 (O_968,N_21455,N_21327);
nor UO_969 (O_969,N_24812,N_24778);
or UO_970 (O_970,N_22127,N_24738);
nor UO_971 (O_971,N_22743,N_23118);
nand UO_972 (O_972,N_24801,N_20416);
and UO_973 (O_973,N_24659,N_20033);
or UO_974 (O_974,N_24437,N_23119);
nor UO_975 (O_975,N_23404,N_21841);
xnor UO_976 (O_976,N_24333,N_20780);
or UO_977 (O_977,N_24329,N_20748);
nand UO_978 (O_978,N_21459,N_24227);
and UO_979 (O_979,N_20491,N_24980);
nand UO_980 (O_980,N_24213,N_21696);
or UO_981 (O_981,N_24371,N_22379);
nor UO_982 (O_982,N_24882,N_23128);
and UO_983 (O_983,N_23957,N_22081);
or UO_984 (O_984,N_23388,N_22361);
or UO_985 (O_985,N_20075,N_21891);
or UO_986 (O_986,N_24016,N_24919);
or UO_987 (O_987,N_20521,N_21596);
and UO_988 (O_988,N_22309,N_20403);
nand UO_989 (O_989,N_21623,N_21413);
and UO_990 (O_990,N_24541,N_22402);
nand UO_991 (O_991,N_20124,N_24848);
nand UO_992 (O_992,N_24327,N_24291);
or UO_993 (O_993,N_22590,N_20437);
nand UO_994 (O_994,N_22825,N_23490);
or UO_995 (O_995,N_20583,N_23788);
nor UO_996 (O_996,N_22759,N_21273);
and UO_997 (O_997,N_20360,N_21179);
or UO_998 (O_998,N_24543,N_23143);
xor UO_999 (O_999,N_24963,N_24132);
nand UO_1000 (O_1000,N_20901,N_24197);
and UO_1001 (O_1001,N_23859,N_21344);
nand UO_1002 (O_1002,N_22446,N_22376);
nand UO_1003 (O_1003,N_23929,N_24089);
or UO_1004 (O_1004,N_21225,N_23798);
nand UO_1005 (O_1005,N_23169,N_21250);
nand UO_1006 (O_1006,N_22377,N_21624);
nor UO_1007 (O_1007,N_24890,N_20123);
nor UO_1008 (O_1008,N_24222,N_23396);
nor UO_1009 (O_1009,N_23924,N_23866);
or UO_1010 (O_1010,N_21411,N_24416);
and UO_1011 (O_1011,N_23718,N_20454);
and UO_1012 (O_1012,N_21774,N_23507);
nand UO_1013 (O_1013,N_22110,N_24461);
or UO_1014 (O_1014,N_22935,N_20380);
nor UO_1015 (O_1015,N_22418,N_21575);
nor UO_1016 (O_1016,N_21608,N_21011);
and UO_1017 (O_1017,N_22136,N_20511);
nor UO_1018 (O_1018,N_24160,N_22403);
or UO_1019 (O_1019,N_24392,N_22920);
nand UO_1020 (O_1020,N_23516,N_22809);
or UO_1021 (O_1021,N_24483,N_20460);
nand UO_1022 (O_1022,N_22512,N_20565);
nand UO_1023 (O_1023,N_23795,N_20545);
nand UO_1024 (O_1024,N_21866,N_21765);
nor UO_1025 (O_1025,N_24534,N_22782);
or UO_1026 (O_1026,N_24957,N_24021);
or UO_1027 (O_1027,N_20674,N_23618);
nand UO_1028 (O_1028,N_24305,N_20006);
or UO_1029 (O_1029,N_21908,N_24582);
or UO_1030 (O_1030,N_24552,N_21540);
and UO_1031 (O_1031,N_21625,N_23713);
xor UO_1032 (O_1032,N_21979,N_20308);
nand UO_1033 (O_1033,N_20339,N_23726);
nor UO_1034 (O_1034,N_20981,N_20290);
or UO_1035 (O_1035,N_20037,N_23294);
or UO_1036 (O_1036,N_23416,N_24399);
nor UO_1037 (O_1037,N_20919,N_20806);
or UO_1038 (O_1038,N_23330,N_22158);
xnor UO_1039 (O_1039,N_22756,N_20699);
nand UO_1040 (O_1040,N_24502,N_23921);
nor UO_1041 (O_1041,N_24814,N_24278);
xnor UO_1042 (O_1042,N_21917,N_21399);
nand UO_1043 (O_1043,N_22167,N_24065);
nor UO_1044 (O_1044,N_24467,N_22436);
xnor UO_1045 (O_1045,N_22270,N_21563);
or UO_1046 (O_1046,N_22978,N_21818);
nor UO_1047 (O_1047,N_22056,N_20877);
xnor UO_1048 (O_1048,N_23769,N_22333);
nor UO_1049 (O_1049,N_23362,N_21586);
nand UO_1050 (O_1050,N_20371,N_24025);
and UO_1051 (O_1051,N_21725,N_20188);
nand UO_1052 (O_1052,N_22498,N_24649);
nand UO_1053 (O_1053,N_23728,N_21163);
or UO_1054 (O_1054,N_24723,N_21665);
nor UO_1055 (O_1055,N_21402,N_22476);
and UO_1056 (O_1056,N_24902,N_22350);
and UO_1057 (O_1057,N_20600,N_23586);
or UO_1058 (O_1058,N_21817,N_23539);
nand UO_1059 (O_1059,N_20163,N_21401);
and UO_1060 (O_1060,N_23524,N_22016);
nor UO_1061 (O_1061,N_20096,N_23860);
and UO_1062 (O_1062,N_22221,N_23275);
nand UO_1063 (O_1063,N_21264,N_21662);
xor UO_1064 (O_1064,N_24834,N_22296);
or UO_1065 (O_1065,N_20908,N_22804);
and UO_1066 (O_1066,N_21096,N_21351);
nand UO_1067 (O_1067,N_24444,N_21157);
nor UO_1068 (O_1068,N_21269,N_23234);
xor UO_1069 (O_1069,N_21388,N_23965);
nor UO_1070 (O_1070,N_21687,N_24526);
nand UO_1071 (O_1071,N_23117,N_20728);
xnor UO_1072 (O_1072,N_22459,N_23233);
or UO_1073 (O_1073,N_24732,N_22509);
xnor UO_1074 (O_1074,N_20601,N_20404);
and UO_1075 (O_1075,N_24969,N_22835);
or UO_1076 (O_1076,N_23324,N_20134);
or UO_1077 (O_1077,N_23002,N_24062);
nor UO_1078 (O_1078,N_23905,N_21126);
nor UO_1079 (O_1079,N_23075,N_22833);
or UO_1080 (O_1080,N_22302,N_21768);
nand UO_1081 (O_1081,N_22566,N_21146);
and UO_1082 (O_1082,N_21303,N_20630);
or UO_1083 (O_1083,N_23941,N_24411);
or UO_1084 (O_1084,N_23182,N_20615);
and UO_1085 (O_1085,N_21153,N_23126);
nand UO_1086 (O_1086,N_20447,N_24380);
xnor UO_1087 (O_1087,N_20691,N_22220);
nand UO_1088 (O_1088,N_20436,N_23171);
or UO_1089 (O_1089,N_22864,N_20838);
nand UO_1090 (O_1090,N_24506,N_21989);
or UO_1091 (O_1091,N_21082,N_23508);
nor UO_1092 (O_1092,N_20423,N_22119);
and UO_1093 (O_1093,N_22860,N_24162);
nand UO_1094 (O_1094,N_24761,N_24958);
nor UO_1095 (O_1095,N_24925,N_23525);
nand UO_1096 (O_1096,N_21139,N_24688);
or UO_1097 (O_1097,N_24895,N_21971);
nand UO_1098 (O_1098,N_20058,N_21374);
nor UO_1099 (O_1099,N_23704,N_21618);
and UO_1100 (O_1100,N_23904,N_21432);
or UO_1101 (O_1101,N_22251,N_22389);
nor UO_1102 (O_1102,N_22125,N_21071);
or UO_1103 (O_1103,N_22355,N_22791);
and UO_1104 (O_1104,N_20961,N_20913);
or UO_1105 (O_1105,N_22534,N_20455);
nor UO_1106 (O_1106,N_23401,N_23283);
nand UO_1107 (O_1107,N_24322,N_20917);
and UO_1108 (O_1108,N_24302,N_20009);
nor UO_1109 (O_1109,N_20247,N_23168);
nor UO_1110 (O_1110,N_23254,N_23761);
nand UO_1111 (O_1111,N_22019,N_22354);
and UO_1112 (O_1112,N_20158,N_22035);
nor UO_1113 (O_1113,N_24782,N_22306);
and UO_1114 (O_1114,N_24744,N_23060);
nand UO_1115 (O_1115,N_23601,N_21614);
and UO_1116 (O_1116,N_21007,N_24012);
nand UO_1117 (O_1117,N_24513,N_23457);
xnor UO_1118 (O_1118,N_21663,N_24352);
and UO_1119 (O_1119,N_21256,N_23714);
and UO_1120 (O_1120,N_23544,N_20695);
nand UO_1121 (O_1121,N_21779,N_24099);
or UO_1122 (O_1122,N_23336,N_22638);
and UO_1123 (O_1123,N_23776,N_21807);
and UO_1124 (O_1124,N_23383,N_23727);
and UO_1125 (O_1125,N_20811,N_24395);
and UO_1126 (O_1126,N_24595,N_24344);
and UO_1127 (O_1127,N_21942,N_20128);
and UO_1128 (O_1128,N_22676,N_22949);
or UO_1129 (O_1129,N_21480,N_22021);
nor UO_1130 (O_1130,N_20230,N_22729);
nand UO_1131 (O_1131,N_20873,N_22201);
xor UO_1132 (O_1132,N_24792,N_22700);
and UO_1133 (O_1133,N_23016,N_21583);
xnor UO_1134 (O_1134,N_23731,N_23291);
nor UO_1135 (O_1135,N_21427,N_23978);
or UO_1136 (O_1136,N_20589,N_20261);
or UO_1137 (O_1137,N_24040,N_23110);
or UO_1138 (O_1138,N_21709,N_22075);
or UO_1139 (O_1139,N_22951,N_20696);
xnor UO_1140 (O_1140,N_23622,N_20742);
or UO_1141 (O_1141,N_23149,N_23484);
and UO_1142 (O_1142,N_22096,N_21010);
nor UO_1143 (O_1143,N_24776,N_20717);
and UO_1144 (O_1144,N_24175,N_21078);
xor UO_1145 (O_1145,N_20377,N_21899);
nor UO_1146 (O_1146,N_22691,N_22922);
nand UO_1147 (O_1147,N_20883,N_20706);
nand UO_1148 (O_1148,N_24817,N_24094);
nor UO_1149 (O_1149,N_22583,N_22287);
or UO_1150 (O_1150,N_22675,N_20569);
or UO_1151 (O_1151,N_22844,N_21972);
and UO_1152 (O_1152,N_23458,N_23833);
and UO_1153 (O_1153,N_22491,N_23939);
and UO_1154 (O_1154,N_21119,N_23033);
nand UO_1155 (O_1155,N_21834,N_20100);
xor UO_1156 (O_1156,N_21029,N_21135);
nor UO_1157 (O_1157,N_20480,N_24072);
and UO_1158 (O_1158,N_24579,N_20161);
nor UO_1159 (O_1159,N_21702,N_23466);
nand UO_1160 (O_1160,N_20591,N_21506);
nor UO_1161 (O_1161,N_20744,N_21636);
xnor UO_1162 (O_1162,N_20730,N_23616);
xnor UO_1163 (O_1163,N_22581,N_22324);
nand UO_1164 (O_1164,N_24472,N_21106);
or UO_1165 (O_1165,N_23063,N_23660);
nand UO_1166 (O_1166,N_23345,N_23381);
nor UO_1167 (O_1167,N_22944,N_21632);
nand UO_1168 (O_1168,N_21913,N_22772);
nand UO_1169 (O_1169,N_21659,N_21813);
or UO_1170 (O_1170,N_21343,N_21054);
or UO_1171 (O_1171,N_23670,N_22849);
nor UO_1172 (O_1172,N_23723,N_23588);
xnor UO_1173 (O_1173,N_20328,N_23074);
or UO_1174 (O_1174,N_22406,N_22539);
nand UO_1175 (O_1175,N_20593,N_22677);
nor UO_1176 (O_1176,N_22307,N_23922);
nor UO_1177 (O_1177,N_24916,N_20107);
nand UO_1178 (O_1178,N_20401,N_22079);
or UO_1179 (O_1179,N_22434,N_20199);
and UO_1180 (O_1180,N_24312,N_22937);
nand UO_1181 (O_1181,N_24488,N_23464);
and UO_1182 (O_1182,N_21278,N_21073);
or UO_1183 (O_1183,N_23068,N_23807);
and UO_1184 (O_1184,N_22980,N_23346);
nand UO_1185 (O_1185,N_21707,N_23678);
nor UO_1186 (O_1186,N_23805,N_24439);
nor UO_1187 (O_1187,N_23064,N_21503);
nor UO_1188 (O_1188,N_22820,N_23163);
or UO_1189 (O_1189,N_20915,N_23007);
nor UO_1190 (O_1190,N_21819,N_22345);
nand UO_1191 (O_1191,N_24497,N_20372);
nand UO_1192 (O_1192,N_20580,N_23858);
or UO_1193 (O_1193,N_21449,N_20213);
nand UO_1194 (O_1194,N_23014,N_23936);
or UO_1195 (O_1195,N_22710,N_24704);
nand UO_1196 (O_1196,N_20831,N_23611);
or UO_1197 (O_1197,N_20118,N_24445);
xor UO_1198 (O_1198,N_23874,N_23192);
nor UO_1199 (O_1199,N_24678,N_20638);
nor UO_1200 (O_1200,N_21857,N_23750);
or UO_1201 (O_1201,N_21870,N_24074);
nor UO_1202 (O_1202,N_22405,N_21853);
and UO_1203 (O_1203,N_21137,N_24083);
nand UO_1204 (O_1204,N_23337,N_24112);
and UO_1205 (O_1205,N_21876,N_23948);
nor UO_1206 (O_1206,N_23806,N_24975);
xnor UO_1207 (O_1207,N_21245,N_23247);
nor UO_1208 (O_1208,N_24521,N_20875);
or UO_1209 (O_1209,N_23222,N_23700);
nand UO_1210 (O_1210,N_22781,N_24859);
or UO_1211 (O_1211,N_22486,N_21446);
nand UO_1212 (O_1212,N_21844,N_23315);
nand UO_1213 (O_1213,N_21764,N_20349);
nor UO_1214 (O_1214,N_23311,N_22188);
and UO_1215 (O_1215,N_20133,N_20260);
nand UO_1216 (O_1216,N_24379,N_22477);
or UO_1217 (O_1217,N_21810,N_21381);
nand UO_1218 (O_1218,N_21294,N_20257);
and UO_1219 (O_1219,N_24956,N_24063);
nor UO_1220 (O_1220,N_21798,N_20382);
nand UO_1221 (O_1221,N_23852,N_22321);
nor UO_1222 (O_1222,N_22588,N_23313);
nand UO_1223 (O_1223,N_20094,N_20997);
nor UO_1224 (O_1224,N_21693,N_20813);
xor UO_1225 (O_1225,N_21038,N_23813);
or UO_1226 (O_1226,N_20882,N_23691);
xnor UO_1227 (O_1227,N_22058,N_24337);
or UO_1228 (O_1228,N_22055,N_22114);
nor UO_1229 (O_1229,N_23495,N_23528);
or UO_1230 (O_1230,N_24420,N_23675);
nor UO_1231 (O_1231,N_22289,N_20669);
nor UO_1232 (O_1232,N_21981,N_23964);
xnor UO_1233 (O_1233,N_23951,N_22279);
and UO_1234 (O_1234,N_22986,N_24632);
nor UO_1235 (O_1235,N_20005,N_20978);
or UO_1236 (O_1236,N_22360,N_24945);
nor UO_1237 (O_1237,N_20494,N_23450);
or UO_1238 (O_1238,N_21730,N_22394);
or UO_1239 (O_1239,N_21098,N_21691);
or UO_1240 (O_1240,N_20733,N_24662);
nor UO_1241 (O_1241,N_23419,N_24565);
and UO_1242 (O_1242,N_21481,N_24696);
nand UO_1243 (O_1243,N_21442,N_22237);
nor UO_1244 (O_1244,N_23176,N_21297);
nor UO_1245 (O_1245,N_21093,N_23540);
and UO_1246 (O_1246,N_24520,N_24053);
nor UO_1247 (O_1247,N_22975,N_20977);
and UO_1248 (O_1248,N_20297,N_22154);
nand UO_1249 (O_1249,N_21363,N_24143);
and UO_1250 (O_1250,N_21685,N_20797);
nand UO_1251 (O_1251,N_22973,N_21613);
and UO_1252 (O_1252,N_22202,N_23600);
xor UO_1253 (O_1253,N_22124,N_22024);
nor UO_1254 (O_1254,N_20657,N_20777);
xor UO_1255 (O_1255,N_20492,N_22177);
and UO_1256 (O_1256,N_22672,N_23386);
and UO_1257 (O_1257,N_23245,N_20990);
or UO_1258 (O_1258,N_21237,N_21534);
nand UO_1259 (O_1259,N_22776,N_21460);
nand UO_1260 (O_1260,N_24250,N_21122);
nand UO_1261 (O_1261,N_24139,N_22886);
and UO_1262 (O_1262,N_22543,N_23445);
or UO_1263 (O_1263,N_23535,N_20888);
nand UO_1264 (O_1264,N_20288,N_23327);
nand UO_1265 (O_1265,N_20634,N_24183);
or UO_1266 (O_1266,N_22214,N_22496);
or UO_1267 (O_1267,N_23823,N_23721);
or UO_1268 (O_1268,N_22301,N_23803);
nand UO_1269 (O_1269,N_23801,N_22168);
nor UO_1270 (O_1270,N_22503,N_24586);
xnor UO_1271 (O_1271,N_23677,N_20715);
xnor UO_1272 (O_1272,N_24216,N_20198);
or UO_1273 (O_1273,N_24457,N_22673);
nor UO_1274 (O_1274,N_22410,N_24280);
nand UO_1275 (O_1275,N_20949,N_24989);
nor UO_1276 (O_1276,N_20182,N_23351);
or UO_1277 (O_1277,N_20825,N_21923);
nor UO_1278 (O_1278,N_24653,N_24475);
nand UO_1279 (O_1279,N_20687,N_23802);
or UO_1280 (O_1280,N_21047,N_22153);
nor UO_1281 (O_1281,N_24645,N_22175);
or UO_1282 (O_1282,N_24745,N_24922);
xor UO_1283 (O_1283,N_22089,N_24482);
or UO_1284 (O_1284,N_21786,N_24047);
xor UO_1285 (O_1285,N_23578,N_20896);
and UO_1286 (O_1286,N_23449,N_20789);
nor UO_1287 (O_1287,N_20850,N_22900);
and UO_1288 (O_1288,N_20388,N_23412);
nor UO_1289 (O_1289,N_20649,N_20965);
or UO_1290 (O_1290,N_20727,N_20903);
nand UO_1291 (O_1291,N_21990,N_24691);
and UO_1292 (O_1292,N_23114,N_21763);
nand UO_1293 (O_1293,N_23278,N_21258);
or UO_1294 (O_1294,N_20890,N_22304);
nor UO_1295 (O_1295,N_21789,N_21454);
and UO_1296 (O_1296,N_24816,N_22537);
nor UO_1297 (O_1297,N_22565,N_22181);
and UO_1298 (O_1298,N_22066,N_22636);
and UO_1299 (O_1299,N_24637,N_23470);
nand UO_1300 (O_1300,N_22637,N_23056);
or UO_1301 (O_1301,N_21761,N_20612);
nor UO_1302 (O_1302,N_22725,N_20419);
and UO_1303 (O_1303,N_23632,N_24754);
nand UO_1304 (O_1304,N_22991,N_22657);
nor UO_1305 (O_1305,N_22501,N_22652);
nor UO_1306 (O_1306,N_20265,N_23217);
nor UO_1307 (O_1307,N_24710,N_20021);
or UO_1308 (O_1308,N_23784,N_20764);
and UO_1309 (O_1309,N_21107,N_20930);
nand UO_1310 (O_1310,N_20064,N_24518);
or UO_1311 (O_1311,N_22022,N_20594);
nor UO_1312 (O_1312,N_21796,N_21086);
nand UO_1313 (O_1313,N_22983,N_21629);
nand UO_1314 (O_1314,N_24791,N_21016);
nand UO_1315 (O_1315,N_23885,N_20422);
nor UO_1316 (O_1316,N_22589,N_20383);
xnor UO_1317 (O_1317,N_21775,N_24248);
nor UO_1318 (O_1318,N_21326,N_23537);
nand UO_1319 (O_1319,N_24596,N_20808);
and UO_1320 (O_1320,N_24317,N_21406);
nand UO_1321 (O_1321,N_24944,N_24911);
nor UO_1322 (O_1322,N_23230,N_24713);
and UO_1323 (O_1323,N_24576,N_23625);
or UO_1324 (O_1324,N_23444,N_24128);
and UO_1325 (O_1325,N_24169,N_24674);
nor UO_1326 (O_1326,N_22853,N_20292);
or UO_1327 (O_1327,N_20884,N_22805);
xor UO_1328 (O_1328,N_24428,N_22003);
and UO_1329 (O_1329,N_22443,N_24574);
xor UO_1330 (O_1330,N_23706,N_24064);
and UO_1331 (O_1331,N_24718,N_22429);
nor UO_1332 (O_1332,N_24184,N_24623);
nor UO_1333 (O_1333,N_20656,N_24236);
and UO_1334 (O_1334,N_21255,N_21783);
or UO_1335 (O_1335,N_24599,N_20203);
nand UO_1336 (O_1336,N_23084,N_23607);
nor UO_1337 (O_1337,N_21198,N_23488);
and UO_1338 (O_1338,N_21275,N_22223);
or UO_1339 (O_1339,N_20554,N_21102);
or UO_1340 (O_1340,N_24281,N_24406);
nand UO_1341 (O_1341,N_22716,N_21576);
nor UO_1342 (O_1342,N_24463,N_23934);
or UO_1343 (O_1343,N_24712,N_20146);
nand UO_1344 (O_1344,N_24332,N_22874);
or UO_1345 (O_1345,N_22684,N_21965);
nor UO_1346 (O_1346,N_23039,N_24553);
nand UO_1347 (O_1347,N_21919,N_21099);
nor UO_1348 (O_1348,N_23966,N_20067);
xor UO_1349 (O_1349,N_21053,N_20775);
nor UO_1350 (O_1350,N_22640,N_23547);
or UO_1351 (O_1351,N_23561,N_20280);
and UO_1352 (O_1352,N_21664,N_24986);
and UO_1353 (O_1353,N_22012,N_22662);
nor UO_1354 (O_1354,N_20794,N_20799);
and UO_1355 (O_1355,N_23898,N_23736);
and UO_1356 (O_1356,N_21305,N_20258);
and UO_1357 (O_1357,N_21484,N_24200);
nor UO_1358 (O_1358,N_20311,N_22005);
xnor UO_1359 (O_1359,N_21974,N_20592);
and UO_1360 (O_1360,N_24022,N_24939);
and UO_1361 (O_1361,N_20074,N_24729);
nand UO_1362 (O_1362,N_20394,N_21282);
nor UO_1363 (O_1363,N_21612,N_22752);
nor UO_1364 (O_1364,N_24705,N_24836);
or UO_1365 (O_1365,N_24799,N_23219);
and UO_1366 (O_1366,N_21049,N_20196);
and UO_1367 (O_1367,N_23725,N_20413);
and UO_1368 (O_1368,N_21516,N_20670);
or UO_1369 (O_1369,N_23170,N_23511);
nand UO_1370 (O_1370,N_23950,N_24675);
nand UO_1371 (O_1371,N_24824,N_24952);
and UO_1372 (O_1372,N_24505,N_23943);
and UO_1373 (O_1373,N_23583,N_21173);
and UO_1374 (O_1374,N_22344,N_24953);
and UO_1375 (O_1375,N_22755,N_22996);
or UO_1376 (O_1376,N_24808,N_24523);
nand UO_1377 (O_1377,N_21338,N_22332);
or UO_1378 (O_1378,N_20772,N_20743);
xnor UO_1379 (O_1379,N_20747,N_20979);
nor UO_1380 (O_1380,N_23221,N_22771);
nand UO_1381 (O_1381,N_21112,N_22741);
and UO_1382 (O_1382,N_21299,N_20164);
nand UO_1383 (O_1383,N_22128,N_21199);
and UO_1384 (O_1384,N_20119,N_21539);
nor UO_1385 (O_1385,N_24993,N_20415);
or UO_1386 (O_1386,N_21134,N_20631);
nor UO_1387 (O_1387,N_23764,N_23868);
or UO_1388 (O_1388,N_23433,N_22631);
nor UO_1389 (O_1389,N_22956,N_23070);
xor UO_1390 (O_1390,N_24262,N_20573);
nand UO_1391 (O_1391,N_24810,N_21013);
or UO_1392 (O_1392,N_20956,N_20218);
or UO_1393 (O_1393,N_22368,N_22183);
or UO_1394 (O_1394,N_24646,N_20463);
and UO_1395 (O_1395,N_23055,N_24864);
and UO_1396 (O_1396,N_20219,N_20845);
nor UO_1397 (O_1397,N_24915,N_23009);
nor UO_1398 (O_1398,N_21962,N_22313);
and UO_1399 (O_1399,N_23279,N_20495);
xnor UO_1400 (O_1400,N_22475,N_21204);
nand UO_1401 (O_1401,N_21280,N_21216);
and UO_1402 (O_1402,N_20268,N_20259);
nand UO_1403 (O_1403,N_23380,N_22668);
and UO_1404 (O_1404,N_24770,N_21875);
nand UO_1405 (O_1405,N_20547,N_24563);
nor UO_1406 (O_1406,N_21145,N_23520);
or UO_1407 (O_1407,N_24735,N_21422);
and UO_1408 (O_1408,N_22569,N_24393);
xor UO_1409 (O_1409,N_20379,N_23639);
nor UO_1410 (O_1410,N_22111,N_22199);
and UO_1411 (O_1411,N_20673,N_20970);
nor UO_1412 (O_1412,N_24233,N_23738);
xor UO_1413 (O_1413,N_21643,N_24878);
or UO_1414 (O_1414,N_22834,N_23991);
nand UO_1415 (O_1415,N_24855,N_21443);
or UO_1416 (O_1416,N_22232,N_24013);
nor UO_1417 (O_1417,N_20867,N_22044);
or UO_1418 (O_1418,N_24932,N_21471);
xor UO_1419 (O_1419,N_21690,N_21661);
xnor UO_1420 (O_1420,N_21114,N_24441);
and UO_1421 (O_1421,N_22367,N_23628);
nand UO_1422 (O_1422,N_21713,N_21324);
and UO_1423 (O_1423,N_22941,N_24589);
or UO_1424 (O_1424,N_23178,N_24821);
and UO_1425 (O_1425,N_23242,N_23749);
or UO_1426 (O_1426,N_23151,N_20553);
or UO_1427 (O_1427,N_22552,N_24519);
or UO_1428 (O_1428,N_21681,N_22918);
nand UO_1429 (O_1429,N_21223,N_20365);
or UO_1430 (O_1430,N_23559,N_22663);
or UO_1431 (O_1431,N_21148,N_21440);
nand UO_1432 (O_1432,N_20291,N_23284);
and UO_1433 (O_1433,N_23634,N_21697);
and UO_1434 (O_1434,N_22171,N_21879);
and UO_1435 (O_1435,N_24603,N_21341);
or UO_1436 (O_1436,N_21568,N_21647);
and UO_1437 (O_1437,N_22892,N_22968);
nand UO_1438 (O_1438,N_20396,N_21293);
or UO_1439 (O_1439,N_23094,N_23796);
nor UO_1440 (O_1440,N_21329,N_24427);
nand UO_1441 (O_1441,N_24601,N_23510);
nand UO_1442 (O_1442,N_24967,N_23530);
nor UO_1443 (O_1443,N_23672,N_21814);
or UO_1444 (O_1444,N_23081,N_21322);
nor UO_1445 (O_1445,N_24593,N_23500);
and UO_1446 (O_1446,N_23040,N_20644);
or UO_1447 (O_1447,N_24124,N_22536);
or UO_1448 (O_1448,N_20769,N_21700);
nand UO_1449 (O_1449,N_20807,N_22104);
nor UO_1450 (O_1450,N_24134,N_24701);
and UO_1451 (O_1451,N_20072,N_20039);
nor UO_1452 (O_1452,N_22031,N_22919);
or UO_1453 (O_1453,N_23184,N_20029);
and UO_1454 (O_1454,N_21584,N_23347);
or UO_1455 (O_1455,N_24006,N_22380);
or UO_1456 (O_1456,N_20304,N_20445);
nand UO_1457 (O_1457,N_22701,N_21190);
nor UO_1458 (O_1458,N_24525,N_20659);
or UO_1459 (O_1459,N_23020,N_24103);
nor UO_1460 (O_1460,N_22758,N_22126);
and UO_1461 (O_1461,N_24837,N_23197);
or UO_1462 (O_1462,N_22086,N_22542);
nand UO_1463 (O_1463,N_24716,N_20648);
nand UO_1464 (O_1464,N_22827,N_24116);
and UO_1465 (O_1465,N_24652,N_21318);
and UO_1466 (O_1466,N_20175,N_23309);
nor UO_1467 (O_1467,N_23742,N_23354);
nor UO_1468 (O_1468,N_20782,N_20070);
and UO_1469 (O_1469,N_22932,N_23992);
or UO_1470 (O_1470,N_22823,N_22604);
xor UO_1471 (O_1471,N_21890,N_20059);
nand UO_1472 (O_1472,N_23724,N_22665);
and UO_1473 (O_1473,N_24432,N_23534);
nand UO_1474 (O_1474,N_24668,N_21319);
nor UO_1475 (O_1475,N_24219,N_24480);
and UO_1476 (O_1476,N_22832,N_21551);
and UO_1477 (O_1477,N_21004,N_22585);
nor UO_1478 (O_1478,N_22850,N_24954);
xnor UO_1479 (O_1479,N_21136,N_21308);
nor UO_1480 (O_1480,N_24168,N_21384);
or UO_1481 (O_1481,N_21431,N_22444);
or UO_1482 (O_1482,N_20502,N_24880);
or UO_1483 (O_1483,N_20095,N_22291);
nand UO_1484 (O_1484,N_22041,N_21105);
xnor UO_1485 (O_1485,N_21877,N_22876);
nor UO_1486 (O_1486,N_23329,N_20336);
nor UO_1487 (O_1487,N_20127,N_23971);
or UO_1488 (O_1488,N_24318,N_23101);
and UO_1489 (O_1489,N_22736,N_24039);
nand UO_1490 (O_1490,N_20579,N_21166);
nor UO_1491 (O_1491,N_20277,N_24272);
nor UO_1492 (O_1492,N_20490,N_22938);
nor UO_1493 (O_1493,N_21840,N_23656);
and UO_1494 (O_1494,N_23052,N_24715);
and UO_1495 (O_1495,N_24243,N_20967);
and UO_1496 (O_1496,N_23043,N_24988);
or UO_1497 (O_1497,N_24903,N_22458);
and UO_1498 (O_1498,N_21438,N_24218);
nand UO_1499 (O_1499,N_22855,N_21236);
and UO_1500 (O_1500,N_20329,N_24114);
nand UO_1501 (O_1501,N_22490,N_22828);
nor UO_1502 (O_1502,N_20737,N_20425);
nand UO_1503 (O_1503,N_24860,N_24917);
nor UO_1504 (O_1504,N_21030,N_22258);
nand UO_1505 (O_1505,N_21572,N_20000);
nand UO_1506 (O_1506,N_20703,N_24608);
nor UO_1507 (O_1507,N_22616,N_24011);
and UO_1508 (O_1508,N_24826,N_21334);
and UO_1509 (O_1509,N_24150,N_20597);
or UO_1510 (O_1510,N_20243,N_22351);
nor UO_1511 (O_1511,N_23712,N_24460);
or UO_1512 (O_1512,N_22687,N_22623);
nor UO_1513 (O_1513,N_23923,N_22017);
nand UO_1514 (O_1514,N_21809,N_20242);
or UO_1515 (O_1515,N_22659,N_20902);
nor UO_1516 (O_1516,N_23927,N_21091);
xor UO_1517 (O_1517,N_20407,N_22470);
nand UO_1518 (O_1518,N_21387,N_20528);
or UO_1519 (O_1519,N_20473,N_22186);
nand UO_1520 (O_1520,N_23000,N_23982);
and UO_1521 (O_1521,N_23790,N_21069);
or UO_1522 (O_1522,N_24644,N_22671);
nand UO_1523 (O_1523,N_21067,N_21380);
or UO_1524 (O_1524,N_20226,N_23899);
and UO_1525 (O_1525,N_21969,N_21208);
nor UO_1526 (O_1526,N_20169,N_23137);
nor UO_1527 (O_1527,N_22499,N_23423);
nand UO_1528 (O_1528,N_24906,N_20898);
nand UO_1529 (O_1529,N_20566,N_22316);
and UO_1530 (O_1530,N_20275,N_22241);
xnor UO_1531 (O_1531,N_21723,N_24138);
nand UO_1532 (O_1532,N_24719,N_22514);
nor UO_1533 (O_1533,N_20700,N_21555);
and UO_1534 (O_1534,N_20572,N_21992);
and UO_1535 (O_1535,N_23779,N_20205);
and UO_1536 (O_1536,N_20474,N_24887);
and UO_1537 (O_1537,N_21019,N_23133);
and UO_1538 (O_1538,N_23322,N_22065);
or UO_1539 (O_1539,N_24624,N_23869);
nor UO_1540 (O_1540,N_23059,N_20556);
nand UO_1541 (O_1541,N_23917,N_21020);
or UO_1542 (O_1542,N_20832,N_21202);
nor UO_1543 (O_1543,N_20305,N_22092);
nand UO_1544 (O_1544,N_23270,N_24037);
nand UO_1545 (O_1545,N_24604,N_22764);
nor UO_1546 (O_1546,N_21220,N_23871);
nor UO_1547 (O_1547,N_20048,N_20364);
nor UO_1548 (O_1548,N_24643,N_23017);
or UO_1549 (O_1549,N_22036,N_20056);
and UO_1550 (O_1550,N_24203,N_21252);
nand UO_1551 (O_1551,N_23031,N_21985);
and UO_1552 (O_1552,N_23485,N_24690);
or UO_1553 (O_1553,N_20486,N_20533);
xnor UO_1554 (O_1554,N_20987,N_20709);
or UO_1555 (O_1555,N_22343,N_22733);
nand UO_1556 (O_1556,N_20632,N_21585);
or UO_1557 (O_1557,N_22145,N_23666);
or UO_1558 (O_1558,N_24466,N_23104);
and UO_1559 (O_1559,N_23986,N_22863);
and UO_1560 (O_1560,N_24580,N_22841);
nand UO_1561 (O_1561,N_20512,N_23042);
nor UO_1562 (O_1562,N_22899,N_24700);
nor UO_1563 (O_1563,N_20157,N_20215);
and UO_1564 (O_1564,N_20220,N_24239);
nand UO_1565 (O_1565,N_21393,N_23012);
nand UO_1566 (O_1566,N_22661,N_21973);
nand UO_1567 (O_1567,N_23812,N_20611);
nand UO_1568 (O_1568,N_24186,N_24029);
nand UO_1569 (O_1569,N_24921,N_20111);
nand UO_1570 (O_1570,N_21941,N_21637);
and UO_1571 (O_1571,N_21496,N_20347);
nand UO_1572 (O_1572,N_23447,N_24285);
and UO_1573 (O_1573,N_22213,N_21918);
and UO_1574 (O_1574,N_23338,N_22533);
nor UO_1575 (O_1575,N_24811,N_24489);
and UO_1576 (O_1576,N_21640,N_24364);
nand UO_1577 (O_1577,N_23290,N_20233);
and UO_1578 (O_1578,N_20889,N_21638);
or UO_1579 (O_1579,N_20356,N_20301);
nor UO_1580 (O_1580,N_23781,N_24087);
nor UO_1581 (O_1581,N_23919,N_21646);
or UO_1582 (O_1582,N_22454,N_21541);
nor UO_1583 (O_1583,N_24549,N_21648);
and UO_1584 (O_1584,N_20156,N_20905);
or UO_1585 (O_1585,N_21425,N_23480);
or UO_1586 (O_1586,N_21546,N_21159);
nand UO_1587 (O_1587,N_20524,N_22883);
or UO_1588 (O_1588,N_22416,N_24034);
nand UO_1589 (O_1589,N_22082,N_22546);
or UO_1590 (O_1590,N_24947,N_20088);
nor UO_1591 (O_1591,N_24905,N_23312);
and UO_1592 (O_1592,N_20089,N_21290);
or UO_1593 (O_1593,N_24620,N_24561);
nor UO_1594 (O_1594,N_24228,N_21174);
nor UO_1595 (O_1595,N_24796,N_24176);
nor UO_1596 (O_1596,N_24269,N_22176);
nor UO_1597 (O_1597,N_23596,N_21021);
nor UO_1598 (O_1598,N_21905,N_24907);
and UO_1599 (O_1599,N_20069,N_22047);
nor UO_1600 (O_1600,N_24617,N_22522);
nor UO_1601 (O_1601,N_24303,N_20200);
or UO_1602 (O_1602,N_23453,N_23577);
nor UO_1603 (O_1603,N_21544,N_22654);
and UO_1604 (O_1604,N_24253,N_22811);
or UO_1605 (O_1605,N_24684,N_21897);
nor UO_1606 (O_1606,N_21880,N_21366);
nand UO_1607 (O_1607,N_20665,N_21265);
nor UO_1608 (O_1608,N_22113,N_20025);
or UO_1609 (O_1609,N_20287,N_20061);
nor UO_1610 (O_1610,N_23397,N_23479);
nor UO_1611 (O_1611,N_21677,N_20019);
nor UO_1612 (O_1612,N_22116,N_21900);
or UO_1613 (O_1613,N_22974,N_23403);
nor UO_1614 (O_1614,N_23983,N_21960);
and UO_1615 (O_1615,N_22030,N_22957);
nor UO_1616 (O_1616,N_21435,N_24019);
nand UO_1617 (O_1617,N_22295,N_23274);
and UO_1618 (O_1618,N_24122,N_21143);
xnor UO_1619 (O_1619,N_22369,N_21552);
nand UO_1620 (O_1620,N_23637,N_24557);
nor UO_1621 (O_1621,N_21892,N_20142);
or UO_1622 (O_1622,N_23954,N_23384);
nand UO_1623 (O_1623,N_24985,N_22813);
and UO_1624 (O_1624,N_23940,N_20181);
and UO_1625 (O_1625,N_23642,N_20176);
nor UO_1626 (O_1626,N_20122,N_22703);
and UO_1627 (O_1627,N_23387,N_21926);
or UO_1628 (O_1628,N_21631,N_21084);
xnor UO_1629 (O_1629,N_21300,N_20729);
nand UO_1630 (O_1630,N_24870,N_23252);
nand UO_1631 (O_1631,N_22790,N_24180);
and UO_1632 (O_1632,N_22121,N_21894);
or UO_1633 (O_1633,N_20034,N_24301);
xor UO_1634 (O_1634,N_22364,N_23189);
nor UO_1635 (O_1635,N_23698,N_22105);
and UO_1636 (O_1636,N_22762,N_24923);
or UO_1637 (O_1637,N_22594,N_24459);
and UO_1638 (O_1638,N_22137,N_24607);
nor UO_1639 (O_1639,N_23875,N_22497);
nand UO_1640 (O_1640,N_21964,N_22327);
xor UO_1641 (O_1641,N_22048,N_21784);
or UO_1642 (O_1642,N_22622,N_21014);
nor UO_1643 (O_1643,N_22015,N_22315);
nor UO_1644 (O_1644,N_24894,N_20279);
xor UO_1645 (O_1645,N_24119,N_22836);
xor UO_1646 (O_1646,N_22083,N_22299);
nor UO_1647 (O_1647,N_21488,N_23425);
nor UO_1648 (O_1648,N_22878,N_20452);
and UO_1649 (O_1649,N_23873,N_20549);
nand UO_1650 (O_1650,N_20983,N_23877);
and UO_1651 (O_1651,N_20862,N_21704);
nand UO_1652 (O_1652,N_23452,N_24152);
and UO_1653 (O_1653,N_22619,N_22040);
nor UO_1654 (O_1654,N_20114,N_21562);
or UO_1655 (O_1655,N_24756,N_22865);
nand UO_1656 (O_1656,N_21826,N_24308);
nand UO_1657 (O_1657,N_20629,N_23624);
xor UO_1658 (O_1658,N_22447,N_21520);
and UO_1659 (O_1659,N_21085,N_21315);
and UO_1660 (O_1660,N_23590,N_22993);
nand UO_1661 (O_1661,N_24345,N_20837);
nor UO_1662 (O_1662,N_24910,N_22162);
and UO_1663 (O_1663,N_21792,N_20223);
and UO_1664 (O_1664,N_24664,N_24838);
nor UO_1665 (O_1665,N_23962,N_24307);
or UO_1666 (O_1666,N_21649,N_22222);
nor UO_1667 (O_1667,N_21769,N_24191);
xor UO_1668 (O_1668,N_20319,N_23004);
nand UO_1669 (O_1669,N_22795,N_20931);
or UO_1670 (O_1670,N_24147,N_20451);
or UO_1671 (O_1671,N_23615,N_22964);
and UO_1672 (O_1672,N_20020,N_22902);
and UO_1673 (O_1673,N_24976,N_23036);
and UO_1674 (O_1674,N_24606,N_21301);
nand UO_1675 (O_1675,N_24283,N_20893);
or UO_1676 (O_1676,N_23920,N_23669);
nor UO_1677 (O_1677,N_24661,N_20373);
and UO_1678 (O_1678,N_20350,N_20564);
xnor UO_1679 (O_1679,N_24876,N_23553);
nand UO_1680 (O_1680,N_20147,N_22715);
nand UO_1681 (O_1681,N_22656,N_23228);
and UO_1682 (O_1682,N_23427,N_21797);
or UO_1683 (O_1683,N_22090,N_22263);
and UO_1684 (O_1684,N_24033,N_23879);
and UO_1685 (O_1685,N_22381,N_24397);
or UO_1686 (O_1686,N_21400,N_20090);
nand UO_1687 (O_1687,N_20125,N_23817);
nor UO_1688 (O_1688,N_22164,N_20325);
xor UO_1689 (O_1689,N_21869,N_20542);
or UO_1690 (O_1690,N_21896,N_20303);
or UO_1691 (O_1691,N_23265,N_23641);
xor UO_1692 (O_1692,N_20899,N_23494);
nor UO_1693 (O_1693,N_24015,N_21087);
or UO_1694 (O_1694,N_24677,N_20658);
nand UO_1695 (O_1695,N_22064,N_22966);
xnor UO_1696 (O_1696,N_20812,N_20868);
nand UO_1697 (O_1697,N_20180,N_24598);
and UO_1698 (O_1698,N_21433,N_23335);
nor UO_1699 (O_1699,N_20724,N_22397);
xor UO_1700 (O_1700,N_22579,N_24004);
or UO_1701 (O_1701,N_21888,N_20577);
and UO_1702 (O_1702,N_22239,N_21523);
nor UO_1703 (O_1703,N_21712,N_21342);
nor UO_1704 (O_1704,N_20273,N_23897);
nor UO_1705 (O_1705,N_22541,N_22912);
and UO_1706 (O_1706,N_20685,N_22599);
xnor UO_1707 (O_1707,N_21519,N_22421);
xnor UO_1708 (O_1708,N_20112,N_24173);
and UO_1709 (O_1709,N_22959,N_24842);
and UO_1710 (O_1710,N_22234,N_24451);
nand UO_1711 (O_1711,N_21560,N_22634);
and UO_1712 (O_1712,N_23368,N_23521);
nor UO_1713 (O_1713,N_23157,N_24546);
nand UO_1714 (O_1714,N_23208,N_22039);
or UO_1715 (O_1715,N_24121,N_21605);
and UO_1716 (O_1716,N_23181,N_20653);
nand UO_1717 (O_1717,N_24793,N_20829);
nor UO_1718 (O_1718,N_21874,N_23013);
and UO_1719 (O_1719,N_23906,N_21474);
or UO_1720 (O_1720,N_24970,N_20770);
or UO_1721 (O_1721,N_21215,N_21672);
and UO_1722 (O_1722,N_22994,N_22272);
nor UO_1723 (O_1723,N_20596,N_24774);
or UO_1724 (O_1724,N_20860,N_20816);
nand UO_1725 (O_1725,N_21901,N_24853);
xnor UO_1726 (O_1726,N_24511,N_22770);
and UO_1727 (O_1727,N_24172,N_21589);
and UO_1728 (O_1728,N_22472,N_22210);
and UO_1729 (O_1729,N_24783,N_20411);
and UO_1730 (O_1730,N_22266,N_22339);
and UO_1731 (O_1731,N_22556,N_24023);
xnor UO_1732 (O_1732,N_21642,N_23125);
nand UO_1733 (O_1733,N_24107,N_21622);
nand UO_1734 (O_1734,N_23405,N_20757);
and UO_1735 (O_1735,N_21795,N_23930);
nor UO_1736 (O_1736,N_24085,N_22601);
nand UO_1737 (O_1737,N_21382,N_24111);
nor UO_1738 (O_1738,N_24687,N_22004);
and UO_1739 (O_1739,N_24960,N_24353);
and UO_1740 (O_1740,N_23080,N_21785);
and UO_1741 (O_1741,N_21197,N_21253);
and UO_1742 (O_1742,N_22196,N_21472);
or UO_1743 (O_1743,N_23343,N_23830);
nand UO_1744 (O_1744,N_23098,N_22101);
nand UO_1745 (O_1745,N_24314,N_24351);
xor UO_1746 (O_1746,N_23360,N_22226);
nand UO_1747 (O_1747,N_24335,N_21392);
nand UO_1748 (O_1748,N_23318,N_23282);
or UO_1749 (O_1749,N_24818,N_24097);
nor UO_1750 (O_1750,N_24750,N_23652);
nand UO_1751 (O_1751,N_20190,N_24926);
and UO_1752 (O_1752,N_22614,N_20688);
and UO_1753 (O_1753,N_20050,N_20578);
or UO_1754 (O_1754,N_21975,N_22655);
nand UO_1755 (O_1755,N_21206,N_23164);
nor UO_1756 (O_1756,N_22936,N_22946);
and UO_1757 (O_1757,N_22026,N_22233);
nor UO_1758 (O_1758,N_20262,N_21267);
or UO_1759 (O_1759,N_20827,N_21045);
or UO_1760 (O_1760,N_21227,N_24077);
nand UO_1761 (O_1761,N_20801,N_22829);
nand UO_1762 (O_1762,N_23420,N_22837);
xnor UO_1763 (O_1763,N_20725,N_21164);
xnor UO_1764 (O_1764,N_22160,N_23599);
or UO_1765 (O_1765,N_22494,N_21140);
nor UO_1766 (O_1766,N_22621,N_22057);
and UO_1767 (O_1767,N_22861,N_23571);
and UO_1768 (O_1768,N_21274,N_21423);
nand UO_1769 (O_1769,N_22778,N_24951);
xor UO_1770 (O_1770,N_20101,N_22607);
and UO_1771 (O_1771,N_21559,N_23473);
nor UO_1772 (O_1772,N_21578,N_21515);
nand UO_1773 (O_1773,N_22592,N_22108);
and UO_1774 (O_1774,N_22971,N_23953);
and UO_1775 (O_1775,N_20950,N_21794);
or UO_1776 (O_1776,N_24569,N_21403);
nand UO_1777 (O_1777,N_20686,N_22754);
or UO_1778 (O_1778,N_23364,N_20662);
nand UO_1779 (O_1779,N_21059,N_20331);
or UO_1780 (O_1780,N_20320,N_21232);
and UO_1781 (O_1781,N_22230,N_24698);
nor UO_1782 (O_1782,N_20221,N_20767);
and UO_1783 (O_1783,N_23815,N_23186);
or UO_1784 (O_1784,N_21191,N_22698);
nand UO_1785 (O_1785,N_21248,N_24149);
or UO_1786 (O_1786,N_20655,N_20434);
xnor UO_1787 (O_1787,N_21949,N_20427);
and UO_1788 (O_1788,N_20082,N_21571);
xnor UO_1789 (O_1789,N_22606,N_20907);
nor UO_1790 (O_1790,N_20391,N_24840);
or UO_1791 (O_1791,N_24070,N_23285);
or UO_1792 (O_1792,N_22129,N_23132);
nor UO_1793 (O_1793,N_21957,N_21961);
nor UO_1794 (O_1794,N_23103,N_22388);
nor UO_1795 (O_1795,N_21952,N_21416);
or UO_1796 (O_1796,N_24276,N_20166);
and UO_1797 (O_1797,N_22567,N_23140);
and UO_1798 (O_1798,N_20621,N_24768);
nor UO_1799 (O_1799,N_23501,N_21012);
nand UO_1800 (O_1800,N_21864,N_20002);
xor UO_1801 (O_1801,N_23408,N_21043);
or UO_1802 (O_1802,N_23942,N_24271);
xor UO_1803 (O_1803,N_21987,N_22212);
nor UO_1804 (O_1804,N_23455,N_21316);
and UO_1805 (O_1805,N_24912,N_23531);
xnor UO_1806 (O_1806,N_23505,N_23008);
nand UO_1807 (O_1807,N_23771,N_21218);
xnor UO_1808 (O_1808,N_22690,N_23442);
xor UO_1809 (O_1809,N_23683,N_21479);
nor UO_1810 (O_1810,N_20751,N_23987);
nand UO_1811 (O_1811,N_23352,N_23938);
xnor UO_1812 (O_1812,N_22080,N_23366);
nand UO_1813 (O_1813,N_20283,N_24790);
or UO_1814 (O_1814,N_20097,N_21154);
or UO_1815 (O_1815,N_20608,N_20136);
or UO_1816 (O_1816,N_22184,N_24940);
and UO_1817 (O_1817,N_21839,N_23454);
and UO_1818 (O_1818,N_21352,N_21738);
or UO_1819 (O_1819,N_22071,N_22611);
or UO_1820 (O_1820,N_23288,N_23415);
or UO_1821 (O_1821,N_20517,N_21436);
or UO_1822 (O_1822,N_24633,N_22926);
nand UO_1823 (O_1823,N_24315,N_23985);
nor UO_1824 (O_1824,N_21386,N_22000);
or UO_1825 (O_1825,N_21529,N_24442);
nor UO_1826 (O_1826,N_22564,N_20527);
nor UO_1827 (O_1827,N_22627,N_23648);
or UO_1828 (O_1828,N_22325,N_20852);
nor UO_1829 (O_1829,N_24886,N_20916);
and UO_1830 (O_1830,N_23030,N_22269);
or UO_1831 (O_1831,N_24082,N_22245);
and UO_1832 (O_1832,N_24125,N_24600);
nand UO_1833 (O_1833,N_23443,N_20539);
xor UO_1834 (O_1834,N_20693,N_21389);
nor UO_1835 (O_1835,N_21259,N_21948);
nand UO_1836 (O_1836,N_24827,N_22009);
or UO_1837 (O_1837,N_20126,N_21024);
and UO_1838 (O_1838,N_22905,N_20998);
nor UO_1839 (O_1839,N_23664,N_20314);
nand UO_1840 (O_1840,N_20678,N_21064);
or UO_1841 (O_1841,N_22699,N_21543);
and UO_1842 (O_1842,N_23145,N_24464);
nand UO_1843 (O_1843,N_22571,N_21171);
or UO_1844 (O_1844,N_23737,N_24537);
or UO_1845 (O_1845,N_21617,N_20567);
nor UO_1846 (O_1846,N_22819,N_22954);
or UO_1847 (O_1847,N_24820,N_24676);
and UO_1848 (O_1848,N_23549,N_20270);
or UO_1849 (O_1849,N_22077,N_22143);
nand UO_1850 (O_1850,N_21967,N_21903);
nor UO_1851 (O_1851,N_23976,N_22540);
and UO_1852 (O_1852,N_20344,N_23572);
or UO_1853 (O_1853,N_21924,N_20514);
nor UO_1854 (O_1854,N_20269,N_20802);
nor UO_1855 (O_1855,N_22373,N_22215);
or UO_1856 (O_1856,N_22107,N_21850);
nor UO_1857 (O_1857,N_23760,N_23467);
nand UO_1858 (O_1858,N_23970,N_20115);
nand UO_1859 (O_1859,N_21510,N_24815);
and UO_1860 (O_1860,N_21599,N_20340);
nor UO_1861 (O_1861,N_20891,N_23320);
nand UO_1862 (O_1862,N_21577,N_24086);
and UO_1863 (O_1863,N_21412,N_22139);
nand UO_1864 (O_1864,N_23483,N_20595);
nor UO_1865 (O_1865,N_21524,N_21620);
nand UO_1866 (O_1866,N_20272,N_20582);
or UO_1867 (O_1867,N_20741,N_23035);
nand UO_1868 (O_1868,N_20904,N_21988);
or UO_1869 (O_1869,N_24736,N_24290);
or UO_1870 (O_1870,N_21587,N_20810);
nor UO_1871 (O_1871,N_21645,N_23260);
nor UO_1872 (O_1872,N_21513,N_23138);
nor UO_1873 (O_1873,N_20120,N_22785);
and UO_1874 (O_1874,N_24156,N_22646);
nand UO_1875 (O_1875,N_24987,N_23112);
and UO_1876 (O_1876,N_20038,N_22929);
and UO_1877 (O_1877,N_22891,N_24185);
xnor UO_1878 (O_1878,N_20274,N_23629);
and UO_1879 (O_1879,N_21567,N_22483);
and UO_1880 (O_1880,N_24931,N_22529);
and UO_1881 (O_1881,N_21295,N_20953);
or UO_1882 (O_1882,N_20942,N_23377);
nor UO_1883 (O_1883,N_20680,N_22464);
or UO_1884 (O_1884,N_24694,N_22265);
or UO_1885 (O_1885,N_20620,N_24823);
and UO_1886 (O_1886,N_24448,N_22284);
or UO_1887 (O_1887,N_22401,N_24438);
or UO_1888 (O_1888,N_22480,N_22955);
nand UO_1889 (O_1889,N_24578,N_24949);
and UO_1890 (O_1890,N_24703,N_22928);
and UO_1891 (O_1891,N_23400,N_20172);
nor UO_1892 (O_1892,N_22884,N_21345);
or UO_1893 (O_1893,N_21068,N_20815);
and UO_1894 (O_1894,N_20749,N_22877);
or UO_1895 (O_1895,N_20563,N_21832);
or UO_1896 (O_1896,N_24656,N_20222);
nand UO_1897 (O_1897,N_24081,N_22165);
nor UO_1898 (O_1898,N_20719,N_21724);
nor UO_1899 (O_1899,N_22093,N_24731);
nand UO_1900 (O_1900,N_24091,N_22359);
or UO_1901 (O_1901,N_22879,N_21627);
nand UO_1902 (O_1902,N_21005,N_24360);
xnor UO_1903 (O_1903,N_20668,N_24414);
nor UO_1904 (O_1904,N_24058,N_20798);
and UO_1905 (O_1905,N_20040,N_21360);
xnor UO_1906 (O_1906,N_20613,N_24681);
or UO_1907 (O_1907,N_21508,N_20327);
or UO_1908 (O_1908,N_22797,N_22478);
xnor UO_1909 (O_1909,N_21100,N_22765);
or UO_1910 (O_1910,N_21530,N_22001);
nand UO_1911 (O_1911,N_22818,N_23220);
nor UO_1912 (O_1912,N_20590,N_24277);
nand UO_1913 (O_1913,N_20267,N_20210);
nor UO_1914 (O_1914,N_24055,N_20955);
and UO_1915 (O_1915,N_22479,N_22683);
or UO_1916 (O_1916,N_24500,N_23267);
nand UO_1917 (O_1917,N_22720,N_24426);
nand UO_1918 (O_1918,N_22362,N_24331);
or UO_1919 (O_1919,N_24654,N_24996);
and UO_1920 (O_1920,N_21008,N_23621);
nand UO_1921 (O_1921,N_21538,N_23697);
nand UO_1922 (O_1922,N_22255,N_22277);
nand UO_1923 (O_1923,N_22896,N_24844);
or UO_1924 (O_1924,N_24803,N_24174);
nand UO_1925 (O_1925,N_22473,N_24101);
and UO_1926 (O_1926,N_22807,N_21800);
nor UO_1927 (O_1927,N_22135,N_21233);
nand UO_1928 (O_1928,N_22358,N_21755);
and UO_1929 (O_1929,N_20876,N_21862);
nor UO_1930 (O_1930,N_24685,N_20471);
nand UO_1931 (O_1931,N_24320,N_21063);
nor UO_1932 (O_1932,N_20387,N_23436);
or UO_1933 (O_1933,N_20791,N_22582);
and UO_1934 (O_1934,N_24642,N_24171);
or UO_1935 (O_1935,N_24686,N_20358);
nor UO_1936 (O_1936,N_22694,N_20498);
xor UO_1937 (O_1937,N_20646,N_21428);
nor UO_1938 (O_1938,N_20461,N_21336);
xor UO_1939 (O_1939,N_23258,N_22553);
or UO_1940 (O_1940,N_24211,N_22799);
or UO_1941 (O_1941,N_23373,N_24343);
or UO_1942 (O_1942,N_20971,N_21744);
and UO_1943 (O_1943,N_24210,N_22987);
or UO_1944 (O_1944,N_21528,N_20650);
or UO_1945 (O_1945,N_22244,N_20508);
and UO_1946 (O_1946,N_23185,N_20765);
or UO_1947 (O_1947,N_20354,N_23246);
nand UO_1948 (O_1948,N_21056,N_22311);
nor UO_1949 (O_1949,N_22605,N_24708);
nor UO_1950 (O_1950,N_22420,N_24001);
or UO_1951 (O_1951,N_21977,N_20500);
xnor UO_1952 (O_1952,N_21561,N_21922);
and UO_1953 (O_1953,N_20778,N_20708);
and UO_1954 (O_1954,N_20306,N_21570);
and UO_1955 (O_1955,N_20856,N_22382);
and UO_1956 (O_1956,N_23876,N_20897);
nand UO_1957 (O_1957,N_20361,N_24398);
nor UO_1958 (O_1958,N_21450,N_24845);
nand UO_1959 (O_1959,N_23696,N_23066);
xnor UO_1960 (O_1960,N_23435,N_22087);
nand UO_1961 (O_1961,N_23289,N_21089);
xnor UO_1962 (O_1962,N_22618,N_23989);
or UO_1963 (O_1963,N_21668,N_22197);
and UO_1964 (O_1964,N_23087,N_20721);
nor UO_1965 (O_1965,N_23314,N_21752);
or UO_1966 (O_1966,N_24340,N_24059);
and UO_1967 (O_1967,N_22848,N_21445);
or UO_1968 (O_1968,N_23023,N_20343);
nor UO_1969 (O_1969,N_22576,N_22530);
nand UO_1970 (O_1970,N_23515,N_23235);
and UO_1971 (O_1971,N_21348,N_24900);
or UO_1972 (O_1972,N_24998,N_21040);
and UO_1973 (O_1973,N_24048,N_22826);
nand UO_1974 (O_1974,N_23895,N_21421);
and UO_1975 (O_1975,N_23886,N_23562);
nor UO_1976 (O_1976,N_24733,N_22545);
or UO_1977 (O_1977,N_20618,N_24336);
or UO_1978 (O_1978,N_23460,N_20619);
xor UO_1979 (O_1979,N_24232,N_20576);
or UO_1980 (O_1980,N_24402,N_20410);
and UO_1981 (O_1981,N_22033,N_20285);
nand UO_1982 (O_1982,N_23229,N_21984);
or UO_1983 (O_1983,N_20857,N_24752);
nand UO_1984 (O_1984,N_22866,N_20187);
nand UO_1985 (O_1985,N_21335,N_24530);
or UO_1986 (O_1986,N_24078,N_20716);
nand UO_1987 (O_1987,N_20661,N_23432);
nand UO_1988 (O_1988,N_22398,N_23949);
nor UO_1989 (O_1989,N_21939,N_20531);
and UO_1990 (O_1990,N_22517,N_23001);
or UO_1991 (O_1991,N_21522,N_24665);
or UO_1992 (O_1992,N_22430,N_20108);
nand UO_1993 (O_1993,N_21683,N_21950);
xnor UO_1994 (O_1994,N_22909,N_24456);
and UO_1995 (O_1995,N_24725,N_20640);
or UO_1996 (O_1996,N_20271,N_22400);
nor UO_1997 (O_1997,N_23661,N_24749);
and UO_1998 (O_1998,N_20936,N_21464);
nor UO_1999 (O_1999,N_20752,N_22500);
nand UO_2000 (O_2000,N_21205,N_21743);
and UO_2001 (O_2001,N_22745,N_21052);
nor UO_2002 (O_2002,N_20010,N_23051);
nand UO_2003 (O_2003,N_23568,N_23564);
nor UO_2004 (O_2004,N_22773,N_24872);
or UO_2005 (O_2005,N_20910,N_21246);
and UO_2006 (O_2006,N_22560,N_23722);
and UO_2007 (O_2007,N_24209,N_21385);
nor UO_2008 (O_2008,N_24423,N_21062);
nand UO_2009 (O_2009,N_23734,N_23502);
nand UO_2010 (O_2010,N_20550,N_24904);
nor UO_2011 (O_2011,N_23773,N_24751);
nand UO_2012 (O_2012,N_21025,N_20887);
xnor UO_2013 (O_2013,N_21694,N_24974);
xor UO_2014 (O_2014,N_20342,N_21239);
and UO_2015 (O_2015,N_22488,N_22155);
and UO_2016 (O_2016,N_20231,N_21158);
and UO_2017 (O_2017,N_22273,N_24054);
nor UO_2018 (O_2018,N_21547,N_23340);
nor UO_2019 (O_2019,N_23838,N_21929);
xor UO_2020 (O_2020,N_20574,N_20246);
and UO_2021 (O_2021,N_20435,N_20584);
nor UO_2022 (O_2022,N_24825,N_22142);
xor UO_2023 (O_2023,N_21773,N_21714);
and UO_2024 (O_2024,N_22095,N_23646);
nand UO_2025 (O_2025,N_22738,N_24966);
nand UO_2026 (O_2026,N_20225,N_20462);
nand UO_2027 (O_2027,N_22449,N_20381);
or UO_2028 (O_2028,N_22872,N_21787);
nand UO_2029 (O_2029,N_22495,N_24455);
and UO_2030 (O_2030,N_24157,N_23644);
and UO_2031 (O_2031,N_23821,N_24930);
and UO_2032 (O_2032,N_24773,N_21860);
nor UO_2033 (O_2033,N_22901,N_24503);
nor UO_2034 (O_2034,N_23931,N_20092);
nand UO_2035 (O_2035,N_20117,N_21820);
xnor UO_2036 (O_2036,N_23213,N_21667);
nand UO_2037 (O_2037,N_23271,N_22995);
nand UO_2038 (O_2038,N_20535,N_23046);
nor UO_2039 (O_2039,N_20626,N_20871);
nor UO_2040 (O_2040,N_23179,N_24071);
nor UO_2041 (O_2041,N_23606,N_23819);
and UO_2042 (O_2042,N_20294,N_24487);
and UO_2043 (O_2043,N_21048,N_24972);
nand UO_2044 (O_2044,N_22643,N_23047);
nor UO_2045 (O_2045,N_21072,N_20754);
nand UO_2046 (O_2046,N_22880,N_23463);
or UO_2047 (O_2047,N_23303,N_22942);
nand UO_2048 (O_2048,N_24093,N_21856);
xnor UO_2049 (O_2049,N_23429,N_20895);
or UO_2050 (O_2050,N_21686,N_22260);
and UO_2051 (O_2051,N_20544,N_23593);
xor UO_2052 (O_2052,N_20091,N_24263);
and UO_2053 (O_2053,N_20872,N_21654);
and UO_2054 (O_2054,N_22732,N_20932);
xor UO_2055 (O_2055,N_23862,N_22574);
nor UO_2056 (O_2056,N_20346,N_23808);
nor UO_2057 (O_2057,N_23687,N_23836);
nor UO_2058 (O_2058,N_21330,N_21138);
or UO_2059 (O_2059,N_23536,N_20102);
nand UO_2060 (O_2060,N_21023,N_20481);
nor UO_2061 (O_2061,N_21757,N_24822);
and UO_2062 (O_2062,N_21226,N_23214);
nand UO_2063 (O_2063,N_23299,N_22386);
and UO_2064 (O_2064,N_23574,N_21823);
nand UO_2065 (O_2065,N_21277,N_20013);
nor UO_2066 (O_2066,N_22558,N_20555);
nor UO_2067 (O_2067,N_21339,N_23272);
nand UO_2068 (O_2068,N_22653,N_23925);
nand UO_2069 (O_2069,N_20063,N_22240);
nor UO_2070 (O_2070,N_22461,N_23619);
and UO_2071 (O_2071,N_23560,N_24292);
nand UO_2072 (O_2072,N_22078,N_20628);
nor UO_2073 (O_2073,N_22340,N_24760);
nand UO_2074 (O_2074,N_20151,N_22570);
nor UO_2075 (O_2075,N_23434,N_20972);
and UO_2076 (O_2076,N_24695,N_23548);
and UO_2077 (O_2077,N_22010,N_23974);
nor UO_2078 (O_2078,N_23555,N_24151);
nor UO_2079 (O_2079,N_23650,N_21468);
nor UO_2080 (O_2080,N_23610,N_22182);
or UO_2081 (O_2081,N_20363,N_24802);
and UO_2082 (O_2082,N_24819,N_22433);
or UO_2083 (O_2083,N_23573,N_24294);
nand UO_2084 (O_2084,N_20885,N_23240);
and UO_2085 (O_2085,N_20874,N_20538);
or UO_2086 (O_2086,N_24240,N_22682);
nand UO_2087 (O_2087,N_20052,N_22159);
nand UO_2088 (O_2088,N_23756,N_21211);
nand UO_2089 (O_2089,N_23481,N_23668);
nand UO_2090 (O_2090,N_23682,N_23437);
nand UO_2091 (O_2091,N_21307,N_23831);
or UO_2092 (O_2092,N_21830,N_22895);
or UO_2093 (O_2093,N_22718,N_21828);
or UO_2094 (O_2094,N_24049,N_22192);
or UO_2095 (O_2095,N_20141,N_21097);
nand UO_2096 (O_2096,N_21147,N_21229);
or UO_2097 (O_2097,N_22346,N_24057);
and UO_2098 (O_2098,N_20370,N_20004);
or UO_2099 (O_2099,N_20249,N_20374);
nor UO_2100 (O_2100,N_23693,N_21180);
nand UO_2101 (O_2101,N_21243,N_20779);
nor UO_2102 (O_2102,N_23743,N_21889);
and UO_2103 (O_2103,N_23591,N_24246);
xnor UO_2104 (O_2104,N_22680,N_24548);
nor UO_2105 (O_2105,N_21804,N_23994);
or UO_2106 (O_2106,N_22916,N_21034);
nand UO_2107 (O_2107,N_23720,N_24990);
and UO_2108 (O_2108,N_22054,N_23276);
nand UO_2109 (O_2109,N_22557,N_22462);
or UO_2110 (O_2110,N_20839,N_20428);
nor UO_2111 (O_2111,N_20682,N_22871);
nor UO_2112 (O_2112,N_24496,N_20338);
nor UO_2113 (O_2113,N_24205,N_21228);
nand UO_2114 (O_2114,N_21306,N_23947);
or UO_2115 (O_2115,N_21554,N_20614);
nand UO_2116 (O_2116,N_23594,N_23851);
nor UO_2117 (O_2117,N_23038,N_21115);
or UO_2118 (O_2118,N_24843,N_22721);
nand UO_2119 (O_2119,N_24231,N_24724);
nor UO_2120 (O_2120,N_20771,N_20324);
or UO_2121 (O_2121,N_23417,N_24494);
or UO_2122 (O_2122,N_20519,N_20762);
nor UO_2123 (O_2123,N_23353,N_21525);
nand UO_2124 (O_2124,N_21287,N_21542);
and UO_2125 (O_2125,N_22894,N_20501);
nor UO_2126 (O_2126,N_24539,N_23091);
or UO_2127 (O_2127,N_21855,N_21321);
or UO_2128 (O_2128,N_24328,N_24384);
nor UO_2129 (O_2129,N_21777,N_24100);
or UO_2130 (O_2130,N_23431,N_21238);
xnor UO_2131 (O_2131,N_24454,N_20322);
nor UO_2132 (O_2132,N_24670,N_24795);
nand UO_2133 (O_2133,N_24268,N_20774);
nand UO_2134 (O_2134,N_21838,N_24306);
nand UO_2135 (O_2135,N_20234,N_23729);
nand UO_2136 (O_2136,N_23472,N_24568);
nand UO_2137 (O_2137,N_22456,N_23695);
or UO_2138 (O_2138,N_20551,N_21976);
nand UO_2139 (O_2139,N_24462,N_23765);
nor UO_2140 (O_2140,N_24199,N_23826);
nand UO_2141 (O_2141,N_21017,N_22467);
or UO_2142 (O_2142,N_20755,N_20131);
and UO_2143 (O_2143,N_20375,N_22391);
nand UO_2144 (O_2144,N_21364,N_23554);
and UO_2145 (O_2145,N_21912,N_22609);
and UO_2146 (O_2146,N_23916,N_21847);
or UO_2147 (O_2147,N_21716,N_22264);
nor UO_2148 (O_2148,N_24003,N_20821);
and UO_2149 (O_2149,N_21088,N_22195);
nor UO_2150 (O_2150,N_21811,N_20448);
and UO_2151 (O_2151,N_21928,N_20323);
and UO_2152 (O_2152,N_23984,N_22378);
or UO_2153 (O_2153,N_20822,N_22783);
xor UO_2154 (O_2154,N_24547,N_24027);
or UO_2155 (O_2155,N_24920,N_23438);
and UO_2156 (O_2156,N_24465,N_24347);
or UO_2157 (O_2157,N_22122,N_21527);
and UO_2158 (O_2158,N_24408,N_23317);
or UO_2159 (O_2159,N_24167,N_21441);
or UO_2160 (O_2160,N_21867,N_21288);
or UO_2161 (O_2161,N_21633,N_24346);
and UO_2162 (O_2162,N_21254,N_21934);
nor UO_2163 (O_2163,N_24927,N_23308);
xnor UO_2164 (O_2164,N_23849,N_21430);
and UO_2165 (O_2165,N_24918,N_23585);
or UO_2166 (O_2166,N_21347,N_21644);
nand UO_2167 (O_2167,N_23310,N_24038);
and UO_2168 (O_2168,N_20217,N_20412);
and UO_2169 (O_2169,N_22578,N_24355);
xor UO_2170 (O_2170,N_23710,N_24730);
xnor UO_2171 (O_2171,N_21141,N_24992);
and UO_2172 (O_2172,N_22085,N_21046);
nand UO_2173 (O_2173,N_23709,N_22123);
xor UO_2174 (O_2174,N_20518,N_24217);
nor UO_2175 (O_2175,N_23166,N_21486);
nor UO_2176 (O_2176,N_24852,N_24135);
nor UO_2177 (O_2177,N_23889,N_22216);
nor UO_2178 (O_2178,N_23855,N_24728);
nor UO_2179 (O_2179,N_23333,N_22505);
nor UO_2180 (O_2180,N_24639,N_20083);
or UO_2181 (O_2181,N_20143,N_22812);
and UO_2182 (O_2182,N_21462,N_23257);
nand UO_2183 (O_2183,N_23062,N_24935);
and UO_2184 (O_2184,N_20109,N_21373);
nor UO_2185 (O_2185,N_23888,N_24165);
nand UO_2186 (O_2186,N_24583,N_22798);
or UO_2187 (O_2187,N_20302,N_23890);
nor UO_2188 (O_2188,N_22962,N_22843);
nor UO_2189 (O_2189,N_24769,N_24899);
nor UO_2190 (O_2190,N_22625,N_22997);
and UO_2191 (O_2191,N_20066,N_22787);
nor UO_2192 (O_2192,N_20610,N_24196);
or UO_2193 (O_2193,N_23342,N_22207);
nand UO_2194 (O_2194,N_24564,N_24181);
and UO_2195 (O_2195,N_24610,N_24592);
or UO_2196 (O_2196,N_23439,N_20300);
or UO_2197 (O_2197,N_23109,N_23356);
or UO_2198 (O_2198,N_23757,N_23144);
and UO_2199 (O_2199,N_20206,N_23739);
nor UO_2200 (O_2200,N_23708,N_23471);
nor UO_2201 (O_2201,N_24417,N_23491);
and UO_2202 (O_2202,N_23782,N_23331);
nor UO_2203 (O_2203,N_21802,N_22131);
xor UO_2204 (O_2204,N_21849,N_21954);
nand UO_2205 (O_2205,N_22383,N_21160);
nand UO_2206 (O_2206,N_21956,N_20804);
and UO_2207 (O_2207,N_22070,N_24898);
nor UO_2208 (O_2208,N_20232,N_22666);
nor UO_2209 (O_2209,N_22334,N_21603);
nand UO_2210 (O_2210,N_20007,N_20384);
nand UO_2211 (O_2211,N_21799,N_24737);
nand UO_2212 (O_2212,N_22440,N_23241);
or UO_2213 (O_2213,N_20149,N_22043);
nand UO_2214 (O_2214,N_22645,N_20186);
or UO_2215 (O_2215,N_22911,N_23010);
or UO_2216 (O_2216,N_20795,N_20239);
or UO_2217 (O_2217,N_24780,N_23827);
nand UO_2218 (O_2218,N_22432,N_24602);
nor UO_2219 (O_2219,N_24764,N_21111);
nand UO_2220 (O_2220,N_24405,N_21476);
nor UO_2221 (O_2221,N_24788,N_22091);
and UO_2222 (O_2222,N_22170,N_20609);
or UO_2223 (O_2223,N_22784,N_21822);
or UO_2224 (O_2224,N_22800,N_21037);
and UO_2225 (O_2225,N_24950,N_21325);
and UO_2226 (O_2226,N_24933,N_24046);
nor UO_2227 (O_2227,N_21619,N_23301);
or UO_2228 (O_2228,N_21276,N_20240);
and UO_2229 (O_2229,N_20450,N_21594);
nor UO_2230 (O_2230,N_24851,N_24471);
nor UO_2231 (O_2231,N_24123,N_20947);
and UO_2232 (O_2232,N_20738,N_22504);
nor UO_2233 (O_2233,N_24193,N_20870);
xor UO_2234 (O_2234,N_24868,N_22407);
xor UO_2235 (O_2235,N_21272,N_22511);
nand UO_2236 (O_2236,N_24234,N_22580);
xor UO_2237 (O_2237,N_23582,N_24316);
and UO_2238 (O_2238,N_20985,N_20263);
and UO_2239 (O_2239,N_22013,N_21652);
nor UO_2240 (O_2240,N_21556,N_24717);
nor UO_2241 (O_2241,N_22235,N_21938);
and UO_2242 (O_2242,N_21626,N_21110);
nand UO_2243 (O_2243,N_21128,N_21615);
nor UO_2244 (O_2244,N_22693,N_20641);
xnor UO_2245 (O_2245,N_22739,N_23997);
nor UO_2246 (O_2246,N_23210,N_20030);
and UO_2247 (O_2247,N_21478,N_24635);
and UO_2248 (O_2248,N_23915,N_20321);
nand UO_2249 (O_2249,N_23822,N_23486);
nor UO_2250 (O_2250,N_20848,N_24779);
or UO_2251 (O_2251,N_23804,N_20487);
and UO_2252 (O_2252,N_21943,N_22424);
and UO_2253 (O_2253,N_20341,N_23090);
nor UO_2254 (O_2254,N_24572,N_22547);
nand UO_2255 (O_2255,N_22148,N_23614);
xnor UO_2256 (O_2256,N_24714,N_20575);
nor UO_2257 (O_2257,N_21512,N_24469);
or UO_2258 (O_2258,N_21042,N_20783);
nor UO_2259 (O_2259,N_21698,N_23504);
nor UO_2260 (O_2260,N_20015,N_20624);
nand UO_2261 (O_2261,N_23767,N_20781);
or UO_2262 (O_2262,N_22422,N_22179);
or UO_2263 (O_2263,N_24636,N_21168);
xnor UO_2264 (O_2264,N_21959,N_21963);
nand UO_2265 (O_2265,N_23857,N_24118);
nor UO_2266 (O_2266,N_21395,N_22939);
nand UO_2267 (O_2267,N_23937,N_20598);
and UO_2268 (O_2268,N_20666,N_21595);
xor UO_2269 (O_2269,N_20395,N_21182);
or UO_2270 (O_2270,N_22842,N_21514);
or UO_2271 (O_2271,N_20750,N_20207);
or UO_2272 (O_2272,N_23514,N_20479);
and UO_2273 (O_2273,N_24800,N_22510);
nor UO_2274 (O_2274,N_24571,N_21737);
or UO_2275 (O_2275,N_24035,N_22451);
nand UO_2276 (O_2276,N_24410,N_24421);
or UO_2277 (O_2277,N_22238,N_21651);
nor UO_2278 (O_2278,N_23556,N_23839);
and UO_2279 (O_2279,N_22988,N_23268);
and UO_2280 (O_2280,N_23503,N_20507);
and UO_2281 (O_2281,N_21333,N_21075);
and UO_2282 (O_2282,N_24605,N_20414);
nor UO_2283 (O_2283,N_21751,N_23369);
nand UO_2284 (O_2284,N_24429,N_24050);
or UO_2285 (O_2285,N_22408,N_20405);
nand UO_2286 (O_2286,N_21728,N_24104);
xor UO_2287 (O_2287,N_24747,N_20076);
xnor UO_2288 (O_2288,N_21372,N_21125);
nor UO_2289 (O_2289,N_24237,N_21545);
xnor UO_2290 (O_2290,N_20836,N_20357);
nand UO_2291 (O_2291,N_21310,N_23913);
nand UO_2292 (O_2292,N_24391,N_21951);
nor UO_2293 (O_2293,N_23174,N_24338);
nand UO_2294 (O_2294,N_24893,N_24660);
nand UO_2295 (O_2295,N_23647,N_23604);
or UO_2296 (O_2296,N_20229,N_22471);
nand UO_2297 (O_2297,N_22484,N_21548);
nor UO_2298 (O_2298,N_23617,N_23701);
and UO_2299 (O_2299,N_22730,N_21861);
nor UO_2300 (O_2300,N_23034,N_21628);
xor UO_2301 (O_2301,N_21044,N_24376);
nand UO_2302 (O_2302,N_21129,N_22247);
nor UO_2303 (O_2303,N_22253,N_22713);
xnor UO_2304 (O_2304,N_23261,N_21781);
nor UO_2305 (O_2305,N_22310,N_23456);
or UO_2306 (O_2306,N_23592,N_24946);
nor UO_2307 (O_2307,N_24254,N_24613);
and UO_2308 (O_2308,N_22711,N_20071);
nor UO_2309 (O_2309,N_20740,N_20244);
and UO_2310 (O_2310,N_23772,N_22246);
and UO_2311 (O_2311,N_23602,N_24404);
and UO_2312 (O_2312,N_23842,N_20406);
nand UO_2313 (O_2313,N_23894,N_24806);
xor UO_2314 (O_2314,N_20430,N_23150);
nand UO_2315 (O_2315,N_22704,N_21721);
and UO_2316 (O_2316,N_21782,N_24208);
nor UO_2317 (O_2317,N_22002,N_20194);
nand UO_2318 (O_2318,N_24365,N_23846);
or UO_2319 (O_2319,N_23832,N_22524);
nor UO_2320 (O_2320,N_20766,N_20193);
and UO_2321 (O_2321,N_24136,N_20139);
and UO_2322 (O_2322,N_20077,N_20335);
and UO_2323 (O_2323,N_22209,N_22283);
nor UO_2324 (O_2324,N_20472,N_20861);
or UO_2325 (O_2325,N_24356,N_24874);
nor UO_2326 (O_2326,N_24597,N_23887);
and UO_2327 (O_2327,N_21247,N_24120);
nor UO_2328 (O_2328,N_22586,N_23799);
xor UO_2329 (O_2329,N_24293,N_21156);
or UO_2330 (O_2330,N_22887,N_24828);
nand UO_2331 (O_2331,N_20032,N_20099);
nand UO_2332 (O_2332,N_21843,N_20697);
xor UO_2333 (O_2333,N_20833,N_22106);
and UO_2334 (O_2334,N_23990,N_20516);
nand UO_2335 (O_2335,N_24226,N_22144);
or UO_2336 (O_2336,N_21092,N_21703);
nor UO_2337 (O_2337,N_22526,N_24709);
and UO_2338 (O_2338,N_23263,N_23148);
xnor UO_2339 (O_2339,N_22084,N_20718);
nand UO_2340 (O_2340,N_21203,N_23758);
and UO_2341 (O_2341,N_20756,N_23061);
or UO_2342 (O_2342,N_24979,N_23911);
nor UO_2343 (O_2343,N_21497,N_23067);
nor UO_2344 (O_2344,N_23475,N_23580);
nor UO_2345 (O_2345,N_22428,N_20911);
and UO_2346 (O_2346,N_20540,N_22134);
nor UO_2347 (O_2347,N_24666,N_21371);
and UO_2348 (O_2348,N_22393,N_23026);
or UO_2349 (O_2349,N_24447,N_23201);
and UO_2350 (O_2350,N_24434,N_23349);
or UO_2351 (O_2351,N_24657,N_20996);
or UO_2352 (O_2352,N_23402,N_23690);
nand UO_2353 (O_2353,N_21658,N_24270);
nor UO_2354 (O_2354,N_22658,N_21118);
nand UO_2355 (O_2355,N_23651,N_23316);
xor UO_2356 (O_2356,N_20392,N_21491);
nor UO_2357 (O_2357,N_23231,N_23292);
nand UO_2358 (O_2358,N_21872,N_24984);
nor UO_2359 (O_2359,N_22193,N_22438);
or UO_2360 (O_2360,N_20714,N_24830);
or UO_2361 (O_2361,N_22353,N_20603);
or UO_2362 (O_2362,N_24587,N_20920);
or UO_2363 (O_2363,N_24304,N_20475);
and UO_2364 (O_2364,N_22999,N_20503);
nor UO_2365 (O_2365,N_21925,N_20027);
nor UO_2366 (O_2366,N_21323,N_22414);
xnor UO_2367 (O_2367,N_24501,N_23901);
nor UO_2368 (O_2368,N_21261,N_24109);
xor UO_2369 (O_2369,N_22550,N_21982);
xnor UO_2370 (O_2370,N_22722,N_21188);
or UO_2371 (O_2371,N_20185,N_24092);
nand UO_2372 (O_2372,N_23095,N_21793);
xnor UO_2373 (O_2373,N_22206,N_24311);
and UO_2374 (O_2374,N_22457,N_20332);
or UO_2375 (O_2375,N_23108,N_20276);
and UO_2376 (O_2376,N_22227,N_23224);
and UO_2377 (O_2377,N_23595,N_24273);
xnor UO_2378 (O_2378,N_23076,N_22068);
nor UO_2379 (O_2379,N_21127,N_24968);
or UO_2380 (O_2380,N_20457,N_24936);
xor UO_2381 (O_2381,N_24220,N_21369);
or UO_2382 (O_2382,N_22669,N_24018);
nor UO_2383 (O_2383,N_21825,N_21535);
nand UO_2384 (O_2384,N_24504,N_21356);
or UO_2385 (O_2385,N_24068,N_20788);
and UO_2386 (O_2386,N_22387,N_20389);
nor UO_2387 (O_2387,N_22204,N_22667);
nand UO_2388 (O_2388,N_23959,N_24288);
xnor UO_2389 (O_2389,N_24555,N_24260);
and UO_2390 (O_2390,N_23187,N_22923);
or UO_2391 (O_2391,N_20116,N_21234);
and UO_2392 (O_2392,N_21066,N_23800);
nor UO_2393 (O_2393,N_24436,N_20245);
nor UO_2394 (O_2394,N_23717,N_20505);
nand UO_2395 (O_2395,N_23498,N_20736);
nand UO_2396 (O_2396,N_24069,N_21898);
and UO_2397 (O_2397,N_23237,N_23685);
or UO_2398 (O_2398,N_20796,N_24742);
nor UO_2399 (O_2399,N_22465,N_23474);
or UO_2400 (O_2400,N_22945,N_21296);
nor UO_2401 (O_2401,N_21916,N_22117);
nor UO_2402 (O_2402,N_22965,N_24528);
or UO_2403 (O_2403,N_21116,N_20759);
and UO_2404 (O_2404,N_23854,N_20168);
nor UO_2405 (O_2405,N_21859,N_22138);
and UO_2406 (O_2406,N_20571,N_20722);
and UO_2407 (O_2407,N_22838,N_20663);
xor UO_2408 (O_2408,N_23326,N_23131);
nor UO_2409 (O_2409,N_20878,N_24313);
and UO_2410 (O_2410,N_24419,N_23409);
nor UO_2411 (O_2411,N_23705,N_20701);
nand UO_2412 (O_2412,N_23332,N_23141);
or UO_2413 (O_2413,N_24961,N_21553);
or UO_2414 (O_2414,N_22231,N_20057);
and UO_2415 (O_2415,N_20880,N_21501);
nor UO_2416 (O_2416,N_21362,N_24640);
xnor UO_2417 (O_2417,N_21083,N_21447);
or UO_2418 (O_2418,N_21242,N_21405);
or UO_2419 (O_2419,N_21660,N_23977);
nor UO_2420 (O_2420,N_23907,N_23569);
nand UO_2421 (O_2421,N_22642,N_20636);
or UO_2422 (O_2422,N_24076,N_23152);
or UO_2423 (O_2423,N_22169,N_21090);
or UO_2424 (O_2424,N_23654,N_20293);
or UO_2425 (O_2425,N_20385,N_20080);
and UO_2426 (O_2426,N_23130,N_23880);
nand UO_2427 (O_2427,N_23598,N_22147);
and UO_2428 (O_2428,N_21150,N_20105);
nand UO_2429 (O_2429,N_22796,N_21235);
nor UO_2430 (O_2430,N_23054,N_22846);
nor UO_2431 (O_2431,N_21848,N_23093);
and UO_2432 (O_2432,N_23609,N_24043);
or UO_2433 (O_2433,N_20828,N_21355);
xor UO_2434 (O_2434,N_20253,N_24492);
or UO_2435 (O_2435,N_20183,N_22156);
xor UO_2436 (O_2436,N_22596,N_22276);
nor UO_2437 (O_2437,N_20449,N_21026);
or UO_2438 (O_2438,N_22620,N_22709);
nand UO_2439 (O_2439,N_23996,N_23256);
nor UO_2440 (O_2440,N_21641,N_21854);
or UO_2441 (O_2441,N_23037,N_23088);
nand UO_2442 (O_2442,N_21878,N_24284);
nor UO_2443 (O_2443,N_24235,N_21753);
nand UO_2444 (O_2444,N_23461,N_23774);
xnor UO_2445 (O_2445,N_20568,N_23251);
nand UO_2446 (O_2446,N_21673,N_22347);
nor UO_2447 (O_2447,N_22023,N_24720);
xnor UO_2448 (O_2448,N_23111,N_23418);
nor UO_2449 (O_2449,N_21745,N_22178);
or UO_2450 (O_2450,N_21194,N_24375);
and UO_2451 (O_2451,N_20295,N_24032);
and UO_2452 (O_2452,N_23468,N_20008);
nor UO_2453 (O_2453,N_24856,N_21196);
or UO_2454 (O_2454,N_24251,N_24575);
or UO_2455 (O_2455,N_22977,N_24841);
or UO_2456 (O_2456,N_24616,N_22963);
nor UO_2457 (O_2457,N_23389,N_22038);
and UO_2458 (O_2458,N_24140,N_22925);
and UO_2459 (O_2459,N_24257,N_23253);
and UO_2460 (O_2460,N_22779,N_23307);
nor UO_2461 (O_2461,N_20256,N_21858);
and UO_2462 (O_2462,N_22774,N_24468);
or UO_2463 (O_2463,N_24658,N_24611);
nand UO_2464 (O_2464,N_21370,N_20964);
or UO_2465 (O_2465,N_24067,N_21039);
nor UO_2466 (O_2466,N_20960,N_24858);
or UO_2467 (O_2467,N_23499,N_21172);
or UO_2468 (O_2468,N_20104,N_22112);
nand UO_2469 (O_2469,N_23653,N_24388);
nand UO_2470 (O_2470,N_21028,N_20863);
xor UO_2471 (O_2471,N_21475,N_22600);
nand UO_2472 (O_2472,N_23630,N_21463);
xor UO_2473 (O_2473,N_23173,N_24339);
nor UO_2474 (O_2474,N_21377,N_23748);
nand UO_2475 (O_2475,N_23339,N_23269);
or UO_2476 (O_2476,N_22544,N_23623);
or UO_2477 (O_2477,N_20110,N_20499);
nor UO_2478 (O_2478,N_21490,N_23032);
or UO_2479 (O_2479,N_24476,N_21945);
xor UO_2480 (O_2480,N_23165,N_24357);
or UO_2481 (O_2481,N_23348,N_21727);
nand UO_2482 (O_2482,N_21281,N_20753);
or UO_2483 (O_2483,N_24669,N_21041);
xnor UO_2484 (O_2484,N_23011,N_21170);
nor UO_2485 (O_2485,N_24102,N_24490);
xor UO_2486 (O_2486,N_20869,N_21251);
or UO_2487 (O_2487,N_20676,N_21219);
nand UO_2488 (O_2488,N_24707,N_20045);
and UO_2489 (O_2489,N_21429,N_22256);
nand UO_2490 (O_2490,N_24090,N_22150);
nor UO_2491 (O_2491,N_22130,N_24896);
xor UO_2492 (O_2492,N_23791,N_22506);
or UO_2493 (O_2493,N_23563,N_24740);
xnor UO_2494 (O_2494,N_24106,N_21461);
or UO_2495 (O_2495,N_22650,N_23575);
nor UO_2496 (O_2496,N_22985,N_23134);
xor UO_2497 (O_2497,N_22174,N_22366);
nor UO_2498 (O_2498,N_20651,N_21887);
nand UO_2499 (O_2499,N_24762,N_22632);
nor UO_2500 (O_2500,N_21045,N_24360);
or UO_2501 (O_2501,N_24490,N_24711);
xnor UO_2502 (O_2502,N_22009,N_22828);
nor UO_2503 (O_2503,N_23315,N_24789);
or UO_2504 (O_2504,N_24795,N_22752);
nand UO_2505 (O_2505,N_23499,N_21236);
nor UO_2506 (O_2506,N_23998,N_23060);
and UO_2507 (O_2507,N_20413,N_21462);
nor UO_2508 (O_2508,N_24767,N_20912);
nor UO_2509 (O_2509,N_20159,N_22824);
xor UO_2510 (O_2510,N_22068,N_21506);
nand UO_2511 (O_2511,N_24245,N_20036);
and UO_2512 (O_2512,N_24726,N_24873);
nand UO_2513 (O_2513,N_20998,N_24480);
nor UO_2514 (O_2514,N_20482,N_21950);
and UO_2515 (O_2515,N_24424,N_21187);
or UO_2516 (O_2516,N_21044,N_22896);
nor UO_2517 (O_2517,N_21743,N_21283);
xor UO_2518 (O_2518,N_22595,N_20424);
or UO_2519 (O_2519,N_20310,N_23330);
xor UO_2520 (O_2520,N_22325,N_23610);
nand UO_2521 (O_2521,N_23832,N_23781);
and UO_2522 (O_2522,N_22963,N_23432);
and UO_2523 (O_2523,N_20394,N_21571);
or UO_2524 (O_2524,N_23911,N_23443);
xnor UO_2525 (O_2525,N_24210,N_24328);
nand UO_2526 (O_2526,N_20559,N_21716);
nand UO_2527 (O_2527,N_24137,N_23736);
nor UO_2528 (O_2528,N_24891,N_20896);
or UO_2529 (O_2529,N_20119,N_22500);
nand UO_2530 (O_2530,N_20599,N_23588);
and UO_2531 (O_2531,N_21946,N_22965);
nand UO_2532 (O_2532,N_22467,N_20665);
and UO_2533 (O_2533,N_21951,N_21129);
or UO_2534 (O_2534,N_20591,N_21669);
and UO_2535 (O_2535,N_23936,N_20261);
nor UO_2536 (O_2536,N_22928,N_23633);
and UO_2537 (O_2537,N_22505,N_23022);
or UO_2538 (O_2538,N_23446,N_21611);
xor UO_2539 (O_2539,N_21212,N_21660);
nor UO_2540 (O_2540,N_20926,N_23625);
xor UO_2541 (O_2541,N_22080,N_20351);
nor UO_2542 (O_2542,N_20717,N_21362);
xnor UO_2543 (O_2543,N_22386,N_21323);
nor UO_2544 (O_2544,N_20597,N_24244);
nand UO_2545 (O_2545,N_23703,N_21867);
and UO_2546 (O_2546,N_23590,N_22654);
nand UO_2547 (O_2547,N_20685,N_20170);
nand UO_2548 (O_2548,N_21808,N_20727);
and UO_2549 (O_2549,N_23362,N_24316);
or UO_2550 (O_2550,N_22073,N_22692);
nor UO_2551 (O_2551,N_21700,N_22032);
xnor UO_2552 (O_2552,N_21716,N_23371);
xor UO_2553 (O_2553,N_22505,N_22378);
nand UO_2554 (O_2554,N_21792,N_24298);
nor UO_2555 (O_2555,N_20267,N_24145);
nor UO_2556 (O_2556,N_22120,N_20670);
and UO_2557 (O_2557,N_20771,N_20172);
nor UO_2558 (O_2558,N_24256,N_22148);
xnor UO_2559 (O_2559,N_22846,N_24590);
nand UO_2560 (O_2560,N_20727,N_21696);
nand UO_2561 (O_2561,N_21506,N_21651);
or UO_2562 (O_2562,N_22772,N_21037);
nor UO_2563 (O_2563,N_24084,N_21171);
nand UO_2564 (O_2564,N_23057,N_22434);
nor UO_2565 (O_2565,N_24336,N_23549);
or UO_2566 (O_2566,N_21540,N_23329);
nor UO_2567 (O_2567,N_20309,N_22112);
and UO_2568 (O_2568,N_23556,N_20465);
nor UO_2569 (O_2569,N_23332,N_23463);
and UO_2570 (O_2570,N_23624,N_21083);
and UO_2571 (O_2571,N_20699,N_23200);
and UO_2572 (O_2572,N_23813,N_22726);
and UO_2573 (O_2573,N_21782,N_22040);
and UO_2574 (O_2574,N_24701,N_24190);
or UO_2575 (O_2575,N_22357,N_20358);
and UO_2576 (O_2576,N_23210,N_21756);
or UO_2577 (O_2577,N_22196,N_23415);
or UO_2578 (O_2578,N_23810,N_22837);
nand UO_2579 (O_2579,N_22082,N_24341);
and UO_2580 (O_2580,N_24769,N_22659);
nand UO_2581 (O_2581,N_20991,N_23699);
nor UO_2582 (O_2582,N_24944,N_22669);
or UO_2583 (O_2583,N_24536,N_22452);
nor UO_2584 (O_2584,N_21923,N_24662);
nand UO_2585 (O_2585,N_20903,N_23878);
nor UO_2586 (O_2586,N_23743,N_21260);
nand UO_2587 (O_2587,N_22563,N_20903);
and UO_2588 (O_2588,N_24189,N_21462);
or UO_2589 (O_2589,N_20570,N_23511);
or UO_2590 (O_2590,N_21518,N_24161);
nand UO_2591 (O_2591,N_23143,N_22201);
or UO_2592 (O_2592,N_21672,N_22610);
or UO_2593 (O_2593,N_24313,N_23534);
and UO_2594 (O_2594,N_24797,N_22253);
or UO_2595 (O_2595,N_21213,N_23904);
nor UO_2596 (O_2596,N_22939,N_22434);
nor UO_2597 (O_2597,N_20747,N_23041);
or UO_2598 (O_2598,N_24591,N_23937);
and UO_2599 (O_2599,N_21850,N_22787);
nor UO_2600 (O_2600,N_21731,N_24872);
nand UO_2601 (O_2601,N_20642,N_24038);
or UO_2602 (O_2602,N_24103,N_21674);
and UO_2603 (O_2603,N_21946,N_22135);
nor UO_2604 (O_2604,N_21635,N_24119);
or UO_2605 (O_2605,N_23258,N_24625);
nor UO_2606 (O_2606,N_24370,N_20786);
or UO_2607 (O_2607,N_20899,N_20841);
nor UO_2608 (O_2608,N_23136,N_22183);
nor UO_2609 (O_2609,N_23274,N_24544);
and UO_2610 (O_2610,N_24225,N_24878);
nand UO_2611 (O_2611,N_24811,N_23492);
and UO_2612 (O_2612,N_20390,N_22117);
or UO_2613 (O_2613,N_21198,N_22624);
nor UO_2614 (O_2614,N_21957,N_23491);
or UO_2615 (O_2615,N_21327,N_22625);
xor UO_2616 (O_2616,N_20018,N_22815);
nor UO_2617 (O_2617,N_23091,N_24049);
nand UO_2618 (O_2618,N_23679,N_24910);
xor UO_2619 (O_2619,N_23040,N_20447);
and UO_2620 (O_2620,N_24677,N_21162);
nor UO_2621 (O_2621,N_22902,N_24054);
nand UO_2622 (O_2622,N_21886,N_24939);
nor UO_2623 (O_2623,N_20698,N_24112);
nor UO_2624 (O_2624,N_22764,N_22029);
nor UO_2625 (O_2625,N_22083,N_20886);
and UO_2626 (O_2626,N_23867,N_21173);
xor UO_2627 (O_2627,N_23454,N_21285);
nand UO_2628 (O_2628,N_22083,N_23094);
nor UO_2629 (O_2629,N_24636,N_23432);
nand UO_2630 (O_2630,N_22858,N_21445);
or UO_2631 (O_2631,N_23943,N_21077);
and UO_2632 (O_2632,N_24821,N_23694);
nor UO_2633 (O_2633,N_23304,N_21143);
nor UO_2634 (O_2634,N_22075,N_22756);
nand UO_2635 (O_2635,N_21082,N_24737);
or UO_2636 (O_2636,N_20795,N_23484);
nor UO_2637 (O_2637,N_20380,N_23282);
nor UO_2638 (O_2638,N_20518,N_24657);
and UO_2639 (O_2639,N_20531,N_22633);
or UO_2640 (O_2640,N_21574,N_23512);
nand UO_2641 (O_2641,N_21975,N_21247);
and UO_2642 (O_2642,N_21894,N_23591);
and UO_2643 (O_2643,N_21937,N_22066);
or UO_2644 (O_2644,N_20760,N_20694);
xor UO_2645 (O_2645,N_24364,N_24053);
nand UO_2646 (O_2646,N_20705,N_21652);
or UO_2647 (O_2647,N_23971,N_24423);
nor UO_2648 (O_2648,N_23763,N_20752);
or UO_2649 (O_2649,N_23223,N_20880);
or UO_2650 (O_2650,N_24491,N_22789);
nor UO_2651 (O_2651,N_22477,N_20027);
nand UO_2652 (O_2652,N_21843,N_21796);
nand UO_2653 (O_2653,N_22988,N_22366);
nand UO_2654 (O_2654,N_22606,N_23059);
or UO_2655 (O_2655,N_24887,N_21473);
or UO_2656 (O_2656,N_23339,N_22024);
and UO_2657 (O_2657,N_23143,N_23560);
nor UO_2658 (O_2658,N_21466,N_24172);
or UO_2659 (O_2659,N_23175,N_21987);
or UO_2660 (O_2660,N_22049,N_20825);
or UO_2661 (O_2661,N_20740,N_21405);
or UO_2662 (O_2662,N_20947,N_23922);
and UO_2663 (O_2663,N_21439,N_20005);
and UO_2664 (O_2664,N_23660,N_22538);
or UO_2665 (O_2665,N_23110,N_20873);
nor UO_2666 (O_2666,N_22922,N_24057);
nand UO_2667 (O_2667,N_21804,N_22560);
nand UO_2668 (O_2668,N_20034,N_23238);
and UO_2669 (O_2669,N_20236,N_21211);
nor UO_2670 (O_2670,N_21849,N_21197);
xor UO_2671 (O_2671,N_24241,N_21011);
nand UO_2672 (O_2672,N_22707,N_23676);
xnor UO_2673 (O_2673,N_21965,N_24727);
nand UO_2674 (O_2674,N_21849,N_24302);
and UO_2675 (O_2675,N_21958,N_20216);
nor UO_2676 (O_2676,N_23099,N_24191);
nand UO_2677 (O_2677,N_24528,N_23893);
nand UO_2678 (O_2678,N_21864,N_22343);
or UO_2679 (O_2679,N_24921,N_22938);
or UO_2680 (O_2680,N_22071,N_20197);
and UO_2681 (O_2681,N_22279,N_20561);
nor UO_2682 (O_2682,N_23776,N_22813);
xor UO_2683 (O_2683,N_23109,N_22809);
xor UO_2684 (O_2684,N_20276,N_24215);
xnor UO_2685 (O_2685,N_20317,N_21736);
xor UO_2686 (O_2686,N_22604,N_24306);
nor UO_2687 (O_2687,N_20414,N_22668);
and UO_2688 (O_2688,N_21640,N_24791);
and UO_2689 (O_2689,N_20543,N_23101);
nor UO_2690 (O_2690,N_22607,N_24179);
and UO_2691 (O_2691,N_21456,N_22214);
xnor UO_2692 (O_2692,N_23287,N_23187);
nand UO_2693 (O_2693,N_24210,N_21317);
xor UO_2694 (O_2694,N_23861,N_22967);
nor UO_2695 (O_2695,N_23523,N_21033);
nor UO_2696 (O_2696,N_23099,N_21798);
nand UO_2697 (O_2697,N_20959,N_24306);
and UO_2698 (O_2698,N_24902,N_20390);
nand UO_2699 (O_2699,N_24497,N_23789);
nand UO_2700 (O_2700,N_21141,N_23289);
nor UO_2701 (O_2701,N_24800,N_20865);
or UO_2702 (O_2702,N_24433,N_20327);
and UO_2703 (O_2703,N_24387,N_21926);
or UO_2704 (O_2704,N_24771,N_24610);
nand UO_2705 (O_2705,N_20738,N_22995);
nand UO_2706 (O_2706,N_23937,N_23174);
and UO_2707 (O_2707,N_22459,N_21958);
or UO_2708 (O_2708,N_22074,N_22232);
nor UO_2709 (O_2709,N_23760,N_24652);
or UO_2710 (O_2710,N_24242,N_24050);
or UO_2711 (O_2711,N_20125,N_23422);
nand UO_2712 (O_2712,N_20065,N_24876);
xor UO_2713 (O_2713,N_20271,N_23743);
xor UO_2714 (O_2714,N_20955,N_21152);
nor UO_2715 (O_2715,N_21226,N_23108);
and UO_2716 (O_2716,N_24889,N_22576);
and UO_2717 (O_2717,N_21524,N_22108);
xnor UO_2718 (O_2718,N_20134,N_22093);
nand UO_2719 (O_2719,N_23241,N_22105);
nand UO_2720 (O_2720,N_22018,N_22455);
nand UO_2721 (O_2721,N_21654,N_24554);
nor UO_2722 (O_2722,N_22262,N_20599);
nand UO_2723 (O_2723,N_22540,N_24939);
and UO_2724 (O_2724,N_24128,N_20744);
nand UO_2725 (O_2725,N_22315,N_24851);
nor UO_2726 (O_2726,N_21488,N_21896);
xnor UO_2727 (O_2727,N_22414,N_20315);
and UO_2728 (O_2728,N_21238,N_21026);
nor UO_2729 (O_2729,N_23788,N_24960);
or UO_2730 (O_2730,N_24044,N_21332);
nor UO_2731 (O_2731,N_21566,N_24535);
nand UO_2732 (O_2732,N_23750,N_24025);
or UO_2733 (O_2733,N_21405,N_20135);
nor UO_2734 (O_2734,N_24679,N_24198);
nand UO_2735 (O_2735,N_21265,N_21132);
nor UO_2736 (O_2736,N_21119,N_23780);
nor UO_2737 (O_2737,N_23925,N_21241);
nor UO_2738 (O_2738,N_20678,N_24039);
nor UO_2739 (O_2739,N_22818,N_20077);
nor UO_2740 (O_2740,N_20949,N_21973);
and UO_2741 (O_2741,N_24168,N_22895);
or UO_2742 (O_2742,N_23795,N_22039);
nand UO_2743 (O_2743,N_20794,N_22818);
nand UO_2744 (O_2744,N_24342,N_20940);
and UO_2745 (O_2745,N_23990,N_24845);
xnor UO_2746 (O_2746,N_23711,N_24231);
or UO_2747 (O_2747,N_24502,N_23053);
or UO_2748 (O_2748,N_23627,N_22041);
nor UO_2749 (O_2749,N_20804,N_22390);
xnor UO_2750 (O_2750,N_24580,N_24413);
xnor UO_2751 (O_2751,N_24674,N_22216);
or UO_2752 (O_2752,N_23998,N_22412);
or UO_2753 (O_2753,N_24593,N_22173);
xnor UO_2754 (O_2754,N_21425,N_21713);
or UO_2755 (O_2755,N_20176,N_23719);
nor UO_2756 (O_2756,N_23496,N_21629);
nand UO_2757 (O_2757,N_23934,N_23717);
or UO_2758 (O_2758,N_20530,N_24132);
nand UO_2759 (O_2759,N_24210,N_22812);
nand UO_2760 (O_2760,N_22624,N_21510);
or UO_2761 (O_2761,N_21595,N_22602);
and UO_2762 (O_2762,N_23903,N_22208);
and UO_2763 (O_2763,N_22942,N_22874);
and UO_2764 (O_2764,N_24215,N_22601);
and UO_2765 (O_2765,N_22824,N_21656);
nor UO_2766 (O_2766,N_22975,N_24211);
or UO_2767 (O_2767,N_24870,N_22056);
and UO_2768 (O_2768,N_22752,N_22275);
or UO_2769 (O_2769,N_23190,N_21295);
nor UO_2770 (O_2770,N_21231,N_23785);
and UO_2771 (O_2771,N_23547,N_24938);
or UO_2772 (O_2772,N_23943,N_24931);
nor UO_2773 (O_2773,N_21482,N_21149);
nor UO_2774 (O_2774,N_23702,N_22478);
nor UO_2775 (O_2775,N_24188,N_21620);
and UO_2776 (O_2776,N_21406,N_22576);
xor UO_2777 (O_2777,N_23906,N_22653);
and UO_2778 (O_2778,N_22413,N_24839);
and UO_2779 (O_2779,N_23788,N_24212);
and UO_2780 (O_2780,N_20757,N_22010);
xnor UO_2781 (O_2781,N_21553,N_20844);
nand UO_2782 (O_2782,N_23490,N_20036);
and UO_2783 (O_2783,N_24215,N_24708);
nand UO_2784 (O_2784,N_24873,N_23230);
or UO_2785 (O_2785,N_23185,N_23078);
or UO_2786 (O_2786,N_20364,N_23630);
and UO_2787 (O_2787,N_20112,N_23410);
and UO_2788 (O_2788,N_21396,N_22374);
or UO_2789 (O_2789,N_22816,N_24104);
nand UO_2790 (O_2790,N_22758,N_24624);
xnor UO_2791 (O_2791,N_24409,N_23558);
nand UO_2792 (O_2792,N_20689,N_23547);
or UO_2793 (O_2793,N_22619,N_22678);
nand UO_2794 (O_2794,N_21973,N_24919);
or UO_2795 (O_2795,N_24005,N_20929);
nor UO_2796 (O_2796,N_24885,N_20278);
or UO_2797 (O_2797,N_22080,N_23475);
nand UO_2798 (O_2798,N_21783,N_21124);
nand UO_2799 (O_2799,N_21971,N_23867);
and UO_2800 (O_2800,N_20772,N_21936);
and UO_2801 (O_2801,N_20478,N_21594);
nor UO_2802 (O_2802,N_20827,N_23147);
and UO_2803 (O_2803,N_20974,N_23667);
nand UO_2804 (O_2804,N_22502,N_20536);
xnor UO_2805 (O_2805,N_21865,N_22208);
xor UO_2806 (O_2806,N_21123,N_22012);
and UO_2807 (O_2807,N_20600,N_22426);
nand UO_2808 (O_2808,N_21872,N_22062);
nand UO_2809 (O_2809,N_22320,N_23219);
nand UO_2810 (O_2810,N_24052,N_22729);
nor UO_2811 (O_2811,N_21823,N_20500);
xor UO_2812 (O_2812,N_24193,N_23780);
xnor UO_2813 (O_2813,N_20949,N_23611);
and UO_2814 (O_2814,N_21577,N_22729);
nand UO_2815 (O_2815,N_21608,N_22762);
nand UO_2816 (O_2816,N_24418,N_23376);
or UO_2817 (O_2817,N_23791,N_24089);
nand UO_2818 (O_2818,N_20457,N_23681);
nand UO_2819 (O_2819,N_22607,N_21245);
xor UO_2820 (O_2820,N_22909,N_24759);
nor UO_2821 (O_2821,N_22842,N_23020);
and UO_2822 (O_2822,N_21795,N_22048);
or UO_2823 (O_2823,N_21414,N_22090);
nor UO_2824 (O_2824,N_21117,N_21084);
nand UO_2825 (O_2825,N_21354,N_23168);
xor UO_2826 (O_2826,N_23749,N_21214);
and UO_2827 (O_2827,N_21641,N_20958);
or UO_2828 (O_2828,N_21818,N_24119);
and UO_2829 (O_2829,N_22863,N_20878);
xor UO_2830 (O_2830,N_23907,N_21231);
xor UO_2831 (O_2831,N_22887,N_22713);
xor UO_2832 (O_2832,N_23999,N_23829);
and UO_2833 (O_2833,N_23844,N_20176);
nand UO_2834 (O_2834,N_23773,N_22323);
and UO_2835 (O_2835,N_23890,N_22718);
nor UO_2836 (O_2836,N_24456,N_23420);
nor UO_2837 (O_2837,N_23522,N_23325);
nor UO_2838 (O_2838,N_23498,N_24928);
and UO_2839 (O_2839,N_21611,N_20375);
and UO_2840 (O_2840,N_23455,N_22091);
nand UO_2841 (O_2841,N_21897,N_22901);
or UO_2842 (O_2842,N_20258,N_24495);
or UO_2843 (O_2843,N_20992,N_24770);
nand UO_2844 (O_2844,N_21468,N_22145);
nor UO_2845 (O_2845,N_23675,N_24865);
nand UO_2846 (O_2846,N_24463,N_24876);
nor UO_2847 (O_2847,N_24643,N_21053);
nand UO_2848 (O_2848,N_21655,N_22780);
or UO_2849 (O_2849,N_21850,N_23389);
or UO_2850 (O_2850,N_22859,N_24276);
nor UO_2851 (O_2851,N_23290,N_20731);
nor UO_2852 (O_2852,N_20921,N_21812);
or UO_2853 (O_2853,N_22061,N_23860);
nand UO_2854 (O_2854,N_22334,N_21020);
nor UO_2855 (O_2855,N_22382,N_22580);
nand UO_2856 (O_2856,N_20794,N_24458);
nor UO_2857 (O_2857,N_21376,N_21996);
nor UO_2858 (O_2858,N_21105,N_24700);
or UO_2859 (O_2859,N_24092,N_22267);
nor UO_2860 (O_2860,N_21263,N_22681);
and UO_2861 (O_2861,N_24296,N_20268);
and UO_2862 (O_2862,N_21746,N_24049);
or UO_2863 (O_2863,N_20877,N_21288);
nand UO_2864 (O_2864,N_20856,N_21319);
nand UO_2865 (O_2865,N_20874,N_21052);
nand UO_2866 (O_2866,N_23110,N_21821);
and UO_2867 (O_2867,N_21579,N_22924);
and UO_2868 (O_2868,N_20848,N_22736);
nand UO_2869 (O_2869,N_23658,N_24989);
xor UO_2870 (O_2870,N_20859,N_20979);
xor UO_2871 (O_2871,N_22039,N_23862);
nor UO_2872 (O_2872,N_23776,N_20593);
nand UO_2873 (O_2873,N_23145,N_21554);
and UO_2874 (O_2874,N_22848,N_23892);
nor UO_2875 (O_2875,N_24512,N_23376);
nor UO_2876 (O_2876,N_24251,N_21985);
and UO_2877 (O_2877,N_24939,N_21794);
or UO_2878 (O_2878,N_20562,N_23055);
nor UO_2879 (O_2879,N_24963,N_24637);
nand UO_2880 (O_2880,N_24244,N_23257);
or UO_2881 (O_2881,N_24316,N_24671);
and UO_2882 (O_2882,N_22263,N_21670);
or UO_2883 (O_2883,N_24016,N_24195);
nor UO_2884 (O_2884,N_24195,N_21388);
nor UO_2885 (O_2885,N_23711,N_23230);
or UO_2886 (O_2886,N_23218,N_21382);
and UO_2887 (O_2887,N_23539,N_21667);
or UO_2888 (O_2888,N_24686,N_21076);
nor UO_2889 (O_2889,N_21565,N_22604);
nor UO_2890 (O_2890,N_23671,N_24644);
nor UO_2891 (O_2891,N_21965,N_22051);
or UO_2892 (O_2892,N_24800,N_21539);
or UO_2893 (O_2893,N_23313,N_24723);
nand UO_2894 (O_2894,N_24253,N_24756);
and UO_2895 (O_2895,N_20452,N_21533);
or UO_2896 (O_2896,N_20691,N_22728);
nor UO_2897 (O_2897,N_21978,N_21100);
xnor UO_2898 (O_2898,N_23814,N_20256);
xor UO_2899 (O_2899,N_21039,N_23808);
and UO_2900 (O_2900,N_24195,N_20767);
or UO_2901 (O_2901,N_22166,N_23889);
nor UO_2902 (O_2902,N_21700,N_20484);
xor UO_2903 (O_2903,N_21814,N_22723);
nand UO_2904 (O_2904,N_20672,N_20955);
nor UO_2905 (O_2905,N_24895,N_20143);
and UO_2906 (O_2906,N_24878,N_21705);
or UO_2907 (O_2907,N_22351,N_24250);
xor UO_2908 (O_2908,N_23676,N_22178);
nor UO_2909 (O_2909,N_21055,N_21931);
nand UO_2910 (O_2910,N_22326,N_22805);
or UO_2911 (O_2911,N_24183,N_23281);
nor UO_2912 (O_2912,N_21492,N_20868);
or UO_2913 (O_2913,N_23205,N_22849);
xnor UO_2914 (O_2914,N_23419,N_22160);
nor UO_2915 (O_2915,N_24088,N_24395);
and UO_2916 (O_2916,N_23644,N_21028);
xor UO_2917 (O_2917,N_21226,N_24678);
or UO_2918 (O_2918,N_20643,N_22845);
or UO_2919 (O_2919,N_24802,N_21670);
xor UO_2920 (O_2920,N_21741,N_21933);
nor UO_2921 (O_2921,N_22720,N_23827);
or UO_2922 (O_2922,N_23483,N_23885);
nand UO_2923 (O_2923,N_21651,N_22888);
nor UO_2924 (O_2924,N_21532,N_21708);
or UO_2925 (O_2925,N_23984,N_24795);
nand UO_2926 (O_2926,N_21469,N_21507);
nand UO_2927 (O_2927,N_22938,N_20870);
nand UO_2928 (O_2928,N_22481,N_22640);
or UO_2929 (O_2929,N_22804,N_23105);
and UO_2930 (O_2930,N_22284,N_22170);
nand UO_2931 (O_2931,N_20652,N_22264);
nand UO_2932 (O_2932,N_20688,N_24323);
nor UO_2933 (O_2933,N_22626,N_23964);
and UO_2934 (O_2934,N_23644,N_20891);
nor UO_2935 (O_2935,N_23840,N_20380);
nand UO_2936 (O_2936,N_20564,N_20272);
nand UO_2937 (O_2937,N_23043,N_24313);
or UO_2938 (O_2938,N_21777,N_22669);
nor UO_2939 (O_2939,N_22341,N_21000);
and UO_2940 (O_2940,N_21217,N_22218);
or UO_2941 (O_2941,N_23260,N_24950);
nand UO_2942 (O_2942,N_24876,N_23938);
or UO_2943 (O_2943,N_20518,N_23254);
nand UO_2944 (O_2944,N_24692,N_24770);
nand UO_2945 (O_2945,N_23393,N_20162);
and UO_2946 (O_2946,N_22422,N_20169);
and UO_2947 (O_2947,N_23737,N_22224);
or UO_2948 (O_2948,N_23102,N_22801);
or UO_2949 (O_2949,N_24615,N_22138);
and UO_2950 (O_2950,N_23964,N_22996);
xor UO_2951 (O_2951,N_21114,N_24893);
and UO_2952 (O_2952,N_21983,N_21910);
or UO_2953 (O_2953,N_24777,N_20035);
or UO_2954 (O_2954,N_22189,N_23064);
nor UO_2955 (O_2955,N_20400,N_21572);
nand UO_2956 (O_2956,N_21865,N_23939);
nand UO_2957 (O_2957,N_23987,N_21792);
xnor UO_2958 (O_2958,N_24224,N_21010);
and UO_2959 (O_2959,N_23650,N_23152);
or UO_2960 (O_2960,N_21396,N_23051);
nor UO_2961 (O_2961,N_21858,N_24742);
or UO_2962 (O_2962,N_20503,N_24366);
and UO_2963 (O_2963,N_24164,N_21604);
nor UO_2964 (O_2964,N_21639,N_22997);
nand UO_2965 (O_2965,N_23728,N_20874);
nor UO_2966 (O_2966,N_21200,N_20354);
or UO_2967 (O_2967,N_20649,N_22771);
and UO_2968 (O_2968,N_21827,N_24304);
or UO_2969 (O_2969,N_20996,N_23091);
or UO_2970 (O_2970,N_24298,N_23639);
nand UO_2971 (O_2971,N_21759,N_23945);
and UO_2972 (O_2972,N_20448,N_22243);
or UO_2973 (O_2973,N_23791,N_24390);
nor UO_2974 (O_2974,N_22841,N_22736);
or UO_2975 (O_2975,N_22616,N_20110);
nand UO_2976 (O_2976,N_22792,N_22811);
nand UO_2977 (O_2977,N_24746,N_21559);
and UO_2978 (O_2978,N_21712,N_22550);
nor UO_2979 (O_2979,N_22443,N_24798);
or UO_2980 (O_2980,N_22287,N_21866);
and UO_2981 (O_2981,N_23537,N_21112);
and UO_2982 (O_2982,N_24689,N_24444);
and UO_2983 (O_2983,N_22070,N_21614);
or UO_2984 (O_2984,N_22661,N_21387);
or UO_2985 (O_2985,N_20653,N_21317);
or UO_2986 (O_2986,N_24503,N_21391);
nor UO_2987 (O_2987,N_22433,N_22504);
nor UO_2988 (O_2988,N_23345,N_20963);
nor UO_2989 (O_2989,N_22705,N_21319);
nand UO_2990 (O_2990,N_24432,N_23814);
nor UO_2991 (O_2991,N_23453,N_24131);
nand UO_2992 (O_2992,N_20925,N_21127);
nand UO_2993 (O_2993,N_22139,N_22051);
or UO_2994 (O_2994,N_21605,N_22704);
or UO_2995 (O_2995,N_22919,N_22786);
or UO_2996 (O_2996,N_22962,N_24218);
and UO_2997 (O_2997,N_21441,N_22566);
or UO_2998 (O_2998,N_22311,N_22771);
nor UO_2999 (O_2999,N_24707,N_21651);
endmodule