module basic_2000_20000_2500_25_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_39,In_758);
nand U1 (N_1,In_212,In_1741);
nor U2 (N_2,In_67,In_1602);
nand U3 (N_3,In_1961,In_1742);
nor U4 (N_4,In_603,In_661);
and U5 (N_5,In_848,In_789);
or U6 (N_6,In_694,In_541);
and U7 (N_7,In_897,In_1829);
or U8 (N_8,In_313,In_1395);
or U9 (N_9,In_1784,In_832);
or U10 (N_10,In_851,In_600);
nor U11 (N_11,In_879,In_1931);
nor U12 (N_12,In_143,In_1558);
and U13 (N_13,In_816,In_785);
or U14 (N_14,In_517,In_357);
nand U15 (N_15,In_1330,In_1086);
xor U16 (N_16,In_1156,In_1247);
xnor U17 (N_17,In_931,In_369);
and U18 (N_18,In_1475,In_1481);
and U19 (N_19,In_1263,In_350);
nor U20 (N_20,In_902,In_1325);
and U21 (N_21,In_1660,In_1903);
or U22 (N_22,In_852,In_1027);
and U23 (N_23,In_1062,In_1268);
xnor U24 (N_24,In_1081,In_1009);
nand U25 (N_25,In_1709,In_178);
xor U26 (N_26,In_1810,In_91);
or U27 (N_27,In_1934,In_1382);
or U28 (N_28,In_415,In_397);
xnor U29 (N_29,In_891,In_76);
and U30 (N_30,In_786,In_386);
nand U31 (N_31,In_1729,In_381);
and U32 (N_32,In_858,In_1805);
xor U33 (N_33,In_493,In_577);
and U34 (N_34,In_1982,In_1289);
and U35 (N_35,In_332,In_294);
xor U36 (N_36,In_177,In_4);
xnor U37 (N_37,In_1985,In_1441);
nor U38 (N_38,In_1643,In_973);
xor U39 (N_39,In_1292,In_1042);
or U40 (N_40,In_1588,In_1762);
nor U41 (N_41,In_187,In_671);
nand U42 (N_42,In_1986,In_1831);
and U43 (N_43,In_1484,In_1275);
nand U44 (N_44,In_1642,In_85);
nor U45 (N_45,In_881,In_1652);
nor U46 (N_46,In_193,In_1527);
nand U47 (N_47,In_261,In_285);
nor U48 (N_48,In_452,In_1241);
nand U49 (N_49,In_481,In_1515);
xor U50 (N_50,In_992,In_251);
nor U51 (N_51,In_225,In_1257);
nand U52 (N_52,In_329,In_1235);
xnor U53 (N_53,In_314,In_213);
nor U54 (N_54,In_245,In_1824);
xnor U55 (N_55,In_861,In_923);
nand U56 (N_56,In_728,In_96);
or U57 (N_57,In_61,In_1743);
or U58 (N_58,In_1057,In_811);
or U59 (N_59,In_1041,In_1299);
xor U60 (N_60,In_1284,In_52);
or U61 (N_61,In_834,In_1685);
nor U62 (N_62,In_1862,In_673);
xor U63 (N_63,In_431,In_627);
nand U64 (N_64,In_706,In_633);
and U65 (N_65,In_530,In_746);
nor U66 (N_66,In_954,In_801);
or U67 (N_67,In_1840,In_782);
and U68 (N_68,In_1113,In_636);
nor U69 (N_69,In_1434,In_169);
and U70 (N_70,In_1625,In_1074);
and U71 (N_71,In_1253,In_641);
xnor U72 (N_72,In_1087,In_1679);
nor U73 (N_73,In_802,In_844);
or U74 (N_74,In_1905,In_1509);
nand U75 (N_75,In_1448,In_62);
or U76 (N_76,In_293,In_911);
and U77 (N_77,In_1783,In_1560);
or U78 (N_78,In_186,In_937);
xnor U79 (N_79,In_148,In_716);
and U80 (N_80,In_48,In_1281);
nor U81 (N_81,In_35,In_1384);
nand U82 (N_82,In_1954,In_841);
xor U83 (N_83,In_1133,In_523);
xnor U84 (N_84,In_1953,In_1803);
nand U85 (N_85,In_1091,In_1834);
and U86 (N_86,In_1970,In_1766);
nand U87 (N_87,In_505,In_978);
or U88 (N_88,In_1635,In_915);
nand U89 (N_89,In_1720,In_1261);
nand U90 (N_90,In_191,In_687);
or U91 (N_91,In_630,In_1442);
xor U92 (N_92,In_404,In_1374);
nor U93 (N_93,In_1344,In_643);
nand U94 (N_94,In_1606,In_270);
nand U95 (N_95,In_1624,In_578);
and U96 (N_96,In_1114,In_1590);
xnor U97 (N_97,In_463,In_131);
or U98 (N_98,In_367,In_232);
nor U99 (N_99,In_714,In_1109);
and U100 (N_100,In_124,In_1266);
or U101 (N_101,In_1872,In_920);
and U102 (N_102,In_24,In_260);
nor U103 (N_103,In_1759,In_885);
xnor U104 (N_104,In_1549,In_1362);
nand U105 (N_105,In_1782,In_1035);
or U106 (N_106,In_133,In_696);
and U107 (N_107,In_908,In_859);
and U108 (N_108,In_818,In_63);
nand U109 (N_109,In_112,In_1820);
nor U110 (N_110,In_1301,In_1052);
nand U111 (N_111,In_435,In_1006);
or U112 (N_112,In_649,In_840);
nor U113 (N_113,In_886,In_1911);
and U114 (N_114,In_1236,In_1376);
nand U115 (N_115,In_953,In_779);
and U116 (N_116,In_70,In_1676);
or U117 (N_117,In_482,In_1956);
xnor U118 (N_118,In_797,In_1496);
or U119 (N_119,In_1693,In_866);
nand U120 (N_120,In_37,In_1227);
xor U121 (N_121,In_146,In_325);
nand U122 (N_122,In_1189,In_1068);
nand U123 (N_123,In_1963,In_1815);
xnor U124 (N_124,In_443,In_149);
or U125 (N_125,In_1288,In_1898);
and U126 (N_126,In_1196,In_814);
xor U127 (N_127,In_762,In_123);
nand U128 (N_128,In_1518,In_916);
nand U129 (N_129,In_719,In_1924);
or U130 (N_130,In_1517,In_1220);
or U131 (N_131,In_228,In_1184);
and U132 (N_132,In_701,In_1134);
or U133 (N_133,In_1490,In_73);
and U134 (N_134,In_1812,In_1244);
and U135 (N_135,In_1525,In_669);
and U136 (N_136,In_1878,In_1798);
or U137 (N_137,In_229,In_152);
or U138 (N_138,In_849,In_1912);
nand U139 (N_139,In_17,In_1663);
and U140 (N_140,In_922,In_581);
and U141 (N_141,In_1700,In_1310);
or U142 (N_142,In_190,In_218);
or U143 (N_143,In_257,In_1445);
or U144 (N_144,In_355,In_1576);
xor U145 (N_145,In_489,In_555);
xor U146 (N_146,In_1192,In_54);
or U147 (N_147,In_1021,In_1402);
nand U148 (N_148,In_557,In_119);
or U149 (N_149,In_766,In_180);
and U150 (N_150,In_1877,In_1180);
or U151 (N_151,In_663,In_929);
nand U152 (N_152,In_1223,In_1233);
xnor U153 (N_153,In_157,In_1753);
and U154 (N_154,In_315,In_1336);
or U155 (N_155,In_726,In_1976);
or U156 (N_156,In_1311,In_1152);
nor U157 (N_157,In_296,In_1464);
or U158 (N_158,In_1415,In_1228);
nor U159 (N_159,In_888,In_1066);
or U160 (N_160,In_1867,In_1339);
xnor U161 (N_161,In_479,In_536);
nor U162 (N_162,In_1044,In_1486);
nor U163 (N_163,In_1162,In_47);
xor U164 (N_164,In_943,In_55);
or U165 (N_165,In_938,In_697);
xnor U166 (N_166,In_952,In_769);
nand U167 (N_167,In_1396,In_60);
xnor U168 (N_168,In_1201,In_259);
xor U169 (N_169,In_7,In_1680);
xor U170 (N_170,In_933,In_1669);
nor U171 (N_171,In_1796,In_934);
nand U172 (N_172,In_1768,In_188);
nor U173 (N_173,In_1639,In_1125);
and U174 (N_174,In_775,In_1927);
nor U175 (N_175,In_1064,In_38);
nor U176 (N_176,In_670,In_566);
xor U177 (N_177,In_356,In_1505);
or U178 (N_178,In_826,In_808);
or U179 (N_179,In_455,In_1168);
xnor U180 (N_180,In_1592,In_1452);
and U181 (N_181,In_488,In_292);
nand U182 (N_182,In_1893,In_1090);
or U183 (N_183,In_1955,In_319);
or U184 (N_184,In_1340,In_471);
or U185 (N_185,In_1966,In_383);
nor U186 (N_186,In_829,In_1410);
nand U187 (N_187,In_9,In_1342);
or U188 (N_188,In_604,In_1422);
or U189 (N_189,In_1175,In_476);
xor U190 (N_190,In_1404,In_29);
nand U191 (N_191,In_1533,In_1391);
and U192 (N_192,In_1230,In_1992);
xor U193 (N_193,In_25,In_1455);
xnor U194 (N_194,In_657,In_15);
xnor U195 (N_195,In_1357,In_1556);
nor U196 (N_196,In_1489,In_1914);
nor U197 (N_197,In_596,In_1430);
nor U198 (N_198,In_1835,In_1072);
nor U199 (N_199,In_1388,In_1032);
xor U200 (N_200,In_1463,In_1545);
xor U201 (N_201,In_1403,In_215);
and U202 (N_202,In_371,In_1826);
nand U203 (N_203,In_884,In_871);
and U204 (N_204,In_1744,In_948);
or U205 (N_205,In_1569,In_1425);
nor U206 (N_206,In_1919,In_552);
xor U207 (N_207,In_800,In_1273);
nor U208 (N_208,In_1651,In_1346);
nor U209 (N_209,In_265,In_1684);
and U210 (N_210,In_1169,In_1722);
xnor U211 (N_211,In_1521,In_1896);
or U212 (N_212,In_1735,In_1731);
and U213 (N_213,In_1389,In_253);
or U214 (N_214,In_790,In_983);
nand U215 (N_215,In_273,In_745);
nand U216 (N_216,In_524,In_1377);
xor U217 (N_217,In_1671,In_318);
nand U218 (N_218,In_617,In_410);
nor U219 (N_219,In_174,In_1933);
and U220 (N_220,In_1078,In_153);
or U221 (N_221,In_1780,In_194);
or U222 (N_222,In_1269,In_772);
and U223 (N_223,In_733,In_1314);
and U224 (N_224,In_1015,In_1587);
or U225 (N_225,In_873,In_184);
nand U226 (N_226,In_221,In_1324);
nand U227 (N_227,In_1777,In_1551);
nand U228 (N_228,In_1423,In_182);
and U229 (N_229,In_1522,In_1502);
nor U230 (N_230,In_804,In_1029);
nand U231 (N_231,In_1980,In_1534);
nor U232 (N_232,In_906,In_450);
nand U233 (N_233,In_1689,In_1013);
xnor U234 (N_234,In_72,In_941);
xor U235 (N_235,In_887,In_864);
nand U236 (N_236,In_89,In_862);
or U237 (N_237,In_351,In_693);
nor U238 (N_238,In_1000,In_1245);
nand U239 (N_239,In_110,In_1922);
or U240 (N_240,In_680,In_1132);
xnor U241 (N_241,In_1984,In_837);
nor U242 (N_242,In_1876,In_1280);
nand U243 (N_243,In_1531,In_1217);
nor U244 (N_244,In_619,In_827);
or U245 (N_245,In_244,In_104);
xnor U246 (N_246,In_1099,In_1547);
nand U247 (N_247,In_1776,In_1667);
xor U248 (N_248,In_546,In_685);
xor U249 (N_249,In_1054,In_1349);
and U250 (N_250,In_1051,In_1668);
xnor U251 (N_251,In_704,In_1839);
nor U252 (N_252,In_903,In_12);
and U253 (N_253,In_195,In_691);
and U254 (N_254,In_799,In_1649);
xnor U255 (N_255,In_477,In_1694);
xnor U256 (N_256,In_1974,In_1364);
and U257 (N_257,In_1707,In_1967);
and U258 (N_258,In_1126,In_1881);
nand U259 (N_259,In_1946,In_979);
or U260 (N_260,In_1987,In_1510);
nand U261 (N_261,In_935,In_1716);
nand U262 (N_262,In_635,In_1016);
or U263 (N_263,In_398,In_51);
xnor U264 (N_264,In_1629,In_1504);
nand U265 (N_265,In_1902,In_497);
nand U266 (N_266,In_1250,In_936);
and U267 (N_267,In_1645,In_1412);
xor U268 (N_268,In_269,In_1644);
or U269 (N_269,In_1355,In_1740);
nand U270 (N_270,In_845,In_1785);
nand U271 (N_271,In_1350,In_173);
nand U272 (N_272,In_1774,In_995);
xnor U273 (N_273,In_1672,In_36);
and U274 (N_274,In_1083,In_258);
and U275 (N_275,In_907,In_1381);
and U276 (N_276,In_773,In_1399);
or U277 (N_277,In_855,In_1120);
nand U278 (N_278,In_1012,In_1014);
xor U279 (N_279,In_1631,In_1234);
or U280 (N_280,In_699,In_139);
nor U281 (N_281,In_1771,In_918);
and U282 (N_282,In_1347,In_1313);
or U283 (N_283,In_1908,In_162);
nand U284 (N_284,In_1176,In_1335);
or U285 (N_285,In_1387,In_407);
xor U286 (N_286,In_729,In_723);
xor U287 (N_287,In_278,In_1371);
nand U288 (N_288,In_1207,In_660);
nand U289 (N_289,In_8,In_831);
or U290 (N_290,In_1159,In_606);
or U291 (N_291,In_612,In_1802);
and U292 (N_292,In_436,In_677);
or U293 (N_293,In_1601,In_1711);
or U294 (N_294,In_1623,In_1127);
nor U295 (N_295,In_342,In_263);
and U296 (N_296,In_107,In_784);
nor U297 (N_297,In_1240,In_1186);
xor U298 (N_298,In_1322,In_761);
or U299 (N_299,In_1345,In_243);
or U300 (N_300,In_155,In_474);
nand U301 (N_301,In_653,In_1191);
or U302 (N_302,In_6,In_770);
or U303 (N_303,In_360,In_1252);
and U304 (N_304,In_28,In_0);
and U305 (N_305,In_893,In_298);
nor U306 (N_306,In_632,In_585);
and U307 (N_307,In_921,In_1630);
xor U308 (N_308,In_1706,In_1855);
nor U309 (N_309,In_1373,In_1101);
xnor U310 (N_310,In_1895,In_589);
nand U311 (N_311,In_1188,In_1461);
or U312 (N_312,In_1365,In_764);
nand U313 (N_313,In_445,In_1929);
nor U314 (N_314,In_242,In_628);
nand U315 (N_315,In_1477,In_1304);
nor U316 (N_316,In_151,In_950);
and U317 (N_317,In_890,In_1677);
nand U318 (N_318,In_521,In_209);
nor U319 (N_319,In_1728,In_1938);
nand U320 (N_320,In_721,In_88);
or U321 (N_321,In_376,In_792);
nor U322 (N_322,In_57,In_125);
and U323 (N_323,In_272,In_1612);
xor U324 (N_324,In_1899,In_1869);
nor U325 (N_325,In_277,In_59);
xnor U326 (N_326,In_1363,In_867);
or U327 (N_327,In_1254,In_1747);
nand U328 (N_328,In_511,In_1714);
nor U329 (N_329,In_1880,In_956);
nand U330 (N_330,In_542,In_1761);
xnor U331 (N_331,In_100,In_533);
and U332 (N_332,In_598,In_711);
xor U333 (N_333,In_365,In_1599);
and U334 (N_334,In_778,In_1559);
nor U335 (N_335,In_1928,In_1750);
nand U336 (N_336,In_1456,In_84);
nor U337 (N_337,In_545,In_828);
nand U338 (N_338,In_501,In_1571);
nor U339 (N_339,In_427,In_506);
and U340 (N_340,In_1851,In_1331);
nor U341 (N_341,In_317,In_925);
or U342 (N_342,In_1237,In_1255);
and U343 (N_343,In_896,In_1333);
nor U344 (N_344,In_1697,In_927);
nand U345 (N_345,In_206,In_1795);
nor U346 (N_346,In_1524,In_1585);
xnor U347 (N_347,In_1203,In_1832);
or U348 (N_348,In_868,In_1633);
and U349 (N_349,In_564,In_163);
nor U350 (N_350,In_960,In_374);
nor U351 (N_351,In_1594,In_13);
nor U352 (N_352,In_199,In_81);
and U353 (N_353,In_1181,In_754);
xor U354 (N_354,In_1951,In_1959);
nor U355 (N_355,In_965,In_1030);
nor U356 (N_356,In_1121,In_771);
and U357 (N_357,In_132,In_639);
and U358 (N_358,In_495,In_166);
xnor U359 (N_359,In_1123,In_1596);
nor U360 (N_360,In_625,In_1249);
and U361 (N_361,In_744,In_835);
xnor U362 (N_362,In_974,In_568);
or U363 (N_363,In_1418,In_1562);
and U364 (N_364,In_1248,In_967);
and U365 (N_365,In_1674,In_428);
xnor U366 (N_366,In_1321,In_1329);
nor U367 (N_367,In_940,In_1546);
or U368 (N_368,In_705,In_1413);
xnor U369 (N_369,In_1307,In_403);
nor U370 (N_370,In_1096,In_1164);
xnor U371 (N_371,In_675,In_1420);
and U372 (N_372,In_985,In_1137);
and U373 (N_373,In_1838,In_608);
xor U374 (N_374,In_1197,In_1246);
nand U375 (N_375,In_850,In_498);
or U376 (N_376,In_79,In_543);
nor U377 (N_377,In_1792,In_1317);
and U378 (N_378,In_1309,In_1295);
nand U379 (N_379,In_1686,In_650);
xnor U380 (N_380,In_880,In_1023);
and U381 (N_381,In_1219,In_1298);
or U382 (N_382,In_485,In_1031);
nor U383 (N_383,In_1047,In_447);
and U384 (N_384,In_1320,In_1804);
and U385 (N_385,In_553,In_1069);
nand U386 (N_386,In_777,In_1721);
xnor U387 (N_387,In_624,In_579);
xnor U388 (N_388,In_392,In_19);
xor U389 (N_389,In_117,In_1925);
and U390 (N_390,In_513,In_550);
and U391 (N_391,In_267,In_1038);
xnor U392 (N_392,In_1765,In_432);
nor U393 (N_393,In_1353,In_565);
xnor U394 (N_394,In_1323,In_1202);
nand U395 (N_395,In_1143,In_930);
nor U396 (N_396,In_526,In_394);
and U397 (N_397,In_1821,In_698);
and U398 (N_398,In_1909,In_1739);
and U399 (N_399,In_105,In_1865);
nand U400 (N_400,In_520,In_684);
xor U401 (N_401,In_361,In_791);
nor U402 (N_402,In_889,In_430);
nor U403 (N_403,In_1119,In_185);
and U404 (N_404,In_514,In_1183);
nor U405 (N_405,In_1470,In_210);
xor U406 (N_406,In_44,In_1089);
nor U407 (N_407,In_420,In_1526);
xnor U408 (N_408,In_373,In_1724);
and U409 (N_409,In_1882,In_3);
nor U410 (N_410,In_1846,In_448);
and U411 (N_411,In_709,In_279);
or U412 (N_412,In_378,In_1787);
nand U413 (N_413,In_563,In_715);
xor U414 (N_414,In_339,In_45);
xnor U415 (N_415,In_413,In_1135);
nand U416 (N_416,In_1675,In_18);
or U417 (N_417,In_454,In_334);
nand U418 (N_418,In_980,In_424);
nand U419 (N_419,In_1405,In_231);
nand U420 (N_420,In_1209,In_1613);
and U421 (N_421,In_1174,In_534);
xnor U422 (N_422,In_1568,In_1411);
and U423 (N_423,In_1226,In_1681);
nor U424 (N_424,In_1968,In_1198);
nor U425 (N_425,In_1904,In_14);
or U426 (N_426,In_256,In_803);
xnor U427 (N_427,In_1210,In_993);
nor U428 (N_428,In_1888,In_853);
nor U429 (N_429,In_99,In_1122);
nand U430 (N_430,In_1375,In_570);
nor U431 (N_431,In_516,In_1758);
xor U432 (N_432,In_307,In_748);
and U433 (N_433,In_1178,In_1102);
and U434 (N_434,In_1161,In_1769);
xor U435 (N_435,In_796,In_142);
or U436 (N_436,In_987,In_1414);
and U437 (N_437,In_358,In_1604);
nand U438 (N_438,In_1930,In_1705);
nand U439 (N_439,In_1332,In_90);
xnor U440 (N_440,In_1258,In_1084);
nor U441 (N_441,In_924,In_1216);
nand U442 (N_442,In_756,In_264);
or U443 (N_443,In_1100,In_327);
and U444 (N_444,In_1428,In_976);
or U445 (N_445,In_882,In_349);
or U446 (N_446,In_1628,In_399);
nor U447 (N_447,In_912,In_1566);
xor U448 (N_448,In_678,In_695);
nand U449 (N_449,In_1971,In_1037);
nand U450 (N_450,In_1608,In_275);
nand U451 (N_451,In_1507,In_137);
nor U452 (N_452,In_1557,In_1398);
and U453 (N_453,In_266,In_580);
nand U454 (N_454,In_1182,In_1767);
xnor U455 (N_455,In_1935,In_1570);
nand U456 (N_456,In_651,In_759);
and U457 (N_457,In_1222,In_652);
xor U458 (N_458,In_741,In_408);
or U459 (N_459,In_1286,In_1055);
nor U460 (N_460,In_1265,In_990);
and U461 (N_461,In_958,In_1467);
and U462 (N_462,In_127,In_1793);
xor U463 (N_463,In_1495,In_1683);
and U464 (N_464,In_1528,In_457);
nor U465 (N_465,In_755,In_1294);
or U466 (N_466,In_344,In_1480);
and U467 (N_467,In_224,In_21);
or U468 (N_468,In_1199,In_631);
and U469 (N_469,In_220,In_1993);
nor U470 (N_470,In_101,In_1943);
nand U471 (N_471,In_751,In_322);
nand U472 (N_472,In_658,In_1020);
and U473 (N_473,In_1147,In_136);
xor U474 (N_474,In_573,In_1341);
nand U475 (N_475,In_688,In_441);
nand U476 (N_476,In_629,In_1138);
nor U477 (N_477,In_1530,In_102);
or U478 (N_478,In_913,In_108);
nor U479 (N_479,In_354,In_611);
and U480 (N_480,In_1861,In_1544);
nor U481 (N_481,In_717,In_402);
nor U482 (N_482,In_308,In_1276);
or U483 (N_483,In_97,In_535);
and U484 (N_484,In_1636,In_703);
nand U485 (N_485,In_1429,In_200);
or U486 (N_486,In_982,In_1703);
nand U487 (N_487,In_393,In_1318);
nand U488 (N_488,In_1842,In_1727);
xnor U489 (N_489,In_372,In_1080);
and U490 (N_490,In_1239,In_1139);
xnor U491 (N_491,In_33,In_981);
nor U492 (N_492,In_1224,In_122);
xor U493 (N_493,In_710,In_348);
or U494 (N_494,In_647,In_150);
and U495 (N_495,In_1973,In_216);
xor U496 (N_496,In_171,In_1807);
nand U497 (N_497,In_926,In_1775);
nand U498 (N_498,In_525,In_310);
nand U499 (N_499,In_1290,In_1165);
nand U500 (N_500,In_1603,In_268);
or U501 (N_501,In_337,In_1704);
and U502 (N_502,In_1338,In_824);
or U503 (N_503,In_1638,In_1756);
xnor U504 (N_504,In_515,In_400);
nor U505 (N_505,In_23,In_1615);
nor U506 (N_506,In_1471,In_749);
nand U507 (N_507,In_1435,In_549);
and U508 (N_508,In_1918,In_1040);
and U509 (N_509,In_364,In_1950);
or U510 (N_510,In_490,In_1243);
xor U511 (N_511,In_1699,In_664);
and U512 (N_512,In_788,In_1607);
nand U513 (N_513,In_1659,In_1438);
and U514 (N_514,In_1488,In_1696);
nor U515 (N_515,In_738,In_567);
or U516 (N_516,In_970,In_503);
nand U517 (N_517,In_949,In_1370);
and U518 (N_518,In_262,In_1781);
and U519 (N_519,In_391,In_686);
or U520 (N_520,In_1885,In_1107);
nand U521 (N_521,In_467,In_1945);
nor U522 (N_522,In_1179,In_1906);
and U523 (N_523,In_1972,In_994);
or U524 (N_524,In_1598,In_874);
xnor U525 (N_525,In_626,In_1958);
and U526 (N_526,In_340,In_910);
or U527 (N_527,In_1011,In_50);
xor U528 (N_528,In_1641,In_158);
and U529 (N_529,In_1028,In_128);
xnor U530 (N_530,In_1474,In_297);
or U531 (N_531,In_421,In_456);
nor U532 (N_532,In_446,In_240);
or U533 (N_533,In_66,In_1948);
and U534 (N_534,In_1725,In_1897);
xor U535 (N_535,In_1212,In_894);
xnor U536 (N_536,In_1451,In_1482);
xor U537 (N_537,In_947,In_1424);
or U538 (N_538,In_1380,In_284);
and U539 (N_539,In_27,In_876);
nand U540 (N_540,In_1891,In_1019);
nand U541 (N_541,In_1901,In_202);
or U542 (N_542,In_1866,In_1287);
nand U543 (N_543,In_1491,In_1890);
or U544 (N_544,In_1308,In_1892);
xor U545 (N_545,In_548,In_1788);
nand U546 (N_546,In_103,In_1506);
nand U547 (N_547,In_370,In_1473);
or U548 (N_548,In_175,In_1837);
nand U549 (N_549,In_783,In_154);
nand U550 (N_550,In_181,In_1368);
nor U551 (N_551,In_1923,In_593);
or U552 (N_552,In_1900,In_233);
nor U553 (N_553,In_1408,In_955);
or U554 (N_554,In_1640,In_1579);
nor U555 (N_555,In_1508,In_434);
nor U556 (N_556,In_623,In_865);
and U557 (N_557,In_998,In_1001);
or U558 (N_558,In_1883,In_966);
xor U559 (N_559,In_594,In_1550);
and U560 (N_560,In_1701,In_547);
or U561 (N_561,In_727,In_722);
and U562 (N_562,In_1554,In_1046);
xnor U563 (N_563,In_964,In_1469);
nand U564 (N_564,In_1348,In_1238);
xor U565 (N_565,In_1617,In_1112);
nor U566 (N_566,In_86,In_854);
and U567 (N_567,In_438,In_1772);
nor U568 (N_568,In_1111,In_204);
nand U569 (N_569,In_1757,In_2);
or U570 (N_570,In_1650,In_856);
nor U571 (N_571,In_1597,In_1008);
or U572 (N_572,In_426,In_1005);
nor U573 (N_573,In_878,In_1478);
xor U574 (N_574,In_290,In_1437);
xnor U575 (N_575,In_914,In_144);
or U576 (N_576,In_1024,In_375);
or U577 (N_577,In_610,In_1379);
nand U578 (N_578,In_462,In_1079);
nand U579 (N_579,In_312,In_1552);
nor U580 (N_580,In_377,In_1516);
and U581 (N_581,In_1279,In_58);
or U582 (N_582,In_1426,In_1520);
xor U583 (N_583,In_1274,In_690);
nor U584 (N_584,In_1145,In_1621);
xor U585 (N_585,In_502,In_1998);
or U586 (N_586,In_939,In_558);
or U587 (N_587,In_969,In_1822);
or U588 (N_588,In_1702,In_118);
nand U589 (N_589,In_1917,In_1067);
nor U590 (N_590,In_1093,In_1397);
or U591 (N_591,In_839,In_207);
and U592 (N_592,In_323,In_1926);
nand U593 (N_593,In_1937,In_551);
xnor U594 (N_594,In_735,In_1231);
xor U595 (N_595,In_1296,In_1664);
xor U596 (N_596,In_328,In_1858);
and U597 (N_597,In_406,In_616);
or U598 (N_598,In_1539,In_1103);
nor U599 (N_599,In_1140,In_1657);
nor U600 (N_600,In_1654,In_366);
xor U601 (N_601,In_1995,In_16);
or U602 (N_602,In_1691,In_1229);
and U603 (N_603,In_560,In_602);
nand U604 (N_604,In_1749,In_962);
and U605 (N_605,In_883,In_1150);
nor U606 (N_606,In_5,In_1886);
nand U607 (N_607,In_1070,In_1555);
xor U608 (N_608,In_1921,In_380);
and U609 (N_609,In_198,In_1653);
and U610 (N_610,In_972,In_1833);
or U611 (N_611,In_164,In_1609);
nor U612 (N_612,In_459,In_1097);
nor U613 (N_613,In_469,In_599);
or U614 (N_614,In_183,In_1048);
or U615 (N_615,In_847,In_607);
or U616 (N_616,In_531,In_1218);
and U617 (N_617,In_997,In_1458);
or U618 (N_618,In_429,In_167);
nand U619 (N_619,In_1626,In_1719);
or U620 (N_620,In_418,In_1334);
nand U621 (N_621,In_1733,In_32);
nor U622 (N_622,In_644,In_532);
and U623 (N_623,In_810,In_389);
and U624 (N_624,In_1367,In_1170);
and U625 (N_625,In_395,In_648);
xnor U626 (N_626,In_659,In_241);
xor U627 (N_627,In_1619,In_1887);
and U628 (N_628,In_1206,In_1200);
and U629 (N_629,In_945,In_1827);
nand U630 (N_630,In_1647,In_1);
and U631 (N_631,In_1864,In_1007);
and U632 (N_632,In_1655,In_1989);
nand U633 (N_633,In_390,In_1786);
nor U634 (N_634,In_211,In_1860);
xnor U635 (N_635,In_321,In_414);
nand U636 (N_636,In_1537,In_65);
and U637 (N_637,In_78,In_1098);
nor U638 (N_638,In_637,In_757);
xor U639 (N_639,In_1043,In_857);
and U640 (N_640,In_1300,In_760);
and U641 (N_641,In_1136,In_271);
and U642 (N_642,In_1994,In_1673);
nor U643 (N_643,In_126,In_1844);
or U644 (N_644,In_26,In_1801);
or U645 (N_645,In_1859,In_80);
xor U646 (N_646,In_1462,In_236);
xnor U647 (N_647,In_156,In_306);
nor U648 (N_648,In_863,In_1789);
or U649 (N_649,In_214,In_1512);
or U650 (N_650,In_1670,In_1541);
or U651 (N_651,In_1836,In_944);
and U652 (N_652,In_472,In_1466);
nand U653 (N_653,In_554,In_1427);
xnor U654 (N_654,In_1519,In_815);
nor U655 (N_655,In_1538,In_466);
xnor U656 (N_656,In_1868,In_1085);
nor U657 (N_657,In_384,In_1717);
and U658 (N_658,In_1149,In_917);
nand U659 (N_659,In_1022,In_901);
nand U660 (N_660,In_1634,In_1561);
or U661 (N_661,In_780,In_781);
and U662 (N_662,In_338,In_1104);
and U663 (N_663,In_1155,In_1799);
xnor U664 (N_664,In_1406,In_1077);
and U665 (N_665,In_1977,In_1975);
nor U666 (N_666,In_1718,In_40);
nand U667 (N_667,In_582,In_1213);
and U668 (N_668,In_444,In_250);
nor U669 (N_669,In_1665,In_975);
and U670 (N_670,In_1116,In_519);
nor U671 (N_671,In_730,In_409);
xor U672 (N_672,In_1088,In_877);
nand U673 (N_673,In_1988,In_892);
nand U674 (N_674,In_1952,In_287);
xnor U675 (N_675,In_1637,In_343);
nor U676 (N_676,In_1589,In_1553);
and U677 (N_677,In_618,In_147);
xnor U678 (N_678,In_1194,In_1312);
and U679 (N_679,In_1773,In_528);
xor U680 (N_680,In_1282,In_458);
xor U681 (N_681,In_1204,In_286);
or U682 (N_682,In_1440,In_247);
or U683 (N_683,In_82,In_451);
and U684 (N_684,In_821,In_425);
xor U685 (N_685,In_1498,In_609);
and U686 (N_686,In_833,In_875);
nor U687 (N_687,In_1256,In_753);
xor U688 (N_688,In_1548,In_440);
xnor U689 (N_689,In_464,In_518);
or U690 (N_690,In_68,In_140);
nor U691 (N_691,In_1916,In_1913);
or U692 (N_692,In_1964,In_1076);
or U693 (N_693,In_1082,In_1151);
nor U694 (N_694,In_283,In_235);
or U695 (N_695,In_1884,In_223);
or U696 (N_696,In_1850,In_1712);
or U697 (N_697,In_574,In_352);
and U698 (N_698,In_1620,In_692);
or U699 (N_699,In_276,In_899);
xnor U700 (N_700,In_1965,In_544);
or U701 (N_701,In_1962,In_1790);
xnor U702 (N_702,In_1849,In_977);
and U703 (N_703,In_249,In_486);
nor U704 (N_704,In_1808,In_1359);
and U705 (N_705,In_1173,In_1421);
or U706 (N_706,In_1746,In_1841);
nand U707 (N_707,In_1595,In_1932);
and U708 (N_708,In_1996,In_320);
and U709 (N_709,In_470,In_230);
or U710 (N_710,In_1723,In_1940);
nand U711 (N_711,In_473,In_597);
xnor U712 (N_712,In_449,In_1460);
xor U713 (N_713,In_1369,In_1358);
xnor U714 (N_714,In_1979,In_475);
nand U715 (N_715,In_1873,In_1409);
xnor U716 (N_716,In_335,In_1271);
xnor U717 (N_717,In_1690,In_1004);
and U718 (N_718,In_77,In_1002);
xor U719 (N_719,In_1025,In_583);
nor U720 (N_720,In_765,In_1845);
xor U721 (N_721,In_42,In_170);
or U722 (N_722,In_1453,In_1171);
xnor U723 (N_723,In_305,In_1529);
or U724 (N_724,In_1503,In_1267);
and U725 (N_725,In_1770,In_1394);
nor U726 (N_726,In_909,In_991);
nand U727 (N_727,In_1319,In_838);
or U728 (N_728,In_959,In_491);
xnor U729 (N_729,In_605,In_1316);
nand U730 (N_730,In_1306,In_1763);
xnor U731 (N_731,In_94,In_1823);
or U732 (N_732,In_10,In_1616);
and U733 (N_733,In_1738,In_807);
xnor U734 (N_734,In_1148,In_556);
or U735 (N_735,In_423,In_1352);
or U736 (N_736,In_109,In_830);
or U737 (N_737,In_1957,In_665);
xor U738 (N_738,In_274,In_946);
nor U739 (N_739,In_634,In_1532);
nor U740 (N_740,In_1622,In_1565);
nor U741 (N_741,In_809,In_1809);
and U742 (N_742,In_507,In_734);
nor U743 (N_743,In_1500,In_1095);
nor U744 (N_744,In_1050,In_681);
nor U745 (N_745,In_281,In_1692);
and U746 (N_746,In_1920,In_1889);
and U747 (N_747,In_1190,In_1949);
nor U748 (N_748,In_1018,In_1487);
nand U749 (N_749,In_1614,In_1073);
and U750 (N_750,In_1293,In_1166);
or U751 (N_751,In_1185,In_461);
xor U752 (N_752,In_1075,In_1439);
nor U753 (N_753,In_141,In_1734);
and U754 (N_754,In_1816,In_1540);
and U755 (N_755,In_905,In_1999);
nor U756 (N_756,In_1354,In_1291);
nand U757 (N_757,In_1666,In_385);
nor U758 (N_758,In_1713,In_590);
nor U759 (N_759,In_1167,In_1848);
nand U760 (N_760,In_165,In_1969);
or U761 (N_761,In_1383,In_988);
or U762 (N_762,In_622,In_825);
nor U763 (N_763,In_1981,In_561);
and U764 (N_764,In_1278,In_1465);
or U765 (N_765,In_957,In_1302);
or U766 (N_766,In_1105,In_1819);
xor U767 (N_767,In_795,In_1144);
nor U768 (N_768,In_1611,In_83);
nor U769 (N_769,In_805,In_1214);
nand U770 (N_770,In_1710,In_1417);
or U771 (N_771,In_820,In_860);
xnor U772 (N_772,In_740,In_646);
nand U773 (N_773,In_1187,In_1752);
and U774 (N_774,In_291,In_1513);
nand U775 (N_775,In_341,In_1656);
xor U776 (N_776,In_1811,In_1907);
nand U777 (N_777,In_111,In_1648);
nor U778 (N_778,In_569,In_1446);
or U779 (N_779,In_1564,In_227);
nand U780 (N_780,In_656,In_1259);
and U781 (N_781,In_1272,In_1045);
xnor U782 (N_782,In_417,In_1351);
and U783 (N_783,In_613,In_1326);
nor U784 (N_784,In_620,In_1852);
nor U785 (N_785,In_1130,In_812);
nor U786 (N_786,In_1662,In_1760);
and U787 (N_787,In_1110,In_433);
or U788 (N_788,In_529,In_1748);
nor U789 (N_789,In_1610,In_1874);
and U790 (N_790,In_129,In_1071);
nand U791 (N_791,In_971,In_1944);
nand U792 (N_792,In_1327,In_919);
or U793 (N_793,In_743,In_1343);
or U794 (N_794,In_11,In_645);
and U795 (N_795,In_904,In_1567);
nor U796 (N_796,In_870,In_326);
nor U797 (N_797,In_1678,In_353);
and U798 (N_798,In_672,In_484);
nand U799 (N_799,In_1386,In_1871);
and U800 (N_800,N_292,N_796);
or U801 (N_801,In_203,In_1863);
nand U802 (N_802,N_355,N_276);
xnor U803 (N_803,In_234,In_1146);
nand U804 (N_804,N_312,N_176);
or U805 (N_805,N_44,N_373);
or U806 (N_806,N_559,N_158);
and U807 (N_807,N_540,In_1360);
nand U808 (N_808,In_64,In_437);
and U809 (N_809,N_175,In_963);
or U810 (N_810,N_127,In_87);
and U811 (N_811,In_134,N_297);
xor U812 (N_812,In_822,N_224);
nor U813 (N_813,N_742,In_1193);
and U814 (N_814,N_74,N_741);
nor U815 (N_815,In_767,N_12);
nor U816 (N_816,N_246,In_1131);
nand U817 (N_817,In_20,N_159);
and U818 (N_818,In_591,N_782);
nor U819 (N_819,In_683,N_442);
nor U820 (N_820,In_1297,In_1794);
xnor U821 (N_821,N_756,In_842);
or U822 (N_822,N_364,N_139);
xor U823 (N_823,N_567,N_20);
and U824 (N_824,N_258,N_481);
nor U825 (N_825,N_681,In_1065);
and U826 (N_826,N_227,In_1737);
nor U827 (N_827,N_183,N_7);
nand U828 (N_828,N_223,In_1260);
nand U829 (N_829,N_541,In_362);
nand U830 (N_830,N_760,N_96);
or U831 (N_831,In_718,N_112);
or U832 (N_832,In_682,In_205);
nor U833 (N_833,In_1401,In_1847);
nand U834 (N_834,N_717,N_478);
or U835 (N_835,N_713,N_537);
or U836 (N_836,In_763,N_33);
or U837 (N_837,N_116,In_405);
nand U838 (N_838,N_59,In_732);
nand U839 (N_839,In_295,In_1061);
xor U840 (N_840,N_456,N_173);
xnor U841 (N_841,In_1875,N_293);
and U842 (N_842,In_986,In_1277);
nand U843 (N_843,In_1658,N_288);
and U844 (N_844,N_745,N_539);
nand U845 (N_845,N_311,In_1797);
or U846 (N_846,N_450,N_383);
nand U847 (N_847,N_122,N_425);
or U848 (N_848,In_1129,N_716);
or U849 (N_849,N_445,N_668);
nand U850 (N_850,N_273,N_707);
nand U851 (N_851,In_401,N_595);
xor U852 (N_852,N_396,N_734);
nor U853 (N_853,N_566,In_192);
nor U854 (N_854,N_181,N_169);
and U855 (N_855,N_198,N_51);
and U856 (N_856,N_697,In_932);
and U857 (N_857,N_665,N_502);
nand U858 (N_858,N_687,N_405);
and U859 (N_859,N_317,In_1141);
and U860 (N_860,In_1542,In_1094);
xnor U861 (N_861,In_1053,N_672);
nor U862 (N_862,In_689,N_339);
nand U863 (N_863,In_494,N_550);
or U864 (N_864,In_289,In_1941);
nand U865 (N_865,N_131,In_1745);
xnor U866 (N_866,In_43,N_324);
nand U867 (N_867,In_480,N_469);
or U868 (N_868,N_392,N_432);
nand U869 (N_869,N_367,N_157);
nor U870 (N_870,N_272,In_1577);
and U871 (N_871,N_786,In_1361);
nor U872 (N_872,In_1003,N_107);
xnor U873 (N_873,In_1118,N_798);
nor U874 (N_874,N_100,In_895);
and U875 (N_875,N_363,N_499);
xnor U876 (N_876,N_587,In_869);
nand U877 (N_877,N_45,N_576);
and U878 (N_878,N_77,N_82);
nand U879 (N_879,In_130,In_872);
or U880 (N_880,N_408,N_757);
nand U881 (N_881,In_309,N_667);
and U882 (N_882,N_736,In_1058);
nand U883 (N_883,N_421,N_692);
nor U884 (N_884,In_1990,In_145);
nand U885 (N_885,N_623,In_638);
or U886 (N_886,N_36,N_728);
nand U887 (N_887,In_571,In_996);
nor U888 (N_888,N_19,N_635);
nor U889 (N_889,N_343,N_261);
and U890 (N_890,N_18,In_1983);
nor U891 (N_891,N_705,In_587);
xor U892 (N_892,N_369,N_301);
or U893 (N_893,N_221,N_578);
and U894 (N_894,N_605,N_362);
nand U895 (N_895,N_72,N_477);
and U896 (N_896,N_91,In_1574);
xnor U897 (N_897,In_752,N_138);
and U898 (N_898,In_22,In_1431);
nor U899 (N_899,N_585,N_265);
nand U900 (N_900,N_586,N_126);
xnor U901 (N_901,N_360,In_1499);
and U902 (N_902,In_346,N_551);
xor U903 (N_903,N_626,N_243);
nor U904 (N_904,N_193,N_303);
nand U905 (N_905,N_233,N_275);
or U906 (N_906,N_712,N_331);
nor U907 (N_907,N_632,In_1632);
nor U908 (N_908,N_443,N_535);
xor U909 (N_909,N_655,In_1270);
xnor U910 (N_910,N_380,In_1205);
xor U911 (N_911,In_527,In_537);
xnor U912 (N_912,In_1232,N_588);
xnor U913 (N_913,In_794,N_67);
nand U914 (N_914,In_1661,N_103);
or U915 (N_915,N_571,In_388);
nor U916 (N_916,In_324,In_301);
or U917 (N_917,In_1960,N_4);
nand U918 (N_918,N_350,N_155);
and U919 (N_919,N_503,N_685);
xnor U920 (N_920,N_57,In_667);
xor U921 (N_921,N_310,N_229);
and U922 (N_922,N_444,N_524);
nand U923 (N_923,N_748,In_1563);
nand U924 (N_924,N_49,N_73);
or U925 (N_925,N_108,N_746);
xnor U926 (N_926,N_9,N_270);
nand U927 (N_927,N_621,N_743);
nand U928 (N_928,N_87,N_81);
nor U929 (N_929,N_110,N_562);
and U930 (N_930,N_279,In_311);
and U931 (N_931,In_416,In_642);
nor U932 (N_932,N_622,N_326);
or U933 (N_933,In_559,In_1117);
or U934 (N_934,In_75,In_1857);
xor U935 (N_935,N_767,N_698);
nand U936 (N_936,N_530,In_1514);
or U937 (N_937,N_708,N_128);
nand U938 (N_938,In_1393,In_1936);
or U939 (N_939,N_280,N_124);
or U940 (N_940,In_1511,In_1142);
or U941 (N_941,N_184,In_640);
or U942 (N_942,In_1017,N_231);
nand U943 (N_943,In_1163,In_347);
nand U944 (N_944,N_93,N_686);
nor U945 (N_945,N_31,N_506);
nor U946 (N_946,N_168,N_426);
nor U947 (N_947,In_1221,In_928);
and U948 (N_948,In_95,N_35);
xor U949 (N_949,N_149,In_168);
nand U950 (N_950,In_817,N_309);
nor U951 (N_951,N_307,N_200);
nand U952 (N_952,N_141,N_511);
nor U953 (N_953,N_454,N_345);
xor U954 (N_954,In_1600,In_725);
xnor U955 (N_955,N_777,N_8);
nor U956 (N_956,In_252,In_1854);
or U957 (N_957,N_412,N_23);
and U958 (N_958,N_483,N_232);
or U959 (N_959,In_1450,N_531);
or U960 (N_960,N_269,N_165);
nor U961 (N_961,N_484,N_661);
nor U962 (N_962,In_396,N_519);
xnor U963 (N_963,N_447,N_439);
and U964 (N_964,N_402,N_218);
xor U965 (N_965,In_248,N_613);
xor U966 (N_966,In_562,N_285);
nor U967 (N_967,In_460,N_298);
and U968 (N_968,N_673,N_780);
or U969 (N_969,N_646,N_291);
xnor U970 (N_970,In_1153,N_267);
and U971 (N_971,N_98,N_147);
nor U972 (N_972,N_117,In_724);
and U973 (N_973,N_446,N_762);
or U974 (N_974,N_654,N_105);
xor U975 (N_975,N_300,In_819);
or U976 (N_976,In_30,N_625);
nand U977 (N_977,N_163,In_1730);
xnor U978 (N_978,N_83,In_1432);
xnor U979 (N_979,N_631,N_467);
nor U980 (N_980,N_55,N_489);
and U981 (N_981,N_68,In_1264);
and U982 (N_982,In_572,In_712);
and U983 (N_983,In_674,In_1039);
nor U984 (N_984,N_664,N_114);
xnor U985 (N_985,In_968,In_1459);
xnor U986 (N_986,In_31,N_744);
and U987 (N_987,N_793,In_56);
nand U988 (N_988,N_66,In_522);
xnor U989 (N_989,N_212,In_120);
xor U990 (N_990,In_1049,In_750);
nor U991 (N_991,N_755,N_709);
xor U992 (N_992,N_507,N_29);
or U993 (N_993,N_774,In_654);
or U994 (N_994,N_694,N_594);
xor U995 (N_995,N_255,N_287);
nand U996 (N_996,N_334,N_188);
nand U997 (N_997,In_34,N_710);
nand U998 (N_998,N_409,In_138);
and U999 (N_999,In_176,N_637);
nor U1000 (N_1000,In_1328,In_1978);
nor U1001 (N_1001,N_118,N_735);
xor U1002 (N_1002,In_1497,N_241);
nand U1003 (N_1003,N_335,N_466);
nor U1004 (N_1004,N_38,N_239);
and U1005 (N_1005,In_1817,N_753);
nor U1006 (N_1006,N_185,In_316);
xnor U1007 (N_1007,N_565,N_611);
nand U1008 (N_1008,N_281,In_1879);
and U1009 (N_1009,N_682,In_1736);
or U1010 (N_1010,In_731,N_388);
or U1011 (N_1011,In_679,In_1732);
or U1012 (N_1012,N_28,N_620);
nand U1013 (N_1013,N_453,N_352);
nand U1014 (N_1014,In_707,N_278);
nand U1015 (N_1015,N_513,N_737);
xor U1016 (N_1016,In_601,In_708);
or U1017 (N_1017,N_50,N_644);
xor U1018 (N_1018,N_171,In_1591);
nand U1019 (N_1019,In_1523,N_479);
xnor U1020 (N_1020,In_1225,N_572);
nand U1021 (N_1021,In_720,In_1128);
or U1022 (N_1022,N_764,N_53);
nand U1023 (N_1023,N_358,N_336);
nand U1024 (N_1024,N_492,N_21);
or U1025 (N_1025,In_700,N_527);
xnor U1026 (N_1026,In_302,N_451);
or U1027 (N_1027,In_1283,N_95);
or U1028 (N_1028,In_668,N_553);
and U1029 (N_1029,N_459,In_1575);
xnor U1030 (N_1030,N_113,N_340);
xor U1031 (N_1031,N_619,In_333);
nor U1032 (N_1032,N_749,N_216);
or U1033 (N_1033,In_584,N_156);
or U1034 (N_1034,N_257,N_154);
and U1035 (N_1035,In_368,N_384);
nor U1036 (N_1036,N_570,In_196);
or U1037 (N_1037,N_522,N_704);
or U1038 (N_1038,N_468,N_612);
xor U1039 (N_1039,N_252,N_13);
nor U1040 (N_1040,In_1708,In_159);
or U1041 (N_1041,N_333,N_251);
and U1042 (N_1042,N_617,N_508);
nor U1043 (N_1043,In_1416,In_1443);
nor U1044 (N_1044,N_164,In_793);
and U1045 (N_1045,N_415,N_313);
nor U1046 (N_1046,N_370,In_239);
nand U1047 (N_1047,N_268,N_220);
xor U1048 (N_1048,N_423,N_690);
xnor U1049 (N_1049,N_377,N_560);
nor U1050 (N_1050,In_468,N_341);
nor U1051 (N_1051,In_576,N_548);
nand U1052 (N_1052,N_14,In_197);
and U1053 (N_1053,N_441,N_574);
nand U1054 (N_1054,N_320,In_1843);
and U1055 (N_1055,In_106,N_614);
xnor U1056 (N_1056,N_486,N_607);
nand U1057 (N_1057,N_327,N_234);
xnor U1058 (N_1058,N_102,N_294);
and U1059 (N_1059,N_675,In_1305);
or U1060 (N_1060,N_608,N_526);
or U1061 (N_1061,N_491,N_202);
nor U1062 (N_1062,N_581,N_778);
nor U1063 (N_1063,N_792,In_114);
xor U1064 (N_1064,N_775,In_1285);
xor U1065 (N_1065,N_214,N_356);
nor U1066 (N_1066,In_999,In_201);
nand U1067 (N_1067,N_648,In_1726);
and U1068 (N_1068,N_591,N_187);
nand U1069 (N_1069,In_900,N_199);
nor U1070 (N_1070,In_776,N_794);
nor U1071 (N_1071,In_288,In_1578);
nor U1072 (N_1072,N_344,In_1646);
xnor U1073 (N_1073,N_399,N_497);
xor U1074 (N_1074,N_235,N_25);
and U1075 (N_1075,N_465,N_589);
nor U1076 (N_1076,In_951,N_386);
nor U1077 (N_1077,N_706,N_30);
nand U1078 (N_1078,In_510,N_427);
nor U1079 (N_1079,N_422,N_43);
xor U1080 (N_1080,In_1688,In_1436);
xor U1081 (N_1081,In_499,N_606);
nand U1082 (N_1082,N_573,N_547);
nor U1083 (N_1083,In_1154,N_514);
nand U1084 (N_1084,N_366,In_208);
xnor U1085 (N_1085,N_6,In_1449);
nor U1086 (N_1086,In_1535,N_207);
and U1087 (N_1087,N_795,In_113);
nor U1088 (N_1088,In_1419,In_1468);
and U1089 (N_1089,N_740,N_61);
nor U1090 (N_1090,N_776,N_410);
nand U1091 (N_1091,In_74,In_1536);
and U1092 (N_1092,N_10,N_659);
or U1093 (N_1093,N_765,In_363);
nor U1094 (N_1094,N_784,N_129);
xnor U1095 (N_1095,N_747,In_736);
nand U1096 (N_1096,In_161,In_1751);
nand U1097 (N_1097,In_1715,N_245);
nor U1098 (N_1098,N_516,N_691);
xor U1099 (N_1099,In_115,In_1618);
nand U1100 (N_1100,N_462,N_599);
xor U1101 (N_1101,In_53,In_379);
or U1102 (N_1102,N_119,N_474);
xor U1103 (N_1103,N_97,N_330);
nor U1104 (N_1104,N_517,In_336);
and U1105 (N_1105,In_1778,In_1215);
and U1106 (N_1106,N_161,N_378);
and U1107 (N_1107,N_282,In_304);
xor U1108 (N_1108,N_437,N_152);
and U1109 (N_1109,N_27,N_46);
and U1110 (N_1110,N_429,N_347);
nand U1111 (N_1111,In_1372,N_99);
nor U1112 (N_1112,N_394,N_418);
and U1113 (N_1113,N_37,N_393);
xnor U1114 (N_1114,N_733,N_144);
nor U1115 (N_1115,N_449,N_580);
and U1116 (N_1116,In_575,N_799);
nand U1117 (N_1117,N_348,N_398);
or U1118 (N_1118,In_615,N_52);
or U1119 (N_1119,In_1160,N_106);
xnor U1120 (N_1120,N_538,N_177);
nand U1121 (N_1121,In_1390,In_345);
nor U1122 (N_1122,In_1059,N_375);
and U1123 (N_1123,N_662,N_306);
or U1124 (N_1124,N_5,N_299);
or U1125 (N_1125,N_47,N_598);
and U1126 (N_1126,N_236,N_361);
xor U1127 (N_1127,N_521,In_1392);
or U1128 (N_1128,N_457,In_1779);
nor U1129 (N_1129,N_332,N_461);
nor U1130 (N_1130,N_274,N_650);
or U1131 (N_1131,N_554,N_219);
nor U1132 (N_1132,In_71,In_747);
nor U1133 (N_1133,In_1492,In_813);
nor U1134 (N_1134,N_0,N_670);
and U1135 (N_1135,In_539,N_463);
xor U1136 (N_1136,In_1543,N_208);
or U1137 (N_1137,In_255,In_655);
and U1138 (N_1138,In_453,In_1262);
and U1139 (N_1139,N_250,N_663);
nor U1140 (N_1140,N_711,In_1056);
xor U1141 (N_1141,In_116,In_1830);
nand U1142 (N_1142,N_135,N_259);
xnor U1143 (N_1143,In_1754,In_500);
and U1144 (N_1144,In_836,N_761);
or U1145 (N_1145,In_1172,N_487);
or U1146 (N_1146,In_1303,N_374);
or U1147 (N_1147,N_379,N_151);
or U1148 (N_1148,In_442,N_592);
xnor U1149 (N_1149,In_98,In_246);
nand U1150 (N_1150,N_726,N_153);
xnor U1151 (N_1151,N_94,In_1479);
nand U1152 (N_1152,N_568,N_115);
nand U1153 (N_1153,In_1211,N_172);
nand U1154 (N_1154,N_525,N_739);
nor U1155 (N_1155,In_1791,In_1593);
nand U1156 (N_1156,N_440,In_1939);
and U1157 (N_1157,In_487,N_316);
nor U1158 (N_1158,N_354,N_143);
nand U1159 (N_1159,N_88,In_1476);
nand U1160 (N_1160,N_215,In_1251);
nand U1161 (N_1161,N_501,N_204);
or U1162 (N_1162,In_1485,In_226);
or U1163 (N_1163,N_78,In_621);
or U1164 (N_1164,In_439,N_69);
or U1165 (N_1165,N_48,N_575);
and U1166 (N_1166,N_84,N_564);
nor U1167 (N_1167,N_249,N_600);
xnor U1168 (N_1168,N_438,In_1501);
nand U1169 (N_1169,N_750,N_387);
xnor U1170 (N_1170,N_797,N_189);
nor U1171 (N_1171,N_719,In_1494);
and U1172 (N_1172,In_1853,N_630);
and U1173 (N_1173,In_1572,In_846);
or U1174 (N_1174,N_640,In_1115);
or U1175 (N_1175,N_264,N_315);
and U1176 (N_1176,N_111,N_390);
xor U1177 (N_1177,N_222,N_528);
nand U1178 (N_1178,N_533,N_2);
nand U1179 (N_1179,In_135,N_684);
nor U1180 (N_1180,N_385,N_217);
nand U1181 (N_1181,N_130,In_1870);
xor U1182 (N_1182,In_419,In_1242);
nand U1183 (N_1183,In_1385,N_322);
nor U1184 (N_1184,N_556,N_63);
and U1185 (N_1185,N_56,N_160);
and U1186 (N_1186,In_595,N_593);
nor U1187 (N_1187,N_314,N_346);
nor U1188 (N_1188,In_676,In_1586);
nor U1189 (N_1189,N_201,N_123);
nand U1190 (N_1190,N_419,N_638);
or U1191 (N_1191,In_254,N_256);
or U1192 (N_1192,N_543,N_357);
xor U1193 (N_1193,N_791,In_1584);
xor U1194 (N_1194,N_558,N_17);
and U1195 (N_1195,N_496,N_542);
xnor U1196 (N_1196,N_70,In_898);
and U1197 (N_1197,N_253,N_420);
xor U1198 (N_1198,N_407,In_465);
xor U1199 (N_1199,N_395,N_101);
and U1200 (N_1200,N_561,N_406);
and U1201 (N_1201,N_783,N_683);
xor U1202 (N_1202,In_412,In_172);
or U1203 (N_1203,N_597,N_510);
nor U1204 (N_1204,N_41,N_460);
nand U1205 (N_1205,N_604,N_166);
xnor U1206 (N_1206,N_602,N_549);
and U1207 (N_1207,N_472,N_651);
or U1208 (N_1208,N_656,In_189);
nand U1209 (N_1209,N_178,In_1444);
nor U1210 (N_1210,In_843,N_338);
and U1211 (N_1211,N_428,N_65);
xnor U1212 (N_1212,N_162,N_475);
xnor U1213 (N_1213,N_353,N_544);
or U1214 (N_1214,N_430,N_195);
or U1215 (N_1215,N_688,N_520);
nor U1216 (N_1216,N_186,In_1687);
nand U1217 (N_1217,N_579,N_752);
or U1218 (N_1218,N_197,N_596);
nand U1219 (N_1219,N_295,N_308);
nand U1220 (N_1220,N_464,N_639);
or U1221 (N_1221,N_495,N_342);
and U1222 (N_1222,N_509,N_391);
xor U1223 (N_1223,In_1060,N_436);
nor U1224 (N_1224,N_205,N_779);
or U1225 (N_1225,In_411,N_376);
or U1226 (N_1226,N_699,N_788);
nor U1227 (N_1227,N_194,N_125);
nand U1228 (N_1228,In_1825,In_504);
or U1229 (N_1229,N_676,N_590);
nand U1230 (N_1230,In_508,N_727);
or U1231 (N_1231,N_660,N_54);
nand U1232 (N_1232,N_413,In_1493);
xnor U1233 (N_1233,N_240,N_624);
xnor U1234 (N_1234,In_1407,In_1177);
xor U1235 (N_1235,In_774,In_1063);
or U1236 (N_1236,N_518,N_39);
or U1237 (N_1237,N_381,N_226);
or U1238 (N_1238,N_79,N_225);
xnor U1239 (N_1239,N_262,N_414);
xnor U1240 (N_1240,N_601,N_787);
or U1241 (N_1241,N_657,N_254);
or U1242 (N_1242,N_473,N_633);
xnor U1243 (N_1243,In_1828,N_206);
nor U1244 (N_1244,In_359,N_180);
nand U1245 (N_1245,N_417,N_546);
xnor U1246 (N_1246,N_758,In_282);
xor U1247 (N_1247,In_238,N_433);
nor U1248 (N_1248,In_1026,In_1582);
xor U1249 (N_1249,N_763,In_422);
xor U1250 (N_1250,N_584,N_552);
xnor U1251 (N_1251,N_493,N_58);
nand U1252 (N_1252,N_244,In_961);
xnor U1253 (N_1253,N_329,N_636);
nand U1254 (N_1254,In_387,In_222);
and U1255 (N_1255,In_1337,In_742);
xor U1256 (N_1256,N_629,N_722);
nor U1257 (N_1257,In_331,N_669);
nand U1258 (N_1258,N_615,In_93);
xnor U1259 (N_1259,N_210,In_588);
nand U1260 (N_1260,In_1573,In_823);
or U1261 (N_1261,N_754,N_40);
and U1262 (N_1262,N_470,In_586);
xor U1263 (N_1263,N_693,N_137);
and U1264 (N_1264,In_1157,N_15);
and U1265 (N_1265,N_71,In_592);
nor U1266 (N_1266,N_731,N_721);
nor U1267 (N_1267,N_536,In_300);
xnor U1268 (N_1268,In_1447,N_191);
nor U1269 (N_1269,N_11,In_1695);
or U1270 (N_1270,In_492,N_494);
and U1271 (N_1271,In_702,In_92);
nand U1272 (N_1272,N_720,N_109);
and U1273 (N_1273,In_737,In_69);
xor U1274 (N_1274,N_62,N_237);
nor U1275 (N_1275,N_248,N_700);
nand U1276 (N_1276,N_136,N_321);
xor U1277 (N_1277,In_299,In_41);
nand U1278 (N_1278,N_290,N_416);
xnor U1279 (N_1279,N_368,In_739);
nand U1280 (N_1280,N_577,N_678);
or U1281 (N_1281,N_401,N_382);
nand U1282 (N_1282,In_666,N_653);
xnor U1283 (N_1283,N_555,In_1818);
and U1284 (N_1284,In_1915,N_397);
and U1285 (N_1285,N_729,In_1813);
nor U1286 (N_1286,N_349,N_609);
nor U1287 (N_1287,N_523,In_787);
and U1288 (N_1288,In_483,In_1356);
xnor U1289 (N_1289,N_458,N_790);
nand U1290 (N_1290,N_271,In_179);
nand U1291 (N_1291,N_730,N_260);
and U1292 (N_1292,N_480,N_167);
xor U1293 (N_1293,N_150,N_674);
or U1294 (N_1294,N_545,N_174);
and U1295 (N_1295,N_610,N_411);
nand U1296 (N_1296,N_86,In_1997);
xnor U1297 (N_1297,In_382,N_723);
nor U1298 (N_1298,In_1400,In_1208);
xnor U1299 (N_1299,N_142,N_789);
xor U1300 (N_1300,N_677,N_715);
and U1301 (N_1301,N_634,N_714);
nand U1302 (N_1302,N_323,N_359);
xor U1303 (N_1303,N_121,In_1682);
and U1304 (N_1304,In_713,In_1755);
xor U1305 (N_1305,N_424,In_121);
or U1306 (N_1306,N_192,N_647);
or U1307 (N_1307,N_725,N_104);
nor U1308 (N_1308,N_196,In_540);
or U1309 (N_1309,N_64,N_781);
and U1310 (N_1310,N_148,In_1698);
nor U1311 (N_1311,N_32,N_696);
nand U1312 (N_1312,N_179,N_703);
xor U1313 (N_1313,N_228,In_989);
nand U1314 (N_1314,N_371,N_400);
xor U1315 (N_1315,In_538,N_488);
or U1316 (N_1316,In_219,N_768);
or U1317 (N_1317,In_1472,In_46);
nor U1318 (N_1318,In_1991,N_140);
nand U1319 (N_1319,N_732,In_1106);
nor U1320 (N_1320,N_145,N_485);
nor U1321 (N_1321,N_771,N_582);
nor U1322 (N_1322,N_627,N_652);
xnor U1323 (N_1323,N_351,N_773);
nor U1324 (N_1324,In_1034,N_238);
nor U1325 (N_1325,N_512,N_263);
xor U1326 (N_1326,In_1605,N_146);
xnor U1327 (N_1327,N_557,N_24);
nand U1328 (N_1328,N_500,N_286);
nor U1329 (N_1329,N_641,N_26);
and U1330 (N_1330,In_1457,In_768);
xor U1331 (N_1331,In_1627,In_942);
and U1332 (N_1332,In_1010,N_247);
and U1333 (N_1333,N_89,N_618);
xnor U1334 (N_1334,In_1158,N_318);
nand U1335 (N_1335,N_515,N_190);
or U1336 (N_1336,N_289,In_1856);
and U1337 (N_1337,N_770,In_1433);
or U1338 (N_1338,N_759,N_404);
nand U1339 (N_1339,N_452,N_3);
nand U1340 (N_1340,N_434,N_435);
and U1341 (N_1341,N_304,In_1806);
and U1342 (N_1342,N_645,In_512);
nand U1343 (N_1343,N_724,N_85);
xor U1344 (N_1344,N_448,In_1800);
nor U1345 (N_1345,N_319,N_403);
xnor U1346 (N_1346,N_76,N_642);
nand U1347 (N_1347,N_671,N_120);
xnor U1348 (N_1348,N_666,N_658);
nor U1349 (N_1349,N_302,N_772);
xor U1350 (N_1350,N_490,N_296);
xnor U1351 (N_1351,N_680,N_42);
nor U1352 (N_1352,In_1454,In_1033);
or U1353 (N_1353,N_209,N_628);
xnor U1354 (N_1354,N_182,N_337);
nor U1355 (N_1355,N_211,In_1814);
nor U1356 (N_1356,In_1910,In_798);
nor U1357 (N_1357,In_1894,N_679);
and U1358 (N_1358,N_325,N_242);
and U1359 (N_1359,N_431,N_213);
and U1360 (N_1360,In_1581,In_1580);
nor U1361 (N_1361,N_284,N_583);
nor U1362 (N_1362,In_984,N_75);
nand U1363 (N_1363,N_134,N_203);
and U1364 (N_1364,In_1092,In_1195);
and U1365 (N_1365,N_643,N_689);
nor U1366 (N_1366,In_217,N_534);
or U1367 (N_1367,N_738,In_614);
nand U1368 (N_1368,N_305,N_92);
xnor U1369 (N_1369,N_132,N_389);
xnor U1370 (N_1370,In_1124,In_1378);
and U1371 (N_1371,N_60,N_455);
nor U1372 (N_1372,N_751,N_498);
nor U1373 (N_1373,N_532,N_482);
or U1374 (N_1374,In_1764,N_16);
nor U1375 (N_1375,N_476,N_230);
and U1376 (N_1376,N_563,N_769);
and U1377 (N_1377,N_766,N_1);
xnor U1378 (N_1378,In_160,In_280);
xor U1379 (N_1379,N_283,N_649);
xor U1380 (N_1380,N_695,N_471);
nand U1381 (N_1381,In_806,In_1583);
or U1382 (N_1382,In_303,N_277);
nand U1383 (N_1383,N_505,In_478);
or U1384 (N_1384,N_266,In_496);
and U1385 (N_1385,N_702,In_1036);
nand U1386 (N_1386,N_529,In_237);
nand U1387 (N_1387,N_701,In_1947);
or U1388 (N_1388,N_22,In_1315);
xor U1389 (N_1389,In_1483,N_170);
and U1390 (N_1390,In_330,N_718);
xor U1391 (N_1391,N_616,N_80);
nor U1392 (N_1392,N_372,In_509);
nor U1393 (N_1393,N_365,In_1366);
and U1394 (N_1394,N_603,In_1942);
nor U1395 (N_1395,In_662,N_569);
or U1396 (N_1396,N_90,N_133);
nor U1397 (N_1397,N_504,N_328);
xor U1398 (N_1398,N_785,In_1108);
and U1399 (N_1399,In_49,N_34);
or U1400 (N_1400,N_124,N_458);
and U1401 (N_1401,N_716,In_1315);
nand U1402 (N_1402,In_1303,In_1154);
nand U1403 (N_1403,In_1581,N_186);
xnor U1404 (N_1404,In_494,In_900);
nor U1405 (N_1405,N_723,In_324);
or U1406 (N_1406,In_1493,N_100);
and U1407 (N_1407,In_201,N_64);
xor U1408 (N_1408,In_192,N_250);
and U1409 (N_1409,In_794,In_1960);
nor U1410 (N_1410,N_305,N_264);
or U1411 (N_1411,In_226,In_1828);
nor U1412 (N_1412,In_1328,N_2);
and U1413 (N_1413,N_390,N_565);
and U1414 (N_1414,N_392,N_351);
or U1415 (N_1415,N_297,In_439);
or U1416 (N_1416,N_127,N_752);
nor U1417 (N_1417,N_322,In_1450);
xnor U1418 (N_1418,N_335,N_291);
or U1419 (N_1419,N_651,N_621);
nor U1420 (N_1420,N_213,N_541);
nand U1421 (N_1421,In_586,N_412);
nor U1422 (N_1422,N_72,N_33);
nand U1423 (N_1423,N_616,N_70);
nand U1424 (N_1424,N_744,N_616);
nor U1425 (N_1425,N_416,N_207);
xor U1426 (N_1426,In_712,N_433);
or U1427 (N_1427,N_601,N_731);
nor U1428 (N_1428,N_30,In_900);
nand U1429 (N_1429,N_748,N_150);
xnor U1430 (N_1430,N_279,In_1017);
or U1431 (N_1431,N_626,In_43);
and U1432 (N_1432,N_346,In_1572);
and U1433 (N_1433,N_545,N_442);
or U1434 (N_1434,N_365,In_928);
nand U1435 (N_1435,In_282,N_447);
and U1436 (N_1436,N_764,N_663);
nor U1437 (N_1437,N_72,N_417);
or U1438 (N_1438,N_86,N_453);
nor U1439 (N_1439,N_152,In_1941);
or U1440 (N_1440,In_1806,In_1581);
nor U1441 (N_1441,N_116,In_591);
nor U1442 (N_1442,N_200,N_744);
nand U1443 (N_1443,N_394,In_662);
xnor U1444 (N_1444,N_461,N_477);
or U1445 (N_1445,N_300,In_654);
or U1446 (N_1446,In_331,N_80);
xnor U1447 (N_1447,In_1447,N_65);
nor U1448 (N_1448,In_487,N_494);
nand U1449 (N_1449,N_709,In_817);
nand U1450 (N_1450,N_669,N_736);
or U1451 (N_1451,N_245,In_1242);
or U1452 (N_1452,N_215,N_522);
nand U1453 (N_1453,N_109,N_193);
or U1454 (N_1454,In_1584,In_1251);
xor U1455 (N_1455,N_645,In_1436);
xnor U1456 (N_1456,N_30,N_349);
or U1457 (N_1457,N_414,N_552);
or U1458 (N_1458,In_145,N_399);
nor U1459 (N_1459,In_1297,N_232);
xor U1460 (N_1460,N_48,In_504);
or U1461 (N_1461,N_426,In_1535);
xor U1462 (N_1462,N_190,In_336);
and U1463 (N_1463,N_437,In_1737);
nor U1464 (N_1464,N_459,N_48);
or U1465 (N_1465,N_272,N_580);
or U1466 (N_1466,In_1501,N_443);
nor U1467 (N_1467,In_1941,In_248);
nand U1468 (N_1468,In_537,N_307);
xnor U1469 (N_1469,N_678,N_74);
nand U1470 (N_1470,N_526,N_438);
or U1471 (N_1471,N_693,N_692);
nand U1472 (N_1472,N_246,N_160);
or U1473 (N_1473,N_317,In_1942);
nor U1474 (N_1474,In_1806,N_93);
or U1475 (N_1475,N_700,In_989);
and U1476 (N_1476,N_734,N_565);
nor U1477 (N_1477,N_569,N_447);
nor U1478 (N_1478,In_1225,N_774);
nor U1479 (N_1479,In_872,In_584);
nor U1480 (N_1480,N_601,N_48);
nor U1481 (N_1481,N_159,N_424);
nor U1482 (N_1482,N_756,N_668);
or U1483 (N_1483,In_330,In_591);
nand U1484 (N_1484,N_8,N_143);
or U1485 (N_1485,N_82,In_819);
and U1486 (N_1486,N_219,N_346);
nor U1487 (N_1487,In_1997,In_192);
and U1488 (N_1488,N_603,N_387);
or U1489 (N_1489,N_57,N_761);
xnor U1490 (N_1490,N_515,In_724);
or U1491 (N_1491,N_609,In_1983);
nand U1492 (N_1492,N_78,In_707);
or U1493 (N_1493,N_236,N_408);
xor U1494 (N_1494,N_736,N_425);
or U1495 (N_1495,N_637,N_42);
nor U1496 (N_1496,N_149,N_510);
nor U1497 (N_1497,N_281,In_731);
nand U1498 (N_1498,In_1034,In_1141);
nor U1499 (N_1499,N_382,N_490);
nand U1500 (N_1500,N_208,N_93);
or U1501 (N_1501,In_382,N_415);
xnor U1502 (N_1502,N_344,In_87);
nand U1503 (N_1503,N_365,N_524);
or U1504 (N_1504,In_500,N_523);
nand U1505 (N_1505,In_584,N_483);
and U1506 (N_1506,N_508,N_408);
nor U1507 (N_1507,In_254,N_32);
and U1508 (N_1508,N_695,In_575);
or U1509 (N_1509,N_445,N_263);
nor U1510 (N_1510,N_715,N_255);
nor U1511 (N_1511,In_460,N_380);
xor U1512 (N_1512,In_161,In_1843);
xor U1513 (N_1513,N_494,N_55);
nand U1514 (N_1514,In_179,In_1575);
and U1515 (N_1515,N_76,N_203);
or U1516 (N_1516,N_663,N_354);
or U1517 (N_1517,N_102,N_595);
nor U1518 (N_1518,In_1600,N_671);
nor U1519 (N_1519,N_492,N_585);
nand U1520 (N_1520,In_1857,N_296);
or U1521 (N_1521,In_362,In_176);
or U1522 (N_1522,In_731,N_546);
nand U1523 (N_1523,N_626,In_106);
xor U1524 (N_1524,N_384,N_558);
nand U1525 (N_1525,N_587,N_378);
or U1526 (N_1526,In_160,N_122);
nand U1527 (N_1527,N_270,N_714);
nor U1528 (N_1528,In_999,N_745);
nor U1529 (N_1529,In_747,N_236);
nor U1530 (N_1530,N_103,In_932);
and U1531 (N_1531,N_40,N_708);
xor U1532 (N_1532,In_1514,N_418);
or U1533 (N_1533,N_742,N_349);
or U1534 (N_1534,In_1936,In_43);
or U1535 (N_1535,In_1755,In_750);
and U1536 (N_1536,N_411,N_717);
xor U1537 (N_1537,N_657,In_379);
xor U1538 (N_1538,N_187,In_1578);
nand U1539 (N_1539,N_643,N_756);
or U1540 (N_1540,N_264,N_419);
nor U1541 (N_1541,N_232,N_526);
and U1542 (N_1542,N_371,N_518);
xor U1543 (N_1543,In_1910,N_348);
nand U1544 (N_1544,N_780,N_639);
and U1545 (N_1545,N_625,N_730);
xnor U1546 (N_1546,In_1337,N_301);
or U1547 (N_1547,In_331,In_679);
nand U1548 (N_1548,N_457,In_540);
and U1549 (N_1549,N_671,N_642);
nand U1550 (N_1550,N_499,N_32);
and U1551 (N_1551,N_502,N_729);
xnor U1552 (N_1552,N_235,N_669);
nand U1553 (N_1553,N_771,N_201);
nor U1554 (N_1554,In_1450,In_1260);
nand U1555 (N_1555,N_679,N_717);
xor U1556 (N_1556,N_634,N_516);
nor U1557 (N_1557,N_444,In_737);
nand U1558 (N_1558,In_246,N_639);
or U1559 (N_1559,N_169,N_646);
xnor U1560 (N_1560,N_411,N_744);
or U1561 (N_1561,N_328,N_388);
nand U1562 (N_1562,N_779,In_737);
nand U1563 (N_1563,N_136,N_653);
nand U1564 (N_1564,N_189,In_559);
nor U1565 (N_1565,N_718,N_226);
and U1566 (N_1566,N_466,N_768);
and U1567 (N_1567,N_34,N_321);
nor U1568 (N_1568,In_640,N_305);
and U1569 (N_1569,N_170,In_396);
nand U1570 (N_1570,In_1053,N_5);
nand U1571 (N_1571,In_1337,N_546);
or U1572 (N_1572,N_710,N_593);
or U1573 (N_1573,N_104,In_1094);
nor U1574 (N_1574,N_22,N_450);
and U1575 (N_1575,N_749,In_1260);
nor U1576 (N_1576,N_694,In_1060);
nor U1577 (N_1577,In_1825,In_591);
nor U1578 (N_1578,N_266,In_331);
xor U1579 (N_1579,In_121,N_381);
nand U1580 (N_1580,In_527,N_403);
nand U1581 (N_1581,In_1661,In_823);
nor U1582 (N_1582,N_333,N_570);
xnor U1583 (N_1583,In_1492,In_575);
and U1584 (N_1584,N_754,N_718);
nand U1585 (N_1585,N_796,N_84);
xor U1586 (N_1586,N_706,N_219);
and U1587 (N_1587,N_161,In_1894);
nor U1588 (N_1588,In_679,N_679);
nor U1589 (N_1589,N_317,N_552);
nand U1590 (N_1590,N_465,In_1511);
nor U1591 (N_1591,N_323,N_536);
xnor U1592 (N_1592,N_727,N_730);
nor U1593 (N_1593,N_92,N_751);
and U1594 (N_1594,N_380,N_526);
nor U1595 (N_1595,N_516,In_1443);
xor U1596 (N_1596,In_562,In_968);
or U1597 (N_1597,N_354,N_332);
or U1598 (N_1598,N_489,N_92);
nor U1599 (N_1599,In_1847,N_342);
or U1600 (N_1600,N_1430,N_1255);
and U1601 (N_1601,N_1347,N_1489);
or U1602 (N_1602,N_1258,N_1356);
nor U1603 (N_1603,N_1394,N_873);
xnor U1604 (N_1604,N_1414,N_1573);
or U1605 (N_1605,N_1509,N_1057);
nand U1606 (N_1606,N_1273,N_1559);
nand U1607 (N_1607,N_1123,N_1235);
nand U1608 (N_1608,N_1391,N_1328);
nand U1609 (N_1609,N_840,N_1408);
nand U1610 (N_1610,N_918,N_838);
nor U1611 (N_1611,N_1493,N_1513);
nor U1612 (N_1612,N_1360,N_919);
xor U1613 (N_1613,N_1148,N_1240);
and U1614 (N_1614,N_1061,N_1449);
or U1615 (N_1615,N_1445,N_1253);
and U1616 (N_1616,N_916,N_935);
nand U1617 (N_1617,N_1369,N_1159);
xnor U1618 (N_1618,N_1309,N_959);
nor U1619 (N_1619,N_1045,N_1434);
xor U1620 (N_1620,N_1571,N_848);
nand U1621 (N_1621,N_882,N_809);
and U1622 (N_1622,N_1024,N_1036);
nor U1623 (N_1623,N_931,N_989);
or U1624 (N_1624,N_1259,N_992);
or U1625 (N_1625,N_962,N_846);
xor U1626 (N_1626,N_1536,N_1237);
xnor U1627 (N_1627,N_1040,N_1247);
or U1628 (N_1628,N_859,N_965);
and U1629 (N_1629,N_1557,N_941);
and U1630 (N_1630,N_1000,N_829);
nor U1631 (N_1631,N_1260,N_908);
nand U1632 (N_1632,N_1572,N_1366);
xor U1633 (N_1633,N_1107,N_868);
xnor U1634 (N_1634,N_1568,N_1421);
xor U1635 (N_1635,N_1400,N_922);
or U1636 (N_1636,N_870,N_1083);
nand U1637 (N_1637,N_1500,N_1021);
nand U1638 (N_1638,N_1196,N_1043);
and U1639 (N_1639,N_1276,N_1348);
or U1640 (N_1640,N_1266,N_1218);
nand U1641 (N_1641,N_1238,N_1515);
nor U1642 (N_1642,N_1569,N_1062);
or U1643 (N_1643,N_1307,N_1297);
and U1644 (N_1644,N_807,N_1404);
or U1645 (N_1645,N_1225,N_1448);
and U1646 (N_1646,N_1130,N_1232);
or U1647 (N_1647,N_1129,N_936);
and U1648 (N_1648,N_1472,N_836);
nand U1649 (N_1649,N_1351,N_1467);
or U1650 (N_1650,N_1164,N_867);
xor U1651 (N_1651,N_1070,N_1383);
nor U1652 (N_1652,N_815,N_1466);
nor U1653 (N_1653,N_1533,N_843);
or U1654 (N_1654,N_1171,N_1189);
or U1655 (N_1655,N_1113,N_1188);
xnor U1656 (N_1656,N_1575,N_818);
or U1657 (N_1657,N_1398,N_1185);
or U1658 (N_1658,N_1461,N_1399);
xnor U1659 (N_1659,N_1127,N_1423);
nor U1660 (N_1660,N_1163,N_1243);
xnor U1661 (N_1661,N_1223,N_1352);
nand U1662 (N_1662,N_860,N_1574);
nand U1663 (N_1663,N_1162,N_1444);
nor U1664 (N_1664,N_1244,N_1068);
nor U1665 (N_1665,N_1194,N_1094);
and U1666 (N_1666,N_834,N_1395);
nand U1667 (N_1667,N_855,N_891);
or U1668 (N_1668,N_1169,N_1089);
or U1669 (N_1669,N_1455,N_1011);
or U1670 (N_1670,N_1405,N_1447);
nor U1671 (N_1671,N_827,N_1517);
nand U1672 (N_1672,N_1424,N_883);
xor U1673 (N_1673,N_1481,N_847);
or U1674 (N_1674,N_1268,N_949);
nor U1675 (N_1675,N_988,N_1242);
or U1676 (N_1676,N_1592,N_912);
or U1677 (N_1677,N_1246,N_1263);
or U1678 (N_1678,N_1510,N_960);
xor U1679 (N_1679,N_1279,N_1026);
nor U1680 (N_1680,N_1087,N_1006);
xor U1681 (N_1681,N_1217,N_1050);
and U1682 (N_1682,N_1155,N_1108);
or U1683 (N_1683,N_845,N_1302);
xor U1684 (N_1684,N_1310,N_1579);
or U1685 (N_1685,N_872,N_1211);
and U1686 (N_1686,N_1402,N_1300);
nand U1687 (N_1687,N_1137,N_1502);
and U1688 (N_1688,N_1042,N_1022);
and U1689 (N_1689,N_910,N_1413);
and U1690 (N_1690,N_1284,N_1009);
and U1691 (N_1691,N_1530,N_879);
nand U1692 (N_1692,N_886,N_1377);
or U1693 (N_1693,N_978,N_1554);
xor U1694 (N_1694,N_1082,N_1578);
nand U1695 (N_1695,N_850,N_964);
nand U1696 (N_1696,N_1028,N_1135);
nor U1697 (N_1697,N_1589,N_1295);
or U1698 (N_1698,N_1035,N_1521);
and U1699 (N_1699,N_1375,N_1522);
or U1700 (N_1700,N_1115,N_950);
xnor U1701 (N_1701,N_1272,N_1463);
nor U1702 (N_1702,N_1325,N_1512);
or U1703 (N_1703,N_1384,N_1261);
xnor U1704 (N_1704,N_1198,N_1373);
nor U1705 (N_1705,N_816,N_1374);
nand U1706 (N_1706,N_1140,N_924);
and U1707 (N_1707,N_1551,N_1496);
and U1708 (N_1708,N_1346,N_1345);
nor U1709 (N_1709,N_1560,N_1393);
xor U1710 (N_1710,N_1128,N_1588);
or U1711 (N_1711,N_975,N_1220);
or U1712 (N_1712,N_1074,N_1296);
xnor U1713 (N_1713,N_1367,N_1314);
nand U1714 (N_1714,N_812,N_1535);
and U1715 (N_1715,N_1230,N_1562);
and U1716 (N_1716,N_979,N_1044);
nand U1717 (N_1717,N_943,N_1204);
or U1718 (N_1718,N_1239,N_839);
nor U1719 (N_1719,N_997,N_1007);
nor U1720 (N_1720,N_1339,N_811);
and U1721 (N_1721,N_972,N_1060);
or U1722 (N_1722,N_1048,N_853);
xnor U1723 (N_1723,N_1165,N_1183);
nor U1724 (N_1724,N_1111,N_925);
nor U1725 (N_1725,N_933,N_1390);
or U1726 (N_1726,N_1321,N_932);
nor U1727 (N_1727,N_917,N_1553);
or U1728 (N_1728,N_1431,N_1208);
nor U1729 (N_1729,N_1432,N_1091);
and U1730 (N_1730,N_1590,N_974);
xor U1731 (N_1731,N_1598,N_1331);
and U1732 (N_1732,N_1547,N_1058);
or U1733 (N_1733,N_1166,N_1131);
nand U1734 (N_1734,N_1497,N_928);
nor U1735 (N_1735,N_874,N_929);
nand U1736 (N_1736,N_888,N_1457);
xnor U1737 (N_1737,N_991,N_948);
nand U1738 (N_1738,N_1299,N_1523);
or U1739 (N_1739,N_1548,N_937);
and U1740 (N_1740,N_1338,N_995);
and U1741 (N_1741,N_1102,N_1032);
nor U1742 (N_1742,N_1187,N_1425);
nand U1743 (N_1743,N_1088,N_1207);
or U1744 (N_1744,N_810,N_1370);
or U1745 (N_1745,N_1516,N_1226);
nand U1746 (N_1746,N_980,N_1095);
or U1747 (N_1747,N_1506,N_1567);
nor U1748 (N_1748,N_864,N_1251);
nor U1749 (N_1749,N_985,N_956);
or U1750 (N_1750,N_1293,N_1052);
xnor U1751 (N_1751,N_1397,N_1145);
nor U1752 (N_1752,N_942,N_1197);
or U1753 (N_1753,N_833,N_1093);
nand U1754 (N_1754,N_1327,N_1139);
nor U1755 (N_1755,N_881,N_1353);
and U1756 (N_1756,N_1486,N_1286);
or U1757 (N_1757,N_1540,N_1122);
nand U1758 (N_1758,N_1531,N_849);
nand U1759 (N_1759,N_1387,N_1080);
and U1760 (N_1760,N_1101,N_1178);
or U1761 (N_1761,N_822,N_999);
or U1762 (N_1762,N_1033,N_808);
or U1763 (N_1763,N_1435,N_1053);
or U1764 (N_1764,N_971,N_1365);
nand U1765 (N_1765,N_1511,N_1236);
xnor U1766 (N_1766,N_1396,N_1474);
or U1767 (N_1767,N_1542,N_866);
nor U1768 (N_1768,N_884,N_1333);
nand U1769 (N_1769,N_1464,N_1460);
nor U1770 (N_1770,N_1470,N_946);
and U1771 (N_1771,N_1478,N_1202);
xor U1772 (N_1772,N_1100,N_1144);
xnor U1773 (N_1773,N_893,N_1018);
or U1774 (N_1774,N_1193,N_1219);
or U1775 (N_1775,N_1334,N_1311);
xnor U1776 (N_1776,N_1228,N_1544);
and U1777 (N_1777,N_1120,N_1459);
or U1778 (N_1778,N_1546,N_1025);
nor U1779 (N_1779,N_1023,N_1281);
nor U1780 (N_1780,N_1063,N_1172);
or U1781 (N_1781,N_926,N_1537);
nor U1782 (N_1782,N_1142,N_894);
and U1783 (N_1783,N_862,N_1599);
xnor U1784 (N_1784,N_1248,N_823);
nor U1785 (N_1785,N_1157,N_1591);
or U1786 (N_1786,N_898,N_1525);
nand U1787 (N_1787,N_1357,N_905);
nor U1788 (N_1788,N_887,N_1287);
and U1789 (N_1789,N_1499,N_1051);
xnor U1790 (N_1790,N_907,N_1231);
xor U1791 (N_1791,N_863,N_1078);
or U1792 (N_1792,N_1555,N_1495);
nand U1793 (N_1793,N_824,N_1426);
nand U1794 (N_1794,N_1566,N_1453);
nand U1795 (N_1795,N_1587,N_1361);
xor U1796 (N_1796,N_1465,N_934);
xor U1797 (N_1797,N_819,N_1419);
and U1798 (N_1798,N_1020,N_1265);
and U1799 (N_1799,N_994,N_1494);
xnor U1800 (N_1800,N_1289,N_820);
and U1801 (N_1801,N_856,N_903);
nand U1802 (N_1802,N_826,N_1301);
and U1803 (N_1803,N_1105,N_967);
nand U1804 (N_1804,N_939,N_1222);
xor U1805 (N_1805,N_920,N_1324);
and U1806 (N_1806,N_1451,N_830);
xor U1807 (N_1807,N_1498,N_1507);
nor U1808 (N_1808,N_1282,N_1143);
or U1809 (N_1809,N_1146,N_1371);
nand U1810 (N_1810,N_1583,N_1149);
nor U1811 (N_1811,N_1337,N_1503);
nor U1812 (N_1812,N_1192,N_958);
or U1813 (N_1813,N_1593,N_1117);
nand U1814 (N_1814,N_875,N_1380);
nand U1815 (N_1815,N_1005,N_1580);
nor U1816 (N_1816,N_1450,N_1104);
nand U1817 (N_1817,N_1097,N_1476);
nand U1818 (N_1818,N_1167,N_1132);
nor U1819 (N_1819,N_1118,N_1473);
and U1820 (N_1820,N_1234,N_1477);
or U1821 (N_1821,N_865,N_1382);
xor U1822 (N_1822,N_1179,N_1595);
nand U1823 (N_1823,N_1565,N_1200);
nand U1824 (N_1824,N_1027,N_955);
nand U1825 (N_1825,N_1176,N_909);
or U1826 (N_1826,N_1436,N_1410);
and U1827 (N_1827,N_1003,N_1594);
xnor U1828 (N_1828,N_1004,N_953);
nand U1829 (N_1829,N_981,N_1529);
nor U1830 (N_1830,N_1429,N_951);
and U1831 (N_1831,N_1359,N_1280);
nand U1832 (N_1832,N_1440,N_869);
nand U1833 (N_1833,N_895,N_1292);
nor U1834 (N_1834,N_1527,N_1277);
or U1835 (N_1835,N_957,N_1514);
or U1836 (N_1836,N_1038,N_1418);
and U1837 (N_1837,N_1195,N_1469);
and U1838 (N_1838,N_968,N_1294);
or U1839 (N_1839,N_1209,N_1283);
nor U1840 (N_1840,N_821,N_885);
nor U1841 (N_1841,N_1274,N_852);
or U1842 (N_1842,N_1256,N_1047);
or U1843 (N_1843,N_1316,N_1597);
xor U1844 (N_1844,N_983,N_1322);
nor U1845 (N_1845,N_1437,N_1319);
nand U1846 (N_1846,N_1160,N_966);
or U1847 (N_1847,N_1141,N_1482);
xnor U1848 (N_1848,N_1072,N_1278);
nor U1849 (N_1849,N_1392,N_1570);
and U1850 (N_1850,N_1581,N_806);
xnor U1851 (N_1851,N_1199,N_1168);
and U1852 (N_1852,N_1584,N_1229);
and U1853 (N_1853,N_1343,N_1147);
or U1854 (N_1854,N_1306,N_1125);
nor U1855 (N_1855,N_1075,N_876);
or U1856 (N_1856,N_900,N_1250);
nor U1857 (N_1857,N_1386,N_993);
or U1858 (N_1858,N_1181,N_1439);
nor U1859 (N_1859,N_1191,N_805);
nor U1860 (N_1860,N_1415,N_1010);
nor U1861 (N_1861,N_890,N_854);
nand U1862 (N_1862,N_1173,N_1015);
nor U1863 (N_1863,N_1019,N_970);
or U1864 (N_1864,N_947,N_842);
xor U1865 (N_1865,N_1427,N_1262);
xor U1866 (N_1866,N_1524,N_899);
or U1867 (N_1867,N_1519,N_1407);
and U1868 (N_1868,N_1285,N_1158);
nand U1869 (N_1869,N_1315,N_1182);
nand U1870 (N_1870,N_945,N_1112);
and U1871 (N_1871,N_1001,N_801);
nand U1872 (N_1872,N_802,N_1151);
xnor U1873 (N_1873,N_1409,N_982);
nor U1874 (N_1874,N_1170,N_1071);
and U1875 (N_1875,N_1030,N_1252);
nor U1876 (N_1876,N_1491,N_1090);
nor U1877 (N_1877,N_1084,N_1354);
xnor U1878 (N_1878,N_1479,N_921);
and U1879 (N_1879,N_1216,N_1073);
nand U1880 (N_1880,N_1326,N_1552);
nand U1881 (N_1881,N_1341,N_1119);
and U1882 (N_1882,N_841,N_1206);
xor U1883 (N_1883,N_990,N_998);
nand U1884 (N_1884,N_1543,N_1308);
or U1885 (N_1885,N_973,N_844);
xor U1886 (N_1886,N_1064,N_1538);
nor U1887 (N_1887,N_1039,N_1561);
and U1888 (N_1888,N_837,N_828);
xnor U1889 (N_1889,N_1154,N_1017);
nor U1890 (N_1890,N_1330,N_1358);
and U1891 (N_1891,N_1098,N_1504);
xor U1892 (N_1892,N_901,N_927);
nand U1893 (N_1893,N_1109,N_1270);
xnor U1894 (N_1894,N_1124,N_1106);
and U1895 (N_1895,N_1008,N_1180);
nor U1896 (N_1896,N_1049,N_963);
nor U1897 (N_1897,N_857,N_1037);
xor U1898 (N_1898,N_1586,N_1086);
and U1899 (N_1899,N_1417,N_1456);
xnor U1900 (N_1900,N_1190,N_803);
or U1901 (N_1901,N_880,N_1518);
nor U1902 (N_1902,N_817,N_1342);
nand U1903 (N_1903,N_1205,N_902);
nor U1904 (N_1904,N_1458,N_1545);
and U1905 (N_1905,N_1318,N_1363);
xor U1906 (N_1906,N_1582,N_1055);
and U1907 (N_1907,N_1099,N_961);
or U1908 (N_1908,N_804,N_1452);
or U1909 (N_1909,N_1317,N_1136);
or U1910 (N_1910,N_1267,N_1385);
nor U1911 (N_1911,N_1362,N_858);
xnor U1912 (N_1912,N_1126,N_1534);
and U1913 (N_1913,N_1133,N_1340);
nand U1914 (N_1914,N_1484,N_1462);
nor U1915 (N_1915,N_906,N_1271);
nand U1916 (N_1916,N_878,N_1520);
or U1917 (N_1917,N_977,N_1313);
or U1918 (N_1918,N_1029,N_1096);
nand U1919 (N_1919,N_1376,N_835);
nor U1920 (N_1920,N_1320,N_1336);
or U1921 (N_1921,N_1233,N_1471);
nand U1922 (N_1922,N_1121,N_1201);
or U1923 (N_1923,N_1556,N_1505);
and U1924 (N_1924,N_1549,N_1203);
and U1925 (N_1925,N_1103,N_889);
nand U1926 (N_1926,N_1254,N_1066);
or U1927 (N_1927,N_832,N_944);
nor U1928 (N_1928,N_976,N_1085);
xnor U1929 (N_1929,N_1221,N_1335);
nand U1930 (N_1930,N_1291,N_1304);
nor U1931 (N_1931,N_1067,N_1116);
and U1932 (N_1932,N_1442,N_1212);
and U1933 (N_1933,N_930,N_1446);
and U1934 (N_1934,N_1303,N_1596);
nand U1935 (N_1935,N_1186,N_1013);
nor U1936 (N_1936,N_1428,N_825);
xnor U1937 (N_1937,N_851,N_1508);
nand U1938 (N_1938,N_1577,N_1152);
or U1939 (N_1939,N_1406,N_1454);
nand U1940 (N_1940,N_1501,N_1564);
nor U1941 (N_1941,N_1487,N_1269);
xnor U1942 (N_1942,N_892,N_987);
nand U1943 (N_1943,N_1480,N_911);
nor U1944 (N_1944,N_1528,N_1485);
nand U1945 (N_1945,N_1438,N_1443);
xor U1946 (N_1946,N_831,N_1092);
xor U1947 (N_1947,N_814,N_1150);
or U1948 (N_1948,N_1016,N_897);
nand U1949 (N_1949,N_1264,N_1389);
and U1950 (N_1950,N_1215,N_871);
or U1951 (N_1951,N_1422,N_1076);
nor U1952 (N_1952,N_1110,N_1041);
xnor U1953 (N_1953,N_1257,N_1177);
nor U1954 (N_1954,N_1312,N_1081);
xor U1955 (N_1955,N_1138,N_1349);
nand U1956 (N_1956,N_984,N_1002);
and U1957 (N_1957,N_1539,N_1401);
or U1958 (N_1958,N_1558,N_1368);
xor U1959 (N_1959,N_1355,N_940);
nand U1960 (N_1960,N_1420,N_1161);
or U1961 (N_1961,N_1403,N_1065);
xor U1962 (N_1962,N_1412,N_1483);
nor U1963 (N_1963,N_1046,N_1492);
nor U1964 (N_1964,N_1550,N_1174);
nand U1965 (N_1965,N_1134,N_877);
nand U1966 (N_1966,N_1213,N_1298);
nor U1967 (N_1967,N_1323,N_1175);
xor U1968 (N_1968,N_1210,N_1012);
or U1969 (N_1969,N_1079,N_813);
nor U1970 (N_1970,N_1245,N_1388);
and U1971 (N_1971,N_1332,N_800);
nand U1972 (N_1972,N_1488,N_954);
nand U1973 (N_1973,N_1014,N_1411);
nand U1974 (N_1974,N_1416,N_1344);
nor U1975 (N_1975,N_915,N_1585);
or U1976 (N_1976,N_1381,N_1364);
and U1977 (N_1977,N_913,N_1526);
xor U1978 (N_1978,N_1290,N_1077);
or U1979 (N_1979,N_1288,N_938);
or U1980 (N_1980,N_1532,N_1433);
xor U1981 (N_1981,N_1378,N_1224);
nand U1982 (N_1982,N_986,N_914);
nor U1983 (N_1983,N_1031,N_1372);
nand U1984 (N_1984,N_1329,N_896);
and U1985 (N_1985,N_1059,N_1241);
or U1986 (N_1986,N_1350,N_1563);
xnor U1987 (N_1987,N_904,N_1056);
nor U1988 (N_1988,N_1054,N_1034);
nor U1989 (N_1989,N_1214,N_1490);
or U1990 (N_1990,N_1576,N_1541);
or U1991 (N_1991,N_1249,N_1305);
and U1992 (N_1992,N_1156,N_923);
nor U1993 (N_1993,N_1069,N_1275);
nor U1994 (N_1994,N_1153,N_1379);
xor U1995 (N_1995,N_1184,N_861);
nand U1996 (N_1996,N_969,N_1475);
nor U1997 (N_1997,N_996,N_1441);
xor U1998 (N_1998,N_1114,N_952);
or U1999 (N_1999,N_1468,N_1227);
nor U2000 (N_2000,N_1463,N_1091);
or U2001 (N_2001,N_911,N_1009);
or U2002 (N_2002,N_923,N_1118);
or U2003 (N_2003,N_1302,N_1502);
and U2004 (N_2004,N_1165,N_1348);
nand U2005 (N_2005,N_1416,N_1489);
nor U2006 (N_2006,N_1032,N_1460);
xnor U2007 (N_2007,N_1107,N_1481);
nor U2008 (N_2008,N_1248,N_1464);
xnor U2009 (N_2009,N_863,N_862);
and U2010 (N_2010,N_1438,N_1054);
and U2011 (N_2011,N_960,N_966);
nand U2012 (N_2012,N_1022,N_1454);
and U2013 (N_2013,N_1054,N_1298);
nor U2014 (N_2014,N_929,N_1260);
nand U2015 (N_2015,N_1028,N_809);
and U2016 (N_2016,N_1516,N_1312);
or U2017 (N_2017,N_1066,N_1344);
nand U2018 (N_2018,N_1441,N_1145);
nand U2019 (N_2019,N_1235,N_1113);
or U2020 (N_2020,N_1155,N_1282);
or U2021 (N_2021,N_1510,N_1094);
and U2022 (N_2022,N_1051,N_1596);
and U2023 (N_2023,N_1562,N_1031);
and U2024 (N_2024,N_1200,N_1364);
xor U2025 (N_2025,N_1564,N_839);
xnor U2026 (N_2026,N_1367,N_1534);
and U2027 (N_2027,N_1230,N_1473);
or U2028 (N_2028,N_1411,N_957);
nor U2029 (N_2029,N_1431,N_947);
or U2030 (N_2030,N_1270,N_1597);
and U2031 (N_2031,N_1090,N_1213);
nand U2032 (N_2032,N_879,N_1000);
and U2033 (N_2033,N_1481,N_830);
and U2034 (N_2034,N_1473,N_998);
or U2035 (N_2035,N_1366,N_1421);
xnor U2036 (N_2036,N_1231,N_1074);
xnor U2037 (N_2037,N_1130,N_1221);
nor U2038 (N_2038,N_1094,N_1533);
nand U2039 (N_2039,N_1451,N_1108);
and U2040 (N_2040,N_1317,N_1222);
or U2041 (N_2041,N_1276,N_1526);
nand U2042 (N_2042,N_1412,N_1101);
xor U2043 (N_2043,N_1151,N_968);
nor U2044 (N_2044,N_805,N_1414);
nand U2045 (N_2045,N_1267,N_1478);
nor U2046 (N_2046,N_1594,N_1039);
xor U2047 (N_2047,N_821,N_1506);
nand U2048 (N_2048,N_1563,N_1141);
and U2049 (N_2049,N_1156,N_1149);
nand U2050 (N_2050,N_1038,N_1111);
nor U2051 (N_2051,N_1251,N_1372);
or U2052 (N_2052,N_1297,N_1392);
nor U2053 (N_2053,N_1455,N_1267);
xor U2054 (N_2054,N_1323,N_1312);
or U2055 (N_2055,N_859,N_916);
nor U2056 (N_2056,N_1356,N_835);
xnor U2057 (N_2057,N_1205,N_1246);
and U2058 (N_2058,N_1159,N_1016);
nor U2059 (N_2059,N_1348,N_961);
nor U2060 (N_2060,N_819,N_1024);
nand U2061 (N_2061,N_1055,N_1053);
and U2062 (N_2062,N_1132,N_1210);
and U2063 (N_2063,N_1175,N_1221);
and U2064 (N_2064,N_888,N_839);
nor U2065 (N_2065,N_1107,N_1463);
nand U2066 (N_2066,N_1523,N_895);
and U2067 (N_2067,N_1117,N_1350);
xor U2068 (N_2068,N_1535,N_1195);
and U2069 (N_2069,N_962,N_1417);
xnor U2070 (N_2070,N_1232,N_1547);
nand U2071 (N_2071,N_1051,N_1236);
or U2072 (N_2072,N_1521,N_1321);
and U2073 (N_2073,N_803,N_971);
or U2074 (N_2074,N_1146,N_1513);
and U2075 (N_2075,N_1453,N_1450);
and U2076 (N_2076,N_1200,N_1057);
nor U2077 (N_2077,N_860,N_1115);
and U2078 (N_2078,N_1549,N_1394);
nor U2079 (N_2079,N_1262,N_836);
xor U2080 (N_2080,N_801,N_1181);
nor U2081 (N_2081,N_1029,N_1112);
or U2082 (N_2082,N_828,N_1477);
nand U2083 (N_2083,N_1312,N_1536);
and U2084 (N_2084,N_1018,N_857);
nor U2085 (N_2085,N_1210,N_1586);
xnor U2086 (N_2086,N_1590,N_1018);
and U2087 (N_2087,N_868,N_1142);
xor U2088 (N_2088,N_1409,N_1200);
xor U2089 (N_2089,N_1575,N_1312);
and U2090 (N_2090,N_1316,N_1014);
nor U2091 (N_2091,N_1099,N_818);
or U2092 (N_2092,N_995,N_1498);
or U2093 (N_2093,N_941,N_1054);
xor U2094 (N_2094,N_879,N_1504);
nor U2095 (N_2095,N_1350,N_1145);
xor U2096 (N_2096,N_930,N_1393);
nand U2097 (N_2097,N_1292,N_1028);
nand U2098 (N_2098,N_991,N_817);
xnor U2099 (N_2099,N_1125,N_808);
and U2100 (N_2100,N_994,N_1161);
xor U2101 (N_2101,N_1184,N_1379);
and U2102 (N_2102,N_1296,N_1246);
nor U2103 (N_2103,N_1255,N_1316);
or U2104 (N_2104,N_894,N_952);
and U2105 (N_2105,N_1182,N_1268);
nor U2106 (N_2106,N_919,N_1019);
nor U2107 (N_2107,N_1484,N_1488);
xnor U2108 (N_2108,N_1514,N_1397);
and U2109 (N_2109,N_1503,N_1193);
nor U2110 (N_2110,N_1422,N_1343);
or U2111 (N_2111,N_964,N_1274);
or U2112 (N_2112,N_1091,N_1466);
or U2113 (N_2113,N_938,N_926);
nor U2114 (N_2114,N_1452,N_1085);
nor U2115 (N_2115,N_1014,N_907);
nor U2116 (N_2116,N_1120,N_917);
xnor U2117 (N_2117,N_1463,N_1114);
or U2118 (N_2118,N_1079,N_1579);
nand U2119 (N_2119,N_1380,N_1330);
nor U2120 (N_2120,N_1076,N_983);
nor U2121 (N_2121,N_1547,N_1470);
nand U2122 (N_2122,N_1555,N_943);
nand U2123 (N_2123,N_1220,N_1374);
or U2124 (N_2124,N_1461,N_1464);
or U2125 (N_2125,N_1043,N_953);
and U2126 (N_2126,N_1333,N_886);
xnor U2127 (N_2127,N_1443,N_1200);
xor U2128 (N_2128,N_834,N_1079);
nor U2129 (N_2129,N_1264,N_1408);
nand U2130 (N_2130,N_865,N_1121);
or U2131 (N_2131,N_1136,N_1120);
or U2132 (N_2132,N_1563,N_1086);
and U2133 (N_2133,N_957,N_1062);
xnor U2134 (N_2134,N_1111,N_1480);
or U2135 (N_2135,N_1295,N_997);
nand U2136 (N_2136,N_869,N_946);
nor U2137 (N_2137,N_1242,N_1471);
xor U2138 (N_2138,N_815,N_1382);
nor U2139 (N_2139,N_1404,N_816);
and U2140 (N_2140,N_1053,N_1388);
nor U2141 (N_2141,N_1207,N_843);
xnor U2142 (N_2142,N_1219,N_927);
and U2143 (N_2143,N_827,N_939);
xor U2144 (N_2144,N_1181,N_1542);
or U2145 (N_2145,N_1464,N_1028);
nand U2146 (N_2146,N_1483,N_1112);
and U2147 (N_2147,N_1301,N_1432);
nand U2148 (N_2148,N_900,N_1028);
xor U2149 (N_2149,N_1539,N_844);
or U2150 (N_2150,N_946,N_943);
or U2151 (N_2151,N_847,N_959);
xor U2152 (N_2152,N_1366,N_1005);
nor U2153 (N_2153,N_1417,N_838);
nand U2154 (N_2154,N_1509,N_1344);
nand U2155 (N_2155,N_1154,N_1005);
nand U2156 (N_2156,N_1165,N_1462);
xor U2157 (N_2157,N_957,N_1552);
nor U2158 (N_2158,N_1152,N_824);
xnor U2159 (N_2159,N_971,N_1039);
nand U2160 (N_2160,N_1436,N_1460);
or U2161 (N_2161,N_896,N_1352);
nor U2162 (N_2162,N_1069,N_1006);
xnor U2163 (N_2163,N_850,N_1561);
xnor U2164 (N_2164,N_1467,N_1376);
or U2165 (N_2165,N_1456,N_1062);
nor U2166 (N_2166,N_920,N_1598);
nand U2167 (N_2167,N_953,N_923);
or U2168 (N_2168,N_994,N_1068);
and U2169 (N_2169,N_886,N_1591);
xor U2170 (N_2170,N_1279,N_898);
nor U2171 (N_2171,N_925,N_1336);
or U2172 (N_2172,N_1282,N_1041);
and U2173 (N_2173,N_1530,N_846);
or U2174 (N_2174,N_847,N_819);
and U2175 (N_2175,N_1077,N_880);
xnor U2176 (N_2176,N_949,N_1306);
or U2177 (N_2177,N_1598,N_1161);
nand U2178 (N_2178,N_1206,N_1533);
or U2179 (N_2179,N_897,N_1266);
nand U2180 (N_2180,N_1094,N_1379);
nor U2181 (N_2181,N_1584,N_1466);
nor U2182 (N_2182,N_860,N_821);
and U2183 (N_2183,N_1111,N_971);
nand U2184 (N_2184,N_944,N_1055);
and U2185 (N_2185,N_1110,N_1222);
or U2186 (N_2186,N_1080,N_1082);
xor U2187 (N_2187,N_1223,N_1135);
nor U2188 (N_2188,N_1207,N_886);
nor U2189 (N_2189,N_984,N_924);
or U2190 (N_2190,N_1082,N_989);
nand U2191 (N_2191,N_941,N_847);
xor U2192 (N_2192,N_1358,N_895);
xnor U2193 (N_2193,N_1254,N_1455);
xnor U2194 (N_2194,N_1153,N_1297);
xor U2195 (N_2195,N_958,N_846);
or U2196 (N_2196,N_1465,N_905);
nor U2197 (N_2197,N_800,N_1294);
or U2198 (N_2198,N_1178,N_1424);
xor U2199 (N_2199,N_893,N_963);
nand U2200 (N_2200,N_1107,N_1591);
nor U2201 (N_2201,N_864,N_1057);
nor U2202 (N_2202,N_1431,N_1071);
nand U2203 (N_2203,N_855,N_955);
xnor U2204 (N_2204,N_1121,N_821);
or U2205 (N_2205,N_1595,N_1371);
and U2206 (N_2206,N_1310,N_963);
nor U2207 (N_2207,N_983,N_1332);
nand U2208 (N_2208,N_1289,N_1176);
or U2209 (N_2209,N_1025,N_834);
nand U2210 (N_2210,N_944,N_1396);
or U2211 (N_2211,N_966,N_1179);
xnor U2212 (N_2212,N_867,N_1182);
and U2213 (N_2213,N_800,N_1142);
nor U2214 (N_2214,N_1261,N_1214);
nand U2215 (N_2215,N_1536,N_1497);
nand U2216 (N_2216,N_1256,N_1104);
nor U2217 (N_2217,N_908,N_1143);
and U2218 (N_2218,N_1344,N_1378);
nor U2219 (N_2219,N_1288,N_954);
xor U2220 (N_2220,N_1067,N_1250);
and U2221 (N_2221,N_1375,N_1124);
nor U2222 (N_2222,N_983,N_1319);
nand U2223 (N_2223,N_916,N_971);
and U2224 (N_2224,N_1487,N_943);
xor U2225 (N_2225,N_1487,N_1072);
nand U2226 (N_2226,N_1461,N_1147);
nand U2227 (N_2227,N_1463,N_979);
or U2228 (N_2228,N_1114,N_879);
nand U2229 (N_2229,N_1347,N_1232);
nand U2230 (N_2230,N_1104,N_900);
nand U2231 (N_2231,N_828,N_1205);
nor U2232 (N_2232,N_888,N_1183);
and U2233 (N_2233,N_1270,N_844);
or U2234 (N_2234,N_1407,N_1462);
nand U2235 (N_2235,N_960,N_963);
or U2236 (N_2236,N_1500,N_1174);
or U2237 (N_2237,N_1434,N_1537);
nor U2238 (N_2238,N_1565,N_1078);
and U2239 (N_2239,N_1500,N_1103);
nor U2240 (N_2240,N_915,N_1002);
nand U2241 (N_2241,N_858,N_924);
xnor U2242 (N_2242,N_868,N_1207);
or U2243 (N_2243,N_824,N_1366);
and U2244 (N_2244,N_1337,N_986);
xor U2245 (N_2245,N_1172,N_922);
or U2246 (N_2246,N_1187,N_1510);
xor U2247 (N_2247,N_1040,N_1004);
xor U2248 (N_2248,N_1295,N_1049);
nor U2249 (N_2249,N_1459,N_1558);
or U2250 (N_2250,N_831,N_1400);
and U2251 (N_2251,N_1532,N_1430);
and U2252 (N_2252,N_884,N_1086);
nor U2253 (N_2253,N_968,N_884);
nor U2254 (N_2254,N_1392,N_1183);
nand U2255 (N_2255,N_818,N_837);
or U2256 (N_2256,N_1086,N_1077);
nor U2257 (N_2257,N_965,N_1446);
nor U2258 (N_2258,N_1533,N_1213);
xnor U2259 (N_2259,N_1588,N_1181);
or U2260 (N_2260,N_1380,N_1596);
or U2261 (N_2261,N_1318,N_889);
xor U2262 (N_2262,N_1409,N_905);
nand U2263 (N_2263,N_1057,N_1132);
nor U2264 (N_2264,N_830,N_1407);
nor U2265 (N_2265,N_1261,N_840);
xor U2266 (N_2266,N_874,N_1493);
nand U2267 (N_2267,N_1154,N_1157);
and U2268 (N_2268,N_913,N_1055);
nand U2269 (N_2269,N_1155,N_906);
nand U2270 (N_2270,N_935,N_1367);
and U2271 (N_2271,N_1217,N_1083);
nor U2272 (N_2272,N_1198,N_1090);
xor U2273 (N_2273,N_1146,N_915);
or U2274 (N_2274,N_1517,N_903);
or U2275 (N_2275,N_877,N_1110);
xnor U2276 (N_2276,N_800,N_1003);
nor U2277 (N_2277,N_909,N_1481);
nand U2278 (N_2278,N_925,N_1471);
nand U2279 (N_2279,N_1472,N_870);
nor U2280 (N_2280,N_1598,N_1262);
nand U2281 (N_2281,N_1426,N_1100);
or U2282 (N_2282,N_931,N_1163);
and U2283 (N_2283,N_1372,N_927);
nor U2284 (N_2284,N_1460,N_954);
nand U2285 (N_2285,N_803,N_1330);
xor U2286 (N_2286,N_1103,N_1347);
and U2287 (N_2287,N_1290,N_1229);
xor U2288 (N_2288,N_1461,N_1188);
xor U2289 (N_2289,N_1352,N_1126);
or U2290 (N_2290,N_963,N_1337);
nand U2291 (N_2291,N_1085,N_1236);
or U2292 (N_2292,N_1479,N_1583);
nand U2293 (N_2293,N_1441,N_1167);
or U2294 (N_2294,N_873,N_1408);
nor U2295 (N_2295,N_1023,N_1450);
nor U2296 (N_2296,N_1272,N_996);
nor U2297 (N_2297,N_1498,N_873);
xnor U2298 (N_2298,N_1548,N_1124);
or U2299 (N_2299,N_1161,N_1458);
and U2300 (N_2300,N_1133,N_809);
and U2301 (N_2301,N_809,N_1217);
xnor U2302 (N_2302,N_862,N_1315);
nand U2303 (N_2303,N_1121,N_1301);
xnor U2304 (N_2304,N_1515,N_1124);
xnor U2305 (N_2305,N_1212,N_1067);
and U2306 (N_2306,N_1200,N_1130);
nor U2307 (N_2307,N_842,N_1159);
nor U2308 (N_2308,N_1160,N_1591);
xnor U2309 (N_2309,N_1245,N_1394);
xor U2310 (N_2310,N_1468,N_1446);
xnor U2311 (N_2311,N_1102,N_884);
or U2312 (N_2312,N_1350,N_1126);
xor U2313 (N_2313,N_1391,N_1270);
or U2314 (N_2314,N_984,N_1073);
and U2315 (N_2315,N_1546,N_1136);
and U2316 (N_2316,N_833,N_1081);
and U2317 (N_2317,N_1227,N_1048);
and U2318 (N_2318,N_1514,N_1143);
and U2319 (N_2319,N_1137,N_1534);
and U2320 (N_2320,N_1234,N_1565);
and U2321 (N_2321,N_1120,N_1111);
nor U2322 (N_2322,N_811,N_1479);
xnor U2323 (N_2323,N_1207,N_1359);
nand U2324 (N_2324,N_1295,N_1461);
xor U2325 (N_2325,N_1520,N_1596);
xnor U2326 (N_2326,N_1541,N_1490);
nor U2327 (N_2327,N_970,N_1011);
nor U2328 (N_2328,N_1546,N_1014);
xor U2329 (N_2329,N_1486,N_1326);
nand U2330 (N_2330,N_1435,N_1110);
and U2331 (N_2331,N_1019,N_1468);
nor U2332 (N_2332,N_824,N_1449);
nor U2333 (N_2333,N_1194,N_1351);
and U2334 (N_2334,N_1383,N_897);
or U2335 (N_2335,N_1471,N_1195);
xnor U2336 (N_2336,N_841,N_1082);
nor U2337 (N_2337,N_1576,N_1444);
nor U2338 (N_2338,N_981,N_1266);
xnor U2339 (N_2339,N_1586,N_1271);
nor U2340 (N_2340,N_1216,N_1276);
or U2341 (N_2341,N_1316,N_1413);
nand U2342 (N_2342,N_1235,N_1463);
nand U2343 (N_2343,N_1127,N_1053);
and U2344 (N_2344,N_1285,N_1216);
xnor U2345 (N_2345,N_854,N_830);
nor U2346 (N_2346,N_1514,N_1462);
nand U2347 (N_2347,N_1130,N_1008);
nand U2348 (N_2348,N_1188,N_870);
nand U2349 (N_2349,N_842,N_1441);
and U2350 (N_2350,N_1388,N_1041);
and U2351 (N_2351,N_1583,N_1414);
and U2352 (N_2352,N_1443,N_958);
xnor U2353 (N_2353,N_1154,N_1475);
or U2354 (N_2354,N_1096,N_1559);
nor U2355 (N_2355,N_1184,N_1572);
nand U2356 (N_2356,N_1019,N_1398);
and U2357 (N_2357,N_1197,N_1304);
and U2358 (N_2358,N_972,N_904);
or U2359 (N_2359,N_1024,N_1069);
nand U2360 (N_2360,N_1028,N_843);
or U2361 (N_2361,N_1339,N_1237);
nand U2362 (N_2362,N_896,N_1101);
nand U2363 (N_2363,N_1232,N_1112);
nand U2364 (N_2364,N_838,N_853);
or U2365 (N_2365,N_1062,N_1545);
or U2366 (N_2366,N_1045,N_1182);
nor U2367 (N_2367,N_1108,N_1464);
or U2368 (N_2368,N_1189,N_1461);
nand U2369 (N_2369,N_840,N_1136);
xnor U2370 (N_2370,N_1017,N_916);
and U2371 (N_2371,N_924,N_1335);
nand U2372 (N_2372,N_1279,N_1195);
or U2373 (N_2373,N_876,N_1183);
xor U2374 (N_2374,N_834,N_1409);
nor U2375 (N_2375,N_809,N_1277);
nand U2376 (N_2376,N_867,N_842);
and U2377 (N_2377,N_1362,N_1337);
nand U2378 (N_2378,N_1049,N_1594);
and U2379 (N_2379,N_1067,N_1003);
and U2380 (N_2380,N_852,N_1216);
xnor U2381 (N_2381,N_846,N_1587);
xnor U2382 (N_2382,N_1267,N_1502);
or U2383 (N_2383,N_1252,N_911);
and U2384 (N_2384,N_1242,N_871);
and U2385 (N_2385,N_826,N_1583);
xor U2386 (N_2386,N_1474,N_1557);
xor U2387 (N_2387,N_948,N_1189);
or U2388 (N_2388,N_1010,N_1508);
nor U2389 (N_2389,N_966,N_1185);
or U2390 (N_2390,N_1288,N_1542);
nor U2391 (N_2391,N_1111,N_833);
and U2392 (N_2392,N_1278,N_1187);
xor U2393 (N_2393,N_1320,N_1139);
xnor U2394 (N_2394,N_901,N_1158);
xnor U2395 (N_2395,N_1236,N_1577);
and U2396 (N_2396,N_1093,N_1186);
xor U2397 (N_2397,N_1161,N_1163);
nand U2398 (N_2398,N_813,N_1563);
and U2399 (N_2399,N_1216,N_1584);
nor U2400 (N_2400,N_1772,N_2259);
nor U2401 (N_2401,N_1742,N_1883);
xor U2402 (N_2402,N_1603,N_1931);
nand U2403 (N_2403,N_2313,N_1741);
xor U2404 (N_2404,N_1915,N_1826);
nor U2405 (N_2405,N_2316,N_2202);
xnor U2406 (N_2406,N_1950,N_1948);
nor U2407 (N_2407,N_1975,N_1893);
nor U2408 (N_2408,N_2383,N_2189);
or U2409 (N_2409,N_2036,N_1843);
xnor U2410 (N_2410,N_2214,N_2197);
or U2411 (N_2411,N_1935,N_2002);
and U2412 (N_2412,N_1808,N_1906);
xnor U2413 (N_2413,N_1832,N_1728);
and U2414 (N_2414,N_2394,N_2335);
nor U2415 (N_2415,N_1994,N_2295);
and U2416 (N_2416,N_2306,N_1890);
xnor U2417 (N_2417,N_2219,N_1690);
and U2418 (N_2418,N_1745,N_2270);
and U2419 (N_2419,N_2044,N_2091);
nand U2420 (N_2420,N_2369,N_2321);
nand U2421 (N_2421,N_1819,N_2042);
and U2422 (N_2422,N_1983,N_1848);
nor U2423 (N_2423,N_2209,N_2255);
nor U2424 (N_2424,N_1946,N_2134);
and U2425 (N_2425,N_1771,N_1961);
nor U2426 (N_2426,N_2376,N_2346);
or U2427 (N_2427,N_1767,N_2319);
nor U2428 (N_2428,N_2297,N_1886);
nor U2429 (N_2429,N_2308,N_1973);
and U2430 (N_2430,N_1662,N_1933);
or U2431 (N_2431,N_2130,N_2194);
xor U2432 (N_2432,N_2039,N_1696);
or U2433 (N_2433,N_2092,N_2048);
xor U2434 (N_2434,N_2291,N_2017);
nor U2435 (N_2435,N_2276,N_1941);
and U2436 (N_2436,N_2244,N_1919);
xor U2437 (N_2437,N_2200,N_2104);
nand U2438 (N_2438,N_1943,N_2196);
or U2439 (N_2439,N_1630,N_1666);
or U2440 (N_2440,N_2298,N_1799);
xor U2441 (N_2441,N_2212,N_2050);
nand U2442 (N_2442,N_1959,N_1650);
xnor U2443 (N_2443,N_1790,N_2234);
xor U2444 (N_2444,N_1709,N_1770);
xor U2445 (N_2445,N_1902,N_2345);
nand U2446 (N_2446,N_2207,N_1929);
xor U2447 (N_2447,N_2094,N_1667);
nand U2448 (N_2448,N_1702,N_1956);
or U2449 (N_2449,N_1844,N_1677);
nor U2450 (N_2450,N_2162,N_2361);
nand U2451 (N_2451,N_1971,N_1699);
nor U2452 (N_2452,N_1715,N_1922);
nor U2453 (N_2453,N_1999,N_2339);
or U2454 (N_2454,N_2303,N_1672);
nand U2455 (N_2455,N_2309,N_2382);
nand U2456 (N_2456,N_1768,N_2347);
and U2457 (N_2457,N_2210,N_1888);
and U2458 (N_2458,N_1618,N_2026);
nand U2459 (N_2459,N_2389,N_2146);
nor U2460 (N_2460,N_2367,N_1987);
or U2461 (N_2461,N_2300,N_1782);
nand U2462 (N_2462,N_1825,N_2368);
nor U2463 (N_2463,N_2153,N_1688);
nor U2464 (N_2464,N_1676,N_2012);
xnor U2465 (N_2465,N_2000,N_2114);
nor U2466 (N_2466,N_2228,N_2386);
and U2467 (N_2467,N_1820,N_1720);
nand U2468 (N_2468,N_1727,N_1789);
nor U2469 (N_2469,N_2180,N_2078);
and U2470 (N_2470,N_1798,N_2187);
or U2471 (N_2471,N_1879,N_2107);
or U2472 (N_2472,N_1854,N_1644);
xnor U2473 (N_2473,N_2222,N_2317);
nand U2474 (N_2474,N_1701,N_2193);
nand U2475 (N_2475,N_1927,N_1997);
nor U2476 (N_2476,N_1884,N_2041);
nor U2477 (N_2477,N_2358,N_1641);
and U2478 (N_2478,N_2058,N_2179);
or U2479 (N_2479,N_1864,N_2384);
nand U2480 (N_2480,N_2084,N_2256);
nand U2481 (N_2481,N_1716,N_1680);
or U2482 (N_2482,N_1862,N_2360);
nand U2483 (N_2483,N_1998,N_1976);
or U2484 (N_2484,N_2066,N_1610);
and U2485 (N_2485,N_1646,N_2342);
nor U2486 (N_2486,N_1964,N_2357);
nor U2487 (N_2487,N_2003,N_1865);
nor U2488 (N_2488,N_1831,N_2023);
nand U2489 (N_2489,N_2217,N_1754);
and U2490 (N_2490,N_1810,N_2030);
and U2491 (N_2491,N_1907,N_1605);
xor U2492 (N_2492,N_2322,N_1981);
nand U2493 (N_2493,N_2129,N_2371);
nor U2494 (N_2494,N_2395,N_1990);
nor U2495 (N_2495,N_1985,N_1800);
xor U2496 (N_2496,N_2333,N_2304);
and U2497 (N_2497,N_2059,N_1734);
xnor U2498 (N_2498,N_1868,N_1803);
nand U2499 (N_2499,N_2109,N_2230);
and U2500 (N_2500,N_1962,N_1801);
and U2501 (N_2501,N_1954,N_2277);
and U2502 (N_2502,N_2315,N_1615);
and U2503 (N_2503,N_1995,N_1796);
xor U2504 (N_2504,N_2213,N_1815);
and U2505 (N_2505,N_1735,N_1881);
nand U2506 (N_2506,N_1938,N_2205);
or U2507 (N_2507,N_2174,N_2353);
nand U2508 (N_2508,N_1600,N_1988);
and U2509 (N_2509,N_1934,N_1762);
nand U2510 (N_2510,N_2172,N_2390);
xnor U2511 (N_2511,N_2211,N_1637);
and U2512 (N_2512,N_1899,N_1953);
nor U2513 (N_2513,N_2126,N_2201);
or U2514 (N_2514,N_1857,N_1664);
nand U2515 (N_2515,N_2103,N_2359);
nor U2516 (N_2516,N_1957,N_1977);
xor U2517 (N_2517,N_1678,N_1923);
or U2518 (N_2518,N_1697,N_1894);
and U2519 (N_2519,N_2152,N_1895);
xor U2520 (N_2520,N_2005,N_2019);
or U2521 (N_2521,N_1773,N_2031);
nand U2522 (N_2522,N_2248,N_2151);
xor U2523 (N_2523,N_2159,N_1694);
nor U2524 (N_2524,N_2198,N_1970);
xnor U2525 (N_2525,N_2073,N_2204);
or U2526 (N_2526,N_1784,N_2133);
nand U2527 (N_2527,N_2334,N_1651);
nor U2528 (N_2528,N_2249,N_2354);
and U2529 (N_2529,N_2254,N_2307);
and U2530 (N_2530,N_1717,N_2370);
nor U2531 (N_2531,N_1858,N_2061);
xnor U2532 (N_2532,N_2349,N_1723);
nor U2533 (N_2533,N_2293,N_2171);
nand U2534 (N_2534,N_1759,N_2034);
xnor U2535 (N_2535,N_1682,N_2267);
or U2536 (N_2536,N_1613,N_2232);
nor U2537 (N_2537,N_1875,N_1670);
nor U2538 (N_2538,N_2138,N_2344);
nand U2539 (N_2539,N_1758,N_1869);
xnor U2540 (N_2540,N_1642,N_1856);
or U2541 (N_2541,N_2013,N_2010);
xor U2542 (N_2542,N_2362,N_1969);
nand U2543 (N_2543,N_2243,N_1960);
nor U2544 (N_2544,N_1905,N_1732);
and U2545 (N_2545,N_1626,N_2074);
nor U2546 (N_2546,N_2252,N_1928);
nand U2547 (N_2547,N_2113,N_1910);
xnor U2548 (N_2548,N_2247,N_2085);
and U2549 (N_2549,N_1827,N_1674);
xnor U2550 (N_2550,N_2258,N_1925);
xnor U2551 (N_2551,N_2242,N_1748);
or U2552 (N_2552,N_2055,N_2191);
nand U2553 (N_2553,N_1795,N_2182);
xor U2554 (N_2554,N_1719,N_2124);
xor U2555 (N_2555,N_2278,N_1836);
xor U2556 (N_2556,N_1623,N_2327);
or U2557 (N_2557,N_1829,N_1628);
and U2558 (N_2558,N_2027,N_2233);
or U2559 (N_2559,N_2337,N_2238);
nand U2560 (N_2560,N_1947,N_2208);
xnor U2561 (N_2561,N_1660,N_2272);
and U2562 (N_2562,N_2150,N_2142);
nand U2563 (N_2563,N_1965,N_1781);
and U2564 (N_2564,N_1698,N_2336);
nand U2565 (N_2565,N_2086,N_1828);
xnor U2566 (N_2566,N_1643,N_1834);
nand U2567 (N_2567,N_1901,N_2090);
nand U2568 (N_2568,N_1774,N_2093);
nor U2569 (N_2569,N_1713,N_1802);
or U2570 (N_2570,N_1867,N_1870);
xor U2571 (N_2571,N_1718,N_2136);
nand U2572 (N_2572,N_1909,N_1652);
nand U2573 (N_2573,N_2241,N_1880);
xnor U2574 (N_2574,N_1982,N_1942);
and U2575 (N_2575,N_2177,N_2266);
or U2576 (N_2576,N_2377,N_2070);
xnor U2577 (N_2577,N_1992,N_2348);
or U2578 (N_2578,N_1740,N_1824);
or U2579 (N_2579,N_1612,N_1840);
xor U2580 (N_2580,N_2016,N_1835);
nand U2581 (N_2581,N_1914,N_2274);
nor U2582 (N_2582,N_1921,N_1917);
xor U2583 (N_2583,N_1611,N_1669);
and U2584 (N_2584,N_1783,N_1945);
and U2585 (N_2585,N_1695,N_1689);
xor U2586 (N_2586,N_1760,N_2236);
nor U2587 (N_2587,N_1638,N_1616);
or U2588 (N_2588,N_1786,N_1703);
xor U2589 (N_2589,N_1793,N_2271);
xor U2590 (N_2590,N_2275,N_1679);
and U2591 (N_2591,N_2154,N_1873);
and U2592 (N_2592,N_1704,N_2137);
or U2593 (N_2593,N_1937,N_1620);
xnor U2594 (N_2594,N_2119,N_1751);
or U2595 (N_2595,N_2149,N_2009);
and U2596 (N_2596,N_1739,N_1749);
or U2597 (N_2597,N_1776,N_2283);
or U2598 (N_2598,N_2169,N_2095);
xnor U2599 (N_2599,N_1996,N_2332);
nor U2600 (N_2600,N_1912,N_2140);
xnor U2601 (N_2601,N_1693,N_2082);
xor U2602 (N_2602,N_2024,N_2340);
nor U2603 (N_2603,N_1968,N_2284);
and U2604 (N_2604,N_1855,N_1871);
nand U2605 (N_2605,N_2101,N_1622);
nand U2606 (N_2606,N_1711,N_1645);
nand U2607 (N_2607,N_1958,N_2393);
nor U2608 (N_2608,N_2015,N_1794);
nand U2609 (N_2609,N_2374,N_1707);
xnor U2610 (N_2610,N_1775,N_1761);
and U2611 (N_2611,N_1809,N_2218);
and U2612 (N_2612,N_2328,N_1980);
xor U2613 (N_2613,N_2183,N_1648);
or U2614 (N_2614,N_2311,N_2077);
or U2615 (N_2615,N_1852,N_2163);
xor U2616 (N_2616,N_1683,N_1898);
nand U2617 (N_2617,N_2399,N_2157);
nor U2618 (N_2618,N_2100,N_2269);
nor U2619 (N_2619,N_2108,N_2088);
or U2620 (N_2620,N_2116,N_2299);
nand U2621 (N_2621,N_2166,N_2178);
nand U2622 (N_2622,N_2117,N_1866);
or U2623 (N_2623,N_2156,N_2155);
nor U2624 (N_2624,N_1668,N_2083);
nor U2625 (N_2625,N_1619,N_1691);
or U2626 (N_2626,N_1814,N_2381);
nor U2627 (N_2627,N_2111,N_2106);
xor U2628 (N_2628,N_2305,N_2047);
or U2629 (N_2629,N_2323,N_2320);
and U2630 (N_2630,N_2290,N_1700);
nand U2631 (N_2631,N_2161,N_1877);
nand U2632 (N_2632,N_2007,N_2318);
nand U2633 (N_2633,N_1708,N_2216);
nand U2634 (N_2634,N_1722,N_2080);
nor U2635 (N_2635,N_1845,N_1896);
xnor U2636 (N_2636,N_1918,N_2186);
nor U2637 (N_2637,N_2115,N_2294);
xnor U2638 (N_2638,N_2184,N_1932);
nor U2639 (N_2639,N_2246,N_2250);
or U2640 (N_2640,N_2122,N_2282);
xnor U2641 (N_2641,N_2287,N_2006);
or U2642 (N_2642,N_1724,N_1617);
or U2643 (N_2643,N_2279,N_2037);
or U2644 (N_2644,N_2018,N_2378);
and U2645 (N_2645,N_1710,N_2221);
xnor U2646 (N_2646,N_1705,N_2056);
nor U2647 (N_2647,N_1816,N_2051);
and U2648 (N_2648,N_1823,N_1939);
xnor U2649 (N_2649,N_1817,N_2069);
nand U2650 (N_2650,N_2063,N_2028);
or U2651 (N_2651,N_2167,N_2067);
and U2652 (N_2652,N_2262,N_1908);
and U2653 (N_2653,N_2231,N_2029);
or U2654 (N_2654,N_1634,N_2364);
or U2655 (N_2655,N_1807,N_2020);
and U2656 (N_2656,N_1882,N_2001);
nand U2657 (N_2657,N_1755,N_2068);
xor U2658 (N_2658,N_1853,N_1654);
nor U2659 (N_2659,N_2160,N_2014);
nor U2660 (N_2660,N_1846,N_2227);
nand U2661 (N_2661,N_1833,N_1659);
nor U2662 (N_2662,N_1665,N_2281);
or U2663 (N_2663,N_1850,N_2173);
and U2664 (N_2664,N_1874,N_1904);
xor U2665 (N_2665,N_1792,N_2225);
nand U2666 (N_2666,N_2072,N_1625);
nor U2667 (N_2667,N_2071,N_2203);
nand U2668 (N_2668,N_1635,N_1752);
or U2669 (N_2669,N_2008,N_2065);
and U2670 (N_2670,N_1614,N_2199);
nor U2671 (N_2671,N_2121,N_1897);
or U2672 (N_2672,N_2288,N_1889);
xor U2673 (N_2673,N_1636,N_1911);
xor U2674 (N_2674,N_1821,N_2025);
or U2675 (N_2675,N_2087,N_1811);
or U2676 (N_2676,N_1764,N_2057);
nand U2677 (N_2677,N_2123,N_1629);
nand U2678 (N_2678,N_1769,N_2188);
xnor U2679 (N_2679,N_2351,N_1812);
nand U2680 (N_2680,N_1859,N_1838);
nor U2681 (N_2681,N_2079,N_1972);
nand U2682 (N_2682,N_2379,N_2396);
and U2683 (N_2683,N_2145,N_2391);
nand U2684 (N_2684,N_1924,N_1730);
and U2685 (N_2685,N_1621,N_2135);
or U2686 (N_2686,N_1765,N_1841);
or U2687 (N_2687,N_2118,N_1737);
or U2688 (N_2688,N_1661,N_1930);
or U2689 (N_2689,N_1967,N_2285);
nand U2690 (N_2690,N_2261,N_1609);
xnor U2691 (N_2691,N_2128,N_2289);
nor U2692 (N_2692,N_2054,N_1989);
xor U2693 (N_2693,N_2190,N_1849);
nand U2694 (N_2694,N_1860,N_1861);
and U2695 (N_2695,N_2168,N_1604);
nand U2696 (N_2696,N_2141,N_1791);
nand U2697 (N_2697,N_1706,N_2240);
xor U2698 (N_2698,N_2338,N_1788);
nand U2699 (N_2699,N_2112,N_2224);
xor U2700 (N_2700,N_2011,N_1876);
and U2701 (N_2701,N_2397,N_1986);
nand U2702 (N_2702,N_1647,N_1916);
nand U2703 (N_2703,N_2110,N_1892);
xnor U2704 (N_2704,N_1822,N_1726);
or U2705 (N_2705,N_2314,N_1671);
nand U2706 (N_2706,N_2223,N_2060);
nor U2707 (N_2707,N_1632,N_1721);
and U2708 (N_2708,N_1631,N_2387);
xor U2709 (N_2709,N_1731,N_2372);
nor U2710 (N_2710,N_1872,N_2245);
xor U2711 (N_2711,N_1778,N_2170);
xor U2712 (N_2712,N_1974,N_1813);
xnor U2713 (N_2713,N_2049,N_1804);
nor U2714 (N_2714,N_2273,N_1797);
or U2715 (N_2715,N_2099,N_1766);
xor U2716 (N_2716,N_1900,N_1863);
nand U2717 (N_2717,N_2096,N_2046);
nor U2718 (N_2718,N_2365,N_1725);
nor U2719 (N_2719,N_2076,N_1714);
nor U2720 (N_2720,N_2280,N_2265);
or U2721 (N_2721,N_2075,N_1805);
xor U2722 (N_2722,N_1851,N_1952);
and U2723 (N_2723,N_1963,N_2021);
and U2724 (N_2724,N_2398,N_2098);
xnor U2725 (N_2725,N_1830,N_2175);
nand U2726 (N_2726,N_1951,N_1847);
and U2727 (N_2727,N_1649,N_2352);
and U2728 (N_2728,N_2032,N_2229);
nor U2729 (N_2729,N_1746,N_1878);
xor U2730 (N_2730,N_2324,N_2220);
and U2731 (N_2731,N_1743,N_1944);
or U2732 (N_2732,N_2350,N_2045);
and U2733 (N_2733,N_2143,N_2165);
nand U2734 (N_2734,N_2325,N_1744);
nor U2735 (N_2735,N_2144,N_2131);
and U2736 (N_2736,N_1949,N_2062);
and U2737 (N_2737,N_2164,N_1920);
xor U2738 (N_2738,N_2380,N_2296);
xor U2739 (N_2739,N_2251,N_1979);
and U2740 (N_2740,N_2355,N_2373);
nand U2741 (N_2741,N_1913,N_1777);
or U2742 (N_2742,N_2312,N_1780);
nand U2743 (N_2743,N_2329,N_1993);
nor U2744 (N_2744,N_1787,N_2192);
nor U2745 (N_2745,N_2081,N_2392);
and U2746 (N_2746,N_1763,N_2038);
or U2747 (N_2747,N_1955,N_1608);
nand U2748 (N_2748,N_2363,N_1738);
and U2749 (N_2749,N_1687,N_2301);
nor U2750 (N_2750,N_1655,N_1984);
xnor U2751 (N_2751,N_1926,N_2052);
or U2752 (N_2752,N_1940,N_2237);
or U2753 (N_2753,N_1684,N_2263);
nand U2754 (N_2754,N_2286,N_1842);
nand U2755 (N_2755,N_1606,N_2292);
nor U2756 (N_2756,N_2195,N_1885);
xnor U2757 (N_2757,N_1818,N_1675);
nor U2758 (N_2758,N_1839,N_2330);
or U2759 (N_2759,N_2302,N_1624);
or U2760 (N_2760,N_2127,N_2257);
and U2761 (N_2761,N_1903,N_2385);
nand U2762 (N_2762,N_2226,N_1656);
nor U2763 (N_2763,N_1653,N_1750);
nor U2764 (N_2764,N_1627,N_1779);
nor U2765 (N_2765,N_1729,N_1673);
and U2766 (N_2766,N_2033,N_2053);
nand U2767 (N_2767,N_2105,N_2215);
or U2768 (N_2768,N_2253,N_1991);
nand U2769 (N_2769,N_2132,N_2102);
or U2770 (N_2770,N_1658,N_2260);
nor U2771 (N_2771,N_2158,N_2264);
and U2772 (N_2772,N_1978,N_2040);
and U2773 (N_2773,N_1966,N_2064);
and U2774 (N_2774,N_2120,N_2268);
and U2775 (N_2775,N_2148,N_1686);
or U2776 (N_2776,N_2147,N_2185);
and U2777 (N_2777,N_2356,N_1891);
and U2778 (N_2778,N_2043,N_2239);
and U2779 (N_2779,N_2022,N_2375);
or U2780 (N_2780,N_2326,N_2366);
nor U2781 (N_2781,N_1756,N_2125);
nor U2782 (N_2782,N_1837,N_2004);
nor U2783 (N_2783,N_1936,N_1633);
and U2784 (N_2784,N_1733,N_1601);
nand U2785 (N_2785,N_1607,N_2235);
and U2786 (N_2786,N_2206,N_1712);
or U2787 (N_2787,N_2341,N_1753);
nor U2788 (N_2788,N_1736,N_2097);
or U2789 (N_2789,N_1887,N_1663);
and U2790 (N_2790,N_2331,N_2089);
nand U2791 (N_2791,N_1602,N_1757);
or U2792 (N_2792,N_1639,N_2035);
nand U2793 (N_2793,N_1681,N_1640);
and U2794 (N_2794,N_1747,N_2181);
or U2795 (N_2795,N_2139,N_2310);
and U2796 (N_2796,N_2388,N_1685);
xnor U2797 (N_2797,N_1806,N_1692);
and U2798 (N_2798,N_1785,N_2343);
nand U2799 (N_2799,N_2176,N_1657);
nor U2800 (N_2800,N_2330,N_1677);
or U2801 (N_2801,N_1999,N_1723);
or U2802 (N_2802,N_2227,N_2373);
nor U2803 (N_2803,N_1948,N_2144);
and U2804 (N_2804,N_2026,N_1831);
or U2805 (N_2805,N_2258,N_1964);
nor U2806 (N_2806,N_2138,N_2190);
and U2807 (N_2807,N_2111,N_2262);
nor U2808 (N_2808,N_2329,N_1750);
xor U2809 (N_2809,N_1965,N_2331);
nor U2810 (N_2810,N_1997,N_2280);
or U2811 (N_2811,N_2139,N_2148);
xnor U2812 (N_2812,N_2050,N_1829);
nand U2813 (N_2813,N_1977,N_2233);
xnor U2814 (N_2814,N_2141,N_1986);
xnor U2815 (N_2815,N_2355,N_1908);
nor U2816 (N_2816,N_2254,N_2202);
xor U2817 (N_2817,N_2241,N_2316);
nand U2818 (N_2818,N_2380,N_2075);
xor U2819 (N_2819,N_1995,N_1820);
nand U2820 (N_2820,N_1606,N_1695);
and U2821 (N_2821,N_1777,N_1696);
or U2822 (N_2822,N_1953,N_1624);
nand U2823 (N_2823,N_2070,N_2313);
xor U2824 (N_2824,N_1824,N_2391);
xnor U2825 (N_2825,N_2200,N_2387);
nand U2826 (N_2826,N_1756,N_2175);
nor U2827 (N_2827,N_1964,N_1693);
nor U2828 (N_2828,N_1810,N_1856);
or U2829 (N_2829,N_1766,N_2046);
or U2830 (N_2830,N_2080,N_1694);
xnor U2831 (N_2831,N_1766,N_2272);
and U2832 (N_2832,N_1924,N_2277);
nand U2833 (N_2833,N_2205,N_2370);
nand U2834 (N_2834,N_2053,N_2238);
nor U2835 (N_2835,N_1988,N_2262);
or U2836 (N_2836,N_2312,N_1637);
or U2837 (N_2837,N_2332,N_1619);
nor U2838 (N_2838,N_2370,N_1650);
and U2839 (N_2839,N_2111,N_1889);
nand U2840 (N_2840,N_2229,N_1873);
xnor U2841 (N_2841,N_2252,N_1902);
nor U2842 (N_2842,N_1881,N_2132);
or U2843 (N_2843,N_2289,N_2101);
xor U2844 (N_2844,N_2161,N_2227);
xor U2845 (N_2845,N_2084,N_2181);
nand U2846 (N_2846,N_1624,N_2379);
nor U2847 (N_2847,N_2079,N_2025);
nor U2848 (N_2848,N_1968,N_2053);
and U2849 (N_2849,N_1978,N_1732);
nor U2850 (N_2850,N_2305,N_2149);
or U2851 (N_2851,N_2177,N_1637);
xnor U2852 (N_2852,N_1954,N_2032);
xor U2853 (N_2853,N_2289,N_2312);
xnor U2854 (N_2854,N_2246,N_2082);
xor U2855 (N_2855,N_1648,N_2112);
or U2856 (N_2856,N_1854,N_2289);
and U2857 (N_2857,N_1619,N_1865);
and U2858 (N_2858,N_1891,N_2143);
or U2859 (N_2859,N_1651,N_2127);
nand U2860 (N_2860,N_1913,N_2068);
xnor U2861 (N_2861,N_1886,N_2255);
nor U2862 (N_2862,N_2091,N_1641);
xor U2863 (N_2863,N_1809,N_1714);
nor U2864 (N_2864,N_1873,N_1670);
or U2865 (N_2865,N_2363,N_1898);
xnor U2866 (N_2866,N_2213,N_1694);
xor U2867 (N_2867,N_2060,N_2393);
nor U2868 (N_2868,N_2174,N_1854);
nand U2869 (N_2869,N_2274,N_1854);
and U2870 (N_2870,N_2316,N_1911);
xor U2871 (N_2871,N_1739,N_2014);
or U2872 (N_2872,N_1911,N_1661);
nand U2873 (N_2873,N_1890,N_2173);
xor U2874 (N_2874,N_1637,N_1649);
nor U2875 (N_2875,N_1945,N_1796);
nor U2876 (N_2876,N_2099,N_1647);
xor U2877 (N_2877,N_1948,N_2352);
xnor U2878 (N_2878,N_1785,N_1832);
xnor U2879 (N_2879,N_2121,N_1604);
and U2880 (N_2880,N_1821,N_1932);
nor U2881 (N_2881,N_1874,N_2258);
nand U2882 (N_2882,N_1821,N_1992);
xnor U2883 (N_2883,N_1935,N_1616);
or U2884 (N_2884,N_1862,N_2122);
or U2885 (N_2885,N_2345,N_2296);
xnor U2886 (N_2886,N_1733,N_2152);
nor U2887 (N_2887,N_1832,N_1622);
nand U2888 (N_2888,N_2244,N_2384);
and U2889 (N_2889,N_1944,N_2334);
xnor U2890 (N_2890,N_2307,N_2120);
xnor U2891 (N_2891,N_1898,N_2159);
nor U2892 (N_2892,N_1763,N_2181);
nor U2893 (N_2893,N_1688,N_1997);
or U2894 (N_2894,N_2301,N_2049);
nand U2895 (N_2895,N_1696,N_1946);
xor U2896 (N_2896,N_2007,N_2319);
or U2897 (N_2897,N_2267,N_2262);
nand U2898 (N_2898,N_1945,N_2194);
xnor U2899 (N_2899,N_1878,N_1795);
nor U2900 (N_2900,N_1866,N_2291);
or U2901 (N_2901,N_1797,N_2018);
xor U2902 (N_2902,N_2157,N_1655);
or U2903 (N_2903,N_2222,N_1710);
nor U2904 (N_2904,N_1800,N_2200);
or U2905 (N_2905,N_2091,N_2037);
or U2906 (N_2906,N_2099,N_1952);
and U2907 (N_2907,N_1610,N_2364);
nor U2908 (N_2908,N_2282,N_1789);
and U2909 (N_2909,N_2052,N_2327);
nand U2910 (N_2910,N_1806,N_2295);
nand U2911 (N_2911,N_1904,N_1725);
nand U2912 (N_2912,N_2077,N_2060);
or U2913 (N_2913,N_1894,N_1732);
and U2914 (N_2914,N_2236,N_2200);
or U2915 (N_2915,N_1772,N_2187);
nor U2916 (N_2916,N_1995,N_2134);
nand U2917 (N_2917,N_2176,N_1941);
nand U2918 (N_2918,N_2311,N_2157);
or U2919 (N_2919,N_2268,N_2132);
nor U2920 (N_2920,N_1697,N_2343);
xnor U2921 (N_2921,N_1845,N_2375);
nor U2922 (N_2922,N_2117,N_2294);
nor U2923 (N_2923,N_1813,N_2218);
and U2924 (N_2924,N_1697,N_1942);
or U2925 (N_2925,N_2138,N_2374);
xnor U2926 (N_2926,N_2087,N_2191);
and U2927 (N_2927,N_2218,N_1656);
nor U2928 (N_2928,N_2299,N_1973);
or U2929 (N_2929,N_1887,N_2181);
xor U2930 (N_2930,N_1944,N_1976);
nand U2931 (N_2931,N_1951,N_1682);
and U2932 (N_2932,N_2376,N_1605);
nand U2933 (N_2933,N_1734,N_1867);
nand U2934 (N_2934,N_2082,N_1845);
and U2935 (N_2935,N_1921,N_2087);
and U2936 (N_2936,N_2203,N_1879);
nand U2937 (N_2937,N_1821,N_1635);
nor U2938 (N_2938,N_2135,N_1993);
nor U2939 (N_2939,N_1761,N_1923);
and U2940 (N_2940,N_2370,N_1910);
or U2941 (N_2941,N_1883,N_1899);
and U2942 (N_2942,N_1651,N_2009);
or U2943 (N_2943,N_1754,N_1731);
nor U2944 (N_2944,N_2305,N_2039);
xor U2945 (N_2945,N_2292,N_2283);
nor U2946 (N_2946,N_1700,N_1840);
nor U2947 (N_2947,N_2258,N_2004);
or U2948 (N_2948,N_1967,N_2049);
xnor U2949 (N_2949,N_2369,N_2216);
or U2950 (N_2950,N_2231,N_1906);
nand U2951 (N_2951,N_2222,N_2004);
and U2952 (N_2952,N_1694,N_1639);
and U2953 (N_2953,N_1805,N_2379);
and U2954 (N_2954,N_1854,N_1648);
nor U2955 (N_2955,N_2394,N_2272);
nor U2956 (N_2956,N_2220,N_2017);
xor U2957 (N_2957,N_2004,N_1605);
xor U2958 (N_2958,N_1661,N_1844);
or U2959 (N_2959,N_2280,N_1692);
nor U2960 (N_2960,N_2397,N_2321);
and U2961 (N_2961,N_1745,N_1710);
xnor U2962 (N_2962,N_1889,N_2193);
or U2963 (N_2963,N_2082,N_1643);
and U2964 (N_2964,N_1795,N_1990);
nor U2965 (N_2965,N_2241,N_1684);
xor U2966 (N_2966,N_1623,N_2282);
and U2967 (N_2967,N_1995,N_2109);
and U2968 (N_2968,N_1925,N_1921);
nor U2969 (N_2969,N_1716,N_1812);
xor U2970 (N_2970,N_2211,N_1685);
xor U2971 (N_2971,N_1774,N_1884);
nor U2972 (N_2972,N_1981,N_1687);
xnor U2973 (N_2973,N_2252,N_2082);
xnor U2974 (N_2974,N_1833,N_2070);
nand U2975 (N_2975,N_2311,N_2058);
nor U2976 (N_2976,N_2346,N_2159);
and U2977 (N_2977,N_1652,N_1686);
and U2978 (N_2978,N_2213,N_1806);
and U2979 (N_2979,N_2045,N_1816);
or U2980 (N_2980,N_2109,N_2117);
nand U2981 (N_2981,N_1750,N_1691);
xnor U2982 (N_2982,N_2177,N_2001);
and U2983 (N_2983,N_2264,N_2351);
nor U2984 (N_2984,N_2386,N_2299);
or U2985 (N_2985,N_2018,N_2261);
xnor U2986 (N_2986,N_2077,N_2297);
nand U2987 (N_2987,N_2326,N_1701);
or U2988 (N_2988,N_2349,N_2329);
nor U2989 (N_2989,N_2034,N_1667);
or U2990 (N_2990,N_1613,N_1635);
nor U2991 (N_2991,N_1881,N_2081);
xor U2992 (N_2992,N_2096,N_1805);
xnor U2993 (N_2993,N_2207,N_2330);
xnor U2994 (N_2994,N_1829,N_2096);
nor U2995 (N_2995,N_2123,N_1829);
nor U2996 (N_2996,N_1733,N_2101);
nor U2997 (N_2997,N_2066,N_1609);
or U2998 (N_2998,N_2265,N_2167);
or U2999 (N_2999,N_2118,N_1999);
nor U3000 (N_3000,N_2275,N_1758);
or U3001 (N_3001,N_2346,N_2024);
xor U3002 (N_3002,N_2395,N_2386);
nand U3003 (N_3003,N_2273,N_2122);
nand U3004 (N_3004,N_1726,N_2183);
nand U3005 (N_3005,N_2288,N_2082);
xnor U3006 (N_3006,N_2044,N_1791);
nand U3007 (N_3007,N_1745,N_1686);
nand U3008 (N_3008,N_1939,N_1685);
or U3009 (N_3009,N_1639,N_1922);
or U3010 (N_3010,N_2385,N_1960);
nor U3011 (N_3011,N_1843,N_1609);
xnor U3012 (N_3012,N_1913,N_2071);
or U3013 (N_3013,N_1957,N_1824);
xor U3014 (N_3014,N_2111,N_1634);
xnor U3015 (N_3015,N_1675,N_1937);
or U3016 (N_3016,N_1717,N_1854);
nand U3017 (N_3017,N_1610,N_1923);
nor U3018 (N_3018,N_1854,N_1901);
nor U3019 (N_3019,N_2191,N_1899);
xnor U3020 (N_3020,N_1819,N_2062);
nand U3021 (N_3021,N_1619,N_1868);
or U3022 (N_3022,N_2198,N_1773);
nand U3023 (N_3023,N_1717,N_1622);
or U3024 (N_3024,N_2390,N_2295);
nand U3025 (N_3025,N_1741,N_1896);
xnor U3026 (N_3026,N_2334,N_2226);
or U3027 (N_3027,N_2043,N_1698);
xor U3028 (N_3028,N_2037,N_2238);
and U3029 (N_3029,N_2302,N_1742);
and U3030 (N_3030,N_2333,N_2364);
nor U3031 (N_3031,N_1781,N_1924);
nor U3032 (N_3032,N_2076,N_2016);
or U3033 (N_3033,N_2158,N_1923);
or U3034 (N_3034,N_2018,N_2148);
nand U3035 (N_3035,N_2275,N_1763);
and U3036 (N_3036,N_2033,N_2068);
or U3037 (N_3037,N_2306,N_1986);
or U3038 (N_3038,N_1659,N_1604);
or U3039 (N_3039,N_1800,N_2003);
and U3040 (N_3040,N_2216,N_2328);
nor U3041 (N_3041,N_1976,N_1974);
or U3042 (N_3042,N_2110,N_2254);
nor U3043 (N_3043,N_2249,N_2168);
and U3044 (N_3044,N_2139,N_2126);
or U3045 (N_3045,N_2011,N_2123);
xnor U3046 (N_3046,N_2291,N_1646);
or U3047 (N_3047,N_1791,N_2385);
nor U3048 (N_3048,N_1738,N_1780);
and U3049 (N_3049,N_2104,N_2291);
or U3050 (N_3050,N_2043,N_2162);
xor U3051 (N_3051,N_2212,N_1749);
and U3052 (N_3052,N_2054,N_2226);
xor U3053 (N_3053,N_2296,N_1713);
nand U3054 (N_3054,N_1657,N_1661);
or U3055 (N_3055,N_2046,N_2055);
or U3056 (N_3056,N_1917,N_1770);
and U3057 (N_3057,N_1655,N_2214);
or U3058 (N_3058,N_2310,N_2130);
xor U3059 (N_3059,N_1854,N_1742);
nor U3060 (N_3060,N_1788,N_2123);
or U3061 (N_3061,N_1938,N_2368);
or U3062 (N_3062,N_2212,N_2252);
or U3063 (N_3063,N_1702,N_2299);
and U3064 (N_3064,N_1642,N_2198);
nand U3065 (N_3065,N_1958,N_2350);
xor U3066 (N_3066,N_2070,N_2035);
nand U3067 (N_3067,N_1973,N_1726);
and U3068 (N_3068,N_2116,N_2160);
xor U3069 (N_3069,N_1774,N_2142);
nor U3070 (N_3070,N_1908,N_2217);
or U3071 (N_3071,N_2026,N_1664);
or U3072 (N_3072,N_1768,N_2018);
nand U3073 (N_3073,N_2268,N_2089);
and U3074 (N_3074,N_1664,N_2048);
nor U3075 (N_3075,N_1757,N_1929);
and U3076 (N_3076,N_1737,N_2359);
or U3077 (N_3077,N_2365,N_1907);
and U3078 (N_3078,N_1730,N_2266);
nand U3079 (N_3079,N_1896,N_2001);
nand U3080 (N_3080,N_2090,N_1865);
or U3081 (N_3081,N_2016,N_1939);
xnor U3082 (N_3082,N_2289,N_2338);
xnor U3083 (N_3083,N_2358,N_1931);
xnor U3084 (N_3084,N_1759,N_1747);
and U3085 (N_3085,N_2063,N_1991);
nor U3086 (N_3086,N_1648,N_2200);
and U3087 (N_3087,N_2080,N_2045);
nand U3088 (N_3088,N_1988,N_2373);
nand U3089 (N_3089,N_2243,N_2082);
nor U3090 (N_3090,N_1917,N_2196);
and U3091 (N_3091,N_1815,N_1787);
and U3092 (N_3092,N_2166,N_2316);
or U3093 (N_3093,N_1988,N_2056);
and U3094 (N_3094,N_2324,N_1878);
xor U3095 (N_3095,N_2314,N_1900);
nand U3096 (N_3096,N_1977,N_1803);
or U3097 (N_3097,N_1925,N_1675);
xnor U3098 (N_3098,N_1775,N_2085);
xnor U3099 (N_3099,N_2335,N_1667);
and U3100 (N_3100,N_2028,N_2001);
nand U3101 (N_3101,N_2270,N_1921);
and U3102 (N_3102,N_2068,N_1950);
or U3103 (N_3103,N_2133,N_1852);
nand U3104 (N_3104,N_1678,N_2113);
xnor U3105 (N_3105,N_1831,N_2189);
nor U3106 (N_3106,N_2206,N_2269);
xor U3107 (N_3107,N_1636,N_1717);
or U3108 (N_3108,N_1782,N_2193);
nand U3109 (N_3109,N_1685,N_2259);
xor U3110 (N_3110,N_2078,N_2319);
xor U3111 (N_3111,N_1629,N_2165);
xor U3112 (N_3112,N_2310,N_2394);
nand U3113 (N_3113,N_1875,N_2295);
and U3114 (N_3114,N_2108,N_2181);
nand U3115 (N_3115,N_2243,N_2122);
or U3116 (N_3116,N_2089,N_2209);
and U3117 (N_3117,N_1892,N_2031);
nor U3118 (N_3118,N_2138,N_1888);
or U3119 (N_3119,N_1797,N_1656);
xor U3120 (N_3120,N_2063,N_1738);
xnor U3121 (N_3121,N_2279,N_2322);
or U3122 (N_3122,N_2214,N_1759);
nor U3123 (N_3123,N_2270,N_2217);
nor U3124 (N_3124,N_2307,N_1840);
or U3125 (N_3125,N_1602,N_2056);
nand U3126 (N_3126,N_2033,N_2102);
xnor U3127 (N_3127,N_1619,N_2388);
or U3128 (N_3128,N_2198,N_1824);
nand U3129 (N_3129,N_1685,N_2242);
and U3130 (N_3130,N_1659,N_1869);
xnor U3131 (N_3131,N_1923,N_1737);
and U3132 (N_3132,N_1961,N_1885);
nand U3133 (N_3133,N_1844,N_1620);
nand U3134 (N_3134,N_1942,N_1749);
nor U3135 (N_3135,N_1613,N_2274);
xor U3136 (N_3136,N_2154,N_1718);
or U3137 (N_3137,N_1848,N_2070);
and U3138 (N_3138,N_1710,N_2163);
and U3139 (N_3139,N_1759,N_1950);
or U3140 (N_3140,N_1970,N_1742);
and U3141 (N_3141,N_2124,N_2178);
and U3142 (N_3142,N_1881,N_1798);
and U3143 (N_3143,N_1862,N_2096);
nor U3144 (N_3144,N_1705,N_2393);
nor U3145 (N_3145,N_1772,N_1933);
and U3146 (N_3146,N_1898,N_2251);
nor U3147 (N_3147,N_1674,N_2259);
or U3148 (N_3148,N_1793,N_2230);
and U3149 (N_3149,N_2210,N_2193);
xor U3150 (N_3150,N_1603,N_1663);
or U3151 (N_3151,N_2208,N_1621);
nor U3152 (N_3152,N_2143,N_2307);
nor U3153 (N_3153,N_1680,N_1949);
nand U3154 (N_3154,N_1701,N_2364);
and U3155 (N_3155,N_2281,N_1921);
xnor U3156 (N_3156,N_2179,N_1640);
nor U3157 (N_3157,N_1898,N_2356);
nor U3158 (N_3158,N_2116,N_1984);
or U3159 (N_3159,N_2388,N_2259);
xor U3160 (N_3160,N_1718,N_1674);
nand U3161 (N_3161,N_2366,N_2382);
nor U3162 (N_3162,N_1661,N_1750);
and U3163 (N_3163,N_1707,N_2114);
or U3164 (N_3164,N_1773,N_1967);
and U3165 (N_3165,N_2378,N_1751);
nand U3166 (N_3166,N_2090,N_1751);
and U3167 (N_3167,N_1810,N_2064);
nor U3168 (N_3168,N_2260,N_1860);
nor U3169 (N_3169,N_1916,N_1960);
xnor U3170 (N_3170,N_1886,N_2201);
or U3171 (N_3171,N_2334,N_1615);
and U3172 (N_3172,N_2250,N_1887);
and U3173 (N_3173,N_2187,N_2126);
xor U3174 (N_3174,N_1977,N_1908);
and U3175 (N_3175,N_1713,N_1891);
or U3176 (N_3176,N_1969,N_2388);
or U3177 (N_3177,N_1998,N_2370);
xnor U3178 (N_3178,N_1909,N_2312);
and U3179 (N_3179,N_1938,N_2303);
and U3180 (N_3180,N_2275,N_2398);
nor U3181 (N_3181,N_1798,N_1800);
xor U3182 (N_3182,N_2361,N_1892);
nand U3183 (N_3183,N_1830,N_1858);
nand U3184 (N_3184,N_2167,N_1601);
or U3185 (N_3185,N_2278,N_2212);
or U3186 (N_3186,N_2086,N_1952);
nor U3187 (N_3187,N_1639,N_2227);
and U3188 (N_3188,N_1945,N_2393);
and U3189 (N_3189,N_1642,N_2027);
nand U3190 (N_3190,N_1706,N_1755);
or U3191 (N_3191,N_2145,N_2059);
nor U3192 (N_3192,N_2374,N_1731);
and U3193 (N_3193,N_1936,N_2359);
xor U3194 (N_3194,N_2212,N_2120);
nor U3195 (N_3195,N_2379,N_1678);
and U3196 (N_3196,N_2315,N_1789);
xnor U3197 (N_3197,N_2313,N_2256);
and U3198 (N_3198,N_1873,N_2355);
and U3199 (N_3199,N_2014,N_1924);
nand U3200 (N_3200,N_3193,N_2716);
or U3201 (N_3201,N_2894,N_2481);
nor U3202 (N_3202,N_2572,N_2406);
and U3203 (N_3203,N_3124,N_2565);
nand U3204 (N_3204,N_2689,N_2457);
and U3205 (N_3205,N_2499,N_2509);
nor U3206 (N_3206,N_2582,N_2775);
nand U3207 (N_3207,N_3022,N_3036);
and U3208 (N_3208,N_2806,N_3165);
nor U3209 (N_3209,N_2829,N_3192);
or U3210 (N_3210,N_2400,N_2488);
nand U3211 (N_3211,N_3043,N_2492);
xnor U3212 (N_3212,N_2997,N_2427);
nor U3213 (N_3213,N_2639,N_2432);
and U3214 (N_3214,N_3015,N_3111);
or U3215 (N_3215,N_2598,N_3176);
xnor U3216 (N_3216,N_2452,N_2464);
nor U3217 (N_3217,N_2984,N_2421);
or U3218 (N_3218,N_2907,N_3011);
and U3219 (N_3219,N_2743,N_2680);
or U3220 (N_3220,N_3026,N_3014);
nor U3221 (N_3221,N_2834,N_2665);
nor U3222 (N_3222,N_2948,N_3175);
nor U3223 (N_3223,N_2512,N_2470);
nand U3224 (N_3224,N_3119,N_3050);
and U3225 (N_3225,N_3006,N_2870);
nand U3226 (N_3226,N_2412,N_3062);
xor U3227 (N_3227,N_2749,N_3144);
nand U3228 (N_3228,N_2890,N_2578);
nor U3229 (N_3229,N_3186,N_2880);
nor U3230 (N_3230,N_2647,N_2947);
nor U3231 (N_3231,N_2570,N_3020);
and U3232 (N_3232,N_2757,N_3084);
nor U3233 (N_3233,N_2416,N_3105);
and U3234 (N_3234,N_2673,N_2623);
nand U3235 (N_3235,N_3117,N_2933);
and U3236 (N_3236,N_2869,N_2720);
or U3237 (N_3237,N_2698,N_2599);
xnor U3238 (N_3238,N_2762,N_2886);
nand U3239 (N_3239,N_3059,N_2558);
or U3240 (N_3240,N_2451,N_2681);
xnor U3241 (N_3241,N_2473,N_3179);
and U3242 (N_3242,N_2646,N_2955);
xor U3243 (N_3243,N_3005,N_2817);
xor U3244 (N_3244,N_2632,N_2779);
and U3245 (N_3245,N_2988,N_3085);
nor U3246 (N_3246,N_2706,N_2917);
nor U3247 (N_3247,N_3003,N_2959);
and U3248 (N_3248,N_3162,N_2508);
nor U3249 (N_3249,N_2874,N_3032);
and U3250 (N_3250,N_3143,N_2825);
or U3251 (N_3251,N_2543,N_3197);
nand U3252 (N_3252,N_2612,N_3095);
or U3253 (N_3253,N_2993,N_3149);
xor U3254 (N_3254,N_2807,N_2966);
and U3255 (N_3255,N_2652,N_3187);
nor U3256 (N_3256,N_2719,N_2651);
xor U3257 (N_3257,N_2745,N_3060);
xor U3258 (N_3258,N_3170,N_2977);
or U3259 (N_3259,N_2641,N_3053);
and U3260 (N_3260,N_2715,N_3129);
nor U3261 (N_3261,N_2844,N_2551);
nor U3262 (N_3262,N_2479,N_2628);
and U3263 (N_3263,N_2969,N_2645);
nand U3264 (N_3264,N_3068,N_2951);
xor U3265 (N_3265,N_2954,N_2631);
or U3266 (N_3266,N_2593,N_3035);
or U3267 (N_3267,N_2677,N_3183);
nand U3268 (N_3268,N_2945,N_2801);
nand U3269 (N_3269,N_2595,N_2401);
xor U3270 (N_3270,N_2973,N_3021);
nand U3271 (N_3271,N_2906,N_2795);
or U3272 (N_3272,N_2580,N_2617);
xor U3273 (N_3273,N_2876,N_2897);
and U3274 (N_3274,N_3133,N_3039);
nand U3275 (N_3275,N_3094,N_2546);
nor U3276 (N_3276,N_2547,N_2782);
nor U3277 (N_3277,N_2515,N_2517);
xnor U3278 (N_3278,N_2956,N_2804);
and U3279 (N_3279,N_3174,N_3097);
nand U3280 (N_3280,N_2530,N_2862);
nand U3281 (N_3281,N_2883,N_2563);
and U3282 (N_3282,N_2932,N_2621);
nor U3283 (N_3283,N_2867,N_2472);
and U3284 (N_3284,N_3077,N_2425);
and U3285 (N_3285,N_2912,N_2848);
nor U3286 (N_3286,N_2992,N_2723);
and U3287 (N_3287,N_2836,N_2591);
and U3288 (N_3288,N_2505,N_3100);
nand U3289 (N_3289,N_2532,N_2971);
nand U3290 (N_3290,N_3132,N_3161);
nor U3291 (N_3291,N_2523,N_2744);
xnor U3292 (N_3292,N_2675,N_2403);
or U3293 (N_3293,N_3109,N_2594);
or U3294 (N_3294,N_2695,N_2797);
xor U3295 (N_3295,N_3024,N_2624);
nor U3296 (N_3296,N_2748,N_2544);
nand U3297 (N_3297,N_2576,N_2989);
xor U3298 (N_3298,N_3103,N_2702);
nand U3299 (N_3299,N_2850,N_2958);
or U3300 (N_3300,N_2697,N_2724);
or U3301 (N_3301,N_2740,N_3028);
nor U3302 (N_3302,N_2751,N_2879);
nand U3303 (N_3303,N_2528,N_2980);
nand U3304 (N_3304,N_2990,N_2629);
and U3305 (N_3305,N_2655,N_2439);
nor U3306 (N_3306,N_2758,N_2468);
nand U3307 (N_3307,N_2601,N_2873);
xor U3308 (N_3308,N_2592,N_2686);
nand U3309 (N_3309,N_2929,N_3093);
nand U3310 (N_3310,N_2991,N_3061);
or U3311 (N_3311,N_2774,N_2960);
and U3312 (N_3312,N_2871,N_2760);
nor U3313 (N_3313,N_3155,N_2810);
and U3314 (N_3314,N_2538,N_3131);
xor U3315 (N_3315,N_2424,N_2767);
and U3316 (N_3316,N_2701,N_2627);
nand U3317 (N_3317,N_2577,N_2889);
nand U3318 (N_3318,N_3089,N_2750);
and U3319 (N_3319,N_2882,N_2409);
nand U3320 (N_3320,N_2562,N_2513);
nand U3321 (N_3321,N_3072,N_2666);
nor U3322 (N_3322,N_3065,N_3071);
and U3323 (N_3323,N_3184,N_2654);
xor U3324 (N_3324,N_2604,N_2430);
and U3325 (N_3325,N_2703,N_2957);
nand U3326 (N_3326,N_2502,N_2986);
nand U3327 (N_3327,N_2765,N_2625);
xnor U3328 (N_3328,N_2575,N_2545);
nand U3329 (N_3329,N_2742,N_2419);
nor U3330 (N_3330,N_2769,N_2461);
nor U3331 (N_3331,N_2794,N_2444);
xnor U3332 (N_3332,N_2438,N_2405);
nor U3333 (N_3333,N_3041,N_2792);
nand U3334 (N_3334,N_2927,N_2483);
and U3335 (N_3335,N_2507,N_3010);
and U3336 (N_3336,N_2459,N_2553);
nor U3337 (N_3337,N_2837,N_3181);
and U3338 (N_3338,N_2462,N_2437);
and U3339 (N_3339,N_2534,N_2476);
nand U3340 (N_3340,N_3090,N_2415);
or U3341 (N_3341,N_2814,N_2976);
or U3342 (N_3342,N_2773,N_2533);
and U3343 (N_3343,N_2633,N_2527);
nor U3344 (N_3344,N_2895,N_2478);
or U3345 (N_3345,N_2846,N_2953);
nand U3346 (N_3346,N_2610,N_2514);
nor U3347 (N_3347,N_2618,N_2501);
or U3348 (N_3348,N_3044,N_2656);
or U3349 (N_3349,N_2660,N_2949);
nor U3350 (N_3350,N_2766,N_2919);
or U3351 (N_3351,N_2474,N_2506);
and U3352 (N_3352,N_2995,N_3152);
and U3353 (N_3353,N_2460,N_3122);
and U3354 (N_3354,N_2410,N_2587);
and U3355 (N_3355,N_2496,N_2985);
nand U3356 (N_3356,N_2443,N_2950);
nor U3357 (N_3357,N_2497,N_2711);
or U3358 (N_3358,N_2830,N_2936);
or U3359 (N_3359,N_2519,N_2710);
nor U3360 (N_3360,N_3154,N_2752);
and U3361 (N_3361,N_3138,N_2448);
or U3362 (N_3362,N_2614,N_2649);
or U3363 (N_3363,N_2926,N_2634);
nor U3364 (N_3364,N_2759,N_3198);
and U3365 (N_3365,N_2608,N_2944);
nand U3366 (N_3366,N_2402,N_2664);
and U3367 (N_3367,N_2418,N_2754);
and U3368 (N_3368,N_2975,N_2809);
or U3369 (N_3369,N_2494,N_3185);
or U3370 (N_3370,N_2796,N_2999);
or U3371 (N_3371,N_2670,N_2861);
xor U3372 (N_3372,N_2454,N_2913);
and U3373 (N_3373,N_2974,N_2676);
and U3374 (N_3374,N_3025,N_3079);
xnor U3375 (N_3375,N_3126,N_3082);
nor U3376 (N_3376,N_3056,N_2480);
or U3377 (N_3377,N_2705,N_3023);
nor U3378 (N_3378,N_2511,N_3130);
or U3379 (N_3379,N_2484,N_2510);
nand U3380 (N_3380,N_2453,N_2735);
nor U3381 (N_3381,N_2613,N_2921);
nor U3382 (N_3382,N_3042,N_3037);
or U3383 (N_3383,N_2682,N_3054);
xnor U3384 (N_3384,N_2783,N_2838);
nor U3385 (N_3385,N_2653,N_3055);
xor U3386 (N_3386,N_2708,N_2832);
nand U3387 (N_3387,N_2812,N_3086);
nor U3388 (N_3388,N_2486,N_2685);
and U3389 (N_3389,N_2531,N_3146);
xor U3390 (N_3390,N_2901,N_2900);
nor U3391 (N_3391,N_2983,N_2722);
nand U3392 (N_3392,N_3167,N_3168);
nand U3393 (N_3393,N_2761,N_2691);
nand U3394 (N_3394,N_2630,N_3078);
nor U3395 (N_3395,N_3178,N_2777);
or U3396 (N_3396,N_2884,N_2855);
nor U3397 (N_3397,N_2994,N_2536);
or U3398 (N_3398,N_2586,N_3169);
nand U3399 (N_3399,N_3004,N_2585);
nor U3400 (N_3400,N_2588,N_2683);
xnor U3401 (N_3401,N_2941,N_2490);
and U3402 (N_3402,N_2658,N_3057);
xnor U3403 (N_3403,N_2542,N_3102);
nand U3404 (N_3404,N_2803,N_2772);
xnor U3405 (N_3405,N_2568,N_2668);
xor U3406 (N_3406,N_3172,N_2477);
nand U3407 (N_3407,N_2902,N_2408);
and U3408 (N_3408,N_2661,N_2690);
xnor U3409 (N_3409,N_2644,N_2996);
xor U3410 (N_3410,N_3074,N_2763);
or U3411 (N_3411,N_3016,N_2539);
nand U3412 (N_3412,N_2877,N_3110);
or U3413 (N_3413,N_2696,N_2564);
xnor U3414 (N_3414,N_3018,N_2747);
or U3415 (N_3415,N_2998,N_2467);
and U3416 (N_3416,N_2915,N_3098);
or U3417 (N_3417,N_2818,N_3134);
xnor U3418 (N_3418,N_2475,N_2916);
or U3419 (N_3419,N_2799,N_3153);
or U3420 (N_3420,N_2866,N_2831);
nand U3421 (N_3421,N_2434,N_2466);
nor U3422 (N_3422,N_2922,N_2860);
nor U3423 (N_3423,N_2560,N_2637);
xnor U3424 (N_3424,N_2442,N_2579);
and U3425 (N_3425,N_2914,N_2805);
and U3426 (N_3426,N_3148,N_2469);
nor U3427 (N_3427,N_2824,N_2800);
nand U3428 (N_3428,N_2819,N_3125);
or U3429 (N_3429,N_2962,N_2465);
xnor U3430 (N_3430,N_2554,N_2943);
xor U3431 (N_3431,N_3038,N_2878);
nand U3432 (N_3432,N_2516,N_2787);
nor U3433 (N_3433,N_2458,N_3151);
or U3434 (N_3434,N_3113,N_2573);
or U3435 (N_3435,N_2892,N_2764);
and U3436 (N_3436,N_2788,N_3066);
xor U3437 (N_3437,N_3017,N_3112);
and U3438 (N_3438,N_3145,N_3140);
and U3439 (N_3439,N_2663,N_3027);
xnor U3440 (N_3440,N_2781,N_3051);
xnor U3441 (N_3441,N_3069,N_3034);
nor U3442 (N_3442,N_2821,N_2569);
xor U3443 (N_3443,N_2640,N_2555);
nor U3444 (N_3444,N_2904,N_2839);
nand U3445 (N_3445,N_3121,N_2662);
nand U3446 (N_3446,N_2935,N_2650);
nand U3447 (N_3447,N_2854,N_2471);
xnor U3448 (N_3448,N_2433,N_3091);
and U3449 (N_3449,N_3101,N_2672);
or U3450 (N_3450,N_3157,N_3139);
xor U3451 (N_3451,N_2657,N_2537);
nor U3452 (N_3452,N_2669,N_2485);
xnor U3453 (N_3453,N_2648,N_3115);
nand U3454 (N_3454,N_2642,N_2768);
and U3455 (N_3455,N_2872,N_2887);
nand U3456 (N_3456,N_2445,N_2753);
xnor U3457 (N_3457,N_3158,N_2606);
xor U3458 (N_3458,N_2784,N_2626);
or U3459 (N_3459,N_3136,N_2487);
nor U3460 (N_3460,N_3083,N_3189);
or U3461 (N_3461,N_2937,N_3092);
nor U3462 (N_3462,N_2571,N_3118);
and U3463 (N_3463,N_2930,N_2728);
xor U3464 (N_3464,N_2611,N_2636);
nor U3465 (N_3465,N_2521,N_2808);
or U3466 (N_3466,N_2482,N_3019);
xor U3467 (N_3467,N_2789,N_2725);
nor U3468 (N_3468,N_2898,N_3029);
nor U3469 (N_3469,N_2940,N_2550);
and U3470 (N_3470,N_3166,N_2833);
and U3471 (N_3471,N_2726,N_2732);
nor U3472 (N_3472,N_2596,N_2423);
nor U3473 (N_3473,N_2712,N_2489);
nor U3474 (N_3474,N_2820,N_2491);
nor U3475 (N_3475,N_2847,N_3076);
nor U3476 (N_3476,N_2671,N_3047);
nand U3477 (N_3477,N_2548,N_3012);
or U3478 (N_3478,N_2731,N_2978);
and U3479 (N_3479,N_2590,N_2557);
or U3480 (N_3480,N_2863,N_2694);
xor U3481 (N_3481,N_2520,N_3045);
nand U3482 (N_3482,N_2456,N_3182);
nand U3483 (N_3483,N_2541,N_2455);
nor U3484 (N_3484,N_2852,N_2549);
nor U3485 (N_3485,N_2778,N_2559);
and U3486 (N_3486,N_2529,N_3164);
or U3487 (N_3487,N_2908,N_2891);
nand U3488 (N_3488,N_3081,N_2659);
and U3489 (N_3489,N_3195,N_2707);
nor U3490 (N_3490,N_2589,N_2620);
or U3491 (N_3491,N_2619,N_3088);
and U3492 (N_3492,N_2843,N_2981);
and U3493 (N_3493,N_2605,N_3052);
or U3494 (N_3494,N_2896,N_2845);
nor U3495 (N_3495,N_2426,N_2780);
nor U3496 (N_3496,N_3137,N_2450);
xor U3497 (N_3497,N_2828,N_2982);
or U3498 (N_3498,N_2964,N_2853);
nand U3499 (N_3499,N_2600,N_2667);
nor U3500 (N_3500,N_2756,N_2822);
xor U3501 (N_3501,N_2910,N_2737);
or U3502 (N_3502,N_2859,N_3160);
xnor U3503 (N_3503,N_2842,N_2811);
and U3504 (N_3504,N_2770,N_3190);
nor U3505 (N_3505,N_2552,N_2518);
and U3506 (N_3506,N_2771,N_2638);
nor U3507 (N_3507,N_2493,N_2584);
nor U3508 (N_3508,N_2905,N_2687);
or U3509 (N_3509,N_2404,N_2858);
nor U3510 (N_3510,N_3048,N_2823);
and U3511 (N_3511,N_2607,N_2911);
nor U3512 (N_3512,N_2721,N_2939);
nor U3513 (N_3513,N_2609,N_2734);
and U3514 (N_3514,N_2961,N_2498);
and U3515 (N_3515,N_2857,N_2500);
nand U3516 (N_3516,N_2597,N_2813);
xor U3517 (N_3517,N_3156,N_3128);
xnor U3518 (N_3518,N_3030,N_2411);
xor U3519 (N_3519,N_3087,N_3171);
nor U3520 (N_3520,N_2524,N_2925);
or U3521 (N_3521,N_2417,N_2709);
nand U3522 (N_3522,N_3046,N_3127);
nor U3523 (N_3523,N_2963,N_2567);
nor U3524 (N_3524,N_2826,N_3007);
and U3525 (N_3525,N_3141,N_3058);
nor U3526 (N_3526,N_3191,N_2463);
xor U3527 (N_3527,N_2965,N_2574);
and U3528 (N_3528,N_2888,N_2616);
or U3529 (N_3529,N_2979,N_2714);
xor U3530 (N_3530,N_3194,N_3135);
xor U3531 (N_3531,N_2918,N_3000);
and U3532 (N_3532,N_2840,N_3080);
nor U3533 (N_3533,N_2704,N_2909);
nand U3534 (N_3534,N_2736,N_2525);
or U3535 (N_3535,N_2688,N_2678);
xnor U3536 (N_3536,N_3147,N_3008);
xor U3537 (N_3537,N_3070,N_2755);
nand U3538 (N_3538,N_2970,N_2504);
xor U3539 (N_3539,N_2864,N_2622);
nand U3540 (N_3540,N_2968,N_2730);
or U3541 (N_3541,N_2713,N_2741);
and U3542 (N_3542,N_2440,N_2583);
or U3543 (N_3543,N_2946,N_2865);
xor U3544 (N_3544,N_2717,N_3163);
or U3545 (N_3545,N_2827,N_3123);
xor U3546 (N_3546,N_2700,N_2972);
nor U3547 (N_3547,N_2407,N_2738);
nand U3548 (N_3548,N_3108,N_2540);
xor U3549 (N_3549,N_2581,N_2449);
and U3550 (N_3550,N_2693,N_2987);
nand U3551 (N_3551,N_2718,N_2802);
nor U3552 (N_3552,N_3064,N_2739);
nor U3553 (N_3553,N_2815,N_2903);
nor U3554 (N_3554,N_2851,N_3002);
and U3555 (N_3555,N_3075,N_2495);
nand U3556 (N_3556,N_3009,N_2934);
and U3557 (N_3557,N_2893,N_2835);
nor U3558 (N_3558,N_2684,N_3114);
or U3559 (N_3559,N_2841,N_2413);
or U3560 (N_3560,N_2556,N_2422);
and U3561 (N_3561,N_3096,N_3107);
nand U3562 (N_3562,N_2436,N_3120);
xor U3563 (N_3563,N_2635,N_3150);
and U3564 (N_3564,N_3040,N_2643);
nand U3565 (N_3565,N_2566,N_2875);
nor U3566 (N_3566,N_2441,N_2733);
xor U3567 (N_3567,N_3063,N_2535);
nand U3568 (N_3568,N_2798,N_2791);
nor U3569 (N_3569,N_3067,N_3073);
or U3570 (N_3570,N_2431,N_2692);
xor U3571 (N_3571,N_2928,N_2920);
nand U3572 (N_3572,N_2931,N_3159);
nor U3573 (N_3573,N_2446,N_2420);
and U3574 (N_3574,N_2674,N_2856);
xor U3575 (N_3575,N_2938,N_2952);
or U3576 (N_3576,N_3013,N_3177);
nor U3577 (N_3577,N_2503,N_2429);
nand U3578 (N_3578,N_2923,N_2790);
nor U3579 (N_3579,N_2967,N_3049);
xor U3580 (N_3580,N_2786,N_3033);
and U3581 (N_3581,N_2885,N_2435);
and U3582 (N_3582,N_2615,N_3104);
and U3583 (N_3583,N_2522,N_2729);
xnor U3584 (N_3584,N_2816,N_2899);
nand U3585 (N_3585,N_3180,N_2561);
and U3586 (N_3586,N_2924,N_2447);
and U3587 (N_3587,N_3106,N_2603);
or U3588 (N_3588,N_3116,N_2868);
and U3589 (N_3589,N_3031,N_2776);
nand U3590 (N_3590,N_3196,N_2785);
and U3591 (N_3591,N_2526,N_2428);
nand U3592 (N_3592,N_2942,N_3001);
and U3593 (N_3593,N_2727,N_2793);
nand U3594 (N_3594,N_2414,N_2602);
nor U3595 (N_3595,N_2881,N_3173);
nor U3596 (N_3596,N_3099,N_3199);
and U3597 (N_3597,N_2699,N_3142);
nor U3598 (N_3598,N_2746,N_2849);
or U3599 (N_3599,N_2679,N_3188);
nor U3600 (N_3600,N_2419,N_2917);
nand U3601 (N_3601,N_3062,N_2713);
nor U3602 (N_3602,N_3171,N_2981);
xor U3603 (N_3603,N_3190,N_2610);
and U3604 (N_3604,N_3044,N_2480);
and U3605 (N_3605,N_3196,N_2557);
xor U3606 (N_3606,N_2415,N_2900);
and U3607 (N_3607,N_2631,N_2623);
xor U3608 (N_3608,N_2997,N_2484);
nand U3609 (N_3609,N_3170,N_2968);
nand U3610 (N_3610,N_2870,N_2835);
or U3611 (N_3611,N_2672,N_2540);
or U3612 (N_3612,N_3146,N_2425);
nand U3613 (N_3613,N_2633,N_2634);
nor U3614 (N_3614,N_3100,N_3197);
nand U3615 (N_3615,N_2530,N_2430);
nand U3616 (N_3616,N_2476,N_3199);
or U3617 (N_3617,N_2636,N_2822);
xor U3618 (N_3618,N_2990,N_2638);
nor U3619 (N_3619,N_2755,N_2498);
or U3620 (N_3620,N_2446,N_2850);
xor U3621 (N_3621,N_3189,N_3038);
and U3622 (N_3622,N_3157,N_2862);
nor U3623 (N_3623,N_3040,N_2864);
nand U3624 (N_3624,N_2947,N_3017);
xnor U3625 (N_3625,N_2626,N_2613);
nand U3626 (N_3626,N_2920,N_2690);
or U3627 (N_3627,N_2959,N_2965);
nor U3628 (N_3628,N_2990,N_2904);
or U3629 (N_3629,N_2467,N_3026);
or U3630 (N_3630,N_2591,N_2588);
or U3631 (N_3631,N_3193,N_3113);
nor U3632 (N_3632,N_3157,N_2692);
xnor U3633 (N_3633,N_2858,N_3138);
nor U3634 (N_3634,N_3059,N_3197);
nor U3635 (N_3635,N_2863,N_3183);
xor U3636 (N_3636,N_2741,N_2705);
and U3637 (N_3637,N_2830,N_2693);
xnor U3638 (N_3638,N_3095,N_3198);
xnor U3639 (N_3639,N_2847,N_3064);
nand U3640 (N_3640,N_2427,N_2555);
nand U3641 (N_3641,N_2531,N_2661);
or U3642 (N_3642,N_2946,N_2817);
nor U3643 (N_3643,N_2589,N_2523);
and U3644 (N_3644,N_3094,N_2960);
nor U3645 (N_3645,N_3140,N_2721);
or U3646 (N_3646,N_3117,N_2978);
nand U3647 (N_3647,N_2656,N_2942);
nor U3648 (N_3648,N_2540,N_3048);
nor U3649 (N_3649,N_2923,N_2874);
nor U3650 (N_3650,N_3039,N_3036);
nor U3651 (N_3651,N_2984,N_2516);
nor U3652 (N_3652,N_3068,N_2612);
or U3653 (N_3653,N_2646,N_2838);
xor U3654 (N_3654,N_2616,N_2774);
and U3655 (N_3655,N_2415,N_2606);
and U3656 (N_3656,N_2886,N_2933);
or U3657 (N_3657,N_3007,N_2579);
nand U3658 (N_3658,N_2915,N_2738);
nand U3659 (N_3659,N_3048,N_2639);
nor U3660 (N_3660,N_3038,N_3056);
nor U3661 (N_3661,N_3165,N_2802);
xor U3662 (N_3662,N_2519,N_3098);
nor U3663 (N_3663,N_2963,N_2635);
xnor U3664 (N_3664,N_2610,N_2866);
or U3665 (N_3665,N_2863,N_2859);
or U3666 (N_3666,N_2922,N_2764);
nor U3667 (N_3667,N_2929,N_2956);
nand U3668 (N_3668,N_2630,N_2651);
or U3669 (N_3669,N_2560,N_2835);
xor U3670 (N_3670,N_2609,N_2798);
and U3671 (N_3671,N_2796,N_2953);
nand U3672 (N_3672,N_2734,N_2668);
nor U3673 (N_3673,N_2670,N_2639);
nor U3674 (N_3674,N_2498,N_2773);
nor U3675 (N_3675,N_2930,N_2699);
or U3676 (N_3676,N_2660,N_3104);
nor U3677 (N_3677,N_2610,N_2844);
and U3678 (N_3678,N_2953,N_2417);
nand U3679 (N_3679,N_2762,N_2651);
or U3680 (N_3680,N_2614,N_2755);
xnor U3681 (N_3681,N_2423,N_2454);
or U3682 (N_3682,N_2741,N_3120);
nor U3683 (N_3683,N_2756,N_3023);
or U3684 (N_3684,N_2528,N_3118);
and U3685 (N_3685,N_2599,N_2491);
nor U3686 (N_3686,N_2742,N_2768);
nor U3687 (N_3687,N_2691,N_2596);
or U3688 (N_3688,N_2411,N_3035);
nor U3689 (N_3689,N_3099,N_2796);
xnor U3690 (N_3690,N_3146,N_2650);
nand U3691 (N_3691,N_2802,N_2760);
xor U3692 (N_3692,N_2662,N_3172);
or U3693 (N_3693,N_2616,N_2842);
and U3694 (N_3694,N_2938,N_3130);
xor U3695 (N_3695,N_3160,N_2761);
or U3696 (N_3696,N_2972,N_2592);
xnor U3697 (N_3697,N_2785,N_2419);
nand U3698 (N_3698,N_2971,N_2582);
or U3699 (N_3699,N_2818,N_2910);
or U3700 (N_3700,N_2998,N_2652);
xor U3701 (N_3701,N_3050,N_2681);
xor U3702 (N_3702,N_2557,N_2840);
and U3703 (N_3703,N_2529,N_2681);
xnor U3704 (N_3704,N_2707,N_3165);
and U3705 (N_3705,N_2423,N_2939);
nand U3706 (N_3706,N_2873,N_2716);
xnor U3707 (N_3707,N_2593,N_2551);
and U3708 (N_3708,N_2825,N_3091);
and U3709 (N_3709,N_2719,N_3000);
or U3710 (N_3710,N_2857,N_3136);
or U3711 (N_3711,N_2611,N_2463);
nand U3712 (N_3712,N_2758,N_3081);
and U3713 (N_3713,N_2908,N_2751);
nand U3714 (N_3714,N_2696,N_3154);
nand U3715 (N_3715,N_2940,N_2857);
nand U3716 (N_3716,N_2857,N_2730);
or U3717 (N_3717,N_2760,N_2781);
xnor U3718 (N_3718,N_2423,N_2734);
nor U3719 (N_3719,N_2966,N_2973);
xnor U3720 (N_3720,N_2832,N_3177);
and U3721 (N_3721,N_2646,N_3070);
nor U3722 (N_3722,N_2702,N_3012);
nand U3723 (N_3723,N_2607,N_2909);
nand U3724 (N_3724,N_3040,N_2622);
or U3725 (N_3725,N_3075,N_2684);
and U3726 (N_3726,N_2838,N_2686);
and U3727 (N_3727,N_2663,N_3125);
xor U3728 (N_3728,N_2671,N_3109);
nor U3729 (N_3729,N_2431,N_2557);
or U3730 (N_3730,N_2777,N_2510);
or U3731 (N_3731,N_3194,N_2504);
or U3732 (N_3732,N_2705,N_2638);
xnor U3733 (N_3733,N_3071,N_3197);
xor U3734 (N_3734,N_3046,N_2552);
nor U3735 (N_3735,N_3122,N_3047);
or U3736 (N_3736,N_3072,N_2572);
and U3737 (N_3737,N_2875,N_2934);
xor U3738 (N_3738,N_2855,N_2947);
nor U3739 (N_3739,N_3119,N_3117);
and U3740 (N_3740,N_2687,N_2793);
and U3741 (N_3741,N_2807,N_2956);
and U3742 (N_3742,N_2813,N_2947);
xor U3743 (N_3743,N_2922,N_3030);
xnor U3744 (N_3744,N_2492,N_2715);
nand U3745 (N_3745,N_2902,N_2979);
nor U3746 (N_3746,N_2880,N_2804);
nand U3747 (N_3747,N_2803,N_3146);
or U3748 (N_3748,N_3121,N_3157);
xnor U3749 (N_3749,N_3046,N_3124);
nor U3750 (N_3750,N_2977,N_2934);
and U3751 (N_3751,N_3012,N_3121);
or U3752 (N_3752,N_2987,N_2834);
xnor U3753 (N_3753,N_2726,N_3188);
nor U3754 (N_3754,N_2923,N_3128);
nand U3755 (N_3755,N_2664,N_2691);
and U3756 (N_3756,N_2896,N_2798);
or U3757 (N_3757,N_2638,N_2836);
or U3758 (N_3758,N_2666,N_3089);
and U3759 (N_3759,N_2932,N_2899);
or U3760 (N_3760,N_2672,N_2884);
xor U3761 (N_3761,N_2584,N_2587);
nand U3762 (N_3762,N_3166,N_2525);
or U3763 (N_3763,N_2882,N_3125);
nand U3764 (N_3764,N_2811,N_2775);
nand U3765 (N_3765,N_2478,N_2898);
nand U3766 (N_3766,N_2840,N_2989);
or U3767 (N_3767,N_3094,N_2506);
nor U3768 (N_3768,N_3061,N_2689);
nand U3769 (N_3769,N_3014,N_2826);
xnor U3770 (N_3770,N_2695,N_2721);
xnor U3771 (N_3771,N_2551,N_2470);
or U3772 (N_3772,N_2842,N_2722);
and U3773 (N_3773,N_3040,N_3124);
nand U3774 (N_3774,N_2876,N_3076);
nor U3775 (N_3775,N_3166,N_2775);
and U3776 (N_3776,N_2584,N_2526);
nand U3777 (N_3777,N_2606,N_3062);
and U3778 (N_3778,N_2700,N_2415);
nand U3779 (N_3779,N_2441,N_2510);
and U3780 (N_3780,N_2789,N_2446);
and U3781 (N_3781,N_3105,N_3161);
and U3782 (N_3782,N_3039,N_3031);
or U3783 (N_3783,N_2628,N_2591);
nor U3784 (N_3784,N_2951,N_3098);
xnor U3785 (N_3785,N_2699,N_2478);
xor U3786 (N_3786,N_2611,N_2688);
and U3787 (N_3787,N_3105,N_3148);
and U3788 (N_3788,N_2401,N_2865);
xnor U3789 (N_3789,N_2767,N_2784);
xnor U3790 (N_3790,N_3034,N_2804);
xor U3791 (N_3791,N_2622,N_2633);
and U3792 (N_3792,N_2485,N_2682);
nor U3793 (N_3793,N_3013,N_2627);
nand U3794 (N_3794,N_2894,N_2969);
nor U3795 (N_3795,N_3077,N_2623);
or U3796 (N_3796,N_3179,N_2577);
nor U3797 (N_3797,N_2685,N_2841);
nor U3798 (N_3798,N_3004,N_2576);
and U3799 (N_3799,N_2638,N_2855);
nor U3800 (N_3800,N_3118,N_2412);
nand U3801 (N_3801,N_2926,N_2792);
nand U3802 (N_3802,N_3081,N_2637);
and U3803 (N_3803,N_3139,N_3099);
nand U3804 (N_3804,N_2722,N_3072);
or U3805 (N_3805,N_2957,N_2462);
or U3806 (N_3806,N_2720,N_2882);
nand U3807 (N_3807,N_2797,N_2854);
and U3808 (N_3808,N_2820,N_2589);
xor U3809 (N_3809,N_2527,N_2913);
nor U3810 (N_3810,N_3022,N_2414);
nand U3811 (N_3811,N_2514,N_2956);
nand U3812 (N_3812,N_3062,N_3030);
xnor U3813 (N_3813,N_2863,N_2728);
nor U3814 (N_3814,N_3050,N_2875);
and U3815 (N_3815,N_2665,N_3026);
nor U3816 (N_3816,N_3006,N_3197);
and U3817 (N_3817,N_2529,N_2611);
or U3818 (N_3818,N_2693,N_2878);
or U3819 (N_3819,N_3011,N_2947);
or U3820 (N_3820,N_2692,N_3113);
nor U3821 (N_3821,N_2957,N_2550);
and U3822 (N_3822,N_3110,N_2735);
nor U3823 (N_3823,N_2743,N_3148);
xor U3824 (N_3824,N_2658,N_2419);
and U3825 (N_3825,N_2561,N_2641);
nor U3826 (N_3826,N_2885,N_2586);
xnor U3827 (N_3827,N_2756,N_2663);
nand U3828 (N_3828,N_2758,N_2823);
or U3829 (N_3829,N_2518,N_2455);
or U3830 (N_3830,N_3097,N_2621);
xor U3831 (N_3831,N_3151,N_2863);
xor U3832 (N_3832,N_2593,N_2955);
xor U3833 (N_3833,N_2469,N_2917);
or U3834 (N_3834,N_2704,N_2906);
nor U3835 (N_3835,N_2972,N_3151);
nand U3836 (N_3836,N_3155,N_2484);
xor U3837 (N_3837,N_3174,N_2648);
or U3838 (N_3838,N_3089,N_2562);
and U3839 (N_3839,N_2468,N_2707);
nor U3840 (N_3840,N_2868,N_2903);
nand U3841 (N_3841,N_2856,N_2846);
nor U3842 (N_3842,N_2944,N_3076);
or U3843 (N_3843,N_2542,N_2839);
nor U3844 (N_3844,N_2680,N_3093);
xor U3845 (N_3845,N_3170,N_2466);
xnor U3846 (N_3846,N_2766,N_2945);
nor U3847 (N_3847,N_2858,N_3121);
nor U3848 (N_3848,N_2449,N_3100);
nand U3849 (N_3849,N_2943,N_2847);
xor U3850 (N_3850,N_3007,N_2598);
xnor U3851 (N_3851,N_2639,N_2592);
and U3852 (N_3852,N_2951,N_3128);
or U3853 (N_3853,N_2905,N_2647);
nand U3854 (N_3854,N_3005,N_2809);
and U3855 (N_3855,N_2434,N_2755);
nor U3856 (N_3856,N_2754,N_2817);
nand U3857 (N_3857,N_2515,N_2519);
and U3858 (N_3858,N_2873,N_3106);
xor U3859 (N_3859,N_3093,N_2616);
nand U3860 (N_3860,N_2480,N_2630);
xnor U3861 (N_3861,N_2494,N_3072);
and U3862 (N_3862,N_2539,N_2522);
nor U3863 (N_3863,N_2680,N_2972);
xnor U3864 (N_3864,N_2844,N_3095);
nor U3865 (N_3865,N_2494,N_2802);
and U3866 (N_3866,N_3108,N_2487);
or U3867 (N_3867,N_2726,N_2489);
nand U3868 (N_3868,N_2518,N_3081);
xnor U3869 (N_3869,N_2970,N_2772);
nor U3870 (N_3870,N_2694,N_3053);
nand U3871 (N_3871,N_2594,N_2658);
nand U3872 (N_3872,N_2472,N_3172);
nor U3873 (N_3873,N_3011,N_2888);
xnor U3874 (N_3874,N_3006,N_2500);
nand U3875 (N_3875,N_3196,N_2881);
or U3876 (N_3876,N_3138,N_2647);
nor U3877 (N_3877,N_2751,N_2435);
xor U3878 (N_3878,N_3035,N_2892);
xnor U3879 (N_3879,N_2510,N_2555);
and U3880 (N_3880,N_3077,N_2935);
nor U3881 (N_3881,N_2563,N_2994);
nand U3882 (N_3882,N_2421,N_3021);
nand U3883 (N_3883,N_3088,N_2832);
and U3884 (N_3884,N_2798,N_2804);
nand U3885 (N_3885,N_2818,N_3107);
or U3886 (N_3886,N_2429,N_2659);
and U3887 (N_3887,N_2702,N_2742);
nor U3888 (N_3888,N_2629,N_3024);
nand U3889 (N_3889,N_2603,N_2528);
or U3890 (N_3890,N_2658,N_2549);
or U3891 (N_3891,N_3140,N_2859);
nor U3892 (N_3892,N_2940,N_2765);
xor U3893 (N_3893,N_2750,N_3032);
and U3894 (N_3894,N_2459,N_3093);
nand U3895 (N_3895,N_2788,N_2640);
xor U3896 (N_3896,N_2623,N_2416);
and U3897 (N_3897,N_2481,N_2727);
xnor U3898 (N_3898,N_2702,N_2686);
nor U3899 (N_3899,N_3027,N_2927);
and U3900 (N_3900,N_2636,N_2504);
nor U3901 (N_3901,N_2701,N_2730);
nand U3902 (N_3902,N_2443,N_3138);
nor U3903 (N_3903,N_2721,N_3007);
and U3904 (N_3904,N_2537,N_2603);
and U3905 (N_3905,N_2782,N_2705);
nor U3906 (N_3906,N_2886,N_3076);
and U3907 (N_3907,N_3089,N_2939);
or U3908 (N_3908,N_3116,N_2545);
xor U3909 (N_3909,N_2870,N_3034);
nand U3910 (N_3910,N_2607,N_2457);
nor U3911 (N_3911,N_3138,N_3187);
and U3912 (N_3912,N_2768,N_2688);
and U3913 (N_3913,N_2828,N_2602);
and U3914 (N_3914,N_2895,N_3051);
and U3915 (N_3915,N_2733,N_2967);
or U3916 (N_3916,N_3166,N_2976);
xnor U3917 (N_3917,N_3138,N_2779);
nor U3918 (N_3918,N_2787,N_2927);
or U3919 (N_3919,N_2951,N_2891);
nor U3920 (N_3920,N_3029,N_2447);
nor U3921 (N_3921,N_2507,N_2747);
or U3922 (N_3922,N_3195,N_3091);
or U3923 (N_3923,N_2901,N_2857);
or U3924 (N_3924,N_2403,N_2468);
xnor U3925 (N_3925,N_2894,N_2626);
and U3926 (N_3926,N_2937,N_2765);
or U3927 (N_3927,N_2823,N_2893);
or U3928 (N_3928,N_2569,N_2621);
nor U3929 (N_3929,N_2888,N_2861);
and U3930 (N_3930,N_3122,N_2593);
or U3931 (N_3931,N_2578,N_2496);
and U3932 (N_3932,N_2809,N_2897);
or U3933 (N_3933,N_2691,N_2594);
xor U3934 (N_3934,N_2911,N_3116);
and U3935 (N_3935,N_2490,N_2473);
xor U3936 (N_3936,N_3112,N_2809);
xnor U3937 (N_3937,N_2534,N_2923);
nor U3938 (N_3938,N_2930,N_3025);
xor U3939 (N_3939,N_2804,N_2572);
nand U3940 (N_3940,N_2787,N_3116);
xnor U3941 (N_3941,N_2450,N_2862);
nor U3942 (N_3942,N_2876,N_2402);
nand U3943 (N_3943,N_2454,N_3004);
or U3944 (N_3944,N_2866,N_2420);
and U3945 (N_3945,N_2416,N_2993);
or U3946 (N_3946,N_2661,N_3173);
or U3947 (N_3947,N_2442,N_3114);
and U3948 (N_3948,N_3070,N_2714);
and U3949 (N_3949,N_2787,N_2417);
xnor U3950 (N_3950,N_3043,N_2731);
and U3951 (N_3951,N_2908,N_3064);
or U3952 (N_3952,N_2756,N_2456);
and U3953 (N_3953,N_3159,N_2516);
nor U3954 (N_3954,N_2999,N_2632);
xnor U3955 (N_3955,N_3001,N_3075);
xnor U3956 (N_3956,N_2420,N_2909);
and U3957 (N_3957,N_2486,N_2402);
nor U3958 (N_3958,N_2856,N_2939);
nand U3959 (N_3959,N_2463,N_2700);
nor U3960 (N_3960,N_3143,N_2670);
nor U3961 (N_3961,N_3142,N_3080);
or U3962 (N_3962,N_2534,N_3052);
nor U3963 (N_3963,N_2682,N_2478);
nor U3964 (N_3964,N_2429,N_2549);
xor U3965 (N_3965,N_2401,N_2868);
xor U3966 (N_3966,N_2776,N_2927);
nand U3967 (N_3967,N_2644,N_2435);
and U3968 (N_3968,N_3155,N_2614);
and U3969 (N_3969,N_2827,N_3119);
nand U3970 (N_3970,N_2400,N_3050);
nor U3971 (N_3971,N_3111,N_2577);
nor U3972 (N_3972,N_2418,N_2464);
or U3973 (N_3973,N_3112,N_2810);
nor U3974 (N_3974,N_2596,N_2941);
nor U3975 (N_3975,N_3143,N_2400);
or U3976 (N_3976,N_3085,N_3007);
nor U3977 (N_3977,N_2556,N_2969);
or U3978 (N_3978,N_2813,N_2808);
nand U3979 (N_3979,N_2893,N_2906);
nand U3980 (N_3980,N_3156,N_2901);
xnor U3981 (N_3981,N_2712,N_3174);
xor U3982 (N_3982,N_2664,N_3013);
nand U3983 (N_3983,N_3115,N_2418);
and U3984 (N_3984,N_3139,N_3172);
nand U3985 (N_3985,N_2574,N_2931);
nor U3986 (N_3986,N_2731,N_2424);
xnor U3987 (N_3987,N_2796,N_2551);
xor U3988 (N_3988,N_3184,N_2548);
or U3989 (N_3989,N_2474,N_3138);
xor U3990 (N_3990,N_3127,N_2929);
or U3991 (N_3991,N_2424,N_3033);
xor U3992 (N_3992,N_3003,N_2753);
nor U3993 (N_3993,N_2566,N_3062);
nor U3994 (N_3994,N_3151,N_2613);
or U3995 (N_3995,N_3159,N_2857);
and U3996 (N_3996,N_3021,N_2728);
nand U3997 (N_3997,N_2945,N_2616);
and U3998 (N_3998,N_2569,N_2694);
or U3999 (N_3999,N_2495,N_2530);
and U4000 (N_4000,N_3310,N_3480);
xor U4001 (N_4001,N_3296,N_3616);
xor U4002 (N_4002,N_3309,N_3784);
xnor U4003 (N_4003,N_3311,N_3628);
and U4004 (N_4004,N_3284,N_3802);
xor U4005 (N_4005,N_3661,N_3958);
xor U4006 (N_4006,N_3876,N_3877);
xnor U4007 (N_4007,N_3439,N_3388);
nand U4008 (N_4008,N_3389,N_3582);
nor U4009 (N_4009,N_3673,N_3472);
or U4010 (N_4010,N_3593,N_3390);
or U4011 (N_4011,N_3627,N_3531);
and U4012 (N_4012,N_3222,N_3468);
and U4013 (N_4013,N_3230,N_3880);
or U4014 (N_4014,N_3568,N_3220);
nor U4015 (N_4015,N_3618,N_3935);
or U4016 (N_4016,N_3791,N_3996);
nand U4017 (N_4017,N_3214,N_3200);
xor U4018 (N_4018,N_3818,N_3423);
xor U4019 (N_4019,N_3779,N_3340);
or U4020 (N_4020,N_3333,N_3552);
and U4021 (N_4021,N_3519,N_3632);
nand U4022 (N_4022,N_3525,N_3303);
nand U4023 (N_4023,N_3831,N_3807);
or U4024 (N_4024,N_3271,N_3883);
nor U4025 (N_4025,N_3923,N_3477);
and U4026 (N_4026,N_3291,N_3799);
and U4027 (N_4027,N_3598,N_3538);
nand U4028 (N_4028,N_3660,N_3548);
nor U4029 (N_4029,N_3959,N_3909);
or U4030 (N_4030,N_3573,N_3971);
xnor U4031 (N_4031,N_3453,N_3621);
nand U4032 (N_4032,N_3858,N_3415);
nand U4033 (N_4033,N_3283,N_3341);
xnor U4034 (N_4034,N_3349,N_3938);
nand U4035 (N_4035,N_3240,N_3308);
or U4036 (N_4036,N_3555,N_3544);
nand U4037 (N_4037,N_3327,N_3307);
or U4038 (N_4038,N_3595,N_3947);
nand U4039 (N_4039,N_3788,N_3956);
and U4040 (N_4040,N_3288,N_3847);
xor U4041 (N_4041,N_3323,N_3738);
or U4042 (N_4042,N_3378,N_3462);
or U4043 (N_4043,N_3526,N_3980);
and U4044 (N_4044,N_3809,N_3910);
nor U4045 (N_4045,N_3920,N_3893);
nand U4046 (N_4046,N_3420,N_3700);
xor U4047 (N_4047,N_3780,N_3225);
or U4048 (N_4048,N_3489,N_3393);
and U4049 (N_4049,N_3437,N_3374);
nor U4050 (N_4050,N_3715,N_3726);
and U4051 (N_4051,N_3435,N_3773);
and U4052 (N_4052,N_3249,N_3617);
nand U4053 (N_4053,N_3662,N_3281);
nor U4054 (N_4054,N_3665,N_3387);
or U4055 (N_4055,N_3392,N_3895);
or U4056 (N_4056,N_3347,N_3916);
nor U4057 (N_4057,N_3745,N_3641);
or U4058 (N_4058,N_3949,N_3451);
or U4059 (N_4059,N_3360,N_3742);
nand U4060 (N_4060,N_3789,N_3457);
xnor U4061 (N_4061,N_3213,N_3238);
xor U4062 (N_4062,N_3533,N_3265);
or U4063 (N_4063,N_3691,N_3348);
or U4064 (N_4064,N_3454,N_3866);
xor U4065 (N_4065,N_3588,N_3962);
and U4066 (N_4066,N_3416,N_3523);
nor U4067 (N_4067,N_3253,N_3889);
xor U4068 (N_4068,N_3912,N_3864);
and U4069 (N_4069,N_3315,N_3482);
nor U4070 (N_4070,N_3888,N_3636);
nand U4071 (N_4071,N_3446,N_3564);
and U4072 (N_4072,N_3794,N_3845);
or U4073 (N_4073,N_3689,N_3695);
nor U4074 (N_4074,N_3272,N_3325);
xor U4075 (N_4075,N_3875,N_3856);
and U4076 (N_4076,N_3223,N_3928);
or U4077 (N_4077,N_3972,N_3776);
or U4078 (N_4078,N_3266,N_3502);
nand U4079 (N_4079,N_3467,N_3837);
nor U4080 (N_4080,N_3269,N_3306);
xnor U4081 (N_4081,N_3343,N_3994);
and U4082 (N_4082,N_3756,N_3406);
xor U4083 (N_4083,N_3841,N_3445);
nor U4084 (N_4084,N_3890,N_3361);
nand U4085 (N_4085,N_3478,N_3395);
xor U4086 (N_4086,N_3550,N_3903);
nand U4087 (N_4087,N_3924,N_3748);
xor U4088 (N_4088,N_3941,N_3512);
and U4089 (N_4089,N_3279,N_3666);
nor U4090 (N_4090,N_3373,N_3603);
xor U4091 (N_4091,N_3687,N_3997);
and U4092 (N_4092,N_3402,N_3797);
xnor U4093 (N_4093,N_3974,N_3945);
and U4094 (N_4094,N_3596,N_3535);
or U4095 (N_4095,N_3359,N_3609);
nand U4096 (N_4096,N_3849,N_3737);
and U4097 (N_4097,N_3473,N_3491);
and U4098 (N_4098,N_3625,N_3287);
xnor U4099 (N_4099,N_3940,N_3647);
or U4100 (N_4100,N_3624,N_3441);
xnor U4101 (N_4101,N_3576,N_3367);
and U4102 (N_4102,N_3954,N_3981);
nand U4103 (N_4103,N_3529,N_3694);
nand U4104 (N_4104,N_3668,N_3973);
nand U4105 (N_4105,N_3202,N_3417);
nor U4106 (N_4106,N_3411,N_3868);
and U4107 (N_4107,N_3886,N_3879);
nor U4108 (N_4108,N_3384,N_3346);
nand U4109 (N_4109,N_3887,N_3905);
xnor U4110 (N_4110,N_3514,N_3982);
nand U4111 (N_4111,N_3711,N_3644);
and U4112 (N_4112,N_3682,N_3551);
or U4113 (N_4113,N_3245,N_3534);
xor U4114 (N_4114,N_3696,N_3236);
xor U4115 (N_4115,N_3563,N_3513);
or U4116 (N_4116,N_3604,N_3581);
xnor U4117 (N_4117,N_3639,N_3561);
nand U4118 (N_4118,N_3842,N_3364);
nand U4119 (N_4119,N_3757,N_3219);
or U4120 (N_4120,N_3207,N_3319);
nand U4121 (N_4121,N_3460,N_3242);
nor U4122 (N_4122,N_3521,N_3256);
or U4123 (N_4123,N_3413,N_3605);
and U4124 (N_4124,N_3764,N_3464);
and U4125 (N_4125,N_3571,N_3444);
nand U4126 (N_4126,N_3226,N_3978);
nor U4127 (N_4127,N_3607,N_3828);
nand U4128 (N_4128,N_3851,N_3710);
and U4129 (N_4129,N_3509,N_3448);
or U4130 (N_4130,N_3730,N_3843);
nand U4131 (N_4131,N_3761,N_3804);
or U4132 (N_4132,N_3298,N_3400);
or U4133 (N_4133,N_3559,N_3721);
nand U4134 (N_4134,N_3999,N_3692);
or U4135 (N_4135,N_3530,N_3232);
xor U4136 (N_4136,N_3485,N_3690);
and U4137 (N_4137,N_3755,N_3570);
and U4138 (N_4138,N_3475,N_3998);
nand U4139 (N_4139,N_3774,N_3369);
or U4140 (N_4140,N_3456,N_3630);
xor U4141 (N_4141,N_3408,N_3925);
xnor U4142 (N_4142,N_3203,N_3931);
or U4143 (N_4143,N_3500,N_3950);
and U4144 (N_4144,N_3878,N_3208);
nor U4145 (N_4145,N_3645,N_3855);
nand U4146 (N_4146,N_3274,N_3718);
and U4147 (N_4147,N_3536,N_3589);
xor U4148 (N_4148,N_3227,N_3684);
and U4149 (N_4149,N_3313,N_3672);
nor U4150 (N_4150,N_3469,N_3587);
xnor U4151 (N_4151,N_3987,N_3305);
and U4152 (N_4152,N_3286,N_3520);
nor U4153 (N_4153,N_3741,N_3251);
or U4154 (N_4154,N_3643,N_3763);
or U4155 (N_4155,N_3729,N_3578);
nor U4156 (N_4156,N_3626,N_3653);
xnor U4157 (N_4157,N_3867,N_3394);
and U4158 (N_4158,N_3900,N_3246);
xnor U4159 (N_4159,N_3629,N_3404);
xor U4160 (N_4160,N_3966,N_3705);
xor U4161 (N_4161,N_3899,N_3270);
xnor U4162 (N_4162,N_3252,N_3591);
nand U4163 (N_4163,N_3833,N_3295);
nand U4164 (N_4164,N_3995,N_3678);
nor U4165 (N_4165,N_3993,N_3952);
nor U4166 (N_4166,N_3262,N_3934);
and U4167 (N_4167,N_3891,N_3777);
nand U4168 (N_4168,N_3902,N_3937);
nor U4169 (N_4169,N_3297,N_3335);
and U4170 (N_4170,N_3820,N_3345);
nand U4171 (N_4171,N_3594,N_3606);
or U4172 (N_4172,N_3583,N_3210);
nor U4173 (N_4173,N_3844,N_3671);
nand U4174 (N_4174,N_3930,N_3725);
xnor U4175 (N_4175,N_3810,N_3686);
nand U4176 (N_4176,N_3433,N_3549);
and U4177 (N_4177,N_3663,N_3352);
xor U4178 (N_4178,N_3259,N_3681);
nand U4179 (N_4179,N_3897,N_3328);
nand U4180 (N_4180,N_3990,N_3209);
nor U4181 (N_4181,N_3719,N_3939);
xnor U4182 (N_4182,N_3635,N_3403);
xnor U4183 (N_4183,N_3407,N_3870);
or U4184 (N_4184,N_3932,N_3892);
or U4185 (N_4185,N_3933,N_3562);
xor U4186 (N_4186,N_3834,N_3574);
xnor U4187 (N_4187,N_3470,N_3450);
nand U4188 (N_4188,N_3599,N_3459);
and U4189 (N_4189,N_3727,N_3339);
nand U4190 (N_4190,N_3546,N_3235);
nor U4191 (N_4191,N_3680,N_3915);
and U4192 (N_4192,N_3495,N_3722);
nor U4193 (N_4193,N_3428,N_3412);
nor U4194 (N_4194,N_3614,N_3613);
nand U4195 (N_4195,N_3946,N_3247);
or U4196 (N_4196,N_3557,N_3273);
and U4197 (N_4197,N_3965,N_3871);
and U4198 (N_4198,N_3803,N_3250);
or U4199 (N_4199,N_3720,N_3419);
or U4200 (N_4200,N_3991,N_3263);
and U4201 (N_4201,N_3753,N_3276);
xnor U4202 (N_4202,N_3267,N_3733);
nor U4203 (N_4203,N_3231,N_3282);
and U4204 (N_4204,N_3747,N_3466);
nand U4205 (N_4205,N_3221,N_3768);
nand U4206 (N_4206,N_3676,N_3703);
xnor U4207 (N_4207,N_3869,N_3398);
and U4208 (N_4208,N_3443,N_3507);
or U4209 (N_4209,N_3264,N_3813);
and U4210 (N_4210,N_3234,N_3829);
xor U4211 (N_4211,N_3430,N_3772);
or U4212 (N_4212,N_3432,N_3859);
or U4213 (N_4213,N_3292,N_3508);
xor U4214 (N_4214,N_3440,N_3642);
xnor U4215 (N_4215,N_3257,N_3382);
xor U4216 (N_4216,N_3438,N_3484);
or U4217 (N_4217,N_3840,N_3385);
or U4218 (N_4218,N_3836,N_3543);
and U4219 (N_4219,N_3960,N_3497);
nand U4220 (N_4220,N_3863,N_3471);
xor U4221 (N_4221,N_3656,N_3860);
nand U4222 (N_4222,N_3664,N_3537);
nand U4223 (N_4223,N_3294,N_3278);
and U4224 (N_4224,N_3754,N_3942);
nand U4225 (N_4225,N_3355,N_3351);
or U4226 (N_4226,N_3948,N_3233);
or U4227 (N_4227,N_3363,N_3850);
or U4228 (N_4228,N_3517,N_3280);
nand U4229 (N_4229,N_3814,N_3724);
nand U4230 (N_4230,N_3494,N_3631);
nor U4231 (N_4231,N_3674,N_3646);
xor U4232 (N_4232,N_3380,N_3806);
and U4233 (N_4233,N_3728,N_3565);
xnor U4234 (N_4234,N_3586,N_3827);
nand U4235 (N_4235,N_3553,N_3637);
and U4236 (N_4236,N_3884,N_3812);
xnor U4237 (N_4237,N_3781,N_3865);
nor U4238 (N_4238,N_3796,N_3356);
or U4239 (N_4239,N_3688,N_3401);
and U4240 (N_4240,N_3312,N_3699);
xor U4241 (N_4241,N_3760,N_3816);
xnor U4242 (N_4242,N_3611,N_3640);
and U4243 (N_4243,N_3683,N_3556);
xnor U4244 (N_4244,N_3775,N_3731);
nand U4245 (N_4245,N_3371,N_3846);
nor U4246 (N_4246,N_3409,N_3967);
xor U4247 (N_4247,N_3427,N_3874);
and U4248 (N_4248,N_3379,N_3904);
or U4249 (N_4249,N_3370,N_3410);
and U4250 (N_4250,N_3329,N_3712);
or U4251 (N_4251,N_3293,N_3449);
nand U4252 (N_4252,N_3669,N_3486);
nand U4253 (N_4253,N_3321,N_3650);
or U4254 (N_4254,N_3707,N_3698);
and U4255 (N_4255,N_3228,N_3602);
nand U4256 (N_4256,N_3391,N_3608);
nor U4257 (N_4257,N_3819,N_3505);
nor U4258 (N_4258,N_3572,N_3330);
or U4259 (N_4259,N_3798,N_3600);
nand U4260 (N_4260,N_3894,N_3334);
xor U4261 (N_4261,N_3824,N_3670);
and U4262 (N_4262,N_3815,N_3968);
or U4263 (N_4263,N_3984,N_3358);
nand U4264 (N_4264,N_3498,N_3717);
nor U4265 (N_4265,N_3597,N_3277);
xnor U4266 (N_4266,N_3396,N_3970);
nand U4267 (N_4267,N_3615,N_3744);
or U4268 (N_4268,N_3414,N_3218);
nand U4269 (N_4269,N_3386,N_3248);
or U4270 (N_4270,N_3988,N_3805);
and U4271 (N_4271,N_3376,N_3832);
and U4272 (N_4272,N_3911,N_3896);
or U4273 (N_4273,N_3260,N_3766);
nand U4274 (N_4274,N_3765,N_3584);
and U4275 (N_4275,N_3314,N_3241);
and U4276 (N_4276,N_3795,N_3811);
nor U4277 (N_4277,N_3927,N_3750);
nor U4278 (N_4278,N_3986,N_3778);
or U4279 (N_4279,N_3979,N_3547);
and U4280 (N_4280,N_3487,N_3872);
nand U4281 (N_4281,N_3357,N_3770);
xor U4282 (N_4282,N_3964,N_3585);
xor U4283 (N_4283,N_3490,N_3455);
xor U4284 (N_4284,N_3704,N_3316);
and U4285 (N_4285,N_3539,N_3590);
xor U4286 (N_4286,N_3337,N_3463);
nor U4287 (N_4287,N_3338,N_3215);
nor U4288 (N_4288,N_3709,N_3655);
nor U4289 (N_4289,N_3771,N_3793);
nand U4290 (N_4290,N_3383,N_3985);
or U4291 (N_4291,N_3504,N_3336);
and U4292 (N_4292,N_3677,N_3580);
and U4293 (N_4293,N_3649,N_3908);
nand U4294 (N_4294,N_3301,N_3476);
and U4295 (N_4295,N_3969,N_3268);
and U4296 (N_4296,N_3921,N_3567);
xnor U4297 (N_4297,N_3289,N_3917);
nand U4298 (N_4298,N_3483,N_3493);
or U4299 (N_4299,N_3751,N_3377);
and U4300 (N_4300,N_3542,N_3652);
nor U4301 (N_4301,N_3638,N_3425);
and U4302 (N_4302,N_3697,N_3826);
and U4303 (N_4303,N_3787,N_3918);
nand U4304 (N_4304,N_3322,N_3381);
and U4305 (N_4305,N_3511,N_3506);
and U4306 (N_4306,N_3975,N_3496);
or U4307 (N_4307,N_3285,N_3790);
nor U4308 (N_4308,N_3332,N_3461);
nand U4309 (N_4309,N_3205,N_3786);
or U4310 (N_4310,N_3667,N_3651);
and U4311 (N_4311,N_3399,N_3955);
nand U4312 (N_4312,N_3299,N_3206);
or U4313 (N_4313,N_3515,N_3619);
xnor U4314 (N_4314,N_3237,N_3622);
nor U4315 (N_4315,N_3421,N_3243);
nand U4316 (N_4316,N_3783,N_3524);
xnor U4317 (N_4317,N_3212,N_3953);
nor U4318 (N_4318,N_3375,N_3612);
or U4319 (N_4319,N_3882,N_3558);
nor U4320 (N_4320,N_3620,N_3488);
xor U4321 (N_4321,N_3579,N_3848);
nor U4322 (N_4322,N_3961,N_3426);
and U4323 (N_4323,N_3976,N_3481);
nor U4324 (N_4324,N_3749,N_3418);
nor U4325 (N_4325,N_3861,N_3634);
or U4326 (N_4326,N_3601,N_3326);
nand U4327 (N_4327,N_3397,N_3424);
nor U4328 (N_4328,N_3901,N_3648);
and U4329 (N_4329,N_3839,N_3881);
and U4330 (N_4330,N_3821,N_3767);
xor U4331 (N_4331,N_3857,N_3769);
or U4332 (N_4332,N_3914,N_3659);
xnor U4333 (N_4333,N_3522,N_3532);
nand U4334 (N_4334,N_3835,N_3782);
and U4335 (N_4335,N_3541,N_3474);
nor U4336 (N_4336,N_3610,N_3342);
xor U4337 (N_4337,N_3290,N_3317);
or U4338 (N_4338,N_3229,N_3762);
xnor U4339 (N_4339,N_3957,N_3479);
or U4340 (N_4340,N_3331,N_3685);
nor U4341 (N_4341,N_3224,N_3800);
nand U4342 (N_4342,N_3943,N_3785);
or U4343 (N_4343,N_3736,N_3254);
or U4344 (N_4344,N_3442,N_3633);
xor U4345 (N_4345,N_3714,N_3708);
nand U4346 (N_4346,N_3977,N_3862);
nand U4347 (N_4347,N_3239,N_3431);
nor U4348 (N_4348,N_3854,N_3658);
or U4349 (N_4349,N_3362,N_3405);
or U4350 (N_4350,N_3906,N_3354);
nor U4351 (N_4351,N_3740,N_3907);
nand U4352 (N_4352,N_3554,N_3706);
xnor U4353 (N_4353,N_3716,N_3510);
and U4354 (N_4354,N_3734,N_3752);
nor U4355 (N_4355,N_3913,N_3853);
nor U4356 (N_4356,N_3429,N_3577);
nand U4357 (N_4357,N_3739,N_3372);
nor U4358 (N_4358,N_3300,N_3992);
xnor U4359 (N_4359,N_3759,N_3304);
nand U4360 (N_4360,N_3365,N_3353);
xnor U4361 (N_4361,N_3919,N_3560);
nand U4362 (N_4362,N_3452,N_3693);
or U4363 (N_4363,N_3702,N_3320);
or U4364 (N_4364,N_3873,N_3929);
and U4365 (N_4365,N_3735,N_3492);
nor U4366 (N_4366,N_3723,N_3566);
nand U4367 (N_4367,N_3302,N_3261);
and U4368 (N_4368,N_3258,N_3528);
or U4369 (N_4369,N_3623,N_3255);
nand U4370 (N_4370,N_3654,N_3575);
xnor U4371 (N_4371,N_3434,N_3545);
nor U4372 (N_4372,N_3808,N_3713);
and U4373 (N_4373,N_3458,N_3885);
and U4374 (N_4374,N_3244,N_3324);
or U4375 (N_4375,N_3540,N_3825);
and U4376 (N_4376,N_3936,N_3679);
nor U4377 (N_4377,N_3499,N_3518);
xor U4378 (N_4378,N_3922,N_3217);
or U4379 (N_4379,N_3822,N_3823);
xor U4380 (N_4380,N_3830,N_3447);
or U4381 (N_4381,N_3792,N_3465);
nand U4382 (N_4382,N_3675,N_3743);
and U4383 (N_4383,N_3503,N_3983);
and U4384 (N_4384,N_3732,N_3366);
nand U4385 (N_4385,N_3758,N_3204);
and U4386 (N_4386,N_3592,N_3527);
nand U4387 (N_4387,N_3852,N_3746);
xnor U4388 (N_4388,N_3275,N_3963);
xnor U4389 (N_4389,N_3368,N_3350);
xor U4390 (N_4390,N_3989,N_3201);
nor U4391 (N_4391,N_3926,N_3344);
nand U4392 (N_4392,N_3951,N_3516);
xor U4393 (N_4393,N_3501,N_3838);
and U4394 (N_4394,N_3216,N_3898);
xnor U4395 (N_4395,N_3569,N_3657);
nor U4396 (N_4396,N_3436,N_3944);
or U4397 (N_4397,N_3318,N_3817);
or U4398 (N_4398,N_3801,N_3701);
xnor U4399 (N_4399,N_3422,N_3211);
xor U4400 (N_4400,N_3359,N_3905);
nor U4401 (N_4401,N_3320,N_3340);
nand U4402 (N_4402,N_3436,N_3662);
and U4403 (N_4403,N_3718,N_3367);
nand U4404 (N_4404,N_3532,N_3737);
nand U4405 (N_4405,N_3682,N_3400);
xnor U4406 (N_4406,N_3591,N_3426);
nor U4407 (N_4407,N_3533,N_3434);
nor U4408 (N_4408,N_3701,N_3798);
xnor U4409 (N_4409,N_3690,N_3568);
and U4410 (N_4410,N_3326,N_3558);
xnor U4411 (N_4411,N_3843,N_3749);
xnor U4412 (N_4412,N_3796,N_3802);
nor U4413 (N_4413,N_3569,N_3656);
xor U4414 (N_4414,N_3375,N_3570);
or U4415 (N_4415,N_3283,N_3908);
or U4416 (N_4416,N_3659,N_3872);
nor U4417 (N_4417,N_3968,N_3670);
and U4418 (N_4418,N_3568,N_3504);
or U4419 (N_4419,N_3842,N_3751);
nor U4420 (N_4420,N_3632,N_3286);
or U4421 (N_4421,N_3846,N_3445);
and U4422 (N_4422,N_3597,N_3475);
xor U4423 (N_4423,N_3870,N_3463);
nor U4424 (N_4424,N_3588,N_3859);
nor U4425 (N_4425,N_3881,N_3740);
or U4426 (N_4426,N_3310,N_3410);
nor U4427 (N_4427,N_3674,N_3527);
xor U4428 (N_4428,N_3544,N_3493);
nand U4429 (N_4429,N_3986,N_3496);
or U4430 (N_4430,N_3427,N_3221);
and U4431 (N_4431,N_3401,N_3881);
nand U4432 (N_4432,N_3951,N_3203);
nor U4433 (N_4433,N_3575,N_3820);
and U4434 (N_4434,N_3957,N_3447);
xor U4435 (N_4435,N_3267,N_3482);
or U4436 (N_4436,N_3793,N_3779);
nor U4437 (N_4437,N_3458,N_3886);
or U4438 (N_4438,N_3613,N_3841);
nand U4439 (N_4439,N_3253,N_3997);
or U4440 (N_4440,N_3903,N_3842);
and U4441 (N_4441,N_3501,N_3259);
nor U4442 (N_4442,N_3788,N_3281);
nand U4443 (N_4443,N_3927,N_3645);
nand U4444 (N_4444,N_3796,N_3715);
and U4445 (N_4445,N_3909,N_3578);
or U4446 (N_4446,N_3676,N_3686);
or U4447 (N_4447,N_3911,N_3881);
or U4448 (N_4448,N_3304,N_3437);
or U4449 (N_4449,N_3755,N_3886);
and U4450 (N_4450,N_3244,N_3823);
and U4451 (N_4451,N_3668,N_3769);
and U4452 (N_4452,N_3858,N_3864);
or U4453 (N_4453,N_3334,N_3481);
nand U4454 (N_4454,N_3768,N_3759);
and U4455 (N_4455,N_3682,N_3421);
xor U4456 (N_4456,N_3744,N_3806);
or U4457 (N_4457,N_3773,N_3415);
nand U4458 (N_4458,N_3454,N_3867);
xor U4459 (N_4459,N_3548,N_3447);
or U4460 (N_4460,N_3515,N_3536);
xnor U4461 (N_4461,N_3456,N_3653);
nor U4462 (N_4462,N_3844,N_3929);
nand U4463 (N_4463,N_3992,N_3715);
xor U4464 (N_4464,N_3999,N_3222);
nand U4465 (N_4465,N_3559,N_3308);
or U4466 (N_4466,N_3227,N_3311);
nand U4467 (N_4467,N_3224,N_3649);
nor U4468 (N_4468,N_3513,N_3800);
and U4469 (N_4469,N_3261,N_3479);
nor U4470 (N_4470,N_3394,N_3322);
nor U4471 (N_4471,N_3342,N_3202);
xnor U4472 (N_4472,N_3987,N_3430);
nor U4473 (N_4473,N_3570,N_3830);
xor U4474 (N_4474,N_3217,N_3740);
and U4475 (N_4475,N_3284,N_3210);
nor U4476 (N_4476,N_3232,N_3592);
and U4477 (N_4477,N_3612,N_3378);
xnor U4478 (N_4478,N_3658,N_3370);
and U4479 (N_4479,N_3753,N_3911);
and U4480 (N_4480,N_3632,N_3320);
nor U4481 (N_4481,N_3795,N_3942);
nor U4482 (N_4482,N_3644,N_3996);
or U4483 (N_4483,N_3761,N_3775);
xor U4484 (N_4484,N_3326,N_3441);
xnor U4485 (N_4485,N_3827,N_3763);
nor U4486 (N_4486,N_3915,N_3662);
nand U4487 (N_4487,N_3334,N_3399);
nand U4488 (N_4488,N_3737,N_3676);
xor U4489 (N_4489,N_3698,N_3376);
or U4490 (N_4490,N_3669,N_3946);
or U4491 (N_4491,N_3892,N_3817);
xnor U4492 (N_4492,N_3249,N_3386);
nor U4493 (N_4493,N_3626,N_3752);
xor U4494 (N_4494,N_3409,N_3465);
or U4495 (N_4495,N_3686,N_3790);
or U4496 (N_4496,N_3582,N_3466);
xor U4497 (N_4497,N_3441,N_3987);
nor U4498 (N_4498,N_3942,N_3519);
or U4499 (N_4499,N_3782,N_3319);
nor U4500 (N_4500,N_3564,N_3288);
xor U4501 (N_4501,N_3630,N_3526);
xnor U4502 (N_4502,N_3264,N_3772);
or U4503 (N_4503,N_3829,N_3773);
or U4504 (N_4504,N_3796,N_3296);
or U4505 (N_4505,N_3598,N_3890);
and U4506 (N_4506,N_3350,N_3838);
nor U4507 (N_4507,N_3287,N_3808);
nor U4508 (N_4508,N_3936,N_3829);
nor U4509 (N_4509,N_3642,N_3737);
nor U4510 (N_4510,N_3872,N_3204);
nor U4511 (N_4511,N_3336,N_3694);
nor U4512 (N_4512,N_3829,N_3298);
and U4513 (N_4513,N_3422,N_3954);
nor U4514 (N_4514,N_3547,N_3606);
and U4515 (N_4515,N_3739,N_3361);
or U4516 (N_4516,N_3953,N_3622);
or U4517 (N_4517,N_3300,N_3349);
xor U4518 (N_4518,N_3707,N_3951);
nand U4519 (N_4519,N_3398,N_3309);
nor U4520 (N_4520,N_3367,N_3669);
xor U4521 (N_4521,N_3693,N_3622);
nor U4522 (N_4522,N_3929,N_3424);
nor U4523 (N_4523,N_3852,N_3245);
nand U4524 (N_4524,N_3885,N_3419);
nor U4525 (N_4525,N_3560,N_3910);
nor U4526 (N_4526,N_3622,N_3308);
or U4527 (N_4527,N_3522,N_3429);
or U4528 (N_4528,N_3440,N_3452);
xor U4529 (N_4529,N_3247,N_3270);
nand U4530 (N_4530,N_3316,N_3688);
or U4531 (N_4531,N_3529,N_3850);
nand U4532 (N_4532,N_3933,N_3744);
and U4533 (N_4533,N_3675,N_3280);
and U4534 (N_4534,N_3736,N_3364);
nand U4535 (N_4535,N_3302,N_3434);
nor U4536 (N_4536,N_3723,N_3817);
or U4537 (N_4537,N_3306,N_3245);
or U4538 (N_4538,N_3772,N_3794);
or U4539 (N_4539,N_3461,N_3717);
or U4540 (N_4540,N_3457,N_3797);
and U4541 (N_4541,N_3670,N_3281);
and U4542 (N_4542,N_3891,N_3491);
xor U4543 (N_4543,N_3654,N_3579);
and U4544 (N_4544,N_3803,N_3883);
and U4545 (N_4545,N_3885,N_3673);
or U4546 (N_4546,N_3687,N_3864);
nand U4547 (N_4547,N_3665,N_3991);
and U4548 (N_4548,N_3892,N_3847);
and U4549 (N_4549,N_3989,N_3211);
and U4550 (N_4550,N_3522,N_3356);
nand U4551 (N_4551,N_3287,N_3264);
xnor U4552 (N_4552,N_3942,N_3294);
or U4553 (N_4553,N_3943,N_3381);
or U4554 (N_4554,N_3475,N_3463);
and U4555 (N_4555,N_3548,N_3811);
or U4556 (N_4556,N_3884,N_3284);
and U4557 (N_4557,N_3667,N_3633);
xnor U4558 (N_4558,N_3649,N_3886);
nor U4559 (N_4559,N_3445,N_3716);
or U4560 (N_4560,N_3718,N_3535);
nor U4561 (N_4561,N_3991,N_3747);
xnor U4562 (N_4562,N_3968,N_3464);
nor U4563 (N_4563,N_3509,N_3601);
nor U4564 (N_4564,N_3983,N_3751);
or U4565 (N_4565,N_3570,N_3351);
nor U4566 (N_4566,N_3511,N_3428);
nor U4567 (N_4567,N_3577,N_3434);
xnor U4568 (N_4568,N_3483,N_3806);
or U4569 (N_4569,N_3918,N_3618);
or U4570 (N_4570,N_3867,N_3396);
or U4571 (N_4571,N_3713,N_3218);
nor U4572 (N_4572,N_3457,N_3901);
or U4573 (N_4573,N_3301,N_3709);
or U4574 (N_4574,N_3256,N_3804);
nand U4575 (N_4575,N_3868,N_3832);
or U4576 (N_4576,N_3650,N_3431);
nor U4577 (N_4577,N_3919,N_3446);
and U4578 (N_4578,N_3949,N_3956);
and U4579 (N_4579,N_3802,N_3969);
and U4580 (N_4580,N_3696,N_3378);
nand U4581 (N_4581,N_3416,N_3472);
nor U4582 (N_4582,N_3686,N_3982);
xor U4583 (N_4583,N_3706,N_3839);
or U4584 (N_4584,N_3689,N_3727);
xnor U4585 (N_4585,N_3424,N_3609);
and U4586 (N_4586,N_3223,N_3435);
nand U4587 (N_4587,N_3432,N_3513);
nand U4588 (N_4588,N_3279,N_3920);
xor U4589 (N_4589,N_3928,N_3815);
xnor U4590 (N_4590,N_3752,N_3796);
or U4591 (N_4591,N_3518,N_3991);
and U4592 (N_4592,N_3246,N_3933);
or U4593 (N_4593,N_3542,N_3699);
or U4594 (N_4594,N_3484,N_3804);
xor U4595 (N_4595,N_3908,N_3464);
nor U4596 (N_4596,N_3552,N_3988);
xor U4597 (N_4597,N_3893,N_3938);
and U4598 (N_4598,N_3358,N_3233);
xnor U4599 (N_4599,N_3855,N_3469);
or U4600 (N_4600,N_3384,N_3389);
nand U4601 (N_4601,N_3427,N_3469);
or U4602 (N_4602,N_3236,N_3717);
nand U4603 (N_4603,N_3515,N_3455);
xor U4604 (N_4604,N_3602,N_3821);
and U4605 (N_4605,N_3677,N_3941);
or U4606 (N_4606,N_3695,N_3481);
or U4607 (N_4607,N_3774,N_3428);
or U4608 (N_4608,N_3566,N_3542);
xor U4609 (N_4609,N_3396,N_3518);
xor U4610 (N_4610,N_3779,N_3943);
xor U4611 (N_4611,N_3496,N_3905);
xor U4612 (N_4612,N_3320,N_3349);
and U4613 (N_4613,N_3290,N_3634);
nand U4614 (N_4614,N_3289,N_3544);
nor U4615 (N_4615,N_3479,N_3433);
nand U4616 (N_4616,N_3387,N_3256);
and U4617 (N_4617,N_3307,N_3722);
nor U4618 (N_4618,N_3278,N_3969);
or U4619 (N_4619,N_3568,N_3694);
nand U4620 (N_4620,N_3791,N_3343);
nor U4621 (N_4621,N_3766,N_3749);
nand U4622 (N_4622,N_3311,N_3314);
nand U4623 (N_4623,N_3672,N_3296);
nor U4624 (N_4624,N_3933,N_3301);
or U4625 (N_4625,N_3466,N_3356);
and U4626 (N_4626,N_3890,N_3847);
and U4627 (N_4627,N_3761,N_3851);
nor U4628 (N_4628,N_3864,N_3204);
and U4629 (N_4629,N_3366,N_3867);
xnor U4630 (N_4630,N_3336,N_3738);
xnor U4631 (N_4631,N_3813,N_3740);
or U4632 (N_4632,N_3427,N_3764);
nor U4633 (N_4633,N_3658,N_3619);
and U4634 (N_4634,N_3265,N_3712);
or U4635 (N_4635,N_3339,N_3922);
and U4636 (N_4636,N_3510,N_3371);
xnor U4637 (N_4637,N_3759,N_3432);
and U4638 (N_4638,N_3867,N_3631);
or U4639 (N_4639,N_3226,N_3582);
nand U4640 (N_4640,N_3759,N_3819);
and U4641 (N_4641,N_3312,N_3705);
and U4642 (N_4642,N_3720,N_3963);
nand U4643 (N_4643,N_3340,N_3363);
nand U4644 (N_4644,N_3524,N_3260);
nand U4645 (N_4645,N_3979,N_3482);
or U4646 (N_4646,N_3798,N_3620);
and U4647 (N_4647,N_3285,N_3217);
nand U4648 (N_4648,N_3939,N_3444);
xnor U4649 (N_4649,N_3611,N_3375);
and U4650 (N_4650,N_3783,N_3518);
and U4651 (N_4651,N_3881,N_3855);
nand U4652 (N_4652,N_3934,N_3410);
nand U4653 (N_4653,N_3220,N_3669);
and U4654 (N_4654,N_3713,N_3604);
xor U4655 (N_4655,N_3855,N_3208);
xnor U4656 (N_4656,N_3746,N_3863);
xor U4657 (N_4657,N_3933,N_3643);
and U4658 (N_4658,N_3809,N_3680);
nand U4659 (N_4659,N_3891,N_3947);
nand U4660 (N_4660,N_3494,N_3268);
nand U4661 (N_4661,N_3682,N_3289);
or U4662 (N_4662,N_3389,N_3668);
nand U4663 (N_4663,N_3876,N_3277);
xor U4664 (N_4664,N_3476,N_3381);
nor U4665 (N_4665,N_3386,N_3430);
xnor U4666 (N_4666,N_3204,N_3429);
and U4667 (N_4667,N_3736,N_3938);
nor U4668 (N_4668,N_3429,N_3319);
nand U4669 (N_4669,N_3289,N_3388);
nor U4670 (N_4670,N_3996,N_3753);
and U4671 (N_4671,N_3240,N_3704);
nor U4672 (N_4672,N_3660,N_3409);
nand U4673 (N_4673,N_3526,N_3984);
nor U4674 (N_4674,N_3514,N_3302);
nand U4675 (N_4675,N_3372,N_3331);
or U4676 (N_4676,N_3971,N_3231);
and U4677 (N_4677,N_3731,N_3202);
nor U4678 (N_4678,N_3224,N_3438);
and U4679 (N_4679,N_3748,N_3703);
nor U4680 (N_4680,N_3405,N_3269);
or U4681 (N_4681,N_3642,N_3621);
and U4682 (N_4682,N_3912,N_3687);
nor U4683 (N_4683,N_3749,N_3781);
nor U4684 (N_4684,N_3427,N_3432);
xnor U4685 (N_4685,N_3649,N_3628);
nor U4686 (N_4686,N_3614,N_3997);
xor U4687 (N_4687,N_3404,N_3607);
nor U4688 (N_4688,N_3610,N_3270);
nor U4689 (N_4689,N_3558,N_3626);
xnor U4690 (N_4690,N_3625,N_3594);
and U4691 (N_4691,N_3756,N_3532);
and U4692 (N_4692,N_3430,N_3309);
nand U4693 (N_4693,N_3321,N_3577);
and U4694 (N_4694,N_3991,N_3724);
nand U4695 (N_4695,N_3793,N_3336);
or U4696 (N_4696,N_3675,N_3403);
or U4697 (N_4697,N_3954,N_3313);
nand U4698 (N_4698,N_3410,N_3459);
or U4699 (N_4699,N_3907,N_3727);
or U4700 (N_4700,N_3878,N_3497);
and U4701 (N_4701,N_3250,N_3791);
and U4702 (N_4702,N_3555,N_3999);
nand U4703 (N_4703,N_3223,N_3710);
and U4704 (N_4704,N_3950,N_3780);
nor U4705 (N_4705,N_3744,N_3888);
xor U4706 (N_4706,N_3264,N_3644);
nand U4707 (N_4707,N_3654,N_3231);
or U4708 (N_4708,N_3494,N_3734);
nand U4709 (N_4709,N_3663,N_3485);
or U4710 (N_4710,N_3295,N_3741);
or U4711 (N_4711,N_3561,N_3414);
nor U4712 (N_4712,N_3540,N_3971);
and U4713 (N_4713,N_3530,N_3635);
and U4714 (N_4714,N_3882,N_3834);
or U4715 (N_4715,N_3615,N_3425);
nor U4716 (N_4716,N_3469,N_3290);
nand U4717 (N_4717,N_3291,N_3672);
xor U4718 (N_4718,N_3257,N_3381);
or U4719 (N_4719,N_3743,N_3355);
and U4720 (N_4720,N_3663,N_3746);
nor U4721 (N_4721,N_3691,N_3575);
nor U4722 (N_4722,N_3263,N_3948);
nand U4723 (N_4723,N_3545,N_3456);
nor U4724 (N_4724,N_3585,N_3747);
xor U4725 (N_4725,N_3583,N_3627);
nand U4726 (N_4726,N_3826,N_3369);
and U4727 (N_4727,N_3557,N_3391);
nand U4728 (N_4728,N_3419,N_3290);
nand U4729 (N_4729,N_3829,N_3735);
xnor U4730 (N_4730,N_3621,N_3229);
nand U4731 (N_4731,N_3806,N_3444);
nand U4732 (N_4732,N_3404,N_3702);
nor U4733 (N_4733,N_3630,N_3909);
xnor U4734 (N_4734,N_3257,N_3396);
and U4735 (N_4735,N_3929,N_3535);
or U4736 (N_4736,N_3663,N_3662);
nor U4737 (N_4737,N_3298,N_3317);
nor U4738 (N_4738,N_3835,N_3635);
xor U4739 (N_4739,N_3895,N_3674);
or U4740 (N_4740,N_3721,N_3793);
nor U4741 (N_4741,N_3303,N_3312);
nand U4742 (N_4742,N_3889,N_3439);
nor U4743 (N_4743,N_3708,N_3493);
or U4744 (N_4744,N_3667,N_3621);
nand U4745 (N_4745,N_3239,N_3969);
xnor U4746 (N_4746,N_3552,N_3706);
xnor U4747 (N_4747,N_3783,N_3706);
or U4748 (N_4748,N_3767,N_3337);
or U4749 (N_4749,N_3881,N_3549);
or U4750 (N_4750,N_3747,N_3376);
and U4751 (N_4751,N_3700,N_3438);
or U4752 (N_4752,N_3438,N_3940);
nor U4753 (N_4753,N_3971,N_3994);
xor U4754 (N_4754,N_3469,N_3770);
xor U4755 (N_4755,N_3935,N_3267);
nand U4756 (N_4756,N_3291,N_3908);
or U4757 (N_4757,N_3616,N_3884);
xnor U4758 (N_4758,N_3896,N_3514);
nor U4759 (N_4759,N_3443,N_3730);
and U4760 (N_4760,N_3811,N_3928);
xor U4761 (N_4761,N_3752,N_3995);
and U4762 (N_4762,N_3761,N_3386);
nor U4763 (N_4763,N_3860,N_3496);
nand U4764 (N_4764,N_3236,N_3342);
or U4765 (N_4765,N_3538,N_3344);
nor U4766 (N_4766,N_3271,N_3258);
and U4767 (N_4767,N_3705,N_3790);
and U4768 (N_4768,N_3866,N_3411);
xor U4769 (N_4769,N_3447,N_3415);
and U4770 (N_4770,N_3686,N_3869);
xor U4771 (N_4771,N_3936,N_3591);
nor U4772 (N_4772,N_3232,N_3999);
and U4773 (N_4773,N_3829,N_3554);
xnor U4774 (N_4774,N_3845,N_3273);
and U4775 (N_4775,N_3619,N_3294);
or U4776 (N_4776,N_3933,N_3471);
nor U4777 (N_4777,N_3860,N_3377);
nand U4778 (N_4778,N_3599,N_3375);
or U4779 (N_4779,N_3793,N_3219);
or U4780 (N_4780,N_3719,N_3769);
xor U4781 (N_4781,N_3262,N_3666);
and U4782 (N_4782,N_3769,N_3695);
or U4783 (N_4783,N_3934,N_3962);
or U4784 (N_4784,N_3546,N_3920);
nand U4785 (N_4785,N_3392,N_3560);
or U4786 (N_4786,N_3224,N_3708);
nand U4787 (N_4787,N_3480,N_3235);
or U4788 (N_4788,N_3261,N_3652);
and U4789 (N_4789,N_3253,N_3576);
xor U4790 (N_4790,N_3892,N_3226);
nor U4791 (N_4791,N_3563,N_3830);
nor U4792 (N_4792,N_3841,N_3771);
nand U4793 (N_4793,N_3226,N_3916);
nor U4794 (N_4794,N_3830,N_3966);
nand U4795 (N_4795,N_3448,N_3825);
xor U4796 (N_4796,N_3965,N_3868);
nand U4797 (N_4797,N_3963,N_3777);
nor U4798 (N_4798,N_3600,N_3613);
xnor U4799 (N_4799,N_3835,N_3354);
nand U4800 (N_4800,N_4779,N_4278);
nor U4801 (N_4801,N_4211,N_4052);
xor U4802 (N_4802,N_4545,N_4064);
and U4803 (N_4803,N_4678,N_4653);
and U4804 (N_4804,N_4160,N_4726);
nand U4805 (N_4805,N_4373,N_4690);
nand U4806 (N_4806,N_4667,N_4352);
nand U4807 (N_4807,N_4047,N_4424);
nand U4808 (N_4808,N_4712,N_4129);
nand U4809 (N_4809,N_4038,N_4378);
nand U4810 (N_4810,N_4055,N_4008);
nand U4811 (N_4811,N_4463,N_4084);
nor U4812 (N_4812,N_4434,N_4670);
or U4813 (N_4813,N_4203,N_4229);
and U4814 (N_4814,N_4236,N_4010);
nand U4815 (N_4815,N_4723,N_4207);
and U4816 (N_4816,N_4391,N_4078);
nor U4817 (N_4817,N_4384,N_4441);
xor U4818 (N_4818,N_4784,N_4113);
nand U4819 (N_4819,N_4320,N_4359);
nand U4820 (N_4820,N_4597,N_4327);
nand U4821 (N_4821,N_4218,N_4367);
nor U4822 (N_4822,N_4529,N_4165);
nand U4823 (N_4823,N_4612,N_4224);
and U4824 (N_4824,N_4354,N_4348);
nand U4825 (N_4825,N_4011,N_4479);
nand U4826 (N_4826,N_4400,N_4628);
xnor U4827 (N_4827,N_4654,N_4213);
nor U4828 (N_4828,N_4114,N_4520);
or U4829 (N_4829,N_4040,N_4000);
xnor U4830 (N_4830,N_4402,N_4554);
nor U4831 (N_4831,N_4250,N_4004);
nand U4832 (N_4832,N_4599,N_4618);
nor U4833 (N_4833,N_4567,N_4413);
nand U4834 (N_4834,N_4194,N_4027);
or U4835 (N_4835,N_4575,N_4738);
nand U4836 (N_4836,N_4157,N_4288);
or U4837 (N_4837,N_4321,N_4731);
or U4838 (N_4838,N_4460,N_4550);
nor U4839 (N_4839,N_4673,N_4684);
and U4840 (N_4840,N_4363,N_4353);
xor U4841 (N_4841,N_4683,N_4528);
nand U4842 (N_4842,N_4467,N_4089);
and U4843 (N_4843,N_4462,N_4499);
nand U4844 (N_4844,N_4765,N_4332);
xor U4845 (N_4845,N_4298,N_4709);
and U4846 (N_4846,N_4660,N_4209);
xor U4847 (N_4847,N_4759,N_4261);
or U4848 (N_4848,N_4007,N_4455);
or U4849 (N_4849,N_4063,N_4539);
xnor U4850 (N_4850,N_4620,N_4590);
nand U4851 (N_4851,N_4217,N_4589);
or U4852 (N_4852,N_4262,N_4243);
xor U4853 (N_4853,N_4118,N_4150);
and U4854 (N_4854,N_4170,N_4631);
nor U4855 (N_4855,N_4741,N_4372);
xnor U4856 (N_4856,N_4360,N_4715);
nor U4857 (N_4857,N_4076,N_4331);
xnor U4858 (N_4858,N_4535,N_4146);
xor U4859 (N_4859,N_4097,N_4502);
xor U4860 (N_4860,N_4613,N_4191);
nor U4861 (N_4861,N_4306,N_4763);
nand U4862 (N_4862,N_4050,N_4214);
nand U4863 (N_4863,N_4205,N_4263);
and U4864 (N_4864,N_4583,N_4592);
or U4865 (N_4865,N_4094,N_4552);
or U4866 (N_4866,N_4451,N_4785);
xor U4867 (N_4867,N_4702,N_4220);
or U4868 (N_4868,N_4130,N_4742);
xor U4869 (N_4869,N_4268,N_4517);
nor U4870 (N_4870,N_4296,N_4031);
xor U4871 (N_4871,N_4423,N_4225);
nand U4872 (N_4872,N_4131,N_4281);
nor U4873 (N_4873,N_4365,N_4440);
nor U4874 (N_4874,N_4798,N_4411);
and U4875 (N_4875,N_4069,N_4501);
nor U4876 (N_4876,N_4248,N_4761);
or U4877 (N_4877,N_4795,N_4641);
xnor U4878 (N_4878,N_4573,N_4208);
xnor U4879 (N_4879,N_4181,N_4270);
xor U4880 (N_4880,N_4062,N_4048);
or U4881 (N_4881,N_4221,N_4231);
nor U4882 (N_4882,N_4565,N_4777);
and U4883 (N_4883,N_4092,N_4238);
xor U4884 (N_4884,N_4143,N_4497);
nand U4885 (N_4885,N_4744,N_4662);
and U4886 (N_4886,N_4188,N_4012);
nand U4887 (N_4887,N_4334,N_4669);
xnor U4888 (N_4888,N_4553,N_4184);
nand U4889 (N_4889,N_4246,N_4161);
or U4890 (N_4890,N_4681,N_4691);
or U4891 (N_4891,N_4021,N_4228);
or U4892 (N_4892,N_4601,N_4791);
nand U4893 (N_4893,N_4075,N_4190);
or U4894 (N_4894,N_4526,N_4685);
and U4895 (N_4895,N_4605,N_4388);
nand U4896 (N_4896,N_4252,N_4736);
and U4897 (N_4897,N_4456,N_4676);
nand U4898 (N_4898,N_4540,N_4587);
or U4899 (N_4899,N_4057,N_4664);
nand U4900 (N_4900,N_4381,N_4090);
nand U4901 (N_4901,N_4557,N_4323);
or U4902 (N_4902,N_4609,N_4408);
xnor U4903 (N_4903,N_4469,N_4254);
xnor U4904 (N_4904,N_4555,N_4340);
nand U4905 (N_4905,N_4346,N_4304);
nand U4906 (N_4906,N_4493,N_4677);
and U4907 (N_4907,N_4235,N_4457);
nor U4908 (N_4908,N_4284,N_4722);
or U4909 (N_4909,N_4755,N_4659);
xnor U4910 (N_4910,N_4748,N_4036);
or U4911 (N_4911,N_4128,N_4632);
or U4912 (N_4912,N_4415,N_4156);
nand U4913 (N_4913,N_4516,N_4171);
and U4914 (N_4914,N_4562,N_4449);
xor U4915 (N_4915,N_4275,N_4571);
and U4916 (N_4916,N_4109,N_4172);
nand U4917 (N_4917,N_4596,N_4148);
and U4918 (N_4918,N_4120,N_4387);
and U4919 (N_4919,N_4368,N_4029);
nor U4920 (N_4920,N_4576,N_4616);
xor U4921 (N_4921,N_4200,N_4087);
nor U4922 (N_4922,N_4705,N_4082);
nor U4923 (N_4923,N_4149,N_4450);
xor U4924 (N_4924,N_4395,N_4427);
or U4925 (N_4925,N_4239,N_4538);
nor U4926 (N_4926,N_4543,N_4778);
xnor U4927 (N_4927,N_4291,N_4470);
xor U4928 (N_4928,N_4285,N_4277);
nand U4929 (N_4929,N_4260,N_4524);
and U4930 (N_4930,N_4672,N_4037);
and U4931 (N_4931,N_4014,N_4333);
or U4932 (N_4932,N_4081,N_4006);
and U4933 (N_4933,N_4637,N_4431);
nor U4934 (N_4934,N_4650,N_4532);
nand U4935 (N_4935,N_4005,N_4189);
nand U4936 (N_4936,N_4490,N_4241);
or U4937 (N_4937,N_4794,N_4775);
and U4938 (N_4938,N_4797,N_4743);
xor U4939 (N_4939,N_4776,N_4175);
and U4940 (N_4940,N_4474,N_4439);
xnor U4941 (N_4941,N_4177,N_4649);
xor U4942 (N_4942,N_4510,N_4152);
or U4943 (N_4943,N_4139,N_4494);
or U4944 (N_4944,N_4174,N_4032);
and U4945 (N_4945,N_4013,N_4369);
or U4946 (N_4946,N_4593,N_4694);
nand U4947 (N_4947,N_4760,N_4397);
nor U4948 (N_4948,N_4077,N_4316);
or U4949 (N_4949,N_4586,N_4735);
nand U4950 (N_4950,N_4247,N_4318);
or U4951 (N_4951,N_4477,N_4046);
xor U4952 (N_4952,N_4399,N_4065);
nor U4953 (N_4953,N_4122,N_4386);
xnor U4954 (N_4954,N_4404,N_4787);
nand U4955 (N_4955,N_4781,N_4717);
or U4956 (N_4956,N_4527,N_4123);
xor U4957 (N_4957,N_4106,N_4508);
nor U4958 (N_4958,N_4215,N_4375);
or U4959 (N_4959,N_4602,N_4519);
xor U4960 (N_4960,N_4624,N_4324);
xor U4961 (N_4961,N_4071,N_4192);
xor U4962 (N_4962,N_4135,N_4251);
nor U4963 (N_4963,N_4648,N_4651);
or U4964 (N_4964,N_4054,N_4196);
nand U4965 (N_4965,N_4671,N_4448);
nand U4966 (N_4966,N_4701,N_4144);
nand U4967 (N_4967,N_4198,N_4083);
xor U4968 (N_4968,N_4603,N_4530);
or U4969 (N_4969,N_4766,N_4230);
nand U4970 (N_4970,N_4015,N_4799);
or U4971 (N_4971,N_4452,N_4138);
nor U4972 (N_4972,N_4729,N_4419);
nor U4973 (N_4973,N_4344,N_4206);
xnor U4974 (N_4974,N_4564,N_4472);
nor U4975 (N_4975,N_4234,N_4614);
and U4976 (N_4976,N_4336,N_4572);
nand U4977 (N_4977,N_4416,N_4356);
nand U4978 (N_4978,N_4574,N_4295);
nand U4979 (N_4979,N_4764,N_4699);
nand U4980 (N_4980,N_4403,N_4745);
xnor U4981 (N_4981,N_4721,N_4266);
xor U4982 (N_4982,N_4405,N_4060);
or U4983 (N_4983,N_4242,N_4183);
nor U4984 (N_4984,N_4500,N_4533);
or U4985 (N_4985,N_4204,N_4219);
or U4986 (N_4986,N_4633,N_4070);
nand U4987 (N_4987,N_4740,N_4115);
nor U4988 (N_4988,N_4433,N_4271);
xnor U4989 (N_4989,N_4039,N_4447);
nand U4990 (N_4990,N_4737,N_4301);
and U4991 (N_4991,N_4394,N_4623);
and U4992 (N_4992,N_4210,N_4410);
and U4993 (N_4993,N_4442,N_4134);
xor U4994 (N_4994,N_4088,N_4119);
nor U4995 (N_4995,N_4317,N_4734);
or U4996 (N_4996,N_4244,N_4259);
and U4997 (N_4997,N_4137,N_4542);
nand U4998 (N_4998,N_4700,N_4513);
xnor U4999 (N_4999,N_4111,N_4361);
xor U5000 (N_5000,N_4329,N_4444);
nand U5001 (N_5001,N_4626,N_4607);
nor U5002 (N_5002,N_4511,N_4293);
or U5003 (N_5003,N_4697,N_4068);
and U5004 (N_5004,N_4313,N_4549);
nor U5005 (N_5005,N_4663,N_4409);
and U5006 (N_5006,N_4199,N_4674);
xor U5007 (N_5007,N_4237,N_4132);
nand U5008 (N_5008,N_4158,N_4269);
and U5009 (N_5009,N_4780,N_4028);
or U5010 (N_5010,N_4746,N_4719);
or U5011 (N_5011,N_4406,N_4757);
nand U5012 (N_5012,N_4556,N_4773);
nor U5013 (N_5013,N_4099,N_4756);
xnor U5014 (N_5014,N_4059,N_4370);
or U5015 (N_5015,N_4026,N_4655);
and U5016 (N_5016,N_4488,N_4461);
or U5017 (N_5017,N_4483,N_4223);
nand U5018 (N_5018,N_4287,N_4311);
nor U5019 (N_5019,N_4617,N_4514);
nand U5020 (N_5020,N_4752,N_4661);
nand U5021 (N_5021,N_4274,N_4292);
nor U5022 (N_5022,N_4125,N_4024);
or U5023 (N_5023,N_4578,N_4117);
nor U5024 (N_5024,N_4053,N_4695);
xor U5025 (N_5025,N_4636,N_4162);
xor U5026 (N_5026,N_4796,N_4300);
nor U5027 (N_5027,N_4468,N_4487);
xnor U5028 (N_5028,N_4001,N_4546);
nand U5029 (N_5029,N_4051,N_4093);
xor U5030 (N_5030,N_4645,N_4257);
nand U5031 (N_5031,N_4226,N_4704);
xnor U5032 (N_5032,N_4591,N_4393);
nor U5033 (N_5033,N_4622,N_4019);
and U5034 (N_5034,N_4627,N_4445);
nand U5035 (N_5035,N_4080,N_4711);
and U5036 (N_5036,N_4561,N_4625);
nor U5037 (N_5037,N_4197,N_4579);
nor U5038 (N_5038,N_4728,N_4446);
nor U5039 (N_5039,N_4345,N_4437);
xor U5040 (N_5040,N_4768,N_4018);
xor U5041 (N_5041,N_4595,N_4429);
nor U5042 (N_5042,N_4767,N_4642);
or U5043 (N_5043,N_4035,N_4716);
xor U5044 (N_5044,N_4147,N_4585);
and U5045 (N_5045,N_4104,N_4072);
or U5046 (N_5046,N_4466,N_4145);
and U5047 (N_5047,N_4558,N_4568);
and U5048 (N_5048,N_4309,N_4272);
or U5049 (N_5049,N_4264,N_4687);
xnor U5050 (N_5050,N_4305,N_4164);
xor U5051 (N_5051,N_4202,N_4392);
and U5052 (N_5052,N_4339,N_4376);
or U5053 (N_5053,N_4710,N_4112);
nor U5054 (N_5054,N_4465,N_4430);
nor U5055 (N_5055,N_4688,N_4294);
and U5056 (N_5056,N_4280,N_4140);
or U5057 (N_5057,N_4049,N_4279);
xnor U5058 (N_5058,N_4116,N_4212);
nand U5059 (N_5059,N_4398,N_4600);
nand U5060 (N_5060,N_4666,N_4030);
and U5061 (N_5061,N_4091,N_4017);
or U5062 (N_5062,N_4426,N_4095);
nand U5063 (N_5063,N_4594,N_4495);
and U5064 (N_5064,N_4482,N_4315);
or U5065 (N_5065,N_4362,N_4136);
or U5066 (N_5066,N_4638,N_4176);
and U5067 (N_5067,N_4707,N_4232);
nand U5068 (N_5068,N_4619,N_4536);
and U5069 (N_5069,N_4185,N_4282);
nand U5070 (N_5070,N_4749,N_4686);
nor U5071 (N_5071,N_4696,N_4267);
or U5072 (N_5072,N_4486,N_4730);
xnor U5073 (N_5073,N_4753,N_4581);
and U5074 (N_5074,N_4350,N_4286);
nor U5075 (N_5075,N_4066,N_4283);
or U5076 (N_5076,N_4703,N_4180);
nand U5077 (N_5077,N_4725,N_4016);
xor U5078 (N_5078,N_4698,N_4163);
nand U5079 (N_5079,N_4382,N_4258);
xnor U5080 (N_5080,N_4377,N_4544);
and U5081 (N_5081,N_4179,N_4222);
nor U5082 (N_5082,N_4154,N_4523);
nor U5083 (N_5083,N_4253,N_4621);
nor U5084 (N_5084,N_4438,N_4630);
and U5085 (N_5085,N_4338,N_4178);
or U5086 (N_5086,N_4380,N_4615);
or U5087 (N_5087,N_4727,N_4314);
nor U5088 (N_5088,N_4056,N_4679);
and U5089 (N_5089,N_4240,N_4560);
and U5090 (N_5090,N_4086,N_4436);
nand U5091 (N_5091,N_4379,N_4634);
nand U5092 (N_5092,N_4713,N_4793);
nand U5093 (N_5093,N_4506,N_4425);
and U5094 (N_5094,N_4216,N_4307);
and U5095 (N_5095,N_4588,N_4769);
xor U5096 (N_5096,N_4682,N_4762);
and U5097 (N_5097,N_4312,N_4127);
nor U5098 (N_5098,N_4227,N_4720);
or U5099 (N_5099,N_4443,N_4141);
or U5100 (N_5100,N_4347,N_4476);
xnor U5101 (N_5101,N_4548,N_4073);
xor U5102 (N_5102,N_4002,N_4193);
or U5103 (N_5103,N_4656,N_4421);
nand U5104 (N_5104,N_4639,N_4335);
nor U5105 (N_5105,N_4041,N_4580);
nor U5106 (N_5106,N_4643,N_4101);
and U5107 (N_5107,N_4102,N_4349);
and U5108 (N_5108,N_4058,N_4747);
xnor U5109 (N_5109,N_4341,N_4414);
and U5110 (N_5110,N_4582,N_4782);
or U5111 (N_5111,N_4480,N_4319);
xor U5112 (N_5112,N_4491,N_4512);
nor U5113 (N_5113,N_4608,N_4322);
nand U5114 (N_5114,N_4042,N_4635);
nor U5115 (N_5115,N_4754,N_4751);
and U5116 (N_5116,N_4173,N_4390);
and U5117 (N_5117,N_4481,N_4774);
or U5118 (N_5118,N_4566,N_4693);
xor U5119 (N_5119,N_4357,N_4233);
and U5120 (N_5120,N_4108,N_4570);
or U5121 (N_5121,N_4358,N_4033);
xor U5122 (N_5122,N_4739,N_4559);
or U5123 (N_5123,N_4182,N_4485);
and U5124 (N_5124,N_4187,N_4107);
nor U5125 (N_5125,N_4045,N_4657);
nand U5126 (N_5126,N_4245,N_4034);
nor U5127 (N_5127,N_4003,N_4020);
and U5128 (N_5128,N_4525,N_4201);
nor U5129 (N_5129,N_4343,N_4124);
xnor U5130 (N_5130,N_4186,N_4708);
and U5131 (N_5131,N_4195,N_4665);
or U5132 (N_5132,N_4142,N_4675);
and U5133 (N_5133,N_4326,N_4299);
nor U5134 (N_5134,N_4297,N_4401);
nor U5135 (N_5135,N_4342,N_4407);
nor U5136 (N_5136,N_4166,N_4733);
nor U5137 (N_5137,N_4289,N_4432);
xnor U5138 (N_5138,N_4133,N_4531);
or U5139 (N_5139,N_4110,N_4484);
and U5140 (N_5140,N_4790,N_4515);
nand U5141 (N_5141,N_4792,N_4692);
nand U5142 (N_5142,N_4509,N_4786);
nand U5143 (N_5143,N_4383,N_4551);
xor U5144 (N_5144,N_4079,N_4169);
or U5145 (N_5145,N_4714,N_4255);
nand U5146 (N_5146,N_4537,N_4428);
nor U5147 (N_5147,N_4459,N_4772);
nand U5148 (N_5148,N_4168,N_4724);
nand U5149 (N_5149,N_4100,N_4009);
and U5150 (N_5150,N_4569,N_4249);
and U5151 (N_5151,N_4126,N_4492);
and U5152 (N_5152,N_4308,N_4658);
nor U5153 (N_5153,N_4507,N_4478);
and U5154 (N_5154,N_4505,N_4718);
and U5155 (N_5155,N_4422,N_4364);
nor U5156 (N_5156,N_4374,N_4153);
or U5157 (N_5157,N_4151,N_4155);
and U5158 (N_5158,N_4518,N_4389);
nand U5159 (N_5159,N_4103,N_4385);
nand U5160 (N_5160,N_4105,N_4771);
nor U5161 (N_5161,N_4680,N_4417);
or U5162 (N_5162,N_4598,N_4610);
nand U5163 (N_5163,N_4453,N_4647);
and U5164 (N_5164,N_4473,N_4435);
and U5165 (N_5165,N_4085,N_4496);
and U5166 (N_5166,N_4412,N_4025);
nand U5167 (N_5167,N_4770,N_4652);
nor U5168 (N_5168,N_4273,N_4044);
nor U5169 (N_5169,N_4328,N_4789);
and U5170 (N_5170,N_4640,N_4366);
xor U5171 (N_5171,N_4629,N_4547);
nand U5172 (N_5172,N_4371,N_4337);
nor U5173 (N_5173,N_4563,N_4454);
and U5174 (N_5174,N_4606,N_4022);
or U5175 (N_5175,N_4396,N_4067);
nand U5176 (N_5176,N_4498,N_4061);
and U5177 (N_5177,N_4265,N_4668);
and U5178 (N_5178,N_4355,N_4159);
and U5179 (N_5179,N_4167,N_4043);
xor U5180 (N_5180,N_4604,N_4584);
or U5181 (N_5181,N_4577,N_4750);
nand U5182 (N_5182,N_4471,N_4310);
nand U5183 (N_5183,N_4475,N_4504);
nor U5184 (N_5184,N_4611,N_4706);
xor U5185 (N_5185,N_4351,N_4689);
nor U5186 (N_5186,N_4522,N_4732);
or U5187 (N_5187,N_4325,N_4420);
nand U5188 (N_5188,N_4256,N_4464);
nand U5189 (N_5189,N_4646,N_4096);
and U5190 (N_5190,N_4758,N_4503);
xor U5191 (N_5191,N_4489,N_4644);
and U5192 (N_5192,N_4302,N_4290);
or U5193 (N_5193,N_4276,N_4098);
xnor U5194 (N_5194,N_4783,N_4788);
xor U5195 (N_5195,N_4541,N_4418);
nand U5196 (N_5196,N_4074,N_4023);
nor U5197 (N_5197,N_4458,N_4534);
nor U5198 (N_5198,N_4330,N_4303);
or U5199 (N_5199,N_4121,N_4521);
and U5200 (N_5200,N_4652,N_4324);
nor U5201 (N_5201,N_4389,N_4294);
nand U5202 (N_5202,N_4469,N_4775);
or U5203 (N_5203,N_4056,N_4223);
or U5204 (N_5204,N_4438,N_4524);
and U5205 (N_5205,N_4490,N_4393);
nand U5206 (N_5206,N_4625,N_4159);
nand U5207 (N_5207,N_4742,N_4640);
and U5208 (N_5208,N_4145,N_4577);
xnor U5209 (N_5209,N_4768,N_4374);
nand U5210 (N_5210,N_4108,N_4772);
or U5211 (N_5211,N_4723,N_4350);
nor U5212 (N_5212,N_4692,N_4003);
or U5213 (N_5213,N_4344,N_4625);
nor U5214 (N_5214,N_4215,N_4705);
nand U5215 (N_5215,N_4526,N_4789);
or U5216 (N_5216,N_4065,N_4283);
xnor U5217 (N_5217,N_4537,N_4522);
or U5218 (N_5218,N_4752,N_4581);
and U5219 (N_5219,N_4445,N_4527);
nand U5220 (N_5220,N_4667,N_4099);
and U5221 (N_5221,N_4411,N_4352);
nand U5222 (N_5222,N_4314,N_4231);
nor U5223 (N_5223,N_4788,N_4350);
xnor U5224 (N_5224,N_4173,N_4001);
and U5225 (N_5225,N_4073,N_4228);
nor U5226 (N_5226,N_4522,N_4388);
or U5227 (N_5227,N_4487,N_4328);
and U5228 (N_5228,N_4673,N_4079);
xor U5229 (N_5229,N_4135,N_4671);
or U5230 (N_5230,N_4149,N_4496);
or U5231 (N_5231,N_4520,N_4233);
or U5232 (N_5232,N_4726,N_4750);
and U5233 (N_5233,N_4765,N_4567);
and U5234 (N_5234,N_4166,N_4773);
nand U5235 (N_5235,N_4481,N_4105);
and U5236 (N_5236,N_4675,N_4421);
xnor U5237 (N_5237,N_4490,N_4161);
nor U5238 (N_5238,N_4688,N_4078);
xnor U5239 (N_5239,N_4671,N_4765);
and U5240 (N_5240,N_4089,N_4163);
or U5241 (N_5241,N_4568,N_4552);
nor U5242 (N_5242,N_4710,N_4351);
xnor U5243 (N_5243,N_4655,N_4003);
nor U5244 (N_5244,N_4387,N_4772);
or U5245 (N_5245,N_4251,N_4484);
or U5246 (N_5246,N_4043,N_4706);
or U5247 (N_5247,N_4448,N_4123);
and U5248 (N_5248,N_4476,N_4494);
nor U5249 (N_5249,N_4020,N_4764);
nor U5250 (N_5250,N_4078,N_4262);
nor U5251 (N_5251,N_4764,N_4571);
or U5252 (N_5252,N_4470,N_4122);
and U5253 (N_5253,N_4002,N_4684);
nor U5254 (N_5254,N_4219,N_4167);
nor U5255 (N_5255,N_4319,N_4372);
or U5256 (N_5256,N_4736,N_4512);
nor U5257 (N_5257,N_4146,N_4464);
nor U5258 (N_5258,N_4032,N_4698);
nor U5259 (N_5259,N_4427,N_4449);
or U5260 (N_5260,N_4731,N_4451);
or U5261 (N_5261,N_4761,N_4370);
and U5262 (N_5262,N_4656,N_4573);
or U5263 (N_5263,N_4377,N_4749);
or U5264 (N_5264,N_4535,N_4274);
and U5265 (N_5265,N_4034,N_4415);
xnor U5266 (N_5266,N_4269,N_4102);
xnor U5267 (N_5267,N_4058,N_4528);
or U5268 (N_5268,N_4566,N_4266);
and U5269 (N_5269,N_4451,N_4295);
nor U5270 (N_5270,N_4365,N_4449);
and U5271 (N_5271,N_4427,N_4378);
nor U5272 (N_5272,N_4768,N_4044);
xor U5273 (N_5273,N_4581,N_4379);
xnor U5274 (N_5274,N_4223,N_4386);
xnor U5275 (N_5275,N_4383,N_4187);
nor U5276 (N_5276,N_4187,N_4013);
xor U5277 (N_5277,N_4663,N_4684);
nor U5278 (N_5278,N_4428,N_4451);
nand U5279 (N_5279,N_4118,N_4026);
or U5280 (N_5280,N_4090,N_4543);
nor U5281 (N_5281,N_4697,N_4418);
xnor U5282 (N_5282,N_4109,N_4663);
or U5283 (N_5283,N_4137,N_4501);
or U5284 (N_5284,N_4528,N_4763);
and U5285 (N_5285,N_4204,N_4495);
nor U5286 (N_5286,N_4360,N_4279);
nor U5287 (N_5287,N_4767,N_4416);
nand U5288 (N_5288,N_4529,N_4620);
xnor U5289 (N_5289,N_4090,N_4031);
and U5290 (N_5290,N_4723,N_4662);
nor U5291 (N_5291,N_4002,N_4781);
nand U5292 (N_5292,N_4572,N_4161);
nand U5293 (N_5293,N_4540,N_4165);
nand U5294 (N_5294,N_4321,N_4738);
nand U5295 (N_5295,N_4417,N_4345);
and U5296 (N_5296,N_4206,N_4706);
and U5297 (N_5297,N_4322,N_4285);
and U5298 (N_5298,N_4705,N_4771);
xnor U5299 (N_5299,N_4658,N_4528);
or U5300 (N_5300,N_4121,N_4222);
nor U5301 (N_5301,N_4716,N_4410);
and U5302 (N_5302,N_4325,N_4470);
and U5303 (N_5303,N_4255,N_4125);
xor U5304 (N_5304,N_4336,N_4005);
and U5305 (N_5305,N_4535,N_4170);
or U5306 (N_5306,N_4287,N_4649);
or U5307 (N_5307,N_4713,N_4397);
nor U5308 (N_5308,N_4126,N_4146);
nor U5309 (N_5309,N_4744,N_4786);
xor U5310 (N_5310,N_4018,N_4593);
nor U5311 (N_5311,N_4022,N_4795);
and U5312 (N_5312,N_4075,N_4778);
nand U5313 (N_5313,N_4013,N_4404);
xor U5314 (N_5314,N_4632,N_4264);
or U5315 (N_5315,N_4538,N_4065);
or U5316 (N_5316,N_4454,N_4558);
and U5317 (N_5317,N_4324,N_4568);
xnor U5318 (N_5318,N_4738,N_4140);
or U5319 (N_5319,N_4247,N_4197);
and U5320 (N_5320,N_4350,N_4214);
or U5321 (N_5321,N_4491,N_4337);
nor U5322 (N_5322,N_4072,N_4147);
xnor U5323 (N_5323,N_4296,N_4310);
and U5324 (N_5324,N_4120,N_4332);
or U5325 (N_5325,N_4004,N_4539);
xnor U5326 (N_5326,N_4779,N_4097);
nand U5327 (N_5327,N_4159,N_4011);
or U5328 (N_5328,N_4237,N_4233);
xnor U5329 (N_5329,N_4475,N_4791);
nand U5330 (N_5330,N_4101,N_4551);
or U5331 (N_5331,N_4529,N_4083);
nor U5332 (N_5332,N_4780,N_4469);
xor U5333 (N_5333,N_4711,N_4181);
nor U5334 (N_5334,N_4712,N_4244);
and U5335 (N_5335,N_4108,N_4661);
and U5336 (N_5336,N_4765,N_4503);
xor U5337 (N_5337,N_4277,N_4084);
nor U5338 (N_5338,N_4639,N_4679);
nor U5339 (N_5339,N_4665,N_4548);
nand U5340 (N_5340,N_4774,N_4125);
nor U5341 (N_5341,N_4356,N_4209);
nand U5342 (N_5342,N_4305,N_4549);
xnor U5343 (N_5343,N_4010,N_4738);
nand U5344 (N_5344,N_4397,N_4581);
nor U5345 (N_5345,N_4478,N_4669);
xor U5346 (N_5346,N_4786,N_4356);
nor U5347 (N_5347,N_4783,N_4376);
xnor U5348 (N_5348,N_4607,N_4572);
nand U5349 (N_5349,N_4416,N_4544);
nor U5350 (N_5350,N_4364,N_4160);
and U5351 (N_5351,N_4785,N_4532);
nand U5352 (N_5352,N_4317,N_4073);
nor U5353 (N_5353,N_4126,N_4369);
nand U5354 (N_5354,N_4441,N_4471);
or U5355 (N_5355,N_4016,N_4557);
or U5356 (N_5356,N_4146,N_4767);
and U5357 (N_5357,N_4564,N_4062);
nor U5358 (N_5358,N_4583,N_4768);
and U5359 (N_5359,N_4287,N_4028);
xnor U5360 (N_5360,N_4678,N_4351);
nor U5361 (N_5361,N_4354,N_4555);
xnor U5362 (N_5362,N_4694,N_4617);
xor U5363 (N_5363,N_4262,N_4216);
nor U5364 (N_5364,N_4123,N_4110);
or U5365 (N_5365,N_4036,N_4399);
and U5366 (N_5366,N_4169,N_4470);
xnor U5367 (N_5367,N_4193,N_4060);
nand U5368 (N_5368,N_4753,N_4484);
or U5369 (N_5369,N_4454,N_4004);
xnor U5370 (N_5370,N_4673,N_4110);
nor U5371 (N_5371,N_4636,N_4137);
nand U5372 (N_5372,N_4722,N_4176);
nand U5373 (N_5373,N_4433,N_4508);
and U5374 (N_5374,N_4314,N_4638);
nand U5375 (N_5375,N_4121,N_4291);
or U5376 (N_5376,N_4407,N_4237);
xnor U5377 (N_5377,N_4420,N_4659);
nor U5378 (N_5378,N_4563,N_4184);
xor U5379 (N_5379,N_4395,N_4220);
and U5380 (N_5380,N_4341,N_4151);
and U5381 (N_5381,N_4366,N_4484);
xnor U5382 (N_5382,N_4664,N_4287);
or U5383 (N_5383,N_4052,N_4585);
xor U5384 (N_5384,N_4188,N_4743);
nand U5385 (N_5385,N_4703,N_4536);
nand U5386 (N_5386,N_4144,N_4681);
nor U5387 (N_5387,N_4715,N_4168);
nor U5388 (N_5388,N_4774,N_4384);
nand U5389 (N_5389,N_4727,N_4449);
xnor U5390 (N_5390,N_4207,N_4116);
and U5391 (N_5391,N_4595,N_4457);
or U5392 (N_5392,N_4646,N_4584);
nor U5393 (N_5393,N_4257,N_4753);
xor U5394 (N_5394,N_4576,N_4407);
and U5395 (N_5395,N_4470,N_4601);
nand U5396 (N_5396,N_4584,N_4259);
nor U5397 (N_5397,N_4391,N_4050);
nor U5398 (N_5398,N_4288,N_4536);
nand U5399 (N_5399,N_4118,N_4193);
and U5400 (N_5400,N_4144,N_4538);
or U5401 (N_5401,N_4043,N_4466);
xor U5402 (N_5402,N_4742,N_4171);
nor U5403 (N_5403,N_4472,N_4289);
or U5404 (N_5404,N_4127,N_4151);
or U5405 (N_5405,N_4245,N_4134);
nand U5406 (N_5406,N_4756,N_4774);
and U5407 (N_5407,N_4522,N_4172);
and U5408 (N_5408,N_4588,N_4633);
xnor U5409 (N_5409,N_4291,N_4450);
or U5410 (N_5410,N_4606,N_4062);
nor U5411 (N_5411,N_4004,N_4011);
and U5412 (N_5412,N_4531,N_4370);
nor U5413 (N_5413,N_4101,N_4277);
nand U5414 (N_5414,N_4437,N_4636);
and U5415 (N_5415,N_4669,N_4284);
nor U5416 (N_5416,N_4612,N_4274);
nor U5417 (N_5417,N_4523,N_4242);
xnor U5418 (N_5418,N_4305,N_4345);
xnor U5419 (N_5419,N_4468,N_4531);
xor U5420 (N_5420,N_4616,N_4060);
xor U5421 (N_5421,N_4294,N_4480);
xnor U5422 (N_5422,N_4250,N_4474);
nor U5423 (N_5423,N_4074,N_4487);
and U5424 (N_5424,N_4767,N_4539);
or U5425 (N_5425,N_4440,N_4133);
nand U5426 (N_5426,N_4625,N_4507);
nor U5427 (N_5427,N_4687,N_4621);
and U5428 (N_5428,N_4395,N_4541);
nand U5429 (N_5429,N_4019,N_4584);
or U5430 (N_5430,N_4427,N_4769);
xor U5431 (N_5431,N_4131,N_4001);
or U5432 (N_5432,N_4513,N_4734);
nor U5433 (N_5433,N_4592,N_4070);
nor U5434 (N_5434,N_4585,N_4798);
or U5435 (N_5435,N_4641,N_4215);
xor U5436 (N_5436,N_4720,N_4405);
nand U5437 (N_5437,N_4382,N_4170);
and U5438 (N_5438,N_4647,N_4281);
and U5439 (N_5439,N_4430,N_4074);
xor U5440 (N_5440,N_4488,N_4154);
nand U5441 (N_5441,N_4597,N_4216);
nand U5442 (N_5442,N_4660,N_4298);
nand U5443 (N_5443,N_4311,N_4490);
and U5444 (N_5444,N_4726,N_4267);
xnor U5445 (N_5445,N_4250,N_4366);
nor U5446 (N_5446,N_4298,N_4229);
nand U5447 (N_5447,N_4732,N_4319);
or U5448 (N_5448,N_4087,N_4478);
and U5449 (N_5449,N_4685,N_4327);
or U5450 (N_5450,N_4025,N_4045);
or U5451 (N_5451,N_4106,N_4276);
nand U5452 (N_5452,N_4432,N_4478);
xor U5453 (N_5453,N_4347,N_4504);
or U5454 (N_5454,N_4271,N_4291);
or U5455 (N_5455,N_4455,N_4243);
and U5456 (N_5456,N_4565,N_4299);
xnor U5457 (N_5457,N_4636,N_4757);
xnor U5458 (N_5458,N_4588,N_4081);
nand U5459 (N_5459,N_4651,N_4159);
nand U5460 (N_5460,N_4546,N_4286);
or U5461 (N_5461,N_4067,N_4268);
xnor U5462 (N_5462,N_4344,N_4769);
xnor U5463 (N_5463,N_4479,N_4101);
or U5464 (N_5464,N_4774,N_4361);
or U5465 (N_5465,N_4240,N_4259);
and U5466 (N_5466,N_4234,N_4017);
and U5467 (N_5467,N_4562,N_4092);
and U5468 (N_5468,N_4009,N_4260);
xor U5469 (N_5469,N_4206,N_4173);
or U5470 (N_5470,N_4629,N_4319);
and U5471 (N_5471,N_4601,N_4049);
nor U5472 (N_5472,N_4491,N_4661);
nand U5473 (N_5473,N_4460,N_4746);
nor U5474 (N_5474,N_4528,N_4420);
or U5475 (N_5475,N_4794,N_4617);
nand U5476 (N_5476,N_4032,N_4196);
nand U5477 (N_5477,N_4148,N_4062);
and U5478 (N_5478,N_4358,N_4767);
nor U5479 (N_5479,N_4184,N_4331);
and U5480 (N_5480,N_4736,N_4644);
xnor U5481 (N_5481,N_4323,N_4495);
nand U5482 (N_5482,N_4217,N_4278);
or U5483 (N_5483,N_4725,N_4194);
or U5484 (N_5484,N_4435,N_4316);
nor U5485 (N_5485,N_4440,N_4273);
nand U5486 (N_5486,N_4078,N_4621);
or U5487 (N_5487,N_4211,N_4299);
nor U5488 (N_5488,N_4783,N_4392);
nand U5489 (N_5489,N_4474,N_4709);
nor U5490 (N_5490,N_4469,N_4120);
and U5491 (N_5491,N_4779,N_4548);
or U5492 (N_5492,N_4204,N_4265);
or U5493 (N_5493,N_4272,N_4361);
and U5494 (N_5494,N_4512,N_4797);
xnor U5495 (N_5495,N_4087,N_4417);
nor U5496 (N_5496,N_4759,N_4595);
or U5497 (N_5497,N_4514,N_4469);
and U5498 (N_5498,N_4741,N_4630);
and U5499 (N_5499,N_4094,N_4080);
nor U5500 (N_5500,N_4309,N_4247);
nand U5501 (N_5501,N_4626,N_4706);
nand U5502 (N_5502,N_4141,N_4796);
nand U5503 (N_5503,N_4609,N_4203);
xor U5504 (N_5504,N_4298,N_4647);
xor U5505 (N_5505,N_4421,N_4699);
xor U5506 (N_5506,N_4270,N_4310);
nand U5507 (N_5507,N_4406,N_4418);
or U5508 (N_5508,N_4027,N_4534);
nor U5509 (N_5509,N_4363,N_4175);
nand U5510 (N_5510,N_4140,N_4676);
xor U5511 (N_5511,N_4187,N_4393);
nor U5512 (N_5512,N_4417,N_4071);
nand U5513 (N_5513,N_4322,N_4049);
and U5514 (N_5514,N_4023,N_4163);
nor U5515 (N_5515,N_4242,N_4050);
or U5516 (N_5516,N_4470,N_4771);
nor U5517 (N_5517,N_4455,N_4323);
xnor U5518 (N_5518,N_4160,N_4125);
xnor U5519 (N_5519,N_4386,N_4687);
or U5520 (N_5520,N_4128,N_4052);
and U5521 (N_5521,N_4447,N_4557);
xnor U5522 (N_5522,N_4707,N_4069);
or U5523 (N_5523,N_4098,N_4465);
and U5524 (N_5524,N_4176,N_4749);
and U5525 (N_5525,N_4550,N_4072);
xnor U5526 (N_5526,N_4129,N_4010);
xnor U5527 (N_5527,N_4472,N_4109);
nand U5528 (N_5528,N_4502,N_4571);
and U5529 (N_5529,N_4536,N_4046);
or U5530 (N_5530,N_4257,N_4078);
or U5531 (N_5531,N_4705,N_4356);
nor U5532 (N_5532,N_4635,N_4085);
or U5533 (N_5533,N_4449,N_4546);
nor U5534 (N_5534,N_4037,N_4315);
nand U5535 (N_5535,N_4613,N_4653);
xor U5536 (N_5536,N_4121,N_4586);
nor U5537 (N_5537,N_4710,N_4745);
xnor U5538 (N_5538,N_4393,N_4687);
nand U5539 (N_5539,N_4233,N_4470);
and U5540 (N_5540,N_4218,N_4580);
nand U5541 (N_5541,N_4623,N_4123);
nand U5542 (N_5542,N_4215,N_4522);
xnor U5543 (N_5543,N_4501,N_4008);
xor U5544 (N_5544,N_4637,N_4390);
nor U5545 (N_5545,N_4025,N_4426);
and U5546 (N_5546,N_4691,N_4404);
or U5547 (N_5547,N_4113,N_4799);
xor U5548 (N_5548,N_4594,N_4627);
or U5549 (N_5549,N_4744,N_4158);
or U5550 (N_5550,N_4143,N_4565);
and U5551 (N_5551,N_4727,N_4632);
and U5552 (N_5552,N_4658,N_4736);
nor U5553 (N_5553,N_4716,N_4074);
nor U5554 (N_5554,N_4639,N_4604);
nand U5555 (N_5555,N_4019,N_4497);
or U5556 (N_5556,N_4237,N_4746);
nor U5557 (N_5557,N_4253,N_4521);
xnor U5558 (N_5558,N_4790,N_4213);
nand U5559 (N_5559,N_4635,N_4669);
nor U5560 (N_5560,N_4595,N_4477);
and U5561 (N_5561,N_4685,N_4315);
and U5562 (N_5562,N_4265,N_4739);
or U5563 (N_5563,N_4719,N_4029);
xnor U5564 (N_5564,N_4726,N_4334);
or U5565 (N_5565,N_4619,N_4439);
xor U5566 (N_5566,N_4120,N_4371);
xor U5567 (N_5567,N_4286,N_4346);
or U5568 (N_5568,N_4185,N_4698);
or U5569 (N_5569,N_4430,N_4280);
and U5570 (N_5570,N_4480,N_4783);
nor U5571 (N_5571,N_4711,N_4024);
or U5572 (N_5572,N_4119,N_4144);
or U5573 (N_5573,N_4117,N_4195);
or U5574 (N_5574,N_4611,N_4192);
xor U5575 (N_5575,N_4611,N_4080);
or U5576 (N_5576,N_4691,N_4796);
or U5577 (N_5577,N_4595,N_4713);
nand U5578 (N_5578,N_4124,N_4006);
and U5579 (N_5579,N_4292,N_4343);
or U5580 (N_5580,N_4275,N_4308);
or U5581 (N_5581,N_4391,N_4587);
xor U5582 (N_5582,N_4017,N_4300);
nand U5583 (N_5583,N_4776,N_4757);
xnor U5584 (N_5584,N_4259,N_4683);
nor U5585 (N_5585,N_4748,N_4613);
or U5586 (N_5586,N_4558,N_4646);
xnor U5587 (N_5587,N_4673,N_4603);
nand U5588 (N_5588,N_4726,N_4624);
or U5589 (N_5589,N_4470,N_4440);
nor U5590 (N_5590,N_4666,N_4250);
or U5591 (N_5591,N_4732,N_4305);
and U5592 (N_5592,N_4131,N_4694);
nor U5593 (N_5593,N_4273,N_4177);
nor U5594 (N_5594,N_4081,N_4110);
or U5595 (N_5595,N_4712,N_4475);
nor U5596 (N_5596,N_4549,N_4642);
xnor U5597 (N_5597,N_4069,N_4574);
xor U5598 (N_5598,N_4726,N_4082);
and U5599 (N_5599,N_4714,N_4565);
nand U5600 (N_5600,N_5172,N_4932);
or U5601 (N_5601,N_5484,N_5081);
nand U5602 (N_5602,N_5076,N_5097);
nor U5603 (N_5603,N_5471,N_4868);
nor U5604 (N_5604,N_5210,N_4820);
or U5605 (N_5605,N_4927,N_4884);
or U5606 (N_5606,N_4917,N_5103);
nor U5607 (N_5607,N_5045,N_4822);
and U5608 (N_5608,N_5021,N_5307);
xnor U5609 (N_5609,N_5430,N_5215);
nor U5610 (N_5610,N_5478,N_5351);
xnor U5611 (N_5611,N_5000,N_5056);
nor U5612 (N_5612,N_5014,N_5335);
nand U5613 (N_5613,N_5320,N_5567);
or U5614 (N_5614,N_4890,N_5362);
xor U5615 (N_5615,N_4894,N_5548);
or U5616 (N_5616,N_4818,N_4805);
and U5617 (N_5617,N_4980,N_5541);
nor U5618 (N_5618,N_5383,N_5507);
nor U5619 (N_5619,N_4965,N_5490);
nand U5620 (N_5620,N_5206,N_4913);
and U5621 (N_5621,N_4836,N_5575);
xor U5622 (N_5622,N_4975,N_4977);
nor U5623 (N_5623,N_4887,N_4986);
xor U5624 (N_5624,N_5528,N_5192);
nand U5625 (N_5625,N_5273,N_4909);
nor U5626 (N_5626,N_4883,N_5209);
and U5627 (N_5627,N_4892,N_5463);
nor U5628 (N_5628,N_5572,N_4831);
nand U5629 (N_5629,N_5070,N_4929);
nand U5630 (N_5630,N_5593,N_5553);
and U5631 (N_5631,N_5361,N_5183);
and U5632 (N_5632,N_5074,N_4912);
xor U5633 (N_5633,N_5433,N_4924);
or U5634 (N_5634,N_5296,N_5378);
nor U5635 (N_5635,N_5105,N_5440);
xor U5636 (N_5636,N_4861,N_5050);
or U5637 (N_5637,N_5256,N_5517);
or U5638 (N_5638,N_4900,N_4899);
xor U5639 (N_5639,N_5522,N_5554);
or U5640 (N_5640,N_4910,N_5495);
nand U5641 (N_5641,N_4840,N_5476);
or U5642 (N_5642,N_5055,N_5002);
nand U5643 (N_5643,N_5315,N_5505);
and U5644 (N_5644,N_5282,N_5068);
xnor U5645 (N_5645,N_5565,N_5322);
nor U5646 (N_5646,N_5480,N_5020);
or U5647 (N_5647,N_5143,N_5584);
nor U5648 (N_5648,N_4863,N_5061);
xnor U5649 (N_5649,N_4806,N_5201);
and U5650 (N_5650,N_4835,N_5487);
and U5651 (N_5651,N_5087,N_5562);
xnor U5652 (N_5652,N_5396,N_5039);
nor U5653 (N_5653,N_5308,N_5346);
nor U5654 (N_5654,N_4915,N_4922);
or U5655 (N_5655,N_5400,N_5560);
and U5656 (N_5656,N_5537,N_5017);
or U5657 (N_5657,N_5341,N_5489);
and U5658 (N_5658,N_5437,N_4838);
or U5659 (N_5659,N_4946,N_5113);
xor U5660 (N_5660,N_5016,N_5295);
or U5661 (N_5661,N_5167,N_5262);
nor U5662 (N_5662,N_4962,N_5218);
nor U5663 (N_5663,N_5424,N_5263);
and U5664 (N_5664,N_5175,N_5112);
nor U5665 (N_5665,N_5136,N_5510);
xnor U5666 (N_5666,N_5391,N_5024);
xor U5667 (N_5667,N_5547,N_5202);
nor U5668 (N_5668,N_4904,N_5423);
nand U5669 (N_5669,N_5312,N_5379);
xor U5670 (N_5670,N_5096,N_5003);
nand U5671 (N_5671,N_5043,N_4878);
and U5672 (N_5672,N_5271,N_5501);
nor U5673 (N_5673,N_5591,N_4874);
or U5674 (N_5674,N_5008,N_4813);
nor U5675 (N_5675,N_5121,N_5082);
nand U5676 (N_5676,N_5534,N_5417);
and U5677 (N_5677,N_5023,N_5291);
or U5678 (N_5678,N_4939,N_5149);
or U5679 (N_5679,N_5561,N_4814);
and U5680 (N_5680,N_5040,N_4837);
nor U5681 (N_5681,N_5098,N_5460);
and U5682 (N_5682,N_5375,N_5146);
or U5683 (N_5683,N_4829,N_5544);
xor U5684 (N_5684,N_5456,N_5369);
nor U5685 (N_5685,N_5037,N_5052);
xnor U5686 (N_5686,N_5334,N_5289);
nor U5687 (N_5687,N_5197,N_5216);
nand U5688 (N_5688,N_5154,N_4921);
xnor U5689 (N_5689,N_5367,N_5111);
xor U5690 (N_5690,N_5598,N_5166);
xnor U5691 (N_5691,N_5570,N_5464);
xnor U5692 (N_5692,N_5515,N_5571);
xnor U5693 (N_5693,N_5481,N_5107);
or U5694 (N_5694,N_5427,N_5546);
nor U5695 (N_5695,N_5477,N_5277);
and U5696 (N_5696,N_4888,N_5304);
or U5697 (N_5697,N_4864,N_5414);
nor U5698 (N_5698,N_4817,N_5110);
nor U5699 (N_5699,N_5599,N_4844);
nor U5700 (N_5700,N_5494,N_5445);
xnor U5701 (N_5701,N_5004,N_5190);
or U5702 (N_5702,N_5413,N_4841);
nand U5703 (N_5703,N_4935,N_4846);
xnor U5704 (N_5704,N_5473,N_5550);
xnor U5705 (N_5705,N_5497,N_4978);
nand U5706 (N_5706,N_5314,N_5503);
and U5707 (N_5707,N_5182,N_5191);
or U5708 (N_5708,N_4880,N_4807);
nand U5709 (N_5709,N_5582,N_5421);
or U5710 (N_5710,N_4891,N_5313);
xnor U5711 (N_5711,N_5329,N_4976);
nor U5712 (N_5712,N_5186,N_5453);
nor U5713 (N_5713,N_5179,N_5587);
nand U5714 (N_5714,N_5441,N_4827);
nor U5715 (N_5715,N_5422,N_5029);
xnor U5716 (N_5716,N_5504,N_5472);
nand U5717 (N_5717,N_5022,N_5316);
and U5718 (N_5718,N_5249,N_5298);
xnor U5719 (N_5719,N_5145,N_4923);
or U5720 (N_5720,N_4987,N_4948);
and U5721 (N_5721,N_5005,N_5426);
xor U5722 (N_5722,N_5493,N_5224);
nor U5723 (N_5723,N_5347,N_5200);
and U5724 (N_5724,N_5164,N_5062);
xor U5725 (N_5725,N_5144,N_5574);
or U5726 (N_5726,N_5229,N_5042);
or U5727 (N_5727,N_5397,N_5538);
nor U5728 (N_5728,N_5011,N_5213);
nor U5729 (N_5729,N_5482,N_5344);
nor U5730 (N_5730,N_5302,N_4854);
or U5731 (N_5731,N_5088,N_5261);
or U5732 (N_5732,N_5454,N_4843);
or U5733 (N_5733,N_5306,N_4947);
nand U5734 (N_5734,N_5118,N_4958);
or U5735 (N_5735,N_5108,N_5284);
nand U5736 (N_5736,N_5390,N_4898);
or U5737 (N_5737,N_5169,N_5188);
or U5738 (N_5738,N_5001,N_5125);
nor U5739 (N_5739,N_5048,N_5388);
xor U5740 (N_5740,N_5009,N_5447);
nand U5741 (N_5741,N_5467,N_5293);
or U5742 (N_5742,N_4984,N_5138);
xnor U5743 (N_5743,N_5533,N_5139);
xnor U5744 (N_5744,N_4824,N_4937);
and U5745 (N_5745,N_5208,N_5207);
or U5746 (N_5746,N_5134,N_5151);
and U5747 (N_5747,N_5231,N_5535);
nor U5748 (N_5748,N_4972,N_5475);
nor U5749 (N_5749,N_5323,N_5095);
and U5750 (N_5750,N_5279,N_5147);
xnor U5751 (N_5751,N_5398,N_4979);
and U5752 (N_5752,N_5246,N_5349);
nor U5753 (N_5753,N_4832,N_5058);
nand U5754 (N_5754,N_4943,N_5434);
nor U5755 (N_5755,N_5506,N_5583);
and U5756 (N_5756,N_4901,N_4886);
nand U5757 (N_5757,N_5485,N_4810);
or U5758 (N_5758,N_5496,N_5157);
or U5759 (N_5759,N_5597,N_5133);
or U5760 (N_5760,N_5558,N_5180);
and U5761 (N_5761,N_4959,N_5331);
and U5762 (N_5762,N_5371,N_5025);
nor U5763 (N_5763,N_4897,N_4803);
nand U5764 (N_5764,N_5049,N_4875);
or U5765 (N_5765,N_5556,N_5270);
nor U5766 (N_5766,N_5226,N_4999);
or U5767 (N_5767,N_5405,N_4881);
or U5768 (N_5768,N_5559,N_5457);
xnor U5769 (N_5769,N_5163,N_5126);
nor U5770 (N_5770,N_5243,N_4916);
xnor U5771 (N_5771,N_4925,N_5168);
xor U5772 (N_5772,N_5115,N_5019);
or U5773 (N_5773,N_5268,N_5137);
nor U5774 (N_5774,N_5358,N_5174);
nor U5775 (N_5775,N_4860,N_5079);
nand U5776 (N_5776,N_5227,N_5235);
nor U5777 (N_5777,N_4938,N_5403);
xor U5778 (N_5778,N_5013,N_5170);
nor U5779 (N_5779,N_5581,N_5381);
and U5780 (N_5780,N_5211,N_4982);
and U5781 (N_5781,N_5193,N_5511);
or U5782 (N_5782,N_5248,N_5435);
and U5783 (N_5783,N_5324,N_5205);
nor U5784 (N_5784,N_5491,N_5438);
or U5785 (N_5785,N_5552,N_5366);
and U5786 (N_5786,N_5116,N_4801);
xor U5787 (N_5787,N_4828,N_5060);
and U5788 (N_5788,N_5189,N_5408);
xnor U5789 (N_5789,N_4834,N_5418);
xor U5790 (N_5790,N_5303,N_5589);
nor U5791 (N_5791,N_5094,N_5032);
nand U5792 (N_5792,N_5236,N_5247);
nand U5793 (N_5793,N_4816,N_5339);
nand U5794 (N_5794,N_4882,N_4981);
or U5795 (N_5795,N_4992,N_5327);
and U5796 (N_5796,N_4988,N_5161);
nor U5797 (N_5797,N_4934,N_5519);
or U5798 (N_5798,N_5269,N_5594);
nor U5799 (N_5799,N_4808,N_5450);
and U5800 (N_5800,N_5075,N_5353);
nand U5801 (N_5801,N_5513,N_5091);
nand U5802 (N_5802,N_4954,N_4871);
nand U5803 (N_5803,N_5204,N_5444);
xor U5804 (N_5804,N_5350,N_5382);
nor U5805 (N_5805,N_5374,N_5276);
xnor U5806 (N_5806,N_5252,N_5240);
or U5807 (N_5807,N_4905,N_5089);
or U5808 (N_5808,N_5027,N_5330);
xnor U5809 (N_5809,N_4953,N_5041);
or U5810 (N_5810,N_5077,N_5274);
nor U5811 (N_5811,N_5580,N_5128);
and U5812 (N_5812,N_5549,N_5285);
and U5813 (N_5813,N_5203,N_5159);
nor U5814 (N_5814,N_5365,N_5498);
or U5815 (N_5815,N_5177,N_5523);
nand U5816 (N_5816,N_5458,N_5539);
nor U5817 (N_5817,N_5419,N_4815);
and U5818 (N_5818,N_5232,N_5286);
and U5819 (N_5819,N_5486,N_5195);
or U5820 (N_5820,N_5474,N_4936);
nand U5821 (N_5821,N_5508,N_5305);
nand U5822 (N_5822,N_5321,N_5266);
and U5823 (N_5823,N_5411,N_5573);
nand U5824 (N_5824,N_5187,N_4819);
and U5825 (N_5825,N_4858,N_5173);
or U5826 (N_5826,N_5083,N_5328);
nor U5827 (N_5827,N_5030,N_5569);
xor U5828 (N_5828,N_5406,N_5563);
xor U5829 (N_5829,N_5380,N_4974);
or U5830 (N_5830,N_5104,N_4902);
xor U5831 (N_5831,N_5551,N_4941);
xor U5832 (N_5832,N_4914,N_5439);
or U5833 (N_5833,N_5527,N_5124);
xnor U5834 (N_5834,N_5036,N_5067);
and U5835 (N_5835,N_5254,N_4918);
and U5836 (N_5836,N_5443,N_4847);
xnor U5837 (N_5837,N_4809,N_5337);
and U5838 (N_5838,N_5373,N_5386);
nor U5839 (N_5839,N_5360,N_5586);
xnor U5840 (N_5840,N_5160,N_5199);
and U5841 (N_5841,N_5150,N_5499);
or U5842 (N_5842,N_5526,N_5198);
nand U5843 (N_5843,N_5233,N_5123);
nand U5844 (N_5844,N_5018,N_5120);
nor U5845 (N_5845,N_5420,N_5015);
nor U5846 (N_5846,N_5148,N_4867);
nor U5847 (N_5847,N_5010,N_5465);
and U5848 (N_5848,N_5214,N_5415);
nor U5849 (N_5849,N_5448,N_5340);
or U5850 (N_5850,N_5102,N_4998);
and U5851 (N_5851,N_5162,N_5479);
and U5852 (N_5852,N_5222,N_4931);
nor U5853 (N_5853,N_4973,N_5370);
and U5854 (N_5854,N_4862,N_5272);
nand U5855 (N_5855,N_4848,N_4963);
xnor U5856 (N_5856,N_5238,N_4990);
nor U5857 (N_5857,N_5318,N_5090);
and U5858 (N_5858,N_5542,N_4957);
and U5859 (N_5859,N_4876,N_5033);
nand U5860 (N_5860,N_5514,N_4949);
nor U5861 (N_5861,N_5431,N_5114);
and U5862 (N_5862,N_5509,N_5127);
xnor U5863 (N_5863,N_5557,N_5117);
or U5864 (N_5864,N_5051,N_5100);
nor U5865 (N_5865,N_4996,N_5387);
and U5866 (N_5866,N_5566,N_4997);
or U5867 (N_5867,N_5185,N_5228);
nor U5868 (N_5868,N_4933,N_5086);
nand U5869 (N_5869,N_4991,N_4951);
xor U5870 (N_5870,N_4865,N_4889);
nor U5871 (N_5871,N_4839,N_4993);
nand U5872 (N_5872,N_5244,N_4872);
xor U5873 (N_5873,N_5392,N_5536);
xnor U5874 (N_5874,N_5326,N_5155);
and U5875 (N_5875,N_5348,N_5336);
xor U5876 (N_5876,N_5064,N_4989);
xnor U5877 (N_5877,N_5035,N_5462);
and U5878 (N_5878,N_5278,N_5059);
nand U5879 (N_5879,N_5389,N_5038);
and U5880 (N_5880,N_5342,N_5455);
nand U5881 (N_5881,N_4920,N_5409);
or U5882 (N_5882,N_5156,N_5141);
or U5883 (N_5883,N_5310,N_5596);
and U5884 (N_5884,N_5122,N_5069);
xnor U5885 (N_5885,N_5309,N_5543);
or U5886 (N_5886,N_5555,N_4955);
nor U5887 (N_5887,N_4812,N_4850);
xnor U5888 (N_5888,N_5301,N_4950);
xnor U5889 (N_5889,N_5354,N_4930);
xor U5890 (N_5890,N_5007,N_5132);
nor U5891 (N_5891,N_5364,N_5545);
nor U5892 (N_5892,N_4800,N_5130);
xor U5893 (N_5893,N_5153,N_5220);
and U5894 (N_5894,N_4908,N_5449);
xor U5895 (N_5895,N_4940,N_5294);
xnor U5896 (N_5896,N_5300,N_5525);
and U5897 (N_5897,N_5401,N_5026);
nand U5898 (N_5898,N_5099,N_5585);
or U5899 (N_5899,N_5520,N_5385);
xor U5900 (N_5900,N_5084,N_4994);
or U5901 (N_5901,N_5568,N_4903);
and U5902 (N_5902,N_5540,N_4842);
nor U5903 (N_5903,N_4960,N_4964);
and U5904 (N_5904,N_5578,N_5028);
and U5905 (N_5905,N_4896,N_5080);
nand U5906 (N_5906,N_5425,N_4873);
xor U5907 (N_5907,N_5230,N_5595);
and U5908 (N_5908,N_5258,N_5343);
and U5909 (N_5909,N_5085,N_5265);
xnor U5910 (N_5910,N_5178,N_5135);
or U5911 (N_5911,N_5529,N_5412);
or U5912 (N_5912,N_4845,N_5524);
or U5913 (N_5913,N_5044,N_5093);
or U5914 (N_5914,N_5280,N_4945);
xnor U5915 (N_5915,N_4804,N_5404);
and U5916 (N_5916,N_5241,N_4966);
nand U5917 (N_5917,N_5181,N_5532);
or U5918 (N_5918,N_5101,N_5275);
and U5919 (N_5919,N_5576,N_5319);
nor U5920 (N_5920,N_4944,N_4859);
nor U5921 (N_5921,N_5176,N_5292);
xor U5922 (N_5922,N_4855,N_5054);
nor U5923 (N_5923,N_5407,N_4969);
nand U5924 (N_5924,N_4866,N_5359);
or U5925 (N_5925,N_4895,N_5264);
xor U5926 (N_5926,N_5259,N_5432);
xnor U5927 (N_5927,N_5394,N_5171);
nand U5928 (N_5928,N_5217,N_5399);
nor U5929 (N_5929,N_4919,N_5516);
xor U5930 (N_5930,N_5325,N_4926);
xnor U5931 (N_5931,N_5512,N_5046);
nand U5932 (N_5932,N_5590,N_5466);
nand U5933 (N_5933,N_5564,N_5281);
or U5934 (N_5934,N_5253,N_5531);
nor U5935 (N_5935,N_5006,N_5131);
nor U5936 (N_5936,N_5129,N_4928);
or U5937 (N_5937,N_5299,N_4885);
nor U5938 (N_5938,N_5521,N_5384);
nand U5939 (N_5939,N_5442,N_5451);
nor U5940 (N_5940,N_5357,N_4967);
nand U5941 (N_5941,N_5311,N_4830);
and U5942 (N_5942,N_5250,N_5245);
nand U5943 (N_5943,N_4911,N_5047);
nand U5944 (N_5944,N_5352,N_5372);
nand U5945 (N_5945,N_5395,N_5219);
or U5946 (N_5946,N_5446,N_5355);
or U5947 (N_5947,N_4851,N_5066);
nand U5948 (N_5948,N_5065,N_5452);
nor U5949 (N_5949,N_4952,N_5518);
xnor U5950 (N_5950,N_5488,N_5345);
and U5951 (N_5951,N_5470,N_5410);
and U5952 (N_5952,N_4942,N_4985);
nor U5953 (N_5953,N_5225,N_4956);
and U5954 (N_5954,N_4971,N_4856);
nor U5955 (N_5955,N_4857,N_4825);
and U5956 (N_5956,N_5500,N_5221);
and U5957 (N_5957,N_5436,N_5333);
nand U5958 (N_5958,N_4983,N_5459);
nor U5959 (N_5959,N_5368,N_4970);
xor U5960 (N_5960,N_5158,N_5165);
and U5961 (N_5961,N_4853,N_5092);
and U5962 (N_5962,N_5251,N_5063);
or U5963 (N_5963,N_5212,N_4893);
and U5964 (N_5964,N_5469,N_5338);
xor U5965 (N_5965,N_5071,N_5577);
nand U5966 (N_5966,N_5530,N_5332);
nor U5967 (N_5967,N_5242,N_4852);
nor U5968 (N_5968,N_5492,N_4823);
xor U5969 (N_5969,N_4879,N_5356);
xnor U5970 (N_5970,N_4821,N_5237);
nand U5971 (N_5971,N_5290,N_5428);
or U5972 (N_5972,N_5078,N_5072);
xor U5973 (N_5973,N_5053,N_5588);
or U5974 (N_5974,N_4907,N_4869);
or U5975 (N_5975,N_5106,N_4833);
and U5976 (N_5976,N_5239,N_4877);
nand U5977 (N_5977,N_5287,N_5109);
nor U5978 (N_5978,N_5152,N_5592);
nand U5979 (N_5979,N_5255,N_5283);
or U5980 (N_5980,N_5057,N_5073);
nor U5981 (N_5981,N_5140,N_5142);
xor U5982 (N_5982,N_5502,N_5234);
and U5983 (N_5983,N_5376,N_5260);
nand U5984 (N_5984,N_5184,N_5579);
nor U5985 (N_5985,N_4802,N_5288);
nand U5986 (N_5986,N_5012,N_5119);
or U5987 (N_5987,N_5377,N_5393);
and U5988 (N_5988,N_5267,N_4961);
or U5989 (N_5989,N_4811,N_5416);
nand U5990 (N_5990,N_4995,N_5034);
or U5991 (N_5991,N_5223,N_4968);
nor U5992 (N_5992,N_5031,N_4849);
and U5993 (N_5993,N_4870,N_5194);
xnor U5994 (N_5994,N_5483,N_5468);
nand U5995 (N_5995,N_5297,N_5429);
and U5996 (N_5996,N_5196,N_5402);
and U5997 (N_5997,N_5363,N_5257);
nor U5998 (N_5998,N_4826,N_5317);
and U5999 (N_5999,N_5461,N_4906);
nand U6000 (N_6000,N_5113,N_5331);
nand U6001 (N_6001,N_4966,N_4969);
or U6002 (N_6002,N_5160,N_5202);
nand U6003 (N_6003,N_5102,N_5154);
xor U6004 (N_6004,N_5051,N_5597);
xnor U6005 (N_6005,N_5582,N_4970);
nor U6006 (N_6006,N_5430,N_5281);
or U6007 (N_6007,N_5470,N_5554);
nand U6008 (N_6008,N_5355,N_4984);
nand U6009 (N_6009,N_5386,N_5555);
and U6010 (N_6010,N_4807,N_5548);
xor U6011 (N_6011,N_5116,N_5405);
xnor U6012 (N_6012,N_5190,N_4819);
xor U6013 (N_6013,N_5090,N_5501);
or U6014 (N_6014,N_5175,N_5127);
nor U6015 (N_6015,N_5570,N_5147);
and U6016 (N_6016,N_4835,N_5398);
nand U6017 (N_6017,N_5471,N_4975);
nand U6018 (N_6018,N_4924,N_5500);
or U6019 (N_6019,N_4896,N_4965);
nor U6020 (N_6020,N_5216,N_5111);
xor U6021 (N_6021,N_5406,N_4809);
or U6022 (N_6022,N_5073,N_4965);
nor U6023 (N_6023,N_5100,N_4889);
and U6024 (N_6024,N_5598,N_5409);
and U6025 (N_6025,N_5128,N_5092);
or U6026 (N_6026,N_4987,N_5299);
and U6027 (N_6027,N_4852,N_4930);
or U6028 (N_6028,N_5092,N_4865);
or U6029 (N_6029,N_5440,N_5247);
or U6030 (N_6030,N_5114,N_5591);
xnor U6031 (N_6031,N_5130,N_5586);
nor U6032 (N_6032,N_5596,N_5021);
nor U6033 (N_6033,N_5389,N_5108);
and U6034 (N_6034,N_5549,N_4997);
or U6035 (N_6035,N_5516,N_5497);
and U6036 (N_6036,N_5038,N_5486);
nor U6037 (N_6037,N_5266,N_5505);
or U6038 (N_6038,N_5393,N_5220);
or U6039 (N_6039,N_4970,N_5351);
or U6040 (N_6040,N_5442,N_5275);
and U6041 (N_6041,N_4958,N_5369);
or U6042 (N_6042,N_4804,N_4895);
or U6043 (N_6043,N_4848,N_5114);
xor U6044 (N_6044,N_5541,N_5389);
xnor U6045 (N_6045,N_4964,N_5443);
nand U6046 (N_6046,N_5028,N_5187);
and U6047 (N_6047,N_5046,N_5344);
and U6048 (N_6048,N_5421,N_4911);
and U6049 (N_6049,N_5172,N_4855);
nor U6050 (N_6050,N_5552,N_5339);
or U6051 (N_6051,N_5184,N_5084);
and U6052 (N_6052,N_5030,N_5400);
xnor U6053 (N_6053,N_5016,N_5579);
xor U6054 (N_6054,N_5229,N_5434);
xor U6055 (N_6055,N_5141,N_4816);
nor U6056 (N_6056,N_5124,N_5075);
nor U6057 (N_6057,N_5106,N_5259);
or U6058 (N_6058,N_5295,N_5186);
nor U6059 (N_6059,N_4910,N_5422);
nand U6060 (N_6060,N_5428,N_5380);
xor U6061 (N_6061,N_5384,N_5062);
or U6062 (N_6062,N_5467,N_4990);
or U6063 (N_6063,N_5474,N_5055);
nand U6064 (N_6064,N_5034,N_5429);
nand U6065 (N_6065,N_5038,N_5557);
nand U6066 (N_6066,N_5059,N_4967);
xor U6067 (N_6067,N_4991,N_5499);
or U6068 (N_6068,N_4975,N_5147);
nor U6069 (N_6069,N_5579,N_4855);
or U6070 (N_6070,N_5232,N_5507);
nand U6071 (N_6071,N_5508,N_5077);
nand U6072 (N_6072,N_5412,N_5284);
and U6073 (N_6073,N_4987,N_4876);
and U6074 (N_6074,N_4946,N_4942);
xnor U6075 (N_6075,N_5589,N_5143);
nor U6076 (N_6076,N_5186,N_5544);
nand U6077 (N_6077,N_5360,N_4839);
and U6078 (N_6078,N_5339,N_5286);
nor U6079 (N_6079,N_5581,N_5059);
nor U6080 (N_6080,N_5430,N_4948);
nor U6081 (N_6081,N_5196,N_4921);
xor U6082 (N_6082,N_5537,N_5268);
xnor U6083 (N_6083,N_4851,N_5317);
xor U6084 (N_6084,N_5051,N_5081);
or U6085 (N_6085,N_5068,N_5240);
xnor U6086 (N_6086,N_4904,N_5359);
or U6087 (N_6087,N_5064,N_5020);
and U6088 (N_6088,N_5186,N_4859);
or U6089 (N_6089,N_5447,N_5558);
and U6090 (N_6090,N_5419,N_5463);
or U6091 (N_6091,N_5124,N_5212);
or U6092 (N_6092,N_4945,N_5595);
or U6093 (N_6093,N_5592,N_5138);
nand U6094 (N_6094,N_4840,N_5428);
or U6095 (N_6095,N_4955,N_4978);
xor U6096 (N_6096,N_4900,N_5435);
nor U6097 (N_6097,N_5108,N_5121);
or U6098 (N_6098,N_5200,N_5282);
and U6099 (N_6099,N_4813,N_5549);
nand U6100 (N_6100,N_5443,N_5314);
or U6101 (N_6101,N_5500,N_5355);
nor U6102 (N_6102,N_4959,N_5441);
xnor U6103 (N_6103,N_5425,N_5122);
xor U6104 (N_6104,N_5159,N_5250);
or U6105 (N_6105,N_5556,N_5096);
and U6106 (N_6106,N_5584,N_4884);
and U6107 (N_6107,N_5535,N_5030);
xor U6108 (N_6108,N_4867,N_4860);
nand U6109 (N_6109,N_5491,N_5288);
nor U6110 (N_6110,N_5081,N_4854);
or U6111 (N_6111,N_5376,N_4903);
or U6112 (N_6112,N_4807,N_5589);
and U6113 (N_6113,N_5586,N_4866);
nor U6114 (N_6114,N_4970,N_5249);
xnor U6115 (N_6115,N_5294,N_5017);
nor U6116 (N_6116,N_5307,N_4828);
or U6117 (N_6117,N_5540,N_5162);
xor U6118 (N_6118,N_5016,N_4845);
or U6119 (N_6119,N_4900,N_4987);
or U6120 (N_6120,N_5130,N_5582);
or U6121 (N_6121,N_5300,N_5129);
or U6122 (N_6122,N_5481,N_5018);
and U6123 (N_6123,N_5202,N_5168);
xor U6124 (N_6124,N_4977,N_5032);
and U6125 (N_6125,N_5215,N_5096);
nor U6126 (N_6126,N_4966,N_5525);
nand U6127 (N_6127,N_4850,N_5113);
and U6128 (N_6128,N_4924,N_5349);
nor U6129 (N_6129,N_5567,N_4857);
nand U6130 (N_6130,N_5516,N_5582);
nor U6131 (N_6131,N_5150,N_5378);
nor U6132 (N_6132,N_5315,N_4933);
and U6133 (N_6133,N_4830,N_5195);
and U6134 (N_6134,N_5059,N_5110);
xor U6135 (N_6135,N_5349,N_5330);
nand U6136 (N_6136,N_5200,N_5031);
and U6137 (N_6137,N_5191,N_5083);
or U6138 (N_6138,N_5303,N_4894);
xor U6139 (N_6139,N_5223,N_4845);
and U6140 (N_6140,N_5127,N_5545);
nor U6141 (N_6141,N_5123,N_5356);
nor U6142 (N_6142,N_4902,N_5440);
and U6143 (N_6143,N_5066,N_5393);
nand U6144 (N_6144,N_5323,N_5450);
nand U6145 (N_6145,N_5323,N_5593);
or U6146 (N_6146,N_5231,N_5479);
nor U6147 (N_6147,N_5114,N_5416);
nor U6148 (N_6148,N_5205,N_5526);
and U6149 (N_6149,N_5239,N_4835);
xor U6150 (N_6150,N_4910,N_5272);
nor U6151 (N_6151,N_4844,N_4926);
or U6152 (N_6152,N_5014,N_5314);
xor U6153 (N_6153,N_4866,N_5218);
xor U6154 (N_6154,N_5507,N_5477);
or U6155 (N_6155,N_5346,N_4917);
nor U6156 (N_6156,N_5093,N_5598);
nand U6157 (N_6157,N_4997,N_5000);
xor U6158 (N_6158,N_4859,N_5437);
nand U6159 (N_6159,N_5240,N_5097);
nand U6160 (N_6160,N_5546,N_5351);
nand U6161 (N_6161,N_5390,N_4803);
and U6162 (N_6162,N_5241,N_5039);
or U6163 (N_6163,N_5486,N_5575);
nor U6164 (N_6164,N_5328,N_5463);
nand U6165 (N_6165,N_5193,N_5155);
or U6166 (N_6166,N_5285,N_5115);
and U6167 (N_6167,N_5126,N_5553);
xor U6168 (N_6168,N_5001,N_5243);
nand U6169 (N_6169,N_5011,N_5486);
nor U6170 (N_6170,N_5129,N_5500);
xor U6171 (N_6171,N_4917,N_5057);
nor U6172 (N_6172,N_5505,N_4817);
nand U6173 (N_6173,N_5073,N_5083);
nand U6174 (N_6174,N_5370,N_4827);
and U6175 (N_6175,N_5325,N_5078);
nand U6176 (N_6176,N_5344,N_5311);
xor U6177 (N_6177,N_5444,N_5539);
and U6178 (N_6178,N_5412,N_4828);
and U6179 (N_6179,N_5010,N_5523);
nor U6180 (N_6180,N_5208,N_4964);
or U6181 (N_6181,N_5597,N_5236);
and U6182 (N_6182,N_4963,N_4874);
or U6183 (N_6183,N_5214,N_4899);
xor U6184 (N_6184,N_5110,N_5161);
or U6185 (N_6185,N_5491,N_5424);
or U6186 (N_6186,N_4866,N_4948);
or U6187 (N_6187,N_5187,N_5594);
xor U6188 (N_6188,N_5175,N_5419);
xor U6189 (N_6189,N_4911,N_5302);
xor U6190 (N_6190,N_5530,N_5030);
and U6191 (N_6191,N_5082,N_5536);
nand U6192 (N_6192,N_5535,N_5084);
nand U6193 (N_6193,N_5517,N_5002);
nand U6194 (N_6194,N_5472,N_5011);
and U6195 (N_6195,N_5283,N_5061);
and U6196 (N_6196,N_4816,N_4969);
and U6197 (N_6197,N_5245,N_5178);
or U6198 (N_6198,N_5306,N_5367);
or U6199 (N_6199,N_5571,N_4914);
nand U6200 (N_6200,N_5549,N_5319);
or U6201 (N_6201,N_5244,N_5421);
and U6202 (N_6202,N_5175,N_5042);
nor U6203 (N_6203,N_5477,N_5282);
and U6204 (N_6204,N_5572,N_4835);
xor U6205 (N_6205,N_5022,N_5205);
nor U6206 (N_6206,N_5358,N_5429);
and U6207 (N_6207,N_4973,N_4845);
or U6208 (N_6208,N_5316,N_4860);
xor U6209 (N_6209,N_5365,N_4889);
xor U6210 (N_6210,N_5305,N_5340);
or U6211 (N_6211,N_5150,N_5008);
and U6212 (N_6212,N_5462,N_5167);
and U6213 (N_6213,N_5383,N_5595);
xnor U6214 (N_6214,N_4884,N_5092);
nand U6215 (N_6215,N_4873,N_4993);
nor U6216 (N_6216,N_5309,N_4876);
xor U6217 (N_6217,N_5359,N_5076);
or U6218 (N_6218,N_5417,N_4852);
and U6219 (N_6219,N_5094,N_4822);
or U6220 (N_6220,N_4909,N_5190);
and U6221 (N_6221,N_5477,N_5269);
or U6222 (N_6222,N_4992,N_5206);
xnor U6223 (N_6223,N_5030,N_5153);
nor U6224 (N_6224,N_5452,N_5355);
or U6225 (N_6225,N_5595,N_5119);
and U6226 (N_6226,N_4918,N_4993);
or U6227 (N_6227,N_5233,N_5405);
nor U6228 (N_6228,N_5137,N_5065);
xor U6229 (N_6229,N_5427,N_5416);
and U6230 (N_6230,N_5151,N_4963);
and U6231 (N_6231,N_5251,N_5213);
xnor U6232 (N_6232,N_5120,N_5046);
xnor U6233 (N_6233,N_5531,N_5586);
and U6234 (N_6234,N_5121,N_5045);
and U6235 (N_6235,N_4842,N_5064);
and U6236 (N_6236,N_4859,N_5051);
nor U6237 (N_6237,N_5161,N_5244);
xnor U6238 (N_6238,N_5081,N_5376);
or U6239 (N_6239,N_5231,N_4986);
or U6240 (N_6240,N_5308,N_4870);
or U6241 (N_6241,N_5211,N_5219);
nand U6242 (N_6242,N_5361,N_5098);
or U6243 (N_6243,N_5228,N_5038);
or U6244 (N_6244,N_4834,N_5459);
nor U6245 (N_6245,N_5586,N_5334);
and U6246 (N_6246,N_5347,N_4908);
and U6247 (N_6247,N_5427,N_5480);
and U6248 (N_6248,N_5416,N_5187);
and U6249 (N_6249,N_4823,N_5491);
or U6250 (N_6250,N_5233,N_5559);
or U6251 (N_6251,N_5134,N_5302);
xor U6252 (N_6252,N_5508,N_5132);
and U6253 (N_6253,N_5240,N_4954);
and U6254 (N_6254,N_4840,N_5439);
or U6255 (N_6255,N_5272,N_5319);
and U6256 (N_6256,N_5083,N_4994);
nand U6257 (N_6257,N_5539,N_5498);
nor U6258 (N_6258,N_5185,N_5107);
nor U6259 (N_6259,N_5409,N_5253);
nor U6260 (N_6260,N_5399,N_5044);
nand U6261 (N_6261,N_5196,N_4939);
nor U6262 (N_6262,N_5577,N_5117);
nand U6263 (N_6263,N_5058,N_5405);
nand U6264 (N_6264,N_5574,N_5472);
nor U6265 (N_6265,N_4902,N_4875);
nor U6266 (N_6266,N_5009,N_5026);
nand U6267 (N_6267,N_5450,N_5220);
or U6268 (N_6268,N_5445,N_5275);
or U6269 (N_6269,N_5099,N_4981);
or U6270 (N_6270,N_5380,N_5072);
nand U6271 (N_6271,N_5224,N_5084);
xor U6272 (N_6272,N_5032,N_5116);
and U6273 (N_6273,N_5204,N_5571);
nor U6274 (N_6274,N_5350,N_4887);
and U6275 (N_6275,N_5589,N_5406);
nand U6276 (N_6276,N_5442,N_5555);
nor U6277 (N_6277,N_5539,N_5599);
xnor U6278 (N_6278,N_5446,N_4859);
nand U6279 (N_6279,N_5547,N_5135);
and U6280 (N_6280,N_5220,N_4876);
nor U6281 (N_6281,N_4996,N_5349);
nand U6282 (N_6282,N_4817,N_5445);
xnor U6283 (N_6283,N_5193,N_4870);
or U6284 (N_6284,N_5250,N_5564);
nand U6285 (N_6285,N_5007,N_4821);
and U6286 (N_6286,N_5388,N_5425);
or U6287 (N_6287,N_4934,N_5048);
or U6288 (N_6288,N_5559,N_5319);
or U6289 (N_6289,N_4883,N_5272);
xor U6290 (N_6290,N_5464,N_5096);
nor U6291 (N_6291,N_5263,N_5052);
xor U6292 (N_6292,N_5081,N_5365);
or U6293 (N_6293,N_5174,N_5420);
xnor U6294 (N_6294,N_5182,N_5432);
nor U6295 (N_6295,N_5254,N_5469);
xnor U6296 (N_6296,N_5220,N_5358);
or U6297 (N_6297,N_5296,N_5467);
xnor U6298 (N_6298,N_5501,N_5152);
xnor U6299 (N_6299,N_5176,N_5554);
xnor U6300 (N_6300,N_5559,N_5398);
xnor U6301 (N_6301,N_5183,N_5074);
nor U6302 (N_6302,N_5362,N_4806);
and U6303 (N_6303,N_5204,N_5427);
or U6304 (N_6304,N_5587,N_5579);
xor U6305 (N_6305,N_5306,N_5209);
nor U6306 (N_6306,N_5179,N_5585);
xnor U6307 (N_6307,N_5584,N_5292);
nand U6308 (N_6308,N_5552,N_5425);
or U6309 (N_6309,N_5537,N_4818);
xnor U6310 (N_6310,N_5373,N_5260);
nand U6311 (N_6311,N_5252,N_4986);
or U6312 (N_6312,N_5523,N_5021);
xnor U6313 (N_6313,N_5472,N_5192);
and U6314 (N_6314,N_5407,N_4877);
nor U6315 (N_6315,N_4977,N_5549);
or U6316 (N_6316,N_5001,N_5554);
and U6317 (N_6317,N_5540,N_4917);
xor U6318 (N_6318,N_5557,N_4893);
and U6319 (N_6319,N_4859,N_5170);
nor U6320 (N_6320,N_5562,N_5221);
nand U6321 (N_6321,N_5494,N_5326);
and U6322 (N_6322,N_4842,N_5103);
or U6323 (N_6323,N_4925,N_4923);
nand U6324 (N_6324,N_5254,N_5345);
nor U6325 (N_6325,N_5157,N_5246);
or U6326 (N_6326,N_4818,N_5223);
xor U6327 (N_6327,N_5574,N_5092);
or U6328 (N_6328,N_5372,N_5404);
nand U6329 (N_6329,N_4857,N_4973);
or U6330 (N_6330,N_5599,N_4840);
and U6331 (N_6331,N_5491,N_4908);
xor U6332 (N_6332,N_4985,N_5495);
and U6333 (N_6333,N_5571,N_4967);
xnor U6334 (N_6334,N_4937,N_5154);
nand U6335 (N_6335,N_5121,N_4860);
nor U6336 (N_6336,N_5438,N_5398);
nor U6337 (N_6337,N_5160,N_5054);
and U6338 (N_6338,N_4891,N_5027);
nor U6339 (N_6339,N_5311,N_5455);
or U6340 (N_6340,N_5323,N_5545);
nand U6341 (N_6341,N_5486,N_5583);
nor U6342 (N_6342,N_4828,N_4904);
nand U6343 (N_6343,N_5400,N_5420);
and U6344 (N_6344,N_5336,N_5046);
nand U6345 (N_6345,N_5475,N_5503);
or U6346 (N_6346,N_4929,N_5515);
nor U6347 (N_6347,N_5500,N_5071);
nand U6348 (N_6348,N_5028,N_5241);
nand U6349 (N_6349,N_4832,N_5307);
xor U6350 (N_6350,N_5568,N_4811);
nand U6351 (N_6351,N_5412,N_4912);
xnor U6352 (N_6352,N_5503,N_5563);
nand U6353 (N_6353,N_4902,N_5304);
xnor U6354 (N_6354,N_4913,N_5054);
nand U6355 (N_6355,N_5592,N_5526);
or U6356 (N_6356,N_5121,N_5010);
nand U6357 (N_6357,N_5300,N_4830);
and U6358 (N_6358,N_5021,N_4921);
nor U6359 (N_6359,N_5035,N_4822);
nor U6360 (N_6360,N_5302,N_5431);
or U6361 (N_6361,N_5044,N_5592);
or U6362 (N_6362,N_4923,N_5219);
nand U6363 (N_6363,N_4826,N_5548);
or U6364 (N_6364,N_4989,N_5000);
or U6365 (N_6365,N_5548,N_5542);
or U6366 (N_6366,N_4862,N_5483);
nand U6367 (N_6367,N_5586,N_5111);
xnor U6368 (N_6368,N_5486,N_4974);
nand U6369 (N_6369,N_4891,N_5578);
or U6370 (N_6370,N_5339,N_5541);
nand U6371 (N_6371,N_4978,N_4928);
nor U6372 (N_6372,N_4806,N_5156);
xor U6373 (N_6373,N_5445,N_5342);
xnor U6374 (N_6374,N_5473,N_5189);
nand U6375 (N_6375,N_5569,N_5556);
or U6376 (N_6376,N_5069,N_5249);
or U6377 (N_6377,N_5430,N_5493);
nand U6378 (N_6378,N_5472,N_5562);
xnor U6379 (N_6379,N_5105,N_4803);
and U6380 (N_6380,N_5036,N_5355);
nand U6381 (N_6381,N_5282,N_5207);
and U6382 (N_6382,N_5111,N_5207);
or U6383 (N_6383,N_4865,N_4945);
xor U6384 (N_6384,N_4966,N_5291);
nor U6385 (N_6385,N_4941,N_5483);
nand U6386 (N_6386,N_5428,N_5548);
nand U6387 (N_6387,N_5349,N_4956);
or U6388 (N_6388,N_4877,N_5313);
nand U6389 (N_6389,N_5008,N_5456);
nor U6390 (N_6390,N_5322,N_5474);
and U6391 (N_6391,N_5134,N_5433);
or U6392 (N_6392,N_4866,N_5410);
or U6393 (N_6393,N_5009,N_5253);
or U6394 (N_6394,N_4855,N_4888);
xor U6395 (N_6395,N_5428,N_5434);
xor U6396 (N_6396,N_5381,N_4802);
or U6397 (N_6397,N_4865,N_4933);
or U6398 (N_6398,N_5214,N_5169);
nand U6399 (N_6399,N_5472,N_5200);
and U6400 (N_6400,N_5747,N_5883);
and U6401 (N_6401,N_6314,N_5653);
or U6402 (N_6402,N_6088,N_6096);
or U6403 (N_6403,N_6054,N_5703);
nor U6404 (N_6404,N_6195,N_5831);
nand U6405 (N_6405,N_5956,N_6152);
nand U6406 (N_6406,N_5977,N_5938);
nor U6407 (N_6407,N_5765,N_5855);
nand U6408 (N_6408,N_6224,N_6352);
or U6409 (N_6409,N_5925,N_6082);
xor U6410 (N_6410,N_5948,N_5662);
or U6411 (N_6411,N_6145,N_6377);
or U6412 (N_6412,N_6131,N_5716);
nand U6413 (N_6413,N_6237,N_5897);
and U6414 (N_6414,N_5699,N_6239);
nand U6415 (N_6415,N_6127,N_5970);
or U6416 (N_6416,N_5908,N_5763);
nor U6417 (N_6417,N_6147,N_6126);
xor U6418 (N_6418,N_6020,N_5713);
nand U6419 (N_6419,N_5993,N_5959);
or U6420 (N_6420,N_5958,N_5992);
and U6421 (N_6421,N_5835,N_5625);
or U6422 (N_6422,N_6039,N_5648);
nand U6423 (N_6423,N_6032,N_6365);
xor U6424 (N_6424,N_5893,N_6109);
nor U6425 (N_6425,N_5787,N_5861);
or U6426 (N_6426,N_5687,N_6396);
or U6427 (N_6427,N_5769,N_6087);
and U6428 (N_6428,N_6036,N_6299);
nand U6429 (N_6429,N_6332,N_5912);
xor U6430 (N_6430,N_5628,N_5878);
xor U6431 (N_6431,N_5966,N_5691);
nand U6432 (N_6432,N_6001,N_6155);
xnor U6433 (N_6433,N_6010,N_5882);
nand U6434 (N_6434,N_6230,N_5936);
and U6435 (N_6435,N_6367,N_5756);
nand U6436 (N_6436,N_6372,N_6395);
nor U6437 (N_6437,N_5999,N_6053);
nor U6438 (N_6438,N_5867,N_6236);
or U6439 (N_6439,N_6258,N_6313);
and U6440 (N_6440,N_6295,N_6186);
xnor U6441 (N_6441,N_5899,N_6385);
and U6442 (N_6442,N_6300,N_5918);
xnor U6443 (N_6443,N_6283,N_6388);
xnor U6444 (N_6444,N_5829,N_6334);
and U6445 (N_6445,N_6103,N_5904);
xor U6446 (N_6446,N_6312,N_5996);
nor U6447 (N_6447,N_6322,N_6264);
and U6448 (N_6448,N_6217,N_5683);
and U6449 (N_6449,N_6046,N_5749);
or U6450 (N_6450,N_5984,N_5907);
or U6451 (N_6451,N_5813,N_6132);
and U6452 (N_6452,N_6059,N_5913);
and U6453 (N_6453,N_5608,N_5668);
xor U6454 (N_6454,N_6221,N_6113);
or U6455 (N_6455,N_5611,N_5737);
nor U6456 (N_6456,N_6292,N_6320);
and U6457 (N_6457,N_5927,N_5660);
or U6458 (N_6458,N_5946,N_5640);
nor U6459 (N_6459,N_5890,N_6285);
nand U6460 (N_6460,N_5681,N_5785);
nor U6461 (N_6461,N_6029,N_5847);
xnor U6462 (N_6462,N_6354,N_5783);
and U6463 (N_6463,N_5857,N_5926);
xor U6464 (N_6464,N_5770,N_6184);
nor U6465 (N_6465,N_6199,N_6319);
nand U6466 (N_6466,N_5862,N_5950);
and U6467 (N_6467,N_6062,N_5606);
nand U6468 (N_6468,N_5663,N_6159);
or U6469 (N_6469,N_5605,N_6247);
and U6470 (N_6470,N_5814,N_6222);
nor U6471 (N_6471,N_5782,N_5824);
or U6472 (N_6472,N_5607,N_6212);
nor U6473 (N_6473,N_5971,N_6187);
and U6474 (N_6474,N_5869,N_5788);
or U6475 (N_6475,N_5851,N_6047);
nor U6476 (N_6476,N_6233,N_5828);
nor U6477 (N_6477,N_5886,N_6343);
nand U6478 (N_6478,N_5807,N_5836);
and U6479 (N_6479,N_5771,N_5885);
or U6480 (N_6480,N_5614,N_6137);
nor U6481 (N_6481,N_5715,N_5643);
xnor U6482 (N_6482,N_6191,N_5953);
or U6483 (N_6483,N_6333,N_5811);
nor U6484 (N_6484,N_5759,N_6148);
and U6485 (N_6485,N_6323,N_5638);
or U6486 (N_6486,N_5932,N_5766);
or U6487 (N_6487,N_5641,N_5916);
nand U6488 (N_6488,N_5994,N_6209);
xor U6489 (N_6489,N_5985,N_5854);
and U6490 (N_6490,N_6038,N_5777);
and U6491 (N_6491,N_6100,N_5838);
and U6492 (N_6492,N_5955,N_6275);
nor U6493 (N_6493,N_5772,N_5945);
nor U6494 (N_6494,N_6269,N_6043);
xor U6495 (N_6495,N_5998,N_6241);
and U6496 (N_6496,N_5613,N_6007);
and U6497 (N_6497,N_5930,N_6041);
and U6498 (N_6498,N_5963,N_5701);
xnor U6499 (N_6499,N_6146,N_5744);
nor U6500 (N_6500,N_6393,N_6390);
xor U6501 (N_6501,N_5919,N_6144);
xnor U6502 (N_6502,N_6071,N_5892);
or U6503 (N_6503,N_6073,N_6302);
or U6504 (N_6504,N_5859,N_6359);
nor U6505 (N_6505,N_6358,N_6143);
or U6506 (N_6506,N_5724,N_5793);
nor U6507 (N_6507,N_5740,N_6339);
xnor U6508 (N_6508,N_5609,N_5627);
and U6509 (N_6509,N_5979,N_6213);
nand U6510 (N_6510,N_5820,N_5942);
xnor U6511 (N_6511,N_5898,N_5610);
nand U6512 (N_6512,N_6242,N_6290);
nand U6513 (N_6513,N_6198,N_6200);
and U6514 (N_6514,N_5712,N_5846);
and U6515 (N_6515,N_5686,N_5839);
and U6516 (N_6516,N_5750,N_6014);
and U6517 (N_6517,N_5937,N_6348);
and U6518 (N_6518,N_6060,N_6092);
or U6519 (N_6519,N_6021,N_5619);
nor U6520 (N_6520,N_6130,N_6154);
xnor U6521 (N_6521,N_5949,N_5990);
or U6522 (N_6522,N_6067,N_5853);
nor U6523 (N_6523,N_5844,N_5733);
nor U6524 (N_6524,N_5791,N_6265);
or U6525 (N_6525,N_5741,N_5708);
xnor U6526 (N_6526,N_6114,N_5832);
nand U6527 (N_6527,N_6211,N_6136);
nand U6528 (N_6528,N_6140,N_6015);
nor U6529 (N_6529,N_6080,N_5626);
nand U6530 (N_6530,N_6316,N_6279);
nor U6531 (N_6531,N_5805,N_6260);
nor U6532 (N_6532,N_5909,N_6360);
nor U6533 (N_6533,N_5714,N_6037);
and U6534 (N_6534,N_6185,N_5794);
nor U6535 (N_6535,N_6263,N_5612);
xor U6536 (N_6536,N_5685,N_5901);
nor U6537 (N_6537,N_5623,N_5721);
nand U6538 (N_6538,N_5666,N_5603);
nor U6539 (N_6539,N_6347,N_6251);
nand U6540 (N_6540,N_5726,N_5997);
and U6541 (N_6541,N_6068,N_5727);
nand U6542 (N_6542,N_6035,N_6381);
xor U6543 (N_6543,N_6086,N_5843);
and U6544 (N_6544,N_5705,N_5808);
nor U6545 (N_6545,N_5818,N_5644);
nor U6546 (N_6546,N_6289,N_6017);
nand U6547 (N_6547,N_5774,N_6050);
or U6548 (N_6548,N_5864,N_5696);
nand U6549 (N_6549,N_5887,N_6350);
nor U6550 (N_6550,N_5986,N_6028);
nand U6551 (N_6551,N_6214,N_5943);
xnor U6552 (N_6552,N_6379,N_6244);
xnor U6553 (N_6553,N_6376,N_5669);
xnor U6554 (N_6554,N_5917,N_6326);
nand U6555 (N_6555,N_5934,N_6123);
or U6556 (N_6556,N_6064,N_6201);
nand U6557 (N_6557,N_5929,N_5694);
and U6558 (N_6558,N_6125,N_6108);
xor U6559 (N_6559,N_6206,N_6169);
and U6560 (N_6560,N_6077,N_6194);
and U6561 (N_6561,N_5654,N_5753);
and U6562 (N_6562,N_6139,N_5764);
xor U6563 (N_6563,N_6386,N_6327);
xnor U6564 (N_6564,N_6133,N_6234);
nor U6565 (N_6565,N_5903,N_6262);
xnor U6566 (N_6566,N_6363,N_6156);
xnor U6567 (N_6567,N_6016,N_5863);
xnor U6568 (N_6568,N_6177,N_6141);
nor U6569 (N_6569,N_6399,N_5841);
xor U6570 (N_6570,N_5856,N_6192);
xnor U6571 (N_6571,N_6164,N_5967);
nor U6572 (N_6572,N_6383,N_5974);
nand U6573 (N_6573,N_6370,N_5815);
and U6574 (N_6574,N_6034,N_6346);
or U6575 (N_6575,N_6368,N_5889);
or U6576 (N_6576,N_6324,N_6303);
nor U6577 (N_6577,N_5884,N_6353);
or U6578 (N_6578,N_6072,N_6150);
nor U6579 (N_6579,N_5827,N_5975);
nand U6580 (N_6580,N_5664,N_5751);
nand U6581 (N_6581,N_5928,N_5707);
nand U6582 (N_6582,N_6189,N_6340);
or U6583 (N_6583,N_6170,N_6120);
and U6584 (N_6584,N_5639,N_6274);
xor U6585 (N_6585,N_5803,N_6066);
and U6586 (N_6586,N_6078,N_6351);
and U6587 (N_6587,N_5631,N_5972);
and U6588 (N_6588,N_5978,N_6305);
and U6589 (N_6589,N_6387,N_6098);
nor U6590 (N_6590,N_6196,N_6294);
or U6591 (N_6591,N_6134,N_6249);
xnor U6592 (N_6592,N_6093,N_6095);
or U6593 (N_6593,N_5939,N_6268);
nand U6594 (N_6594,N_5888,N_6138);
xnor U6595 (N_6595,N_5840,N_5849);
nand U6596 (N_6596,N_6012,N_5902);
and U6597 (N_6597,N_5761,N_6124);
nand U6598 (N_6598,N_6118,N_6374);
nor U6599 (N_6599,N_5657,N_6297);
or U6600 (N_6600,N_5776,N_5935);
or U6601 (N_6601,N_6119,N_5702);
or U6602 (N_6602,N_5632,N_5800);
and U6603 (N_6603,N_5693,N_6380);
nand U6604 (N_6604,N_5768,N_6208);
xor U6605 (N_6605,N_5743,N_5752);
and U6606 (N_6606,N_6031,N_5722);
and U6607 (N_6607,N_5602,N_5822);
nor U6608 (N_6608,N_6129,N_6165);
nand U6609 (N_6609,N_6040,N_5758);
nand U6610 (N_6610,N_5674,N_5717);
xor U6611 (N_6611,N_6336,N_5624);
and U6612 (N_6612,N_5601,N_6135);
and U6613 (N_6613,N_6398,N_6063);
and U6614 (N_6614,N_6307,N_5915);
or U6615 (N_6615,N_6005,N_6003);
xnor U6616 (N_6616,N_6219,N_6278);
and U6617 (N_6617,N_5621,N_6277);
nand U6618 (N_6618,N_6267,N_5672);
nor U6619 (N_6619,N_6161,N_6330);
or U6620 (N_6620,N_5731,N_6254);
or U6621 (N_6621,N_5940,N_6094);
xnor U6622 (N_6622,N_6030,N_5637);
xor U6623 (N_6623,N_5826,N_6178);
nor U6624 (N_6624,N_5665,N_6061);
and U6625 (N_6625,N_5629,N_5786);
nor U6626 (N_6626,N_6057,N_5636);
nand U6627 (N_6627,N_6105,N_6171);
or U6628 (N_6628,N_5634,N_6345);
xnor U6629 (N_6629,N_6309,N_6231);
and U6630 (N_6630,N_6070,N_5690);
nor U6631 (N_6631,N_5630,N_5905);
nand U6632 (N_6632,N_5812,N_6253);
nand U6633 (N_6633,N_6325,N_5842);
and U6634 (N_6634,N_6227,N_6378);
or U6635 (N_6635,N_5987,N_6321);
nor U6636 (N_6636,N_6104,N_5921);
and U6637 (N_6637,N_5989,N_5865);
or U6638 (N_6638,N_6301,N_5645);
xor U6639 (N_6639,N_5894,N_5679);
and U6640 (N_6640,N_6287,N_6122);
xnor U6641 (N_6641,N_5745,N_6250);
nand U6642 (N_6642,N_6157,N_6284);
nand U6643 (N_6643,N_6293,N_6190);
xor U6644 (N_6644,N_6252,N_5700);
or U6645 (N_6645,N_5675,N_6115);
nand U6646 (N_6646,N_6162,N_5806);
or U6647 (N_6647,N_6022,N_5834);
nand U6648 (N_6648,N_5684,N_5848);
and U6649 (N_6649,N_5868,N_6291);
nand U6650 (N_6650,N_6090,N_5615);
or U6651 (N_6651,N_6218,N_5760);
nand U6652 (N_6652,N_6153,N_5649);
xor U6653 (N_6653,N_5661,N_5875);
xor U6654 (N_6654,N_5757,N_6202);
and U6655 (N_6655,N_6025,N_6308);
xor U6656 (N_6656,N_6270,N_5973);
nor U6657 (N_6657,N_5964,N_6013);
and U6658 (N_6658,N_6052,N_6331);
nand U6659 (N_6659,N_5646,N_5981);
nand U6660 (N_6660,N_6344,N_5656);
nor U6661 (N_6661,N_5647,N_5866);
or U6662 (N_6662,N_5697,N_5952);
xor U6663 (N_6663,N_5845,N_6329);
and U6664 (N_6664,N_5695,N_6280);
nand U6665 (N_6665,N_5906,N_5962);
nor U6666 (N_6666,N_6175,N_6366);
nand U6667 (N_6667,N_5742,N_6328);
xnor U6668 (N_6668,N_5947,N_5732);
xnor U6669 (N_6669,N_5746,N_6205);
xnor U6670 (N_6670,N_6166,N_5725);
or U6671 (N_6671,N_5704,N_5873);
or U6672 (N_6672,N_5976,N_6226);
or U6673 (N_6673,N_5980,N_6364);
xnor U6674 (N_6674,N_6009,N_5735);
nor U6675 (N_6675,N_5604,N_6232);
xnor U6676 (N_6676,N_6207,N_6311);
nand U6677 (N_6677,N_6282,N_5659);
and U6678 (N_6678,N_5830,N_6272);
and U6679 (N_6679,N_5655,N_6048);
nand U6680 (N_6680,N_5652,N_5819);
or U6681 (N_6681,N_6304,N_6117);
xnor U6682 (N_6682,N_5635,N_5874);
xor U6683 (N_6683,N_6042,N_5891);
nand U6684 (N_6684,N_6341,N_6128);
nand U6685 (N_6685,N_6188,N_6392);
and U6686 (N_6686,N_6179,N_6197);
xnor U6687 (N_6687,N_6079,N_5991);
nand U6688 (N_6688,N_6288,N_5692);
and U6689 (N_6689,N_5804,N_6255);
and U6690 (N_6690,N_6369,N_6055);
xor U6691 (N_6691,N_6315,N_5775);
or U6692 (N_6692,N_5858,N_6158);
or U6693 (N_6693,N_6389,N_5651);
nand U6694 (N_6694,N_5723,N_5730);
and U6695 (N_6695,N_5870,N_5728);
nand U6696 (N_6696,N_5642,N_5957);
and U6697 (N_6697,N_6203,N_5982);
nor U6698 (N_6698,N_6357,N_6121);
nand U6699 (N_6699,N_6110,N_5738);
nand U6700 (N_6700,N_5880,N_6167);
nand U6701 (N_6701,N_5739,N_5680);
nand U6702 (N_6702,N_6318,N_5821);
and U6703 (N_6703,N_6044,N_5670);
and U6704 (N_6704,N_6210,N_5881);
nand U6705 (N_6705,N_6019,N_6225);
xor U6706 (N_6706,N_6271,N_6228);
xnor U6707 (N_6707,N_6384,N_5689);
and U6708 (N_6708,N_5924,N_5837);
nor U6709 (N_6709,N_5798,N_6083);
nand U6710 (N_6710,N_6394,N_6023);
nand U6711 (N_6711,N_5781,N_6089);
nor U6712 (N_6712,N_6342,N_5754);
nor U6713 (N_6713,N_5677,N_5922);
and U6714 (N_6714,N_6002,N_6204);
or U6715 (N_6715,N_5778,N_5796);
or U6716 (N_6716,N_6182,N_5850);
nand U6717 (N_6717,N_5809,N_6391);
and U6718 (N_6718,N_5789,N_5673);
nand U6719 (N_6719,N_6337,N_5944);
nand U6720 (N_6720,N_5709,N_6049);
xnor U6721 (N_6721,N_5816,N_5682);
xnor U6722 (N_6722,N_6229,N_6116);
nand U6723 (N_6723,N_6168,N_5734);
xor U6724 (N_6724,N_6276,N_5895);
or U6725 (N_6725,N_6261,N_5871);
nand U6726 (N_6726,N_6102,N_5876);
or U6727 (N_6727,N_6142,N_5988);
or U6728 (N_6728,N_5931,N_5622);
nand U6729 (N_6729,N_5698,N_5923);
and U6730 (N_6730,N_6349,N_6298);
xnor U6731 (N_6731,N_6018,N_6076);
and U6732 (N_6732,N_5933,N_6084);
xnor U6733 (N_6733,N_6317,N_6273);
and U6734 (N_6734,N_5762,N_6051);
xor U6735 (N_6735,N_6151,N_6355);
nor U6736 (N_6736,N_6246,N_6174);
nor U6737 (N_6737,N_6215,N_5706);
or U6738 (N_6738,N_6008,N_6006);
or U6739 (N_6739,N_5633,N_5790);
or U6740 (N_6740,N_6361,N_5667);
or U6741 (N_6741,N_5961,N_5823);
xor U6742 (N_6742,N_6160,N_6243);
nand U6743 (N_6743,N_5620,N_5658);
and U6744 (N_6744,N_5954,N_5920);
nand U6745 (N_6745,N_5600,N_5780);
nand U6746 (N_6746,N_5710,N_6306);
or U6747 (N_6747,N_6257,N_5792);
nand U6748 (N_6748,N_6296,N_5914);
xnor U6749 (N_6749,N_6173,N_6149);
nor U6750 (N_6750,N_6180,N_6172);
nand U6751 (N_6751,N_5617,N_5720);
xor U6752 (N_6752,N_5773,N_5736);
xnor U6753 (N_6753,N_5900,N_6111);
and U6754 (N_6754,N_6091,N_5779);
and U6755 (N_6755,N_5784,N_5951);
nor U6756 (N_6756,N_6235,N_6163);
and U6757 (N_6757,N_6220,N_6081);
and U6758 (N_6758,N_6112,N_6065);
or U6759 (N_6759,N_6238,N_5995);
and U6760 (N_6760,N_6075,N_5729);
nor U6761 (N_6761,N_5676,N_5941);
or U6762 (N_6762,N_5896,N_5872);
xor U6763 (N_6763,N_5616,N_5833);
or U6764 (N_6764,N_5860,N_6382);
nand U6765 (N_6765,N_6027,N_5960);
nand U6766 (N_6766,N_6256,N_5968);
nor U6767 (N_6767,N_6176,N_5767);
nand U6768 (N_6768,N_6056,N_5825);
or U6769 (N_6769,N_6101,N_6085);
xnor U6770 (N_6770,N_6011,N_6335);
or U6771 (N_6771,N_6097,N_6266);
or U6772 (N_6772,N_5965,N_6245);
xnor U6773 (N_6773,N_5618,N_6033);
nor U6774 (N_6774,N_6373,N_6338);
and U6775 (N_6775,N_6106,N_5817);
xnor U6776 (N_6776,N_6107,N_5877);
or U6777 (N_6777,N_6281,N_6004);
nor U6778 (N_6778,N_6216,N_6026);
nand U6779 (N_6779,N_6259,N_6024);
nand U6780 (N_6780,N_5802,N_5969);
or U6781 (N_6781,N_6397,N_5671);
or U6782 (N_6782,N_6248,N_5799);
xor U6783 (N_6783,N_6183,N_6286);
xnor U6784 (N_6784,N_5650,N_5748);
nor U6785 (N_6785,N_5983,N_6099);
and U6786 (N_6786,N_5910,N_5911);
nor U6787 (N_6787,N_5711,N_6069);
or U6788 (N_6788,N_5810,N_5879);
or U6789 (N_6789,N_6375,N_6074);
nand U6790 (N_6790,N_6181,N_5718);
nand U6791 (N_6791,N_5688,N_5755);
nand U6792 (N_6792,N_5852,N_6045);
nand U6793 (N_6793,N_5801,N_6240);
or U6794 (N_6794,N_6223,N_6000);
or U6795 (N_6795,N_6193,N_5795);
or U6796 (N_6796,N_6362,N_5797);
nor U6797 (N_6797,N_5719,N_6058);
nor U6798 (N_6798,N_6356,N_5678);
nor U6799 (N_6799,N_6310,N_6371);
and U6800 (N_6800,N_5881,N_6226);
nor U6801 (N_6801,N_5787,N_6150);
nand U6802 (N_6802,N_5649,N_5722);
or U6803 (N_6803,N_5779,N_6347);
and U6804 (N_6804,N_6093,N_5880);
or U6805 (N_6805,N_5627,N_5894);
xor U6806 (N_6806,N_5709,N_6246);
or U6807 (N_6807,N_5653,N_5700);
xor U6808 (N_6808,N_6254,N_6194);
and U6809 (N_6809,N_5708,N_6212);
nand U6810 (N_6810,N_6213,N_6015);
xnor U6811 (N_6811,N_5992,N_5784);
and U6812 (N_6812,N_6063,N_5806);
nor U6813 (N_6813,N_6171,N_5616);
nor U6814 (N_6814,N_6115,N_6332);
xnor U6815 (N_6815,N_6093,N_5858);
nor U6816 (N_6816,N_6347,N_6183);
or U6817 (N_6817,N_5702,N_6103);
nor U6818 (N_6818,N_5882,N_5726);
xor U6819 (N_6819,N_5768,N_6153);
or U6820 (N_6820,N_5639,N_6026);
nand U6821 (N_6821,N_5834,N_5656);
or U6822 (N_6822,N_5801,N_5997);
nor U6823 (N_6823,N_5647,N_6321);
nor U6824 (N_6824,N_5612,N_5702);
or U6825 (N_6825,N_6154,N_5930);
and U6826 (N_6826,N_6351,N_5693);
nand U6827 (N_6827,N_6123,N_6338);
nand U6828 (N_6828,N_5843,N_6089);
xor U6829 (N_6829,N_5978,N_6213);
and U6830 (N_6830,N_6155,N_5838);
xnor U6831 (N_6831,N_6054,N_5657);
or U6832 (N_6832,N_5715,N_6048);
xnor U6833 (N_6833,N_6023,N_5799);
nand U6834 (N_6834,N_5904,N_6369);
or U6835 (N_6835,N_6333,N_5981);
nand U6836 (N_6836,N_5883,N_5809);
xor U6837 (N_6837,N_5675,N_5792);
nand U6838 (N_6838,N_5900,N_6120);
nand U6839 (N_6839,N_5604,N_5996);
xnor U6840 (N_6840,N_6296,N_5866);
xnor U6841 (N_6841,N_5674,N_5670);
or U6842 (N_6842,N_5874,N_6093);
nand U6843 (N_6843,N_6012,N_5628);
xnor U6844 (N_6844,N_6134,N_5961);
xor U6845 (N_6845,N_5761,N_5668);
nand U6846 (N_6846,N_5953,N_6333);
nand U6847 (N_6847,N_5935,N_6112);
or U6848 (N_6848,N_6271,N_5816);
nor U6849 (N_6849,N_6121,N_6021);
nand U6850 (N_6850,N_5755,N_5958);
nand U6851 (N_6851,N_5860,N_6191);
and U6852 (N_6852,N_5745,N_5673);
nor U6853 (N_6853,N_6365,N_6316);
nor U6854 (N_6854,N_6173,N_5608);
xor U6855 (N_6855,N_6158,N_6131);
and U6856 (N_6856,N_6300,N_6374);
and U6857 (N_6857,N_6095,N_6044);
nor U6858 (N_6858,N_6166,N_5818);
or U6859 (N_6859,N_5909,N_5972);
or U6860 (N_6860,N_6296,N_6139);
nor U6861 (N_6861,N_5758,N_6003);
nand U6862 (N_6862,N_6183,N_5797);
nor U6863 (N_6863,N_6049,N_6198);
xor U6864 (N_6864,N_5609,N_6137);
nand U6865 (N_6865,N_5940,N_6346);
nand U6866 (N_6866,N_6033,N_5901);
xnor U6867 (N_6867,N_6082,N_5783);
or U6868 (N_6868,N_6337,N_5635);
nand U6869 (N_6869,N_6046,N_5632);
and U6870 (N_6870,N_5997,N_5704);
xor U6871 (N_6871,N_6293,N_5852);
nor U6872 (N_6872,N_5622,N_5937);
nand U6873 (N_6873,N_5775,N_5912);
xor U6874 (N_6874,N_5620,N_5774);
and U6875 (N_6875,N_6243,N_5864);
nand U6876 (N_6876,N_6368,N_6035);
nand U6877 (N_6877,N_5885,N_6272);
nor U6878 (N_6878,N_6221,N_5642);
or U6879 (N_6879,N_6135,N_5846);
and U6880 (N_6880,N_6150,N_5713);
nor U6881 (N_6881,N_5908,N_5802);
and U6882 (N_6882,N_5813,N_5656);
nor U6883 (N_6883,N_6292,N_5985);
nor U6884 (N_6884,N_6097,N_5695);
and U6885 (N_6885,N_5643,N_6071);
and U6886 (N_6886,N_6218,N_5924);
nand U6887 (N_6887,N_5923,N_6017);
nand U6888 (N_6888,N_6006,N_5649);
nor U6889 (N_6889,N_6069,N_5975);
and U6890 (N_6890,N_5936,N_6343);
nand U6891 (N_6891,N_6040,N_6001);
nor U6892 (N_6892,N_6322,N_5641);
xor U6893 (N_6893,N_6189,N_6378);
and U6894 (N_6894,N_6216,N_5954);
and U6895 (N_6895,N_6239,N_5714);
or U6896 (N_6896,N_6343,N_6361);
xor U6897 (N_6897,N_5608,N_5611);
nand U6898 (N_6898,N_6055,N_6033);
or U6899 (N_6899,N_5859,N_6144);
nand U6900 (N_6900,N_6319,N_6291);
nor U6901 (N_6901,N_6257,N_6315);
and U6902 (N_6902,N_5989,N_6190);
xnor U6903 (N_6903,N_5953,N_6127);
nor U6904 (N_6904,N_6043,N_6348);
xnor U6905 (N_6905,N_5955,N_5601);
and U6906 (N_6906,N_5780,N_6314);
nor U6907 (N_6907,N_6386,N_5656);
xor U6908 (N_6908,N_5610,N_6244);
nor U6909 (N_6909,N_5797,N_5903);
and U6910 (N_6910,N_5843,N_6272);
nor U6911 (N_6911,N_6303,N_5816);
and U6912 (N_6912,N_6384,N_6107);
nand U6913 (N_6913,N_6370,N_6393);
xor U6914 (N_6914,N_5846,N_5970);
xor U6915 (N_6915,N_6016,N_5748);
nand U6916 (N_6916,N_6032,N_5833);
xnor U6917 (N_6917,N_6013,N_6320);
nor U6918 (N_6918,N_6287,N_5861);
and U6919 (N_6919,N_6070,N_6260);
nor U6920 (N_6920,N_6287,N_6215);
or U6921 (N_6921,N_5821,N_6238);
nor U6922 (N_6922,N_5846,N_6093);
nor U6923 (N_6923,N_6373,N_6330);
or U6924 (N_6924,N_6009,N_6267);
nand U6925 (N_6925,N_6350,N_6101);
nor U6926 (N_6926,N_6159,N_5757);
nand U6927 (N_6927,N_6122,N_6360);
and U6928 (N_6928,N_5849,N_6116);
nor U6929 (N_6929,N_5648,N_5855);
or U6930 (N_6930,N_6333,N_5951);
nor U6931 (N_6931,N_5700,N_6374);
nand U6932 (N_6932,N_6046,N_5862);
nand U6933 (N_6933,N_6118,N_6324);
nor U6934 (N_6934,N_5655,N_6142);
nand U6935 (N_6935,N_6102,N_5600);
xor U6936 (N_6936,N_5977,N_5941);
xnor U6937 (N_6937,N_6076,N_6032);
and U6938 (N_6938,N_6003,N_6226);
xnor U6939 (N_6939,N_5984,N_6372);
xor U6940 (N_6940,N_5944,N_6224);
or U6941 (N_6941,N_5967,N_6067);
xor U6942 (N_6942,N_5697,N_5988);
or U6943 (N_6943,N_5659,N_6179);
xnor U6944 (N_6944,N_5952,N_5861);
and U6945 (N_6945,N_6259,N_6327);
or U6946 (N_6946,N_5972,N_5651);
and U6947 (N_6947,N_6362,N_5779);
xnor U6948 (N_6948,N_6193,N_6265);
and U6949 (N_6949,N_6393,N_6334);
nand U6950 (N_6950,N_5602,N_6378);
and U6951 (N_6951,N_6302,N_6249);
xor U6952 (N_6952,N_5924,N_6226);
xnor U6953 (N_6953,N_6383,N_6029);
xor U6954 (N_6954,N_6066,N_6017);
nor U6955 (N_6955,N_5990,N_5624);
and U6956 (N_6956,N_6068,N_5753);
nor U6957 (N_6957,N_6303,N_5999);
xnor U6958 (N_6958,N_5755,N_6220);
nor U6959 (N_6959,N_6235,N_5667);
or U6960 (N_6960,N_5851,N_6112);
nor U6961 (N_6961,N_5806,N_5712);
nor U6962 (N_6962,N_6178,N_5743);
nor U6963 (N_6963,N_5654,N_5744);
nand U6964 (N_6964,N_5810,N_6117);
or U6965 (N_6965,N_6130,N_6095);
nor U6966 (N_6966,N_6135,N_6372);
xnor U6967 (N_6967,N_5777,N_5869);
or U6968 (N_6968,N_5606,N_6251);
nand U6969 (N_6969,N_6269,N_5665);
nor U6970 (N_6970,N_5963,N_6337);
nand U6971 (N_6971,N_6156,N_5915);
nor U6972 (N_6972,N_6270,N_6145);
xor U6973 (N_6973,N_5790,N_6337);
and U6974 (N_6974,N_5671,N_5925);
nand U6975 (N_6975,N_6109,N_5774);
nand U6976 (N_6976,N_5746,N_6057);
and U6977 (N_6977,N_5706,N_6368);
xor U6978 (N_6978,N_6336,N_5743);
and U6979 (N_6979,N_5671,N_6378);
or U6980 (N_6980,N_5644,N_6036);
and U6981 (N_6981,N_5804,N_6228);
and U6982 (N_6982,N_6053,N_6300);
nand U6983 (N_6983,N_5614,N_6148);
xor U6984 (N_6984,N_5911,N_5641);
or U6985 (N_6985,N_6345,N_5860);
nand U6986 (N_6986,N_5887,N_6202);
or U6987 (N_6987,N_6242,N_6381);
or U6988 (N_6988,N_5782,N_5808);
nand U6989 (N_6989,N_6201,N_6389);
and U6990 (N_6990,N_5768,N_5688);
or U6991 (N_6991,N_5795,N_6305);
xnor U6992 (N_6992,N_5854,N_6310);
xnor U6993 (N_6993,N_5734,N_6143);
and U6994 (N_6994,N_5646,N_6282);
or U6995 (N_6995,N_6148,N_6038);
nor U6996 (N_6996,N_6297,N_6231);
or U6997 (N_6997,N_6265,N_6366);
nand U6998 (N_6998,N_6189,N_5998);
xor U6999 (N_6999,N_5823,N_5941);
and U7000 (N_7000,N_6267,N_5781);
or U7001 (N_7001,N_6270,N_6176);
or U7002 (N_7002,N_6304,N_5837);
nand U7003 (N_7003,N_6046,N_6169);
xnor U7004 (N_7004,N_6120,N_5667);
nand U7005 (N_7005,N_5972,N_6248);
nand U7006 (N_7006,N_5728,N_5620);
nand U7007 (N_7007,N_6028,N_5815);
and U7008 (N_7008,N_6346,N_5633);
nand U7009 (N_7009,N_6261,N_6395);
and U7010 (N_7010,N_6189,N_6146);
nand U7011 (N_7011,N_5964,N_5933);
nand U7012 (N_7012,N_5900,N_5791);
xor U7013 (N_7013,N_6377,N_5700);
and U7014 (N_7014,N_5756,N_6182);
nand U7015 (N_7015,N_5831,N_6028);
xnor U7016 (N_7016,N_6333,N_5620);
or U7017 (N_7017,N_5670,N_5736);
or U7018 (N_7018,N_6060,N_6337);
nor U7019 (N_7019,N_6259,N_5744);
nand U7020 (N_7020,N_5962,N_5700);
xnor U7021 (N_7021,N_6163,N_6211);
nand U7022 (N_7022,N_5884,N_5810);
or U7023 (N_7023,N_5626,N_6216);
and U7024 (N_7024,N_5757,N_5971);
and U7025 (N_7025,N_6382,N_6307);
xor U7026 (N_7026,N_6381,N_6052);
or U7027 (N_7027,N_6394,N_5874);
xnor U7028 (N_7028,N_6086,N_6242);
nand U7029 (N_7029,N_5953,N_5933);
or U7030 (N_7030,N_6370,N_5875);
or U7031 (N_7031,N_5623,N_6109);
xor U7032 (N_7032,N_5954,N_6118);
xnor U7033 (N_7033,N_5898,N_6160);
xnor U7034 (N_7034,N_6200,N_6040);
xnor U7035 (N_7035,N_6223,N_6345);
xor U7036 (N_7036,N_5754,N_6290);
or U7037 (N_7037,N_5737,N_6267);
nor U7038 (N_7038,N_5737,N_5852);
xnor U7039 (N_7039,N_5655,N_5731);
nor U7040 (N_7040,N_5607,N_6306);
nor U7041 (N_7041,N_6164,N_5771);
nor U7042 (N_7042,N_6155,N_6204);
and U7043 (N_7043,N_5743,N_6191);
xnor U7044 (N_7044,N_5974,N_6191);
nor U7045 (N_7045,N_6103,N_6167);
or U7046 (N_7046,N_5842,N_6345);
and U7047 (N_7047,N_5941,N_5963);
xnor U7048 (N_7048,N_5820,N_6159);
nor U7049 (N_7049,N_5698,N_5693);
or U7050 (N_7050,N_6141,N_5966);
and U7051 (N_7051,N_6347,N_5710);
or U7052 (N_7052,N_6185,N_6286);
or U7053 (N_7053,N_6129,N_6072);
nor U7054 (N_7054,N_6286,N_5736);
nand U7055 (N_7055,N_6161,N_5780);
nor U7056 (N_7056,N_5835,N_6098);
and U7057 (N_7057,N_5867,N_5790);
and U7058 (N_7058,N_5934,N_5969);
nor U7059 (N_7059,N_6204,N_6196);
nor U7060 (N_7060,N_5919,N_5892);
and U7061 (N_7061,N_5926,N_6135);
and U7062 (N_7062,N_6093,N_6226);
xor U7063 (N_7063,N_6125,N_6250);
xnor U7064 (N_7064,N_5954,N_6184);
nor U7065 (N_7065,N_5615,N_6330);
xnor U7066 (N_7066,N_6239,N_6391);
nand U7067 (N_7067,N_5655,N_6173);
and U7068 (N_7068,N_5992,N_5733);
or U7069 (N_7069,N_6249,N_5945);
or U7070 (N_7070,N_5680,N_5692);
xor U7071 (N_7071,N_6190,N_5736);
or U7072 (N_7072,N_6133,N_5730);
and U7073 (N_7073,N_5670,N_5852);
and U7074 (N_7074,N_5899,N_6163);
or U7075 (N_7075,N_6035,N_6161);
and U7076 (N_7076,N_5882,N_6168);
xor U7077 (N_7077,N_6020,N_6193);
and U7078 (N_7078,N_6013,N_5864);
nor U7079 (N_7079,N_5999,N_5725);
nor U7080 (N_7080,N_5930,N_6096);
xnor U7081 (N_7081,N_6215,N_6379);
xor U7082 (N_7082,N_6207,N_5845);
nor U7083 (N_7083,N_6280,N_5891);
xor U7084 (N_7084,N_6397,N_6031);
nor U7085 (N_7085,N_5761,N_5921);
nor U7086 (N_7086,N_6076,N_6093);
or U7087 (N_7087,N_6105,N_5801);
and U7088 (N_7088,N_5689,N_5841);
nor U7089 (N_7089,N_6265,N_5711);
nor U7090 (N_7090,N_5863,N_6176);
xor U7091 (N_7091,N_6217,N_6233);
xor U7092 (N_7092,N_6016,N_6310);
or U7093 (N_7093,N_5692,N_6236);
and U7094 (N_7094,N_6225,N_6082);
xor U7095 (N_7095,N_5842,N_5651);
nor U7096 (N_7096,N_6132,N_6339);
nor U7097 (N_7097,N_6283,N_5916);
or U7098 (N_7098,N_5647,N_5721);
or U7099 (N_7099,N_5792,N_6256);
nor U7100 (N_7100,N_5806,N_6141);
or U7101 (N_7101,N_5761,N_6280);
nor U7102 (N_7102,N_5926,N_6141);
xor U7103 (N_7103,N_6115,N_5666);
nand U7104 (N_7104,N_6094,N_6395);
or U7105 (N_7105,N_5624,N_6197);
nor U7106 (N_7106,N_5673,N_5956);
nand U7107 (N_7107,N_5743,N_6040);
and U7108 (N_7108,N_6122,N_5601);
and U7109 (N_7109,N_5919,N_5739);
nor U7110 (N_7110,N_6216,N_5755);
or U7111 (N_7111,N_5938,N_6141);
xnor U7112 (N_7112,N_6242,N_6033);
nand U7113 (N_7113,N_5863,N_6066);
nor U7114 (N_7114,N_5838,N_5650);
xnor U7115 (N_7115,N_5871,N_6280);
xnor U7116 (N_7116,N_5797,N_5928);
and U7117 (N_7117,N_5855,N_5717);
and U7118 (N_7118,N_5850,N_5800);
nand U7119 (N_7119,N_5849,N_5817);
xnor U7120 (N_7120,N_5773,N_5843);
or U7121 (N_7121,N_5914,N_5962);
nand U7122 (N_7122,N_6185,N_5686);
and U7123 (N_7123,N_6292,N_6138);
nor U7124 (N_7124,N_5902,N_6050);
xor U7125 (N_7125,N_6095,N_5941);
nor U7126 (N_7126,N_5603,N_6275);
and U7127 (N_7127,N_6134,N_5769);
or U7128 (N_7128,N_5901,N_5682);
or U7129 (N_7129,N_6192,N_6099);
xnor U7130 (N_7130,N_6050,N_5741);
nor U7131 (N_7131,N_5840,N_6289);
nand U7132 (N_7132,N_5681,N_6271);
and U7133 (N_7133,N_5962,N_5785);
and U7134 (N_7134,N_6108,N_5797);
and U7135 (N_7135,N_6120,N_5782);
and U7136 (N_7136,N_6327,N_5731);
or U7137 (N_7137,N_6066,N_6126);
or U7138 (N_7138,N_5963,N_5901);
or U7139 (N_7139,N_5758,N_5952);
nand U7140 (N_7140,N_5629,N_6101);
and U7141 (N_7141,N_5736,N_6091);
xnor U7142 (N_7142,N_6154,N_6255);
nand U7143 (N_7143,N_5862,N_6012);
nor U7144 (N_7144,N_6083,N_6230);
nand U7145 (N_7145,N_6047,N_6380);
and U7146 (N_7146,N_6314,N_5694);
xor U7147 (N_7147,N_5604,N_5946);
and U7148 (N_7148,N_5799,N_6084);
nor U7149 (N_7149,N_5840,N_6129);
xnor U7150 (N_7150,N_5793,N_6340);
or U7151 (N_7151,N_6078,N_6161);
xnor U7152 (N_7152,N_5864,N_5811);
nor U7153 (N_7153,N_5920,N_6058);
nor U7154 (N_7154,N_6266,N_6325);
nor U7155 (N_7155,N_5940,N_5864);
nor U7156 (N_7156,N_6029,N_5845);
nand U7157 (N_7157,N_5713,N_5809);
nand U7158 (N_7158,N_5758,N_6071);
xor U7159 (N_7159,N_5864,N_6377);
nand U7160 (N_7160,N_6335,N_6341);
nand U7161 (N_7161,N_5796,N_5801);
nand U7162 (N_7162,N_6171,N_6002);
or U7163 (N_7163,N_5827,N_6384);
nand U7164 (N_7164,N_6073,N_5871);
and U7165 (N_7165,N_6122,N_6025);
nand U7166 (N_7166,N_6336,N_6088);
xnor U7167 (N_7167,N_6252,N_5723);
or U7168 (N_7168,N_6109,N_6197);
nor U7169 (N_7169,N_5850,N_5994);
nor U7170 (N_7170,N_6325,N_6097);
xor U7171 (N_7171,N_6062,N_6122);
and U7172 (N_7172,N_5979,N_6057);
and U7173 (N_7173,N_5860,N_6131);
nor U7174 (N_7174,N_5969,N_5645);
or U7175 (N_7175,N_5807,N_6249);
or U7176 (N_7176,N_5758,N_6086);
xor U7177 (N_7177,N_5604,N_5831);
nor U7178 (N_7178,N_6264,N_6323);
nor U7179 (N_7179,N_6042,N_5624);
or U7180 (N_7180,N_5621,N_6173);
xnor U7181 (N_7181,N_6248,N_5783);
nand U7182 (N_7182,N_5965,N_6271);
nand U7183 (N_7183,N_5677,N_5917);
nand U7184 (N_7184,N_5770,N_5993);
and U7185 (N_7185,N_6395,N_6101);
xnor U7186 (N_7186,N_6234,N_5823);
and U7187 (N_7187,N_5614,N_5924);
nand U7188 (N_7188,N_5798,N_5933);
or U7189 (N_7189,N_6243,N_6240);
or U7190 (N_7190,N_6250,N_6046);
nand U7191 (N_7191,N_6392,N_6281);
and U7192 (N_7192,N_6164,N_6010);
or U7193 (N_7193,N_6390,N_5764);
and U7194 (N_7194,N_6300,N_6174);
or U7195 (N_7195,N_6192,N_6142);
xnor U7196 (N_7196,N_6126,N_6358);
nor U7197 (N_7197,N_6260,N_5827);
nand U7198 (N_7198,N_5899,N_6127);
nor U7199 (N_7199,N_5714,N_5616);
nor U7200 (N_7200,N_6712,N_7176);
nand U7201 (N_7201,N_6769,N_6409);
xnor U7202 (N_7202,N_6724,N_6721);
xor U7203 (N_7203,N_6833,N_6420);
nand U7204 (N_7204,N_6454,N_6857);
and U7205 (N_7205,N_7051,N_6498);
and U7206 (N_7206,N_6475,N_6743);
and U7207 (N_7207,N_6938,N_6914);
or U7208 (N_7208,N_6937,N_6872);
nand U7209 (N_7209,N_6876,N_7171);
and U7210 (N_7210,N_6535,N_7187);
nor U7211 (N_7211,N_6871,N_7159);
or U7212 (N_7212,N_6696,N_6494);
nor U7213 (N_7213,N_6901,N_6666);
nor U7214 (N_7214,N_6843,N_6840);
nor U7215 (N_7215,N_6439,N_6661);
nor U7216 (N_7216,N_7118,N_6802);
xor U7217 (N_7217,N_6610,N_7195);
nand U7218 (N_7218,N_7029,N_7158);
nand U7219 (N_7219,N_6408,N_7155);
nor U7220 (N_7220,N_7149,N_6601);
xor U7221 (N_7221,N_6456,N_6824);
nor U7222 (N_7222,N_7121,N_6866);
or U7223 (N_7223,N_6903,N_7024);
nor U7224 (N_7224,N_6782,N_6413);
nor U7225 (N_7225,N_6839,N_7168);
nand U7226 (N_7226,N_6697,N_6997);
xnor U7227 (N_7227,N_7143,N_6734);
nor U7228 (N_7228,N_6879,N_6440);
nor U7229 (N_7229,N_6629,N_6924);
or U7230 (N_7230,N_7002,N_7045);
xnor U7231 (N_7231,N_6943,N_6583);
nand U7232 (N_7232,N_6771,N_6756);
or U7233 (N_7233,N_7095,N_6928);
nor U7234 (N_7234,N_6720,N_7164);
nor U7235 (N_7235,N_6676,N_6902);
xor U7236 (N_7236,N_6524,N_6741);
nand U7237 (N_7237,N_6457,N_6599);
or U7238 (N_7238,N_6591,N_6622);
nand U7239 (N_7239,N_6795,N_7181);
or U7240 (N_7240,N_6774,N_7009);
and U7241 (N_7241,N_6500,N_6966);
nand U7242 (N_7242,N_6698,N_7094);
or U7243 (N_7243,N_6639,N_6617);
nor U7244 (N_7244,N_6953,N_6746);
xnor U7245 (N_7245,N_6681,N_6468);
and U7246 (N_7246,N_6964,N_6547);
nor U7247 (N_7247,N_6702,N_6611);
and U7248 (N_7248,N_6765,N_6781);
nand U7249 (N_7249,N_6506,N_6404);
nor U7250 (N_7250,N_6899,N_6921);
xor U7251 (N_7251,N_6814,N_6633);
and U7252 (N_7252,N_6554,N_6642);
xnor U7253 (N_7253,N_7132,N_7136);
nand U7254 (N_7254,N_7092,N_6910);
nand U7255 (N_7255,N_6608,N_6678);
nand U7256 (N_7256,N_6729,N_6564);
and U7257 (N_7257,N_6527,N_6847);
xor U7258 (N_7258,N_7161,N_6799);
nand U7259 (N_7259,N_7062,N_6888);
nand U7260 (N_7260,N_6869,N_6770);
and U7261 (N_7261,N_6897,N_6875);
or U7262 (N_7262,N_6913,N_6455);
nor U7263 (N_7263,N_6425,N_7022);
nor U7264 (N_7264,N_7070,N_7173);
xor U7265 (N_7265,N_6415,N_6733);
nor U7266 (N_7266,N_6801,N_7055);
and U7267 (N_7267,N_6448,N_6882);
or U7268 (N_7268,N_7080,N_6406);
and U7269 (N_7269,N_6537,N_7056);
xor U7270 (N_7270,N_6837,N_6859);
nand U7271 (N_7271,N_6740,N_7157);
nand U7272 (N_7272,N_6985,N_6571);
or U7273 (N_7273,N_6735,N_7113);
or U7274 (N_7274,N_6932,N_6447);
and U7275 (N_7275,N_6446,N_6464);
xnor U7276 (N_7276,N_6727,N_6512);
nand U7277 (N_7277,N_6556,N_6715);
xor U7278 (N_7278,N_6626,N_6686);
and U7279 (N_7279,N_6555,N_6958);
and U7280 (N_7280,N_6768,N_7172);
or U7281 (N_7281,N_7154,N_6585);
and U7282 (N_7282,N_6878,N_7166);
or U7283 (N_7283,N_6852,N_6905);
or U7284 (N_7284,N_6714,N_6432);
or U7285 (N_7285,N_7048,N_7046);
or U7286 (N_7286,N_6424,N_7099);
xnor U7287 (N_7287,N_7003,N_6561);
or U7288 (N_7288,N_7035,N_6788);
or U7289 (N_7289,N_6907,N_7087);
or U7290 (N_7290,N_6660,N_6429);
or U7291 (N_7291,N_7047,N_6865);
or U7292 (N_7292,N_6808,N_7190);
or U7293 (N_7293,N_6423,N_6652);
and U7294 (N_7294,N_6753,N_6792);
nand U7295 (N_7295,N_7042,N_6478);
nor U7296 (N_7296,N_7145,N_6559);
nor U7297 (N_7297,N_7067,N_6541);
nor U7298 (N_7298,N_6656,N_6900);
nand U7299 (N_7299,N_7138,N_6606);
or U7300 (N_7300,N_6908,N_6552);
xnor U7301 (N_7301,N_7030,N_6476);
or U7302 (N_7302,N_6594,N_6936);
xnor U7303 (N_7303,N_7069,N_7081);
nor U7304 (N_7304,N_6526,N_6543);
or U7305 (N_7305,N_6993,N_6628);
nor U7306 (N_7306,N_6465,N_6728);
and U7307 (N_7307,N_6811,N_7130);
xnor U7308 (N_7308,N_6980,N_6680);
xnor U7309 (N_7309,N_6864,N_6893);
nand U7310 (N_7310,N_7000,N_6722);
and U7311 (N_7311,N_6472,N_6523);
nand U7312 (N_7312,N_6576,N_6574);
or U7313 (N_7313,N_6977,N_6605);
nand U7314 (N_7314,N_7065,N_7185);
nor U7315 (N_7315,N_6671,N_6744);
and U7316 (N_7316,N_6402,N_6563);
or U7317 (N_7317,N_6813,N_6780);
and U7318 (N_7318,N_7049,N_6492);
or U7319 (N_7319,N_7119,N_6818);
nor U7320 (N_7320,N_6663,N_6826);
nand U7321 (N_7321,N_6590,N_6776);
and U7322 (N_7322,N_6688,N_6950);
and U7323 (N_7323,N_7058,N_6403);
xor U7324 (N_7324,N_7020,N_6533);
xor U7325 (N_7325,N_6568,N_6850);
nor U7326 (N_7326,N_7129,N_6796);
and U7327 (N_7327,N_6613,N_6436);
xor U7328 (N_7328,N_7085,N_6920);
xor U7329 (N_7329,N_6961,N_6469);
nand U7330 (N_7330,N_7091,N_6787);
or U7331 (N_7331,N_6790,N_6760);
or U7332 (N_7332,N_6548,N_7192);
or U7333 (N_7333,N_7004,N_6705);
nor U7334 (N_7334,N_6948,N_6607);
and U7335 (N_7335,N_6895,N_6834);
and U7336 (N_7336,N_6942,N_6630);
nand U7337 (N_7337,N_7139,N_6484);
and U7338 (N_7338,N_6677,N_6983);
xor U7339 (N_7339,N_6836,N_6965);
xnor U7340 (N_7340,N_6445,N_6603);
and U7341 (N_7341,N_6699,N_6586);
nand U7342 (N_7342,N_7117,N_6994);
and U7343 (N_7343,N_7013,N_7183);
nand U7344 (N_7344,N_6416,N_6690);
nand U7345 (N_7345,N_6502,N_6772);
xnor U7346 (N_7346,N_6507,N_6957);
nand U7347 (N_7347,N_7196,N_6679);
xnor U7348 (N_7348,N_6670,N_6479);
and U7349 (N_7349,N_7034,N_7019);
and U7350 (N_7350,N_7112,N_7131);
and U7351 (N_7351,N_7014,N_6732);
nand U7352 (N_7352,N_6870,N_6967);
nand U7353 (N_7353,N_6867,N_6549);
and U7354 (N_7354,N_6922,N_6545);
nand U7355 (N_7355,N_6810,N_7137);
nand U7356 (N_7356,N_6856,N_6815);
nor U7357 (N_7357,N_6604,N_7197);
and U7358 (N_7358,N_6933,N_6831);
nand U7359 (N_7359,N_7005,N_6832);
xor U7360 (N_7360,N_6968,N_6877);
xnor U7361 (N_7361,N_6410,N_7147);
and U7362 (N_7362,N_6805,N_6481);
xor U7363 (N_7363,N_6505,N_6520);
or U7364 (N_7364,N_7169,N_6466);
nand U7365 (N_7365,N_6971,N_6598);
xor U7366 (N_7366,N_6650,N_6767);
nor U7367 (N_7367,N_6575,N_6725);
nor U7368 (N_7368,N_6946,N_6995);
nand U7369 (N_7369,N_7098,N_6917);
xor U7370 (N_7370,N_6615,N_7180);
or U7371 (N_7371,N_7152,N_6491);
and U7372 (N_7372,N_7036,N_7107);
xor U7373 (N_7373,N_6822,N_6437);
or U7374 (N_7374,N_7186,N_6657);
nor U7375 (N_7375,N_6509,N_6996);
and U7376 (N_7376,N_6861,N_6855);
xor U7377 (N_7377,N_7052,N_6742);
xor U7378 (N_7378,N_6989,N_6817);
xor U7379 (N_7379,N_6962,N_6894);
nand U7380 (N_7380,N_6625,N_7144);
and U7381 (N_7381,N_6664,N_6739);
or U7382 (N_7382,N_6749,N_6773);
and U7383 (N_7383,N_6981,N_6929);
nand U7384 (N_7384,N_6751,N_7068);
nand U7385 (N_7385,N_6499,N_6578);
nor U7386 (N_7386,N_6915,N_7106);
xor U7387 (N_7387,N_6627,N_6421);
xor U7388 (N_7388,N_6777,N_6784);
nor U7389 (N_7389,N_6597,N_7165);
xnor U7390 (N_7390,N_6700,N_6779);
xor U7391 (N_7391,N_6763,N_6898);
nand U7392 (N_7392,N_6819,N_6667);
and U7393 (N_7393,N_6930,N_6460);
nor U7394 (N_7394,N_6992,N_6659);
xnor U7395 (N_7395,N_6412,N_6546);
or U7396 (N_7396,N_7015,N_6544);
or U7397 (N_7397,N_7148,N_7153);
nor U7398 (N_7398,N_6430,N_6600);
nor U7399 (N_7399,N_7054,N_6584);
and U7400 (N_7400,N_6827,N_6495);
xor U7401 (N_7401,N_6703,N_6534);
and U7402 (N_7402,N_6912,N_6593);
or U7403 (N_7403,N_6828,N_6419);
xnor U7404 (N_7404,N_7075,N_6637);
or U7405 (N_7405,N_6634,N_6441);
and U7406 (N_7406,N_6518,N_6785);
nor U7407 (N_7407,N_7059,N_6969);
xnor U7408 (N_7408,N_6638,N_6462);
nand U7409 (N_7409,N_6612,N_7007);
or U7410 (N_7410,N_6874,N_7011);
xor U7411 (N_7411,N_6496,N_6434);
nor U7412 (N_7412,N_6467,N_6528);
nor U7413 (N_7413,N_6538,N_6890);
xor U7414 (N_7414,N_6803,N_6820);
and U7415 (N_7415,N_7043,N_6991);
xnor U7416 (N_7416,N_6884,N_6658);
nand U7417 (N_7417,N_6738,N_7109);
or U7418 (N_7418,N_6689,N_7199);
xor U7419 (N_7419,N_7066,N_6687);
nand U7420 (N_7420,N_6504,N_6845);
and U7421 (N_7421,N_6934,N_6775);
xor U7422 (N_7422,N_7041,N_7124);
xnor U7423 (N_7423,N_6816,N_7167);
and U7424 (N_7424,N_6668,N_6654);
xnor U7425 (N_7425,N_6405,N_6759);
xnor U7426 (N_7426,N_6530,N_6949);
nor U7427 (N_7427,N_6830,N_7017);
and U7428 (N_7428,N_6411,N_6842);
nor U7429 (N_7429,N_7110,N_6999);
xor U7430 (N_7430,N_6477,N_6955);
and U7431 (N_7431,N_6672,N_6806);
or U7432 (N_7432,N_6595,N_6669);
and U7433 (N_7433,N_6570,N_6487);
nor U7434 (N_7434,N_6987,N_6517);
nor U7435 (N_7435,N_6614,N_6510);
or U7436 (N_7436,N_7134,N_6655);
nor U7437 (N_7437,N_6974,N_6453);
or U7438 (N_7438,N_6461,N_6553);
and U7439 (N_7439,N_6757,N_6794);
xnor U7440 (N_7440,N_6588,N_6452);
xnor U7441 (N_7441,N_6522,N_6880);
nor U7442 (N_7442,N_6508,N_6926);
xnor U7443 (N_7443,N_6809,N_6947);
nor U7444 (N_7444,N_6736,N_6674);
xor U7445 (N_7445,N_6560,N_6645);
nand U7446 (N_7446,N_6501,N_6986);
nor U7447 (N_7447,N_6973,N_6963);
and U7448 (N_7448,N_6719,N_6918);
and U7449 (N_7449,N_7053,N_6400);
nand U7450 (N_7450,N_6786,N_6750);
and U7451 (N_7451,N_6998,N_6835);
or U7452 (N_7452,N_6887,N_7188);
xnor U7453 (N_7453,N_7097,N_6592);
or U7454 (N_7454,N_6923,N_6407);
nand U7455 (N_7455,N_6952,N_7115);
or U7456 (N_7456,N_6730,N_6891);
xnor U7457 (N_7457,N_7101,N_6916);
nor U7458 (N_7458,N_7064,N_6511);
nor U7459 (N_7459,N_6644,N_6927);
nand U7460 (N_7460,N_6401,N_6791);
nor U7461 (N_7461,N_6521,N_6566);
and U7462 (N_7462,N_6470,N_6704);
xnor U7463 (N_7463,N_6532,N_6976);
nor U7464 (N_7464,N_6482,N_7120);
and U7465 (N_7465,N_6619,N_6450);
or U7466 (N_7466,N_6431,N_6685);
or U7467 (N_7467,N_6940,N_6881);
nand U7468 (N_7468,N_7150,N_6474);
nand U7469 (N_7469,N_6463,N_7104);
nor U7470 (N_7470,N_6648,N_6990);
and U7471 (N_7471,N_6959,N_6683);
and U7472 (N_7472,N_6709,N_6550);
and U7473 (N_7473,N_7074,N_7076);
nor U7474 (N_7474,N_6649,N_6418);
or U7475 (N_7475,N_7026,N_6539);
xnor U7476 (N_7476,N_6641,N_6444);
nand U7477 (N_7477,N_6825,N_7037);
or U7478 (N_7478,N_7142,N_6737);
and U7479 (N_7479,N_6896,N_6904);
and U7480 (N_7480,N_6778,N_6620);
nor U7481 (N_7481,N_6789,N_7111);
and U7482 (N_7482,N_7105,N_6931);
xor U7483 (N_7483,N_6647,N_6417);
xnor U7484 (N_7484,N_7008,N_6486);
nand U7485 (N_7485,N_6414,N_6982);
and U7486 (N_7486,N_6713,N_7170);
or U7487 (N_7487,N_6567,N_6525);
nor U7488 (N_7488,N_7012,N_6988);
and U7489 (N_7489,N_6941,N_7140);
nor U7490 (N_7490,N_7103,N_6565);
xnor U7491 (N_7491,N_6675,N_6844);
nand U7492 (N_7492,N_6752,N_7032);
or U7493 (N_7493,N_7084,N_6562);
xnor U7494 (N_7494,N_6694,N_7040);
nor U7495 (N_7495,N_7108,N_7063);
or U7496 (N_7496,N_7090,N_6692);
xnor U7497 (N_7497,N_6489,N_6673);
xnor U7498 (N_7498,N_7060,N_6651);
xor U7499 (N_7499,N_6939,N_7156);
or U7500 (N_7500,N_7086,N_6662);
nand U7501 (N_7501,N_6761,N_6572);
or U7502 (N_7502,N_6783,N_6954);
or U7503 (N_7503,N_7198,N_6862);
nor U7504 (N_7504,N_6580,N_6854);
or U7505 (N_7505,N_6889,N_6793);
and U7506 (N_7506,N_6438,N_6762);
xor U7507 (N_7507,N_6945,N_6459);
nor U7508 (N_7508,N_7141,N_6707);
nand U7509 (N_7509,N_7163,N_7038);
and U7510 (N_7510,N_7071,N_6573);
or U7511 (N_7511,N_7096,N_6427);
nand U7512 (N_7512,N_6706,N_7078);
nand U7513 (N_7513,N_7114,N_6800);
nor U7514 (N_7514,N_7057,N_6823);
or U7515 (N_7515,N_6868,N_6540);
or U7516 (N_7516,N_7151,N_6755);
nand U7517 (N_7517,N_7044,N_6925);
or U7518 (N_7518,N_6911,N_6691);
xnor U7519 (N_7519,N_6616,N_6892);
nor U7520 (N_7520,N_6551,N_6860);
or U7521 (N_7521,N_6458,N_7050);
or U7522 (N_7522,N_6848,N_6646);
nand U7523 (N_7523,N_6631,N_7073);
nand U7524 (N_7524,N_6978,N_6636);
nor U7525 (N_7525,N_6529,N_6851);
nand U7526 (N_7526,N_7184,N_7178);
and U7527 (N_7527,N_6748,N_6754);
nand U7528 (N_7528,N_7128,N_6718);
nor U7529 (N_7529,N_6701,N_6602);
xor U7530 (N_7530,N_6726,N_6853);
and U7531 (N_7531,N_6632,N_6684);
or U7532 (N_7532,N_7189,N_7116);
and U7533 (N_7533,N_6536,N_7122);
or U7534 (N_7534,N_6873,N_6695);
nor U7535 (N_7535,N_6483,N_6886);
xnor U7536 (N_7536,N_7033,N_6587);
xor U7537 (N_7537,N_6863,N_6635);
nand U7538 (N_7538,N_7175,N_7016);
xor U7539 (N_7539,N_6480,N_6451);
xnor U7540 (N_7540,N_6531,N_6764);
or U7541 (N_7541,N_6621,N_7179);
and U7542 (N_7542,N_6807,N_7088);
nor U7543 (N_7543,N_6731,N_7162);
xor U7544 (N_7544,N_6618,N_7127);
nor U7545 (N_7545,N_6970,N_6935);
nand U7546 (N_7546,N_6577,N_7093);
nor U7547 (N_7547,N_6558,N_7102);
and U7548 (N_7548,N_6426,N_6443);
or U7549 (N_7549,N_6710,N_6665);
xor U7550 (N_7550,N_6693,N_7077);
nor U7551 (N_7551,N_7135,N_7133);
nand U7552 (N_7552,N_7194,N_7182);
nand U7553 (N_7553,N_7082,N_6919);
and U7554 (N_7554,N_6435,N_6488);
xor U7555 (N_7555,N_6471,N_6643);
xor U7556 (N_7556,N_6589,N_6542);
xor U7557 (N_7557,N_6960,N_6849);
nor U7558 (N_7558,N_7027,N_6797);
and U7559 (N_7559,N_6944,N_7079);
or U7560 (N_7560,N_6747,N_6979);
nor U7561 (N_7561,N_7039,N_6838);
nand U7562 (N_7562,N_7023,N_6442);
nor U7563 (N_7563,N_7177,N_6490);
or U7564 (N_7564,N_6829,N_6708);
and U7565 (N_7565,N_6515,N_7160);
xnor U7566 (N_7566,N_6711,N_6579);
and U7567 (N_7567,N_6581,N_6582);
xnor U7568 (N_7568,N_7001,N_7031);
nor U7569 (N_7569,N_6846,N_7100);
and U7570 (N_7570,N_6841,N_7061);
and U7571 (N_7571,N_6433,N_7018);
or U7572 (N_7572,N_7123,N_6906);
nand U7573 (N_7573,N_6493,N_6503);
xor U7574 (N_7574,N_6513,N_6653);
nor U7575 (N_7575,N_6975,N_6449);
and U7576 (N_7576,N_7126,N_6717);
nand U7577 (N_7577,N_7083,N_6609);
and U7578 (N_7578,N_6804,N_6745);
or U7579 (N_7579,N_7028,N_6519);
or U7580 (N_7580,N_7025,N_6516);
nand U7581 (N_7581,N_6766,N_7174);
or U7582 (N_7582,N_6758,N_6972);
nand U7583 (N_7583,N_6909,N_6885);
xor U7584 (N_7584,N_7146,N_6514);
and U7585 (N_7585,N_6623,N_7010);
nand U7586 (N_7586,N_6812,N_6428);
nand U7587 (N_7587,N_6485,N_7072);
and U7588 (N_7588,N_6497,N_7089);
xnor U7589 (N_7589,N_6821,N_6956);
or U7590 (N_7590,N_6984,N_6716);
xor U7591 (N_7591,N_6473,N_7191);
nand U7592 (N_7592,N_7193,N_6596);
nand U7593 (N_7593,N_6569,N_6640);
nor U7594 (N_7594,N_6798,N_6682);
nor U7595 (N_7595,N_6858,N_7021);
nand U7596 (N_7596,N_6723,N_6951);
nand U7597 (N_7597,N_6422,N_6883);
xnor U7598 (N_7598,N_7006,N_6624);
nor U7599 (N_7599,N_6557,N_7125);
or U7600 (N_7600,N_6796,N_6737);
xor U7601 (N_7601,N_6559,N_6423);
nor U7602 (N_7602,N_6923,N_6561);
nor U7603 (N_7603,N_6762,N_6982);
and U7604 (N_7604,N_6653,N_6752);
nand U7605 (N_7605,N_6767,N_7056);
nor U7606 (N_7606,N_6674,N_6854);
xnor U7607 (N_7607,N_6953,N_7071);
nor U7608 (N_7608,N_6917,N_6585);
xnor U7609 (N_7609,N_6691,N_6552);
and U7610 (N_7610,N_7067,N_7040);
and U7611 (N_7611,N_6707,N_7014);
or U7612 (N_7612,N_6591,N_6431);
and U7613 (N_7613,N_7144,N_7059);
or U7614 (N_7614,N_6558,N_6977);
nor U7615 (N_7615,N_6748,N_6678);
or U7616 (N_7616,N_6839,N_7090);
nand U7617 (N_7617,N_6955,N_6588);
nand U7618 (N_7618,N_6847,N_7103);
and U7619 (N_7619,N_7187,N_7193);
nor U7620 (N_7620,N_6837,N_6429);
nand U7621 (N_7621,N_6954,N_7007);
xnor U7622 (N_7622,N_6762,N_6433);
xnor U7623 (N_7623,N_6567,N_6929);
nor U7624 (N_7624,N_6622,N_6689);
or U7625 (N_7625,N_6400,N_6648);
nand U7626 (N_7626,N_6743,N_6799);
nor U7627 (N_7627,N_6718,N_6427);
xnor U7628 (N_7628,N_6503,N_7005);
nor U7629 (N_7629,N_7076,N_7014);
xor U7630 (N_7630,N_6944,N_6925);
xor U7631 (N_7631,N_7156,N_6721);
nand U7632 (N_7632,N_6428,N_6454);
nor U7633 (N_7633,N_7152,N_7169);
xor U7634 (N_7634,N_7002,N_6415);
nor U7635 (N_7635,N_6420,N_6461);
nor U7636 (N_7636,N_7066,N_6917);
nand U7637 (N_7637,N_7147,N_6599);
or U7638 (N_7638,N_6808,N_6813);
nand U7639 (N_7639,N_7024,N_6694);
nand U7640 (N_7640,N_6826,N_6424);
xor U7641 (N_7641,N_7077,N_7148);
xor U7642 (N_7642,N_7188,N_6670);
xor U7643 (N_7643,N_6967,N_6546);
and U7644 (N_7644,N_6491,N_6745);
xnor U7645 (N_7645,N_6680,N_6414);
and U7646 (N_7646,N_6988,N_6657);
or U7647 (N_7647,N_6509,N_7192);
or U7648 (N_7648,N_6550,N_6973);
and U7649 (N_7649,N_6553,N_6910);
xnor U7650 (N_7650,N_6675,N_6960);
and U7651 (N_7651,N_7077,N_6598);
xnor U7652 (N_7652,N_6476,N_6493);
nand U7653 (N_7653,N_6890,N_6859);
nand U7654 (N_7654,N_6439,N_6465);
nand U7655 (N_7655,N_7020,N_7135);
nor U7656 (N_7656,N_7064,N_6919);
or U7657 (N_7657,N_6974,N_6464);
or U7658 (N_7658,N_7155,N_6972);
and U7659 (N_7659,N_7195,N_7066);
or U7660 (N_7660,N_7009,N_6657);
nand U7661 (N_7661,N_7151,N_6842);
and U7662 (N_7662,N_6922,N_6763);
and U7663 (N_7663,N_6820,N_6511);
nor U7664 (N_7664,N_6406,N_6506);
nand U7665 (N_7665,N_6818,N_6522);
nand U7666 (N_7666,N_6557,N_7060);
xor U7667 (N_7667,N_6646,N_6419);
nor U7668 (N_7668,N_6763,N_7093);
or U7669 (N_7669,N_7064,N_7129);
nand U7670 (N_7670,N_6865,N_6674);
and U7671 (N_7671,N_7089,N_7155);
and U7672 (N_7672,N_7136,N_6673);
nand U7673 (N_7673,N_6950,N_6549);
or U7674 (N_7674,N_7195,N_6691);
nor U7675 (N_7675,N_6466,N_6878);
and U7676 (N_7676,N_7147,N_6614);
or U7677 (N_7677,N_6844,N_6753);
nand U7678 (N_7678,N_6479,N_6757);
nor U7679 (N_7679,N_6652,N_6811);
or U7680 (N_7680,N_7024,N_6701);
nand U7681 (N_7681,N_6833,N_6478);
nand U7682 (N_7682,N_6511,N_6555);
or U7683 (N_7683,N_6845,N_7052);
and U7684 (N_7684,N_6849,N_6906);
or U7685 (N_7685,N_6782,N_6604);
or U7686 (N_7686,N_6411,N_6464);
xor U7687 (N_7687,N_6508,N_6681);
nor U7688 (N_7688,N_7186,N_6558);
xor U7689 (N_7689,N_6488,N_7026);
or U7690 (N_7690,N_7006,N_7153);
nand U7691 (N_7691,N_6844,N_6967);
nand U7692 (N_7692,N_6554,N_6686);
nand U7693 (N_7693,N_7013,N_6870);
or U7694 (N_7694,N_6511,N_6651);
and U7695 (N_7695,N_6628,N_7112);
and U7696 (N_7696,N_6809,N_6523);
xor U7697 (N_7697,N_6515,N_6420);
xor U7698 (N_7698,N_6974,N_6919);
nor U7699 (N_7699,N_7107,N_6415);
or U7700 (N_7700,N_6586,N_7193);
and U7701 (N_7701,N_6575,N_7001);
xnor U7702 (N_7702,N_6629,N_6525);
nor U7703 (N_7703,N_6703,N_6430);
nand U7704 (N_7704,N_6712,N_7025);
xor U7705 (N_7705,N_6839,N_6617);
or U7706 (N_7706,N_6732,N_6424);
xor U7707 (N_7707,N_6663,N_6574);
or U7708 (N_7708,N_6667,N_6579);
nand U7709 (N_7709,N_7005,N_7074);
and U7710 (N_7710,N_7067,N_6865);
nand U7711 (N_7711,N_6884,N_6456);
nor U7712 (N_7712,N_7057,N_7019);
nand U7713 (N_7713,N_7125,N_6447);
xnor U7714 (N_7714,N_6801,N_6794);
or U7715 (N_7715,N_6664,N_6565);
nand U7716 (N_7716,N_6618,N_6582);
xor U7717 (N_7717,N_6776,N_6646);
or U7718 (N_7718,N_6548,N_7155);
or U7719 (N_7719,N_6783,N_6465);
nor U7720 (N_7720,N_6649,N_6468);
xnor U7721 (N_7721,N_6558,N_6860);
nand U7722 (N_7722,N_6882,N_6732);
nor U7723 (N_7723,N_6459,N_7115);
or U7724 (N_7724,N_7191,N_6899);
or U7725 (N_7725,N_6590,N_6850);
xnor U7726 (N_7726,N_6635,N_6933);
xor U7727 (N_7727,N_7181,N_6921);
nand U7728 (N_7728,N_7157,N_6456);
or U7729 (N_7729,N_6930,N_7131);
nand U7730 (N_7730,N_6763,N_6650);
or U7731 (N_7731,N_6437,N_7119);
and U7732 (N_7732,N_7069,N_6548);
or U7733 (N_7733,N_6414,N_6884);
nand U7734 (N_7734,N_6412,N_6737);
and U7735 (N_7735,N_7052,N_6585);
or U7736 (N_7736,N_6471,N_6561);
or U7737 (N_7737,N_7126,N_6768);
and U7738 (N_7738,N_6794,N_6864);
xor U7739 (N_7739,N_7058,N_6412);
nor U7740 (N_7740,N_6864,N_6704);
nand U7741 (N_7741,N_6742,N_7069);
nand U7742 (N_7742,N_7118,N_7005);
or U7743 (N_7743,N_7189,N_6600);
xnor U7744 (N_7744,N_6621,N_6714);
xnor U7745 (N_7745,N_7056,N_6586);
and U7746 (N_7746,N_7194,N_6937);
nand U7747 (N_7747,N_6437,N_6542);
and U7748 (N_7748,N_6479,N_6822);
and U7749 (N_7749,N_6510,N_6418);
xnor U7750 (N_7750,N_6756,N_6437);
and U7751 (N_7751,N_7141,N_7116);
nand U7752 (N_7752,N_6493,N_7094);
and U7753 (N_7753,N_6511,N_6608);
xor U7754 (N_7754,N_6548,N_6438);
or U7755 (N_7755,N_7043,N_7047);
and U7756 (N_7756,N_7198,N_7176);
nand U7757 (N_7757,N_6498,N_7160);
and U7758 (N_7758,N_6628,N_7137);
or U7759 (N_7759,N_6780,N_6940);
or U7760 (N_7760,N_6564,N_7130);
xnor U7761 (N_7761,N_6455,N_7033);
nand U7762 (N_7762,N_6434,N_7186);
nand U7763 (N_7763,N_6751,N_6819);
and U7764 (N_7764,N_6580,N_6868);
nor U7765 (N_7765,N_6721,N_6467);
or U7766 (N_7766,N_6974,N_6746);
and U7767 (N_7767,N_6702,N_6501);
and U7768 (N_7768,N_6946,N_6953);
xnor U7769 (N_7769,N_6976,N_7129);
xnor U7770 (N_7770,N_6800,N_6736);
nor U7771 (N_7771,N_6955,N_7128);
nor U7772 (N_7772,N_7047,N_6832);
nor U7773 (N_7773,N_6583,N_6999);
nand U7774 (N_7774,N_7031,N_6524);
and U7775 (N_7775,N_6997,N_6777);
nand U7776 (N_7776,N_6965,N_6967);
xor U7777 (N_7777,N_7020,N_7134);
xor U7778 (N_7778,N_6880,N_6547);
or U7779 (N_7779,N_6831,N_6692);
or U7780 (N_7780,N_7051,N_6974);
nor U7781 (N_7781,N_6870,N_6957);
nand U7782 (N_7782,N_7076,N_6851);
or U7783 (N_7783,N_7140,N_6869);
or U7784 (N_7784,N_6586,N_6415);
or U7785 (N_7785,N_7002,N_6714);
and U7786 (N_7786,N_6402,N_6650);
xnor U7787 (N_7787,N_6819,N_6783);
nand U7788 (N_7788,N_7042,N_6705);
xor U7789 (N_7789,N_6727,N_6714);
and U7790 (N_7790,N_6802,N_7195);
nor U7791 (N_7791,N_6909,N_7033);
and U7792 (N_7792,N_6875,N_6980);
nand U7793 (N_7793,N_6593,N_6884);
nor U7794 (N_7794,N_6914,N_7183);
xor U7795 (N_7795,N_7159,N_6607);
or U7796 (N_7796,N_7138,N_6402);
nand U7797 (N_7797,N_6927,N_6698);
nor U7798 (N_7798,N_6846,N_7147);
nor U7799 (N_7799,N_6481,N_6473);
or U7800 (N_7800,N_6990,N_6947);
nand U7801 (N_7801,N_6531,N_6453);
nor U7802 (N_7802,N_7110,N_7065);
or U7803 (N_7803,N_7172,N_6884);
nand U7804 (N_7804,N_6724,N_6938);
xor U7805 (N_7805,N_7151,N_6997);
xor U7806 (N_7806,N_6585,N_6842);
nor U7807 (N_7807,N_6937,N_7156);
or U7808 (N_7808,N_7199,N_7179);
nand U7809 (N_7809,N_6748,N_7107);
and U7810 (N_7810,N_6764,N_6702);
nor U7811 (N_7811,N_6614,N_6498);
nor U7812 (N_7812,N_7089,N_6713);
nor U7813 (N_7813,N_6481,N_6438);
or U7814 (N_7814,N_7139,N_7120);
and U7815 (N_7815,N_7086,N_6932);
and U7816 (N_7816,N_7005,N_6495);
nor U7817 (N_7817,N_6518,N_6519);
nor U7818 (N_7818,N_6849,N_7113);
nor U7819 (N_7819,N_7066,N_7006);
nand U7820 (N_7820,N_6460,N_6634);
and U7821 (N_7821,N_7132,N_7058);
or U7822 (N_7822,N_6532,N_7100);
or U7823 (N_7823,N_6899,N_7134);
and U7824 (N_7824,N_6944,N_6656);
nand U7825 (N_7825,N_6426,N_6495);
nand U7826 (N_7826,N_6825,N_6787);
xnor U7827 (N_7827,N_6672,N_6737);
and U7828 (N_7828,N_6874,N_6741);
and U7829 (N_7829,N_6780,N_7062);
nor U7830 (N_7830,N_6828,N_7002);
nor U7831 (N_7831,N_6637,N_7035);
nor U7832 (N_7832,N_6585,N_6788);
or U7833 (N_7833,N_6761,N_6817);
nand U7834 (N_7834,N_7023,N_6466);
and U7835 (N_7835,N_6915,N_6736);
or U7836 (N_7836,N_6744,N_6426);
nor U7837 (N_7837,N_7081,N_6431);
and U7838 (N_7838,N_6932,N_6583);
nand U7839 (N_7839,N_6410,N_6719);
nand U7840 (N_7840,N_7194,N_6552);
and U7841 (N_7841,N_6770,N_6773);
and U7842 (N_7842,N_6966,N_6773);
or U7843 (N_7843,N_6603,N_7126);
nor U7844 (N_7844,N_7011,N_6435);
xnor U7845 (N_7845,N_6561,N_6625);
and U7846 (N_7846,N_7100,N_7097);
or U7847 (N_7847,N_7126,N_6746);
or U7848 (N_7848,N_6768,N_6465);
xnor U7849 (N_7849,N_7182,N_6669);
and U7850 (N_7850,N_6702,N_6758);
nand U7851 (N_7851,N_7081,N_6981);
nor U7852 (N_7852,N_7067,N_6909);
nor U7853 (N_7853,N_6561,N_6965);
and U7854 (N_7854,N_6818,N_6870);
or U7855 (N_7855,N_7046,N_6581);
or U7856 (N_7856,N_6846,N_7086);
xor U7857 (N_7857,N_6489,N_6729);
and U7858 (N_7858,N_6525,N_6925);
xnor U7859 (N_7859,N_6549,N_7189);
and U7860 (N_7860,N_6577,N_7004);
nand U7861 (N_7861,N_6603,N_7027);
xnor U7862 (N_7862,N_6671,N_6730);
and U7863 (N_7863,N_6666,N_6553);
and U7864 (N_7864,N_6667,N_7078);
nor U7865 (N_7865,N_6928,N_6711);
and U7866 (N_7866,N_6903,N_6502);
nor U7867 (N_7867,N_6901,N_6661);
nor U7868 (N_7868,N_6974,N_6465);
nor U7869 (N_7869,N_7156,N_6537);
nor U7870 (N_7870,N_6534,N_6932);
xnor U7871 (N_7871,N_6666,N_6996);
nor U7872 (N_7872,N_7067,N_6418);
or U7873 (N_7873,N_6448,N_6734);
xnor U7874 (N_7874,N_6662,N_6526);
nor U7875 (N_7875,N_7026,N_6836);
and U7876 (N_7876,N_7047,N_6980);
xor U7877 (N_7877,N_6782,N_6417);
and U7878 (N_7878,N_7125,N_6702);
nand U7879 (N_7879,N_6842,N_6819);
xor U7880 (N_7880,N_6934,N_6935);
nor U7881 (N_7881,N_6782,N_6556);
nand U7882 (N_7882,N_7152,N_7175);
or U7883 (N_7883,N_7099,N_6432);
or U7884 (N_7884,N_6616,N_7002);
xor U7885 (N_7885,N_6430,N_6976);
nor U7886 (N_7886,N_6820,N_6930);
nand U7887 (N_7887,N_6867,N_6985);
or U7888 (N_7888,N_6721,N_6738);
and U7889 (N_7889,N_6771,N_6452);
xnor U7890 (N_7890,N_6940,N_6655);
nand U7891 (N_7891,N_6542,N_7037);
and U7892 (N_7892,N_6896,N_7091);
xor U7893 (N_7893,N_6795,N_6993);
or U7894 (N_7894,N_6832,N_6618);
and U7895 (N_7895,N_6781,N_6811);
or U7896 (N_7896,N_6931,N_6639);
or U7897 (N_7897,N_6918,N_7135);
and U7898 (N_7898,N_6672,N_6482);
nand U7899 (N_7899,N_6429,N_6461);
and U7900 (N_7900,N_6819,N_6402);
nor U7901 (N_7901,N_6701,N_7132);
nand U7902 (N_7902,N_6730,N_7132);
xor U7903 (N_7903,N_6657,N_6817);
nor U7904 (N_7904,N_6726,N_7113);
or U7905 (N_7905,N_6621,N_7084);
xnor U7906 (N_7906,N_6520,N_6822);
nand U7907 (N_7907,N_6710,N_6464);
nor U7908 (N_7908,N_6820,N_7024);
and U7909 (N_7909,N_6640,N_6975);
xnor U7910 (N_7910,N_6412,N_7194);
and U7911 (N_7911,N_6558,N_6710);
xnor U7912 (N_7912,N_6643,N_6439);
and U7913 (N_7913,N_6796,N_6600);
nand U7914 (N_7914,N_7046,N_7185);
and U7915 (N_7915,N_6716,N_6439);
nand U7916 (N_7916,N_6458,N_7096);
nand U7917 (N_7917,N_7091,N_7197);
xor U7918 (N_7918,N_7071,N_6699);
nor U7919 (N_7919,N_6533,N_6409);
or U7920 (N_7920,N_7136,N_6912);
nor U7921 (N_7921,N_6710,N_6695);
nand U7922 (N_7922,N_6617,N_6498);
and U7923 (N_7923,N_6557,N_7050);
and U7924 (N_7924,N_6738,N_6683);
nand U7925 (N_7925,N_7092,N_6510);
and U7926 (N_7926,N_6400,N_7024);
xor U7927 (N_7927,N_6738,N_6420);
or U7928 (N_7928,N_6449,N_6977);
or U7929 (N_7929,N_6452,N_6605);
nand U7930 (N_7930,N_7063,N_7173);
xnor U7931 (N_7931,N_6790,N_6954);
or U7932 (N_7932,N_6795,N_6474);
or U7933 (N_7933,N_6903,N_6549);
nor U7934 (N_7934,N_7110,N_6947);
or U7935 (N_7935,N_6429,N_6762);
xnor U7936 (N_7936,N_6814,N_6628);
xor U7937 (N_7937,N_6732,N_6694);
or U7938 (N_7938,N_6948,N_6753);
and U7939 (N_7939,N_6558,N_7006);
xnor U7940 (N_7940,N_6802,N_6404);
and U7941 (N_7941,N_7071,N_7105);
xnor U7942 (N_7942,N_6776,N_6991);
or U7943 (N_7943,N_6452,N_6966);
nand U7944 (N_7944,N_6898,N_6822);
nand U7945 (N_7945,N_6449,N_7148);
nor U7946 (N_7946,N_7107,N_6762);
xor U7947 (N_7947,N_6759,N_6808);
xnor U7948 (N_7948,N_7126,N_6968);
xor U7949 (N_7949,N_7054,N_6600);
nor U7950 (N_7950,N_6418,N_7174);
and U7951 (N_7951,N_6946,N_6934);
nor U7952 (N_7952,N_6971,N_6651);
and U7953 (N_7953,N_6632,N_6628);
or U7954 (N_7954,N_7112,N_6878);
nand U7955 (N_7955,N_6782,N_6477);
nand U7956 (N_7956,N_7155,N_6513);
and U7957 (N_7957,N_6950,N_6929);
or U7958 (N_7958,N_7028,N_6498);
nand U7959 (N_7959,N_7094,N_7048);
or U7960 (N_7960,N_6408,N_6555);
or U7961 (N_7961,N_6774,N_6645);
or U7962 (N_7962,N_7024,N_6636);
nor U7963 (N_7963,N_6446,N_6488);
or U7964 (N_7964,N_6761,N_6550);
nand U7965 (N_7965,N_7016,N_6589);
and U7966 (N_7966,N_6699,N_6401);
nand U7967 (N_7967,N_6408,N_6508);
or U7968 (N_7968,N_6579,N_6656);
nor U7969 (N_7969,N_6407,N_6834);
nand U7970 (N_7970,N_6742,N_7106);
and U7971 (N_7971,N_6965,N_7086);
or U7972 (N_7972,N_6658,N_6914);
nand U7973 (N_7973,N_6415,N_6559);
nand U7974 (N_7974,N_6681,N_6929);
or U7975 (N_7975,N_6547,N_7133);
xor U7976 (N_7976,N_7121,N_6561);
nor U7977 (N_7977,N_6874,N_6968);
nor U7978 (N_7978,N_7043,N_6493);
xor U7979 (N_7979,N_6598,N_6763);
xnor U7980 (N_7980,N_7111,N_6573);
or U7981 (N_7981,N_6943,N_6929);
xnor U7982 (N_7982,N_6559,N_6489);
or U7983 (N_7983,N_6833,N_6804);
and U7984 (N_7984,N_7057,N_6709);
nand U7985 (N_7985,N_6919,N_6752);
or U7986 (N_7986,N_6550,N_6919);
nand U7987 (N_7987,N_6710,N_6948);
xnor U7988 (N_7988,N_7148,N_7195);
nand U7989 (N_7989,N_7060,N_6984);
nand U7990 (N_7990,N_6853,N_6993);
xnor U7991 (N_7991,N_7128,N_6496);
and U7992 (N_7992,N_7101,N_7025);
xnor U7993 (N_7993,N_7061,N_7068);
nor U7994 (N_7994,N_6874,N_7065);
and U7995 (N_7995,N_6673,N_6583);
and U7996 (N_7996,N_6676,N_6785);
nand U7997 (N_7997,N_6998,N_6868);
or U7998 (N_7998,N_7012,N_7117);
and U7999 (N_7999,N_6931,N_7168);
or U8000 (N_8000,N_7673,N_7916);
or U8001 (N_8001,N_7489,N_7754);
xor U8002 (N_8002,N_7914,N_7412);
nor U8003 (N_8003,N_7960,N_7347);
and U8004 (N_8004,N_7784,N_7574);
xor U8005 (N_8005,N_7456,N_7505);
nor U8006 (N_8006,N_7256,N_7342);
xnor U8007 (N_8007,N_7742,N_7952);
and U8008 (N_8008,N_7668,N_7895);
nand U8009 (N_8009,N_7885,N_7555);
and U8010 (N_8010,N_7706,N_7504);
nor U8011 (N_8011,N_7813,N_7702);
and U8012 (N_8012,N_7277,N_7604);
nand U8013 (N_8013,N_7569,N_7486);
nand U8014 (N_8014,N_7631,N_7925);
and U8015 (N_8015,N_7319,N_7829);
or U8016 (N_8016,N_7619,N_7200);
nand U8017 (N_8017,N_7202,N_7451);
xor U8018 (N_8018,N_7561,N_7876);
or U8019 (N_8019,N_7220,N_7490);
or U8020 (N_8020,N_7753,N_7766);
nor U8021 (N_8021,N_7287,N_7933);
xnor U8022 (N_8022,N_7307,N_7877);
and U8023 (N_8023,N_7691,N_7414);
or U8024 (N_8024,N_7971,N_7441);
nor U8025 (N_8025,N_7799,N_7312);
nand U8026 (N_8026,N_7399,N_7758);
or U8027 (N_8027,N_7208,N_7499);
nor U8028 (N_8028,N_7320,N_7643);
nand U8029 (N_8029,N_7212,N_7756);
nor U8030 (N_8030,N_7720,N_7411);
nor U8031 (N_8031,N_7874,N_7313);
and U8032 (N_8032,N_7944,N_7355);
and U8033 (N_8033,N_7567,N_7258);
or U8034 (N_8034,N_7275,N_7420);
nand U8035 (N_8035,N_7217,N_7632);
xor U8036 (N_8036,N_7357,N_7472);
or U8037 (N_8037,N_7438,N_7390);
nand U8038 (N_8038,N_7846,N_7301);
xor U8039 (N_8039,N_7783,N_7601);
nand U8040 (N_8040,N_7889,N_7857);
nor U8041 (N_8041,N_7350,N_7645);
nand U8042 (N_8042,N_7733,N_7309);
nand U8043 (N_8043,N_7810,N_7366);
or U8044 (N_8044,N_7209,N_7460);
xnor U8045 (N_8045,N_7264,N_7927);
nand U8046 (N_8046,N_7329,N_7918);
or U8047 (N_8047,N_7726,N_7586);
nand U8048 (N_8048,N_7432,N_7470);
nand U8049 (N_8049,N_7576,N_7234);
nor U8050 (N_8050,N_7518,N_7406);
xor U8051 (N_8051,N_7435,N_7932);
nor U8052 (N_8052,N_7279,N_7239);
nor U8053 (N_8053,N_7238,N_7884);
nor U8054 (N_8054,N_7910,N_7980);
or U8055 (N_8055,N_7607,N_7224);
and U8056 (N_8056,N_7936,N_7636);
xnor U8057 (N_8057,N_7969,N_7730);
and U8058 (N_8058,N_7278,N_7848);
xnor U8059 (N_8059,N_7345,N_7340);
xor U8060 (N_8060,N_7901,N_7516);
or U8061 (N_8061,N_7622,N_7316);
nor U8062 (N_8062,N_7304,N_7640);
xnor U8063 (N_8063,N_7739,N_7442);
and U8064 (N_8064,N_7803,N_7262);
xnor U8065 (N_8065,N_7628,N_7699);
or U8066 (N_8066,N_7694,N_7232);
xnor U8067 (N_8067,N_7807,N_7805);
nand U8068 (N_8068,N_7658,N_7377);
xnor U8069 (N_8069,N_7364,N_7245);
nand U8070 (N_8070,N_7983,N_7911);
xnor U8071 (N_8071,N_7426,N_7249);
nand U8072 (N_8072,N_7428,N_7687);
and U8073 (N_8073,N_7346,N_7326);
and U8074 (N_8074,N_7981,N_7297);
and U8075 (N_8075,N_7423,N_7235);
xor U8076 (N_8076,N_7721,N_7370);
xor U8077 (N_8077,N_7533,N_7948);
nor U8078 (N_8078,N_7809,N_7674);
or U8079 (N_8079,N_7882,N_7873);
xnor U8080 (N_8080,N_7651,N_7798);
xor U8081 (N_8081,N_7664,N_7868);
or U8082 (N_8082,N_7255,N_7341);
xnor U8083 (N_8083,N_7861,N_7429);
nor U8084 (N_8084,N_7851,N_7416);
xnor U8085 (N_8085,N_7701,N_7539);
nand U8086 (N_8086,N_7782,N_7265);
xnor U8087 (N_8087,N_7253,N_7482);
or U8088 (N_8088,N_7457,N_7388);
nor U8089 (N_8089,N_7828,N_7290);
and U8090 (N_8090,N_7644,N_7703);
or U8091 (N_8091,N_7716,N_7402);
nor U8092 (N_8092,N_7509,N_7566);
or U8093 (N_8093,N_7833,N_7719);
nand U8094 (N_8094,N_7820,N_7988);
and U8095 (N_8095,N_7863,N_7424);
and U8096 (N_8096,N_7514,N_7707);
xnor U8097 (N_8097,N_7440,N_7930);
xnor U8098 (N_8098,N_7856,N_7656);
or U8099 (N_8099,N_7334,N_7921);
nand U8100 (N_8100,N_7693,N_7998);
nand U8101 (N_8101,N_7718,N_7315);
or U8102 (N_8102,N_7790,N_7878);
or U8103 (N_8103,N_7285,N_7384);
nand U8104 (N_8104,N_7915,N_7800);
or U8105 (N_8105,N_7284,N_7477);
nor U8106 (N_8106,N_7449,N_7547);
nand U8107 (N_8107,N_7450,N_7862);
or U8108 (N_8108,N_7544,N_7240);
nand U8109 (N_8109,N_7273,N_7661);
and U8110 (N_8110,N_7271,N_7589);
nand U8111 (N_8111,N_7478,N_7538);
nand U8112 (N_8112,N_7379,N_7898);
xor U8113 (N_8113,N_7425,N_7582);
and U8114 (N_8114,N_7751,N_7962);
xnor U8115 (N_8115,N_7904,N_7348);
nor U8116 (N_8116,N_7639,N_7503);
and U8117 (N_8117,N_7413,N_7527);
nand U8118 (N_8118,N_7242,N_7943);
nand U8119 (N_8119,N_7532,N_7573);
xnor U8120 (N_8120,N_7864,N_7880);
nand U8121 (N_8121,N_7204,N_7825);
and U8122 (N_8122,N_7463,N_7570);
or U8123 (N_8123,N_7536,N_7627);
nand U8124 (N_8124,N_7793,N_7717);
or U8125 (N_8125,N_7421,N_7996);
xnor U8126 (N_8126,N_7688,N_7966);
xor U8127 (N_8127,N_7458,N_7373);
xnor U8128 (N_8128,N_7343,N_7445);
xor U8129 (N_8129,N_7900,N_7507);
nand U8130 (N_8130,N_7681,N_7974);
nand U8131 (N_8131,N_7741,N_7684);
nor U8132 (N_8132,N_7854,N_7690);
and U8133 (N_8133,N_7587,N_7893);
nand U8134 (N_8134,N_7487,N_7830);
or U8135 (N_8135,N_7203,N_7992);
or U8136 (N_8136,N_7252,N_7484);
xnor U8137 (N_8137,N_7774,N_7723);
nor U8138 (N_8138,N_7579,N_7953);
xor U8139 (N_8139,N_7697,N_7955);
or U8140 (N_8140,N_7906,N_7332);
nand U8141 (N_8141,N_7819,N_7838);
nor U8142 (N_8142,N_7993,N_7372);
and U8143 (N_8143,N_7609,N_7363);
nor U8144 (N_8144,N_7225,N_7443);
xor U8145 (N_8145,N_7709,N_7608);
nor U8146 (N_8146,N_7931,N_7975);
or U8147 (N_8147,N_7466,N_7920);
and U8148 (N_8148,N_7599,N_7229);
xnor U8149 (N_8149,N_7219,N_7374);
xnor U8150 (N_8150,N_7352,N_7792);
nand U8151 (N_8151,N_7559,N_7705);
nor U8152 (N_8152,N_7655,N_7840);
xnor U8153 (N_8153,N_7560,N_7606);
nor U8154 (N_8154,N_7528,N_7750);
or U8155 (N_8155,N_7317,N_7853);
nand U8156 (N_8156,N_7365,N_7427);
and U8157 (N_8157,N_7474,N_7985);
xor U8158 (N_8158,N_7994,N_7529);
xnor U8159 (N_8159,N_7710,N_7376);
nand U8160 (N_8160,N_7328,N_7760);
or U8161 (N_8161,N_7339,N_7801);
nand U8162 (N_8162,N_7437,N_7625);
or U8163 (N_8163,N_7821,N_7353);
xnor U8164 (N_8164,N_7642,N_7879);
nand U8165 (N_8165,N_7795,N_7841);
nor U8166 (N_8166,N_7727,N_7811);
xor U8167 (N_8167,N_7909,N_7712);
nand U8168 (N_8168,N_7945,N_7497);
or U8169 (N_8169,N_7831,N_7613);
and U8170 (N_8170,N_7501,N_7999);
and U8171 (N_8171,N_7737,N_7223);
nand U8172 (N_8172,N_7454,N_7715);
or U8173 (N_8173,N_7548,N_7236);
or U8174 (N_8174,N_7652,N_7294);
and U8175 (N_8175,N_7475,N_7660);
or U8176 (N_8176,N_7585,N_7976);
nor U8177 (N_8177,N_7806,N_7724);
xor U8178 (N_8178,N_7657,N_7939);
nand U8179 (N_8179,N_7344,N_7410);
and U8180 (N_8180,N_7769,N_7823);
and U8181 (N_8181,N_7237,N_7483);
or U8182 (N_8182,N_7896,N_7387);
and U8183 (N_8183,N_7292,N_7666);
or U8184 (N_8184,N_7354,N_7708);
nor U8185 (N_8185,N_7816,N_7205);
and U8186 (N_8186,N_7797,N_7335);
nand U8187 (N_8187,N_7762,N_7796);
or U8188 (N_8188,N_7653,N_7241);
nand U8189 (N_8189,N_7508,N_7700);
and U8190 (N_8190,N_7564,N_7448);
nor U8191 (N_8191,N_7446,N_7471);
nand U8192 (N_8192,N_7493,N_7211);
nand U8193 (N_8193,N_7526,N_7407);
xor U8194 (N_8194,N_7648,N_7722);
and U8195 (N_8195,N_7704,N_7260);
and U8196 (N_8196,N_7485,N_7540);
nor U8197 (N_8197,N_7515,N_7629);
or U8198 (N_8198,N_7360,N_7865);
xor U8199 (N_8199,N_7929,N_7369);
and U8200 (N_8200,N_7593,N_7779);
and U8201 (N_8201,N_7459,N_7283);
nand U8202 (N_8202,N_7665,N_7323);
nor U8203 (N_8203,N_7937,N_7984);
nand U8204 (N_8204,N_7595,N_7512);
or U8205 (N_8205,N_7736,N_7675);
nor U8206 (N_8206,N_7812,N_7767);
nor U8207 (N_8207,N_7250,N_7822);
nor U8208 (N_8208,N_7788,N_7633);
and U8209 (N_8209,N_7391,N_7940);
xnor U8210 (N_8210,N_7965,N_7913);
or U8211 (N_8211,N_7480,N_7630);
and U8212 (N_8212,N_7725,N_7554);
nor U8213 (N_8213,N_7386,N_7867);
nor U8214 (N_8214,N_7226,N_7280);
xnor U8215 (N_8215,N_7957,N_7967);
nand U8216 (N_8216,N_7958,N_7467);
and U8217 (N_8217,N_7327,N_7747);
nor U8218 (N_8218,N_7537,N_7520);
and U8219 (N_8219,N_7695,N_7872);
xnor U8220 (N_8220,N_7973,N_7844);
nor U8221 (N_8221,N_7543,N_7670);
nand U8222 (N_8222,N_7611,N_7761);
or U8223 (N_8223,N_7776,N_7362);
nand U8224 (N_8224,N_7522,N_7845);
and U8225 (N_8225,N_7511,N_7447);
nor U8226 (N_8226,N_7519,N_7917);
or U8227 (N_8227,N_7358,N_7650);
or U8228 (N_8228,N_7602,N_7979);
nor U8229 (N_8229,N_7257,N_7689);
nor U8230 (N_8230,N_7274,N_7883);
nand U8231 (N_8231,N_7468,N_7214);
and U8232 (N_8232,N_7254,N_7903);
and U8233 (N_8233,N_7531,N_7588);
xnor U8234 (N_8234,N_7562,N_7247);
or U8235 (N_8235,N_7455,N_7295);
nor U8236 (N_8236,N_7565,N_7771);
xor U8237 (N_8237,N_7382,N_7899);
nand U8238 (N_8238,N_7785,N_7433);
and U8239 (N_8239,N_7781,N_7575);
nor U8240 (N_8240,N_7298,N_7698);
nand U8241 (N_8241,N_7336,N_7772);
or U8242 (N_8242,N_7215,N_7246);
or U8243 (N_8243,N_7941,N_7759);
xnor U8244 (N_8244,N_7963,N_7635);
nand U8245 (N_8245,N_7870,N_7680);
or U8246 (N_8246,N_7299,N_7623);
xor U8247 (N_8247,N_7852,N_7495);
and U8248 (N_8248,N_7321,N_7732);
xnor U8249 (N_8249,N_7886,N_7318);
or U8250 (N_8250,N_7462,N_7902);
nor U8251 (N_8251,N_7938,N_7907);
and U8252 (N_8252,N_7453,N_7481);
xnor U8253 (N_8253,N_7525,N_7912);
or U8254 (N_8254,N_7836,N_7734);
xnor U8255 (N_8255,N_7972,N_7530);
xor U8256 (N_8256,N_7634,N_7371);
nor U8257 (N_8257,N_7881,N_7594);
or U8258 (N_8258,N_7558,N_7266);
or U8259 (N_8259,N_7310,N_7415);
nand U8260 (N_8260,N_7677,N_7305);
nor U8261 (N_8261,N_7534,N_7649);
or U8262 (N_8262,N_7682,N_7934);
nand U8263 (N_8263,N_7638,N_7991);
and U8264 (N_8264,N_7465,N_7667);
or U8265 (N_8265,N_7524,N_7926);
and U8266 (N_8266,N_7464,N_7696);
and U8267 (N_8267,N_7590,N_7891);
nand U8268 (N_8268,N_7637,N_7578);
and U8269 (N_8269,N_7678,N_7614);
nand U8270 (N_8270,N_7672,N_7206);
nor U8271 (N_8271,N_7815,N_7461);
xor U8272 (N_8272,N_7887,N_7408);
nor U8273 (N_8273,N_7397,N_7671);
nor U8274 (N_8274,N_7654,N_7331);
nand U8275 (N_8275,N_7647,N_7418);
xnor U8276 (N_8276,N_7230,N_7591);
nand U8277 (N_8277,N_7804,N_7977);
nand U8278 (N_8278,N_7735,N_7479);
and U8279 (N_8279,N_7871,N_7968);
nor U8280 (N_8280,N_7289,N_7227);
or U8281 (N_8281,N_7404,N_7905);
nor U8282 (N_8282,N_7251,N_7598);
and U8283 (N_8283,N_7282,N_7286);
nor U8284 (N_8284,N_7683,N_7835);
xnor U8285 (N_8285,N_7866,N_7949);
nand U8286 (N_8286,N_7603,N_7248);
and U8287 (N_8287,N_7859,N_7947);
nor U8288 (N_8288,N_7763,N_7584);
and U8289 (N_8289,N_7431,N_7349);
xor U8290 (N_8290,N_7288,N_7296);
nor U8291 (N_8291,N_7616,N_7403);
nor U8292 (N_8292,N_7597,N_7492);
xor U8293 (N_8293,N_7535,N_7686);
xor U8294 (N_8294,N_7860,N_7995);
and U8295 (N_8295,N_7213,N_7990);
nand U8296 (N_8296,N_7385,N_7263);
nor U8297 (N_8297,N_7476,N_7961);
xnor U8298 (N_8298,N_7351,N_7314);
nand U8299 (N_8299,N_7814,N_7714);
and U8300 (N_8300,N_7333,N_7581);
nor U8301 (N_8301,N_7592,N_7568);
nand U8302 (N_8302,N_7729,N_7434);
or U8303 (N_8303,N_7291,N_7243);
and U8304 (N_8304,N_7610,N_7617);
and U8305 (N_8305,N_7325,N_7268);
or U8306 (N_8306,N_7378,N_7620);
and U8307 (N_8307,N_7843,N_7794);
nand U8308 (N_8308,N_7261,N_7400);
and U8309 (N_8309,N_7942,N_7626);
or U8310 (N_8310,N_7837,N_7713);
or U8311 (N_8311,N_7970,N_7989);
or U8312 (N_8312,N_7791,N_7618);
or U8313 (N_8313,N_7430,N_7389);
or U8314 (N_8314,N_7546,N_7338);
nor U8315 (N_8315,N_7605,N_7201);
xnor U8316 (N_8316,N_7749,N_7818);
nor U8317 (N_8317,N_7473,N_7600);
xnor U8318 (N_8318,N_7897,N_7875);
or U8319 (N_8319,N_7523,N_7778);
nand U8320 (N_8320,N_7571,N_7808);
xor U8321 (N_8321,N_7302,N_7768);
nor U8322 (N_8322,N_7281,N_7502);
or U8323 (N_8323,N_7777,N_7839);
nor U8324 (N_8324,N_7221,N_7744);
xnor U8325 (N_8325,N_7383,N_7692);
or U8326 (N_8326,N_7272,N_7773);
xor U8327 (N_8327,N_7394,N_7923);
nor U8328 (N_8328,N_7827,N_7826);
nand U8329 (N_8329,N_7924,N_7375);
nand U8330 (N_8330,N_7517,N_7303);
and U8331 (N_8331,N_7858,N_7919);
or U8332 (N_8332,N_7308,N_7405);
or U8333 (N_8333,N_7469,N_7842);
nand U8334 (N_8334,N_7954,N_7577);
or U8335 (N_8335,N_7210,N_7824);
or U8336 (N_8336,N_7367,N_7337);
nor U8337 (N_8337,N_7491,N_7817);
nand U8338 (N_8338,N_7552,N_7269);
nor U8339 (N_8339,N_7436,N_7765);
or U8340 (N_8340,N_7545,N_7787);
xor U8341 (N_8341,N_7986,N_7521);
and U8342 (N_8342,N_7422,N_7646);
nand U8343 (N_8343,N_7513,N_7832);
or U8344 (N_8344,N_7580,N_7745);
and U8345 (N_8345,N_7946,N_7306);
xor U8346 (N_8346,N_7496,N_7869);
nand U8347 (N_8347,N_7951,N_7802);
or U8348 (N_8348,N_7401,N_7956);
nand U8349 (N_8349,N_7596,N_7615);
or U8350 (N_8350,N_7572,N_7922);
and U8351 (N_8351,N_7556,N_7359);
nand U8352 (N_8352,N_7270,N_7669);
xor U8353 (N_8353,N_7659,N_7786);
nand U8354 (N_8354,N_7935,N_7356);
and U8355 (N_8355,N_7894,N_7506);
nand U8356 (N_8356,N_7452,N_7850);
and U8357 (N_8357,N_7324,N_7711);
or U8358 (N_8358,N_7293,N_7216);
nor U8359 (N_8359,N_7380,N_7959);
or U8360 (N_8360,N_7557,N_7322);
nor U8361 (N_8361,N_7276,N_7381);
or U8362 (N_8362,N_7928,N_7419);
nand U8363 (N_8363,N_7662,N_7409);
nand U8364 (N_8364,N_7764,N_7982);
or U8365 (N_8365,N_7488,N_7740);
and U8366 (N_8366,N_7494,N_7855);
or U8367 (N_8367,N_7392,N_7510);
and U8368 (N_8368,N_7498,N_7641);
and U8369 (N_8369,N_7755,N_7621);
nand U8370 (N_8370,N_7950,N_7233);
xor U8371 (N_8371,N_7542,N_7398);
or U8372 (N_8372,N_7624,N_7789);
and U8373 (N_8373,N_7228,N_7849);
nor U8374 (N_8374,N_7997,N_7311);
nand U8375 (N_8375,N_7892,N_7222);
or U8376 (N_8376,N_7847,N_7218);
nor U8377 (N_8377,N_7888,N_7444);
and U8378 (N_8378,N_7541,N_7676);
xnor U8379 (N_8379,N_7550,N_7890);
and U8380 (N_8380,N_7563,N_7834);
and U8381 (N_8381,N_7964,N_7553);
xnor U8382 (N_8382,N_7259,N_7738);
or U8383 (N_8383,N_7612,N_7207);
or U8384 (N_8384,N_7330,N_7396);
nand U8385 (N_8385,N_7780,N_7731);
nor U8386 (N_8386,N_7500,N_7361);
nand U8387 (N_8387,N_7987,N_7978);
nand U8388 (N_8388,N_7417,N_7368);
nand U8389 (N_8389,N_7549,N_7908);
and U8390 (N_8390,N_7267,N_7393);
nor U8391 (N_8391,N_7583,N_7770);
nand U8392 (N_8392,N_7231,N_7746);
nand U8393 (N_8393,N_7551,N_7663);
xnor U8394 (N_8394,N_7300,N_7728);
nor U8395 (N_8395,N_7757,N_7752);
nor U8396 (N_8396,N_7685,N_7748);
or U8397 (N_8397,N_7743,N_7244);
and U8398 (N_8398,N_7395,N_7679);
nor U8399 (N_8399,N_7439,N_7775);
nand U8400 (N_8400,N_7855,N_7455);
and U8401 (N_8401,N_7739,N_7627);
xnor U8402 (N_8402,N_7597,N_7470);
or U8403 (N_8403,N_7326,N_7982);
nand U8404 (N_8404,N_7924,N_7343);
and U8405 (N_8405,N_7684,N_7567);
or U8406 (N_8406,N_7396,N_7445);
nor U8407 (N_8407,N_7450,N_7580);
xor U8408 (N_8408,N_7843,N_7858);
xor U8409 (N_8409,N_7998,N_7589);
or U8410 (N_8410,N_7992,N_7425);
nand U8411 (N_8411,N_7572,N_7941);
or U8412 (N_8412,N_7885,N_7376);
and U8413 (N_8413,N_7452,N_7985);
nand U8414 (N_8414,N_7691,N_7679);
xor U8415 (N_8415,N_7720,N_7923);
xor U8416 (N_8416,N_7357,N_7752);
and U8417 (N_8417,N_7548,N_7774);
and U8418 (N_8418,N_7996,N_7894);
nor U8419 (N_8419,N_7525,N_7949);
xor U8420 (N_8420,N_7339,N_7253);
nand U8421 (N_8421,N_7804,N_7481);
nand U8422 (N_8422,N_7930,N_7300);
or U8423 (N_8423,N_7782,N_7344);
xor U8424 (N_8424,N_7836,N_7956);
xnor U8425 (N_8425,N_7294,N_7493);
xnor U8426 (N_8426,N_7792,N_7801);
nand U8427 (N_8427,N_7896,N_7332);
or U8428 (N_8428,N_7709,N_7424);
nor U8429 (N_8429,N_7588,N_7273);
nand U8430 (N_8430,N_7669,N_7695);
nand U8431 (N_8431,N_7965,N_7497);
nor U8432 (N_8432,N_7831,N_7982);
xnor U8433 (N_8433,N_7927,N_7812);
or U8434 (N_8434,N_7367,N_7265);
nor U8435 (N_8435,N_7397,N_7328);
nor U8436 (N_8436,N_7728,N_7223);
nand U8437 (N_8437,N_7513,N_7619);
xor U8438 (N_8438,N_7528,N_7280);
xnor U8439 (N_8439,N_7410,N_7356);
nand U8440 (N_8440,N_7839,N_7856);
nand U8441 (N_8441,N_7845,N_7868);
xor U8442 (N_8442,N_7523,N_7591);
or U8443 (N_8443,N_7286,N_7317);
and U8444 (N_8444,N_7672,N_7518);
and U8445 (N_8445,N_7372,N_7269);
nor U8446 (N_8446,N_7967,N_7665);
or U8447 (N_8447,N_7278,N_7630);
nor U8448 (N_8448,N_7419,N_7471);
and U8449 (N_8449,N_7795,N_7524);
nor U8450 (N_8450,N_7225,N_7657);
xor U8451 (N_8451,N_7487,N_7491);
nand U8452 (N_8452,N_7930,N_7606);
or U8453 (N_8453,N_7477,N_7476);
nand U8454 (N_8454,N_7890,N_7971);
nor U8455 (N_8455,N_7745,N_7457);
or U8456 (N_8456,N_7546,N_7472);
nor U8457 (N_8457,N_7835,N_7307);
nor U8458 (N_8458,N_7822,N_7888);
or U8459 (N_8459,N_7622,N_7557);
nor U8460 (N_8460,N_7823,N_7843);
and U8461 (N_8461,N_7615,N_7528);
and U8462 (N_8462,N_7808,N_7574);
nor U8463 (N_8463,N_7500,N_7410);
nand U8464 (N_8464,N_7688,N_7581);
nand U8465 (N_8465,N_7513,N_7933);
nand U8466 (N_8466,N_7859,N_7626);
or U8467 (N_8467,N_7704,N_7513);
nand U8468 (N_8468,N_7564,N_7452);
or U8469 (N_8469,N_7825,N_7815);
or U8470 (N_8470,N_7788,N_7760);
or U8471 (N_8471,N_7553,N_7735);
nand U8472 (N_8472,N_7660,N_7890);
nand U8473 (N_8473,N_7604,N_7420);
nor U8474 (N_8474,N_7354,N_7626);
nor U8475 (N_8475,N_7200,N_7792);
and U8476 (N_8476,N_7234,N_7957);
or U8477 (N_8477,N_7884,N_7784);
nor U8478 (N_8478,N_7662,N_7303);
and U8479 (N_8479,N_7266,N_7396);
nor U8480 (N_8480,N_7675,N_7767);
nand U8481 (N_8481,N_7586,N_7338);
xor U8482 (N_8482,N_7355,N_7405);
nor U8483 (N_8483,N_7386,N_7228);
nor U8484 (N_8484,N_7482,N_7825);
and U8485 (N_8485,N_7698,N_7482);
nor U8486 (N_8486,N_7760,N_7666);
nand U8487 (N_8487,N_7823,N_7862);
or U8488 (N_8488,N_7738,N_7592);
and U8489 (N_8489,N_7815,N_7384);
or U8490 (N_8490,N_7585,N_7726);
xnor U8491 (N_8491,N_7863,N_7292);
nor U8492 (N_8492,N_7645,N_7625);
and U8493 (N_8493,N_7383,N_7800);
xor U8494 (N_8494,N_7927,N_7667);
xor U8495 (N_8495,N_7559,N_7978);
xnor U8496 (N_8496,N_7587,N_7771);
nand U8497 (N_8497,N_7752,N_7470);
xor U8498 (N_8498,N_7970,N_7813);
nor U8499 (N_8499,N_7962,N_7828);
or U8500 (N_8500,N_7988,N_7255);
nand U8501 (N_8501,N_7609,N_7704);
nand U8502 (N_8502,N_7343,N_7285);
and U8503 (N_8503,N_7620,N_7460);
and U8504 (N_8504,N_7614,N_7766);
and U8505 (N_8505,N_7687,N_7730);
and U8506 (N_8506,N_7801,N_7648);
nor U8507 (N_8507,N_7926,N_7536);
nand U8508 (N_8508,N_7823,N_7468);
or U8509 (N_8509,N_7488,N_7205);
or U8510 (N_8510,N_7374,N_7710);
or U8511 (N_8511,N_7230,N_7580);
nand U8512 (N_8512,N_7668,N_7741);
and U8513 (N_8513,N_7535,N_7522);
xnor U8514 (N_8514,N_7606,N_7610);
nand U8515 (N_8515,N_7773,N_7626);
and U8516 (N_8516,N_7570,N_7205);
nor U8517 (N_8517,N_7447,N_7498);
nand U8518 (N_8518,N_7220,N_7824);
and U8519 (N_8519,N_7552,N_7212);
xnor U8520 (N_8520,N_7523,N_7541);
nand U8521 (N_8521,N_7803,N_7971);
xor U8522 (N_8522,N_7489,N_7388);
xor U8523 (N_8523,N_7396,N_7908);
xor U8524 (N_8524,N_7282,N_7237);
or U8525 (N_8525,N_7458,N_7871);
or U8526 (N_8526,N_7518,N_7425);
or U8527 (N_8527,N_7697,N_7786);
or U8528 (N_8528,N_7452,N_7894);
nor U8529 (N_8529,N_7436,N_7273);
nor U8530 (N_8530,N_7876,N_7920);
or U8531 (N_8531,N_7307,N_7765);
or U8532 (N_8532,N_7314,N_7715);
nor U8533 (N_8533,N_7261,N_7315);
and U8534 (N_8534,N_7779,N_7848);
or U8535 (N_8535,N_7222,N_7908);
xnor U8536 (N_8536,N_7803,N_7425);
xor U8537 (N_8537,N_7483,N_7667);
nor U8538 (N_8538,N_7204,N_7601);
xnor U8539 (N_8539,N_7487,N_7762);
nand U8540 (N_8540,N_7219,N_7524);
nor U8541 (N_8541,N_7607,N_7893);
xor U8542 (N_8542,N_7947,N_7919);
or U8543 (N_8543,N_7929,N_7510);
and U8544 (N_8544,N_7526,N_7960);
nand U8545 (N_8545,N_7328,N_7591);
or U8546 (N_8546,N_7547,N_7859);
and U8547 (N_8547,N_7532,N_7386);
and U8548 (N_8548,N_7318,N_7549);
and U8549 (N_8549,N_7495,N_7537);
nand U8550 (N_8550,N_7975,N_7457);
nor U8551 (N_8551,N_7737,N_7885);
and U8552 (N_8552,N_7924,N_7719);
xnor U8553 (N_8553,N_7947,N_7591);
xnor U8554 (N_8554,N_7634,N_7767);
and U8555 (N_8555,N_7472,N_7224);
nor U8556 (N_8556,N_7525,N_7356);
nand U8557 (N_8557,N_7395,N_7221);
nor U8558 (N_8558,N_7762,N_7864);
nor U8559 (N_8559,N_7622,N_7609);
nor U8560 (N_8560,N_7489,N_7602);
nand U8561 (N_8561,N_7244,N_7560);
nand U8562 (N_8562,N_7586,N_7291);
and U8563 (N_8563,N_7252,N_7693);
nand U8564 (N_8564,N_7623,N_7223);
nand U8565 (N_8565,N_7848,N_7547);
nand U8566 (N_8566,N_7231,N_7805);
or U8567 (N_8567,N_7261,N_7529);
xnor U8568 (N_8568,N_7885,N_7702);
or U8569 (N_8569,N_7706,N_7341);
xnor U8570 (N_8570,N_7288,N_7819);
nand U8571 (N_8571,N_7219,N_7614);
nor U8572 (N_8572,N_7763,N_7597);
nand U8573 (N_8573,N_7223,N_7634);
nand U8574 (N_8574,N_7607,N_7687);
and U8575 (N_8575,N_7933,N_7376);
nor U8576 (N_8576,N_7772,N_7965);
nor U8577 (N_8577,N_7209,N_7771);
xnor U8578 (N_8578,N_7930,N_7328);
nand U8579 (N_8579,N_7964,N_7892);
xor U8580 (N_8580,N_7699,N_7205);
or U8581 (N_8581,N_7608,N_7210);
or U8582 (N_8582,N_7943,N_7219);
and U8583 (N_8583,N_7961,N_7898);
xor U8584 (N_8584,N_7311,N_7582);
nor U8585 (N_8585,N_7852,N_7307);
or U8586 (N_8586,N_7662,N_7325);
or U8587 (N_8587,N_7300,N_7833);
or U8588 (N_8588,N_7297,N_7646);
nand U8589 (N_8589,N_7240,N_7652);
nand U8590 (N_8590,N_7408,N_7666);
nand U8591 (N_8591,N_7380,N_7935);
or U8592 (N_8592,N_7830,N_7510);
nand U8593 (N_8593,N_7942,N_7460);
xor U8594 (N_8594,N_7843,N_7554);
nor U8595 (N_8595,N_7302,N_7643);
xor U8596 (N_8596,N_7576,N_7826);
xnor U8597 (N_8597,N_7896,N_7935);
xor U8598 (N_8598,N_7258,N_7990);
xnor U8599 (N_8599,N_7853,N_7742);
xor U8600 (N_8600,N_7822,N_7707);
xor U8601 (N_8601,N_7565,N_7449);
xnor U8602 (N_8602,N_7796,N_7429);
xor U8603 (N_8603,N_7242,N_7732);
nand U8604 (N_8604,N_7707,N_7814);
nor U8605 (N_8605,N_7736,N_7639);
xor U8606 (N_8606,N_7952,N_7877);
xor U8607 (N_8607,N_7457,N_7825);
nor U8608 (N_8608,N_7396,N_7292);
nand U8609 (N_8609,N_7877,N_7325);
or U8610 (N_8610,N_7242,N_7404);
nor U8611 (N_8611,N_7529,N_7966);
xor U8612 (N_8612,N_7637,N_7392);
nand U8613 (N_8613,N_7238,N_7565);
xnor U8614 (N_8614,N_7904,N_7454);
xnor U8615 (N_8615,N_7935,N_7639);
nand U8616 (N_8616,N_7353,N_7954);
xor U8617 (N_8617,N_7944,N_7836);
nand U8618 (N_8618,N_7623,N_7603);
nor U8619 (N_8619,N_7467,N_7824);
and U8620 (N_8620,N_7648,N_7905);
and U8621 (N_8621,N_7899,N_7482);
or U8622 (N_8622,N_7779,N_7499);
or U8623 (N_8623,N_7905,N_7405);
xor U8624 (N_8624,N_7693,N_7455);
xor U8625 (N_8625,N_7941,N_7726);
nand U8626 (N_8626,N_7837,N_7284);
and U8627 (N_8627,N_7739,N_7805);
nand U8628 (N_8628,N_7398,N_7264);
xnor U8629 (N_8629,N_7242,N_7691);
nand U8630 (N_8630,N_7415,N_7747);
xnor U8631 (N_8631,N_7331,N_7294);
nor U8632 (N_8632,N_7993,N_7909);
and U8633 (N_8633,N_7495,N_7643);
xor U8634 (N_8634,N_7343,N_7733);
or U8635 (N_8635,N_7997,N_7864);
xnor U8636 (N_8636,N_7317,N_7981);
nor U8637 (N_8637,N_7305,N_7420);
or U8638 (N_8638,N_7521,N_7910);
or U8639 (N_8639,N_7785,N_7783);
and U8640 (N_8640,N_7946,N_7750);
nand U8641 (N_8641,N_7986,N_7863);
and U8642 (N_8642,N_7661,N_7219);
xor U8643 (N_8643,N_7896,N_7527);
xnor U8644 (N_8644,N_7239,N_7241);
or U8645 (N_8645,N_7864,N_7902);
or U8646 (N_8646,N_7711,N_7253);
nand U8647 (N_8647,N_7216,N_7781);
and U8648 (N_8648,N_7715,N_7296);
or U8649 (N_8649,N_7639,N_7285);
xor U8650 (N_8650,N_7274,N_7309);
nor U8651 (N_8651,N_7820,N_7951);
and U8652 (N_8652,N_7222,N_7764);
xor U8653 (N_8653,N_7869,N_7692);
xor U8654 (N_8654,N_7538,N_7727);
nor U8655 (N_8655,N_7533,N_7943);
and U8656 (N_8656,N_7839,N_7952);
xor U8657 (N_8657,N_7657,N_7794);
nand U8658 (N_8658,N_7509,N_7275);
nor U8659 (N_8659,N_7822,N_7228);
nor U8660 (N_8660,N_7414,N_7704);
or U8661 (N_8661,N_7935,N_7351);
xor U8662 (N_8662,N_7873,N_7567);
nand U8663 (N_8663,N_7527,N_7710);
or U8664 (N_8664,N_7345,N_7955);
xor U8665 (N_8665,N_7529,N_7260);
nand U8666 (N_8666,N_7950,N_7915);
and U8667 (N_8667,N_7896,N_7496);
or U8668 (N_8668,N_7708,N_7324);
and U8669 (N_8669,N_7961,N_7803);
and U8670 (N_8670,N_7259,N_7565);
and U8671 (N_8671,N_7639,N_7977);
nand U8672 (N_8672,N_7311,N_7628);
nor U8673 (N_8673,N_7248,N_7985);
and U8674 (N_8674,N_7227,N_7579);
nand U8675 (N_8675,N_7469,N_7938);
nor U8676 (N_8676,N_7500,N_7946);
nand U8677 (N_8677,N_7714,N_7269);
or U8678 (N_8678,N_7601,N_7591);
and U8679 (N_8679,N_7634,N_7292);
xor U8680 (N_8680,N_7853,N_7696);
or U8681 (N_8681,N_7754,N_7790);
xor U8682 (N_8682,N_7411,N_7590);
nor U8683 (N_8683,N_7282,N_7968);
xor U8684 (N_8684,N_7390,N_7514);
or U8685 (N_8685,N_7453,N_7835);
nor U8686 (N_8686,N_7803,N_7742);
nor U8687 (N_8687,N_7401,N_7315);
xor U8688 (N_8688,N_7826,N_7823);
xor U8689 (N_8689,N_7572,N_7584);
xor U8690 (N_8690,N_7377,N_7973);
and U8691 (N_8691,N_7970,N_7967);
or U8692 (N_8692,N_7426,N_7395);
or U8693 (N_8693,N_7775,N_7938);
nand U8694 (N_8694,N_7803,N_7904);
nor U8695 (N_8695,N_7836,N_7843);
nor U8696 (N_8696,N_7643,N_7323);
nor U8697 (N_8697,N_7564,N_7914);
nand U8698 (N_8698,N_7544,N_7843);
and U8699 (N_8699,N_7428,N_7361);
nand U8700 (N_8700,N_7890,N_7607);
and U8701 (N_8701,N_7233,N_7635);
or U8702 (N_8702,N_7795,N_7239);
or U8703 (N_8703,N_7482,N_7846);
or U8704 (N_8704,N_7685,N_7482);
xnor U8705 (N_8705,N_7672,N_7538);
nand U8706 (N_8706,N_7362,N_7722);
nor U8707 (N_8707,N_7545,N_7227);
or U8708 (N_8708,N_7678,N_7370);
and U8709 (N_8709,N_7610,N_7859);
nor U8710 (N_8710,N_7460,N_7693);
nand U8711 (N_8711,N_7587,N_7549);
nor U8712 (N_8712,N_7454,N_7804);
or U8713 (N_8713,N_7657,N_7899);
or U8714 (N_8714,N_7960,N_7202);
nand U8715 (N_8715,N_7992,N_7945);
or U8716 (N_8716,N_7483,N_7315);
nor U8717 (N_8717,N_7490,N_7617);
nor U8718 (N_8718,N_7449,N_7827);
and U8719 (N_8719,N_7341,N_7827);
and U8720 (N_8720,N_7516,N_7987);
nand U8721 (N_8721,N_7729,N_7275);
nand U8722 (N_8722,N_7267,N_7937);
and U8723 (N_8723,N_7921,N_7613);
or U8724 (N_8724,N_7811,N_7804);
nand U8725 (N_8725,N_7727,N_7306);
xnor U8726 (N_8726,N_7966,N_7586);
xnor U8727 (N_8727,N_7606,N_7581);
nor U8728 (N_8728,N_7771,N_7761);
nor U8729 (N_8729,N_7909,N_7269);
and U8730 (N_8730,N_7474,N_7934);
nand U8731 (N_8731,N_7512,N_7949);
or U8732 (N_8732,N_7598,N_7406);
nor U8733 (N_8733,N_7624,N_7958);
nor U8734 (N_8734,N_7442,N_7471);
nor U8735 (N_8735,N_7203,N_7736);
and U8736 (N_8736,N_7704,N_7711);
nor U8737 (N_8737,N_7540,N_7576);
nand U8738 (N_8738,N_7627,N_7341);
or U8739 (N_8739,N_7287,N_7806);
nand U8740 (N_8740,N_7264,N_7813);
nand U8741 (N_8741,N_7383,N_7736);
or U8742 (N_8742,N_7566,N_7888);
xor U8743 (N_8743,N_7314,N_7877);
nor U8744 (N_8744,N_7658,N_7811);
or U8745 (N_8745,N_7294,N_7241);
and U8746 (N_8746,N_7627,N_7657);
and U8747 (N_8747,N_7640,N_7892);
and U8748 (N_8748,N_7985,N_7849);
and U8749 (N_8749,N_7402,N_7636);
xnor U8750 (N_8750,N_7366,N_7663);
xor U8751 (N_8751,N_7991,N_7335);
xor U8752 (N_8752,N_7636,N_7645);
nor U8753 (N_8753,N_7801,N_7516);
and U8754 (N_8754,N_7698,N_7317);
nor U8755 (N_8755,N_7787,N_7727);
or U8756 (N_8756,N_7299,N_7844);
and U8757 (N_8757,N_7604,N_7351);
xor U8758 (N_8758,N_7754,N_7663);
nor U8759 (N_8759,N_7672,N_7936);
and U8760 (N_8760,N_7303,N_7266);
or U8761 (N_8761,N_7370,N_7231);
nand U8762 (N_8762,N_7333,N_7739);
nor U8763 (N_8763,N_7289,N_7279);
and U8764 (N_8764,N_7659,N_7678);
xnor U8765 (N_8765,N_7854,N_7824);
or U8766 (N_8766,N_7394,N_7436);
nand U8767 (N_8767,N_7778,N_7462);
nand U8768 (N_8768,N_7514,N_7212);
nor U8769 (N_8769,N_7257,N_7385);
and U8770 (N_8770,N_7406,N_7227);
and U8771 (N_8771,N_7233,N_7945);
xnor U8772 (N_8772,N_7754,N_7340);
and U8773 (N_8773,N_7360,N_7437);
or U8774 (N_8774,N_7650,N_7229);
or U8775 (N_8775,N_7990,N_7616);
nor U8776 (N_8776,N_7255,N_7393);
xnor U8777 (N_8777,N_7651,N_7881);
nor U8778 (N_8778,N_7520,N_7839);
or U8779 (N_8779,N_7659,N_7203);
xnor U8780 (N_8780,N_7938,N_7427);
nor U8781 (N_8781,N_7256,N_7530);
nand U8782 (N_8782,N_7918,N_7517);
or U8783 (N_8783,N_7980,N_7339);
and U8784 (N_8784,N_7742,N_7747);
and U8785 (N_8785,N_7610,N_7825);
and U8786 (N_8786,N_7798,N_7626);
and U8787 (N_8787,N_7377,N_7311);
nor U8788 (N_8788,N_7596,N_7606);
xor U8789 (N_8789,N_7230,N_7584);
xor U8790 (N_8790,N_7541,N_7908);
or U8791 (N_8791,N_7418,N_7228);
nand U8792 (N_8792,N_7875,N_7945);
nor U8793 (N_8793,N_7217,N_7607);
and U8794 (N_8794,N_7480,N_7541);
xnor U8795 (N_8795,N_7979,N_7792);
nor U8796 (N_8796,N_7590,N_7916);
nor U8797 (N_8797,N_7662,N_7423);
xnor U8798 (N_8798,N_7908,N_7339);
nor U8799 (N_8799,N_7268,N_7857);
and U8800 (N_8800,N_8260,N_8309);
or U8801 (N_8801,N_8476,N_8473);
nor U8802 (N_8802,N_8168,N_8154);
xnor U8803 (N_8803,N_8676,N_8758);
xnor U8804 (N_8804,N_8101,N_8080);
nand U8805 (N_8805,N_8798,N_8112);
xor U8806 (N_8806,N_8070,N_8714);
xor U8807 (N_8807,N_8507,N_8323);
nor U8808 (N_8808,N_8413,N_8647);
nand U8809 (N_8809,N_8698,N_8635);
xnor U8810 (N_8810,N_8582,N_8001);
nor U8811 (N_8811,N_8567,N_8304);
nor U8812 (N_8812,N_8445,N_8409);
xnor U8813 (N_8813,N_8663,N_8143);
or U8814 (N_8814,N_8435,N_8297);
nor U8815 (N_8815,N_8633,N_8623);
nor U8816 (N_8816,N_8419,N_8495);
nand U8817 (N_8817,N_8064,N_8439);
nor U8818 (N_8818,N_8328,N_8670);
nor U8819 (N_8819,N_8406,N_8162);
and U8820 (N_8820,N_8580,N_8277);
or U8821 (N_8821,N_8730,N_8648);
nor U8822 (N_8822,N_8308,N_8382);
or U8823 (N_8823,N_8303,N_8478);
nand U8824 (N_8824,N_8751,N_8528);
xnor U8825 (N_8825,N_8604,N_8142);
and U8826 (N_8826,N_8174,N_8606);
xor U8827 (N_8827,N_8190,N_8431);
nor U8828 (N_8828,N_8680,N_8315);
nand U8829 (N_8829,N_8270,N_8205);
xnor U8830 (N_8830,N_8152,N_8498);
and U8831 (N_8831,N_8385,N_8570);
and U8832 (N_8832,N_8492,N_8776);
and U8833 (N_8833,N_8150,N_8373);
and U8834 (N_8834,N_8756,N_8223);
xor U8835 (N_8835,N_8600,N_8561);
or U8836 (N_8836,N_8319,N_8017);
or U8837 (N_8837,N_8133,N_8559);
and U8838 (N_8838,N_8306,N_8464);
xor U8839 (N_8839,N_8192,N_8639);
nand U8840 (N_8840,N_8265,N_8029);
nand U8841 (N_8841,N_8114,N_8593);
nor U8842 (N_8842,N_8259,N_8653);
and U8843 (N_8843,N_8049,N_8622);
xor U8844 (N_8844,N_8025,N_8766);
and U8845 (N_8845,N_8658,N_8674);
and U8846 (N_8846,N_8273,N_8396);
nor U8847 (N_8847,N_8734,N_8624);
xnor U8848 (N_8848,N_8264,N_8295);
and U8849 (N_8849,N_8448,N_8657);
nand U8850 (N_8850,N_8208,N_8719);
nor U8851 (N_8851,N_8778,N_8748);
nand U8852 (N_8852,N_8553,N_8386);
nor U8853 (N_8853,N_8089,N_8481);
or U8854 (N_8854,N_8075,N_8677);
nand U8855 (N_8855,N_8661,N_8603);
nand U8856 (N_8856,N_8221,N_8146);
xnor U8857 (N_8857,N_8428,N_8337);
nand U8858 (N_8858,N_8185,N_8348);
or U8859 (N_8859,N_8762,N_8510);
and U8860 (N_8860,N_8280,N_8131);
or U8861 (N_8861,N_8708,N_8384);
or U8862 (N_8862,N_8166,N_8254);
nand U8863 (N_8863,N_8668,N_8556);
or U8864 (N_8864,N_8235,N_8506);
or U8865 (N_8865,N_8342,N_8576);
and U8866 (N_8866,N_8753,N_8151);
xor U8867 (N_8867,N_8740,N_8249);
or U8868 (N_8868,N_8334,N_8052);
nand U8869 (N_8869,N_8388,N_8057);
xnor U8870 (N_8870,N_8551,N_8522);
nand U8871 (N_8871,N_8568,N_8736);
nand U8872 (N_8872,N_8521,N_8482);
xor U8873 (N_8873,N_8098,N_8126);
xor U8874 (N_8874,N_8330,N_8581);
nand U8875 (N_8875,N_8183,N_8302);
or U8876 (N_8876,N_8372,N_8283);
nand U8877 (N_8877,N_8312,N_8028);
nor U8878 (N_8878,N_8662,N_8757);
or U8879 (N_8879,N_8161,N_8038);
and U8880 (N_8880,N_8686,N_8368);
xnor U8881 (N_8881,N_8298,N_8588);
nand U8882 (N_8882,N_8353,N_8761);
nand U8883 (N_8883,N_8789,N_8095);
xor U8884 (N_8884,N_8710,N_8742);
nor U8885 (N_8885,N_8641,N_8232);
nand U8886 (N_8886,N_8013,N_8520);
and U8887 (N_8887,N_8546,N_8485);
or U8888 (N_8888,N_8007,N_8147);
and U8889 (N_8889,N_8116,N_8631);
xor U8890 (N_8890,N_8014,N_8438);
and U8891 (N_8891,N_8401,N_8160);
or U8892 (N_8892,N_8016,N_8104);
or U8893 (N_8893,N_8292,N_8043);
and U8894 (N_8894,N_8324,N_8547);
nand U8895 (N_8895,N_8646,N_8313);
nor U8896 (N_8896,N_8602,N_8056);
xnor U8897 (N_8897,N_8375,N_8466);
and U8898 (N_8898,N_8307,N_8728);
nand U8899 (N_8899,N_8035,N_8031);
nor U8900 (N_8900,N_8491,N_8155);
nand U8901 (N_8901,N_8595,N_8526);
nand U8902 (N_8902,N_8241,N_8799);
xnor U8903 (N_8903,N_8027,N_8063);
nor U8904 (N_8904,N_8794,N_8629);
or U8905 (N_8905,N_8705,N_8020);
xnor U8906 (N_8906,N_8477,N_8347);
xnor U8907 (N_8907,N_8276,N_8138);
nor U8908 (N_8908,N_8018,N_8096);
nor U8909 (N_8909,N_8159,N_8412);
and U8910 (N_8910,N_8768,N_8442);
nand U8911 (N_8911,N_8461,N_8113);
and U8912 (N_8912,N_8533,N_8077);
nor U8913 (N_8913,N_8225,N_8655);
and U8914 (N_8914,N_8772,N_8474);
xor U8915 (N_8915,N_8779,N_8355);
xnor U8916 (N_8916,N_8215,N_8525);
and U8917 (N_8917,N_8123,N_8673);
and U8918 (N_8918,N_8248,N_8572);
nor U8919 (N_8919,N_8311,N_8314);
xor U8920 (N_8920,N_8763,N_8177);
nor U8921 (N_8921,N_8187,N_8224);
or U8922 (N_8922,N_8496,N_8699);
nand U8923 (N_8923,N_8499,N_8108);
and U8924 (N_8924,N_8380,N_8605);
and U8925 (N_8925,N_8410,N_8701);
or U8926 (N_8926,N_8238,N_8744);
nor U8927 (N_8927,N_8091,N_8227);
xor U8928 (N_8928,N_8269,N_8207);
nand U8929 (N_8929,N_8251,N_8395);
and U8930 (N_8930,N_8760,N_8444);
nand U8931 (N_8931,N_8599,N_8274);
nor U8932 (N_8932,N_8634,N_8246);
nor U8933 (N_8933,N_8777,N_8217);
xnor U8934 (N_8934,N_8747,N_8745);
nor U8935 (N_8935,N_8394,N_8539);
xnor U8936 (N_8936,N_8709,N_8361);
and U8937 (N_8937,N_8134,N_8642);
or U8938 (N_8938,N_8212,N_8695);
nor U8939 (N_8939,N_8128,N_8073);
nand U8940 (N_8940,N_8229,N_8233);
nor U8941 (N_8941,N_8790,N_8284);
nand U8942 (N_8942,N_8344,N_8237);
or U8943 (N_8943,N_8079,N_8360);
or U8944 (N_8944,N_8687,N_8666);
nand U8945 (N_8945,N_8069,N_8203);
nand U8946 (N_8946,N_8716,N_8791);
xor U8947 (N_8947,N_8544,N_8211);
and U8948 (N_8948,N_8738,N_8103);
xor U8949 (N_8949,N_8068,N_8718);
nor U8950 (N_8950,N_8500,N_8693);
xnor U8951 (N_8951,N_8426,N_8508);
and U8952 (N_8952,N_8149,N_8268);
and U8953 (N_8953,N_8329,N_8282);
xor U8954 (N_8954,N_8601,N_8487);
xor U8955 (N_8955,N_8332,N_8338);
or U8956 (N_8956,N_8540,N_8182);
nor U8957 (N_8957,N_8130,N_8144);
nor U8958 (N_8958,N_8316,N_8737);
and U8959 (N_8959,N_8471,N_8451);
nor U8960 (N_8960,N_8099,N_8189);
nand U8961 (N_8961,N_8377,N_8354);
nor U8962 (N_8962,N_8796,N_8383);
xor U8963 (N_8963,N_8058,N_8222);
xnor U8964 (N_8964,N_8290,N_8141);
nor U8965 (N_8965,N_8659,N_8357);
xnor U8966 (N_8966,N_8735,N_8021);
nand U8967 (N_8967,N_8076,N_8370);
nor U8968 (N_8968,N_8792,N_8449);
and U8969 (N_8969,N_8534,N_8102);
xor U8970 (N_8970,N_8170,N_8455);
xor U8971 (N_8971,N_8702,N_8511);
or U8972 (N_8972,N_8584,N_8258);
and U8973 (N_8973,N_8618,N_8093);
xnor U8974 (N_8974,N_8242,N_8543);
xnor U8975 (N_8975,N_8721,N_8483);
and U8976 (N_8976,N_8783,N_8715);
and U8977 (N_8977,N_8032,N_8517);
xor U8978 (N_8978,N_8122,N_8202);
xnor U8979 (N_8979,N_8503,N_8530);
or U8980 (N_8980,N_8367,N_8044);
nor U8981 (N_8981,N_8468,N_8720);
xor U8982 (N_8982,N_8771,N_8011);
nor U8983 (N_8983,N_8691,N_8486);
and U8984 (N_8984,N_8411,N_8059);
xor U8985 (N_8985,N_8397,N_8341);
and U8986 (N_8986,N_8643,N_8061);
nand U8987 (N_8987,N_8392,N_8550);
nand U8988 (N_8988,N_8664,N_8132);
nor U8989 (N_8989,N_8741,N_8594);
nor U8990 (N_8990,N_8405,N_8769);
xnor U8991 (N_8991,N_8271,N_8425);
nand U8992 (N_8992,N_8671,N_8243);
or U8993 (N_8993,N_8711,N_8226);
xnor U8994 (N_8994,N_8678,N_8041);
nor U8995 (N_8995,N_8610,N_8675);
xor U8996 (N_8996,N_8196,N_8033);
and U8997 (N_8997,N_8590,N_8683);
and U8998 (N_8998,N_8281,N_8545);
and U8999 (N_8999,N_8045,N_8681);
nand U9000 (N_9000,N_8739,N_8219);
or U9001 (N_9001,N_8030,N_8430);
or U9002 (N_9002,N_8775,N_8188);
and U9003 (N_9003,N_8300,N_8071);
nor U9004 (N_9004,N_8793,N_8275);
nor U9005 (N_9005,N_8327,N_8110);
nand U9006 (N_9006,N_8684,N_8023);
nand U9007 (N_9007,N_8621,N_8598);
xor U9008 (N_9008,N_8404,N_8630);
nor U9009 (N_9009,N_8053,N_8501);
xor U9010 (N_9010,N_8107,N_8084);
and U9011 (N_9011,N_8432,N_8596);
nand U9012 (N_9012,N_8349,N_8585);
or U9013 (N_9013,N_8351,N_8786);
xnor U9014 (N_9014,N_8400,N_8176);
and U9015 (N_9015,N_8169,N_8644);
nor U9016 (N_9016,N_8555,N_8434);
and U9017 (N_9017,N_8039,N_8105);
and U9018 (N_9018,N_8012,N_8797);
nand U9019 (N_9019,N_8690,N_8565);
xor U9020 (N_9020,N_8542,N_8163);
nor U9021 (N_9021,N_8459,N_8389);
and U9022 (N_9022,N_8453,N_8239);
nand U9023 (N_9023,N_8206,N_8247);
xor U9024 (N_9024,N_8139,N_8352);
nor U9025 (N_9025,N_8175,N_8607);
and U9026 (N_9026,N_8713,N_8460);
or U9027 (N_9027,N_8181,N_8310);
and U9028 (N_9028,N_8272,N_8552);
nor U9029 (N_9029,N_8733,N_8649);
and U9030 (N_9030,N_8632,N_8443);
nand U9031 (N_9031,N_8078,N_8376);
or U9032 (N_9032,N_8415,N_8256);
nand U9033 (N_9033,N_8153,N_8296);
nor U9034 (N_9034,N_8364,N_8346);
nor U9035 (N_9035,N_8454,N_8119);
nand U9036 (N_9036,N_8617,N_8578);
and U9037 (N_9037,N_8234,N_8467);
nor U9038 (N_9038,N_8563,N_8158);
and U9039 (N_9039,N_8682,N_8577);
and U9040 (N_9040,N_8650,N_8278);
xnor U9041 (N_9041,N_8515,N_8788);
and U9042 (N_9042,N_8047,N_8216);
nor U9043 (N_9043,N_8450,N_8746);
or U9044 (N_9044,N_8672,N_8723);
and U9045 (N_9045,N_8480,N_8692);
nand U9046 (N_9046,N_8731,N_8494);
nor U9047 (N_9047,N_8117,N_8529);
and U9048 (N_9048,N_8179,N_8365);
nand U9049 (N_9049,N_8145,N_8764);
nand U9050 (N_9050,N_8362,N_8497);
nand U9051 (N_9051,N_8722,N_8009);
xnor U9052 (N_9052,N_8088,N_8350);
nand U9053 (N_9053,N_8512,N_8437);
and U9054 (N_9054,N_8560,N_8255);
nor U9055 (N_9055,N_8253,N_8121);
nand U9056 (N_9056,N_8263,N_8082);
xnor U9057 (N_9057,N_8667,N_8502);
nor U9058 (N_9058,N_8537,N_8299);
nand U9059 (N_9059,N_8785,N_8050);
nor U9060 (N_9060,N_8172,N_8120);
nor U9061 (N_9061,N_8509,N_8024);
nor U9062 (N_9062,N_8051,N_8773);
nor U9063 (N_9063,N_8042,N_8291);
nor U9064 (N_9064,N_8293,N_8106);
nor U9065 (N_9065,N_8257,N_8262);
or U9066 (N_9066,N_8195,N_8005);
nand U9067 (N_9067,N_8782,N_8245);
nand U9068 (N_9068,N_8067,N_8331);
nor U9069 (N_9069,N_8597,N_8562);
and U9070 (N_9070,N_8317,N_8055);
and U9071 (N_9071,N_8345,N_8575);
xnor U9072 (N_9072,N_8066,N_8479);
nand U9073 (N_9073,N_8532,N_8574);
xnor U9074 (N_9074,N_8531,N_8685);
nor U9075 (N_9075,N_8127,N_8408);
or U9076 (N_9076,N_8571,N_8228);
and U9077 (N_9077,N_8090,N_8703);
nand U9078 (N_9078,N_8171,N_8416);
or U9079 (N_9079,N_8759,N_8087);
or U9080 (N_9080,N_8640,N_8427);
nor U9081 (N_9081,N_8441,N_8320);
and U9082 (N_9082,N_8614,N_8339);
nand U9083 (N_9083,N_8034,N_8200);
or U9084 (N_9084,N_8191,N_8704);
nor U9085 (N_9085,N_8457,N_8637);
or U9086 (N_9086,N_8638,N_8109);
and U9087 (N_9087,N_8240,N_8743);
nor U9088 (N_9088,N_8421,N_8165);
nand U9089 (N_9089,N_8554,N_8472);
and U9090 (N_9090,N_8573,N_8725);
nand U9091 (N_9091,N_8326,N_8767);
and U9092 (N_9092,N_8201,N_8463);
and U9093 (N_9093,N_8403,N_8636);
or U9094 (N_9094,N_8514,N_8436);
or U9095 (N_9095,N_8213,N_8288);
nand U9096 (N_9096,N_8002,N_8689);
and U9097 (N_9097,N_8148,N_8538);
nand U9098 (N_9098,N_8214,N_8186);
xor U9099 (N_9099,N_8627,N_8135);
xnor U9100 (N_9100,N_8518,N_8727);
nand U9101 (N_9101,N_8340,N_8669);
nand U9102 (N_9102,N_8398,N_8178);
nand U9103 (N_9103,N_8688,N_8083);
or U9104 (N_9104,N_8513,N_8006);
and U9105 (N_9105,N_8423,N_8452);
nor U9106 (N_9106,N_8440,N_8335);
or U9107 (N_9107,N_8231,N_8037);
xor U9108 (N_9108,N_8591,N_8516);
and U9109 (N_9109,N_8420,N_8611);
nand U9110 (N_9110,N_8566,N_8000);
and U9111 (N_9111,N_8765,N_8564);
nand U9112 (N_9112,N_8418,N_8008);
nand U9113 (N_9113,N_8780,N_8665);
or U9114 (N_9114,N_8004,N_8125);
and U9115 (N_9115,N_8615,N_8321);
nand U9116 (N_9116,N_8301,N_8527);
and U9117 (N_9117,N_8536,N_8010);
and U9118 (N_9118,N_8363,N_8287);
or U9119 (N_9119,N_8579,N_8157);
or U9120 (N_9120,N_8285,N_8267);
nand U9121 (N_9121,N_8322,N_8366);
nor U9122 (N_9122,N_8399,N_8755);
xor U9123 (N_9123,N_8305,N_8054);
nor U9124 (N_9124,N_8129,N_8065);
nand U9125 (N_9125,N_8333,N_8336);
or U9126 (N_9126,N_8456,N_8724);
and U9127 (N_9127,N_8374,N_8749);
and U9128 (N_9128,N_8019,N_8173);
and U9129 (N_9129,N_8589,N_8469);
nor U9130 (N_9130,N_8535,N_8569);
nor U9131 (N_9131,N_8040,N_8210);
and U9132 (N_9132,N_8726,N_8609);
nand U9133 (N_9133,N_8294,N_8371);
xnor U9134 (N_9134,N_8484,N_8085);
xor U9135 (N_9135,N_8387,N_8696);
or U9136 (N_9136,N_8359,N_8656);
nor U9137 (N_9137,N_8470,N_8003);
nor U9138 (N_9138,N_8094,N_8729);
xor U9139 (N_9139,N_8180,N_8343);
nand U9140 (N_9140,N_8493,N_8795);
nand U9141 (N_9141,N_8608,N_8198);
nand U9142 (N_9142,N_8424,N_8592);
nand U9143 (N_9143,N_8379,N_8422);
or U9144 (N_9144,N_8697,N_8097);
xor U9145 (N_9145,N_8124,N_8465);
nor U9146 (N_9146,N_8458,N_8706);
nand U9147 (N_9147,N_8524,N_8325);
nand U9148 (N_9148,N_8252,N_8679);
and U9149 (N_9149,N_8750,N_8447);
xor U9150 (N_9150,N_8587,N_8164);
and U9151 (N_9151,N_8700,N_8197);
nand U9152 (N_9152,N_8462,N_8712);
nor U9153 (N_9153,N_8549,N_8184);
xnor U9154 (N_9154,N_8378,N_8136);
xor U9155 (N_9155,N_8717,N_8261);
xnor U9156 (N_9156,N_8092,N_8548);
nand U9157 (N_9157,N_8628,N_8414);
nor U9158 (N_9158,N_8022,N_8036);
nand U9159 (N_9159,N_8060,N_8504);
or U9160 (N_9160,N_8072,N_8358);
nand U9161 (N_9161,N_8787,N_8654);
and U9162 (N_9162,N_8752,N_8115);
nand U9163 (N_9163,N_8475,N_8612);
xnor U9164 (N_9164,N_8194,N_8620);
xnor U9165 (N_9165,N_8209,N_8381);
and U9166 (N_9166,N_8137,N_8015);
nor U9167 (N_9167,N_8489,N_8433);
and U9168 (N_9168,N_8167,N_8393);
xnor U9169 (N_9169,N_8770,N_8583);
or U9170 (N_9170,N_8707,N_8558);
and U9171 (N_9171,N_8732,N_8784);
nand U9172 (N_9172,N_8626,N_8118);
nor U9173 (N_9173,N_8062,N_8086);
or U9174 (N_9174,N_8193,N_8048);
or U9175 (N_9175,N_8523,N_8356);
nand U9176 (N_9176,N_8557,N_8446);
nand U9177 (N_9177,N_8391,N_8100);
nand U9178 (N_9178,N_8046,N_8619);
or U9179 (N_9179,N_8645,N_8754);
xor U9180 (N_9180,N_8111,N_8429);
nor U9181 (N_9181,N_8266,N_8279);
and U9182 (N_9182,N_8199,N_8081);
nor U9183 (N_9183,N_8407,N_8781);
nand U9184 (N_9184,N_8488,N_8230);
and U9185 (N_9185,N_8218,N_8220);
nand U9186 (N_9186,N_8140,N_8318);
nand U9187 (N_9187,N_8244,N_8369);
or U9188 (N_9188,N_8289,N_8074);
nand U9189 (N_9189,N_8774,N_8286);
or U9190 (N_9190,N_8616,N_8417);
nor U9191 (N_9191,N_8505,N_8402);
and U9192 (N_9192,N_8694,N_8519);
xnor U9193 (N_9193,N_8236,N_8586);
and U9194 (N_9194,N_8660,N_8541);
and U9195 (N_9195,N_8652,N_8250);
nand U9196 (N_9196,N_8204,N_8390);
or U9197 (N_9197,N_8026,N_8490);
nand U9198 (N_9198,N_8625,N_8613);
and U9199 (N_9199,N_8156,N_8651);
or U9200 (N_9200,N_8561,N_8659);
xnor U9201 (N_9201,N_8342,N_8679);
and U9202 (N_9202,N_8111,N_8401);
xor U9203 (N_9203,N_8115,N_8339);
nor U9204 (N_9204,N_8158,N_8497);
nand U9205 (N_9205,N_8783,N_8144);
xor U9206 (N_9206,N_8154,N_8308);
and U9207 (N_9207,N_8096,N_8217);
or U9208 (N_9208,N_8114,N_8052);
nand U9209 (N_9209,N_8661,N_8238);
nand U9210 (N_9210,N_8548,N_8459);
or U9211 (N_9211,N_8691,N_8331);
and U9212 (N_9212,N_8494,N_8785);
nand U9213 (N_9213,N_8542,N_8504);
nand U9214 (N_9214,N_8425,N_8226);
and U9215 (N_9215,N_8699,N_8482);
nand U9216 (N_9216,N_8170,N_8772);
nand U9217 (N_9217,N_8360,N_8608);
nand U9218 (N_9218,N_8484,N_8444);
or U9219 (N_9219,N_8475,N_8793);
xor U9220 (N_9220,N_8521,N_8780);
and U9221 (N_9221,N_8655,N_8635);
xor U9222 (N_9222,N_8538,N_8686);
nor U9223 (N_9223,N_8330,N_8767);
xor U9224 (N_9224,N_8124,N_8694);
nor U9225 (N_9225,N_8634,N_8730);
and U9226 (N_9226,N_8761,N_8303);
nor U9227 (N_9227,N_8751,N_8212);
and U9228 (N_9228,N_8419,N_8096);
or U9229 (N_9229,N_8088,N_8019);
nand U9230 (N_9230,N_8530,N_8316);
nand U9231 (N_9231,N_8145,N_8796);
or U9232 (N_9232,N_8675,N_8312);
and U9233 (N_9233,N_8040,N_8070);
or U9234 (N_9234,N_8560,N_8205);
xor U9235 (N_9235,N_8096,N_8559);
nand U9236 (N_9236,N_8579,N_8471);
or U9237 (N_9237,N_8688,N_8101);
nor U9238 (N_9238,N_8300,N_8740);
nand U9239 (N_9239,N_8606,N_8397);
nor U9240 (N_9240,N_8298,N_8016);
nand U9241 (N_9241,N_8581,N_8373);
and U9242 (N_9242,N_8082,N_8783);
xor U9243 (N_9243,N_8016,N_8696);
nand U9244 (N_9244,N_8255,N_8570);
or U9245 (N_9245,N_8374,N_8764);
and U9246 (N_9246,N_8051,N_8746);
nor U9247 (N_9247,N_8250,N_8679);
or U9248 (N_9248,N_8410,N_8033);
and U9249 (N_9249,N_8119,N_8740);
xnor U9250 (N_9250,N_8719,N_8590);
nand U9251 (N_9251,N_8769,N_8644);
xnor U9252 (N_9252,N_8289,N_8147);
or U9253 (N_9253,N_8258,N_8209);
and U9254 (N_9254,N_8012,N_8104);
or U9255 (N_9255,N_8368,N_8763);
or U9256 (N_9256,N_8037,N_8219);
and U9257 (N_9257,N_8556,N_8626);
and U9258 (N_9258,N_8301,N_8484);
xor U9259 (N_9259,N_8243,N_8579);
xor U9260 (N_9260,N_8439,N_8258);
and U9261 (N_9261,N_8138,N_8645);
nand U9262 (N_9262,N_8265,N_8301);
and U9263 (N_9263,N_8727,N_8720);
nor U9264 (N_9264,N_8470,N_8733);
or U9265 (N_9265,N_8254,N_8788);
and U9266 (N_9266,N_8016,N_8735);
and U9267 (N_9267,N_8377,N_8351);
or U9268 (N_9268,N_8694,N_8046);
and U9269 (N_9269,N_8639,N_8245);
nand U9270 (N_9270,N_8042,N_8422);
or U9271 (N_9271,N_8196,N_8746);
nor U9272 (N_9272,N_8452,N_8174);
xor U9273 (N_9273,N_8535,N_8663);
nor U9274 (N_9274,N_8084,N_8056);
or U9275 (N_9275,N_8522,N_8227);
nand U9276 (N_9276,N_8194,N_8099);
xnor U9277 (N_9277,N_8492,N_8561);
or U9278 (N_9278,N_8519,N_8149);
xnor U9279 (N_9279,N_8157,N_8728);
nand U9280 (N_9280,N_8089,N_8315);
xnor U9281 (N_9281,N_8508,N_8400);
and U9282 (N_9282,N_8497,N_8736);
or U9283 (N_9283,N_8473,N_8297);
and U9284 (N_9284,N_8045,N_8314);
and U9285 (N_9285,N_8051,N_8527);
and U9286 (N_9286,N_8480,N_8753);
nand U9287 (N_9287,N_8799,N_8147);
xor U9288 (N_9288,N_8659,N_8432);
or U9289 (N_9289,N_8174,N_8111);
nor U9290 (N_9290,N_8642,N_8252);
nand U9291 (N_9291,N_8498,N_8323);
nand U9292 (N_9292,N_8704,N_8108);
xor U9293 (N_9293,N_8181,N_8315);
or U9294 (N_9294,N_8324,N_8475);
or U9295 (N_9295,N_8786,N_8062);
nand U9296 (N_9296,N_8307,N_8679);
or U9297 (N_9297,N_8347,N_8125);
nand U9298 (N_9298,N_8073,N_8174);
nand U9299 (N_9299,N_8328,N_8251);
nand U9300 (N_9300,N_8571,N_8793);
xnor U9301 (N_9301,N_8202,N_8292);
nor U9302 (N_9302,N_8069,N_8555);
xor U9303 (N_9303,N_8433,N_8286);
nand U9304 (N_9304,N_8547,N_8056);
nor U9305 (N_9305,N_8238,N_8050);
nand U9306 (N_9306,N_8716,N_8252);
or U9307 (N_9307,N_8043,N_8481);
and U9308 (N_9308,N_8124,N_8711);
nor U9309 (N_9309,N_8382,N_8555);
xor U9310 (N_9310,N_8175,N_8316);
nand U9311 (N_9311,N_8661,N_8106);
or U9312 (N_9312,N_8047,N_8431);
or U9313 (N_9313,N_8775,N_8791);
xor U9314 (N_9314,N_8788,N_8346);
nor U9315 (N_9315,N_8780,N_8580);
nor U9316 (N_9316,N_8411,N_8405);
or U9317 (N_9317,N_8772,N_8737);
xnor U9318 (N_9318,N_8497,N_8291);
nand U9319 (N_9319,N_8222,N_8257);
and U9320 (N_9320,N_8667,N_8467);
nand U9321 (N_9321,N_8542,N_8441);
nand U9322 (N_9322,N_8665,N_8773);
or U9323 (N_9323,N_8636,N_8551);
nor U9324 (N_9324,N_8099,N_8623);
or U9325 (N_9325,N_8655,N_8681);
xnor U9326 (N_9326,N_8285,N_8503);
or U9327 (N_9327,N_8357,N_8095);
and U9328 (N_9328,N_8726,N_8713);
nand U9329 (N_9329,N_8052,N_8444);
xor U9330 (N_9330,N_8162,N_8665);
nand U9331 (N_9331,N_8166,N_8047);
and U9332 (N_9332,N_8449,N_8266);
nand U9333 (N_9333,N_8041,N_8167);
or U9334 (N_9334,N_8034,N_8273);
xnor U9335 (N_9335,N_8581,N_8467);
or U9336 (N_9336,N_8328,N_8136);
xor U9337 (N_9337,N_8749,N_8198);
xor U9338 (N_9338,N_8198,N_8241);
xnor U9339 (N_9339,N_8685,N_8136);
nor U9340 (N_9340,N_8257,N_8514);
xor U9341 (N_9341,N_8722,N_8786);
nor U9342 (N_9342,N_8045,N_8499);
nor U9343 (N_9343,N_8337,N_8513);
nand U9344 (N_9344,N_8759,N_8260);
nor U9345 (N_9345,N_8159,N_8490);
and U9346 (N_9346,N_8796,N_8724);
nand U9347 (N_9347,N_8020,N_8726);
xnor U9348 (N_9348,N_8202,N_8142);
and U9349 (N_9349,N_8140,N_8774);
xor U9350 (N_9350,N_8552,N_8573);
and U9351 (N_9351,N_8144,N_8668);
and U9352 (N_9352,N_8215,N_8378);
and U9353 (N_9353,N_8160,N_8459);
and U9354 (N_9354,N_8277,N_8634);
nor U9355 (N_9355,N_8084,N_8581);
and U9356 (N_9356,N_8184,N_8088);
nand U9357 (N_9357,N_8628,N_8033);
nor U9358 (N_9358,N_8789,N_8679);
or U9359 (N_9359,N_8120,N_8515);
and U9360 (N_9360,N_8798,N_8243);
nor U9361 (N_9361,N_8215,N_8457);
xnor U9362 (N_9362,N_8793,N_8760);
or U9363 (N_9363,N_8506,N_8488);
nand U9364 (N_9364,N_8302,N_8041);
and U9365 (N_9365,N_8040,N_8377);
nand U9366 (N_9366,N_8400,N_8530);
xnor U9367 (N_9367,N_8730,N_8033);
xnor U9368 (N_9368,N_8047,N_8386);
or U9369 (N_9369,N_8103,N_8150);
nor U9370 (N_9370,N_8314,N_8399);
nand U9371 (N_9371,N_8330,N_8425);
and U9372 (N_9372,N_8183,N_8118);
xnor U9373 (N_9373,N_8640,N_8782);
or U9374 (N_9374,N_8620,N_8475);
or U9375 (N_9375,N_8326,N_8743);
xnor U9376 (N_9376,N_8314,N_8363);
nand U9377 (N_9377,N_8008,N_8232);
nor U9378 (N_9378,N_8306,N_8402);
and U9379 (N_9379,N_8443,N_8355);
nor U9380 (N_9380,N_8422,N_8710);
nor U9381 (N_9381,N_8316,N_8583);
and U9382 (N_9382,N_8215,N_8571);
or U9383 (N_9383,N_8480,N_8793);
nor U9384 (N_9384,N_8186,N_8372);
nand U9385 (N_9385,N_8748,N_8387);
xor U9386 (N_9386,N_8017,N_8076);
nor U9387 (N_9387,N_8311,N_8002);
xnor U9388 (N_9388,N_8552,N_8738);
xor U9389 (N_9389,N_8530,N_8261);
xor U9390 (N_9390,N_8000,N_8236);
nand U9391 (N_9391,N_8794,N_8123);
nand U9392 (N_9392,N_8153,N_8134);
xor U9393 (N_9393,N_8760,N_8696);
nand U9394 (N_9394,N_8673,N_8137);
nor U9395 (N_9395,N_8280,N_8612);
nor U9396 (N_9396,N_8756,N_8777);
xor U9397 (N_9397,N_8340,N_8422);
xor U9398 (N_9398,N_8113,N_8223);
and U9399 (N_9399,N_8400,N_8472);
or U9400 (N_9400,N_8011,N_8449);
and U9401 (N_9401,N_8109,N_8314);
and U9402 (N_9402,N_8404,N_8740);
nand U9403 (N_9403,N_8269,N_8507);
and U9404 (N_9404,N_8601,N_8050);
xor U9405 (N_9405,N_8434,N_8185);
or U9406 (N_9406,N_8500,N_8328);
or U9407 (N_9407,N_8787,N_8015);
and U9408 (N_9408,N_8019,N_8115);
xnor U9409 (N_9409,N_8253,N_8743);
nand U9410 (N_9410,N_8746,N_8161);
nor U9411 (N_9411,N_8449,N_8412);
or U9412 (N_9412,N_8465,N_8542);
or U9413 (N_9413,N_8303,N_8638);
nor U9414 (N_9414,N_8674,N_8270);
or U9415 (N_9415,N_8414,N_8355);
nand U9416 (N_9416,N_8584,N_8396);
nor U9417 (N_9417,N_8434,N_8652);
and U9418 (N_9418,N_8545,N_8139);
and U9419 (N_9419,N_8594,N_8722);
or U9420 (N_9420,N_8233,N_8243);
nor U9421 (N_9421,N_8717,N_8744);
nor U9422 (N_9422,N_8554,N_8191);
nor U9423 (N_9423,N_8282,N_8606);
nand U9424 (N_9424,N_8428,N_8457);
or U9425 (N_9425,N_8415,N_8405);
nor U9426 (N_9426,N_8629,N_8393);
xor U9427 (N_9427,N_8084,N_8275);
nand U9428 (N_9428,N_8323,N_8167);
xor U9429 (N_9429,N_8610,N_8005);
and U9430 (N_9430,N_8510,N_8312);
nor U9431 (N_9431,N_8249,N_8158);
xnor U9432 (N_9432,N_8610,N_8076);
or U9433 (N_9433,N_8336,N_8760);
and U9434 (N_9434,N_8306,N_8049);
nor U9435 (N_9435,N_8035,N_8713);
xor U9436 (N_9436,N_8599,N_8442);
nand U9437 (N_9437,N_8353,N_8679);
nor U9438 (N_9438,N_8715,N_8291);
nor U9439 (N_9439,N_8581,N_8472);
xor U9440 (N_9440,N_8248,N_8047);
nand U9441 (N_9441,N_8015,N_8149);
nand U9442 (N_9442,N_8530,N_8794);
nor U9443 (N_9443,N_8209,N_8295);
or U9444 (N_9444,N_8240,N_8562);
xnor U9445 (N_9445,N_8472,N_8704);
and U9446 (N_9446,N_8613,N_8118);
xnor U9447 (N_9447,N_8460,N_8137);
and U9448 (N_9448,N_8024,N_8640);
nor U9449 (N_9449,N_8615,N_8383);
nand U9450 (N_9450,N_8563,N_8318);
nor U9451 (N_9451,N_8308,N_8110);
and U9452 (N_9452,N_8149,N_8653);
and U9453 (N_9453,N_8036,N_8429);
nand U9454 (N_9454,N_8423,N_8331);
xnor U9455 (N_9455,N_8049,N_8595);
and U9456 (N_9456,N_8571,N_8341);
nand U9457 (N_9457,N_8369,N_8754);
nor U9458 (N_9458,N_8408,N_8447);
nand U9459 (N_9459,N_8060,N_8680);
or U9460 (N_9460,N_8332,N_8053);
and U9461 (N_9461,N_8243,N_8755);
xnor U9462 (N_9462,N_8519,N_8314);
xor U9463 (N_9463,N_8568,N_8565);
or U9464 (N_9464,N_8040,N_8397);
nand U9465 (N_9465,N_8550,N_8428);
or U9466 (N_9466,N_8490,N_8129);
or U9467 (N_9467,N_8758,N_8768);
nand U9468 (N_9468,N_8003,N_8417);
nand U9469 (N_9469,N_8355,N_8516);
nand U9470 (N_9470,N_8752,N_8730);
nand U9471 (N_9471,N_8578,N_8769);
or U9472 (N_9472,N_8217,N_8622);
nor U9473 (N_9473,N_8283,N_8172);
xor U9474 (N_9474,N_8205,N_8143);
nand U9475 (N_9475,N_8548,N_8664);
nand U9476 (N_9476,N_8177,N_8650);
and U9477 (N_9477,N_8181,N_8061);
xor U9478 (N_9478,N_8363,N_8534);
or U9479 (N_9479,N_8285,N_8659);
nor U9480 (N_9480,N_8481,N_8427);
nand U9481 (N_9481,N_8430,N_8746);
or U9482 (N_9482,N_8712,N_8007);
and U9483 (N_9483,N_8451,N_8232);
nor U9484 (N_9484,N_8216,N_8635);
nor U9485 (N_9485,N_8533,N_8073);
xnor U9486 (N_9486,N_8701,N_8044);
and U9487 (N_9487,N_8064,N_8717);
and U9488 (N_9488,N_8754,N_8065);
or U9489 (N_9489,N_8675,N_8234);
nand U9490 (N_9490,N_8586,N_8563);
and U9491 (N_9491,N_8235,N_8634);
and U9492 (N_9492,N_8053,N_8536);
xor U9493 (N_9493,N_8651,N_8561);
xnor U9494 (N_9494,N_8575,N_8299);
or U9495 (N_9495,N_8279,N_8052);
nor U9496 (N_9496,N_8160,N_8249);
or U9497 (N_9497,N_8748,N_8089);
and U9498 (N_9498,N_8567,N_8641);
nand U9499 (N_9499,N_8039,N_8433);
or U9500 (N_9500,N_8419,N_8470);
nor U9501 (N_9501,N_8679,N_8149);
and U9502 (N_9502,N_8194,N_8040);
nand U9503 (N_9503,N_8013,N_8449);
and U9504 (N_9504,N_8029,N_8423);
or U9505 (N_9505,N_8560,N_8796);
nor U9506 (N_9506,N_8447,N_8085);
or U9507 (N_9507,N_8670,N_8351);
nor U9508 (N_9508,N_8325,N_8516);
xnor U9509 (N_9509,N_8365,N_8688);
or U9510 (N_9510,N_8451,N_8212);
or U9511 (N_9511,N_8741,N_8082);
xnor U9512 (N_9512,N_8463,N_8539);
nor U9513 (N_9513,N_8557,N_8296);
or U9514 (N_9514,N_8567,N_8786);
and U9515 (N_9515,N_8783,N_8175);
or U9516 (N_9516,N_8025,N_8275);
and U9517 (N_9517,N_8618,N_8780);
or U9518 (N_9518,N_8009,N_8331);
xor U9519 (N_9519,N_8378,N_8757);
xnor U9520 (N_9520,N_8202,N_8279);
and U9521 (N_9521,N_8141,N_8764);
xnor U9522 (N_9522,N_8231,N_8719);
or U9523 (N_9523,N_8279,N_8183);
xor U9524 (N_9524,N_8527,N_8225);
nor U9525 (N_9525,N_8052,N_8782);
and U9526 (N_9526,N_8739,N_8005);
nor U9527 (N_9527,N_8160,N_8730);
nor U9528 (N_9528,N_8290,N_8412);
and U9529 (N_9529,N_8615,N_8084);
xor U9530 (N_9530,N_8297,N_8013);
or U9531 (N_9531,N_8125,N_8001);
xnor U9532 (N_9532,N_8383,N_8168);
xor U9533 (N_9533,N_8027,N_8799);
and U9534 (N_9534,N_8558,N_8082);
xor U9535 (N_9535,N_8000,N_8532);
nor U9536 (N_9536,N_8798,N_8374);
xor U9537 (N_9537,N_8386,N_8212);
nor U9538 (N_9538,N_8458,N_8763);
nor U9539 (N_9539,N_8515,N_8367);
nor U9540 (N_9540,N_8214,N_8057);
xnor U9541 (N_9541,N_8748,N_8498);
and U9542 (N_9542,N_8424,N_8722);
or U9543 (N_9543,N_8695,N_8756);
xor U9544 (N_9544,N_8796,N_8143);
nor U9545 (N_9545,N_8459,N_8580);
nor U9546 (N_9546,N_8666,N_8475);
nor U9547 (N_9547,N_8160,N_8733);
and U9548 (N_9548,N_8441,N_8691);
xor U9549 (N_9549,N_8703,N_8265);
and U9550 (N_9550,N_8713,N_8782);
nand U9551 (N_9551,N_8129,N_8399);
or U9552 (N_9552,N_8007,N_8609);
and U9553 (N_9553,N_8372,N_8481);
and U9554 (N_9554,N_8096,N_8389);
xnor U9555 (N_9555,N_8203,N_8470);
or U9556 (N_9556,N_8442,N_8566);
nor U9557 (N_9557,N_8730,N_8789);
nor U9558 (N_9558,N_8658,N_8738);
and U9559 (N_9559,N_8587,N_8134);
xnor U9560 (N_9560,N_8717,N_8745);
xor U9561 (N_9561,N_8713,N_8287);
nand U9562 (N_9562,N_8085,N_8142);
and U9563 (N_9563,N_8437,N_8778);
xor U9564 (N_9564,N_8662,N_8760);
and U9565 (N_9565,N_8364,N_8004);
xnor U9566 (N_9566,N_8228,N_8006);
or U9567 (N_9567,N_8636,N_8053);
and U9568 (N_9568,N_8220,N_8711);
nor U9569 (N_9569,N_8742,N_8736);
nand U9570 (N_9570,N_8041,N_8611);
nand U9571 (N_9571,N_8352,N_8025);
nand U9572 (N_9572,N_8165,N_8194);
nand U9573 (N_9573,N_8245,N_8163);
nor U9574 (N_9574,N_8642,N_8387);
and U9575 (N_9575,N_8061,N_8326);
nor U9576 (N_9576,N_8262,N_8454);
nand U9577 (N_9577,N_8324,N_8080);
nand U9578 (N_9578,N_8672,N_8700);
and U9579 (N_9579,N_8489,N_8255);
and U9580 (N_9580,N_8741,N_8162);
and U9581 (N_9581,N_8565,N_8046);
nand U9582 (N_9582,N_8092,N_8160);
and U9583 (N_9583,N_8613,N_8125);
and U9584 (N_9584,N_8431,N_8697);
xnor U9585 (N_9585,N_8697,N_8145);
nor U9586 (N_9586,N_8014,N_8224);
nor U9587 (N_9587,N_8323,N_8541);
and U9588 (N_9588,N_8054,N_8696);
nor U9589 (N_9589,N_8130,N_8158);
xnor U9590 (N_9590,N_8646,N_8669);
or U9591 (N_9591,N_8531,N_8755);
xnor U9592 (N_9592,N_8513,N_8003);
or U9593 (N_9593,N_8717,N_8599);
or U9594 (N_9594,N_8100,N_8617);
xnor U9595 (N_9595,N_8096,N_8070);
nor U9596 (N_9596,N_8230,N_8535);
nor U9597 (N_9597,N_8756,N_8232);
nor U9598 (N_9598,N_8154,N_8217);
or U9599 (N_9599,N_8390,N_8042);
and U9600 (N_9600,N_9509,N_8836);
nand U9601 (N_9601,N_8813,N_9190);
and U9602 (N_9602,N_9086,N_9236);
or U9603 (N_9603,N_9211,N_8973);
nand U9604 (N_9604,N_9201,N_9482);
nand U9605 (N_9605,N_9500,N_8966);
and U9606 (N_9606,N_9127,N_8829);
or U9607 (N_9607,N_8903,N_9251);
nor U9608 (N_9608,N_8939,N_9538);
and U9609 (N_9609,N_9252,N_9158);
and U9610 (N_9610,N_8875,N_8948);
nor U9611 (N_9611,N_9097,N_9392);
xor U9612 (N_9612,N_9167,N_9088);
nand U9613 (N_9613,N_8997,N_9147);
xor U9614 (N_9614,N_9273,N_9060);
and U9615 (N_9615,N_9467,N_8885);
and U9616 (N_9616,N_9434,N_9452);
nand U9617 (N_9617,N_8984,N_9476);
nor U9618 (N_9618,N_9094,N_9305);
and U9619 (N_9619,N_9474,N_9132);
nand U9620 (N_9620,N_9160,N_9488);
and U9621 (N_9621,N_9159,N_9485);
xnor U9622 (N_9622,N_9347,N_8932);
nor U9623 (N_9623,N_9085,N_9282);
and U9624 (N_9624,N_8860,N_9469);
nor U9625 (N_9625,N_9552,N_9002);
nand U9626 (N_9626,N_8857,N_8974);
xnor U9627 (N_9627,N_8808,N_9335);
nand U9628 (N_9628,N_9442,N_8917);
xnor U9629 (N_9629,N_8902,N_9243);
and U9630 (N_9630,N_9365,N_9134);
nor U9631 (N_9631,N_9143,N_8874);
and U9632 (N_9632,N_9173,N_9261);
or U9633 (N_9633,N_9334,N_8819);
xor U9634 (N_9634,N_9470,N_8924);
nand U9635 (N_9635,N_9383,N_9553);
and U9636 (N_9636,N_9116,N_9161);
and U9637 (N_9637,N_8823,N_9358);
xor U9638 (N_9638,N_9055,N_9399);
or U9639 (N_9639,N_9265,N_9397);
and U9640 (N_9640,N_8852,N_9585);
nand U9641 (N_9641,N_9458,N_9189);
or U9642 (N_9642,N_8834,N_8987);
nor U9643 (N_9643,N_8867,N_9306);
and U9644 (N_9644,N_8981,N_9440);
nor U9645 (N_9645,N_8806,N_9234);
nor U9646 (N_9646,N_8927,N_9247);
xnor U9647 (N_9647,N_9390,N_9516);
or U9648 (N_9648,N_9348,N_9572);
xnor U9649 (N_9649,N_9519,N_9180);
xor U9650 (N_9650,N_9249,N_9367);
xnor U9651 (N_9651,N_9491,N_8858);
and U9652 (N_9652,N_8950,N_9048);
and U9653 (N_9653,N_9130,N_9520);
nor U9654 (N_9654,N_9276,N_9402);
and U9655 (N_9655,N_8910,N_8863);
nand U9656 (N_9656,N_9256,N_9483);
xnor U9657 (N_9657,N_9414,N_9437);
nor U9658 (N_9658,N_9475,N_8810);
or U9659 (N_9659,N_8856,N_9576);
nor U9660 (N_9660,N_9394,N_9416);
nor U9661 (N_9661,N_9092,N_9341);
nor U9662 (N_9662,N_9340,N_8911);
and U9663 (N_9663,N_9217,N_9562);
or U9664 (N_9664,N_9037,N_9556);
xnor U9665 (N_9665,N_9121,N_9300);
xor U9666 (N_9666,N_8814,N_9494);
and U9667 (N_9667,N_8926,N_9559);
or U9668 (N_9668,N_9096,N_9209);
xnor U9669 (N_9669,N_9331,N_8989);
and U9670 (N_9670,N_9401,N_9408);
nand U9671 (N_9671,N_9487,N_8812);
xor U9672 (N_9672,N_9275,N_9356);
and U9673 (N_9673,N_9117,N_9035);
nand U9674 (N_9674,N_9398,N_9181);
or U9675 (N_9675,N_9326,N_9508);
xor U9676 (N_9676,N_9245,N_9110);
nor U9677 (N_9677,N_9449,N_9595);
or U9678 (N_9678,N_9468,N_9241);
xor U9679 (N_9679,N_9125,N_9281);
nand U9680 (N_9680,N_9566,N_9280);
or U9681 (N_9681,N_9030,N_9565);
and U9682 (N_9682,N_9304,N_8822);
or U9683 (N_9683,N_8871,N_9561);
xor U9684 (N_9684,N_8953,N_9598);
xor U9685 (N_9685,N_9391,N_8825);
nand U9686 (N_9686,N_9427,N_8805);
or U9687 (N_9687,N_8920,N_9202);
and U9688 (N_9688,N_9593,N_9316);
nor U9689 (N_9689,N_9428,N_9523);
nand U9690 (N_9690,N_9221,N_9345);
xor U9691 (N_9691,N_9518,N_9109);
or U9692 (N_9692,N_9283,N_9033);
and U9693 (N_9693,N_9011,N_8968);
nor U9694 (N_9694,N_9128,N_9270);
nor U9695 (N_9695,N_8892,N_9318);
xor U9696 (N_9696,N_9403,N_9235);
or U9697 (N_9697,N_9029,N_9406);
nor U9698 (N_9698,N_9082,N_9481);
nand U9699 (N_9699,N_9303,N_9596);
nand U9700 (N_9700,N_9286,N_9230);
and U9701 (N_9701,N_9302,N_9371);
nand U9702 (N_9702,N_9263,N_9266);
nor U9703 (N_9703,N_9580,N_8941);
or U9704 (N_9704,N_9239,N_9171);
or U9705 (N_9705,N_9050,N_8914);
nor U9706 (N_9706,N_9175,N_9226);
nand U9707 (N_9707,N_9176,N_9591);
xnor U9708 (N_9708,N_8821,N_9380);
and U9709 (N_9709,N_9400,N_8969);
xor U9710 (N_9710,N_9229,N_8832);
xor U9711 (N_9711,N_9438,N_9417);
xnor U9712 (N_9712,N_9207,N_9279);
or U9713 (N_9713,N_9444,N_9063);
nor U9714 (N_9714,N_9199,N_9289);
nor U9715 (N_9715,N_8846,N_9111);
or U9716 (N_9716,N_9351,N_9307);
and U9717 (N_9717,N_9079,N_9006);
or U9718 (N_9718,N_9095,N_9058);
nor U9719 (N_9719,N_8835,N_8986);
nand U9720 (N_9720,N_9373,N_9502);
nand U9721 (N_9721,N_9578,N_9000);
or U9722 (N_9722,N_9329,N_8942);
and U9723 (N_9723,N_9374,N_9203);
nand U9724 (N_9724,N_9536,N_9455);
and U9725 (N_9725,N_9407,N_9191);
xor U9726 (N_9726,N_9119,N_9216);
nor U9727 (N_9727,N_9013,N_9533);
nand U9728 (N_9728,N_8862,N_9459);
nand U9729 (N_9729,N_9232,N_8868);
and U9730 (N_9730,N_9075,N_9047);
and U9731 (N_9731,N_8853,N_9359);
nand U9732 (N_9732,N_9584,N_9010);
and U9733 (N_9733,N_8919,N_9321);
or U9734 (N_9734,N_9228,N_9569);
and U9735 (N_9735,N_8931,N_9140);
and U9736 (N_9736,N_9466,N_9511);
nor U9737 (N_9737,N_9100,N_9432);
nand U9738 (N_9738,N_9093,N_9457);
or U9739 (N_9739,N_9193,N_9368);
and U9740 (N_9740,N_8830,N_9162);
xnor U9741 (N_9741,N_9378,N_9142);
nand U9742 (N_9742,N_8965,N_9170);
or U9743 (N_9743,N_9376,N_9545);
and U9744 (N_9744,N_8881,N_9543);
nor U9745 (N_9745,N_8837,N_8958);
and U9746 (N_9746,N_9489,N_9113);
or U9747 (N_9747,N_9103,N_9053);
xor U9748 (N_9748,N_8933,N_9083);
xnor U9749 (N_9749,N_9138,N_9108);
or U9750 (N_9750,N_8886,N_9599);
nor U9751 (N_9751,N_8946,N_9168);
nor U9752 (N_9752,N_9114,N_9105);
or U9753 (N_9753,N_8955,N_8993);
and U9754 (N_9754,N_9024,N_9349);
nor U9755 (N_9755,N_9126,N_9573);
and U9756 (N_9756,N_8851,N_9453);
nand U9757 (N_9757,N_8901,N_9285);
xnor U9758 (N_9758,N_8807,N_9106);
xor U9759 (N_9759,N_9003,N_8930);
or U9760 (N_9760,N_8967,N_9311);
nor U9761 (N_9761,N_9152,N_9353);
xnor U9762 (N_9762,N_9194,N_9492);
or U9763 (N_9763,N_9074,N_9213);
and U9764 (N_9764,N_9587,N_9192);
xnor U9765 (N_9765,N_9278,N_9290);
nand U9766 (N_9766,N_9588,N_8957);
and U9767 (N_9767,N_9415,N_8938);
xnor U9768 (N_9768,N_9350,N_9393);
or U9769 (N_9769,N_9410,N_8944);
or U9770 (N_9770,N_9156,N_9594);
nand U9771 (N_9771,N_9522,N_9525);
and U9772 (N_9772,N_9429,N_9507);
xor U9773 (N_9773,N_9071,N_9515);
or U9774 (N_9774,N_9355,N_9412);
and U9775 (N_9775,N_9059,N_9541);
nand U9776 (N_9776,N_9505,N_8897);
and U9777 (N_9777,N_8859,N_9214);
xor U9778 (N_9778,N_8827,N_9436);
nand U9779 (N_9779,N_9342,N_9026);
nor U9780 (N_9780,N_9008,N_9527);
nor U9781 (N_9781,N_9395,N_9014);
nor U9782 (N_9782,N_9557,N_9233);
and U9783 (N_9783,N_9439,N_9589);
nand U9784 (N_9784,N_9555,N_9291);
xor U9785 (N_9785,N_9066,N_9090);
nor U9786 (N_9786,N_9568,N_9220);
nor U9787 (N_9787,N_9133,N_9041);
nand U9788 (N_9788,N_9366,N_9308);
and U9789 (N_9789,N_8870,N_9240);
or U9790 (N_9790,N_9043,N_9051);
xor U9791 (N_9791,N_9195,N_9313);
nand U9792 (N_9792,N_9069,N_9045);
or U9793 (N_9793,N_9582,N_9441);
nand U9794 (N_9794,N_9549,N_8865);
and U9795 (N_9795,N_8896,N_9091);
xor U9796 (N_9796,N_9567,N_9099);
xnor U9797 (N_9797,N_8880,N_8992);
nor U9798 (N_9798,N_9339,N_9430);
nand U9799 (N_9799,N_8884,N_9472);
and U9800 (N_9800,N_9284,N_8848);
and U9801 (N_9801,N_9295,N_9223);
xnor U9802 (N_9802,N_9361,N_9550);
xor U9803 (N_9803,N_8828,N_9163);
nand U9804 (N_9804,N_9465,N_9381);
xnor U9805 (N_9805,N_9179,N_9120);
nand U9806 (N_9806,N_9344,N_9477);
or U9807 (N_9807,N_9539,N_9293);
nor U9808 (N_9808,N_9040,N_9360);
or U9809 (N_9809,N_9149,N_9046);
or U9810 (N_9810,N_9362,N_9034);
and U9811 (N_9811,N_9486,N_9333);
xor U9812 (N_9812,N_9471,N_9150);
nor U9813 (N_9813,N_9309,N_9001);
nor U9814 (N_9814,N_9462,N_9418);
nand U9815 (N_9815,N_9148,N_9178);
nor U9816 (N_9816,N_8913,N_9205);
xor U9817 (N_9817,N_9153,N_9154);
or U9818 (N_9818,N_9583,N_9560);
nor U9819 (N_9819,N_9237,N_9253);
nand U9820 (N_9820,N_9107,N_9330);
nor U9821 (N_9821,N_9274,N_8899);
and U9822 (N_9822,N_9087,N_9445);
or U9823 (N_9823,N_8850,N_9165);
and U9824 (N_9824,N_9049,N_8929);
nand U9825 (N_9825,N_8925,N_9422);
nand U9826 (N_9826,N_9136,N_9548);
xor U9827 (N_9827,N_9254,N_9257);
or U9828 (N_9828,N_9218,N_9023);
nor U9829 (N_9829,N_9231,N_8954);
or U9830 (N_9830,N_8817,N_8908);
nand U9831 (N_9831,N_9077,N_8841);
and U9832 (N_9832,N_8869,N_8937);
and U9833 (N_9833,N_9346,N_8873);
xnor U9834 (N_9834,N_9364,N_9208);
xor U9835 (N_9835,N_9297,N_8912);
nor U9836 (N_9836,N_9139,N_9141);
xnor U9837 (N_9837,N_9473,N_9038);
xor U9838 (N_9838,N_8818,N_9215);
or U9839 (N_9839,N_8838,N_9387);
or U9840 (N_9840,N_9187,N_9224);
or U9841 (N_9841,N_8970,N_9352);
and U9842 (N_9842,N_9497,N_9463);
or U9843 (N_9843,N_9532,N_9574);
or U9844 (N_9844,N_9423,N_8844);
xnor U9845 (N_9845,N_9370,N_8890);
nor U9846 (N_9846,N_8855,N_8839);
nand U9847 (N_9847,N_9563,N_9404);
nor U9848 (N_9848,N_8861,N_9384);
nand U9849 (N_9849,N_9112,N_9062);
or U9850 (N_9850,N_8824,N_8945);
nand U9851 (N_9851,N_9337,N_8833);
and U9852 (N_9852,N_9597,N_9496);
and U9853 (N_9853,N_9478,N_8879);
and U9854 (N_9854,N_9296,N_9388);
xnor U9855 (N_9855,N_9310,N_8962);
xnor U9856 (N_9856,N_9185,N_9413);
or U9857 (N_9857,N_9460,N_9592);
nand U9858 (N_9858,N_9081,N_8876);
or U9859 (N_9859,N_9448,N_8840);
xnor U9860 (N_9860,N_9219,N_9064);
or U9861 (N_9861,N_9177,N_9018);
nor U9862 (N_9862,N_9183,N_9259);
or U9863 (N_9863,N_9551,N_8894);
nand U9864 (N_9864,N_8878,N_9061);
or U9865 (N_9865,N_9210,N_9506);
nand U9866 (N_9866,N_9503,N_9020);
nor U9867 (N_9867,N_9535,N_9484);
nand U9868 (N_9868,N_9579,N_8800);
xnor U9869 (N_9869,N_9227,N_9514);
or U9870 (N_9870,N_8849,N_9528);
nand U9871 (N_9871,N_9426,N_9479);
nor U9872 (N_9872,N_9004,N_8843);
nand U9873 (N_9873,N_9169,N_8887);
nand U9874 (N_9874,N_9577,N_8891);
xor U9875 (N_9875,N_8998,N_9129);
xnor U9876 (N_9876,N_9571,N_9570);
or U9877 (N_9877,N_9451,N_9332);
xor U9878 (N_9878,N_9104,N_9039);
nand U9879 (N_9879,N_9294,N_9212);
or U9880 (N_9880,N_9070,N_9581);
nor U9881 (N_9881,N_9385,N_9490);
nand U9882 (N_9882,N_8905,N_8801);
xor U9883 (N_9883,N_9424,N_9225);
and U9884 (N_9884,N_8988,N_9327);
xor U9885 (N_9885,N_9419,N_8951);
nor U9886 (N_9886,N_9547,N_9015);
and U9887 (N_9887,N_8854,N_9124);
and U9888 (N_9888,N_9089,N_9196);
nor U9889 (N_9889,N_9363,N_9546);
nand U9890 (N_9890,N_9495,N_9174);
xnor U9891 (N_9891,N_8900,N_9513);
and U9892 (N_9892,N_9073,N_8845);
nor U9893 (N_9893,N_9206,N_9078);
xnor U9894 (N_9894,N_8883,N_8882);
nand U9895 (N_9895,N_8979,N_9433);
nand U9896 (N_9896,N_8956,N_9493);
and U9897 (N_9897,N_9564,N_8922);
nand U9898 (N_9898,N_8915,N_8802);
or U9899 (N_9899,N_9299,N_9287);
and U9900 (N_9900,N_8940,N_9575);
and U9901 (N_9901,N_8877,N_8975);
nand U9902 (N_9902,N_9268,N_9056);
nand U9903 (N_9903,N_9328,N_9072);
or U9904 (N_9904,N_8889,N_9242);
xnor U9905 (N_9905,N_9379,N_9322);
xor U9906 (N_9906,N_9007,N_9032);
nor U9907 (N_9907,N_9068,N_8864);
and U9908 (N_9908,N_8906,N_9512);
xor U9909 (N_9909,N_9372,N_8928);
or U9910 (N_9910,N_9080,N_9531);
xnor U9911 (N_9911,N_9464,N_9324);
or U9912 (N_9912,N_9017,N_9197);
or U9913 (N_9913,N_9317,N_9016);
or U9914 (N_9914,N_9264,N_9146);
xnor U9915 (N_9915,N_9431,N_9036);
and U9916 (N_9916,N_9200,N_8816);
nor U9917 (N_9917,N_8826,N_9336);
or U9918 (N_9918,N_9396,N_8980);
nor U9919 (N_9919,N_8803,N_9021);
or U9920 (N_9920,N_9524,N_9298);
and U9921 (N_9921,N_8971,N_9145);
xnor U9922 (N_9922,N_8895,N_9246);
or U9923 (N_9923,N_9338,N_9262);
and U9924 (N_9924,N_9131,N_9454);
nand U9925 (N_9925,N_9277,N_9558);
xor U9926 (N_9926,N_8964,N_9377);
or U9927 (N_9927,N_8804,N_8866);
nor U9928 (N_9928,N_8907,N_9405);
nand U9929 (N_9929,N_8923,N_9102);
xnor U9930 (N_9930,N_9325,N_9375);
nor U9931 (N_9931,N_9315,N_8972);
or U9932 (N_9932,N_8960,N_9320);
nor U9933 (N_9933,N_9354,N_9590);
xor U9934 (N_9934,N_8976,N_9184);
nor U9935 (N_9935,N_8996,N_9301);
and U9936 (N_9936,N_8977,N_8909);
xor U9937 (N_9937,N_9042,N_8963);
nor U9938 (N_9938,N_8961,N_9122);
or U9939 (N_9939,N_9172,N_8898);
nand U9940 (N_9940,N_8921,N_9319);
nor U9941 (N_9941,N_9118,N_9425);
xor U9942 (N_9942,N_9498,N_9222);
nand U9943 (N_9943,N_8893,N_8991);
and U9944 (N_9944,N_9447,N_8947);
nand U9945 (N_9945,N_9540,N_9292);
nor U9946 (N_9946,N_9186,N_8935);
xnor U9947 (N_9947,N_9098,N_9537);
xor U9948 (N_9948,N_9057,N_9501);
nand U9949 (N_9949,N_9054,N_9255);
and U9950 (N_9950,N_8943,N_9272);
or U9951 (N_9951,N_9517,N_9382);
nor U9952 (N_9952,N_9155,N_8934);
nand U9953 (N_9953,N_9389,N_9312);
xnor U9954 (N_9954,N_9166,N_9435);
nand U9955 (N_9955,N_9065,N_9409);
nor U9956 (N_9956,N_8952,N_8995);
and U9957 (N_9957,N_9499,N_9238);
and U9958 (N_9958,N_8983,N_9267);
nand U9959 (N_9959,N_9031,N_9504);
nor U9960 (N_9960,N_9529,N_9204);
or U9961 (N_9961,N_9542,N_9269);
and U9962 (N_9962,N_9101,N_9443);
nor U9963 (N_9963,N_9343,N_9250);
xnor U9964 (N_9964,N_9369,N_9022);
or U9965 (N_9965,N_9012,N_9067);
xnor U9966 (N_9966,N_8959,N_9135);
and U9967 (N_9967,N_9084,N_8904);
and U9968 (N_9968,N_8842,N_8888);
and U9969 (N_9969,N_9323,N_8999);
nor U9970 (N_9970,N_9123,N_9258);
and U9971 (N_9971,N_9044,N_9288);
xnor U9972 (N_9972,N_9534,N_9188);
nor U9973 (N_9973,N_8916,N_9456);
xnor U9974 (N_9974,N_9137,N_8815);
or U9975 (N_9975,N_9420,N_9386);
or U9976 (N_9976,N_9446,N_8936);
nor U9977 (N_9977,N_8811,N_9052);
nor U9978 (N_9978,N_9526,N_9357);
nand U9979 (N_9979,N_8985,N_9450);
and U9980 (N_9980,N_8994,N_9480);
or U9981 (N_9981,N_9009,N_9025);
nand U9982 (N_9982,N_9164,N_9244);
or U9983 (N_9983,N_9314,N_9019);
and U9984 (N_9984,N_9530,N_8978);
and U9985 (N_9985,N_9115,N_9510);
and U9986 (N_9986,N_9544,N_9005);
and U9987 (N_9987,N_9076,N_8809);
xnor U9988 (N_9988,N_9411,N_9144);
xor U9989 (N_9989,N_9157,N_8982);
xor U9990 (N_9990,N_8847,N_9198);
nor U9991 (N_9991,N_8949,N_8831);
or U9992 (N_9992,N_9248,N_9271);
nor U9993 (N_9993,N_9028,N_8820);
nand U9994 (N_9994,N_9554,N_8990);
xor U9995 (N_9995,N_9521,N_8872);
nor U9996 (N_9996,N_9461,N_9151);
nor U9997 (N_9997,N_9027,N_9586);
or U9998 (N_9998,N_9182,N_8918);
nor U9999 (N_9999,N_9421,N_9260);
xnor U10000 (N_10000,N_9598,N_8866);
or U10001 (N_10001,N_9416,N_9213);
nand U10002 (N_10002,N_9530,N_9582);
and U10003 (N_10003,N_9506,N_9181);
nand U10004 (N_10004,N_8850,N_9044);
xor U10005 (N_10005,N_9225,N_9475);
and U10006 (N_10006,N_9205,N_8816);
xnor U10007 (N_10007,N_9232,N_9344);
xor U10008 (N_10008,N_9287,N_9382);
or U10009 (N_10009,N_9211,N_9306);
or U10010 (N_10010,N_9183,N_8858);
nor U10011 (N_10011,N_9559,N_9351);
or U10012 (N_10012,N_9491,N_9143);
or U10013 (N_10013,N_9390,N_9425);
or U10014 (N_10014,N_8898,N_9024);
xor U10015 (N_10015,N_9256,N_9150);
and U10016 (N_10016,N_8963,N_8922);
or U10017 (N_10017,N_8927,N_9054);
xor U10018 (N_10018,N_8905,N_9205);
xor U10019 (N_10019,N_8872,N_8814);
nor U10020 (N_10020,N_9173,N_9305);
or U10021 (N_10021,N_9124,N_9310);
or U10022 (N_10022,N_9430,N_9243);
nand U10023 (N_10023,N_9535,N_9508);
and U10024 (N_10024,N_9412,N_9064);
nor U10025 (N_10025,N_9366,N_9560);
and U10026 (N_10026,N_9428,N_8955);
xnor U10027 (N_10027,N_9569,N_8982);
nor U10028 (N_10028,N_8910,N_9451);
or U10029 (N_10029,N_8898,N_8929);
and U10030 (N_10030,N_9356,N_8800);
xnor U10031 (N_10031,N_9234,N_9174);
nand U10032 (N_10032,N_8831,N_9176);
and U10033 (N_10033,N_9052,N_9224);
and U10034 (N_10034,N_9398,N_9104);
or U10035 (N_10035,N_9155,N_9033);
or U10036 (N_10036,N_9258,N_9096);
and U10037 (N_10037,N_9164,N_9365);
and U10038 (N_10038,N_9207,N_8909);
xor U10039 (N_10039,N_9156,N_9172);
nand U10040 (N_10040,N_9041,N_9504);
xnor U10041 (N_10041,N_8908,N_9362);
nor U10042 (N_10042,N_8981,N_8983);
and U10043 (N_10043,N_9365,N_8824);
nand U10044 (N_10044,N_9527,N_9208);
xnor U10045 (N_10045,N_9349,N_9322);
xnor U10046 (N_10046,N_8878,N_9353);
nor U10047 (N_10047,N_9266,N_9300);
or U10048 (N_10048,N_9162,N_9085);
or U10049 (N_10049,N_8927,N_8894);
nor U10050 (N_10050,N_9346,N_9483);
nor U10051 (N_10051,N_9378,N_9147);
and U10052 (N_10052,N_9561,N_9492);
and U10053 (N_10053,N_8980,N_9339);
nor U10054 (N_10054,N_9390,N_9552);
xnor U10055 (N_10055,N_9267,N_9539);
nand U10056 (N_10056,N_9230,N_9558);
xnor U10057 (N_10057,N_9414,N_9121);
nor U10058 (N_10058,N_9468,N_9509);
or U10059 (N_10059,N_8912,N_8843);
and U10060 (N_10060,N_9319,N_9371);
nand U10061 (N_10061,N_8879,N_9059);
nor U10062 (N_10062,N_9044,N_8814);
or U10063 (N_10063,N_8887,N_9066);
nor U10064 (N_10064,N_9075,N_8931);
xor U10065 (N_10065,N_8842,N_8962);
xnor U10066 (N_10066,N_9069,N_8887);
xnor U10067 (N_10067,N_9385,N_9117);
and U10068 (N_10068,N_8913,N_8967);
nor U10069 (N_10069,N_8869,N_8847);
nand U10070 (N_10070,N_9136,N_9253);
nor U10071 (N_10071,N_9547,N_9360);
nand U10072 (N_10072,N_9362,N_9525);
nand U10073 (N_10073,N_9505,N_9016);
nand U10074 (N_10074,N_9536,N_9328);
nor U10075 (N_10075,N_9381,N_9460);
nor U10076 (N_10076,N_9300,N_8816);
nor U10077 (N_10077,N_9204,N_9314);
nor U10078 (N_10078,N_9489,N_8978);
or U10079 (N_10079,N_9006,N_9212);
xnor U10080 (N_10080,N_9392,N_9490);
nor U10081 (N_10081,N_9573,N_9095);
and U10082 (N_10082,N_9267,N_8906);
xnor U10083 (N_10083,N_9346,N_9467);
and U10084 (N_10084,N_9320,N_9411);
or U10085 (N_10085,N_9250,N_9421);
nand U10086 (N_10086,N_9072,N_9392);
or U10087 (N_10087,N_9211,N_9439);
nand U10088 (N_10088,N_9211,N_8922);
and U10089 (N_10089,N_8975,N_9531);
or U10090 (N_10090,N_9059,N_8825);
nand U10091 (N_10091,N_9400,N_8854);
and U10092 (N_10092,N_9372,N_8932);
nand U10093 (N_10093,N_9118,N_8856);
or U10094 (N_10094,N_9186,N_8822);
nand U10095 (N_10095,N_9323,N_9365);
nand U10096 (N_10096,N_9068,N_8843);
xor U10097 (N_10097,N_8805,N_9351);
and U10098 (N_10098,N_8888,N_9497);
or U10099 (N_10099,N_9088,N_9121);
or U10100 (N_10100,N_8821,N_9304);
xor U10101 (N_10101,N_9187,N_9333);
xor U10102 (N_10102,N_9547,N_9305);
or U10103 (N_10103,N_8863,N_8935);
nor U10104 (N_10104,N_9053,N_9121);
nand U10105 (N_10105,N_9199,N_9025);
nand U10106 (N_10106,N_9144,N_9378);
nor U10107 (N_10107,N_9140,N_9030);
nor U10108 (N_10108,N_9160,N_8872);
or U10109 (N_10109,N_8809,N_9553);
xor U10110 (N_10110,N_9163,N_9574);
nor U10111 (N_10111,N_9032,N_9468);
nand U10112 (N_10112,N_9213,N_8897);
nand U10113 (N_10113,N_8888,N_9502);
xnor U10114 (N_10114,N_9144,N_9475);
nand U10115 (N_10115,N_9328,N_9500);
nand U10116 (N_10116,N_8882,N_8845);
nor U10117 (N_10117,N_9439,N_9359);
and U10118 (N_10118,N_8995,N_9068);
and U10119 (N_10119,N_8956,N_9477);
nor U10120 (N_10120,N_9474,N_9204);
xor U10121 (N_10121,N_8872,N_9325);
or U10122 (N_10122,N_9289,N_9155);
or U10123 (N_10123,N_9154,N_9050);
nor U10124 (N_10124,N_8965,N_9493);
xor U10125 (N_10125,N_9267,N_9320);
xnor U10126 (N_10126,N_9492,N_9426);
xor U10127 (N_10127,N_9002,N_9033);
nor U10128 (N_10128,N_9255,N_9356);
and U10129 (N_10129,N_9166,N_9022);
xnor U10130 (N_10130,N_9595,N_9072);
nor U10131 (N_10131,N_9480,N_9515);
nor U10132 (N_10132,N_9563,N_9506);
xor U10133 (N_10133,N_9139,N_9137);
nor U10134 (N_10134,N_9592,N_9598);
nor U10135 (N_10135,N_9550,N_9422);
xor U10136 (N_10136,N_9130,N_9015);
and U10137 (N_10137,N_9052,N_8806);
and U10138 (N_10138,N_9413,N_8914);
and U10139 (N_10139,N_8934,N_8804);
nand U10140 (N_10140,N_9582,N_9508);
xor U10141 (N_10141,N_8878,N_9122);
nor U10142 (N_10142,N_8827,N_9083);
or U10143 (N_10143,N_9399,N_8969);
or U10144 (N_10144,N_9275,N_9015);
xnor U10145 (N_10145,N_9011,N_9385);
xnor U10146 (N_10146,N_8882,N_9383);
nor U10147 (N_10147,N_9559,N_9047);
nand U10148 (N_10148,N_9072,N_9377);
nor U10149 (N_10149,N_9188,N_9143);
nor U10150 (N_10150,N_9135,N_9302);
or U10151 (N_10151,N_9564,N_8808);
and U10152 (N_10152,N_9520,N_8982);
nor U10153 (N_10153,N_8816,N_9438);
nor U10154 (N_10154,N_9505,N_8881);
xor U10155 (N_10155,N_9415,N_8953);
nor U10156 (N_10156,N_8934,N_9009);
xnor U10157 (N_10157,N_9529,N_9542);
xnor U10158 (N_10158,N_9573,N_9314);
xor U10159 (N_10159,N_9013,N_9203);
xnor U10160 (N_10160,N_9266,N_9167);
or U10161 (N_10161,N_9107,N_9020);
xnor U10162 (N_10162,N_9361,N_9284);
and U10163 (N_10163,N_8898,N_9281);
xnor U10164 (N_10164,N_9105,N_8909);
or U10165 (N_10165,N_9096,N_8860);
nand U10166 (N_10166,N_8888,N_9072);
nor U10167 (N_10167,N_9248,N_9586);
or U10168 (N_10168,N_8943,N_8931);
or U10169 (N_10169,N_9089,N_8962);
nor U10170 (N_10170,N_9060,N_8884);
nor U10171 (N_10171,N_9348,N_8860);
and U10172 (N_10172,N_8802,N_9259);
or U10173 (N_10173,N_9254,N_8954);
and U10174 (N_10174,N_8950,N_8937);
xor U10175 (N_10175,N_8869,N_8866);
or U10176 (N_10176,N_9157,N_8814);
and U10177 (N_10177,N_9266,N_8951);
nand U10178 (N_10178,N_9077,N_8910);
and U10179 (N_10179,N_9046,N_9103);
nor U10180 (N_10180,N_9375,N_9250);
xor U10181 (N_10181,N_9056,N_9286);
or U10182 (N_10182,N_9247,N_9422);
or U10183 (N_10183,N_9579,N_8815);
nand U10184 (N_10184,N_8804,N_8833);
nand U10185 (N_10185,N_9474,N_9254);
nor U10186 (N_10186,N_9287,N_8803);
nor U10187 (N_10187,N_9433,N_8938);
xnor U10188 (N_10188,N_9574,N_9553);
or U10189 (N_10189,N_9355,N_9394);
nor U10190 (N_10190,N_9178,N_9598);
nand U10191 (N_10191,N_9564,N_8828);
or U10192 (N_10192,N_8924,N_9326);
nor U10193 (N_10193,N_9214,N_9330);
xnor U10194 (N_10194,N_9481,N_8841);
xor U10195 (N_10195,N_8979,N_9029);
nand U10196 (N_10196,N_9549,N_9512);
and U10197 (N_10197,N_8848,N_9352);
xnor U10198 (N_10198,N_8906,N_9309);
and U10199 (N_10199,N_9359,N_8846);
nor U10200 (N_10200,N_8872,N_9398);
nor U10201 (N_10201,N_9411,N_9145);
or U10202 (N_10202,N_9325,N_8858);
and U10203 (N_10203,N_9379,N_9275);
nor U10204 (N_10204,N_9302,N_9038);
nor U10205 (N_10205,N_9187,N_8829);
or U10206 (N_10206,N_9532,N_9459);
xnor U10207 (N_10207,N_9499,N_9221);
nor U10208 (N_10208,N_9227,N_9475);
nor U10209 (N_10209,N_8835,N_8809);
nand U10210 (N_10210,N_9431,N_8891);
or U10211 (N_10211,N_8860,N_8961);
nor U10212 (N_10212,N_9361,N_8944);
nand U10213 (N_10213,N_8937,N_9586);
or U10214 (N_10214,N_9093,N_9346);
or U10215 (N_10215,N_9052,N_9440);
or U10216 (N_10216,N_9049,N_8899);
and U10217 (N_10217,N_9285,N_9404);
nand U10218 (N_10218,N_9369,N_9452);
xor U10219 (N_10219,N_9111,N_8826);
and U10220 (N_10220,N_9043,N_9150);
nor U10221 (N_10221,N_9235,N_9494);
and U10222 (N_10222,N_9577,N_9402);
nand U10223 (N_10223,N_9283,N_9238);
or U10224 (N_10224,N_9156,N_9487);
xor U10225 (N_10225,N_9480,N_8885);
nor U10226 (N_10226,N_9095,N_9514);
nor U10227 (N_10227,N_9193,N_9256);
and U10228 (N_10228,N_9461,N_8953);
or U10229 (N_10229,N_9210,N_9522);
xnor U10230 (N_10230,N_9009,N_9522);
nor U10231 (N_10231,N_8861,N_9323);
xnor U10232 (N_10232,N_9356,N_9451);
xor U10233 (N_10233,N_9557,N_9199);
nor U10234 (N_10234,N_9211,N_9576);
nor U10235 (N_10235,N_8851,N_9471);
xor U10236 (N_10236,N_9229,N_9237);
or U10237 (N_10237,N_9580,N_8867);
nor U10238 (N_10238,N_9380,N_9530);
nand U10239 (N_10239,N_9406,N_9528);
and U10240 (N_10240,N_9471,N_8920);
and U10241 (N_10241,N_9571,N_9448);
or U10242 (N_10242,N_8941,N_9217);
nor U10243 (N_10243,N_8920,N_9536);
or U10244 (N_10244,N_8892,N_9031);
nor U10245 (N_10245,N_9410,N_9348);
nor U10246 (N_10246,N_8981,N_8819);
nand U10247 (N_10247,N_9518,N_9234);
nand U10248 (N_10248,N_9199,N_8956);
or U10249 (N_10249,N_8908,N_8831);
or U10250 (N_10250,N_8963,N_9541);
and U10251 (N_10251,N_9046,N_9522);
xor U10252 (N_10252,N_8805,N_9421);
and U10253 (N_10253,N_9392,N_9426);
nand U10254 (N_10254,N_9518,N_8843);
nand U10255 (N_10255,N_9146,N_9220);
or U10256 (N_10256,N_9109,N_9042);
nor U10257 (N_10257,N_9557,N_9447);
xnor U10258 (N_10258,N_9482,N_9103);
xnor U10259 (N_10259,N_9079,N_9372);
nor U10260 (N_10260,N_9181,N_9427);
nand U10261 (N_10261,N_9413,N_9157);
nand U10262 (N_10262,N_9037,N_9021);
and U10263 (N_10263,N_9075,N_9051);
nor U10264 (N_10264,N_9002,N_9111);
nand U10265 (N_10265,N_9531,N_9098);
nand U10266 (N_10266,N_9228,N_9520);
xor U10267 (N_10267,N_8894,N_8855);
nor U10268 (N_10268,N_9495,N_9286);
or U10269 (N_10269,N_9460,N_9500);
xnor U10270 (N_10270,N_8978,N_9122);
nor U10271 (N_10271,N_9348,N_9008);
or U10272 (N_10272,N_9562,N_8856);
and U10273 (N_10273,N_9446,N_8934);
and U10274 (N_10274,N_8852,N_9026);
nor U10275 (N_10275,N_9248,N_9117);
xnor U10276 (N_10276,N_9345,N_9353);
and U10277 (N_10277,N_8994,N_8924);
or U10278 (N_10278,N_8991,N_8927);
nand U10279 (N_10279,N_8819,N_8801);
nor U10280 (N_10280,N_9043,N_8845);
nor U10281 (N_10281,N_9147,N_8947);
or U10282 (N_10282,N_9394,N_8875);
or U10283 (N_10283,N_9415,N_9072);
or U10284 (N_10284,N_8975,N_8839);
nor U10285 (N_10285,N_9192,N_9142);
and U10286 (N_10286,N_9529,N_8839);
nand U10287 (N_10287,N_9315,N_8852);
nor U10288 (N_10288,N_8964,N_8880);
nand U10289 (N_10289,N_8837,N_9364);
nor U10290 (N_10290,N_9309,N_9205);
or U10291 (N_10291,N_9528,N_9074);
xor U10292 (N_10292,N_9247,N_9373);
nor U10293 (N_10293,N_8943,N_9427);
and U10294 (N_10294,N_9263,N_8906);
xnor U10295 (N_10295,N_9559,N_8999);
or U10296 (N_10296,N_9376,N_9306);
or U10297 (N_10297,N_9498,N_9145);
nand U10298 (N_10298,N_9374,N_9422);
nand U10299 (N_10299,N_9342,N_8884);
nand U10300 (N_10300,N_9377,N_9199);
and U10301 (N_10301,N_9243,N_8830);
or U10302 (N_10302,N_9132,N_9569);
nor U10303 (N_10303,N_9013,N_9433);
nand U10304 (N_10304,N_9283,N_8831);
or U10305 (N_10305,N_9520,N_9411);
or U10306 (N_10306,N_9576,N_9438);
nand U10307 (N_10307,N_9372,N_9240);
nor U10308 (N_10308,N_9174,N_9260);
nand U10309 (N_10309,N_9470,N_9335);
nor U10310 (N_10310,N_9504,N_9045);
nand U10311 (N_10311,N_9594,N_9420);
or U10312 (N_10312,N_9164,N_9304);
nor U10313 (N_10313,N_9097,N_8804);
nor U10314 (N_10314,N_9099,N_9314);
or U10315 (N_10315,N_9357,N_8954);
nand U10316 (N_10316,N_9404,N_9382);
or U10317 (N_10317,N_9229,N_9161);
or U10318 (N_10318,N_8963,N_9292);
nand U10319 (N_10319,N_9056,N_8937);
or U10320 (N_10320,N_9118,N_9519);
xnor U10321 (N_10321,N_9585,N_9377);
nor U10322 (N_10322,N_9043,N_9014);
nor U10323 (N_10323,N_8815,N_8926);
nand U10324 (N_10324,N_9008,N_9220);
or U10325 (N_10325,N_8840,N_8828);
xnor U10326 (N_10326,N_9304,N_9390);
nand U10327 (N_10327,N_9215,N_9154);
nor U10328 (N_10328,N_9418,N_9334);
or U10329 (N_10329,N_9237,N_9466);
xor U10330 (N_10330,N_9549,N_9029);
and U10331 (N_10331,N_8894,N_9399);
nand U10332 (N_10332,N_9202,N_9475);
and U10333 (N_10333,N_9454,N_9237);
nor U10334 (N_10334,N_9561,N_8996);
nor U10335 (N_10335,N_9124,N_9077);
and U10336 (N_10336,N_9593,N_9271);
and U10337 (N_10337,N_9445,N_9442);
nand U10338 (N_10338,N_9067,N_9125);
xor U10339 (N_10339,N_9283,N_9575);
nand U10340 (N_10340,N_9402,N_9560);
xor U10341 (N_10341,N_9592,N_9184);
and U10342 (N_10342,N_8969,N_9207);
nor U10343 (N_10343,N_8968,N_8865);
nor U10344 (N_10344,N_9218,N_9150);
xnor U10345 (N_10345,N_8861,N_9351);
nand U10346 (N_10346,N_9164,N_9289);
xnor U10347 (N_10347,N_8867,N_8884);
nand U10348 (N_10348,N_9177,N_9283);
and U10349 (N_10349,N_8875,N_9078);
xor U10350 (N_10350,N_8886,N_8933);
or U10351 (N_10351,N_8940,N_8956);
xnor U10352 (N_10352,N_8967,N_9538);
nand U10353 (N_10353,N_9037,N_9496);
nand U10354 (N_10354,N_9419,N_8928);
nor U10355 (N_10355,N_9320,N_9393);
xor U10356 (N_10356,N_8915,N_9163);
or U10357 (N_10357,N_8925,N_9043);
xnor U10358 (N_10358,N_9162,N_9068);
and U10359 (N_10359,N_9311,N_9443);
nor U10360 (N_10360,N_9204,N_9098);
or U10361 (N_10361,N_9470,N_9270);
or U10362 (N_10362,N_9009,N_9438);
xor U10363 (N_10363,N_9393,N_8825);
or U10364 (N_10364,N_8910,N_9069);
nand U10365 (N_10365,N_9130,N_9562);
and U10366 (N_10366,N_9235,N_9112);
nand U10367 (N_10367,N_9474,N_9498);
nand U10368 (N_10368,N_9529,N_9203);
nand U10369 (N_10369,N_9506,N_9153);
nand U10370 (N_10370,N_9559,N_9118);
nand U10371 (N_10371,N_9331,N_9563);
and U10372 (N_10372,N_9424,N_8809);
and U10373 (N_10373,N_8860,N_9465);
nand U10374 (N_10374,N_8907,N_8954);
nor U10375 (N_10375,N_8995,N_9313);
xor U10376 (N_10376,N_9374,N_9222);
or U10377 (N_10377,N_9412,N_8898);
xnor U10378 (N_10378,N_9571,N_9273);
nand U10379 (N_10379,N_9014,N_9382);
or U10380 (N_10380,N_9194,N_9431);
or U10381 (N_10381,N_8986,N_9039);
or U10382 (N_10382,N_9407,N_9336);
xnor U10383 (N_10383,N_9067,N_9545);
or U10384 (N_10384,N_9532,N_9188);
nor U10385 (N_10385,N_9217,N_9000);
or U10386 (N_10386,N_9397,N_9588);
or U10387 (N_10387,N_9182,N_9044);
or U10388 (N_10388,N_8993,N_8858);
or U10389 (N_10389,N_8866,N_8978);
nor U10390 (N_10390,N_9045,N_9116);
nor U10391 (N_10391,N_9321,N_9483);
xor U10392 (N_10392,N_9447,N_8952);
or U10393 (N_10393,N_9388,N_9278);
or U10394 (N_10394,N_9554,N_9355);
xnor U10395 (N_10395,N_8855,N_9312);
xnor U10396 (N_10396,N_9122,N_9345);
xor U10397 (N_10397,N_8941,N_9254);
nand U10398 (N_10398,N_9171,N_8801);
nand U10399 (N_10399,N_9298,N_8858);
xor U10400 (N_10400,N_9883,N_10312);
nand U10401 (N_10401,N_9787,N_10198);
xnor U10402 (N_10402,N_9656,N_10001);
nand U10403 (N_10403,N_9614,N_9747);
or U10404 (N_10404,N_9710,N_9625);
or U10405 (N_10405,N_10153,N_9693);
or U10406 (N_10406,N_9696,N_9873);
or U10407 (N_10407,N_9954,N_10028);
or U10408 (N_10408,N_9781,N_9805);
nor U10409 (N_10409,N_10229,N_10351);
and U10410 (N_10410,N_9819,N_10343);
and U10411 (N_10411,N_10238,N_9928);
and U10412 (N_10412,N_10019,N_10133);
and U10413 (N_10413,N_9990,N_10048);
and U10414 (N_10414,N_9639,N_9922);
nand U10415 (N_10415,N_10239,N_10345);
or U10416 (N_10416,N_10381,N_10163);
and U10417 (N_10417,N_9973,N_9833);
and U10418 (N_10418,N_10127,N_10247);
xnor U10419 (N_10419,N_10214,N_10282);
nor U10420 (N_10420,N_9706,N_10279);
or U10421 (N_10421,N_10287,N_10297);
or U10422 (N_10422,N_10313,N_10038);
nand U10423 (N_10423,N_10068,N_10066);
xor U10424 (N_10424,N_9882,N_10232);
and U10425 (N_10425,N_9750,N_10215);
or U10426 (N_10426,N_9764,N_10237);
nor U10427 (N_10427,N_9689,N_9790);
and U10428 (N_10428,N_10029,N_9619);
and U10429 (N_10429,N_9923,N_10358);
xnor U10430 (N_10430,N_10188,N_10074);
nand U10431 (N_10431,N_9729,N_9856);
or U10432 (N_10432,N_9815,N_10393);
xor U10433 (N_10433,N_10035,N_9649);
xnor U10434 (N_10434,N_9801,N_10046);
or U10435 (N_10435,N_10105,N_9676);
nor U10436 (N_10436,N_9866,N_10058);
xor U10437 (N_10437,N_9769,N_10132);
and U10438 (N_10438,N_10075,N_10385);
or U10439 (N_10439,N_9921,N_10146);
nor U10440 (N_10440,N_10037,N_10080);
nor U10441 (N_10441,N_10257,N_10373);
nor U10442 (N_10442,N_9776,N_10069);
xor U10443 (N_10443,N_10272,N_10114);
nor U10444 (N_10444,N_9924,N_10150);
and U10445 (N_10445,N_9711,N_9838);
nand U10446 (N_10446,N_9820,N_10225);
nand U10447 (N_10447,N_10295,N_10368);
or U10448 (N_10448,N_10228,N_10321);
xnor U10449 (N_10449,N_9733,N_10226);
nor U10450 (N_10450,N_9888,N_9969);
nand U10451 (N_10451,N_10333,N_9862);
and U10452 (N_10452,N_10298,N_10040);
and U10453 (N_10453,N_10332,N_9697);
nand U10454 (N_10454,N_10087,N_9908);
xor U10455 (N_10455,N_9932,N_10118);
and U10456 (N_10456,N_10361,N_9653);
or U10457 (N_10457,N_10253,N_10383);
or U10458 (N_10458,N_9878,N_10022);
nor U10459 (N_10459,N_10128,N_10149);
xor U10460 (N_10460,N_9905,N_9739);
nor U10461 (N_10461,N_10026,N_10376);
nor U10462 (N_10462,N_10258,N_9887);
nor U10463 (N_10463,N_9961,N_10121);
xor U10464 (N_10464,N_10330,N_10387);
and U10465 (N_10465,N_10086,N_10005);
nor U10466 (N_10466,N_9813,N_10168);
nand U10467 (N_10467,N_10267,N_10325);
or U10468 (N_10468,N_10220,N_9677);
nand U10469 (N_10469,N_10241,N_10085);
and U10470 (N_10470,N_9647,N_9846);
nand U10471 (N_10471,N_9864,N_10224);
xor U10472 (N_10472,N_10236,N_9616);
xnor U10473 (N_10473,N_9687,N_10172);
nor U10474 (N_10474,N_9914,N_10205);
nand U10475 (N_10475,N_10284,N_10120);
nor U10476 (N_10476,N_10350,N_10342);
and U10477 (N_10477,N_10095,N_9621);
nor U10478 (N_10478,N_9944,N_9986);
nor U10479 (N_10479,N_9977,N_9763);
or U10480 (N_10480,N_10144,N_10165);
or U10481 (N_10481,N_9708,N_9952);
nand U10482 (N_10482,N_10310,N_10043);
or U10483 (N_10483,N_9731,N_9782);
nand U10484 (N_10484,N_9774,N_10203);
or U10485 (N_10485,N_10071,N_10062);
and U10486 (N_10486,N_10396,N_10307);
nand U10487 (N_10487,N_9675,N_9811);
or U10488 (N_10488,N_10015,N_9876);
nand U10489 (N_10489,N_9860,N_9655);
and U10490 (N_10490,N_10006,N_10033);
xor U10491 (N_10491,N_10036,N_10178);
and U10492 (N_10492,N_9768,N_10108);
and U10493 (N_10493,N_10211,N_9610);
nor U10494 (N_10494,N_9725,N_10347);
nor U10495 (N_10495,N_9648,N_10157);
or U10496 (N_10496,N_9985,N_9628);
xnor U10497 (N_10497,N_10125,N_9946);
and U10498 (N_10498,N_10223,N_10335);
xor U10499 (N_10499,N_10030,N_9857);
nand U10500 (N_10500,N_10138,N_10334);
and U10501 (N_10501,N_10327,N_9831);
nand U10502 (N_10502,N_10185,N_9943);
nand U10503 (N_10503,N_10079,N_9945);
xnor U10504 (N_10504,N_10249,N_9915);
xor U10505 (N_10505,N_9827,N_10156);
nand U10506 (N_10506,N_9780,N_10174);
nand U10507 (N_10507,N_10131,N_10115);
xnor U10508 (N_10508,N_9691,N_9816);
or U10509 (N_10509,N_9828,N_9717);
nor U10510 (N_10510,N_9902,N_10049);
or U10511 (N_10511,N_10076,N_9615);
nand U10512 (N_10512,N_10367,N_10265);
xnor U10513 (N_10513,N_9971,N_10260);
xor U10514 (N_10514,N_9715,N_10377);
nand U10515 (N_10515,N_10291,N_9669);
nand U10516 (N_10516,N_10092,N_10057);
and U10517 (N_10517,N_9812,N_9798);
or U10518 (N_10518,N_9761,N_10060);
and U10519 (N_10519,N_9877,N_10160);
nand U10520 (N_10520,N_9868,N_10397);
nand U10521 (N_10521,N_10166,N_9658);
nor U10522 (N_10522,N_9855,N_10235);
nor U10523 (N_10523,N_10240,N_9775);
xor U10524 (N_10524,N_9757,N_10338);
nor U10525 (N_10525,N_10013,N_10285);
and U10526 (N_10526,N_9636,N_9916);
or U10527 (N_10527,N_10191,N_10374);
and U10528 (N_10528,N_9839,N_9665);
nor U10529 (N_10529,N_9728,N_9972);
and U10530 (N_10530,N_10317,N_10130);
nor U10531 (N_10531,N_10276,N_10204);
nand U10532 (N_10532,N_9832,N_9875);
or U10533 (N_10533,N_9901,N_10097);
nand U10534 (N_10534,N_10341,N_9705);
or U10535 (N_10535,N_9630,N_10143);
xnor U10536 (N_10536,N_10230,N_10182);
and U10537 (N_10537,N_10094,N_10304);
nor U10538 (N_10538,N_9858,N_10113);
xor U10539 (N_10539,N_10009,N_9632);
nor U10540 (N_10540,N_10164,N_10045);
and U10541 (N_10541,N_10104,N_10077);
xor U10542 (N_10542,N_9698,N_9641);
and U10543 (N_10543,N_9983,N_10308);
nor U10544 (N_10544,N_9984,N_9891);
nand U10545 (N_10545,N_10122,N_9744);
xnor U10546 (N_10546,N_10109,N_9841);
or U10547 (N_10547,N_9848,N_10096);
nand U10548 (N_10548,N_9918,N_9679);
xnor U10549 (N_10549,N_9817,N_10251);
nor U10550 (N_10550,N_9652,N_9889);
and U10551 (N_10551,N_10281,N_10100);
nand U10552 (N_10552,N_10202,N_10388);
or U10553 (N_10553,N_9970,N_10159);
nor U10554 (N_10554,N_9942,N_9657);
and U10555 (N_10555,N_10289,N_9904);
nand U10556 (N_10556,N_10306,N_9783);
nand U10557 (N_10557,N_10123,N_10021);
or U10558 (N_10558,N_9886,N_10088);
or U10559 (N_10559,N_9951,N_9633);
nand U10560 (N_10560,N_9784,N_10370);
xnor U10561 (N_10561,N_9881,N_9822);
nand U10562 (N_10562,N_9722,N_9859);
nand U10563 (N_10563,N_10231,N_9853);
nand U10564 (N_10564,N_10041,N_10371);
nor U10565 (N_10565,N_9746,N_9899);
or U10566 (N_10566,N_9796,N_10273);
nor U10567 (N_10567,N_9745,N_9861);
nand U10568 (N_10568,N_10020,N_10320);
nand U10569 (N_10569,N_10359,N_10380);
xor U10570 (N_10570,N_9823,N_10129);
xor U10571 (N_10571,N_10158,N_10101);
and U10572 (N_10572,N_9770,N_9893);
nand U10573 (N_10573,N_9695,N_9974);
nand U10574 (N_10574,N_10314,N_9950);
and U10575 (N_10575,N_9803,N_9723);
nor U10576 (N_10576,N_9701,N_9953);
nor U10577 (N_10577,N_9663,N_9992);
xnor U10578 (N_10578,N_9793,N_10252);
or U10579 (N_10579,N_10365,N_10389);
and U10580 (N_10580,N_9907,N_10233);
xor U10581 (N_10581,N_10318,N_10025);
nand U10582 (N_10582,N_9699,N_10213);
nor U10583 (N_10583,N_10246,N_9753);
xnor U10584 (N_10584,N_9879,N_9773);
nor U10585 (N_10585,N_10274,N_10216);
or U10586 (N_10586,N_10296,N_9683);
or U10587 (N_10587,N_9991,N_10288);
xor U10588 (N_10588,N_9939,N_9791);
nand U10589 (N_10589,N_10061,N_9936);
nor U10590 (N_10590,N_9849,N_10208);
and U10591 (N_10591,N_10145,N_10179);
xnor U10592 (N_10592,N_10135,N_10116);
nand U10593 (N_10593,N_9792,N_9933);
xor U10594 (N_10594,N_10323,N_10003);
nand U10595 (N_10595,N_9690,N_10269);
nor U10596 (N_10596,N_10169,N_9981);
xnor U10597 (N_10597,N_10275,N_9667);
nand U10598 (N_10598,N_9987,N_9692);
or U10599 (N_10599,N_9627,N_10250);
and U10600 (N_10600,N_10315,N_10336);
and U10601 (N_10601,N_10192,N_9777);
xnor U10602 (N_10602,N_9824,N_9988);
xor U10603 (N_10603,N_10089,N_10360);
xor U10604 (N_10604,N_9994,N_9642);
and U10605 (N_10605,N_9623,N_9741);
and U10606 (N_10606,N_9799,N_9821);
nor U10607 (N_10607,N_9925,N_9968);
xor U10608 (N_10608,N_10091,N_9959);
or U10609 (N_10609,N_9929,N_9847);
and U10610 (N_10610,N_10243,N_9718);
and U10611 (N_10611,N_10364,N_9870);
nand U10612 (N_10612,N_10050,N_10271);
and U10613 (N_10613,N_10299,N_9617);
nor U10614 (N_10614,N_10090,N_10084);
or U10615 (N_10615,N_9938,N_9626);
nor U10616 (N_10616,N_9712,N_9962);
nor U10617 (N_10617,N_9960,N_9949);
xor U10618 (N_10618,N_9818,N_10254);
nand U10619 (N_10619,N_10126,N_9756);
nand U10620 (N_10620,N_10177,N_10098);
or U10621 (N_10621,N_10277,N_9967);
nor U10622 (N_10622,N_10139,N_10052);
xnor U10623 (N_10623,N_9802,N_9748);
and U10624 (N_10624,N_9937,N_9732);
and U10625 (N_10625,N_9797,N_9975);
or U10626 (N_10626,N_10300,N_10234);
or U10627 (N_10627,N_9976,N_9894);
nor U10628 (N_10628,N_9844,N_9620);
nand U10629 (N_10629,N_9727,N_10355);
xnor U10630 (N_10630,N_10196,N_10319);
and U10631 (N_10631,N_10248,N_10171);
xor U10632 (N_10632,N_10176,N_9854);
and U10633 (N_10633,N_10245,N_10102);
nand U10634 (N_10634,N_9618,N_10184);
or U10635 (N_10635,N_10209,N_10034);
nand U10636 (N_10636,N_10346,N_9721);
xor U10637 (N_10637,N_10366,N_9863);
xnor U10638 (N_10638,N_10137,N_10268);
nor U10639 (N_10639,N_10000,N_10344);
nand U10640 (N_10640,N_10072,N_9659);
and U10641 (N_10641,N_10378,N_10190);
and U10642 (N_10642,N_9851,N_10170);
nand U10643 (N_10643,N_10212,N_10199);
xnor U10644 (N_10644,N_9704,N_9997);
or U10645 (N_10645,N_10175,N_10339);
xor U10646 (N_10646,N_9806,N_9867);
xor U10647 (N_10647,N_9910,N_10051);
or U10648 (N_10648,N_9606,N_10195);
or U10649 (N_10649,N_10055,N_10111);
xor U10650 (N_10650,N_10067,N_9835);
and U10651 (N_10651,N_10112,N_9605);
and U10652 (N_10652,N_10141,N_9825);
xnor U10653 (N_10653,N_10270,N_10316);
or U10654 (N_10654,N_9809,N_9635);
nand U10655 (N_10655,N_10024,N_9752);
xnor U10656 (N_10656,N_10099,N_9685);
and U10657 (N_10657,N_9840,N_10002);
nand U10658 (N_10658,N_10027,N_9919);
xor U10659 (N_10659,N_10218,N_9650);
and U10660 (N_10660,N_10242,N_9754);
and U10661 (N_10661,N_9643,N_10183);
or U10662 (N_10662,N_10244,N_9670);
and U10663 (N_10663,N_9965,N_10264);
xnor U10664 (N_10664,N_10197,N_9800);
and U10665 (N_10665,N_10375,N_9682);
xor U10666 (N_10666,N_9958,N_10011);
nor U10667 (N_10667,N_10107,N_9941);
or U10668 (N_10668,N_10379,N_9808);
xor U10669 (N_10669,N_9743,N_10073);
nand U10670 (N_10670,N_9765,N_9948);
nor U10671 (N_10671,N_9850,N_10386);
nor U10672 (N_10672,N_9688,N_9785);
or U10673 (N_10673,N_10017,N_9637);
and U10674 (N_10674,N_9651,N_9998);
xor U10675 (N_10675,N_9661,N_10348);
or U10676 (N_10676,N_9814,N_10014);
and U10677 (N_10677,N_10152,N_9779);
and U10678 (N_10678,N_9999,N_9980);
xnor U10679 (N_10679,N_10065,N_9601);
nor U10680 (N_10680,N_10210,N_10010);
xor U10681 (N_10681,N_10259,N_9672);
xor U10682 (N_10682,N_10290,N_10309);
xor U10683 (N_10683,N_10142,N_10004);
nor U10684 (N_10684,N_9640,N_9957);
or U10685 (N_10685,N_9720,N_9654);
or U10686 (N_10686,N_9871,N_9843);
xor U10687 (N_10687,N_10256,N_9603);
xnor U10688 (N_10688,N_9934,N_9830);
nor U10689 (N_10689,N_10056,N_9837);
nand U10690 (N_10690,N_10227,N_10187);
or U10691 (N_10691,N_10357,N_10193);
nand U10692 (N_10692,N_9995,N_9629);
nor U10693 (N_10693,N_9707,N_9694);
nand U10694 (N_10694,N_10217,N_10221);
or U10695 (N_10695,N_10007,N_10110);
xnor U10696 (N_10696,N_9892,N_9760);
nand U10697 (N_10697,N_10391,N_9989);
and U10698 (N_10698,N_9740,N_10322);
nand U10699 (N_10699,N_9885,N_9947);
nor U10700 (N_10700,N_10261,N_9979);
nor U10701 (N_10701,N_9869,N_9766);
nor U10702 (N_10702,N_9713,N_10194);
nand U10703 (N_10703,N_10161,N_9730);
nor U10704 (N_10704,N_9681,N_10293);
xor U10705 (N_10705,N_9845,N_10392);
xnor U10706 (N_10706,N_10186,N_9964);
or U10707 (N_10707,N_10362,N_10219);
and U10708 (N_10708,N_9664,N_10039);
nor U10709 (N_10709,N_10044,N_9709);
and U10710 (N_10710,N_9671,N_10390);
or U10711 (N_10711,N_9612,N_9926);
nand U10712 (N_10712,N_10200,N_10255);
and U10713 (N_10713,N_9872,N_9909);
or U10714 (N_10714,N_9622,N_10349);
nor U10715 (N_10715,N_9920,N_10286);
xnor U10716 (N_10716,N_9645,N_9684);
or U10717 (N_10717,N_10337,N_10103);
and U10718 (N_10718,N_10032,N_9810);
nor U10719 (N_10719,N_10093,N_9714);
and U10720 (N_10720,N_9634,N_10262);
and U10721 (N_10721,N_10222,N_10356);
nor U10722 (N_10722,N_9982,N_10280);
nand U10723 (N_10723,N_9789,N_10070);
xnor U10724 (N_10724,N_9911,N_9607);
nor U10725 (N_10725,N_9963,N_10384);
and U10726 (N_10726,N_10023,N_9880);
or U10727 (N_10727,N_9759,N_10326);
and U10728 (N_10728,N_9956,N_9624);
nand U10729 (N_10729,N_9726,N_10147);
or U10730 (N_10730,N_10294,N_9940);
nor U10731 (N_10731,N_9604,N_9666);
and U10732 (N_10732,N_9738,N_10162);
or U10733 (N_10733,N_9702,N_9734);
xnor U10734 (N_10734,N_9611,N_9966);
or U10735 (N_10735,N_10134,N_10047);
xor U10736 (N_10736,N_10059,N_10119);
nor U10737 (N_10737,N_10124,N_10201);
xnor U10738 (N_10738,N_10053,N_10302);
nand U10739 (N_10739,N_10167,N_10399);
xnor U10740 (N_10740,N_10283,N_10353);
and U10741 (N_10741,N_9749,N_9737);
or U10742 (N_10742,N_10207,N_9836);
nand U10743 (N_10743,N_9724,N_10382);
xor U10744 (N_10744,N_9631,N_9716);
and U10745 (N_10745,N_9786,N_9703);
nand U10746 (N_10746,N_9742,N_9807);
xnor U10747 (N_10747,N_9897,N_10018);
nor U10748 (N_10748,N_9834,N_9842);
nand U10749 (N_10749,N_9638,N_9767);
or U10750 (N_10750,N_10354,N_10395);
and U10751 (N_10751,N_10266,N_9686);
and U10752 (N_10752,N_9602,N_9678);
xnor U10753 (N_10753,N_10173,N_10352);
or U10754 (N_10754,N_9993,N_9826);
nand U10755 (N_10755,N_9662,N_10398);
or U10756 (N_10756,N_10054,N_9895);
nor U10757 (N_10757,N_10305,N_9900);
and U10758 (N_10758,N_10106,N_9668);
and U10759 (N_10759,N_9613,N_10331);
nand U10760 (N_10760,N_10136,N_10292);
or U10761 (N_10761,N_9913,N_10083);
or U10762 (N_10762,N_9865,N_10394);
nand U10763 (N_10763,N_10154,N_9927);
nand U10764 (N_10764,N_9795,N_10324);
and U10765 (N_10765,N_9955,N_10064);
and U10766 (N_10766,N_9735,N_10189);
and U10767 (N_10767,N_9931,N_10042);
nor U10768 (N_10768,N_9788,N_10278);
and U10769 (N_10769,N_10369,N_9874);
nand U10770 (N_10770,N_9906,N_9804);
nor U10771 (N_10771,N_10363,N_10008);
or U10772 (N_10772,N_10263,N_9700);
and U10773 (N_10773,N_9935,N_9609);
and U10774 (N_10774,N_10031,N_10016);
nand U10775 (N_10775,N_10151,N_10063);
and U10776 (N_10776,N_9898,N_9646);
nand U10777 (N_10777,N_9794,N_9600);
xor U10778 (N_10778,N_9674,N_9660);
or U10779 (N_10779,N_9673,N_10155);
and U10780 (N_10780,N_10078,N_9930);
xor U10781 (N_10781,N_9758,N_9852);
or U10782 (N_10782,N_10180,N_9917);
xnor U10783 (N_10783,N_9719,N_10081);
or U10784 (N_10784,N_10117,N_9778);
nand U10785 (N_10785,N_10311,N_9644);
nor U10786 (N_10786,N_9755,N_10206);
xor U10787 (N_10787,N_9912,N_9884);
or U10788 (N_10788,N_10340,N_10372);
or U10789 (N_10789,N_9772,N_10328);
and U10790 (N_10790,N_10148,N_9829);
nand U10791 (N_10791,N_9762,N_9608);
xnor U10792 (N_10792,N_10303,N_10301);
nor U10793 (N_10793,N_9896,N_9751);
xor U10794 (N_10794,N_9680,N_9771);
nor U10795 (N_10795,N_9890,N_10012);
or U10796 (N_10796,N_9736,N_9903);
and U10797 (N_10797,N_10329,N_10082);
and U10798 (N_10798,N_10181,N_9996);
nand U10799 (N_10799,N_9978,N_10140);
nand U10800 (N_10800,N_10098,N_10328);
or U10801 (N_10801,N_9851,N_9964);
and U10802 (N_10802,N_9988,N_10394);
and U10803 (N_10803,N_9922,N_10364);
and U10804 (N_10804,N_9886,N_9829);
xor U10805 (N_10805,N_9669,N_9769);
nor U10806 (N_10806,N_10310,N_9614);
xnor U10807 (N_10807,N_9883,N_9794);
nand U10808 (N_10808,N_10081,N_9614);
xnor U10809 (N_10809,N_9952,N_9722);
nor U10810 (N_10810,N_9721,N_9766);
and U10811 (N_10811,N_10206,N_9998);
or U10812 (N_10812,N_10216,N_9870);
and U10813 (N_10813,N_9624,N_9618);
nor U10814 (N_10814,N_9853,N_9870);
xnor U10815 (N_10815,N_10316,N_10087);
nor U10816 (N_10816,N_9643,N_10359);
or U10817 (N_10817,N_9965,N_10102);
nor U10818 (N_10818,N_10200,N_10066);
and U10819 (N_10819,N_9987,N_10048);
and U10820 (N_10820,N_9620,N_10109);
and U10821 (N_10821,N_9918,N_10221);
nand U10822 (N_10822,N_9901,N_10295);
and U10823 (N_10823,N_9982,N_9772);
xnor U10824 (N_10824,N_9890,N_9729);
xor U10825 (N_10825,N_9796,N_10220);
nand U10826 (N_10826,N_10044,N_9929);
nor U10827 (N_10827,N_9915,N_9922);
nand U10828 (N_10828,N_10047,N_10121);
nand U10829 (N_10829,N_10362,N_10107);
nor U10830 (N_10830,N_9898,N_10251);
nand U10831 (N_10831,N_10211,N_10287);
nand U10832 (N_10832,N_9891,N_10285);
xor U10833 (N_10833,N_10004,N_9763);
or U10834 (N_10834,N_10199,N_10030);
nor U10835 (N_10835,N_9605,N_9619);
nor U10836 (N_10836,N_10162,N_9604);
and U10837 (N_10837,N_9708,N_10215);
nand U10838 (N_10838,N_10093,N_10294);
or U10839 (N_10839,N_9749,N_9767);
or U10840 (N_10840,N_10284,N_10370);
nor U10841 (N_10841,N_9794,N_10375);
nor U10842 (N_10842,N_9901,N_9636);
and U10843 (N_10843,N_10103,N_10007);
and U10844 (N_10844,N_9788,N_9938);
nor U10845 (N_10845,N_10302,N_10205);
and U10846 (N_10846,N_9986,N_10039);
xnor U10847 (N_10847,N_10197,N_10229);
nand U10848 (N_10848,N_10152,N_9880);
nor U10849 (N_10849,N_9757,N_9746);
and U10850 (N_10850,N_10248,N_9945);
nor U10851 (N_10851,N_10111,N_10310);
or U10852 (N_10852,N_9879,N_10022);
nand U10853 (N_10853,N_9637,N_9964);
nor U10854 (N_10854,N_10099,N_10089);
or U10855 (N_10855,N_9830,N_10059);
nor U10856 (N_10856,N_10342,N_9855);
and U10857 (N_10857,N_9983,N_9721);
nor U10858 (N_10858,N_10157,N_9817);
xnor U10859 (N_10859,N_10330,N_9878);
nor U10860 (N_10860,N_10136,N_9963);
or U10861 (N_10861,N_9746,N_10278);
nand U10862 (N_10862,N_9720,N_10099);
nand U10863 (N_10863,N_9991,N_9971);
nand U10864 (N_10864,N_10322,N_10206);
and U10865 (N_10865,N_9752,N_10285);
xnor U10866 (N_10866,N_10023,N_9925);
nand U10867 (N_10867,N_9940,N_10090);
and U10868 (N_10868,N_9665,N_9893);
or U10869 (N_10869,N_10139,N_9600);
and U10870 (N_10870,N_10229,N_10394);
nand U10871 (N_10871,N_10167,N_10081);
nor U10872 (N_10872,N_10217,N_9890);
and U10873 (N_10873,N_9808,N_9705);
nor U10874 (N_10874,N_10393,N_10371);
nand U10875 (N_10875,N_10016,N_10363);
nand U10876 (N_10876,N_10039,N_10069);
and U10877 (N_10877,N_10241,N_10341);
nand U10878 (N_10878,N_9965,N_9937);
xnor U10879 (N_10879,N_10337,N_9900);
nor U10880 (N_10880,N_10084,N_9890);
or U10881 (N_10881,N_9941,N_9869);
or U10882 (N_10882,N_9831,N_10055);
nand U10883 (N_10883,N_10240,N_10079);
nor U10884 (N_10884,N_9977,N_9745);
xnor U10885 (N_10885,N_10368,N_9796);
nand U10886 (N_10886,N_9630,N_10382);
xor U10887 (N_10887,N_10237,N_9882);
nand U10888 (N_10888,N_10246,N_9628);
or U10889 (N_10889,N_9824,N_9882);
nand U10890 (N_10890,N_10294,N_9807);
xnor U10891 (N_10891,N_10179,N_9660);
nor U10892 (N_10892,N_9753,N_9913);
nor U10893 (N_10893,N_9910,N_10391);
nand U10894 (N_10894,N_10140,N_9725);
nor U10895 (N_10895,N_10357,N_10107);
nor U10896 (N_10896,N_9763,N_9953);
nand U10897 (N_10897,N_9702,N_9713);
or U10898 (N_10898,N_10396,N_9990);
xnor U10899 (N_10899,N_10321,N_10234);
or U10900 (N_10900,N_9776,N_9783);
or U10901 (N_10901,N_9999,N_10394);
nand U10902 (N_10902,N_10293,N_10189);
xnor U10903 (N_10903,N_10223,N_10138);
nor U10904 (N_10904,N_9682,N_9649);
xor U10905 (N_10905,N_10068,N_10295);
nor U10906 (N_10906,N_9731,N_9625);
and U10907 (N_10907,N_10360,N_10377);
nand U10908 (N_10908,N_10093,N_10135);
nor U10909 (N_10909,N_9952,N_9782);
xor U10910 (N_10910,N_10080,N_9906);
or U10911 (N_10911,N_10382,N_9647);
xnor U10912 (N_10912,N_9860,N_9831);
and U10913 (N_10913,N_10140,N_9911);
and U10914 (N_10914,N_10168,N_10135);
xnor U10915 (N_10915,N_10336,N_10034);
nor U10916 (N_10916,N_9724,N_9962);
nand U10917 (N_10917,N_10268,N_9684);
or U10918 (N_10918,N_9726,N_10275);
xnor U10919 (N_10919,N_9775,N_10266);
or U10920 (N_10920,N_9660,N_10139);
nor U10921 (N_10921,N_9867,N_10137);
and U10922 (N_10922,N_10003,N_10138);
xor U10923 (N_10923,N_10218,N_10034);
xnor U10924 (N_10924,N_10364,N_10249);
nand U10925 (N_10925,N_10230,N_10134);
and U10926 (N_10926,N_9626,N_10146);
or U10927 (N_10927,N_9891,N_10106);
xnor U10928 (N_10928,N_10252,N_10096);
nor U10929 (N_10929,N_10098,N_10045);
or U10930 (N_10930,N_9935,N_10315);
and U10931 (N_10931,N_9648,N_9644);
and U10932 (N_10932,N_9788,N_10276);
xor U10933 (N_10933,N_10229,N_9934);
or U10934 (N_10934,N_9607,N_9830);
nand U10935 (N_10935,N_9985,N_9877);
and U10936 (N_10936,N_9967,N_9637);
nor U10937 (N_10937,N_10245,N_10396);
nor U10938 (N_10938,N_10398,N_9831);
or U10939 (N_10939,N_10295,N_9662);
and U10940 (N_10940,N_10005,N_9944);
nand U10941 (N_10941,N_10030,N_9746);
xor U10942 (N_10942,N_10036,N_9999);
and U10943 (N_10943,N_10311,N_9748);
and U10944 (N_10944,N_10147,N_10142);
or U10945 (N_10945,N_9642,N_10284);
and U10946 (N_10946,N_9982,N_10311);
nand U10947 (N_10947,N_10060,N_10191);
nor U10948 (N_10948,N_10388,N_9754);
xnor U10949 (N_10949,N_9704,N_10385);
nor U10950 (N_10950,N_9895,N_10374);
nor U10951 (N_10951,N_9955,N_10110);
nand U10952 (N_10952,N_10187,N_9785);
nand U10953 (N_10953,N_10360,N_9920);
nor U10954 (N_10954,N_10266,N_10029);
and U10955 (N_10955,N_10106,N_10187);
and U10956 (N_10956,N_10350,N_10387);
or U10957 (N_10957,N_10263,N_10173);
or U10958 (N_10958,N_9975,N_9926);
nor U10959 (N_10959,N_9752,N_9917);
nor U10960 (N_10960,N_10250,N_10035);
xor U10961 (N_10961,N_9656,N_10331);
nor U10962 (N_10962,N_10250,N_9683);
and U10963 (N_10963,N_10326,N_9676);
nand U10964 (N_10964,N_10028,N_10066);
nand U10965 (N_10965,N_9719,N_10079);
xor U10966 (N_10966,N_10338,N_9856);
or U10967 (N_10967,N_9847,N_10093);
and U10968 (N_10968,N_9873,N_10358);
nor U10969 (N_10969,N_9646,N_10026);
xnor U10970 (N_10970,N_9624,N_9613);
nand U10971 (N_10971,N_10243,N_10337);
and U10972 (N_10972,N_9663,N_10235);
xnor U10973 (N_10973,N_10037,N_10341);
nor U10974 (N_10974,N_9756,N_10103);
xor U10975 (N_10975,N_10344,N_10193);
xor U10976 (N_10976,N_10394,N_9747);
or U10977 (N_10977,N_10330,N_9884);
or U10978 (N_10978,N_10366,N_9851);
nor U10979 (N_10979,N_10075,N_9939);
xor U10980 (N_10980,N_10016,N_9840);
nand U10981 (N_10981,N_9853,N_9801);
xnor U10982 (N_10982,N_9706,N_10384);
nor U10983 (N_10983,N_10068,N_9750);
and U10984 (N_10984,N_9749,N_9714);
and U10985 (N_10985,N_10111,N_10106);
xor U10986 (N_10986,N_9964,N_10166);
or U10987 (N_10987,N_10119,N_10394);
and U10988 (N_10988,N_10201,N_9994);
nand U10989 (N_10989,N_10089,N_9968);
and U10990 (N_10990,N_9621,N_9653);
or U10991 (N_10991,N_9730,N_10299);
and U10992 (N_10992,N_10216,N_10055);
xnor U10993 (N_10993,N_9918,N_10367);
nand U10994 (N_10994,N_10345,N_10381);
nand U10995 (N_10995,N_9945,N_9925);
nand U10996 (N_10996,N_10105,N_10177);
nand U10997 (N_10997,N_10275,N_10096);
xor U10998 (N_10998,N_9907,N_10113);
nor U10999 (N_10999,N_10164,N_9748);
nand U11000 (N_11000,N_9602,N_9626);
or U11001 (N_11001,N_9906,N_10199);
and U11002 (N_11002,N_10145,N_10233);
nand U11003 (N_11003,N_9600,N_9781);
nor U11004 (N_11004,N_9962,N_9831);
and U11005 (N_11005,N_9672,N_9653);
xor U11006 (N_11006,N_9852,N_10026);
or U11007 (N_11007,N_10328,N_10278);
xor U11008 (N_11008,N_9990,N_9780);
nor U11009 (N_11009,N_9735,N_10279);
and U11010 (N_11010,N_10094,N_9616);
xnor U11011 (N_11011,N_9645,N_9619);
nand U11012 (N_11012,N_9641,N_10213);
or U11013 (N_11013,N_9955,N_10343);
nand U11014 (N_11014,N_9614,N_10301);
xor U11015 (N_11015,N_9770,N_9877);
nor U11016 (N_11016,N_10374,N_10251);
nor U11017 (N_11017,N_9985,N_10376);
nor U11018 (N_11018,N_10189,N_10105);
or U11019 (N_11019,N_9730,N_10317);
nand U11020 (N_11020,N_9862,N_10188);
nand U11021 (N_11021,N_10208,N_10258);
xor U11022 (N_11022,N_10024,N_10040);
or U11023 (N_11023,N_10129,N_10122);
nor U11024 (N_11024,N_10363,N_10322);
or U11025 (N_11025,N_10320,N_10247);
xor U11026 (N_11026,N_10309,N_9817);
and U11027 (N_11027,N_10383,N_9945);
xor U11028 (N_11028,N_9891,N_9867);
and U11029 (N_11029,N_10053,N_9734);
and U11030 (N_11030,N_9673,N_9868);
or U11031 (N_11031,N_10115,N_10233);
or U11032 (N_11032,N_10371,N_10384);
and U11033 (N_11033,N_10361,N_10225);
nand U11034 (N_11034,N_10334,N_10176);
xnor U11035 (N_11035,N_10351,N_9962);
nor U11036 (N_11036,N_9838,N_10301);
nand U11037 (N_11037,N_10241,N_9945);
nor U11038 (N_11038,N_9942,N_9738);
nor U11039 (N_11039,N_9768,N_9761);
and U11040 (N_11040,N_9910,N_10093);
xor U11041 (N_11041,N_10230,N_9935);
nor U11042 (N_11042,N_10057,N_10053);
and U11043 (N_11043,N_10093,N_9923);
and U11044 (N_11044,N_10243,N_9783);
nand U11045 (N_11045,N_9950,N_9714);
nor U11046 (N_11046,N_10079,N_10377);
and U11047 (N_11047,N_10283,N_10206);
or U11048 (N_11048,N_9665,N_10363);
and U11049 (N_11049,N_10165,N_9618);
and U11050 (N_11050,N_10000,N_10250);
and U11051 (N_11051,N_9738,N_10089);
and U11052 (N_11052,N_10170,N_10221);
nand U11053 (N_11053,N_9739,N_10151);
nor U11054 (N_11054,N_10159,N_9855);
nand U11055 (N_11055,N_9976,N_9826);
nor U11056 (N_11056,N_10171,N_9774);
xor U11057 (N_11057,N_10168,N_10254);
or U11058 (N_11058,N_10331,N_9706);
xor U11059 (N_11059,N_10187,N_9622);
xnor U11060 (N_11060,N_10190,N_10281);
xor U11061 (N_11061,N_9726,N_10209);
or U11062 (N_11062,N_9855,N_9658);
nand U11063 (N_11063,N_10352,N_10287);
xor U11064 (N_11064,N_10211,N_10358);
and U11065 (N_11065,N_9923,N_9771);
nor U11066 (N_11066,N_10067,N_9911);
nor U11067 (N_11067,N_10128,N_10237);
nor U11068 (N_11068,N_9854,N_10275);
or U11069 (N_11069,N_10355,N_9931);
and U11070 (N_11070,N_9679,N_10063);
nand U11071 (N_11071,N_10286,N_10295);
or U11072 (N_11072,N_9879,N_10169);
nor U11073 (N_11073,N_10295,N_9610);
xor U11074 (N_11074,N_10261,N_10297);
and U11075 (N_11075,N_9854,N_9719);
or U11076 (N_11076,N_10110,N_9926);
xor U11077 (N_11077,N_10347,N_9704);
xnor U11078 (N_11078,N_10399,N_10055);
or U11079 (N_11079,N_9641,N_9779);
and U11080 (N_11080,N_9629,N_9993);
or U11081 (N_11081,N_9710,N_9832);
or U11082 (N_11082,N_10178,N_9787);
nand U11083 (N_11083,N_9875,N_10067);
nor U11084 (N_11084,N_9974,N_10162);
xnor U11085 (N_11085,N_10191,N_10275);
nor U11086 (N_11086,N_10367,N_10391);
or U11087 (N_11087,N_10012,N_10154);
or U11088 (N_11088,N_10323,N_10316);
nand U11089 (N_11089,N_9908,N_9817);
or U11090 (N_11090,N_10149,N_9914);
xnor U11091 (N_11091,N_10360,N_9742);
or U11092 (N_11092,N_10387,N_10253);
nor U11093 (N_11093,N_9974,N_10386);
nor U11094 (N_11094,N_10266,N_9886);
nor U11095 (N_11095,N_9968,N_9986);
xnor U11096 (N_11096,N_10227,N_10087);
nand U11097 (N_11097,N_9929,N_10220);
nand U11098 (N_11098,N_10358,N_10187);
or U11099 (N_11099,N_10046,N_10194);
and U11100 (N_11100,N_10206,N_9631);
nor U11101 (N_11101,N_10144,N_10188);
nand U11102 (N_11102,N_9877,N_10066);
or U11103 (N_11103,N_10129,N_9651);
and U11104 (N_11104,N_9896,N_9934);
xor U11105 (N_11105,N_10158,N_10037);
nor U11106 (N_11106,N_9661,N_9930);
and U11107 (N_11107,N_10257,N_9996);
xnor U11108 (N_11108,N_10322,N_10084);
or U11109 (N_11109,N_10255,N_9605);
xor U11110 (N_11110,N_9642,N_10391);
and U11111 (N_11111,N_10178,N_9909);
nand U11112 (N_11112,N_10144,N_9744);
and U11113 (N_11113,N_9817,N_10031);
or U11114 (N_11114,N_9668,N_9611);
xnor U11115 (N_11115,N_9656,N_10151);
and U11116 (N_11116,N_9924,N_10167);
nor U11117 (N_11117,N_10110,N_9689);
nor U11118 (N_11118,N_9916,N_9656);
or U11119 (N_11119,N_9890,N_9685);
and U11120 (N_11120,N_10076,N_9946);
nand U11121 (N_11121,N_9676,N_9721);
xnor U11122 (N_11122,N_9826,N_10380);
nor U11123 (N_11123,N_10113,N_9949);
and U11124 (N_11124,N_9647,N_10112);
nand U11125 (N_11125,N_10060,N_9699);
nand U11126 (N_11126,N_9703,N_9744);
nor U11127 (N_11127,N_10042,N_10139);
nand U11128 (N_11128,N_10358,N_9976);
and U11129 (N_11129,N_10003,N_9805);
nor U11130 (N_11130,N_9885,N_9972);
or U11131 (N_11131,N_9956,N_9812);
or U11132 (N_11132,N_10234,N_9908);
nor U11133 (N_11133,N_10238,N_10107);
or U11134 (N_11134,N_9816,N_10363);
nand U11135 (N_11135,N_9830,N_10290);
and U11136 (N_11136,N_10254,N_10011);
nand U11137 (N_11137,N_10096,N_9729);
and U11138 (N_11138,N_10357,N_9724);
and U11139 (N_11139,N_10058,N_9989);
xnor U11140 (N_11140,N_10176,N_9816);
and U11141 (N_11141,N_10330,N_10198);
nor U11142 (N_11142,N_10025,N_9976);
nand U11143 (N_11143,N_9923,N_9802);
nor U11144 (N_11144,N_9800,N_10083);
nand U11145 (N_11145,N_10125,N_10014);
nor U11146 (N_11146,N_9655,N_9988);
xor U11147 (N_11147,N_9849,N_9938);
or U11148 (N_11148,N_9886,N_10237);
and U11149 (N_11149,N_9841,N_10049);
and U11150 (N_11150,N_10329,N_10245);
nand U11151 (N_11151,N_10164,N_9640);
nand U11152 (N_11152,N_10100,N_9757);
or U11153 (N_11153,N_10013,N_9684);
or U11154 (N_11154,N_10331,N_10284);
and U11155 (N_11155,N_10268,N_9749);
nand U11156 (N_11156,N_10157,N_9809);
nor U11157 (N_11157,N_9606,N_9716);
and U11158 (N_11158,N_10255,N_9648);
and U11159 (N_11159,N_9714,N_9678);
xor U11160 (N_11160,N_10223,N_9621);
xor U11161 (N_11161,N_10155,N_9974);
and U11162 (N_11162,N_9775,N_9721);
and U11163 (N_11163,N_9702,N_9966);
nand U11164 (N_11164,N_9914,N_10040);
nand U11165 (N_11165,N_9711,N_10116);
and U11166 (N_11166,N_9628,N_10362);
nor U11167 (N_11167,N_10226,N_10376);
or U11168 (N_11168,N_9876,N_10080);
nand U11169 (N_11169,N_10047,N_10075);
nand U11170 (N_11170,N_9731,N_9795);
or U11171 (N_11171,N_10374,N_9933);
or U11172 (N_11172,N_10312,N_10169);
xor U11173 (N_11173,N_10058,N_10375);
or U11174 (N_11174,N_10166,N_9932);
or U11175 (N_11175,N_9884,N_10255);
and U11176 (N_11176,N_10092,N_10250);
or U11177 (N_11177,N_9677,N_9882);
nor U11178 (N_11178,N_10074,N_9996);
nand U11179 (N_11179,N_9717,N_10232);
xnor U11180 (N_11180,N_10277,N_10028);
or U11181 (N_11181,N_10088,N_9830);
or U11182 (N_11182,N_9636,N_9789);
nand U11183 (N_11183,N_10155,N_10361);
xnor U11184 (N_11184,N_10039,N_9875);
and U11185 (N_11185,N_10338,N_10190);
xnor U11186 (N_11186,N_9908,N_9949);
xnor U11187 (N_11187,N_9609,N_9920);
xor U11188 (N_11188,N_10344,N_9883);
nor U11189 (N_11189,N_10219,N_9726);
or U11190 (N_11190,N_10311,N_9723);
nand U11191 (N_11191,N_9929,N_10330);
nand U11192 (N_11192,N_10296,N_10051);
nor U11193 (N_11193,N_9794,N_9763);
or U11194 (N_11194,N_9883,N_10265);
and U11195 (N_11195,N_10114,N_10080);
or U11196 (N_11196,N_9911,N_10256);
nand U11197 (N_11197,N_10151,N_9966);
or U11198 (N_11198,N_10223,N_9890);
and U11199 (N_11199,N_10309,N_10316);
nor U11200 (N_11200,N_10971,N_11074);
nor U11201 (N_11201,N_11050,N_10848);
nor U11202 (N_11202,N_10824,N_10610);
and U11203 (N_11203,N_11151,N_11189);
nor U11204 (N_11204,N_10537,N_10573);
nor U11205 (N_11205,N_10995,N_10810);
or U11206 (N_11206,N_10613,N_11055);
xnor U11207 (N_11207,N_10794,N_10567);
and U11208 (N_11208,N_10885,N_10570);
nor U11209 (N_11209,N_10747,N_10770);
nand U11210 (N_11210,N_10727,N_10898);
xnor U11211 (N_11211,N_10990,N_10560);
nand U11212 (N_11212,N_11065,N_11007);
or U11213 (N_11213,N_10685,N_11030);
and U11214 (N_11214,N_11168,N_10498);
xnor U11215 (N_11215,N_11076,N_10458);
xor U11216 (N_11216,N_10452,N_10923);
nor U11217 (N_11217,N_10638,N_10936);
nor U11218 (N_11218,N_10787,N_10412);
xnor U11219 (N_11219,N_10797,N_11122);
nand U11220 (N_11220,N_11057,N_10840);
and U11221 (N_11221,N_10562,N_10514);
nor U11222 (N_11222,N_10531,N_10738);
nor U11223 (N_11223,N_10623,N_10825);
nor U11224 (N_11224,N_10664,N_10521);
nor U11225 (N_11225,N_10742,N_11047);
nand U11226 (N_11226,N_10547,N_10808);
nand U11227 (N_11227,N_10748,N_10558);
or U11228 (N_11228,N_11099,N_10981);
and U11229 (N_11229,N_11004,N_11022);
and U11230 (N_11230,N_10687,N_11128);
and U11231 (N_11231,N_10652,N_10832);
nor U11232 (N_11232,N_10488,N_10499);
and U11233 (N_11233,N_10597,N_10855);
or U11234 (N_11234,N_10965,N_10993);
and U11235 (N_11235,N_11166,N_10453);
xor U11236 (N_11236,N_11023,N_10809);
nor U11237 (N_11237,N_10639,N_10674);
and U11238 (N_11238,N_10921,N_10725);
and U11239 (N_11239,N_10582,N_10774);
or U11240 (N_11240,N_10868,N_10900);
xnor U11241 (N_11241,N_10649,N_11193);
xor U11242 (N_11242,N_10670,N_11124);
or U11243 (N_11243,N_10622,N_10489);
nand U11244 (N_11244,N_10625,N_11001);
xor U11245 (N_11245,N_11160,N_10451);
xnor U11246 (N_11246,N_10538,N_10791);
or U11247 (N_11247,N_10549,N_11186);
and U11248 (N_11248,N_10543,N_11086);
nor U11249 (N_11249,N_10927,N_10686);
and U11250 (N_11250,N_11080,N_10946);
nand U11251 (N_11251,N_10873,N_11083);
or U11252 (N_11252,N_10944,N_10910);
and U11253 (N_11253,N_10853,N_10542);
xor U11254 (N_11254,N_10804,N_10539);
xor U11255 (N_11255,N_11053,N_10765);
and U11256 (N_11256,N_11103,N_10554);
or U11257 (N_11257,N_11015,N_10906);
xnor U11258 (N_11258,N_10572,N_11087);
nor U11259 (N_11259,N_11040,N_10533);
nor U11260 (N_11260,N_10651,N_10422);
nand U11261 (N_11261,N_11106,N_10614);
xnor U11262 (N_11262,N_10595,N_10475);
xor U11263 (N_11263,N_10999,N_10964);
and U11264 (N_11264,N_10856,N_10411);
nand U11265 (N_11265,N_10659,N_10786);
and U11266 (N_11266,N_10561,N_11070);
and U11267 (N_11267,N_11131,N_10783);
xnor U11268 (N_11268,N_10496,N_10520);
nor U11269 (N_11269,N_10550,N_10681);
and U11270 (N_11270,N_11085,N_10829);
or U11271 (N_11271,N_11028,N_11036);
nand U11272 (N_11272,N_11044,N_10979);
nor U11273 (N_11273,N_10544,N_10933);
xnor U11274 (N_11274,N_10878,N_10517);
nand U11275 (N_11275,N_10506,N_10860);
and U11276 (N_11276,N_11164,N_10996);
nand U11277 (N_11277,N_10581,N_10896);
nand U11278 (N_11278,N_10821,N_10519);
or U11279 (N_11279,N_10468,N_10704);
xor U11280 (N_11280,N_10799,N_10823);
and U11281 (N_11281,N_11051,N_10780);
nand U11282 (N_11282,N_10525,N_10590);
nor U11283 (N_11283,N_11126,N_10857);
xnor U11284 (N_11284,N_10526,N_10974);
xor U11285 (N_11285,N_10769,N_10679);
nor U11286 (N_11286,N_10424,N_10417);
nand U11287 (N_11287,N_10509,N_10492);
or U11288 (N_11288,N_10830,N_10414);
nor U11289 (N_11289,N_10881,N_10487);
and U11290 (N_11290,N_10564,N_10958);
nor U11291 (N_11291,N_10793,N_10925);
nor U11292 (N_11292,N_10715,N_10819);
nor U11293 (N_11293,N_11066,N_10407);
nor U11294 (N_11294,N_10655,N_11109);
nand U11295 (N_11295,N_10998,N_11125);
xnor U11296 (N_11296,N_10973,N_11174);
nand U11297 (N_11297,N_10888,N_10696);
nor U11298 (N_11298,N_10739,N_11120);
nor U11299 (N_11299,N_10680,N_10763);
nor U11300 (N_11300,N_11115,N_10557);
nand U11301 (N_11301,N_11182,N_10922);
nand U11302 (N_11302,N_10419,N_11187);
or U11303 (N_11303,N_10400,N_10456);
nor U11304 (N_11304,N_10800,N_11180);
nand U11305 (N_11305,N_10816,N_10524);
or U11306 (N_11306,N_11133,N_10629);
or U11307 (N_11307,N_10694,N_10482);
nor U11308 (N_11308,N_10477,N_10504);
xnor U11309 (N_11309,N_11056,N_10476);
nor U11310 (N_11310,N_10445,N_10940);
xnor U11311 (N_11311,N_11017,N_10527);
nand U11312 (N_11312,N_11042,N_11197);
nor U11313 (N_11313,N_10919,N_10720);
and U11314 (N_11314,N_10471,N_11154);
xor U11315 (N_11315,N_11153,N_10512);
xnor U11316 (N_11316,N_10632,N_10448);
nand U11317 (N_11317,N_10728,N_10437);
or U11318 (N_11318,N_10712,N_10796);
nand U11319 (N_11319,N_11048,N_10884);
xor U11320 (N_11320,N_10457,N_10608);
and U11321 (N_11321,N_11091,N_10510);
nor U11322 (N_11322,N_10569,N_11037);
or U11323 (N_11323,N_10460,N_10425);
nor U11324 (N_11324,N_10501,N_10603);
nand U11325 (N_11325,N_11069,N_11142);
and U11326 (N_11326,N_10784,N_10523);
nand U11327 (N_11327,N_10441,N_10917);
nor U11328 (N_11328,N_11146,N_10935);
nor U11329 (N_11329,N_10650,N_10483);
xor U11330 (N_11330,N_10740,N_11198);
xor U11331 (N_11331,N_10751,N_10676);
and U11332 (N_11332,N_10426,N_10536);
or U11333 (N_11333,N_10931,N_11046);
nand U11334 (N_11334,N_11071,N_10469);
xor U11335 (N_11335,N_10478,N_10630);
nand U11336 (N_11336,N_10644,N_10418);
nand U11337 (N_11337,N_11184,N_10886);
nor U11338 (N_11338,N_10427,N_11096);
nor U11339 (N_11339,N_10421,N_11090);
xnor U11340 (N_11340,N_10963,N_10930);
or U11341 (N_11341,N_10677,N_10773);
nand U11342 (N_11342,N_11190,N_10594);
or U11343 (N_11343,N_10463,N_10907);
and U11344 (N_11344,N_10897,N_10513);
nand U11345 (N_11345,N_11008,N_10975);
or U11346 (N_11346,N_11104,N_11029);
nor U11347 (N_11347,N_10473,N_10953);
xor U11348 (N_11348,N_10420,N_11110);
and U11349 (N_11349,N_11199,N_11191);
and U11350 (N_11350,N_10802,N_10874);
nor U11351 (N_11351,N_11163,N_10472);
nor U11352 (N_11352,N_11033,N_10502);
and U11353 (N_11353,N_10838,N_10682);
xnor U11354 (N_11354,N_10503,N_10444);
nor U11355 (N_11355,N_11075,N_11107);
or U11356 (N_11356,N_11060,N_10675);
nor U11357 (N_11357,N_11116,N_10972);
nand U11358 (N_11358,N_10699,N_10852);
and U11359 (N_11359,N_10495,N_10586);
nor U11360 (N_11360,N_10491,N_10508);
and U11361 (N_11361,N_10969,N_10841);
nor U11362 (N_11362,N_10869,N_11171);
nand U11363 (N_11363,N_10455,N_10654);
nand U11364 (N_11364,N_11192,N_10929);
and U11365 (N_11365,N_10436,N_11097);
or U11366 (N_11366,N_10815,N_10534);
or U11367 (N_11367,N_10835,N_10661);
nand U11368 (N_11368,N_10845,N_10693);
and U11369 (N_11369,N_11195,N_10788);
xnor U11370 (N_11370,N_10552,N_10833);
xor U11371 (N_11371,N_10920,N_10474);
or U11372 (N_11372,N_11135,N_11167);
nor U11373 (N_11373,N_10530,N_10859);
nor U11374 (N_11374,N_10813,N_10689);
and U11375 (N_11375,N_10698,N_10647);
xnor U11376 (N_11376,N_10913,N_10605);
nand U11377 (N_11377,N_10924,N_10532);
or U11378 (N_11378,N_10620,N_10721);
xor U11379 (N_11379,N_10901,N_10575);
nand U11380 (N_11380,N_10673,N_10870);
nor U11381 (N_11381,N_11144,N_10580);
and U11382 (N_11382,N_10609,N_10977);
xnor U11383 (N_11383,N_10970,N_11119);
xnor U11384 (N_11384,N_10589,N_11121);
and U11385 (N_11385,N_10961,N_10954);
or U11386 (N_11386,N_11059,N_10548);
and U11387 (N_11387,N_11155,N_10541);
xor U11388 (N_11388,N_11019,N_10507);
xor U11389 (N_11389,N_10684,N_10805);
xnor U11390 (N_11390,N_10643,N_10872);
and U11391 (N_11391,N_10671,N_10565);
or U11392 (N_11392,N_10828,N_11134);
nand U11393 (N_11393,N_10743,N_10672);
xnor U11394 (N_11394,N_11009,N_10745);
nand U11395 (N_11395,N_11118,N_10827);
nor U11396 (N_11396,N_10415,N_10741);
and U11397 (N_11397,N_10576,N_10776);
nand U11398 (N_11398,N_10812,N_10493);
nor U11399 (N_11399,N_10540,N_11170);
nor U11400 (N_11400,N_10571,N_11188);
nand U11401 (N_11401,N_10811,N_10706);
nand U11402 (N_11402,N_10432,N_10546);
and U11403 (N_11403,N_10467,N_10967);
nand U11404 (N_11404,N_10834,N_10904);
xnor U11405 (N_11405,N_11039,N_10653);
nand U11406 (N_11406,N_10911,N_10749);
and U11407 (N_11407,N_10665,N_10591);
xnor U11408 (N_11408,N_10775,N_10405);
nand U11409 (N_11409,N_11123,N_10750);
or U11410 (N_11410,N_10968,N_11010);
xor U11411 (N_11411,N_10500,N_11088);
xnor U11412 (N_11412,N_10635,N_11035);
xnor U11413 (N_11413,N_11161,N_11077);
and U11414 (N_11414,N_10717,N_10984);
nand U11415 (N_11415,N_11005,N_10559);
and U11416 (N_11416,N_10615,N_10733);
and U11417 (N_11417,N_11178,N_10962);
nor U11418 (N_11418,N_10563,N_10657);
and U11419 (N_11419,N_10807,N_11100);
xor U11420 (N_11420,N_11145,N_11043);
or U11421 (N_11421,N_11058,N_11112);
nand U11422 (N_11422,N_11052,N_10566);
and U11423 (N_11423,N_10918,N_10875);
xor U11424 (N_11424,N_10994,N_10950);
xor U11425 (N_11425,N_10777,N_10450);
nand U11426 (N_11426,N_11049,N_10462);
nor U11427 (N_11427,N_10866,N_10636);
or U11428 (N_11428,N_10716,N_10801);
xnor U11429 (N_11429,N_11108,N_10883);
or U11430 (N_11430,N_10642,N_10849);
nor U11431 (N_11431,N_10817,N_10779);
or U11432 (N_11432,N_10583,N_10584);
xnor U11433 (N_11433,N_10666,N_11084);
and U11434 (N_11434,N_10645,N_11073);
xnor U11435 (N_11435,N_10756,N_10723);
and U11436 (N_11436,N_10772,N_11063);
nand U11437 (N_11437,N_10732,N_11194);
xor U11438 (N_11438,N_11067,N_11013);
nor U11439 (N_11439,N_10734,N_11137);
nand U11440 (N_11440,N_10934,N_10928);
and U11441 (N_11441,N_10978,N_10789);
and U11442 (N_11442,N_10795,N_10839);
nand U11443 (N_11443,N_11179,N_10568);
and U11444 (N_11444,N_10701,N_10843);
xor U11445 (N_11445,N_10966,N_10406);
or U11446 (N_11446,N_11177,N_10430);
nor U11447 (N_11447,N_10863,N_11003);
nand U11448 (N_11448,N_11102,N_11072);
nor U11449 (N_11449,N_10757,N_11141);
and U11450 (N_11450,N_10604,N_10939);
xor U11451 (N_11451,N_10577,N_11196);
xnor U11452 (N_11452,N_11175,N_10588);
nor U11453 (N_11453,N_10844,N_10470);
nor U11454 (N_11454,N_10447,N_10556);
and U11455 (N_11455,N_10465,N_10408);
nor U11456 (N_11456,N_10410,N_10952);
xor U11457 (N_11457,N_10709,N_10862);
and U11458 (N_11458,N_10461,N_10992);
and U11459 (N_11459,N_10606,N_10908);
nand U11460 (N_11460,N_10585,N_10616);
nand U11461 (N_11461,N_10663,N_10646);
xnor U11462 (N_11462,N_11000,N_10767);
xnor U11463 (N_11463,N_10454,N_10850);
xnor U11464 (N_11464,N_10440,N_11129);
nor U11465 (N_11465,N_10518,N_11127);
and U11466 (N_11466,N_10837,N_10707);
xor U11467 (N_11467,N_10915,N_10618);
xnor U11468 (N_11468,N_10882,N_10481);
xnor U11469 (N_11469,N_10718,N_10818);
xor U11470 (N_11470,N_11025,N_10867);
xnor U11471 (N_11471,N_10637,N_10433);
nor U11472 (N_11472,N_10435,N_10428);
nor U11473 (N_11473,N_10683,N_10755);
or U11474 (N_11474,N_10988,N_11089);
or U11475 (N_11475,N_10624,N_11098);
or U11476 (N_11476,N_11054,N_10710);
or U11477 (N_11477,N_10485,N_11027);
nand U11478 (N_11478,N_11114,N_10889);
xor U11479 (N_11479,N_10627,N_10690);
nor U11480 (N_11480,N_10985,N_11011);
and U11481 (N_11481,N_11152,N_10439);
or U11482 (N_11482,N_11159,N_10758);
and U11483 (N_11483,N_11078,N_10402);
nor U11484 (N_11484,N_10497,N_10768);
nand U11485 (N_11485,N_10887,N_10617);
or U11486 (N_11486,N_10714,N_10658);
or U11487 (N_11487,N_11113,N_11062);
xor U11488 (N_11488,N_11138,N_10865);
xnor U11489 (N_11489,N_10941,N_10842);
or U11490 (N_11490,N_10790,N_10692);
or U11491 (N_11491,N_10737,N_10434);
xnor U11492 (N_11492,N_10724,N_10416);
or U11493 (N_11493,N_10895,N_11024);
and U11494 (N_11494,N_10806,N_10633);
xor U11495 (N_11495,N_10551,N_10753);
nand U11496 (N_11496,N_11079,N_10631);
xor U11497 (N_11497,N_11181,N_10942);
nand U11498 (N_11498,N_11140,N_10822);
xor U11499 (N_11499,N_10648,N_10555);
nand U11500 (N_11500,N_10484,N_11014);
or U11501 (N_11501,N_11034,N_10754);
or U11502 (N_11502,N_10621,N_10997);
nand U11503 (N_11503,N_10916,N_10516);
nand U11504 (N_11504,N_10700,N_10957);
and U11505 (N_11505,N_11064,N_10893);
or U11506 (N_11506,N_10814,N_11169);
nor U11507 (N_11507,N_10719,N_10667);
nor U11508 (N_11508,N_10836,N_10449);
nand U11509 (N_11509,N_10600,N_10820);
nand U11510 (N_11510,N_10892,N_11038);
and U11511 (N_11511,N_11185,N_10535);
and U11512 (N_11512,N_10697,N_10669);
and U11513 (N_11513,N_10932,N_10660);
nor U11514 (N_11514,N_11183,N_10599);
xnor U11515 (N_11515,N_10596,N_10785);
or U11516 (N_11516,N_10744,N_10778);
or U11517 (N_11517,N_11158,N_10731);
or U11518 (N_11518,N_10826,N_10735);
nor U11519 (N_11519,N_10401,N_10713);
or U11520 (N_11520,N_10986,N_10947);
and U11521 (N_11521,N_10879,N_10914);
nand U11522 (N_11522,N_10601,N_10607);
xor U11523 (N_11523,N_11172,N_10983);
or U11524 (N_11524,N_10634,N_10522);
or U11525 (N_11525,N_10762,N_10443);
and U11526 (N_11526,N_10423,N_10545);
nand U11527 (N_11527,N_11149,N_10959);
and U11528 (N_11528,N_10956,N_10909);
xnor U11529 (N_11529,N_10708,N_10851);
and U11530 (N_11530,N_10987,N_10876);
nor U11531 (N_11531,N_11093,N_11032);
xnor U11532 (N_11532,N_10592,N_10766);
xor U11533 (N_11533,N_10553,N_11061);
and U11534 (N_11534,N_10691,N_10578);
xnor U11535 (N_11535,N_10409,N_10949);
and U11536 (N_11536,N_11148,N_11117);
and U11537 (N_11537,N_10429,N_10702);
nor U11538 (N_11538,N_10459,N_10515);
and U11539 (N_11539,N_10529,N_11082);
and U11540 (N_11540,N_10494,N_11002);
or U11541 (N_11541,N_10943,N_10899);
xnor U11542 (N_11542,N_11094,N_11031);
nand U11543 (N_11543,N_10688,N_10880);
or U11544 (N_11544,N_10890,N_10528);
and U11545 (N_11545,N_10640,N_11157);
nor U11546 (N_11546,N_10937,N_10431);
or U11547 (N_11547,N_10877,N_10511);
nand U11548 (N_11548,N_10480,N_11139);
and U11549 (N_11549,N_10760,N_10960);
nor U11550 (N_11550,N_11132,N_10695);
xnor U11551 (N_11551,N_10579,N_10759);
xor U11552 (N_11552,N_10764,N_11045);
nor U11553 (N_11553,N_11068,N_10490);
nor U11554 (N_11554,N_10991,N_11162);
xor U11555 (N_11555,N_10926,N_10861);
or U11556 (N_11556,N_10442,N_10611);
xor U11557 (N_11557,N_11092,N_10722);
nand U11558 (N_11558,N_10711,N_10854);
and U11559 (N_11559,N_10466,N_11143);
nor U11560 (N_11560,N_11176,N_10782);
nor U11561 (N_11561,N_11101,N_10479);
or U11562 (N_11562,N_10404,N_11165);
and U11563 (N_11563,N_10982,N_10792);
nor U11564 (N_11564,N_11150,N_10703);
nor U11565 (N_11565,N_11105,N_10746);
or U11566 (N_11566,N_11136,N_10668);
xnor U11567 (N_11567,N_10871,N_10619);
xnor U11568 (N_11568,N_10938,N_11095);
or U11569 (N_11569,N_10612,N_10976);
nor U11570 (N_11570,N_10951,N_10403);
and U11571 (N_11571,N_10593,N_10574);
or U11572 (N_11572,N_10955,N_11016);
xor U11573 (N_11573,N_10847,N_10464);
and U11574 (N_11574,N_10903,N_10626);
xor U11575 (N_11575,N_10894,N_10705);
or U11576 (N_11576,N_10587,N_10803);
or U11577 (N_11577,N_10781,N_10864);
nand U11578 (N_11578,N_10831,N_11156);
or U11579 (N_11579,N_10730,N_10736);
or U11580 (N_11580,N_10438,N_10891);
or U11581 (N_11581,N_11081,N_11020);
and U11582 (N_11582,N_10446,N_10761);
and U11583 (N_11583,N_10912,N_10729);
nand U11584 (N_11584,N_11173,N_11111);
nor U11585 (N_11585,N_10902,N_10752);
or U11586 (N_11586,N_10905,N_11147);
and U11587 (N_11587,N_10678,N_11012);
nor U11588 (N_11588,N_10771,N_10726);
and U11589 (N_11589,N_10662,N_11041);
or U11590 (N_11590,N_10628,N_10641);
and U11591 (N_11591,N_11026,N_10798);
xor U11592 (N_11592,N_10846,N_10989);
nor U11593 (N_11593,N_10505,N_11130);
nand U11594 (N_11594,N_10656,N_10948);
and U11595 (N_11595,N_10980,N_11018);
and U11596 (N_11596,N_11021,N_10598);
xnor U11597 (N_11597,N_10413,N_10858);
and U11598 (N_11598,N_10945,N_10486);
or U11599 (N_11599,N_11006,N_10602);
xnor U11600 (N_11600,N_11032,N_10928);
and U11601 (N_11601,N_10643,N_10714);
xor U11602 (N_11602,N_10696,N_10462);
or U11603 (N_11603,N_10462,N_10686);
xor U11604 (N_11604,N_10941,N_11049);
or U11605 (N_11605,N_10718,N_10485);
or U11606 (N_11606,N_11146,N_10585);
nand U11607 (N_11607,N_11178,N_10955);
nor U11608 (N_11608,N_10756,N_10684);
or U11609 (N_11609,N_11091,N_10666);
or U11610 (N_11610,N_10977,N_11047);
or U11611 (N_11611,N_10914,N_10430);
nand U11612 (N_11612,N_10930,N_10469);
xnor U11613 (N_11613,N_10749,N_11144);
and U11614 (N_11614,N_10823,N_10939);
or U11615 (N_11615,N_11082,N_10625);
nor U11616 (N_11616,N_10446,N_11122);
or U11617 (N_11617,N_10466,N_10683);
and U11618 (N_11618,N_10546,N_10775);
nor U11619 (N_11619,N_10647,N_10539);
and U11620 (N_11620,N_11138,N_10756);
nor U11621 (N_11621,N_10441,N_11118);
or U11622 (N_11622,N_10605,N_10998);
and U11623 (N_11623,N_11065,N_10903);
or U11624 (N_11624,N_11011,N_10801);
or U11625 (N_11625,N_10550,N_11126);
xor U11626 (N_11626,N_10690,N_10415);
xnor U11627 (N_11627,N_11039,N_10505);
xor U11628 (N_11628,N_10580,N_10567);
nor U11629 (N_11629,N_11071,N_10813);
and U11630 (N_11630,N_10508,N_11178);
xor U11631 (N_11631,N_10435,N_10967);
xnor U11632 (N_11632,N_10649,N_10425);
nand U11633 (N_11633,N_11083,N_10584);
xnor U11634 (N_11634,N_10756,N_11174);
and U11635 (N_11635,N_10887,N_11109);
xnor U11636 (N_11636,N_10670,N_10848);
xnor U11637 (N_11637,N_10501,N_11106);
nand U11638 (N_11638,N_10753,N_10954);
nand U11639 (N_11639,N_10675,N_10728);
or U11640 (N_11640,N_10552,N_10436);
nand U11641 (N_11641,N_11023,N_10790);
nand U11642 (N_11642,N_10512,N_10702);
or U11643 (N_11643,N_11165,N_11011);
xnor U11644 (N_11644,N_10515,N_10765);
nand U11645 (N_11645,N_11138,N_10662);
xor U11646 (N_11646,N_10944,N_10419);
xor U11647 (N_11647,N_10965,N_10428);
nor U11648 (N_11648,N_11124,N_10496);
or U11649 (N_11649,N_11163,N_11093);
or U11650 (N_11650,N_10450,N_11103);
and U11651 (N_11651,N_10735,N_11060);
or U11652 (N_11652,N_10848,N_10641);
or U11653 (N_11653,N_10711,N_10570);
or U11654 (N_11654,N_10811,N_10582);
and U11655 (N_11655,N_10959,N_11076);
nand U11656 (N_11656,N_10746,N_10458);
nor U11657 (N_11657,N_11038,N_10490);
or U11658 (N_11658,N_10633,N_10510);
and U11659 (N_11659,N_10723,N_11102);
nand U11660 (N_11660,N_10961,N_11053);
xnor U11661 (N_11661,N_10685,N_11037);
and U11662 (N_11662,N_11123,N_10914);
or U11663 (N_11663,N_11118,N_10781);
nand U11664 (N_11664,N_11063,N_11174);
xor U11665 (N_11665,N_10482,N_11158);
nor U11666 (N_11666,N_11044,N_10531);
and U11667 (N_11667,N_10730,N_10932);
and U11668 (N_11668,N_11139,N_10924);
nand U11669 (N_11669,N_10435,N_10491);
or U11670 (N_11670,N_11047,N_10775);
nor U11671 (N_11671,N_10692,N_11135);
nand U11672 (N_11672,N_10601,N_11033);
nand U11673 (N_11673,N_10856,N_11127);
nor U11674 (N_11674,N_10955,N_10909);
xor U11675 (N_11675,N_10860,N_11071);
xnor U11676 (N_11676,N_10919,N_11132);
nor U11677 (N_11677,N_10865,N_10838);
xor U11678 (N_11678,N_11010,N_10493);
xnor U11679 (N_11679,N_11082,N_10454);
or U11680 (N_11680,N_10872,N_11049);
nand U11681 (N_11681,N_10701,N_10511);
and U11682 (N_11682,N_10731,N_10942);
nand U11683 (N_11683,N_10597,N_10658);
nor U11684 (N_11684,N_11143,N_10535);
xor U11685 (N_11685,N_10920,N_10770);
xor U11686 (N_11686,N_10808,N_10406);
and U11687 (N_11687,N_11187,N_10739);
xor U11688 (N_11688,N_10631,N_10812);
and U11689 (N_11689,N_11036,N_10506);
and U11690 (N_11690,N_10473,N_10761);
xor U11691 (N_11691,N_11077,N_11104);
nor U11692 (N_11692,N_10928,N_10445);
xor U11693 (N_11693,N_10706,N_10900);
nand U11694 (N_11694,N_10777,N_10669);
nand U11695 (N_11695,N_10456,N_10669);
and U11696 (N_11696,N_10750,N_10894);
or U11697 (N_11697,N_10868,N_10866);
and U11698 (N_11698,N_10480,N_10544);
or U11699 (N_11699,N_10468,N_10496);
or U11700 (N_11700,N_10495,N_10400);
nor U11701 (N_11701,N_11153,N_10778);
and U11702 (N_11702,N_10742,N_10887);
nand U11703 (N_11703,N_11152,N_10995);
nand U11704 (N_11704,N_10944,N_11150);
nand U11705 (N_11705,N_10739,N_10998);
or U11706 (N_11706,N_10474,N_11084);
or U11707 (N_11707,N_10583,N_11058);
and U11708 (N_11708,N_10671,N_10998);
or U11709 (N_11709,N_10819,N_11004);
nor U11710 (N_11710,N_10761,N_10835);
or U11711 (N_11711,N_10791,N_10595);
nor U11712 (N_11712,N_11127,N_10599);
and U11713 (N_11713,N_10619,N_11091);
xnor U11714 (N_11714,N_10741,N_10431);
nand U11715 (N_11715,N_10859,N_11066);
xnor U11716 (N_11716,N_11019,N_10447);
nor U11717 (N_11717,N_10412,N_11103);
and U11718 (N_11718,N_10800,N_10824);
nand U11719 (N_11719,N_10957,N_10432);
or U11720 (N_11720,N_10679,N_10535);
nor U11721 (N_11721,N_10555,N_10790);
xor U11722 (N_11722,N_10600,N_10689);
nand U11723 (N_11723,N_10803,N_10879);
nor U11724 (N_11724,N_11024,N_10425);
and U11725 (N_11725,N_10897,N_11137);
nand U11726 (N_11726,N_10869,N_10680);
nand U11727 (N_11727,N_10951,N_10671);
and U11728 (N_11728,N_10615,N_10963);
and U11729 (N_11729,N_11038,N_11090);
nor U11730 (N_11730,N_10532,N_10400);
nor U11731 (N_11731,N_10587,N_10967);
nand U11732 (N_11732,N_10493,N_11041);
nor U11733 (N_11733,N_10634,N_10603);
nor U11734 (N_11734,N_10914,N_10858);
nand U11735 (N_11735,N_10798,N_10648);
nor U11736 (N_11736,N_10748,N_10728);
and U11737 (N_11737,N_10448,N_10678);
nand U11738 (N_11738,N_10527,N_10728);
xnor U11739 (N_11739,N_10926,N_11098);
and U11740 (N_11740,N_11181,N_11083);
or U11741 (N_11741,N_10730,N_10450);
and U11742 (N_11742,N_11047,N_10589);
xor U11743 (N_11743,N_10708,N_10435);
nor U11744 (N_11744,N_10493,N_10444);
nor U11745 (N_11745,N_10742,N_10549);
or U11746 (N_11746,N_10733,N_11112);
and U11747 (N_11747,N_11131,N_11167);
or U11748 (N_11748,N_10692,N_10731);
or U11749 (N_11749,N_10695,N_11113);
and U11750 (N_11750,N_10717,N_10798);
or U11751 (N_11751,N_10954,N_10531);
xor U11752 (N_11752,N_11198,N_10754);
xor U11753 (N_11753,N_11005,N_11101);
xnor U11754 (N_11754,N_10815,N_11052);
nand U11755 (N_11755,N_10794,N_10818);
xnor U11756 (N_11756,N_10942,N_10563);
nor U11757 (N_11757,N_10565,N_10804);
xnor U11758 (N_11758,N_11000,N_10433);
nand U11759 (N_11759,N_11174,N_10601);
and U11760 (N_11760,N_10669,N_10804);
xnor U11761 (N_11761,N_11080,N_10851);
xor U11762 (N_11762,N_10550,N_10563);
nor U11763 (N_11763,N_11145,N_11077);
and U11764 (N_11764,N_10849,N_10698);
nand U11765 (N_11765,N_10538,N_11073);
nand U11766 (N_11766,N_10535,N_10987);
nand U11767 (N_11767,N_10775,N_10976);
nand U11768 (N_11768,N_10913,N_10861);
or U11769 (N_11769,N_11134,N_11023);
xor U11770 (N_11770,N_10507,N_10713);
nand U11771 (N_11771,N_10892,N_10883);
nor U11772 (N_11772,N_10750,N_11170);
nand U11773 (N_11773,N_11038,N_10544);
or U11774 (N_11774,N_10651,N_10462);
nor U11775 (N_11775,N_11115,N_10487);
or U11776 (N_11776,N_11086,N_11195);
nor U11777 (N_11777,N_10538,N_10813);
nor U11778 (N_11778,N_11158,N_10781);
nand U11779 (N_11779,N_10904,N_10769);
nand U11780 (N_11780,N_11047,N_10822);
nor U11781 (N_11781,N_11144,N_10692);
xor U11782 (N_11782,N_10471,N_10441);
xnor U11783 (N_11783,N_10602,N_11104);
or U11784 (N_11784,N_10970,N_10484);
and U11785 (N_11785,N_10509,N_11040);
and U11786 (N_11786,N_10603,N_10793);
nor U11787 (N_11787,N_10564,N_10805);
or U11788 (N_11788,N_11151,N_10439);
and U11789 (N_11789,N_11193,N_10457);
and U11790 (N_11790,N_10571,N_10424);
nand U11791 (N_11791,N_10539,N_10486);
and U11792 (N_11792,N_10620,N_10664);
nor U11793 (N_11793,N_10489,N_10497);
nand U11794 (N_11794,N_11047,N_10406);
or U11795 (N_11795,N_11110,N_10427);
xor U11796 (N_11796,N_10682,N_10896);
xor U11797 (N_11797,N_10511,N_11195);
nor U11798 (N_11798,N_10782,N_10762);
nand U11799 (N_11799,N_10792,N_10928);
and U11800 (N_11800,N_10756,N_10832);
xnor U11801 (N_11801,N_10984,N_10511);
or U11802 (N_11802,N_10478,N_10702);
nand U11803 (N_11803,N_10701,N_10992);
or U11804 (N_11804,N_11142,N_10535);
or U11805 (N_11805,N_11001,N_10544);
or U11806 (N_11806,N_10917,N_10511);
or U11807 (N_11807,N_10712,N_11152);
xor U11808 (N_11808,N_11139,N_10496);
nand U11809 (N_11809,N_10992,N_10990);
xnor U11810 (N_11810,N_11079,N_10543);
nand U11811 (N_11811,N_10843,N_10470);
and U11812 (N_11812,N_11002,N_10619);
or U11813 (N_11813,N_10526,N_11146);
or U11814 (N_11814,N_10609,N_10956);
and U11815 (N_11815,N_10443,N_10475);
nand U11816 (N_11816,N_10954,N_10726);
and U11817 (N_11817,N_10400,N_10567);
or U11818 (N_11818,N_10510,N_11072);
nand U11819 (N_11819,N_11116,N_10954);
nand U11820 (N_11820,N_10816,N_11196);
nand U11821 (N_11821,N_10401,N_10552);
or U11822 (N_11822,N_10637,N_10959);
nand U11823 (N_11823,N_11031,N_10903);
xor U11824 (N_11824,N_10654,N_10809);
nand U11825 (N_11825,N_10932,N_10985);
or U11826 (N_11826,N_11179,N_11170);
nor U11827 (N_11827,N_10817,N_10934);
xnor U11828 (N_11828,N_11191,N_10640);
or U11829 (N_11829,N_10843,N_10508);
xor U11830 (N_11830,N_10688,N_10537);
and U11831 (N_11831,N_10610,N_10836);
nand U11832 (N_11832,N_11050,N_10458);
nand U11833 (N_11833,N_10443,N_10426);
xnor U11834 (N_11834,N_10905,N_11195);
nor U11835 (N_11835,N_11012,N_10604);
nor U11836 (N_11836,N_11124,N_10948);
nor U11837 (N_11837,N_10424,N_10943);
xor U11838 (N_11838,N_10576,N_10557);
nor U11839 (N_11839,N_10681,N_11179);
xor U11840 (N_11840,N_10510,N_10609);
or U11841 (N_11841,N_10828,N_10559);
nand U11842 (N_11842,N_10479,N_10413);
xor U11843 (N_11843,N_10952,N_10713);
nor U11844 (N_11844,N_10983,N_11113);
or U11845 (N_11845,N_10814,N_10963);
or U11846 (N_11846,N_11041,N_10675);
nand U11847 (N_11847,N_11165,N_11161);
nand U11848 (N_11848,N_11077,N_10951);
xnor U11849 (N_11849,N_10759,N_11174);
and U11850 (N_11850,N_10673,N_11181);
xor U11851 (N_11851,N_10961,N_11032);
or U11852 (N_11852,N_10608,N_10662);
and U11853 (N_11853,N_10977,N_11087);
or U11854 (N_11854,N_10848,N_10689);
and U11855 (N_11855,N_10721,N_10542);
and U11856 (N_11856,N_10781,N_10894);
xor U11857 (N_11857,N_10908,N_10984);
and U11858 (N_11858,N_10755,N_10832);
nor U11859 (N_11859,N_10480,N_11125);
and U11860 (N_11860,N_10471,N_10433);
nand U11861 (N_11861,N_10600,N_10726);
nor U11862 (N_11862,N_10869,N_10714);
nand U11863 (N_11863,N_10734,N_10855);
nand U11864 (N_11864,N_10986,N_10725);
nand U11865 (N_11865,N_11081,N_10569);
xor U11866 (N_11866,N_10755,N_10571);
and U11867 (N_11867,N_10636,N_11064);
nor U11868 (N_11868,N_10736,N_10562);
nand U11869 (N_11869,N_10790,N_10600);
xor U11870 (N_11870,N_10768,N_11137);
or U11871 (N_11871,N_11191,N_11120);
nand U11872 (N_11872,N_10884,N_11138);
nand U11873 (N_11873,N_10784,N_10564);
and U11874 (N_11874,N_10412,N_10611);
xnor U11875 (N_11875,N_10514,N_10931);
and U11876 (N_11876,N_10956,N_11182);
nand U11877 (N_11877,N_11004,N_10405);
nor U11878 (N_11878,N_10421,N_10435);
and U11879 (N_11879,N_11105,N_10678);
xor U11880 (N_11880,N_10639,N_11061);
xnor U11881 (N_11881,N_10660,N_11128);
nand U11882 (N_11882,N_10878,N_10725);
xor U11883 (N_11883,N_10883,N_10819);
nand U11884 (N_11884,N_11186,N_10873);
or U11885 (N_11885,N_10614,N_11102);
and U11886 (N_11886,N_11165,N_11194);
nand U11887 (N_11887,N_10644,N_10440);
nand U11888 (N_11888,N_10777,N_10552);
or U11889 (N_11889,N_11080,N_10898);
nor U11890 (N_11890,N_10542,N_11187);
or U11891 (N_11891,N_10472,N_10991);
nand U11892 (N_11892,N_10642,N_10754);
xnor U11893 (N_11893,N_10971,N_10402);
and U11894 (N_11894,N_10687,N_10485);
xnor U11895 (N_11895,N_10502,N_10497);
and U11896 (N_11896,N_11003,N_10905);
nand U11897 (N_11897,N_10965,N_10472);
or U11898 (N_11898,N_10816,N_11028);
and U11899 (N_11899,N_10416,N_11170);
nand U11900 (N_11900,N_10458,N_11195);
nand U11901 (N_11901,N_11178,N_10459);
xnor U11902 (N_11902,N_11036,N_10717);
and U11903 (N_11903,N_11064,N_10678);
xor U11904 (N_11904,N_11016,N_10511);
nor U11905 (N_11905,N_10634,N_11000);
and U11906 (N_11906,N_10771,N_10755);
xnor U11907 (N_11907,N_10641,N_11038);
and U11908 (N_11908,N_10628,N_10905);
nand U11909 (N_11909,N_10602,N_11054);
nor U11910 (N_11910,N_11016,N_10806);
xor U11911 (N_11911,N_10923,N_10675);
nor U11912 (N_11912,N_11118,N_10425);
and U11913 (N_11913,N_11124,N_10800);
nor U11914 (N_11914,N_10439,N_10728);
nor U11915 (N_11915,N_10455,N_11053);
xor U11916 (N_11916,N_10838,N_10958);
and U11917 (N_11917,N_10738,N_11150);
xor U11918 (N_11918,N_11160,N_10720);
xor U11919 (N_11919,N_10615,N_11160);
or U11920 (N_11920,N_10426,N_10975);
xor U11921 (N_11921,N_10738,N_11101);
or U11922 (N_11922,N_10461,N_10509);
xnor U11923 (N_11923,N_11130,N_10491);
nor U11924 (N_11924,N_10625,N_10819);
and U11925 (N_11925,N_10864,N_10734);
and U11926 (N_11926,N_10534,N_11174);
or U11927 (N_11927,N_10969,N_10650);
and U11928 (N_11928,N_10477,N_10408);
xor U11929 (N_11929,N_11196,N_10441);
or U11930 (N_11930,N_10412,N_10768);
nand U11931 (N_11931,N_11138,N_10448);
xnor U11932 (N_11932,N_10508,N_10942);
or U11933 (N_11933,N_10829,N_10946);
nand U11934 (N_11934,N_10959,N_10683);
and U11935 (N_11935,N_10496,N_10418);
xor U11936 (N_11936,N_10996,N_10897);
xnor U11937 (N_11937,N_10683,N_10993);
nand U11938 (N_11938,N_11124,N_10975);
nand U11939 (N_11939,N_10833,N_10792);
nor U11940 (N_11940,N_10576,N_10992);
and U11941 (N_11941,N_10743,N_10863);
nand U11942 (N_11942,N_10419,N_10777);
or U11943 (N_11943,N_10748,N_10944);
or U11944 (N_11944,N_10608,N_10587);
or U11945 (N_11945,N_11153,N_10747);
xnor U11946 (N_11946,N_10440,N_10601);
xor U11947 (N_11947,N_10808,N_10742);
xnor U11948 (N_11948,N_10995,N_10718);
xnor U11949 (N_11949,N_10702,N_11043);
xor U11950 (N_11950,N_10759,N_10555);
nor U11951 (N_11951,N_10928,N_11111);
nor U11952 (N_11952,N_10699,N_10537);
and U11953 (N_11953,N_11041,N_10907);
nand U11954 (N_11954,N_10648,N_10513);
nand U11955 (N_11955,N_10584,N_10818);
or U11956 (N_11956,N_10554,N_11080);
nor U11957 (N_11957,N_10834,N_10828);
nor U11958 (N_11958,N_10427,N_11135);
nor U11959 (N_11959,N_10937,N_10569);
nand U11960 (N_11960,N_10854,N_10858);
xor U11961 (N_11961,N_10512,N_11198);
or U11962 (N_11962,N_11042,N_10930);
nor U11963 (N_11963,N_11160,N_10518);
or U11964 (N_11964,N_10785,N_11165);
nor U11965 (N_11965,N_10455,N_10795);
and U11966 (N_11966,N_10725,N_10727);
xor U11967 (N_11967,N_10723,N_10420);
nor U11968 (N_11968,N_11027,N_10553);
xnor U11969 (N_11969,N_10866,N_10815);
and U11970 (N_11970,N_10903,N_10947);
and U11971 (N_11971,N_10638,N_11011);
xnor U11972 (N_11972,N_10494,N_10673);
nand U11973 (N_11973,N_11181,N_10889);
nand U11974 (N_11974,N_11049,N_10717);
nor U11975 (N_11975,N_11133,N_10647);
or U11976 (N_11976,N_10622,N_10923);
and U11977 (N_11977,N_10970,N_10853);
nand U11978 (N_11978,N_10863,N_10775);
xor U11979 (N_11979,N_10592,N_10524);
nor U11980 (N_11980,N_10525,N_11110);
or U11981 (N_11981,N_10634,N_10497);
and U11982 (N_11982,N_11057,N_10747);
and U11983 (N_11983,N_10627,N_10713);
or U11984 (N_11984,N_10981,N_11164);
nor U11985 (N_11985,N_10766,N_10532);
xnor U11986 (N_11986,N_10644,N_11071);
xnor U11987 (N_11987,N_10520,N_11114);
nand U11988 (N_11988,N_10830,N_11116);
or U11989 (N_11989,N_11091,N_10520);
and U11990 (N_11990,N_11134,N_10946);
and U11991 (N_11991,N_11199,N_10830);
nor U11992 (N_11992,N_10795,N_10749);
nand U11993 (N_11993,N_10834,N_10467);
xnor U11994 (N_11994,N_11088,N_10780);
and U11995 (N_11995,N_10599,N_10773);
or U11996 (N_11996,N_10700,N_10575);
and U11997 (N_11997,N_10873,N_10793);
or U11998 (N_11998,N_10605,N_11138);
or U11999 (N_11999,N_10401,N_11023);
nor U12000 (N_12000,N_11908,N_11276);
or U12001 (N_12001,N_11549,N_11900);
and U12002 (N_12002,N_11997,N_11505);
xnor U12003 (N_12003,N_11879,N_11575);
nor U12004 (N_12004,N_11256,N_11412);
nor U12005 (N_12005,N_11421,N_11802);
nand U12006 (N_12006,N_11286,N_11393);
or U12007 (N_12007,N_11752,N_11295);
nor U12008 (N_12008,N_11413,N_11605);
nand U12009 (N_12009,N_11436,N_11509);
nand U12010 (N_12010,N_11785,N_11202);
nor U12011 (N_12011,N_11811,N_11401);
or U12012 (N_12012,N_11688,N_11614);
xor U12013 (N_12013,N_11270,N_11278);
and U12014 (N_12014,N_11526,N_11717);
nand U12015 (N_12015,N_11613,N_11408);
or U12016 (N_12016,N_11260,N_11967);
or U12017 (N_12017,N_11359,N_11956);
nand U12018 (N_12018,N_11544,N_11981);
nand U12019 (N_12019,N_11827,N_11379);
or U12020 (N_12020,N_11642,N_11714);
or U12021 (N_12021,N_11620,N_11643);
and U12022 (N_12022,N_11800,N_11964);
nand U12023 (N_12023,N_11573,N_11693);
nand U12024 (N_12024,N_11859,N_11257);
and U12025 (N_12025,N_11508,N_11637);
nor U12026 (N_12026,N_11905,N_11488);
or U12027 (N_12027,N_11816,N_11340);
nor U12028 (N_12028,N_11266,N_11467);
xnor U12029 (N_12029,N_11944,N_11601);
xnor U12030 (N_12030,N_11722,N_11640);
nand U12031 (N_12031,N_11825,N_11864);
xnor U12032 (N_12032,N_11846,N_11561);
nand U12033 (N_12033,N_11796,N_11881);
and U12034 (N_12034,N_11272,N_11855);
xnor U12035 (N_12035,N_11226,N_11659);
nor U12036 (N_12036,N_11928,N_11685);
or U12037 (N_12037,N_11747,N_11756);
nor U12038 (N_12038,N_11655,N_11541);
or U12039 (N_12039,N_11400,N_11267);
or U12040 (N_12040,N_11857,N_11294);
and U12041 (N_12041,N_11686,N_11904);
or U12042 (N_12042,N_11471,N_11862);
and U12043 (N_12043,N_11410,N_11603);
xnor U12044 (N_12044,N_11580,N_11919);
nand U12045 (N_12045,N_11959,N_11521);
xor U12046 (N_12046,N_11389,N_11237);
or U12047 (N_12047,N_11607,N_11872);
nand U12048 (N_12048,N_11938,N_11470);
nor U12049 (N_12049,N_11725,N_11795);
xor U12050 (N_12050,N_11845,N_11480);
nor U12051 (N_12051,N_11560,N_11238);
and U12052 (N_12052,N_11483,N_11492);
nand U12053 (N_12053,N_11983,N_11491);
nor U12054 (N_12054,N_11709,N_11497);
nand U12055 (N_12055,N_11679,N_11995);
xor U12056 (N_12056,N_11434,N_11478);
and U12057 (N_12057,N_11984,N_11899);
nor U12058 (N_12058,N_11847,N_11622);
nor U12059 (N_12059,N_11391,N_11596);
and U12060 (N_12060,N_11883,N_11626);
nor U12061 (N_12061,N_11265,N_11874);
and U12062 (N_12062,N_11791,N_11769);
and U12063 (N_12063,N_11441,N_11748);
nand U12064 (N_12064,N_11479,N_11820);
nand U12065 (N_12065,N_11332,N_11826);
xnor U12066 (N_12066,N_11702,N_11821);
xor U12067 (N_12067,N_11435,N_11543);
nor U12068 (N_12068,N_11680,N_11388);
and U12069 (N_12069,N_11598,N_11630);
xnor U12070 (N_12070,N_11735,N_11581);
nor U12071 (N_12071,N_11366,N_11297);
or U12072 (N_12072,N_11527,N_11368);
or U12073 (N_12073,N_11418,N_11411);
or U12074 (N_12074,N_11718,N_11563);
nor U12075 (N_12075,N_11358,N_11784);
or U12076 (N_12076,N_11566,N_11739);
xor U12077 (N_12077,N_11797,N_11831);
nand U12078 (N_12078,N_11477,N_11998);
or U12079 (N_12079,N_11886,N_11455);
xor U12080 (N_12080,N_11667,N_11308);
nand U12081 (N_12081,N_11962,N_11210);
nand U12082 (N_12082,N_11442,N_11300);
or U12083 (N_12083,N_11588,N_11871);
nor U12084 (N_12084,N_11406,N_11394);
xnor U12085 (N_12085,N_11392,N_11474);
or U12086 (N_12086,N_11570,N_11382);
and U12087 (N_12087,N_11325,N_11910);
or U12088 (N_12088,N_11242,N_11447);
nor U12089 (N_12089,N_11681,N_11324);
and U12090 (N_12090,N_11292,N_11363);
nor U12091 (N_12091,N_11692,N_11909);
and U12092 (N_12092,N_11213,N_11375);
nor U12093 (N_12093,N_11774,N_11235);
and U12094 (N_12094,N_11536,N_11458);
nor U12095 (N_12095,N_11662,N_11621);
and U12096 (N_12096,N_11212,N_11933);
or U12097 (N_12097,N_11416,N_11969);
and U12098 (N_12098,N_11571,N_11429);
nand U12099 (N_12099,N_11398,N_11307);
xnor U12100 (N_12100,N_11925,N_11824);
xor U12101 (N_12101,N_11339,N_11887);
or U12102 (N_12102,N_11990,N_11283);
and U12103 (N_12103,N_11425,N_11780);
xnor U12104 (N_12104,N_11431,N_11200);
nor U12105 (N_12105,N_11243,N_11860);
xnor U12106 (N_12106,N_11931,N_11801);
nor U12107 (N_12107,N_11843,N_11830);
xor U12108 (N_12108,N_11208,N_11635);
nor U12109 (N_12109,N_11728,N_11405);
and U12110 (N_12110,N_11277,N_11893);
nor U12111 (N_12111,N_11609,N_11562);
nor U12112 (N_12112,N_11891,N_11350);
xnor U12113 (N_12113,N_11499,N_11633);
nand U12114 (N_12114,N_11745,N_11828);
nor U12115 (N_12115,N_11306,N_11889);
xnor U12116 (N_12116,N_11422,N_11616);
or U12117 (N_12117,N_11281,N_11371);
or U12118 (N_12118,N_11973,N_11740);
or U12119 (N_12119,N_11840,N_11542);
xnor U12120 (N_12120,N_11947,N_11656);
nand U12121 (N_12121,N_11654,N_11695);
or U12122 (N_12122,N_11807,N_11285);
or U12123 (N_12123,N_11729,N_11395);
and U12124 (N_12124,N_11676,N_11383);
or U12125 (N_12125,N_11316,N_11448);
nand U12126 (N_12126,N_11645,N_11290);
or U12127 (N_12127,N_11517,N_11803);
and U12128 (N_12128,N_11568,N_11914);
nand U12129 (N_12129,N_11761,N_11749);
and U12130 (N_12130,N_11450,N_11611);
or U12131 (N_12131,N_11721,N_11514);
nand U12132 (N_12132,N_11794,N_11445);
nand U12133 (N_12133,N_11439,N_11582);
nor U12134 (N_12134,N_11641,N_11484);
and U12135 (N_12135,N_11357,N_11610);
and U12136 (N_12136,N_11848,N_11913);
and U12137 (N_12137,N_11446,N_11775);
or U12138 (N_12138,N_11757,N_11917);
xnor U12139 (N_12139,N_11666,N_11958);
and U12140 (N_12140,N_11951,N_11220);
or U12141 (N_12141,N_11473,N_11806);
nor U12142 (N_12142,N_11251,N_11792);
xor U12143 (N_12143,N_11772,N_11303);
and U12144 (N_12144,N_11629,N_11804);
xnor U12145 (N_12145,N_11215,N_11895);
nand U12146 (N_12146,N_11742,N_11519);
and U12147 (N_12147,N_11952,N_11589);
xor U12148 (N_12148,N_11953,N_11945);
nand U12149 (N_12149,N_11852,N_11664);
xor U12150 (N_12150,N_11229,N_11660);
and U12151 (N_12151,N_11354,N_11593);
and U12152 (N_12152,N_11250,N_11978);
nand U12153 (N_12153,N_11254,N_11898);
xor U12154 (N_12154,N_11330,N_11515);
or U12155 (N_12155,N_11644,N_11236);
and U12156 (N_12156,N_11287,N_11551);
or U12157 (N_12157,N_11911,N_11624);
nand U12158 (N_12158,N_11485,N_11533);
xor U12159 (N_12159,N_11975,N_11451);
nor U12160 (N_12160,N_11837,N_11767);
xor U12161 (N_12161,N_11602,N_11334);
nor U12162 (N_12162,N_11433,N_11789);
or U12163 (N_12163,N_11758,N_11916);
nor U12164 (N_12164,N_11502,N_11720);
xnor U12165 (N_12165,N_11397,N_11513);
xor U12166 (N_12166,N_11832,N_11310);
nand U12167 (N_12167,N_11348,N_11489);
and U12168 (N_12168,N_11259,N_11986);
nor U12169 (N_12169,N_11738,N_11462);
xor U12170 (N_12170,N_11464,N_11960);
and U12171 (N_12171,N_11225,N_11759);
or U12172 (N_12172,N_11475,N_11961);
or U12173 (N_12173,N_11999,N_11569);
or U12174 (N_12174,N_11301,N_11396);
nor U12175 (N_12175,N_11343,N_11538);
or U12176 (N_12176,N_11487,N_11716);
and U12177 (N_12177,N_11352,N_11888);
or U12178 (N_12178,N_11691,N_11545);
or U12179 (N_12179,N_11674,N_11903);
nand U12180 (N_12180,N_11815,N_11380);
nand U12181 (N_12181,N_11902,N_11449);
xor U12182 (N_12182,N_11884,N_11506);
or U12183 (N_12183,N_11894,N_11510);
nand U12184 (N_12184,N_11833,N_11230);
and U12185 (N_12185,N_11341,N_11356);
and U12186 (N_12186,N_11374,N_11617);
and U12187 (N_12187,N_11778,N_11858);
nand U12188 (N_12188,N_11781,N_11378);
or U12189 (N_12189,N_11604,N_11298);
xnor U12190 (N_12190,N_11675,N_11579);
nand U12191 (N_12191,N_11574,N_11255);
nor U12192 (N_12192,N_11317,N_11972);
nand U12193 (N_12193,N_11284,N_11773);
xnor U12194 (N_12194,N_11639,N_11322);
nand U12195 (N_12195,N_11896,N_11223);
nor U12196 (N_12196,N_11572,N_11577);
and U12197 (N_12197,N_11424,N_11595);
nor U12198 (N_12198,N_11790,N_11980);
nor U12199 (N_12199,N_11469,N_11939);
or U12200 (N_12200,N_11700,N_11694);
or U12201 (N_12201,N_11943,N_11466);
nand U12202 (N_12202,N_11634,N_11765);
xnor U12203 (N_12203,N_11746,N_11524);
or U12204 (N_12204,N_11428,N_11460);
or U12205 (N_12205,N_11232,N_11658);
nand U12206 (N_12206,N_11623,N_11590);
or U12207 (N_12207,N_11291,N_11876);
nand U12208 (N_12208,N_11733,N_11211);
nor U12209 (N_12209,N_11377,N_11668);
nor U12210 (N_12210,N_11786,N_11732);
xor U12211 (N_12211,N_11937,N_11203);
xor U12212 (N_12212,N_11987,N_11351);
nand U12213 (N_12213,N_11776,N_11530);
nand U12214 (N_12214,N_11920,N_11892);
and U12215 (N_12215,N_11628,N_11443);
and U12216 (N_12216,N_11841,N_11856);
nor U12217 (N_12217,N_11949,N_11882);
or U12218 (N_12218,N_11402,N_11355);
nand U12219 (N_12219,N_11583,N_11534);
nand U12220 (N_12220,N_11525,N_11793);
xnor U12221 (N_12221,N_11457,N_11531);
nor U12222 (N_12222,N_11968,N_11708);
nor U12223 (N_12223,N_11690,N_11650);
xnor U12224 (N_12224,N_11565,N_11696);
nand U12225 (N_12225,N_11724,N_11713);
xor U12226 (N_12226,N_11314,N_11665);
xor U12227 (N_12227,N_11741,N_11734);
and U12228 (N_12228,N_11697,N_11880);
nor U12229 (N_12229,N_11594,N_11535);
nand U12230 (N_12230,N_11906,N_11954);
nand U12231 (N_12231,N_11218,N_11822);
or U12232 (N_12232,N_11219,N_11423);
nand U12233 (N_12233,N_11770,N_11494);
or U12234 (N_12234,N_11241,N_11730);
xnor U12235 (N_12235,N_11653,N_11842);
xor U12236 (N_12236,N_11966,N_11222);
and U12237 (N_12237,N_11438,N_11403);
xor U12238 (N_12238,N_11851,N_11651);
and U12239 (N_12239,N_11586,N_11591);
nor U12240 (N_12240,N_11768,N_11647);
or U12241 (N_12241,N_11988,N_11345);
and U12242 (N_12242,N_11263,N_11600);
xor U12243 (N_12243,N_11315,N_11963);
and U12244 (N_12244,N_11553,N_11244);
and U12245 (N_12245,N_11673,N_11247);
nand U12246 (N_12246,N_11737,N_11453);
and U12247 (N_12247,N_11548,N_11468);
nand U12248 (N_12248,N_11985,N_11540);
xor U12249 (N_12249,N_11459,N_11618);
nand U12250 (N_12250,N_11472,N_11723);
nand U12251 (N_12251,N_11865,N_11946);
nor U12252 (N_12252,N_11912,N_11979);
nand U12253 (N_12253,N_11924,N_11606);
and U12254 (N_12254,N_11989,N_11711);
nand U12255 (N_12255,N_11362,N_11427);
nand U12256 (N_12256,N_11940,N_11704);
or U12257 (N_12257,N_11373,N_11216);
or U12258 (N_12258,N_11915,N_11992);
nor U12259 (N_12259,N_11559,N_11682);
xnor U12260 (N_12260,N_11870,N_11537);
and U12261 (N_12261,N_11201,N_11547);
and U12262 (N_12262,N_11707,N_11936);
and U12263 (N_12263,N_11875,N_11361);
or U12264 (N_12264,N_11209,N_11677);
or U12265 (N_12265,N_11687,N_11764);
nor U12266 (N_12266,N_11753,N_11576);
or U12267 (N_12267,N_11783,N_11261);
and U12268 (N_12268,N_11918,N_11942);
xnor U12269 (N_12269,N_11839,N_11736);
nand U12270 (N_12270,N_11252,N_11965);
xnor U12271 (N_12271,N_11715,N_11437);
and U12272 (N_12272,N_11376,N_11342);
and U12273 (N_12273,N_11585,N_11444);
or U12274 (N_12274,N_11670,N_11763);
xnor U12275 (N_12275,N_11353,N_11663);
and U12276 (N_12276,N_11399,N_11935);
xor U12277 (N_12277,N_11550,N_11333);
and U12278 (N_12278,N_11850,N_11727);
nand U12279 (N_12279,N_11977,N_11744);
nor U12280 (N_12280,N_11901,N_11743);
and U12281 (N_12281,N_11328,N_11557);
nand U12282 (N_12282,N_11957,N_11482);
xor U12283 (N_12283,N_11710,N_11689);
and U12284 (N_12284,N_11490,N_11554);
nand U12285 (N_12285,N_11854,N_11853);
and U12286 (N_12286,N_11974,N_11275);
and U12287 (N_12287,N_11941,N_11234);
xor U12288 (N_12288,N_11930,N_11615);
and U12289 (N_12289,N_11529,N_11302);
or U12290 (N_12290,N_11246,N_11288);
xor U12291 (N_12291,N_11381,N_11866);
nand U12292 (N_12292,N_11955,N_11264);
or U12293 (N_12293,N_11347,N_11520);
nor U12294 (N_12294,N_11669,N_11982);
and U12295 (N_12295,N_11592,N_11779);
and U12296 (N_12296,N_11344,N_11671);
xnor U12297 (N_12297,N_11360,N_11861);
nor U12298 (N_12298,N_11233,N_11432);
nand U12299 (N_12299,N_11836,N_11221);
nand U12300 (N_12300,N_11309,N_11305);
nor U12301 (N_12301,N_11932,N_11672);
and U12302 (N_12302,N_11788,N_11269);
nor U12303 (N_12303,N_11817,N_11321);
nand U12304 (N_12304,N_11934,N_11948);
or U12305 (N_12305,N_11838,N_11372);
and U12306 (N_12306,N_11849,N_11552);
xnor U12307 (N_12307,N_11522,N_11558);
nor U12308 (N_12308,N_11312,N_11258);
or U12309 (N_12309,N_11227,N_11329);
or U12310 (N_12310,N_11214,N_11678);
nor U12311 (N_12311,N_11684,N_11731);
or U12312 (N_12312,N_11498,N_11703);
xnor U12313 (N_12313,N_11625,N_11699);
nand U12314 (N_12314,N_11868,N_11993);
or U12315 (N_12315,N_11504,N_11760);
nor U12316 (N_12316,N_11239,N_11555);
nand U12317 (N_12317,N_11755,N_11337);
xor U12318 (N_12318,N_11805,N_11407);
nor U12319 (N_12319,N_11349,N_11890);
and U12320 (N_12320,N_11248,N_11346);
nor U12321 (N_12321,N_11228,N_11835);
nand U12322 (N_12322,N_11863,N_11546);
and U12323 (N_12323,N_11578,N_11818);
or U12324 (N_12324,N_11313,N_11528);
xor U12325 (N_12325,N_11829,N_11486);
xnor U12326 (N_12326,N_11262,N_11701);
nand U12327 (N_12327,N_11296,N_11907);
nor U12328 (N_12328,N_11463,N_11873);
nor U12329 (N_12329,N_11496,N_11387);
and U12330 (N_12330,N_11646,N_11465);
nor U12331 (N_12331,N_11495,N_11205);
nor U12332 (N_12332,N_11409,N_11384);
xnor U12333 (N_12333,N_11299,N_11414);
nand U12334 (N_12334,N_11819,N_11319);
xnor U12335 (N_12335,N_11500,N_11231);
nand U12336 (N_12336,N_11390,N_11304);
or U12337 (N_12337,N_11619,N_11599);
nor U12338 (N_12338,N_11273,N_11782);
nor U12339 (N_12339,N_11454,N_11217);
and U12340 (N_12340,N_11501,N_11632);
nor U12341 (N_12341,N_11564,N_11608);
nand U12342 (N_12342,N_11249,N_11511);
xnor U12343 (N_12343,N_11750,N_11207);
nor U12344 (N_12344,N_11706,N_11336);
or U12345 (N_12345,N_11777,N_11523);
nor U12346 (N_12346,N_11810,N_11762);
nor U12347 (N_12347,N_11417,N_11419);
and U12348 (N_12348,N_11420,N_11950);
nor U12349 (N_12349,N_11289,N_11921);
or U12350 (N_12350,N_11507,N_11240);
nor U12351 (N_12351,N_11476,N_11869);
and U12352 (N_12352,N_11877,N_11657);
and U12353 (N_12353,N_11512,N_11456);
nor U12354 (N_12354,N_11652,N_11518);
and U12355 (N_12355,N_11369,N_11799);
nor U12356 (N_12356,N_11976,N_11293);
or U12357 (N_12357,N_11922,N_11516);
nor U12358 (N_12358,N_11338,N_11683);
xor U12359 (N_12359,N_11994,N_11282);
xnor U12360 (N_12360,N_11430,N_11970);
or U12361 (N_12361,N_11280,N_11971);
xor U12362 (N_12362,N_11636,N_11751);
nor U12363 (N_12363,N_11991,N_11204);
xor U12364 (N_12364,N_11584,N_11834);
nand U12365 (N_12365,N_11923,N_11426);
xnor U12366 (N_12366,N_11766,N_11698);
and U12367 (N_12367,N_11926,N_11493);
and U12368 (N_12368,N_11452,N_11440);
nand U12369 (N_12369,N_11814,N_11331);
nor U12370 (N_12370,N_11927,N_11808);
nand U12371 (N_12371,N_11318,N_11370);
and U12372 (N_12372,N_11224,N_11627);
xnor U12373 (N_12373,N_11996,N_11206);
xor U12374 (N_12374,N_11415,N_11567);
or U12375 (N_12375,N_11798,N_11771);
nor U12376 (N_12376,N_11335,N_11253);
nor U12377 (N_12377,N_11787,N_11885);
nand U12378 (N_12378,N_11705,N_11364);
nand U12379 (N_12379,N_11320,N_11612);
nand U12380 (N_12380,N_11268,N_11311);
or U12381 (N_12381,N_11279,N_11812);
and U12382 (N_12382,N_11327,N_11631);
xor U12383 (N_12383,N_11556,N_11481);
and U12384 (N_12384,N_11754,N_11823);
nor U12385 (N_12385,N_11404,N_11326);
nor U12386 (N_12386,N_11587,N_11649);
xnor U12387 (N_12387,N_11726,N_11878);
nand U12388 (N_12388,N_11897,N_11367);
and U12389 (N_12389,N_11597,N_11638);
and U12390 (N_12390,N_11532,N_11867);
or U12391 (N_12391,N_11929,N_11385);
or U12392 (N_12392,N_11539,N_11648);
nor U12393 (N_12393,N_11661,N_11712);
and U12394 (N_12394,N_11274,N_11809);
nand U12395 (N_12395,N_11719,N_11386);
xnor U12396 (N_12396,N_11844,N_11323);
xor U12397 (N_12397,N_11365,N_11813);
xor U12398 (N_12398,N_11503,N_11271);
nand U12399 (N_12399,N_11245,N_11461);
and U12400 (N_12400,N_11755,N_11339);
nand U12401 (N_12401,N_11504,N_11795);
nor U12402 (N_12402,N_11659,N_11873);
or U12403 (N_12403,N_11258,N_11918);
nand U12404 (N_12404,N_11339,N_11484);
xor U12405 (N_12405,N_11971,N_11316);
and U12406 (N_12406,N_11212,N_11707);
nand U12407 (N_12407,N_11345,N_11862);
or U12408 (N_12408,N_11585,N_11728);
nor U12409 (N_12409,N_11248,N_11843);
or U12410 (N_12410,N_11989,N_11829);
nor U12411 (N_12411,N_11913,N_11557);
and U12412 (N_12412,N_11426,N_11510);
nor U12413 (N_12413,N_11773,N_11738);
nand U12414 (N_12414,N_11448,N_11995);
nor U12415 (N_12415,N_11341,N_11893);
nor U12416 (N_12416,N_11689,N_11915);
nor U12417 (N_12417,N_11612,N_11651);
nor U12418 (N_12418,N_11503,N_11228);
and U12419 (N_12419,N_11661,N_11614);
xnor U12420 (N_12420,N_11581,N_11746);
or U12421 (N_12421,N_11939,N_11998);
nand U12422 (N_12422,N_11517,N_11683);
xor U12423 (N_12423,N_11820,N_11779);
nor U12424 (N_12424,N_11631,N_11846);
or U12425 (N_12425,N_11957,N_11661);
nand U12426 (N_12426,N_11255,N_11356);
nor U12427 (N_12427,N_11398,N_11994);
or U12428 (N_12428,N_11932,N_11960);
nor U12429 (N_12429,N_11869,N_11975);
or U12430 (N_12430,N_11697,N_11292);
or U12431 (N_12431,N_11950,N_11364);
xor U12432 (N_12432,N_11224,N_11378);
nor U12433 (N_12433,N_11212,N_11291);
nand U12434 (N_12434,N_11768,N_11667);
and U12435 (N_12435,N_11916,N_11991);
xnor U12436 (N_12436,N_11770,N_11209);
or U12437 (N_12437,N_11317,N_11523);
and U12438 (N_12438,N_11402,N_11365);
and U12439 (N_12439,N_11983,N_11667);
or U12440 (N_12440,N_11889,N_11808);
or U12441 (N_12441,N_11623,N_11912);
or U12442 (N_12442,N_11325,N_11883);
nand U12443 (N_12443,N_11661,N_11600);
xor U12444 (N_12444,N_11618,N_11366);
nor U12445 (N_12445,N_11858,N_11686);
nand U12446 (N_12446,N_11632,N_11465);
xor U12447 (N_12447,N_11609,N_11947);
xnor U12448 (N_12448,N_11920,N_11450);
and U12449 (N_12449,N_11356,N_11737);
nand U12450 (N_12450,N_11274,N_11611);
nor U12451 (N_12451,N_11905,N_11463);
xnor U12452 (N_12452,N_11802,N_11569);
xnor U12453 (N_12453,N_11775,N_11627);
nand U12454 (N_12454,N_11323,N_11640);
and U12455 (N_12455,N_11458,N_11254);
xnor U12456 (N_12456,N_11363,N_11656);
or U12457 (N_12457,N_11577,N_11318);
nand U12458 (N_12458,N_11855,N_11991);
nor U12459 (N_12459,N_11759,N_11824);
xor U12460 (N_12460,N_11701,N_11734);
nor U12461 (N_12461,N_11337,N_11499);
or U12462 (N_12462,N_11939,N_11286);
and U12463 (N_12463,N_11494,N_11857);
nor U12464 (N_12464,N_11664,N_11372);
nand U12465 (N_12465,N_11655,N_11751);
or U12466 (N_12466,N_11247,N_11451);
xor U12467 (N_12467,N_11858,N_11715);
and U12468 (N_12468,N_11959,N_11704);
nand U12469 (N_12469,N_11260,N_11264);
or U12470 (N_12470,N_11998,N_11524);
or U12471 (N_12471,N_11445,N_11902);
xnor U12472 (N_12472,N_11755,N_11615);
or U12473 (N_12473,N_11238,N_11995);
nand U12474 (N_12474,N_11748,N_11688);
or U12475 (N_12475,N_11466,N_11307);
nor U12476 (N_12476,N_11207,N_11885);
xor U12477 (N_12477,N_11604,N_11671);
and U12478 (N_12478,N_11724,N_11312);
xor U12479 (N_12479,N_11272,N_11767);
nand U12480 (N_12480,N_11777,N_11236);
xor U12481 (N_12481,N_11417,N_11475);
and U12482 (N_12482,N_11431,N_11971);
nor U12483 (N_12483,N_11700,N_11762);
nor U12484 (N_12484,N_11843,N_11478);
and U12485 (N_12485,N_11379,N_11605);
nor U12486 (N_12486,N_11308,N_11573);
or U12487 (N_12487,N_11295,N_11671);
xnor U12488 (N_12488,N_11318,N_11904);
nand U12489 (N_12489,N_11977,N_11612);
xor U12490 (N_12490,N_11311,N_11329);
nand U12491 (N_12491,N_11822,N_11414);
nor U12492 (N_12492,N_11951,N_11673);
xnor U12493 (N_12493,N_11495,N_11488);
xor U12494 (N_12494,N_11407,N_11868);
nor U12495 (N_12495,N_11581,N_11227);
or U12496 (N_12496,N_11723,N_11877);
and U12497 (N_12497,N_11365,N_11403);
or U12498 (N_12498,N_11971,N_11985);
nor U12499 (N_12499,N_11802,N_11561);
nand U12500 (N_12500,N_11873,N_11497);
and U12501 (N_12501,N_11599,N_11302);
and U12502 (N_12502,N_11975,N_11947);
nor U12503 (N_12503,N_11213,N_11843);
nand U12504 (N_12504,N_11862,N_11966);
xnor U12505 (N_12505,N_11445,N_11857);
xnor U12506 (N_12506,N_11607,N_11666);
and U12507 (N_12507,N_11596,N_11260);
nor U12508 (N_12508,N_11744,N_11285);
xor U12509 (N_12509,N_11784,N_11930);
nor U12510 (N_12510,N_11766,N_11996);
xor U12511 (N_12511,N_11964,N_11726);
and U12512 (N_12512,N_11952,N_11370);
nand U12513 (N_12513,N_11746,N_11815);
xor U12514 (N_12514,N_11819,N_11761);
and U12515 (N_12515,N_11232,N_11804);
nor U12516 (N_12516,N_11916,N_11242);
or U12517 (N_12517,N_11836,N_11999);
and U12518 (N_12518,N_11748,N_11557);
nand U12519 (N_12519,N_11906,N_11401);
nand U12520 (N_12520,N_11264,N_11913);
and U12521 (N_12521,N_11314,N_11307);
and U12522 (N_12522,N_11637,N_11829);
nand U12523 (N_12523,N_11668,N_11595);
xor U12524 (N_12524,N_11334,N_11990);
or U12525 (N_12525,N_11290,N_11322);
and U12526 (N_12526,N_11795,N_11261);
nand U12527 (N_12527,N_11968,N_11645);
or U12528 (N_12528,N_11793,N_11937);
or U12529 (N_12529,N_11685,N_11609);
nand U12530 (N_12530,N_11373,N_11506);
or U12531 (N_12531,N_11905,N_11960);
or U12532 (N_12532,N_11795,N_11605);
nand U12533 (N_12533,N_11949,N_11970);
nand U12534 (N_12534,N_11414,N_11841);
nor U12535 (N_12535,N_11544,N_11427);
or U12536 (N_12536,N_11520,N_11462);
nand U12537 (N_12537,N_11261,N_11361);
nand U12538 (N_12538,N_11747,N_11276);
nand U12539 (N_12539,N_11636,N_11840);
nand U12540 (N_12540,N_11480,N_11284);
or U12541 (N_12541,N_11923,N_11203);
and U12542 (N_12542,N_11460,N_11235);
or U12543 (N_12543,N_11524,N_11499);
xnor U12544 (N_12544,N_11826,N_11981);
or U12545 (N_12545,N_11521,N_11639);
nand U12546 (N_12546,N_11645,N_11361);
nor U12547 (N_12547,N_11917,N_11554);
xnor U12548 (N_12548,N_11529,N_11879);
and U12549 (N_12549,N_11521,N_11614);
nor U12550 (N_12550,N_11351,N_11350);
nand U12551 (N_12551,N_11777,N_11673);
or U12552 (N_12552,N_11828,N_11537);
xor U12553 (N_12553,N_11657,N_11557);
or U12554 (N_12554,N_11828,N_11564);
nand U12555 (N_12555,N_11637,N_11272);
and U12556 (N_12556,N_11944,N_11629);
xnor U12557 (N_12557,N_11238,N_11242);
nor U12558 (N_12558,N_11233,N_11838);
nand U12559 (N_12559,N_11975,N_11659);
nor U12560 (N_12560,N_11940,N_11708);
xor U12561 (N_12561,N_11229,N_11907);
or U12562 (N_12562,N_11920,N_11788);
nor U12563 (N_12563,N_11203,N_11384);
and U12564 (N_12564,N_11852,N_11971);
nor U12565 (N_12565,N_11218,N_11664);
nand U12566 (N_12566,N_11467,N_11483);
and U12567 (N_12567,N_11610,N_11557);
nand U12568 (N_12568,N_11514,N_11758);
or U12569 (N_12569,N_11784,N_11677);
nand U12570 (N_12570,N_11295,N_11247);
and U12571 (N_12571,N_11998,N_11856);
or U12572 (N_12572,N_11905,N_11264);
nor U12573 (N_12573,N_11278,N_11352);
or U12574 (N_12574,N_11393,N_11490);
xnor U12575 (N_12575,N_11950,N_11645);
nor U12576 (N_12576,N_11671,N_11312);
xnor U12577 (N_12577,N_11228,N_11206);
nor U12578 (N_12578,N_11436,N_11611);
xor U12579 (N_12579,N_11629,N_11555);
and U12580 (N_12580,N_11939,N_11523);
xor U12581 (N_12581,N_11794,N_11307);
or U12582 (N_12582,N_11354,N_11255);
or U12583 (N_12583,N_11275,N_11273);
nand U12584 (N_12584,N_11574,N_11865);
and U12585 (N_12585,N_11510,N_11302);
nand U12586 (N_12586,N_11332,N_11447);
and U12587 (N_12587,N_11939,N_11501);
and U12588 (N_12588,N_11667,N_11921);
and U12589 (N_12589,N_11912,N_11659);
or U12590 (N_12590,N_11852,N_11355);
nand U12591 (N_12591,N_11447,N_11466);
nand U12592 (N_12592,N_11702,N_11662);
and U12593 (N_12593,N_11839,N_11598);
nor U12594 (N_12594,N_11642,N_11639);
xor U12595 (N_12595,N_11242,N_11841);
nand U12596 (N_12596,N_11935,N_11869);
nand U12597 (N_12597,N_11749,N_11215);
nor U12598 (N_12598,N_11743,N_11997);
nand U12599 (N_12599,N_11426,N_11712);
xnor U12600 (N_12600,N_11670,N_11405);
or U12601 (N_12601,N_11395,N_11932);
xor U12602 (N_12602,N_11877,N_11346);
xnor U12603 (N_12603,N_11861,N_11791);
and U12604 (N_12604,N_11329,N_11206);
nor U12605 (N_12605,N_11279,N_11980);
nor U12606 (N_12606,N_11543,N_11672);
xnor U12607 (N_12607,N_11203,N_11202);
xor U12608 (N_12608,N_11243,N_11688);
and U12609 (N_12609,N_11472,N_11464);
xnor U12610 (N_12610,N_11951,N_11429);
nor U12611 (N_12611,N_11927,N_11343);
and U12612 (N_12612,N_11655,N_11464);
nand U12613 (N_12613,N_11442,N_11513);
nor U12614 (N_12614,N_11888,N_11724);
and U12615 (N_12615,N_11281,N_11393);
nand U12616 (N_12616,N_11552,N_11447);
and U12617 (N_12617,N_11901,N_11281);
or U12618 (N_12618,N_11674,N_11515);
xor U12619 (N_12619,N_11614,N_11440);
nand U12620 (N_12620,N_11936,N_11376);
and U12621 (N_12621,N_11803,N_11729);
nand U12622 (N_12622,N_11418,N_11387);
xor U12623 (N_12623,N_11999,N_11949);
nand U12624 (N_12624,N_11758,N_11413);
nand U12625 (N_12625,N_11350,N_11641);
nand U12626 (N_12626,N_11891,N_11444);
and U12627 (N_12627,N_11602,N_11829);
xnor U12628 (N_12628,N_11381,N_11476);
and U12629 (N_12629,N_11759,N_11522);
nand U12630 (N_12630,N_11265,N_11370);
and U12631 (N_12631,N_11757,N_11954);
or U12632 (N_12632,N_11735,N_11914);
nand U12633 (N_12633,N_11839,N_11307);
nor U12634 (N_12634,N_11428,N_11565);
or U12635 (N_12635,N_11938,N_11478);
xor U12636 (N_12636,N_11570,N_11645);
or U12637 (N_12637,N_11614,N_11645);
nor U12638 (N_12638,N_11424,N_11407);
and U12639 (N_12639,N_11965,N_11469);
nand U12640 (N_12640,N_11259,N_11239);
and U12641 (N_12641,N_11838,N_11562);
nand U12642 (N_12642,N_11414,N_11877);
and U12643 (N_12643,N_11619,N_11271);
or U12644 (N_12644,N_11572,N_11753);
nand U12645 (N_12645,N_11957,N_11963);
nor U12646 (N_12646,N_11282,N_11276);
and U12647 (N_12647,N_11672,N_11306);
nor U12648 (N_12648,N_11553,N_11918);
xnor U12649 (N_12649,N_11855,N_11582);
and U12650 (N_12650,N_11669,N_11941);
or U12651 (N_12651,N_11516,N_11409);
nand U12652 (N_12652,N_11963,N_11830);
nand U12653 (N_12653,N_11966,N_11555);
xor U12654 (N_12654,N_11959,N_11349);
or U12655 (N_12655,N_11631,N_11234);
nor U12656 (N_12656,N_11964,N_11351);
nand U12657 (N_12657,N_11550,N_11590);
nand U12658 (N_12658,N_11529,N_11955);
and U12659 (N_12659,N_11980,N_11687);
nor U12660 (N_12660,N_11432,N_11414);
xor U12661 (N_12661,N_11247,N_11205);
or U12662 (N_12662,N_11808,N_11743);
or U12663 (N_12663,N_11613,N_11396);
and U12664 (N_12664,N_11206,N_11620);
nor U12665 (N_12665,N_11943,N_11944);
nand U12666 (N_12666,N_11637,N_11484);
nand U12667 (N_12667,N_11652,N_11448);
nor U12668 (N_12668,N_11246,N_11271);
xor U12669 (N_12669,N_11670,N_11790);
and U12670 (N_12670,N_11915,N_11876);
and U12671 (N_12671,N_11290,N_11348);
xor U12672 (N_12672,N_11524,N_11450);
nand U12673 (N_12673,N_11584,N_11462);
xnor U12674 (N_12674,N_11357,N_11849);
and U12675 (N_12675,N_11441,N_11558);
and U12676 (N_12676,N_11324,N_11964);
and U12677 (N_12677,N_11274,N_11393);
and U12678 (N_12678,N_11757,N_11974);
or U12679 (N_12679,N_11694,N_11504);
xor U12680 (N_12680,N_11348,N_11543);
and U12681 (N_12681,N_11214,N_11414);
nor U12682 (N_12682,N_11565,N_11582);
xor U12683 (N_12683,N_11425,N_11778);
nand U12684 (N_12684,N_11723,N_11609);
xor U12685 (N_12685,N_11886,N_11387);
xor U12686 (N_12686,N_11241,N_11823);
or U12687 (N_12687,N_11976,N_11376);
nand U12688 (N_12688,N_11872,N_11579);
nor U12689 (N_12689,N_11392,N_11707);
nor U12690 (N_12690,N_11332,N_11693);
nor U12691 (N_12691,N_11883,N_11254);
and U12692 (N_12692,N_11380,N_11673);
or U12693 (N_12693,N_11798,N_11379);
and U12694 (N_12694,N_11609,N_11616);
or U12695 (N_12695,N_11334,N_11253);
nand U12696 (N_12696,N_11763,N_11642);
nand U12697 (N_12697,N_11935,N_11393);
and U12698 (N_12698,N_11883,N_11390);
xnor U12699 (N_12699,N_11743,N_11235);
or U12700 (N_12700,N_11928,N_11682);
nor U12701 (N_12701,N_11266,N_11473);
xnor U12702 (N_12702,N_11421,N_11241);
nand U12703 (N_12703,N_11469,N_11214);
or U12704 (N_12704,N_11203,N_11896);
or U12705 (N_12705,N_11539,N_11759);
nor U12706 (N_12706,N_11701,N_11255);
nor U12707 (N_12707,N_11330,N_11867);
nor U12708 (N_12708,N_11444,N_11201);
xor U12709 (N_12709,N_11848,N_11329);
xnor U12710 (N_12710,N_11685,N_11218);
or U12711 (N_12711,N_11683,N_11668);
and U12712 (N_12712,N_11964,N_11308);
nor U12713 (N_12713,N_11726,N_11217);
and U12714 (N_12714,N_11551,N_11665);
nor U12715 (N_12715,N_11390,N_11614);
nor U12716 (N_12716,N_11349,N_11204);
and U12717 (N_12717,N_11875,N_11257);
xnor U12718 (N_12718,N_11440,N_11604);
nor U12719 (N_12719,N_11581,N_11646);
or U12720 (N_12720,N_11656,N_11853);
xnor U12721 (N_12721,N_11558,N_11824);
nor U12722 (N_12722,N_11907,N_11969);
and U12723 (N_12723,N_11368,N_11662);
or U12724 (N_12724,N_11555,N_11978);
and U12725 (N_12725,N_11487,N_11516);
or U12726 (N_12726,N_11653,N_11984);
nor U12727 (N_12727,N_11456,N_11464);
nor U12728 (N_12728,N_11717,N_11586);
or U12729 (N_12729,N_11617,N_11857);
nand U12730 (N_12730,N_11261,N_11594);
nand U12731 (N_12731,N_11507,N_11569);
xnor U12732 (N_12732,N_11789,N_11667);
or U12733 (N_12733,N_11887,N_11929);
and U12734 (N_12734,N_11354,N_11333);
or U12735 (N_12735,N_11731,N_11911);
xor U12736 (N_12736,N_11814,N_11592);
nand U12737 (N_12737,N_11818,N_11229);
xnor U12738 (N_12738,N_11843,N_11907);
nand U12739 (N_12739,N_11856,N_11433);
xnor U12740 (N_12740,N_11282,N_11583);
nor U12741 (N_12741,N_11566,N_11884);
xnor U12742 (N_12742,N_11491,N_11235);
nor U12743 (N_12743,N_11860,N_11983);
nor U12744 (N_12744,N_11908,N_11213);
xnor U12745 (N_12745,N_11805,N_11566);
nand U12746 (N_12746,N_11829,N_11943);
nor U12747 (N_12747,N_11565,N_11882);
nor U12748 (N_12748,N_11957,N_11331);
or U12749 (N_12749,N_11797,N_11524);
xnor U12750 (N_12750,N_11584,N_11695);
nand U12751 (N_12751,N_11745,N_11964);
nor U12752 (N_12752,N_11914,N_11345);
and U12753 (N_12753,N_11777,N_11556);
nor U12754 (N_12754,N_11848,N_11412);
xnor U12755 (N_12755,N_11715,N_11239);
nand U12756 (N_12756,N_11878,N_11299);
and U12757 (N_12757,N_11525,N_11442);
nor U12758 (N_12758,N_11473,N_11213);
xnor U12759 (N_12759,N_11723,N_11775);
or U12760 (N_12760,N_11332,N_11948);
nor U12761 (N_12761,N_11391,N_11326);
nand U12762 (N_12762,N_11224,N_11578);
and U12763 (N_12763,N_11211,N_11726);
nor U12764 (N_12764,N_11933,N_11222);
and U12765 (N_12765,N_11383,N_11601);
or U12766 (N_12766,N_11267,N_11662);
xnor U12767 (N_12767,N_11594,N_11322);
nor U12768 (N_12768,N_11941,N_11287);
nor U12769 (N_12769,N_11302,N_11260);
nor U12770 (N_12770,N_11697,N_11492);
xor U12771 (N_12771,N_11808,N_11318);
or U12772 (N_12772,N_11588,N_11667);
nor U12773 (N_12773,N_11666,N_11649);
nand U12774 (N_12774,N_11666,N_11678);
xor U12775 (N_12775,N_11572,N_11765);
xor U12776 (N_12776,N_11637,N_11397);
or U12777 (N_12777,N_11299,N_11424);
xor U12778 (N_12778,N_11767,N_11627);
nor U12779 (N_12779,N_11837,N_11329);
or U12780 (N_12780,N_11657,N_11819);
or U12781 (N_12781,N_11889,N_11720);
xnor U12782 (N_12782,N_11341,N_11677);
or U12783 (N_12783,N_11523,N_11759);
xor U12784 (N_12784,N_11953,N_11234);
or U12785 (N_12785,N_11890,N_11955);
nor U12786 (N_12786,N_11445,N_11996);
and U12787 (N_12787,N_11779,N_11955);
nor U12788 (N_12788,N_11637,N_11387);
nand U12789 (N_12789,N_11985,N_11528);
or U12790 (N_12790,N_11426,N_11689);
nor U12791 (N_12791,N_11475,N_11521);
and U12792 (N_12792,N_11633,N_11495);
nand U12793 (N_12793,N_11688,N_11799);
xnor U12794 (N_12794,N_11336,N_11833);
xnor U12795 (N_12795,N_11851,N_11960);
nor U12796 (N_12796,N_11365,N_11594);
nand U12797 (N_12797,N_11512,N_11817);
and U12798 (N_12798,N_11647,N_11425);
and U12799 (N_12799,N_11535,N_11475);
xnor U12800 (N_12800,N_12257,N_12155);
xnor U12801 (N_12801,N_12528,N_12048);
nand U12802 (N_12802,N_12077,N_12093);
and U12803 (N_12803,N_12704,N_12401);
nor U12804 (N_12804,N_12335,N_12381);
and U12805 (N_12805,N_12172,N_12341);
or U12806 (N_12806,N_12793,N_12151);
and U12807 (N_12807,N_12089,N_12109);
nand U12808 (N_12808,N_12445,N_12512);
xor U12809 (N_12809,N_12452,N_12671);
or U12810 (N_12810,N_12090,N_12281);
nor U12811 (N_12811,N_12137,N_12477);
and U12812 (N_12812,N_12010,N_12513);
nor U12813 (N_12813,N_12763,N_12150);
and U12814 (N_12814,N_12292,N_12453);
nand U12815 (N_12815,N_12365,N_12400);
nor U12816 (N_12816,N_12421,N_12687);
and U12817 (N_12817,N_12777,N_12626);
nor U12818 (N_12818,N_12439,N_12361);
nor U12819 (N_12819,N_12773,N_12118);
nor U12820 (N_12820,N_12429,N_12614);
nand U12821 (N_12821,N_12588,N_12627);
xnor U12822 (N_12822,N_12099,N_12273);
nand U12823 (N_12823,N_12555,N_12568);
and U12824 (N_12824,N_12009,N_12480);
xor U12825 (N_12825,N_12698,N_12725);
nor U12826 (N_12826,N_12611,N_12218);
nor U12827 (N_12827,N_12536,N_12530);
or U12828 (N_12828,N_12641,N_12045);
xor U12829 (N_12829,N_12438,N_12746);
xnor U12830 (N_12830,N_12500,N_12427);
nand U12831 (N_12831,N_12117,N_12116);
and U12832 (N_12832,N_12322,N_12410);
nand U12833 (N_12833,N_12367,N_12022);
xnor U12834 (N_12834,N_12720,N_12070);
xnor U12835 (N_12835,N_12209,N_12402);
and U12836 (N_12836,N_12545,N_12379);
nand U12837 (N_12837,N_12355,N_12663);
xnor U12838 (N_12838,N_12289,N_12646);
nand U12839 (N_12839,N_12463,N_12315);
xnor U12840 (N_12840,N_12509,N_12543);
nor U12841 (N_12841,N_12111,N_12354);
xor U12842 (N_12842,N_12208,N_12694);
nor U12843 (N_12843,N_12318,N_12211);
or U12844 (N_12844,N_12526,N_12046);
and U12845 (N_12845,N_12443,N_12572);
nand U12846 (N_12846,N_12397,N_12144);
and U12847 (N_12847,N_12140,N_12073);
xor U12848 (N_12848,N_12252,N_12675);
xor U12849 (N_12849,N_12722,N_12470);
or U12850 (N_12850,N_12221,N_12479);
and U12851 (N_12851,N_12344,N_12206);
or U12852 (N_12852,N_12595,N_12409);
or U12853 (N_12853,N_12290,N_12524);
nor U12854 (N_12854,N_12241,N_12043);
nand U12855 (N_12855,N_12059,N_12128);
nor U12856 (N_12856,N_12630,N_12785);
xor U12857 (N_12857,N_12624,N_12781);
xor U12858 (N_12858,N_12200,N_12605);
xnor U12859 (N_12859,N_12504,N_12661);
xnor U12860 (N_12860,N_12072,N_12245);
nand U12861 (N_12861,N_12134,N_12210);
or U12862 (N_12862,N_12343,N_12550);
or U12863 (N_12863,N_12305,N_12436);
nor U12864 (N_12864,N_12237,N_12228);
nor U12865 (N_12865,N_12013,N_12780);
nor U12866 (N_12866,N_12069,N_12057);
nor U12867 (N_12867,N_12593,N_12225);
and U12868 (N_12868,N_12390,N_12712);
nand U12869 (N_12869,N_12638,N_12597);
nand U12870 (N_12870,N_12475,N_12520);
and U12871 (N_12871,N_12581,N_12407);
or U12872 (N_12872,N_12681,N_12548);
nand U12873 (N_12873,N_12388,N_12363);
nor U12874 (N_12874,N_12166,N_12564);
nor U12875 (N_12875,N_12551,N_12458);
and U12876 (N_12876,N_12522,N_12266);
nand U12877 (N_12877,N_12177,N_12146);
or U12878 (N_12878,N_12008,N_12123);
nand U12879 (N_12879,N_12589,N_12461);
or U12880 (N_12880,N_12263,N_12411);
nor U12881 (N_12881,N_12766,N_12213);
and U12882 (N_12882,N_12613,N_12747);
nor U12883 (N_12883,N_12690,N_12672);
nor U12884 (N_12884,N_12575,N_12538);
and U12885 (N_12885,N_12478,N_12387);
nand U12886 (N_12886,N_12404,N_12507);
nand U12887 (N_12887,N_12311,N_12269);
nand U12888 (N_12888,N_12102,N_12629);
nand U12889 (N_12889,N_12255,N_12792);
xor U12890 (N_12890,N_12312,N_12492);
nand U12891 (N_12891,N_12599,N_12424);
nor U12892 (N_12892,N_12718,N_12721);
and U12893 (N_12893,N_12101,N_12351);
or U12894 (N_12894,N_12087,N_12679);
xor U12895 (N_12895,N_12639,N_12382);
nor U12896 (N_12896,N_12161,N_12352);
or U12897 (N_12897,N_12247,N_12431);
and U12898 (N_12898,N_12533,N_12015);
or U12899 (N_12899,N_12251,N_12384);
nor U12900 (N_12900,N_12062,N_12360);
nor U12901 (N_12901,N_12496,N_12441);
or U12902 (N_12902,N_12164,N_12339);
or U12903 (N_12903,N_12095,N_12167);
nor U12904 (N_12904,N_12112,N_12029);
nand U12905 (N_12905,N_12065,N_12449);
nand U12906 (N_12906,N_12236,N_12193);
xnor U12907 (N_12907,N_12414,N_12081);
xor U12908 (N_12908,N_12017,N_12303);
and U12909 (N_12909,N_12521,N_12770);
nor U12910 (N_12910,N_12573,N_12465);
nor U12911 (N_12911,N_12234,N_12444);
nand U12912 (N_12912,N_12306,N_12708);
nor U12913 (N_12913,N_12272,N_12580);
xnor U12914 (N_12914,N_12403,N_12563);
or U12915 (N_12915,N_12511,N_12506);
nand U12916 (N_12916,N_12019,N_12216);
nand U12917 (N_12917,N_12784,N_12645);
and U12918 (N_12918,N_12552,N_12497);
and U12919 (N_12919,N_12764,N_12032);
and U12920 (N_12920,N_12499,N_12615);
and U12921 (N_12921,N_12488,N_12745);
or U12922 (N_12922,N_12217,N_12625);
xnor U12923 (N_12923,N_12709,N_12620);
nor U12924 (N_12924,N_12654,N_12783);
xnor U12925 (N_12925,N_12232,N_12136);
or U12926 (N_12926,N_12034,N_12767);
xnor U12927 (N_12927,N_12796,N_12347);
xor U12928 (N_12928,N_12106,N_12456);
xor U12929 (N_12929,N_12602,N_12420);
nand U12930 (N_12930,N_12024,N_12201);
or U12931 (N_12931,N_12787,N_12519);
nand U12932 (N_12932,N_12130,N_12316);
xnor U12933 (N_12933,N_12394,N_12143);
xnor U12934 (N_12934,N_12612,N_12560);
xor U12935 (N_12935,N_12481,N_12359);
xnor U12936 (N_12936,N_12190,N_12121);
or U12937 (N_12937,N_12031,N_12353);
nor U12938 (N_12938,N_12650,N_12229);
or U12939 (N_12939,N_12212,N_12570);
and U12940 (N_12940,N_12425,N_12776);
xnor U12941 (N_12941,N_12584,N_12622);
xnor U12942 (N_12942,N_12219,N_12765);
nor U12943 (N_12943,N_12254,N_12689);
nor U12944 (N_12944,N_12670,N_12544);
and U12945 (N_12945,N_12691,N_12494);
and U12946 (N_12946,N_12020,N_12405);
nor U12947 (N_12947,N_12744,N_12755);
or U12948 (N_12948,N_12398,N_12334);
or U12949 (N_12949,N_12797,N_12537);
or U12950 (N_12950,N_12790,N_12280);
nor U12951 (N_12951,N_12297,N_12231);
nand U12952 (N_12952,N_12191,N_12386);
or U12953 (N_12953,N_12185,N_12084);
xnor U12954 (N_12954,N_12711,N_12261);
and U12955 (N_12955,N_12418,N_12758);
nor U12956 (N_12956,N_12642,N_12768);
nor U12957 (N_12957,N_12320,N_12267);
and U12958 (N_12958,N_12139,N_12393);
xnor U12959 (N_12959,N_12082,N_12759);
nor U12960 (N_12960,N_12737,N_12184);
nand U12961 (N_12961,N_12732,N_12001);
xnor U12962 (N_12962,N_12056,N_12702);
or U12963 (N_12963,N_12727,N_12050);
nor U12964 (N_12964,N_12396,N_12486);
and U12965 (N_12965,N_12331,N_12577);
or U12966 (N_12966,N_12743,N_12433);
nand U12967 (N_12967,N_12742,N_12607);
and U12968 (N_12968,N_12508,N_12233);
nand U12969 (N_12969,N_12214,N_12035);
or U12970 (N_12970,N_12124,N_12250);
nand U12971 (N_12971,N_12340,N_12462);
and U12972 (N_12972,N_12493,N_12422);
xnor U12973 (N_12973,N_12142,N_12149);
and U12974 (N_12974,N_12535,N_12215);
nand U12975 (N_12975,N_12058,N_12284);
and U12976 (N_12976,N_12385,N_12364);
nor U12977 (N_12977,N_12205,N_12557);
xor U12978 (N_12978,N_12176,N_12476);
xor U12979 (N_12979,N_12002,N_12358);
nor U12980 (N_12980,N_12468,N_12419);
nor U12981 (N_12981,N_12634,N_12715);
nand U12982 (N_12982,N_12180,N_12567);
nor U12983 (N_12983,N_12415,N_12086);
nand U12984 (N_12984,N_12561,N_12196);
nand U12985 (N_12985,N_12649,N_12483);
nor U12986 (N_12986,N_12517,N_12304);
xor U12987 (N_12987,N_12288,N_12258);
and U12988 (N_12988,N_12502,N_12094);
nand U12989 (N_12989,N_12591,N_12348);
or U12990 (N_12990,N_12484,N_12673);
xnor U12991 (N_12991,N_12556,N_12651);
nor U12992 (N_12992,N_12350,N_12697);
nor U12993 (N_12993,N_12063,N_12126);
xor U12994 (N_12994,N_12736,N_12706);
nor U12995 (N_12995,N_12616,N_12194);
and U12996 (N_12996,N_12110,N_12738);
or U12997 (N_12997,N_12623,N_12440);
or U12998 (N_12998,N_12734,N_12383);
or U12999 (N_12999,N_12757,N_12088);
nor U13000 (N_13000,N_12637,N_12587);
xor U13001 (N_13001,N_12230,N_12378);
nand U13002 (N_13002,N_12631,N_12222);
nand U13003 (N_13003,N_12523,N_12170);
nor U13004 (N_13004,N_12064,N_12047);
and U13005 (N_13005,N_12539,N_12558);
nor U13006 (N_13006,N_12075,N_12033);
nor U13007 (N_13007,N_12447,N_12515);
and U13008 (N_13008,N_12085,N_12761);
and U13009 (N_13009,N_12603,N_12157);
nor U13010 (N_13010,N_12152,N_12158);
or U13011 (N_13011,N_12505,N_12677);
and U13012 (N_13012,N_12684,N_12310);
or U13013 (N_13013,N_12338,N_12685);
or U13014 (N_13014,N_12138,N_12547);
and U13015 (N_13015,N_12324,N_12699);
xnor U13016 (N_13016,N_12171,N_12710);
nor U13017 (N_13017,N_12371,N_12326);
xor U13018 (N_13018,N_12666,N_12719);
or U13019 (N_13019,N_12774,N_12187);
nand U13020 (N_13020,N_12100,N_12644);
or U13021 (N_13021,N_12264,N_12789);
nand U13022 (N_13022,N_12606,N_12569);
and U13023 (N_13023,N_12571,N_12313);
nor U13024 (N_13024,N_12283,N_12183);
nor U13025 (N_13025,N_12204,N_12103);
nor U13026 (N_13026,N_12771,N_12643);
xor U13027 (N_13027,N_12399,N_12660);
nor U13028 (N_13028,N_12270,N_12598);
xor U13029 (N_13029,N_12299,N_12105);
nor U13030 (N_13030,N_12052,N_12346);
or U13031 (N_13031,N_12068,N_12518);
nand U13032 (N_13032,N_12071,N_12053);
nand U13033 (N_13033,N_12559,N_12540);
nand U13034 (N_13034,N_12246,N_12042);
and U13035 (N_13035,N_12782,N_12582);
nor U13036 (N_13036,N_12798,N_12795);
nor U13037 (N_13037,N_12125,N_12662);
nor U13038 (N_13038,N_12275,N_12485);
nor U13039 (N_13039,N_12647,N_12027);
and U13040 (N_13040,N_12092,N_12119);
and U13041 (N_13041,N_12426,N_12448);
xnor U13042 (N_13042,N_12145,N_12374);
xor U13043 (N_13043,N_12114,N_12491);
or U13044 (N_13044,N_12362,N_12735);
nand U13045 (N_13045,N_12450,N_12680);
nor U13046 (N_13046,N_12472,N_12207);
xnor U13047 (N_13047,N_12389,N_12132);
nor U13048 (N_13048,N_12610,N_12242);
xor U13049 (N_13049,N_12621,N_12701);
nand U13050 (N_13050,N_12750,N_12489);
and U13051 (N_13051,N_12395,N_12669);
or U13052 (N_13052,N_12298,N_12633);
nor U13053 (N_13053,N_12163,N_12778);
xor U13054 (N_13054,N_12514,N_12244);
or U13055 (N_13055,N_12030,N_12655);
or U13056 (N_13056,N_12113,N_12723);
nor U13057 (N_13057,N_12159,N_12023);
or U13058 (N_13058,N_12665,N_12705);
nor U13059 (N_13059,N_12223,N_12271);
or U13060 (N_13060,N_12014,N_12286);
xor U13061 (N_13061,N_12529,N_12464);
xnor U13062 (N_13062,N_12703,N_12579);
nand U13063 (N_13063,N_12067,N_12285);
and U13064 (N_13064,N_12423,N_12686);
and U13065 (N_13065,N_12287,N_12772);
or U13066 (N_13066,N_12717,N_12129);
or U13067 (N_13067,N_12724,N_12178);
nor U13068 (N_13068,N_12696,N_12018);
xnor U13069 (N_13069,N_12713,N_12542);
and U13070 (N_13070,N_12455,N_12098);
and U13071 (N_13071,N_12296,N_12253);
nor U13072 (N_13072,N_12576,N_12037);
nand U13073 (N_13073,N_12549,N_12268);
nand U13074 (N_13074,N_12091,N_12762);
and U13075 (N_13075,N_12446,N_12372);
nor U13076 (N_13076,N_12238,N_12668);
or U13077 (N_13077,N_12202,N_12366);
nand U13078 (N_13078,N_12688,N_12203);
xor U13079 (N_13079,N_12307,N_12333);
and U13080 (N_13080,N_12451,N_12181);
and U13081 (N_13081,N_12133,N_12175);
and U13082 (N_13082,N_12600,N_12332);
or U13083 (N_13083,N_12107,N_12754);
nor U13084 (N_13084,N_12026,N_12160);
and U13085 (N_13085,N_12122,N_12005);
or U13086 (N_13086,N_12748,N_12156);
nand U13087 (N_13087,N_12430,N_12726);
nand U13088 (N_13088,N_12276,N_12659);
nand U13089 (N_13089,N_12262,N_12503);
nand U13090 (N_13090,N_12553,N_12308);
or U13091 (N_13091,N_12127,N_12235);
nor U13092 (N_13092,N_12751,N_12674);
or U13093 (N_13093,N_12585,N_12741);
and U13094 (N_13094,N_12370,N_12168);
and U13095 (N_13095,N_12274,N_12749);
and U13096 (N_13096,N_12601,N_12028);
and U13097 (N_13097,N_12682,N_12357);
xnor U13098 (N_13098,N_12259,N_12590);
or U13099 (N_13099,N_12729,N_12049);
or U13100 (N_13100,N_12162,N_12323);
and U13101 (N_13101,N_12248,N_12435);
xor U13102 (N_13102,N_12534,N_12329);
nor U13103 (N_13103,N_12291,N_12012);
xnor U13104 (N_13104,N_12131,N_12004);
or U13105 (N_13105,N_12195,N_12076);
or U13106 (N_13106,N_12716,N_12025);
and U13107 (N_13107,N_12731,N_12760);
nor U13108 (N_13108,N_12391,N_12473);
nor U13109 (N_13109,N_12220,N_12636);
nand U13110 (N_13110,N_12021,N_12574);
nor U13111 (N_13111,N_12482,N_12546);
nand U13112 (N_13112,N_12011,N_12728);
xnor U13113 (N_13113,N_12779,N_12460);
and U13114 (N_13114,N_12182,N_12469);
nor U13115 (N_13115,N_12173,N_12300);
or U13116 (N_13116,N_12487,N_12608);
nor U13117 (N_13117,N_12532,N_12279);
xor U13118 (N_13118,N_12769,N_12562);
or U13119 (N_13119,N_12240,N_12527);
and U13120 (N_13120,N_12619,N_12041);
xor U13121 (N_13121,N_12437,N_12406);
nand U13122 (N_13122,N_12380,N_12592);
nand U13123 (N_13123,N_12256,N_12617);
and U13124 (N_13124,N_12525,N_12038);
or U13125 (N_13125,N_12786,N_12120);
xor U13126 (N_13126,N_12501,N_12432);
nand U13127 (N_13127,N_12328,N_12189);
xnor U13128 (N_13128,N_12293,N_12154);
or U13129 (N_13129,N_12061,N_12199);
and U13130 (N_13130,N_12578,N_12282);
nand U13131 (N_13131,N_12799,N_12330);
nand U13132 (N_13132,N_12249,N_12700);
nand U13133 (N_13133,N_12442,N_12096);
and U13134 (N_13134,N_12733,N_12554);
xor U13135 (N_13135,N_12007,N_12147);
nor U13136 (N_13136,N_12115,N_12775);
or U13137 (N_13137,N_12060,N_12078);
or U13138 (N_13138,N_12392,N_12565);
nand U13139 (N_13139,N_12036,N_12474);
or U13140 (N_13140,N_12197,N_12664);
nand U13141 (N_13141,N_12108,N_12676);
nor U13142 (N_13142,N_12104,N_12051);
or U13143 (N_13143,N_12490,N_12321);
nand U13144 (N_13144,N_12408,N_12635);
or U13145 (N_13145,N_12653,N_12596);
xnor U13146 (N_13146,N_12434,N_12459);
xor U13147 (N_13147,N_12466,N_12179);
xnor U13148 (N_13148,N_12016,N_12656);
or U13149 (N_13149,N_12428,N_12658);
and U13150 (N_13150,N_12707,N_12135);
nand U13151 (N_13151,N_12342,N_12667);
nand U13152 (N_13152,N_12467,N_12714);
nand U13153 (N_13153,N_12510,N_12294);
and U13154 (N_13154,N_12097,N_12153);
nor U13155 (N_13155,N_12730,N_12498);
xor U13156 (N_13156,N_12278,N_12457);
nor U13157 (N_13157,N_12186,N_12416);
nand U13158 (N_13158,N_12148,N_12788);
xnor U13159 (N_13159,N_12740,N_12794);
xor U13160 (N_13160,N_12080,N_12586);
and U13161 (N_13161,N_12337,N_12618);
xor U13162 (N_13162,N_12753,N_12566);
xor U13163 (N_13163,N_12198,N_12006);
xnor U13164 (N_13164,N_12652,N_12188);
xor U13165 (N_13165,N_12260,N_12531);
and U13166 (N_13166,N_12756,N_12678);
xor U13167 (N_13167,N_12169,N_12417);
xor U13168 (N_13168,N_12693,N_12683);
nand U13169 (N_13169,N_12044,N_12226);
or U13170 (N_13170,N_12628,N_12368);
xnor U13171 (N_13171,N_12336,N_12632);
or U13172 (N_13172,N_12377,N_12495);
xnor U13173 (N_13173,N_12752,N_12692);
xnor U13174 (N_13174,N_12541,N_12224);
nor U13175 (N_13175,N_12039,N_12739);
or U13176 (N_13176,N_12054,N_12327);
and U13177 (N_13177,N_12192,N_12301);
or U13178 (N_13178,N_12583,N_12165);
or U13179 (N_13179,N_12345,N_12413);
and U13180 (N_13180,N_12319,N_12695);
xnor U13181 (N_13181,N_12648,N_12325);
nand U13182 (N_13182,N_12003,N_12040);
nand U13183 (N_13183,N_12265,N_12349);
or U13184 (N_13184,N_12373,N_12412);
xnor U13185 (N_13185,N_12609,N_12074);
nor U13186 (N_13186,N_12079,N_12604);
nor U13187 (N_13187,N_12239,N_12369);
xor U13188 (N_13188,N_12243,N_12376);
xor U13189 (N_13189,N_12657,N_12295);
and U13190 (N_13190,N_12277,N_12454);
and U13191 (N_13191,N_12356,N_12375);
and U13192 (N_13192,N_12302,N_12000);
or U13193 (N_13193,N_12314,N_12141);
xnor U13194 (N_13194,N_12066,N_12516);
nand U13195 (N_13195,N_12055,N_12640);
nand U13196 (N_13196,N_12317,N_12471);
or U13197 (N_13197,N_12594,N_12083);
and U13198 (N_13198,N_12227,N_12791);
or U13199 (N_13199,N_12309,N_12174);
or U13200 (N_13200,N_12551,N_12170);
xnor U13201 (N_13201,N_12743,N_12337);
or U13202 (N_13202,N_12485,N_12460);
and U13203 (N_13203,N_12159,N_12680);
or U13204 (N_13204,N_12199,N_12101);
or U13205 (N_13205,N_12520,N_12431);
nor U13206 (N_13206,N_12468,N_12162);
nor U13207 (N_13207,N_12310,N_12072);
xnor U13208 (N_13208,N_12183,N_12722);
nand U13209 (N_13209,N_12727,N_12331);
nand U13210 (N_13210,N_12038,N_12076);
nor U13211 (N_13211,N_12455,N_12076);
nand U13212 (N_13212,N_12535,N_12754);
nand U13213 (N_13213,N_12762,N_12582);
xnor U13214 (N_13214,N_12103,N_12091);
nand U13215 (N_13215,N_12549,N_12213);
and U13216 (N_13216,N_12082,N_12074);
nand U13217 (N_13217,N_12597,N_12226);
and U13218 (N_13218,N_12270,N_12144);
or U13219 (N_13219,N_12576,N_12088);
and U13220 (N_13220,N_12698,N_12365);
and U13221 (N_13221,N_12258,N_12083);
or U13222 (N_13222,N_12662,N_12564);
nor U13223 (N_13223,N_12721,N_12682);
nor U13224 (N_13224,N_12358,N_12218);
and U13225 (N_13225,N_12650,N_12302);
nand U13226 (N_13226,N_12441,N_12612);
or U13227 (N_13227,N_12108,N_12563);
and U13228 (N_13228,N_12114,N_12086);
xor U13229 (N_13229,N_12351,N_12461);
or U13230 (N_13230,N_12772,N_12493);
nor U13231 (N_13231,N_12156,N_12475);
or U13232 (N_13232,N_12126,N_12673);
and U13233 (N_13233,N_12463,N_12281);
nand U13234 (N_13234,N_12195,N_12662);
xor U13235 (N_13235,N_12286,N_12529);
and U13236 (N_13236,N_12410,N_12754);
and U13237 (N_13237,N_12703,N_12791);
xnor U13238 (N_13238,N_12555,N_12237);
xor U13239 (N_13239,N_12197,N_12608);
nor U13240 (N_13240,N_12741,N_12278);
nor U13241 (N_13241,N_12420,N_12364);
nor U13242 (N_13242,N_12341,N_12797);
and U13243 (N_13243,N_12798,N_12604);
and U13244 (N_13244,N_12324,N_12783);
and U13245 (N_13245,N_12551,N_12485);
nand U13246 (N_13246,N_12124,N_12463);
and U13247 (N_13247,N_12377,N_12703);
nand U13248 (N_13248,N_12778,N_12150);
and U13249 (N_13249,N_12477,N_12177);
or U13250 (N_13250,N_12619,N_12528);
or U13251 (N_13251,N_12021,N_12191);
or U13252 (N_13252,N_12241,N_12479);
or U13253 (N_13253,N_12441,N_12318);
or U13254 (N_13254,N_12153,N_12353);
nand U13255 (N_13255,N_12164,N_12402);
nand U13256 (N_13256,N_12489,N_12470);
and U13257 (N_13257,N_12231,N_12776);
nor U13258 (N_13258,N_12079,N_12340);
nand U13259 (N_13259,N_12214,N_12721);
and U13260 (N_13260,N_12681,N_12719);
nor U13261 (N_13261,N_12193,N_12462);
xor U13262 (N_13262,N_12560,N_12026);
nor U13263 (N_13263,N_12196,N_12300);
and U13264 (N_13264,N_12719,N_12307);
nand U13265 (N_13265,N_12551,N_12167);
nand U13266 (N_13266,N_12147,N_12571);
and U13267 (N_13267,N_12139,N_12203);
and U13268 (N_13268,N_12254,N_12434);
or U13269 (N_13269,N_12119,N_12004);
and U13270 (N_13270,N_12144,N_12524);
xor U13271 (N_13271,N_12239,N_12108);
nand U13272 (N_13272,N_12796,N_12242);
or U13273 (N_13273,N_12623,N_12494);
nand U13274 (N_13274,N_12389,N_12350);
xnor U13275 (N_13275,N_12006,N_12695);
or U13276 (N_13276,N_12169,N_12789);
and U13277 (N_13277,N_12455,N_12377);
and U13278 (N_13278,N_12100,N_12421);
xnor U13279 (N_13279,N_12796,N_12327);
and U13280 (N_13280,N_12665,N_12330);
or U13281 (N_13281,N_12084,N_12369);
or U13282 (N_13282,N_12035,N_12145);
and U13283 (N_13283,N_12584,N_12601);
xor U13284 (N_13284,N_12530,N_12373);
nand U13285 (N_13285,N_12100,N_12299);
nor U13286 (N_13286,N_12182,N_12403);
xnor U13287 (N_13287,N_12038,N_12107);
and U13288 (N_13288,N_12064,N_12574);
and U13289 (N_13289,N_12096,N_12492);
and U13290 (N_13290,N_12287,N_12605);
or U13291 (N_13291,N_12018,N_12327);
and U13292 (N_13292,N_12751,N_12472);
nand U13293 (N_13293,N_12664,N_12083);
and U13294 (N_13294,N_12381,N_12264);
nor U13295 (N_13295,N_12406,N_12369);
and U13296 (N_13296,N_12069,N_12438);
nor U13297 (N_13297,N_12665,N_12750);
nor U13298 (N_13298,N_12716,N_12459);
or U13299 (N_13299,N_12116,N_12084);
or U13300 (N_13300,N_12333,N_12413);
nand U13301 (N_13301,N_12566,N_12710);
or U13302 (N_13302,N_12126,N_12563);
nor U13303 (N_13303,N_12403,N_12103);
or U13304 (N_13304,N_12290,N_12626);
and U13305 (N_13305,N_12446,N_12200);
and U13306 (N_13306,N_12627,N_12149);
nor U13307 (N_13307,N_12499,N_12253);
nor U13308 (N_13308,N_12443,N_12428);
or U13309 (N_13309,N_12131,N_12650);
and U13310 (N_13310,N_12666,N_12301);
xor U13311 (N_13311,N_12071,N_12578);
or U13312 (N_13312,N_12130,N_12385);
or U13313 (N_13313,N_12512,N_12744);
nor U13314 (N_13314,N_12229,N_12068);
and U13315 (N_13315,N_12677,N_12159);
nor U13316 (N_13316,N_12136,N_12673);
xor U13317 (N_13317,N_12475,N_12446);
nor U13318 (N_13318,N_12553,N_12197);
or U13319 (N_13319,N_12036,N_12337);
nand U13320 (N_13320,N_12630,N_12033);
xnor U13321 (N_13321,N_12011,N_12069);
xnor U13322 (N_13322,N_12659,N_12466);
and U13323 (N_13323,N_12020,N_12346);
or U13324 (N_13324,N_12316,N_12106);
nand U13325 (N_13325,N_12205,N_12045);
and U13326 (N_13326,N_12581,N_12315);
and U13327 (N_13327,N_12784,N_12514);
nor U13328 (N_13328,N_12410,N_12274);
or U13329 (N_13329,N_12106,N_12740);
and U13330 (N_13330,N_12298,N_12729);
nand U13331 (N_13331,N_12636,N_12531);
or U13332 (N_13332,N_12174,N_12331);
and U13333 (N_13333,N_12098,N_12142);
xnor U13334 (N_13334,N_12280,N_12729);
nor U13335 (N_13335,N_12192,N_12415);
nor U13336 (N_13336,N_12330,N_12094);
xnor U13337 (N_13337,N_12658,N_12765);
or U13338 (N_13338,N_12061,N_12481);
and U13339 (N_13339,N_12077,N_12483);
nand U13340 (N_13340,N_12514,N_12509);
xnor U13341 (N_13341,N_12661,N_12615);
nand U13342 (N_13342,N_12655,N_12771);
or U13343 (N_13343,N_12373,N_12311);
nor U13344 (N_13344,N_12595,N_12773);
or U13345 (N_13345,N_12499,N_12660);
and U13346 (N_13346,N_12712,N_12286);
or U13347 (N_13347,N_12208,N_12446);
nand U13348 (N_13348,N_12711,N_12485);
xor U13349 (N_13349,N_12548,N_12764);
and U13350 (N_13350,N_12410,N_12010);
or U13351 (N_13351,N_12262,N_12130);
nor U13352 (N_13352,N_12584,N_12273);
xnor U13353 (N_13353,N_12502,N_12026);
nor U13354 (N_13354,N_12482,N_12086);
xnor U13355 (N_13355,N_12134,N_12586);
or U13356 (N_13356,N_12789,N_12023);
nor U13357 (N_13357,N_12666,N_12542);
nand U13358 (N_13358,N_12676,N_12465);
nor U13359 (N_13359,N_12348,N_12799);
and U13360 (N_13360,N_12414,N_12009);
nand U13361 (N_13361,N_12308,N_12519);
nand U13362 (N_13362,N_12663,N_12395);
or U13363 (N_13363,N_12386,N_12290);
nor U13364 (N_13364,N_12769,N_12323);
xnor U13365 (N_13365,N_12128,N_12678);
nand U13366 (N_13366,N_12209,N_12052);
xor U13367 (N_13367,N_12606,N_12435);
nor U13368 (N_13368,N_12030,N_12459);
or U13369 (N_13369,N_12764,N_12086);
nor U13370 (N_13370,N_12087,N_12022);
nand U13371 (N_13371,N_12202,N_12023);
and U13372 (N_13372,N_12405,N_12016);
and U13373 (N_13373,N_12038,N_12014);
nand U13374 (N_13374,N_12096,N_12323);
or U13375 (N_13375,N_12561,N_12062);
nand U13376 (N_13376,N_12374,N_12683);
and U13377 (N_13377,N_12499,N_12468);
nand U13378 (N_13378,N_12568,N_12203);
xor U13379 (N_13379,N_12598,N_12787);
nor U13380 (N_13380,N_12293,N_12786);
or U13381 (N_13381,N_12335,N_12499);
nor U13382 (N_13382,N_12431,N_12506);
or U13383 (N_13383,N_12656,N_12698);
and U13384 (N_13384,N_12172,N_12432);
or U13385 (N_13385,N_12717,N_12089);
and U13386 (N_13386,N_12245,N_12531);
or U13387 (N_13387,N_12377,N_12073);
nand U13388 (N_13388,N_12212,N_12134);
and U13389 (N_13389,N_12245,N_12214);
nor U13390 (N_13390,N_12636,N_12210);
and U13391 (N_13391,N_12673,N_12717);
nand U13392 (N_13392,N_12744,N_12721);
nand U13393 (N_13393,N_12509,N_12779);
or U13394 (N_13394,N_12219,N_12647);
nor U13395 (N_13395,N_12375,N_12470);
nor U13396 (N_13396,N_12215,N_12307);
nand U13397 (N_13397,N_12133,N_12348);
nor U13398 (N_13398,N_12033,N_12128);
and U13399 (N_13399,N_12550,N_12170);
nand U13400 (N_13400,N_12352,N_12359);
nand U13401 (N_13401,N_12716,N_12730);
xnor U13402 (N_13402,N_12792,N_12621);
nand U13403 (N_13403,N_12308,N_12005);
nor U13404 (N_13404,N_12789,N_12270);
and U13405 (N_13405,N_12506,N_12249);
nor U13406 (N_13406,N_12439,N_12778);
nor U13407 (N_13407,N_12595,N_12238);
and U13408 (N_13408,N_12125,N_12735);
or U13409 (N_13409,N_12781,N_12711);
or U13410 (N_13410,N_12482,N_12387);
and U13411 (N_13411,N_12068,N_12376);
or U13412 (N_13412,N_12673,N_12523);
xnor U13413 (N_13413,N_12654,N_12759);
nor U13414 (N_13414,N_12294,N_12159);
and U13415 (N_13415,N_12357,N_12686);
and U13416 (N_13416,N_12688,N_12698);
and U13417 (N_13417,N_12487,N_12453);
or U13418 (N_13418,N_12517,N_12652);
or U13419 (N_13419,N_12141,N_12796);
nand U13420 (N_13420,N_12546,N_12638);
and U13421 (N_13421,N_12000,N_12099);
or U13422 (N_13422,N_12778,N_12723);
xnor U13423 (N_13423,N_12210,N_12471);
xnor U13424 (N_13424,N_12286,N_12390);
xor U13425 (N_13425,N_12174,N_12719);
nor U13426 (N_13426,N_12054,N_12299);
or U13427 (N_13427,N_12612,N_12071);
xnor U13428 (N_13428,N_12168,N_12076);
nand U13429 (N_13429,N_12319,N_12106);
xor U13430 (N_13430,N_12777,N_12572);
nor U13431 (N_13431,N_12420,N_12705);
and U13432 (N_13432,N_12276,N_12066);
or U13433 (N_13433,N_12073,N_12126);
and U13434 (N_13434,N_12505,N_12230);
nor U13435 (N_13435,N_12197,N_12139);
nand U13436 (N_13436,N_12101,N_12697);
or U13437 (N_13437,N_12437,N_12693);
nor U13438 (N_13438,N_12547,N_12089);
and U13439 (N_13439,N_12492,N_12670);
and U13440 (N_13440,N_12141,N_12233);
and U13441 (N_13441,N_12430,N_12541);
xnor U13442 (N_13442,N_12076,N_12181);
and U13443 (N_13443,N_12300,N_12203);
or U13444 (N_13444,N_12725,N_12792);
nand U13445 (N_13445,N_12238,N_12632);
nor U13446 (N_13446,N_12438,N_12351);
or U13447 (N_13447,N_12489,N_12683);
nand U13448 (N_13448,N_12318,N_12723);
nor U13449 (N_13449,N_12599,N_12644);
or U13450 (N_13450,N_12422,N_12271);
nor U13451 (N_13451,N_12764,N_12386);
or U13452 (N_13452,N_12166,N_12394);
nand U13453 (N_13453,N_12157,N_12406);
and U13454 (N_13454,N_12513,N_12143);
or U13455 (N_13455,N_12086,N_12766);
or U13456 (N_13456,N_12139,N_12771);
nand U13457 (N_13457,N_12231,N_12749);
xor U13458 (N_13458,N_12471,N_12681);
nor U13459 (N_13459,N_12163,N_12780);
and U13460 (N_13460,N_12644,N_12561);
and U13461 (N_13461,N_12369,N_12064);
xnor U13462 (N_13462,N_12442,N_12534);
nor U13463 (N_13463,N_12715,N_12582);
xor U13464 (N_13464,N_12724,N_12693);
and U13465 (N_13465,N_12203,N_12311);
and U13466 (N_13466,N_12227,N_12394);
xnor U13467 (N_13467,N_12631,N_12011);
nor U13468 (N_13468,N_12459,N_12599);
xor U13469 (N_13469,N_12788,N_12221);
nand U13470 (N_13470,N_12523,N_12797);
nand U13471 (N_13471,N_12175,N_12789);
xor U13472 (N_13472,N_12204,N_12789);
xor U13473 (N_13473,N_12039,N_12289);
and U13474 (N_13474,N_12033,N_12185);
xnor U13475 (N_13475,N_12533,N_12616);
nand U13476 (N_13476,N_12229,N_12618);
and U13477 (N_13477,N_12762,N_12758);
or U13478 (N_13478,N_12683,N_12301);
and U13479 (N_13479,N_12511,N_12244);
nand U13480 (N_13480,N_12565,N_12184);
xnor U13481 (N_13481,N_12668,N_12371);
and U13482 (N_13482,N_12149,N_12226);
nor U13483 (N_13483,N_12748,N_12086);
and U13484 (N_13484,N_12148,N_12138);
xor U13485 (N_13485,N_12384,N_12504);
and U13486 (N_13486,N_12481,N_12088);
nor U13487 (N_13487,N_12375,N_12279);
nor U13488 (N_13488,N_12389,N_12518);
xnor U13489 (N_13489,N_12368,N_12667);
nor U13490 (N_13490,N_12347,N_12699);
nand U13491 (N_13491,N_12459,N_12798);
nand U13492 (N_13492,N_12359,N_12624);
or U13493 (N_13493,N_12761,N_12358);
xor U13494 (N_13494,N_12081,N_12154);
or U13495 (N_13495,N_12404,N_12134);
xnor U13496 (N_13496,N_12377,N_12358);
and U13497 (N_13497,N_12482,N_12248);
or U13498 (N_13498,N_12752,N_12245);
xor U13499 (N_13499,N_12228,N_12756);
xor U13500 (N_13500,N_12514,N_12796);
xnor U13501 (N_13501,N_12764,N_12177);
nor U13502 (N_13502,N_12034,N_12366);
nand U13503 (N_13503,N_12517,N_12187);
nand U13504 (N_13504,N_12598,N_12368);
nor U13505 (N_13505,N_12506,N_12350);
nor U13506 (N_13506,N_12783,N_12066);
or U13507 (N_13507,N_12206,N_12022);
nor U13508 (N_13508,N_12353,N_12401);
xor U13509 (N_13509,N_12156,N_12263);
nor U13510 (N_13510,N_12075,N_12702);
or U13511 (N_13511,N_12577,N_12236);
nand U13512 (N_13512,N_12104,N_12071);
or U13513 (N_13513,N_12351,N_12118);
and U13514 (N_13514,N_12796,N_12083);
or U13515 (N_13515,N_12519,N_12221);
and U13516 (N_13516,N_12285,N_12342);
nor U13517 (N_13517,N_12441,N_12615);
nor U13518 (N_13518,N_12515,N_12065);
and U13519 (N_13519,N_12341,N_12659);
nor U13520 (N_13520,N_12064,N_12538);
nor U13521 (N_13521,N_12251,N_12346);
nor U13522 (N_13522,N_12219,N_12485);
nand U13523 (N_13523,N_12392,N_12750);
or U13524 (N_13524,N_12681,N_12424);
nand U13525 (N_13525,N_12106,N_12190);
and U13526 (N_13526,N_12095,N_12364);
or U13527 (N_13527,N_12415,N_12058);
or U13528 (N_13528,N_12604,N_12366);
nand U13529 (N_13529,N_12001,N_12594);
xnor U13530 (N_13530,N_12374,N_12760);
xnor U13531 (N_13531,N_12344,N_12593);
and U13532 (N_13532,N_12522,N_12643);
xor U13533 (N_13533,N_12601,N_12776);
and U13534 (N_13534,N_12010,N_12143);
or U13535 (N_13535,N_12068,N_12353);
or U13536 (N_13536,N_12491,N_12347);
nand U13537 (N_13537,N_12600,N_12510);
or U13538 (N_13538,N_12482,N_12195);
xor U13539 (N_13539,N_12491,N_12463);
or U13540 (N_13540,N_12198,N_12738);
nand U13541 (N_13541,N_12169,N_12630);
nor U13542 (N_13542,N_12584,N_12261);
and U13543 (N_13543,N_12189,N_12507);
nor U13544 (N_13544,N_12595,N_12050);
xnor U13545 (N_13545,N_12436,N_12347);
xnor U13546 (N_13546,N_12086,N_12234);
nand U13547 (N_13547,N_12277,N_12493);
nor U13548 (N_13548,N_12305,N_12109);
xnor U13549 (N_13549,N_12750,N_12297);
nor U13550 (N_13550,N_12682,N_12306);
nor U13551 (N_13551,N_12144,N_12382);
and U13552 (N_13552,N_12282,N_12686);
nand U13553 (N_13553,N_12731,N_12178);
nor U13554 (N_13554,N_12109,N_12381);
xnor U13555 (N_13555,N_12386,N_12460);
xnor U13556 (N_13556,N_12445,N_12151);
xor U13557 (N_13557,N_12149,N_12155);
and U13558 (N_13558,N_12590,N_12653);
xor U13559 (N_13559,N_12519,N_12576);
or U13560 (N_13560,N_12527,N_12267);
and U13561 (N_13561,N_12120,N_12787);
xnor U13562 (N_13562,N_12787,N_12114);
or U13563 (N_13563,N_12441,N_12793);
nand U13564 (N_13564,N_12062,N_12634);
nand U13565 (N_13565,N_12448,N_12747);
xor U13566 (N_13566,N_12648,N_12306);
and U13567 (N_13567,N_12645,N_12320);
and U13568 (N_13568,N_12535,N_12672);
xnor U13569 (N_13569,N_12286,N_12061);
xnor U13570 (N_13570,N_12151,N_12053);
nand U13571 (N_13571,N_12220,N_12229);
xor U13572 (N_13572,N_12690,N_12293);
nor U13573 (N_13573,N_12769,N_12209);
or U13574 (N_13574,N_12762,N_12185);
nor U13575 (N_13575,N_12603,N_12411);
and U13576 (N_13576,N_12143,N_12003);
nor U13577 (N_13577,N_12168,N_12148);
nor U13578 (N_13578,N_12216,N_12654);
nor U13579 (N_13579,N_12161,N_12670);
nand U13580 (N_13580,N_12625,N_12271);
xor U13581 (N_13581,N_12307,N_12184);
and U13582 (N_13582,N_12271,N_12555);
nand U13583 (N_13583,N_12476,N_12120);
xor U13584 (N_13584,N_12320,N_12034);
xor U13585 (N_13585,N_12251,N_12716);
and U13586 (N_13586,N_12106,N_12664);
and U13587 (N_13587,N_12131,N_12426);
and U13588 (N_13588,N_12638,N_12019);
nand U13589 (N_13589,N_12069,N_12035);
xnor U13590 (N_13590,N_12526,N_12568);
xor U13591 (N_13591,N_12791,N_12329);
or U13592 (N_13592,N_12266,N_12158);
nand U13593 (N_13593,N_12453,N_12212);
nor U13594 (N_13594,N_12183,N_12533);
and U13595 (N_13595,N_12662,N_12140);
or U13596 (N_13596,N_12316,N_12728);
nand U13597 (N_13597,N_12722,N_12567);
xnor U13598 (N_13598,N_12595,N_12344);
and U13599 (N_13599,N_12640,N_12551);
and U13600 (N_13600,N_13032,N_13339);
and U13601 (N_13601,N_13035,N_13100);
and U13602 (N_13602,N_13120,N_13315);
xnor U13603 (N_13603,N_12844,N_13252);
and U13604 (N_13604,N_13162,N_13343);
xnor U13605 (N_13605,N_13396,N_13084);
nand U13606 (N_13606,N_13561,N_13182);
nor U13607 (N_13607,N_13390,N_13360);
nor U13608 (N_13608,N_13481,N_13246);
or U13609 (N_13609,N_13357,N_12828);
or U13610 (N_13610,N_13526,N_12934);
or U13611 (N_13611,N_13143,N_12911);
nand U13612 (N_13612,N_12964,N_12865);
nor U13613 (N_13613,N_13308,N_13046);
xnor U13614 (N_13614,N_12870,N_12922);
xor U13615 (N_13615,N_13301,N_13091);
or U13616 (N_13616,N_12990,N_13082);
xor U13617 (N_13617,N_13057,N_13061);
nor U13618 (N_13618,N_13412,N_13038);
nor U13619 (N_13619,N_12923,N_12950);
nor U13620 (N_13620,N_13423,N_13011);
and U13621 (N_13621,N_13063,N_12856);
nand U13622 (N_13622,N_13025,N_12997);
or U13623 (N_13623,N_13362,N_13273);
nand U13624 (N_13624,N_12993,N_13587);
nand U13625 (N_13625,N_12904,N_13494);
nand U13626 (N_13626,N_12988,N_13004);
xnor U13627 (N_13627,N_13275,N_13070);
or U13628 (N_13628,N_13575,N_13230);
nor U13629 (N_13629,N_12814,N_13271);
xnor U13630 (N_13630,N_13260,N_13433);
or U13631 (N_13631,N_13580,N_13332);
and U13632 (N_13632,N_12836,N_13147);
or U13633 (N_13633,N_13438,N_13139);
xnor U13634 (N_13634,N_12889,N_13333);
xnor U13635 (N_13635,N_12945,N_12987);
xnor U13636 (N_13636,N_13242,N_13165);
xor U13637 (N_13637,N_12872,N_12864);
nor U13638 (N_13638,N_13487,N_13078);
nand U13639 (N_13639,N_13248,N_13180);
or U13640 (N_13640,N_13312,N_13116);
or U13641 (N_13641,N_13124,N_12924);
or U13642 (N_13642,N_13527,N_13037);
xor U13643 (N_13643,N_12921,N_13524);
xnor U13644 (N_13644,N_12850,N_13566);
and U13645 (N_13645,N_13572,N_13316);
and U13646 (N_13646,N_13015,N_13207);
nor U13647 (N_13647,N_13356,N_13555);
and U13648 (N_13648,N_13536,N_13504);
nor U13649 (N_13649,N_13384,N_13266);
nor U13650 (N_13650,N_12937,N_13073);
xnor U13651 (N_13651,N_13382,N_12959);
and U13652 (N_13652,N_13101,N_13530);
nand U13653 (N_13653,N_13269,N_13518);
nand U13654 (N_13654,N_13469,N_13379);
and U13655 (N_13655,N_13202,N_13355);
nor U13656 (N_13656,N_12809,N_13102);
and U13657 (N_13657,N_13065,N_13464);
and U13658 (N_13658,N_12825,N_13499);
nor U13659 (N_13659,N_13021,N_13553);
nor U13660 (N_13660,N_13565,N_13589);
xor U13661 (N_13661,N_13346,N_13562);
or U13662 (N_13662,N_12813,N_12855);
xnor U13663 (N_13663,N_13259,N_12832);
xor U13664 (N_13664,N_12891,N_13130);
xnor U13665 (N_13665,N_12886,N_12831);
and U13666 (N_13666,N_13321,N_12866);
or U13667 (N_13667,N_13176,N_12994);
and U13668 (N_13668,N_12970,N_13571);
nor U13669 (N_13669,N_13008,N_13159);
or U13670 (N_13670,N_13445,N_12810);
and U13671 (N_13671,N_13532,N_13185);
xnor U13672 (N_13672,N_13576,N_12868);
or U13673 (N_13673,N_12874,N_13245);
and U13674 (N_13674,N_13533,N_13123);
nor U13675 (N_13675,N_13054,N_13493);
nand U13676 (N_13676,N_12883,N_13393);
or U13677 (N_13677,N_12927,N_13387);
nand U13678 (N_13678,N_13178,N_13585);
nand U13679 (N_13679,N_12913,N_13164);
and U13680 (N_13680,N_12956,N_13331);
nor U13681 (N_13681,N_13388,N_13090);
nor U13682 (N_13682,N_12821,N_12820);
xor U13683 (N_13683,N_13407,N_13426);
xnor U13684 (N_13684,N_12857,N_13599);
nand U13685 (N_13685,N_13089,N_12806);
xor U13686 (N_13686,N_13206,N_13535);
xor U13687 (N_13687,N_13363,N_13353);
nor U13688 (N_13688,N_12816,N_13386);
nor U13689 (N_13689,N_13294,N_13148);
nand U13690 (N_13690,N_13432,N_12852);
nand U13691 (N_13691,N_13459,N_13117);
nor U13692 (N_13692,N_13276,N_13471);
and U13693 (N_13693,N_13431,N_13344);
or U13694 (N_13694,N_13278,N_12819);
and U13695 (N_13695,N_13436,N_13220);
or U13696 (N_13696,N_13106,N_13036);
nand U13697 (N_13697,N_12869,N_13027);
xor U13698 (N_13698,N_13413,N_13597);
nand U13699 (N_13699,N_13411,N_13502);
xnor U13700 (N_13700,N_12878,N_13099);
xor U13701 (N_13701,N_13068,N_13175);
nand U13702 (N_13702,N_13500,N_13244);
xor U13703 (N_13703,N_13018,N_13395);
nor U13704 (N_13704,N_13479,N_13033);
nand U13705 (N_13705,N_13152,N_13199);
nor U13706 (N_13706,N_12811,N_13087);
nand U13707 (N_13707,N_12926,N_12902);
xnor U13708 (N_13708,N_13476,N_13560);
xnor U13709 (N_13709,N_12953,N_13492);
nor U13710 (N_13710,N_13028,N_13593);
or U13711 (N_13711,N_13149,N_13108);
nand U13712 (N_13712,N_12962,N_13019);
and U13713 (N_13713,N_13531,N_13095);
xnor U13714 (N_13714,N_13171,N_13534);
xnor U13715 (N_13715,N_13286,N_13132);
nor U13716 (N_13716,N_13461,N_13127);
nand U13717 (N_13717,N_13482,N_13409);
nand U13718 (N_13718,N_13138,N_13240);
nand U13719 (N_13719,N_13277,N_13193);
xnor U13720 (N_13720,N_13056,N_12834);
xnor U13721 (N_13721,N_13591,N_13086);
and U13722 (N_13722,N_12933,N_13201);
and U13723 (N_13723,N_13369,N_13341);
nand U13724 (N_13724,N_12955,N_13263);
or U13725 (N_13725,N_12817,N_13421);
nand U13726 (N_13726,N_13398,N_13003);
or U13727 (N_13727,N_12971,N_13249);
and U13728 (N_13728,N_13510,N_13214);
or U13729 (N_13729,N_13247,N_13558);
nor U13730 (N_13730,N_13596,N_12888);
xnor U13731 (N_13731,N_13170,N_13236);
nand U13732 (N_13732,N_13505,N_12925);
nor U13733 (N_13733,N_13062,N_12838);
nor U13734 (N_13734,N_12835,N_12966);
and U13735 (N_13735,N_13463,N_13320);
xnor U13736 (N_13736,N_13153,N_13034);
xor U13737 (N_13737,N_13598,N_13352);
or U13738 (N_13738,N_13402,N_12824);
and U13739 (N_13739,N_13231,N_13428);
xor U13740 (N_13740,N_13354,N_12973);
and U13741 (N_13741,N_12960,N_13458);
nor U13742 (N_13742,N_13173,N_13543);
xnor U13743 (N_13743,N_12875,N_13071);
nand U13744 (N_13744,N_13342,N_12845);
xor U13745 (N_13745,N_12967,N_12808);
and U13746 (N_13746,N_13590,N_13416);
nand U13747 (N_13747,N_12939,N_13523);
and U13748 (N_13748,N_13514,N_12860);
nand U13749 (N_13749,N_13313,N_13323);
nand U13750 (N_13750,N_13026,N_13468);
or U13751 (N_13751,N_13140,N_12903);
xnor U13752 (N_13752,N_13298,N_12918);
xnor U13753 (N_13753,N_13299,N_12910);
and U13754 (N_13754,N_13072,N_13020);
or U13755 (N_13755,N_12989,N_13043);
nand U13756 (N_13756,N_13578,N_13389);
and U13757 (N_13757,N_13133,N_13528);
nand U13758 (N_13758,N_13049,N_13234);
xnor U13759 (N_13759,N_13371,N_13425);
xor U13760 (N_13760,N_13009,N_13155);
nand U13761 (N_13761,N_12848,N_13290);
or U13762 (N_13762,N_13196,N_13097);
nand U13763 (N_13763,N_13408,N_13174);
xnor U13764 (N_13764,N_13473,N_13373);
or U13765 (N_13765,N_12839,N_13039);
or U13766 (N_13766,N_13592,N_13168);
nand U13767 (N_13767,N_13268,N_13282);
and U13768 (N_13768,N_13465,N_13564);
and U13769 (N_13769,N_13550,N_13309);
nor U13770 (N_13770,N_13417,N_13349);
nor U13771 (N_13771,N_12944,N_13573);
and U13772 (N_13772,N_12827,N_13262);
nor U13773 (N_13773,N_13048,N_13114);
nand U13774 (N_13774,N_12840,N_12928);
and U13775 (N_13775,N_13005,N_13434);
xor U13776 (N_13776,N_13053,N_13151);
and U13777 (N_13777,N_13258,N_13347);
nand U13778 (N_13778,N_12841,N_12912);
nand U13779 (N_13779,N_13013,N_12807);
or U13780 (N_13780,N_12965,N_13489);
xor U13781 (N_13781,N_13284,N_13215);
xnor U13782 (N_13782,N_13203,N_13288);
or U13783 (N_13783,N_13204,N_12893);
and U13784 (N_13784,N_13563,N_13546);
or U13785 (N_13785,N_13574,N_13154);
or U13786 (N_13786,N_13257,N_13150);
nand U13787 (N_13787,N_13454,N_13483);
and U13788 (N_13788,N_13270,N_13000);
and U13789 (N_13789,N_13305,N_13420);
and U13790 (N_13790,N_12906,N_12974);
nand U13791 (N_13791,N_12949,N_13474);
nand U13792 (N_13792,N_13541,N_13075);
xor U13793 (N_13793,N_13595,N_13583);
and U13794 (N_13794,N_13366,N_13517);
nor U13795 (N_13795,N_13452,N_13179);
nor U13796 (N_13796,N_12829,N_13584);
nand U13797 (N_13797,N_13238,N_12861);
nor U13798 (N_13798,N_13397,N_13291);
nor U13799 (N_13799,N_13239,N_12983);
nor U13800 (N_13800,N_13399,N_13287);
and U13801 (N_13801,N_13237,N_13444);
nand U13802 (N_13802,N_13547,N_13250);
nand U13803 (N_13803,N_13272,N_13455);
nand U13804 (N_13804,N_12854,N_13448);
xor U13805 (N_13805,N_13449,N_12853);
and U13806 (N_13806,N_13163,N_12896);
nand U13807 (N_13807,N_13111,N_13058);
and U13808 (N_13808,N_13450,N_12900);
or U13809 (N_13809,N_13241,N_12991);
xor U13810 (N_13810,N_13085,N_12802);
nor U13811 (N_13811,N_13030,N_13302);
xnor U13812 (N_13812,N_12805,N_12867);
nand U13813 (N_13813,N_12929,N_13289);
or U13814 (N_13814,N_13158,N_13340);
nand U13815 (N_13815,N_13538,N_13223);
nand U13816 (N_13816,N_13121,N_12882);
xor U13817 (N_13817,N_13427,N_13410);
nand U13818 (N_13818,N_13024,N_12954);
nand U13819 (N_13819,N_12876,N_13295);
xor U13820 (N_13820,N_13310,N_12909);
xnor U13821 (N_13821,N_13418,N_13227);
or U13822 (N_13822,N_13283,N_12919);
nand U13823 (N_13823,N_13079,N_12963);
nor U13824 (N_13824,N_13217,N_13370);
and U13825 (N_13825,N_13226,N_13520);
or U13826 (N_13826,N_13172,N_12986);
xor U13827 (N_13827,N_13484,N_13092);
xor U13828 (N_13828,N_13014,N_12972);
or U13829 (N_13829,N_13156,N_13225);
xor U13830 (N_13830,N_13549,N_12940);
and U13831 (N_13831,N_13136,N_12932);
and U13832 (N_13832,N_13443,N_13374);
or U13833 (N_13833,N_12935,N_13330);
xnor U13834 (N_13834,N_12894,N_12892);
and U13835 (N_13835,N_13447,N_13401);
and U13836 (N_13836,N_13183,N_13016);
and U13837 (N_13837,N_12843,N_13146);
or U13838 (N_13838,N_13462,N_13304);
nor U13839 (N_13839,N_13190,N_13317);
and U13840 (N_13840,N_13010,N_12826);
nand U13841 (N_13841,N_13337,N_13128);
and U13842 (N_13842,N_13345,N_13588);
xor U13843 (N_13843,N_13088,N_13335);
xor U13844 (N_13844,N_13012,N_12914);
and U13845 (N_13845,N_13096,N_13069);
or U13846 (N_13846,N_13144,N_13177);
nor U13847 (N_13847,N_13385,N_13569);
nand U13848 (N_13848,N_13351,N_12985);
and U13849 (N_13849,N_13050,N_13328);
and U13850 (N_13850,N_13052,N_13324);
or U13851 (N_13851,N_13364,N_13451);
xnor U13852 (N_13852,N_13570,N_13582);
xor U13853 (N_13853,N_12837,N_13540);
nor U13854 (N_13854,N_13235,N_13205);
nor U13855 (N_13855,N_12975,N_13394);
xor U13856 (N_13856,N_12815,N_13135);
and U13857 (N_13857,N_13265,N_12862);
and U13858 (N_13858,N_13184,N_13400);
and U13859 (N_13859,N_12951,N_13210);
nor U13860 (N_13860,N_13509,N_13567);
and U13861 (N_13861,N_13544,N_13194);
xnor U13862 (N_13862,N_13006,N_13545);
nor U13863 (N_13863,N_12952,N_13359);
xnor U13864 (N_13864,N_13161,N_13212);
or U13865 (N_13865,N_13511,N_13551);
and U13866 (N_13866,N_13319,N_13478);
nand U13867 (N_13867,N_13115,N_12908);
or U13868 (N_13868,N_13415,N_12823);
and U13869 (N_13869,N_13105,N_13232);
xnor U13870 (N_13870,N_12905,N_13594);
xor U13871 (N_13871,N_13098,N_13189);
nor U13872 (N_13872,N_13113,N_13441);
nor U13873 (N_13873,N_13446,N_13074);
and U13874 (N_13874,N_13375,N_13281);
nor U13875 (N_13875,N_13495,N_13083);
nand U13876 (N_13876,N_13023,N_13466);
nand U13877 (N_13877,N_13200,N_13485);
nor U13878 (N_13878,N_13219,N_13213);
and U13879 (N_13879,N_13093,N_13392);
nand U13880 (N_13880,N_13292,N_13537);
and U13881 (N_13881,N_12938,N_13059);
xnor U13882 (N_13882,N_12992,N_13022);
or U13883 (N_13883,N_13253,N_13055);
nor U13884 (N_13884,N_13334,N_13306);
xor U13885 (N_13885,N_12984,N_13066);
nor U13886 (N_13886,N_13002,N_13134);
nand U13887 (N_13887,N_13045,N_13228);
nor U13888 (N_13888,N_13125,N_13103);
nor U13889 (N_13889,N_13255,N_13579);
nor U13890 (N_13890,N_13405,N_13336);
nor U13891 (N_13891,N_13539,N_13381);
xor U13892 (N_13892,N_13361,N_13166);
nor U13893 (N_13893,N_13435,N_13104);
nand U13894 (N_13894,N_12887,N_13141);
and U13895 (N_13895,N_13503,N_13129);
or U13896 (N_13896,N_13208,N_12931);
xnor U13897 (N_13897,N_12917,N_13197);
xor U13898 (N_13898,N_13243,N_13437);
or U13899 (N_13899,N_12968,N_13047);
or U13900 (N_13900,N_13522,N_12948);
xor U13901 (N_13901,N_13460,N_13122);
or U13902 (N_13902,N_13498,N_12946);
nor U13903 (N_13903,N_12885,N_13512);
or U13904 (N_13904,N_13109,N_13142);
nand U13905 (N_13905,N_12998,N_13188);
xor U13906 (N_13906,N_13192,N_13322);
nand U13907 (N_13907,N_13060,N_12901);
nor U13908 (N_13908,N_13521,N_13274);
nand U13909 (N_13909,N_13515,N_13507);
nand U13910 (N_13910,N_12936,N_12979);
nand U13911 (N_13911,N_13329,N_12830);
nand U13912 (N_13912,N_13251,N_13112);
nor U13913 (N_13913,N_13131,N_13229);
xnor U13914 (N_13914,N_12842,N_13211);
nand U13915 (N_13915,N_13529,N_13195);
and U13916 (N_13916,N_13224,N_13490);
or U13917 (N_13917,N_12858,N_13169);
nor U13918 (N_13918,N_13300,N_13118);
xnor U13919 (N_13919,N_12847,N_12812);
and U13920 (N_13920,N_13470,N_13554);
and U13921 (N_13921,N_12957,N_12942);
xnor U13922 (N_13922,N_13497,N_13457);
or U13923 (N_13923,N_13456,N_13557);
nor U13924 (N_13924,N_13525,N_13187);
and U13925 (N_13925,N_12859,N_13296);
nor U13926 (N_13926,N_13264,N_12915);
and U13927 (N_13927,N_12980,N_13181);
nand U13928 (N_13928,N_13513,N_13519);
or U13929 (N_13929,N_13233,N_13279);
xnor U13930 (N_13930,N_12863,N_12999);
and U13931 (N_13931,N_12941,N_13496);
nor U13932 (N_13932,N_13042,N_13477);
or U13933 (N_13933,N_13209,N_12930);
nor U13934 (N_13934,N_13107,N_12947);
nand U13935 (N_13935,N_13067,N_13391);
or U13936 (N_13936,N_13314,N_13160);
nor U13937 (N_13937,N_12916,N_13508);
or U13938 (N_13938,N_13221,N_12881);
nor U13939 (N_13939,N_13542,N_13029);
or U13940 (N_13940,N_13186,N_13419);
nand U13941 (N_13941,N_12873,N_13442);
nand U13942 (N_13942,N_13350,N_13559);
and U13943 (N_13943,N_13311,N_12943);
and U13944 (N_13944,N_12996,N_13577);
xor U13945 (N_13945,N_13261,N_13077);
and U13946 (N_13946,N_13440,N_13403);
xnor U13947 (N_13947,N_12969,N_13424);
nand U13948 (N_13948,N_13348,N_13094);
nand U13949 (N_13949,N_13044,N_13372);
xor U13950 (N_13950,N_12976,N_13378);
nor U13951 (N_13951,N_13383,N_12898);
xor U13952 (N_13952,N_13007,N_13472);
and U13953 (N_13953,N_13556,N_13552);
nand U13954 (N_13954,N_13198,N_13254);
nand U13955 (N_13955,N_13506,N_13501);
and U13956 (N_13956,N_13001,N_12981);
nor U13957 (N_13957,N_13430,N_13318);
nand U13958 (N_13958,N_13081,N_13256);
nand U13959 (N_13959,N_12899,N_12978);
and U13960 (N_13960,N_13145,N_13080);
nand U13961 (N_13961,N_13467,N_13157);
nand U13962 (N_13962,N_13293,N_12897);
nand U13963 (N_13963,N_12890,N_13404);
nor U13964 (N_13964,N_12961,N_13414);
xor U13965 (N_13965,N_13307,N_13581);
xnor U13966 (N_13966,N_13422,N_13367);
or U13967 (N_13967,N_13167,N_12818);
xnor U13968 (N_13968,N_12851,N_13586);
xor U13969 (N_13969,N_13218,N_13064);
nor U13970 (N_13970,N_13475,N_13480);
nand U13971 (N_13971,N_12800,N_12849);
or U13972 (N_13972,N_12895,N_13376);
and U13973 (N_13973,N_12958,N_12833);
nor U13974 (N_13974,N_13137,N_13358);
and U13975 (N_13975,N_13516,N_12880);
nor U13976 (N_13976,N_13119,N_13325);
nor U13977 (N_13977,N_12846,N_13338);
or U13978 (N_13978,N_13377,N_13368);
or U13979 (N_13979,N_12884,N_13216);
and U13980 (N_13980,N_13051,N_13326);
xnor U13981 (N_13981,N_13280,N_13040);
xor U13982 (N_13982,N_13017,N_13297);
xnor U13983 (N_13983,N_13076,N_13222);
xor U13984 (N_13984,N_13191,N_12995);
or U13985 (N_13985,N_12879,N_12822);
xor U13986 (N_13986,N_12803,N_13303);
xor U13987 (N_13987,N_12920,N_13110);
nand U13988 (N_13988,N_13041,N_13285);
and U13989 (N_13989,N_12982,N_13327);
nor U13990 (N_13990,N_12801,N_13491);
and U13991 (N_13991,N_13486,N_13453);
xnor U13992 (N_13992,N_12871,N_13439);
nor U13993 (N_13993,N_12907,N_13380);
nor U13994 (N_13994,N_12804,N_12877);
or U13995 (N_13995,N_13126,N_13031);
or U13996 (N_13996,N_13267,N_12977);
nand U13997 (N_13997,N_13488,N_13568);
and U13998 (N_13998,N_13365,N_13548);
nor U13999 (N_13999,N_13406,N_13429);
and U14000 (N_14000,N_13446,N_13096);
or U14001 (N_14001,N_13073,N_13050);
nand U14002 (N_14002,N_12858,N_13321);
xor U14003 (N_14003,N_13525,N_12960);
and U14004 (N_14004,N_13021,N_13427);
xor U14005 (N_14005,N_13194,N_13376);
xnor U14006 (N_14006,N_13599,N_13497);
and U14007 (N_14007,N_13185,N_13490);
or U14008 (N_14008,N_13478,N_12977);
nand U14009 (N_14009,N_13543,N_13300);
or U14010 (N_14010,N_13505,N_12851);
xor U14011 (N_14011,N_13071,N_13074);
nor U14012 (N_14012,N_13207,N_13485);
nor U14013 (N_14013,N_13580,N_13053);
nand U14014 (N_14014,N_13276,N_12813);
xnor U14015 (N_14015,N_13369,N_12982);
or U14016 (N_14016,N_13421,N_13179);
nor U14017 (N_14017,N_13502,N_13545);
nor U14018 (N_14018,N_13492,N_13425);
and U14019 (N_14019,N_13592,N_13144);
xnor U14020 (N_14020,N_13401,N_12820);
and U14021 (N_14021,N_13380,N_13401);
nand U14022 (N_14022,N_13176,N_13122);
or U14023 (N_14023,N_13369,N_12999);
nand U14024 (N_14024,N_13597,N_13023);
and U14025 (N_14025,N_13520,N_12949);
and U14026 (N_14026,N_13210,N_13599);
and U14027 (N_14027,N_13569,N_13193);
or U14028 (N_14028,N_13230,N_13380);
and U14029 (N_14029,N_13335,N_13343);
xor U14030 (N_14030,N_13499,N_13415);
or U14031 (N_14031,N_13361,N_12853);
xor U14032 (N_14032,N_13362,N_13439);
or U14033 (N_14033,N_13009,N_12861);
and U14034 (N_14034,N_13340,N_13330);
xor U14035 (N_14035,N_13552,N_13588);
nor U14036 (N_14036,N_12829,N_13137);
nor U14037 (N_14037,N_13267,N_12872);
nand U14038 (N_14038,N_13402,N_12808);
nand U14039 (N_14039,N_13430,N_13247);
nor U14040 (N_14040,N_12891,N_13386);
xnor U14041 (N_14041,N_13423,N_13474);
nor U14042 (N_14042,N_13532,N_13094);
xnor U14043 (N_14043,N_12926,N_13164);
nor U14044 (N_14044,N_13078,N_13117);
or U14045 (N_14045,N_13458,N_13235);
and U14046 (N_14046,N_13023,N_13109);
nor U14047 (N_14047,N_13199,N_13524);
nand U14048 (N_14048,N_13241,N_13035);
and U14049 (N_14049,N_13496,N_13131);
nor U14050 (N_14050,N_13078,N_13129);
nor U14051 (N_14051,N_13117,N_13502);
nor U14052 (N_14052,N_13252,N_13542);
and U14053 (N_14053,N_13284,N_13026);
nand U14054 (N_14054,N_13533,N_13109);
nor U14055 (N_14055,N_12889,N_13252);
nor U14056 (N_14056,N_13405,N_13249);
xnor U14057 (N_14057,N_13467,N_13381);
or U14058 (N_14058,N_12870,N_13142);
nor U14059 (N_14059,N_13580,N_12952);
xnor U14060 (N_14060,N_13514,N_13032);
nor U14061 (N_14061,N_13599,N_12940);
or U14062 (N_14062,N_13120,N_13035);
or U14063 (N_14063,N_12888,N_13516);
nor U14064 (N_14064,N_13579,N_13502);
and U14065 (N_14065,N_13115,N_13257);
nand U14066 (N_14066,N_13524,N_13010);
xor U14067 (N_14067,N_12827,N_13158);
or U14068 (N_14068,N_12825,N_12935);
xor U14069 (N_14069,N_13130,N_13380);
or U14070 (N_14070,N_13008,N_13275);
nand U14071 (N_14071,N_13250,N_13536);
nand U14072 (N_14072,N_13192,N_13489);
or U14073 (N_14073,N_13193,N_13147);
nor U14074 (N_14074,N_13265,N_12935);
or U14075 (N_14075,N_13245,N_13384);
nand U14076 (N_14076,N_13015,N_13067);
or U14077 (N_14077,N_12940,N_13504);
xor U14078 (N_14078,N_13220,N_13209);
xor U14079 (N_14079,N_13172,N_13221);
xor U14080 (N_14080,N_13233,N_13535);
nor U14081 (N_14081,N_13130,N_13563);
nand U14082 (N_14082,N_12946,N_13332);
nand U14083 (N_14083,N_13241,N_12888);
and U14084 (N_14084,N_12909,N_12980);
or U14085 (N_14085,N_12989,N_13111);
nor U14086 (N_14086,N_12966,N_12879);
and U14087 (N_14087,N_13395,N_12802);
or U14088 (N_14088,N_13594,N_13263);
nand U14089 (N_14089,N_12990,N_13255);
or U14090 (N_14090,N_13543,N_13202);
xnor U14091 (N_14091,N_13474,N_13490);
xor U14092 (N_14092,N_13268,N_13176);
nand U14093 (N_14093,N_13251,N_13475);
xnor U14094 (N_14094,N_13428,N_13093);
and U14095 (N_14095,N_13101,N_12843);
and U14096 (N_14096,N_12995,N_13249);
xor U14097 (N_14097,N_13021,N_13181);
nand U14098 (N_14098,N_13234,N_12808);
xnor U14099 (N_14099,N_13430,N_13272);
xnor U14100 (N_14100,N_13225,N_13502);
nor U14101 (N_14101,N_13064,N_12884);
nor U14102 (N_14102,N_13229,N_13111);
nor U14103 (N_14103,N_13227,N_13365);
xor U14104 (N_14104,N_12953,N_13187);
nor U14105 (N_14105,N_13454,N_13221);
or U14106 (N_14106,N_13526,N_13019);
nor U14107 (N_14107,N_12943,N_13078);
xor U14108 (N_14108,N_13323,N_13226);
nor U14109 (N_14109,N_13348,N_13066);
xor U14110 (N_14110,N_13398,N_13181);
xnor U14111 (N_14111,N_13257,N_12890);
nand U14112 (N_14112,N_12864,N_13022);
nand U14113 (N_14113,N_12933,N_13536);
nand U14114 (N_14114,N_13342,N_12844);
or U14115 (N_14115,N_12883,N_13334);
or U14116 (N_14116,N_13513,N_13023);
or U14117 (N_14117,N_13145,N_12898);
xor U14118 (N_14118,N_13417,N_12900);
nand U14119 (N_14119,N_13142,N_13554);
or U14120 (N_14120,N_13260,N_13174);
xnor U14121 (N_14121,N_13434,N_13238);
nand U14122 (N_14122,N_12935,N_12880);
and U14123 (N_14123,N_13535,N_12828);
xnor U14124 (N_14124,N_12920,N_13199);
nand U14125 (N_14125,N_13368,N_13125);
or U14126 (N_14126,N_13453,N_12895);
and U14127 (N_14127,N_13557,N_13014);
or U14128 (N_14128,N_13391,N_13249);
and U14129 (N_14129,N_12974,N_12932);
and U14130 (N_14130,N_13549,N_12933);
and U14131 (N_14131,N_13403,N_13328);
and U14132 (N_14132,N_13413,N_12801);
or U14133 (N_14133,N_12829,N_12851);
nand U14134 (N_14134,N_12828,N_13339);
nand U14135 (N_14135,N_13452,N_13059);
and U14136 (N_14136,N_13331,N_13476);
xor U14137 (N_14137,N_13032,N_13416);
and U14138 (N_14138,N_13432,N_13256);
nor U14139 (N_14139,N_13014,N_13225);
and U14140 (N_14140,N_13091,N_13304);
nand U14141 (N_14141,N_12983,N_12929);
nor U14142 (N_14142,N_13522,N_13083);
nand U14143 (N_14143,N_13589,N_12936);
or U14144 (N_14144,N_13013,N_13257);
and U14145 (N_14145,N_13414,N_13532);
nand U14146 (N_14146,N_13426,N_13573);
or U14147 (N_14147,N_13039,N_13582);
or U14148 (N_14148,N_13200,N_13441);
nor U14149 (N_14149,N_13103,N_13023);
and U14150 (N_14150,N_13024,N_12888);
and U14151 (N_14151,N_13092,N_13426);
and U14152 (N_14152,N_13313,N_13591);
and U14153 (N_14153,N_13312,N_13242);
nand U14154 (N_14154,N_13268,N_13513);
and U14155 (N_14155,N_13511,N_12822);
or U14156 (N_14156,N_12802,N_12830);
and U14157 (N_14157,N_13323,N_13387);
and U14158 (N_14158,N_13133,N_13432);
nand U14159 (N_14159,N_13002,N_13351);
xor U14160 (N_14160,N_13094,N_13245);
nand U14161 (N_14161,N_12992,N_13119);
and U14162 (N_14162,N_12990,N_13586);
xor U14163 (N_14163,N_13178,N_13268);
xor U14164 (N_14164,N_13579,N_13098);
and U14165 (N_14165,N_12818,N_13338);
nand U14166 (N_14166,N_13218,N_13388);
and U14167 (N_14167,N_13238,N_13330);
nand U14168 (N_14168,N_13374,N_13174);
xor U14169 (N_14169,N_13087,N_13399);
nand U14170 (N_14170,N_13294,N_13512);
xor U14171 (N_14171,N_13094,N_12916);
and U14172 (N_14172,N_13140,N_12897);
nor U14173 (N_14173,N_13379,N_12995);
and U14174 (N_14174,N_13190,N_13279);
nand U14175 (N_14175,N_13512,N_12840);
nor U14176 (N_14176,N_13069,N_13478);
nand U14177 (N_14177,N_13466,N_13520);
nor U14178 (N_14178,N_12966,N_12834);
nor U14179 (N_14179,N_12894,N_13506);
or U14180 (N_14180,N_13173,N_12841);
and U14181 (N_14181,N_12999,N_13142);
or U14182 (N_14182,N_13175,N_12948);
or U14183 (N_14183,N_12945,N_13126);
nand U14184 (N_14184,N_12850,N_13350);
or U14185 (N_14185,N_13214,N_12931);
and U14186 (N_14186,N_13589,N_13168);
nor U14187 (N_14187,N_12929,N_13506);
xor U14188 (N_14188,N_13403,N_13485);
xnor U14189 (N_14189,N_12957,N_13498);
or U14190 (N_14190,N_13171,N_13246);
or U14191 (N_14191,N_13260,N_12914);
nor U14192 (N_14192,N_13340,N_13021);
and U14193 (N_14193,N_13056,N_13524);
xnor U14194 (N_14194,N_13068,N_13558);
nor U14195 (N_14195,N_13496,N_13022);
xnor U14196 (N_14196,N_13122,N_13107);
nand U14197 (N_14197,N_13241,N_12839);
nor U14198 (N_14198,N_13335,N_13406);
or U14199 (N_14199,N_13339,N_12975);
and U14200 (N_14200,N_13092,N_12902);
nor U14201 (N_14201,N_13029,N_13173);
and U14202 (N_14202,N_13510,N_13042);
and U14203 (N_14203,N_13357,N_13502);
nor U14204 (N_14204,N_12820,N_13142);
or U14205 (N_14205,N_13362,N_13453);
or U14206 (N_14206,N_13497,N_13229);
xnor U14207 (N_14207,N_13395,N_13451);
or U14208 (N_14208,N_12979,N_13268);
xor U14209 (N_14209,N_13121,N_13140);
nand U14210 (N_14210,N_12841,N_13106);
or U14211 (N_14211,N_13398,N_13517);
nand U14212 (N_14212,N_13278,N_13480);
and U14213 (N_14213,N_13346,N_12817);
xor U14214 (N_14214,N_13001,N_13539);
and U14215 (N_14215,N_12989,N_13445);
nor U14216 (N_14216,N_13466,N_12940);
nand U14217 (N_14217,N_13537,N_13403);
xor U14218 (N_14218,N_13538,N_13286);
and U14219 (N_14219,N_13251,N_13592);
or U14220 (N_14220,N_12874,N_13409);
xor U14221 (N_14221,N_13441,N_13510);
or U14222 (N_14222,N_13558,N_13368);
nor U14223 (N_14223,N_13438,N_12975);
nand U14224 (N_14224,N_13047,N_13012);
xor U14225 (N_14225,N_13182,N_13383);
or U14226 (N_14226,N_12887,N_13257);
nor U14227 (N_14227,N_13257,N_13468);
nand U14228 (N_14228,N_13440,N_13375);
nand U14229 (N_14229,N_13040,N_13520);
nand U14230 (N_14230,N_13336,N_13442);
and U14231 (N_14231,N_12839,N_13256);
nand U14232 (N_14232,N_13571,N_12806);
or U14233 (N_14233,N_13436,N_13068);
and U14234 (N_14234,N_13120,N_13107);
and U14235 (N_14235,N_13441,N_13571);
or U14236 (N_14236,N_13263,N_13488);
nand U14237 (N_14237,N_12873,N_13444);
xnor U14238 (N_14238,N_12847,N_13296);
and U14239 (N_14239,N_13114,N_13150);
xor U14240 (N_14240,N_13175,N_13065);
nand U14241 (N_14241,N_13080,N_12844);
nand U14242 (N_14242,N_13420,N_13535);
and U14243 (N_14243,N_13202,N_12806);
or U14244 (N_14244,N_13431,N_13307);
nand U14245 (N_14245,N_13386,N_13102);
nand U14246 (N_14246,N_13453,N_13372);
and U14247 (N_14247,N_13007,N_12809);
or U14248 (N_14248,N_13505,N_13178);
xnor U14249 (N_14249,N_13344,N_13560);
and U14250 (N_14250,N_13238,N_12852);
xnor U14251 (N_14251,N_12825,N_12801);
or U14252 (N_14252,N_13081,N_13563);
or U14253 (N_14253,N_13361,N_13373);
and U14254 (N_14254,N_12906,N_12872);
and U14255 (N_14255,N_12878,N_13059);
xor U14256 (N_14256,N_13153,N_13269);
or U14257 (N_14257,N_13158,N_13184);
xor U14258 (N_14258,N_13293,N_13578);
nand U14259 (N_14259,N_13241,N_13491);
nor U14260 (N_14260,N_12991,N_13516);
or U14261 (N_14261,N_13448,N_12859);
nand U14262 (N_14262,N_12964,N_12984);
and U14263 (N_14263,N_13459,N_12972);
xor U14264 (N_14264,N_12811,N_12859);
or U14265 (N_14265,N_13583,N_13239);
nand U14266 (N_14266,N_12977,N_13349);
xnor U14267 (N_14267,N_12912,N_13264);
nand U14268 (N_14268,N_13041,N_12901);
nand U14269 (N_14269,N_13154,N_12978);
xnor U14270 (N_14270,N_12980,N_13164);
nand U14271 (N_14271,N_13425,N_13350);
xor U14272 (N_14272,N_13026,N_13203);
and U14273 (N_14273,N_12999,N_13160);
nor U14274 (N_14274,N_13396,N_12866);
and U14275 (N_14275,N_13475,N_13338);
nor U14276 (N_14276,N_13232,N_12896);
nand U14277 (N_14277,N_13193,N_12851);
or U14278 (N_14278,N_12915,N_13351);
and U14279 (N_14279,N_13550,N_12826);
xnor U14280 (N_14280,N_13174,N_13469);
and U14281 (N_14281,N_13132,N_13492);
nand U14282 (N_14282,N_13301,N_12878);
xnor U14283 (N_14283,N_13048,N_13018);
or U14284 (N_14284,N_13186,N_13179);
xnor U14285 (N_14285,N_13097,N_13149);
xor U14286 (N_14286,N_13365,N_12984);
nor U14287 (N_14287,N_12928,N_13514);
or U14288 (N_14288,N_12907,N_12901);
and U14289 (N_14289,N_13072,N_13094);
nor U14290 (N_14290,N_13027,N_12952);
or U14291 (N_14291,N_12967,N_12972);
and U14292 (N_14292,N_12852,N_13159);
or U14293 (N_14293,N_12805,N_13468);
and U14294 (N_14294,N_13158,N_13051);
nand U14295 (N_14295,N_13249,N_13264);
and U14296 (N_14296,N_12938,N_13036);
or U14297 (N_14297,N_13118,N_12826);
nor U14298 (N_14298,N_12908,N_12861);
nor U14299 (N_14299,N_13114,N_13512);
xor U14300 (N_14300,N_12956,N_13575);
xor U14301 (N_14301,N_12961,N_13330);
and U14302 (N_14302,N_13260,N_13249);
xor U14303 (N_14303,N_13160,N_13504);
or U14304 (N_14304,N_13570,N_13071);
xor U14305 (N_14305,N_13461,N_13055);
or U14306 (N_14306,N_13203,N_13445);
nor U14307 (N_14307,N_13497,N_13458);
xnor U14308 (N_14308,N_13017,N_12803);
nand U14309 (N_14309,N_13405,N_13026);
xnor U14310 (N_14310,N_13330,N_13203);
and U14311 (N_14311,N_12887,N_12822);
nor U14312 (N_14312,N_13397,N_13466);
nor U14313 (N_14313,N_12884,N_13418);
nand U14314 (N_14314,N_13599,N_12988);
xor U14315 (N_14315,N_13229,N_13583);
or U14316 (N_14316,N_13262,N_13281);
or U14317 (N_14317,N_12998,N_13495);
nand U14318 (N_14318,N_13186,N_13159);
or U14319 (N_14319,N_13394,N_13090);
nand U14320 (N_14320,N_13415,N_13565);
nor U14321 (N_14321,N_13004,N_13431);
nand U14322 (N_14322,N_12853,N_13483);
or U14323 (N_14323,N_13365,N_13045);
nor U14324 (N_14324,N_13306,N_13038);
or U14325 (N_14325,N_13035,N_12994);
or U14326 (N_14326,N_12940,N_13570);
nand U14327 (N_14327,N_13104,N_12842);
nand U14328 (N_14328,N_12944,N_13282);
nand U14329 (N_14329,N_13504,N_12992);
or U14330 (N_14330,N_13446,N_13515);
and U14331 (N_14331,N_13021,N_13419);
and U14332 (N_14332,N_13454,N_13351);
and U14333 (N_14333,N_13126,N_13146);
xor U14334 (N_14334,N_13037,N_13462);
or U14335 (N_14335,N_13436,N_13553);
nor U14336 (N_14336,N_13440,N_13284);
xor U14337 (N_14337,N_13482,N_13248);
nor U14338 (N_14338,N_13405,N_13247);
nor U14339 (N_14339,N_13428,N_13510);
nand U14340 (N_14340,N_13483,N_13035);
nand U14341 (N_14341,N_13272,N_13102);
xor U14342 (N_14342,N_13341,N_13058);
nor U14343 (N_14343,N_13103,N_13187);
xor U14344 (N_14344,N_13445,N_12894);
or U14345 (N_14345,N_12966,N_12946);
or U14346 (N_14346,N_13444,N_13535);
nand U14347 (N_14347,N_13014,N_13422);
nand U14348 (N_14348,N_13576,N_13434);
nor U14349 (N_14349,N_13206,N_13244);
nand U14350 (N_14350,N_13198,N_13331);
or U14351 (N_14351,N_13155,N_13203);
nand U14352 (N_14352,N_12852,N_13410);
nor U14353 (N_14353,N_13075,N_12927);
and U14354 (N_14354,N_13248,N_13013);
and U14355 (N_14355,N_13552,N_13520);
nor U14356 (N_14356,N_13059,N_13583);
xor U14357 (N_14357,N_13192,N_13295);
nand U14358 (N_14358,N_12839,N_13195);
and U14359 (N_14359,N_13132,N_12818);
xor U14360 (N_14360,N_13277,N_13079);
or U14361 (N_14361,N_13022,N_13307);
or U14362 (N_14362,N_12977,N_13414);
nand U14363 (N_14363,N_13437,N_13072);
nor U14364 (N_14364,N_12975,N_13460);
or U14365 (N_14365,N_13076,N_13449);
nor U14366 (N_14366,N_13472,N_13335);
nor U14367 (N_14367,N_13087,N_13227);
or U14368 (N_14368,N_13320,N_13375);
nor U14369 (N_14369,N_13414,N_13503);
or U14370 (N_14370,N_13285,N_13457);
xor U14371 (N_14371,N_13509,N_12805);
or U14372 (N_14372,N_13569,N_13202);
xnor U14373 (N_14373,N_12851,N_12929);
or U14374 (N_14374,N_12843,N_13369);
and U14375 (N_14375,N_13470,N_13109);
xor U14376 (N_14376,N_13498,N_13479);
nor U14377 (N_14377,N_12842,N_13129);
and U14378 (N_14378,N_12879,N_13089);
xor U14379 (N_14379,N_13130,N_13150);
or U14380 (N_14380,N_13369,N_13352);
xor U14381 (N_14381,N_12884,N_13447);
xnor U14382 (N_14382,N_12981,N_12959);
nor U14383 (N_14383,N_12995,N_12852);
nor U14384 (N_14384,N_12887,N_13210);
xnor U14385 (N_14385,N_13455,N_12908);
or U14386 (N_14386,N_13393,N_13461);
nand U14387 (N_14387,N_13042,N_13490);
and U14388 (N_14388,N_13072,N_13218);
or U14389 (N_14389,N_13346,N_13226);
xnor U14390 (N_14390,N_13399,N_13168);
or U14391 (N_14391,N_13314,N_13460);
nor U14392 (N_14392,N_13093,N_12921);
nor U14393 (N_14393,N_13551,N_12866);
or U14394 (N_14394,N_13118,N_13424);
xnor U14395 (N_14395,N_13010,N_12983);
nand U14396 (N_14396,N_13386,N_12911);
nand U14397 (N_14397,N_13120,N_12954);
nand U14398 (N_14398,N_13570,N_13294);
or U14399 (N_14399,N_13382,N_13364);
and U14400 (N_14400,N_13608,N_14080);
xnor U14401 (N_14401,N_13701,N_13823);
xnor U14402 (N_14402,N_14102,N_13687);
or U14403 (N_14403,N_13861,N_14327);
nor U14404 (N_14404,N_13659,N_13621);
nor U14405 (N_14405,N_14017,N_14346);
and U14406 (N_14406,N_14030,N_13658);
xnor U14407 (N_14407,N_13824,N_13997);
and U14408 (N_14408,N_14399,N_14397);
and U14409 (N_14409,N_14147,N_14103);
nand U14410 (N_14410,N_13698,N_14288);
nor U14411 (N_14411,N_14013,N_14055);
or U14412 (N_14412,N_13994,N_14201);
and U14413 (N_14413,N_13802,N_14333);
and U14414 (N_14414,N_13919,N_13875);
xor U14415 (N_14415,N_13971,N_14348);
nand U14416 (N_14416,N_14294,N_13893);
and U14417 (N_14417,N_13848,N_14139);
nor U14418 (N_14418,N_13764,N_14140);
xor U14419 (N_14419,N_14276,N_14023);
nor U14420 (N_14420,N_14290,N_14190);
or U14421 (N_14421,N_13776,N_13839);
and U14422 (N_14422,N_13882,N_13617);
nand U14423 (N_14423,N_13863,N_13881);
and U14424 (N_14424,N_13601,N_13954);
or U14425 (N_14425,N_13715,N_13744);
nor U14426 (N_14426,N_13970,N_14071);
nand U14427 (N_14427,N_13772,N_13936);
or U14428 (N_14428,N_13792,N_13725);
nand U14429 (N_14429,N_13998,N_14186);
xor U14430 (N_14430,N_14090,N_14221);
xnor U14431 (N_14431,N_13800,N_14217);
nor U14432 (N_14432,N_14143,N_14001);
or U14433 (N_14433,N_13742,N_14029);
and U14434 (N_14434,N_13728,N_14342);
or U14435 (N_14435,N_13915,N_13610);
nand U14436 (N_14436,N_13736,N_14255);
nor U14437 (N_14437,N_14341,N_13921);
xnor U14438 (N_14438,N_13969,N_13688);
nand U14439 (N_14439,N_14265,N_14301);
or U14440 (N_14440,N_13706,N_13778);
or U14441 (N_14441,N_13837,N_13850);
and U14442 (N_14442,N_14227,N_13884);
or U14443 (N_14443,N_14195,N_13849);
nor U14444 (N_14444,N_14137,N_14353);
and U14445 (N_14445,N_14377,N_13633);
xor U14446 (N_14446,N_14376,N_14228);
or U14447 (N_14447,N_14066,N_14150);
and U14448 (N_14448,N_14157,N_13791);
nor U14449 (N_14449,N_13755,N_14014);
and U14450 (N_14450,N_14188,N_13923);
nor U14451 (N_14451,N_14329,N_14165);
nand U14452 (N_14452,N_13825,N_14061);
or U14453 (N_14453,N_14269,N_13991);
and U14454 (N_14454,N_14254,N_13628);
or U14455 (N_14455,N_14105,N_14101);
xor U14456 (N_14456,N_13751,N_14088);
nand U14457 (N_14457,N_14126,N_14379);
nor U14458 (N_14458,N_14374,N_14251);
nand U14459 (N_14459,N_13827,N_13868);
xnor U14460 (N_14460,N_14096,N_13932);
nor U14461 (N_14461,N_13902,N_14002);
or U14462 (N_14462,N_14205,N_14142);
and U14463 (N_14463,N_13950,N_14378);
and U14464 (N_14464,N_13714,N_14282);
nor U14465 (N_14465,N_13908,N_13762);
and U14466 (N_14466,N_13870,N_13815);
xor U14467 (N_14467,N_14020,N_14077);
xnor U14468 (N_14468,N_14039,N_13880);
nor U14469 (N_14469,N_13724,N_14218);
xor U14470 (N_14470,N_13966,N_14056);
or U14471 (N_14471,N_14193,N_13841);
nand U14472 (N_14472,N_13903,N_13780);
nand U14473 (N_14473,N_14177,N_14166);
or U14474 (N_14474,N_14115,N_14111);
nand U14475 (N_14475,N_14344,N_13912);
nor U14476 (N_14476,N_13968,N_14054);
nor U14477 (N_14477,N_14268,N_14160);
nor U14478 (N_14478,N_13729,N_13924);
and U14479 (N_14479,N_14113,N_14075);
nand U14480 (N_14480,N_13851,N_14280);
and U14481 (N_14481,N_14381,N_14152);
and U14482 (N_14482,N_14073,N_14295);
nand U14483 (N_14483,N_13951,N_13809);
nand U14484 (N_14484,N_14220,N_13944);
or U14485 (N_14485,N_14035,N_14311);
or U14486 (N_14486,N_13948,N_14314);
or U14487 (N_14487,N_13874,N_13620);
nand U14488 (N_14488,N_13907,N_13666);
nor U14489 (N_14489,N_14273,N_14128);
nor U14490 (N_14490,N_13883,N_13734);
nand U14491 (N_14491,N_13747,N_14340);
xnor U14492 (N_14492,N_13675,N_13856);
and U14493 (N_14493,N_13929,N_13726);
nor U14494 (N_14494,N_14212,N_14230);
nor U14495 (N_14495,N_13871,N_13731);
and U14496 (N_14496,N_13935,N_13739);
nand U14497 (N_14497,N_13808,N_13749);
xor U14498 (N_14498,N_13964,N_14312);
nor U14499 (N_14499,N_13829,N_13679);
nor U14500 (N_14500,N_13822,N_14242);
nor U14501 (N_14501,N_13836,N_13672);
nand U14502 (N_14502,N_14367,N_13801);
nand U14503 (N_14503,N_14070,N_13619);
or U14504 (N_14504,N_14004,N_13989);
xnor U14505 (N_14505,N_13959,N_14026);
or U14506 (N_14506,N_13806,N_14097);
or U14507 (N_14507,N_14027,N_13980);
and U14508 (N_14508,N_13978,N_13866);
nand U14509 (N_14509,N_13766,N_13899);
xnor U14510 (N_14510,N_14326,N_14145);
xor U14511 (N_14511,N_14369,N_13697);
xor U14512 (N_14512,N_13773,N_14279);
nand U14513 (N_14513,N_14125,N_13993);
or U14514 (N_14514,N_13926,N_13692);
and U14515 (N_14515,N_13770,N_13631);
or U14516 (N_14516,N_14007,N_14064);
nand U14517 (N_14517,N_13663,N_13888);
xnor U14518 (N_14518,N_13995,N_13833);
nor U14519 (N_14519,N_13654,N_14078);
nor U14520 (N_14520,N_13717,N_13661);
nand U14521 (N_14521,N_13757,N_13947);
nand U14522 (N_14522,N_14345,N_13957);
nand U14523 (N_14523,N_14386,N_14383);
or U14524 (N_14524,N_13600,N_14296);
xnor U14525 (N_14525,N_14133,N_14068);
xnor U14526 (N_14526,N_14196,N_13955);
or U14527 (N_14527,N_13605,N_14094);
xor U14528 (N_14528,N_14175,N_13958);
and U14529 (N_14529,N_13974,N_14163);
or U14530 (N_14530,N_14063,N_13913);
or U14531 (N_14531,N_14391,N_14363);
nand U14532 (N_14532,N_13961,N_13612);
or U14533 (N_14533,N_13816,N_13844);
nand U14534 (N_14534,N_14236,N_14049);
nand U14535 (N_14535,N_13615,N_14176);
xor U14536 (N_14536,N_14067,N_14325);
nor U14537 (N_14537,N_14098,N_14283);
nor U14538 (N_14538,N_13603,N_13695);
nor U14539 (N_14539,N_13665,N_13673);
xor U14540 (N_14540,N_13650,N_14112);
nor U14541 (N_14541,N_14100,N_13982);
nor U14542 (N_14542,N_13738,N_13669);
nand U14543 (N_14543,N_14322,N_13604);
or U14544 (N_14544,N_13639,N_14202);
or U14545 (N_14545,N_13842,N_14006);
nand U14546 (N_14546,N_13645,N_14321);
and U14547 (N_14547,N_14046,N_14167);
and U14548 (N_14548,N_13803,N_14123);
nand U14549 (N_14549,N_14239,N_14134);
and U14550 (N_14550,N_14349,N_14079);
or U14551 (N_14551,N_13775,N_14306);
nand U14552 (N_14552,N_14108,N_13740);
xnor U14553 (N_14553,N_14159,N_14260);
nand U14554 (N_14554,N_14339,N_13684);
or U14555 (N_14555,N_13756,N_13693);
nand U14556 (N_14556,N_14118,N_14084);
and U14557 (N_14557,N_14315,N_13664);
nand U14558 (N_14558,N_14174,N_14398);
or U14559 (N_14559,N_14074,N_14267);
nor U14560 (N_14560,N_13973,N_14060);
and U14561 (N_14561,N_14194,N_14008);
nand U14562 (N_14562,N_14036,N_13840);
nand U14563 (N_14563,N_14215,N_14203);
and U14564 (N_14564,N_14278,N_14204);
nor U14565 (N_14565,N_14132,N_14182);
and U14566 (N_14566,N_13834,N_14146);
xor U14567 (N_14567,N_14237,N_14121);
xor U14568 (N_14568,N_14323,N_13753);
xor U14569 (N_14569,N_13911,N_13644);
nand U14570 (N_14570,N_14024,N_13767);
nand U14571 (N_14571,N_14360,N_14253);
or U14572 (N_14572,N_14387,N_13723);
or U14573 (N_14573,N_13709,N_13641);
nor U14574 (N_14574,N_14081,N_13676);
nor U14575 (N_14575,N_14334,N_13795);
and U14576 (N_14576,N_13683,N_13838);
xnor U14577 (N_14577,N_14178,N_14395);
nand U14578 (N_14578,N_14200,N_14037);
nor U14579 (N_14579,N_13820,N_13777);
or U14580 (N_14580,N_14375,N_13930);
nor U14581 (N_14581,N_13831,N_14168);
or U14582 (N_14582,N_14116,N_13963);
nor U14583 (N_14583,N_13981,N_14258);
and U14584 (N_14584,N_13745,N_14138);
xor U14585 (N_14585,N_14235,N_13647);
nor U14586 (N_14586,N_14244,N_14241);
nor U14587 (N_14587,N_13784,N_13771);
nor U14588 (N_14588,N_14358,N_14292);
or U14589 (N_14589,N_13962,N_14148);
xnor U14590 (N_14590,N_14038,N_14209);
nor U14591 (N_14591,N_13832,N_13638);
or U14592 (N_14592,N_14033,N_13786);
xor U14593 (N_14593,N_13797,N_13805);
nor U14594 (N_14594,N_14328,N_14277);
xor U14595 (N_14595,N_13854,N_13889);
xor U14596 (N_14596,N_14124,N_13873);
and U14597 (N_14597,N_13678,N_13886);
and U14598 (N_14598,N_14337,N_13732);
and U14599 (N_14599,N_13922,N_13652);
and U14600 (N_14600,N_13960,N_14156);
nor U14601 (N_14601,N_13904,N_13626);
xnor U14602 (N_14602,N_14214,N_13790);
or U14603 (N_14603,N_14229,N_13914);
or U14604 (N_14604,N_14319,N_14380);
nor U14605 (N_14605,N_13804,N_14104);
nor U14606 (N_14606,N_14048,N_14274);
xor U14607 (N_14607,N_14366,N_13972);
or U14608 (N_14608,N_13928,N_14361);
and U14609 (N_14609,N_14044,N_14347);
nand U14610 (N_14610,N_13779,N_13716);
and U14611 (N_14611,N_13986,N_13872);
and U14612 (N_14612,N_14305,N_13817);
or U14613 (N_14613,N_13819,N_13690);
or U14614 (N_14614,N_13763,N_14117);
xor U14615 (N_14615,N_14021,N_13789);
or U14616 (N_14616,N_13668,N_14372);
and U14617 (N_14617,N_13656,N_14354);
nand U14618 (N_14618,N_14370,N_13651);
nor U14619 (N_14619,N_13794,N_13918);
nor U14620 (N_14620,N_14385,N_13705);
nor U14621 (N_14621,N_13761,N_14318);
or U14622 (N_14622,N_14371,N_14316);
or U14623 (N_14623,N_13905,N_14181);
xnor U14624 (N_14624,N_13746,N_13938);
nand U14625 (N_14625,N_14216,N_13774);
xor U14626 (N_14626,N_13999,N_13718);
and U14627 (N_14627,N_13941,N_14155);
xor U14628 (N_14628,N_14382,N_14083);
nand U14629 (N_14629,N_14261,N_13892);
and U14630 (N_14630,N_14362,N_13703);
xor U14631 (N_14631,N_13879,N_13934);
or U14632 (N_14632,N_14271,N_13636);
nor U14633 (N_14633,N_13632,N_13634);
nor U14634 (N_14634,N_14106,N_13818);
xnor U14635 (N_14635,N_13783,N_13735);
xor U14636 (N_14636,N_13689,N_13845);
nand U14637 (N_14637,N_14234,N_13758);
nor U14638 (N_14638,N_14313,N_14355);
nand U14639 (N_14639,N_14359,N_13616);
nand U14640 (N_14640,N_13864,N_13956);
and U14641 (N_14641,N_14127,N_13720);
or U14642 (N_14642,N_14052,N_14058);
nand U14643 (N_14643,N_14042,N_14245);
or U14644 (N_14644,N_14357,N_13655);
xnor U14645 (N_14645,N_13660,N_14252);
nand U14646 (N_14646,N_13630,N_13796);
or U14647 (N_14647,N_13933,N_14297);
nand U14648 (N_14648,N_13846,N_14053);
nor U14649 (N_14649,N_13730,N_13712);
and U14650 (N_14650,N_14032,N_13711);
xnor U14651 (N_14651,N_14085,N_14016);
nor U14652 (N_14652,N_14022,N_14233);
nor U14653 (N_14653,N_14223,N_14162);
and U14654 (N_14654,N_14208,N_14368);
nor U14655 (N_14655,N_13890,N_14302);
xnor U14656 (N_14656,N_14257,N_14041);
and U14657 (N_14657,N_13965,N_14110);
nand U14658 (N_14658,N_14210,N_14180);
or U14659 (N_14659,N_14119,N_13876);
or U14660 (N_14660,N_13860,N_13925);
nor U14661 (N_14661,N_14011,N_13984);
nand U14662 (N_14662,N_13857,N_14135);
xor U14663 (N_14663,N_13646,N_14184);
xnor U14664 (N_14664,N_14247,N_13887);
or U14665 (N_14665,N_13897,N_13682);
or U14666 (N_14666,N_14019,N_13865);
nor U14667 (N_14667,N_13674,N_14350);
nor U14668 (N_14668,N_14087,N_14183);
nand U14669 (N_14669,N_13699,N_13781);
nor U14670 (N_14670,N_13623,N_13785);
and U14671 (N_14671,N_14224,N_13611);
and U14672 (N_14672,N_14352,N_13686);
or U14673 (N_14673,N_13622,N_13942);
xnor U14674 (N_14674,N_14343,N_13992);
nand U14675 (N_14675,N_13694,N_14091);
or U14676 (N_14676,N_13977,N_13657);
nor U14677 (N_14677,N_14093,N_13649);
nor U14678 (N_14678,N_13901,N_13653);
and U14679 (N_14679,N_14264,N_13885);
nor U14680 (N_14680,N_13867,N_13702);
nor U14681 (N_14681,N_14213,N_13607);
or U14682 (N_14682,N_13606,N_14000);
nand U14683 (N_14683,N_13637,N_13741);
nand U14684 (N_14684,N_14231,N_14169);
nand U14685 (N_14685,N_13677,N_14249);
nand U14686 (N_14686,N_14129,N_14062);
or U14687 (N_14687,N_13798,N_14226);
nand U14688 (N_14688,N_14051,N_14050);
nor U14689 (N_14689,N_14173,N_13855);
and U14690 (N_14690,N_14310,N_14043);
and U14691 (N_14691,N_13906,N_13642);
or U14692 (N_14692,N_14298,N_13920);
nand U14693 (N_14693,N_14388,N_14263);
nand U14694 (N_14694,N_13927,N_14338);
nand U14695 (N_14695,N_14161,N_14065);
or U14696 (N_14696,N_14222,N_13862);
nor U14697 (N_14697,N_14356,N_13710);
and U14698 (N_14698,N_14324,N_14364);
and U14699 (N_14699,N_13917,N_14320);
nand U14700 (N_14700,N_13618,N_13629);
xor U14701 (N_14701,N_14270,N_13953);
nand U14702 (N_14702,N_14396,N_13852);
xnor U14703 (N_14703,N_13946,N_13869);
nor U14704 (N_14704,N_14309,N_13900);
nand U14705 (N_14705,N_13609,N_13943);
nor U14706 (N_14706,N_14018,N_13713);
nor U14707 (N_14707,N_14172,N_14072);
nor U14708 (N_14708,N_14299,N_14069);
xnor U14709 (N_14709,N_13979,N_14120);
xor U14710 (N_14710,N_14191,N_13768);
nand U14711 (N_14711,N_14131,N_14076);
and U14712 (N_14712,N_14005,N_14304);
or U14713 (N_14713,N_14211,N_14232);
and U14714 (N_14714,N_13704,N_14206);
xor U14715 (N_14715,N_13909,N_14246);
nor U14716 (N_14716,N_14266,N_13967);
and U14717 (N_14717,N_13891,N_14144);
nor U14718 (N_14718,N_13737,N_13945);
and U14719 (N_14719,N_14332,N_13648);
xor U14720 (N_14720,N_13613,N_13624);
xnor U14721 (N_14721,N_14095,N_13910);
or U14722 (N_14722,N_13733,N_14015);
or U14723 (N_14723,N_13985,N_14107);
nor U14724 (N_14724,N_13662,N_14028);
or U14725 (N_14725,N_13895,N_14009);
or U14726 (N_14726,N_14272,N_13614);
and U14727 (N_14727,N_14393,N_13765);
nand U14728 (N_14728,N_14240,N_14286);
and U14729 (N_14729,N_14010,N_13719);
and U14730 (N_14730,N_14192,N_13681);
and U14731 (N_14731,N_14199,N_13826);
nor U14732 (N_14732,N_14045,N_14390);
or U14733 (N_14733,N_13807,N_14238);
xnor U14734 (N_14734,N_13787,N_13667);
nand U14735 (N_14735,N_14198,N_13625);
nand U14736 (N_14736,N_13937,N_14034);
xnor U14737 (N_14737,N_13940,N_14164);
or U14738 (N_14738,N_13894,N_13635);
nor U14739 (N_14739,N_14109,N_13811);
or U14740 (N_14740,N_13916,N_13988);
nor U14741 (N_14741,N_14307,N_14082);
or U14742 (N_14742,N_14099,N_13685);
nand U14743 (N_14743,N_13722,N_14330);
nor U14744 (N_14744,N_14335,N_14122);
xnor U14745 (N_14745,N_14130,N_13812);
or U14746 (N_14746,N_14281,N_13752);
or U14747 (N_14747,N_13640,N_14394);
nor U14748 (N_14748,N_14248,N_13983);
nor U14749 (N_14749,N_14365,N_13975);
xnor U14750 (N_14750,N_13931,N_13877);
xor U14751 (N_14751,N_13990,N_13760);
or U14752 (N_14752,N_13949,N_13830);
or U14753 (N_14753,N_14185,N_13759);
xnor U14754 (N_14754,N_14040,N_14256);
nor U14755 (N_14755,N_14057,N_14336);
nor U14756 (N_14756,N_14136,N_13627);
xor U14757 (N_14757,N_14003,N_13976);
nand U14758 (N_14758,N_14059,N_13671);
nand U14759 (N_14759,N_14219,N_14025);
nand U14760 (N_14760,N_14197,N_13810);
nor U14761 (N_14761,N_14114,N_13750);
or U14762 (N_14762,N_13748,N_13835);
xor U14763 (N_14763,N_14285,N_13788);
xor U14764 (N_14764,N_13843,N_14089);
and U14765 (N_14765,N_14158,N_14092);
or U14766 (N_14766,N_13987,N_14259);
xor U14767 (N_14767,N_13896,N_14012);
nor U14768 (N_14768,N_13952,N_14207);
or U14769 (N_14769,N_14047,N_14300);
or U14770 (N_14770,N_13828,N_13821);
nor U14771 (N_14771,N_14275,N_13898);
and U14772 (N_14772,N_13691,N_13643);
nand U14773 (N_14773,N_13769,N_14351);
xor U14774 (N_14774,N_13847,N_14243);
nor U14775 (N_14775,N_13782,N_13670);
and U14776 (N_14776,N_14141,N_14189);
xor U14777 (N_14777,N_14293,N_13754);
and U14778 (N_14778,N_14171,N_14086);
and U14779 (N_14779,N_13793,N_13707);
nor U14780 (N_14780,N_14373,N_13799);
and U14781 (N_14781,N_14303,N_14151);
or U14782 (N_14782,N_13696,N_14308);
nand U14783 (N_14783,N_13813,N_14317);
xor U14784 (N_14784,N_13939,N_14384);
nor U14785 (N_14785,N_14389,N_13680);
nand U14786 (N_14786,N_14225,N_13602);
xnor U14787 (N_14787,N_14289,N_13878);
nand U14788 (N_14788,N_14154,N_13853);
and U14789 (N_14789,N_13700,N_14291);
or U14790 (N_14790,N_14392,N_13858);
and U14791 (N_14791,N_14031,N_13708);
nor U14792 (N_14792,N_14331,N_14262);
or U14793 (N_14793,N_13721,N_14170);
or U14794 (N_14794,N_13727,N_13859);
nand U14795 (N_14795,N_14153,N_13743);
nor U14796 (N_14796,N_14284,N_14179);
xnor U14797 (N_14797,N_14187,N_14287);
nand U14798 (N_14798,N_14149,N_13814);
nand U14799 (N_14799,N_14250,N_13996);
or U14800 (N_14800,N_14044,N_14012);
and U14801 (N_14801,N_14107,N_14170);
nor U14802 (N_14802,N_13807,N_13852);
and U14803 (N_14803,N_13708,N_14105);
or U14804 (N_14804,N_13621,N_13969);
nand U14805 (N_14805,N_13913,N_13943);
and U14806 (N_14806,N_14349,N_13789);
nor U14807 (N_14807,N_14159,N_13678);
and U14808 (N_14808,N_14361,N_14066);
and U14809 (N_14809,N_14024,N_13748);
and U14810 (N_14810,N_13985,N_13701);
xnor U14811 (N_14811,N_14127,N_13703);
and U14812 (N_14812,N_13706,N_14297);
nor U14813 (N_14813,N_13986,N_14159);
nor U14814 (N_14814,N_13803,N_13708);
xnor U14815 (N_14815,N_13996,N_14326);
or U14816 (N_14816,N_13951,N_13812);
nand U14817 (N_14817,N_13758,N_14072);
nor U14818 (N_14818,N_13928,N_13666);
and U14819 (N_14819,N_13688,N_13963);
nand U14820 (N_14820,N_14356,N_14027);
and U14821 (N_14821,N_13863,N_14020);
nand U14822 (N_14822,N_14342,N_14161);
nor U14823 (N_14823,N_13787,N_13611);
xor U14824 (N_14824,N_14390,N_13930);
or U14825 (N_14825,N_14173,N_13814);
nand U14826 (N_14826,N_14118,N_14017);
and U14827 (N_14827,N_13697,N_14094);
nand U14828 (N_14828,N_13999,N_14174);
nand U14829 (N_14829,N_14141,N_14030);
and U14830 (N_14830,N_14342,N_13684);
or U14831 (N_14831,N_14176,N_13924);
nor U14832 (N_14832,N_13637,N_13914);
xnor U14833 (N_14833,N_13958,N_14278);
xor U14834 (N_14834,N_14354,N_14046);
nor U14835 (N_14835,N_13913,N_13840);
xnor U14836 (N_14836,N_14147,N_14218);
or U14837 (N_14837,N_13966,N_13684);
nand U14838 (N_14838,N_14387,N_14110);
or U14839 (N_14839,N_14228,N_13747);
nand U14840 (N_14840,N_14371,N_13894);
nand U14841 (N_14841,N_14211,N_14353);
and U14842 (N_14842,N_14053,N_13974);
or U14843 (N_14843,N_14019,N_13823);
nor U14844 (N_14844,N_14318,N_14393);
and U14845 (N_14845,N_13658,N_14390);
nand U14846 (N_14846,N_14017,N_14376);
nor U14847 (N_14847,N_14265,N_13716);
or U14848 (N_14848,N_14278,N_13817);
nor U14849 (N_14849,N_14286,N_13862);
nor U14850 (N_14850,N_13693,N_14171);
nand U14851 (N_14851,N_13781,N_13923);
or U14852 (N_14852,N_13887,N_13891);
or U14853 (N_14853,N_13998,N_14194);
xor U14854 (N_14854,N_13988,N_13670);
or U14855 (N_14855,N_13820,N_14235);
nand U14856 (N_14856,N_14056,N_13854);
or U14857 (N_14857,N_14152,N_14083);
xor U14858 (N_14858,N_14308,N_14217);
xnor U14859 (N_14859,N_14239,N_13990);
xnor U14860 (N_14860,N_13835,N_14292);
xor U14861 (N_14861,N_14215,N_13615);
and U14862 (N_14862,N_13878,N_14057);
nor U14863 (N_14863,N_14160,N_14219);
nor U14864 (N_14864,N_13941,N_13866);
xor U14865 (N_14865,N_14123,N_13697);
nor U14866 (N_14866,N_13735,N_14223);
nor U14867 (N_14867,N_14369,N_14252);
nand U14868 (N_14868,N_14028,N_14015);
xor U14869 (N_14869,N_13689,N_13966);
or U14870 (N_14870,N_14336,N_13653);
nand U14871 (N_14871,N_13875,N_13874);
nor U14872 (N_14872,N_14207,N_13972);
or U14873 (N_14873,N_13682,N_13700);
nand U14874 (N_14874,N_14363,N_14086);
nor U14875 (N_14875,N_13933,N_14260);
nand U14876 (N_14876,N_14055,N_14304);
or U14877 (N_14877,N_14253,N_14076);
or U14878 (N_14878,N_13825,N_13995);
xor U14879 (N_14879,N_14214,N_14127);
nor U14880 (N_14880,N_13632,N_14094);
xnor U14881 (N_14881,N_13982,N_14346);
nand U14882 (N_14882,N_13679,N_14330);
xor U14883 (N_14883,N_13608,N_13611);
or U14884 (N_14884,N_14210,N_14276);
nor U14885 (N_14885,N_14353,N_13723);
or U14886 (N_14886,N_13973,N_13666);
or U14887 (N_14887,N_14227,N_14256);
nand U14888 (N_14888,N_13724,N_14276);
xor U14889 (N_14889,N_14078,N_13938);
nand U14890 (N_14890,N_14232,N_14194);
or U14891 (N_14891,N_14245,N_13809);
xor U14892 (N_14892,N_14295,N_14021);
nand U14893 (N_14893,N_14252,N_13688);
nor U14894 (N_14894,N_13961,N_14223);
nor U14895 (N_14895,N_13726,N_13690);
nor U14896 (N_14896,N_13910,N_13662);
xnor U14897 (N_14897,N_13701,N_13833);
nand U14898 (N_14898,N_14285,N_13627);
nand U14899 (N_14899,N_14042,N_14359);
nand U14900 (N_14900,N_13695,N_13754);
or U14901 (N_14901,N_14267,N_13739);
or U14902 (N_14902,N_13640,N_13753);
and U14903 (N_14903,N_13828,N_13907);
and U14904 (N_14904,N_13902,N_14305);
nand U14905 (N_14905,N_13639,N_14386);
or U14906 (N_14906,N_14231,N_13753);
nor U14907 (N_14907,N_14187,N_13992);
nor U14908 (N_14908,N_13810,N_13606);
or U14909 (N_14909,N_14022,N_14094);
or U14910 (N_14910,N_14253,N_14259);
nand U14911 (N_14911,N_14244,N_14351);
nor U14912 (N_14912,N_14170,N_14121);
and U14913 (N_14913,N_14141,N_14097);
or U14914 (N_14914,N_13748,N_13818);
or U14915 (N_14915,N_14006,N_13825);
nor U14916 (N_14916,N_13922,N_13817);
or U14917 (N_14917,N_13623,N_13703);
xnor U14918 (N_14918,N_13958,N_14052);
xor U14919 (N_14919,N_14360,N_13941);
nand U14920 (N_14920,N_14080,N_14007);
nand U14921 (N_14921,N_13751,N_14134);
and U14922 (N_14922,N_13857,N_13640);
xnor U14923 (N_14923,N_14315,N_13979);
xnor U14924 (N_14924,N_13928,N_13789);
xnor U14925 (N_14925,N_13888,N_13647);
nand U14926 (N_14926,N_14287,N_13894);
xnor U14927 (N_14927,N_13684,N_13814);
or U14928 (N_14928,N_14139,N_14215);
nor U14929 (N_14929,N_13929,N_13910);
or U14930 (N_14930,N_13855,N_14002);
or U14931 (N_14931,N_14301,N_14316);
or U14932 (N_14932,N_13746,N_14252);
nand U14933 (N_14933,N_14055,N_13957);
or U14934 (N_14934,N_14386,N_13656);
nor U14935 (N_14935,N_14122,N_14263);
nor U14936 (N_14936,N_14193,N_13869);
xnor U14937 (N_14937,N_14257,N_13649);
nor U14938 (N_14938,N_14021,N_14038);
and U14939 (N_14939,N_14258,N_13830);
and U14940 (N_14940,N_13842,N_13714);
or U14941 (N_14941,N_13877,N_14385);
and U14942 (N_14942,N_13834,N_13958);
and U14943 (N_14943,N_13930,N_13867);
nand U14944 (N_14944,N_14298,N_13826);
and U14945 (N_14945,N_13801,N_14123);
xor U14946 (N_14946,N_13869,N_13705);
or U14947 (N_14947,N_13909,N_13754);
or U14948 (N_14948,N_14184,N_13951);
nor U14949 (N_14949,N_14116,N_13635);
and U14950 (N_14950,N_14185,N_13914);
xor U14951 (N_14951,N_14148,N_13787);
xnor U14952 (N_14952,N_14394,N_13891);
nor U14953 (N_14953,N_14002,N_14186);
nand U14954 (N_14954,N_14101,N_14163);
nor U14955 (N_14955,N_14348,N_13740);
or U14956 (N_14956,N_13992,N_13917);
nor U14957 (N_14957,N_13926,N_13763);
or U14958 (N_14958,N_13805,N_13628);
nand U14959 (N_14959,N_14075,N_14036);
and U14960 (N_14960,N_13919,N_14221);
nand U14961 (N_14961,N_13850,N_14312);
xnor U14962 (N_14962,N_13953,N_14161);
or U14963 (N_14963,N_13620,N_13810);
and U14964 (N_14964,N_14208,N_13911);
xnor U14965 (N_14965,N_14346,N_14192);
and U14966 (N_14966,N_14390,N_14261);
nor U14967 (N_14967,N_14363,N_13725);
or U14968 (N_14968,N_14376,N_14226);
nor U14969 (N_14969,N_13678,N_13910);
nor U14970 (N_14970,N_14189,N_13650);
or U14971 (N_14971,N_14179,N_14097);
or U14972 (N_14972,N_13823,N_14330);
nand U14973 (N_14973,N_14364,N_14210);
nor U14974 (N_14974,N_14099,N_13736);
and U14975 (N_14975,N_14009,N_13898);
and U14976 (N_14976,N_14228,N_14033);
nor U14977 (N_14977,N_13898,N_14302);
nand U14978 (N_14978,N_13735,N_14159);
or U14979 (N_14979,N_13845,N_13822);
nand U14980 (N_14980,N_13672,N_13861);
nand U14981 (N_14981,N_14176,N_13776);
or U14982 (N_14982,N_13930,N_14144);
nor U14983 (N_14983,N_14127,N_13853);
nand U14984 (N_14984,N_13763,N_14209);
and U14985 (N_14985,N_13940,N_13785);
nor U14986 (N_14986,N_14133,N_13929);
or U14987 (N_14987,N_13867,N_13785);
xnor U14988 (N_14988,N_13760,N_14184);
nand U14989 (N_14989,N_13690,N_13860);
and U14990 (N_14990,N_14331,N_13841);
nor U14991 (N_14991,N_13731,N_13966);
nand U14992 (N_14992,N_13993,N_14178);
or U14993 (N_14993,N_13638,N_14061);
or U14994 (N_14994,N_14199,N_14101);
xnor U14995 (N_14995,N_14155,N_14019);
or U14996 (N_14996,N_14197,N_13892);
or U14997 (N_14997,N_14354,N_14208);
nor U14998 (N_14998,N_13832,N_13895);
nand U14999 (N_14999,N_13783,N_13721);
xor U15000 (N_15000,N_13636,N_13949);
nand U15001 (N_15001,N_13776,N_14061);
nand U15002 (N_15002,N_14183,N_13908);
nand U15003 (N_15003,N_14139,N_13630);
or U15004 (N_15004,N_14209,N_13870);
or U15005 (N_15005,N_14276,N_13793);
nor U15006 (N_15006,N_14057,N_13820);
nand U15007 (N_15007,N_14118,N_13844);
xnor U15008 (N_15008,N_14240,N_14242);
xor U15009 (N_15009,N_14262,N_14109);
or U15010 (N_15010,N_14217,N_14366);
xnor U15011 (N_15011,N_14259,N_13677);
nor U15012 (N_15012,N_13695,N_14209);
and U15013 (N_15013,N_13804,N_13917);
nor U15014 (N_15014,N_13647,N_14099);
nor U15015 (N_15015,N_14241,N_14183);
or U15016 (N_15016,N_13657,N_14212);
nor U15017 (N_15017,N_14276,N_14399);
and U15018 (N_15018,N_13629,N_14356);
xnor U15019 (N_15019,N_13843,N_13606);
xnor U15020 (N_15020,N_13994,N_14035);
nand U15021 (N_15021,N_13668,N_14197);
xnor U15022 (N_15022,N_13709,N_13707);
nand U15023 (N_15023,N_14260,N_14392);
xnor U15024 (N_15024,N_14001,N_14017);
nand U15025 (N_15025,N_13964,N_13929);
and U15026 (N_15026,N_13875,N_14262);
xor U15027 (N_15027,N_13698,N_13760);
or U15028 (N_15028,N_14150,N_13932);
or U15029 (N_15029,N_13955,N_14380);
or U15030 (N_15030,N_14232,N_13686);
xor U15031 (N_15031,N_13920,N_13928);
and U15032 (N_15032,N_14001,N_13794);
xor U15033 (N_15033,N_14068,N_14240);
nor U15034 (N_15034,N_13630,N_14275);
or U15035 (N_15035,N_13714,N_13954);
and U15036 (N_15036,N_14024,N_14364);
nand U15037 (N_15037,N_13802,N_13973);
nand U15038 (N_15038,N_14114,N_13956);
and U15039 (N_15039,N_14386,N_13796);
nor U15040 (N_15040,N_13729,N_13900);
xor U15041 (N_15041,N_14233,N_13649);
nand U15042 (N_15042,N_14327,N_14050);
nand U15043 (N_15043,N_14287,N_14000);
or U15044 (N_15044,N_14372,N_13771);
nand U15045 (N_15045,N_13896,N_13709);
nor U15046 (N_15046,N_13618,N_13788);
xor U15047 (N_15047,N_14106,N_14366);
nand U15048 (N_15048,N_14293,N_13734);
nor U15049 (N_15049,N_13868,N_14373);
nand U15050 (N_15050,N_13952,N_13678);
nor U15051 (N_15051,N_14308,N_13976);
nand U15052 (N_15052,N_13769,N_13602);
xor U15053 (N_15053,N_14387,N_14309);
nor U15054 (N_15054,N_14373,N_13899);
or U15055 (N_15055,N_14189,N_13953);
and U15056 (N_15056,N_14082,N_13815);
nand U15057 (N_15057,N_14055,N_14134);
nor U15058 (N_15058,N_14151,N_14248);
nand U15059 (N_15059,N_14175,N_14117);
xnor U15060 (N_15060,N_13928,N_14260);
nor U15061 (N_15061,N_13727,N_14319);
nor U15062 (N_15062,N_14262,N_13967);
nor U15063 (N_15063,N_13788,N_14138);
and U15064 (N_15064,N_13930,N_14059);
nor U15065 (N_15065,N_13609,N_14184);
nand U15066 (N_15066,N_14372,N_13603);
nor U15067 (N_15067,N_13740,N_13752);
and U15068 (N_15068,N_13983,N_13891);
nor U15069 (N_15069,N_14389,N_14071);
nand U15070 (N_15070,N_13649,N_13650);
or U15071 (N_15071,N_13664,N_14038);
xnor U15072 (N_15072,N_13825,N_14344);
or U15073 (N_15073,N_13646,N_14316);
nor U15074 (N_15074,N_14157,N_13938);
or U15075 (N_15075,N_13758,N_14177);
or U15076 (N_15076,N_13681,N_14183);
and U15077 (N_15077,N_13746,N_14393);
or U15078 (N_15078,N_14395,N_14186);
nand U15079 (N_15079,N_14352,N_13786);
nand U15080 (N_15080,N_13630,N_14007);
or U15081 (N_15081,N_14119,N_14382);
xor U15082 (N_15082,N_13897,N_14205);
or U15083 (N_15083,N_13706,N_13877);
nor U15084 (N_15084,N_13831,N_14387);
nand U15085 (N_15085,N_13928,N_13628);
nand U15086 (N_15086,N_13672,N_13760);
xor U15087 (N_15087,N_13754,N_13899);
or U15088 (N_15088,N_14050,N_14111);
nand U15089 (N_15089,N_13684,N_13762);
or U15090 (N_15090,N_14179,N_14020);
and U15091 (N_15091,N_13898,N_13795);
and U15092 (N_15092,N_13805,N_13827);
and U15093 (N_15093,N_13722,N_14257);
xor U15094 (N_15094,N_13970,N_13617);
and U15095 (N_15095,N_14381,N_13954);
nand U15096 (N_15096,N_14357,N_13863);
and U15097 (N_15097,N_14047,N_13919);
xnor U15098 (N_15098,N_14067,N_14002);
or U15099 (N_15099,N_14196,N_13664);
and U15100 (N_15100,N_14056,N_14309);
and U15101 (N_15101,N_14358,N_14355);
or U15102 (N_15102,N_14257,N_14153);
nor U15103 (N_15103,N_14252,N_14137);
and U15104 (N_15104,N_13716,N_13947);
nor U15105 (N_15105,N_13862,N_13864);
or U15106 (N_15106,N_13933,N_13974);
xnor U15107 (N_15107,N_14344,N_14176);
xor U15108 (N_15108,N_13663,N_14041);
nand U15109 (N_15109,N_13600,N_13705);
xor U15110 (N_15110,N_14276,N_13723);
and U15111 (N_15111,N_13855,N_14356);
nor U15112 (N_15112,N_13730,N_14372);
nand U15113 (N_15113,N_14113,N_14237);
nand U15114 (N_15114,N_13729,N_13759);
and U15115 (N_15115,N_13629,N_13779);
and U15116 (N_15116,N_13732,N_14108);
nand U15117 (N_15117,N_14105,N_14115);
and U15118 (N_15118,N_13813,N_13832);
xnor U15119 (N_15119,N_13922,N_13887);
or U15120 (N_15120,N_14059,N_14304);
and U15121 (N_15121,N_14374,N_14353);
and U15122 (N_15122,N_13681,N_13892);
or U15123 (N_15123,N_13893,N_13866);
nand U15124 (N_15124,N_13916,N_13996);
or U15125 (N_15125,N_14105,N_14296);
nor U15126 (N_15126,N_13700,N_13653);
or U15127 (N_15127,N_13855,N_13984);
and U15128 (N_15128,N_14205,N_13766);
or U15129 (N_15129,N_13952,N_13920);
nand U15130 (N_15130,N_14230,N_14296);
xor U15131 (N_15131,N_13757,N_14100);
nor U15132 (N_15132,N_14052,N_13636);
nand U15133 (N_15133,N_14285,N_14199);
nand U15134 (N_15134,N_14018,N_13744);
xor U15135 (N_15135,N_13765,N_14160);
nand U15136 (N_15136,N_14266,N_13638);
and U15137 (N_15137,N_13657,N_13619);
nand U15138 (N_15138,N_13792,N_13921);
nand U15139 (N_15139,N_14201,N_14133);
nand U15140 (N_15140,N_14242,N_14133);
and U15141 (N_15141,N_13979,N_13942);
nand U15142 (N_15142,N_13706,N_13856);
and U15143 (N_15143,N_13670,N_14161);
xor U15144 (N_15144,N_13669,N_13821);
nand U15145 (N_15145,N_14080,N_13946);
nand U15146 (N_15146,N_13602,N_14378);
xor U15147 (N_15147,N_13903,N_14346);
xnor U15148 (N_15148,N_14328,N_13697);
nor U15149 (N_15149,N_13659,N_14364);
nor U15150 (N_15150,N_14114,N_13734);
or U15151 (N_15151,N_14021,N_13884);
xor U15152 (N_15152,N_13756,N_14371);
nand U15153 (N_15153,N_14302,N_13755);
nor U15154 (N_15154,N_14199,N_14185);
or U15155 (N_15155,N_13743,N_13708);
or U15156 (N_15156,N_13901,N_14251);
xnor U15157 (N_15157,N_14255,N_14309);
xor U15158 (N_15158,N_14211,N_13938);
or U15159 (N_15159,N_14028,N_13744);
nand U15160 (N_15160,N_14010,N_13835);
and U15161 (N_15161,N_13884,N_14170);
or U15162 (N_15162,N_13908,N_14075);
and U15163 (N_15163,N_14132,N_14277);
or U15164 (N_15164,N_14235,N_13731);
nor U15165 (N_15165,N_13859,N_13669);
nand U15166 (N_15166,N_14370,N_13941);
xor U15167 (N_15167,N_13925,N_14004);
and U15168 (N_15168,N_13693,N_14317);
and U15169 (N_15169,N_14261,N_13720);
xnor U15170 (N_15170,N_13693,N_13953);
xor U15171 (N_15171,N_14341,N_13731);
nor U15172 (N_15172,N_14001,N_13680);
or U15173 (N_15173,N_14362,N_13991);
nor U15174 (N_15174,N_14047,N_13682);
xnor U15175 (N_15175,N_14083,N_14075);
nand U15176 (N_15176,N_14022,N_13799);
nand U15177 (N_15177,N_13706,N_13798);
and U15178 (N_15178,N_14129,N_13769);
xnor U15179 (N_15179,N_14383,N_14307);
xor U15180 (N_15180,N_13931,N_13950);
xnor U15181 (N_15181,N_13780,N_13855);
or U15182 (N_15182,N_14168,N_13669);
or U15183 (N_15183,N_13963,N_14217);
xor U15184 (N_15184,N_13853,N_13979);
or U15185 (N_15185,N_14337,N_14211);
and U15186 (N_15186,N_14293,N_14082);
nand U15187 (N_15187,N_14079,N_14212);
xor U15188 (N_15188,N_14072,N_13882);
or U15189 (N_15189,N_14394,N_13675);
and U15190 (N_15190,N_14202,N_14298);
nor U15191 (N_15191,N_14038,N_14182);
xnor U15192 (N_15192,N_13805,N_13779);
or U15193 (N_15193,N_14021,N_13710);
or U15194 (N_15194,N_13940,N_14062);
or U15195 (N_15195,N_14064,N_13932);
nand U15196 (N_15196,N_14179,N_14283);
or U15197 (N_15197,N_13667,N_13872);
nand U15198 (N_15198,N_13920,N_13708);
nand U15199 (N_15199,N_13908,N_14277);
and U15200 (N_15200,N_14728,N_14919);
xor U15201 (N_15201,N_15005,N_14450);
nor U15202 (N_15202,N_15101,N_15053);
and U15203 (N_15203,N_15042,N_14480);
nand U15204 (N_15204,N_14811,N_14851);
or U15205 (N_15205,N_14866,N_14446);
nand U15206 (N_15206,N_14910,N_14889);
or U15207 (N_15207,N_14602,N_14463);
and U15208 (N_15208,N_14568,N_14922);
xor U15209 (N_15209,N_14458,N_15084);
nand U15210 (N_15210,N_15013,N_15122);
xor U15211 (N_15211,N_15108,N_14794);
or U15212 (N_15212,N_14503,N_14803);
xnor U15213 (N_15213,N_14756,N_15052);
or U15214 (N_15214,N_14507,N_14600);
and U15215 (N_15215,N_14896,N_14716);
or U15216 (N_15216,N_14758,N_14850);
or U15217 (N_15217,N_14893,N_14683);
and U15218 (N_15218,N_15006,N_14938);
and U15219 (N_15219,N_14406,N_15123);
xnor U15220 (N_15220,N_14501,N_15025);
nor U15221 (N_15221,N_14781,N_14820);
xor U15222 (N_15222,N_15009,N_15125);
xnor U15223 (N_15223,N_15104,N_14906);
nor U15224 (N_15224,N_14802,N_14936);
nand U15225 (N_15225,N_14885,N_14512);
and U15226 (N_15226,N_15197,N_15070);
xnor U15227 (N_15227,N_14527,N_14477);
xnor U15228 (N_15228,N_14598,N_14740);
and U15229 (N_15229,N_14572,N_14681);
or U15230 (N_15230,N_14551,N_14879);
xnor U15231 (N_15231,N_14881,N_14427);
nand U15232 (N_15232,N_14968,N_14675);
xnor U15233 (N_15233,N_14679,N_15124);
nand U15234 (N_15234,N_14935,N_15198);
nand U15235 (N_15235,N_14953,N_15174);
and U15236 (N_15236,N_14791,N_15026);
and U15237 (N_15237,N_15173,N_14495);
nand U15238 (N_15238,N_15160,N_15003);
nor U15239 (N_15239,N_14698,N_14974);
and U15240 (N_15240,N_15170,N_14521);
nand U15241 (N_15241,N_15179,N_14497);
nor U15242 (N_15242,N_14606,N_14932);
nor U15243 (N_15243,N_15154,N_14731);
xor U15244 (N_15244,N_14877,N_14928);
nor U15245 (N_15245,N_14601,N_14933);
or U15246 (N_15246,N_14711,N_15119);
or U15247 (N_15247,N_14854,N_14920);
and U15248 (N_15248,N_14641,N_15061);
or U15249 (N_15249,N_15151,N_14868);
and U15250 (N_15250,N_14437,N_14487);
xor U15251 (N_15251,N_14636,N_14952);
and U15252 (N_15252,N_14682,N_14685);
nand U15253 (N_15253,N_14482,N_15021);
and U15254 (N_15254,N_15004,N_14415);
and U15255 (N_15255,N_14614,N_14703);
xor U15256 (N_15256,N_15157,N_15008);
and U15257 (N_15257,N_14648,N_15071);
and U15258 (N_15258,N_14806,N_14823);
and U15259 (N_15259,N_14900,N_14566);
or U15260 (N_15260,N_14849,N_15103);
nor U15261 (N_15261,N_14701,N_15128);
or U15262 (N_15262,N_14543,N_14765);
nor U15263 (N_15263,N_14515,N_14493);
xnor U15264 (N_15264,N_15059,N_14770);
nor U15265 (N_15265,N_15145,N_14502);
and U15266 (N_15266,N_14671,N_14821);
xnor U15267 (N_15267,N_14419,N_14736);
xnor U15268 (N_15268,N_14545,N_15001);
and U15269 (N_15269,N_14757,N_15060);
or U15270 (N_15270,N_14622,N_15153);
and U15271 (N_15271,N_15097,N_14788);
xnor U15272 (N_15272,N_14976,N_14407);
and U15273 (N_15273,N_14471,N_14633);
xor U15274 (N_15274,N_14474,N_14750);
nand U15275 (N_15275,N_15164,N_14635);
xor U15276 (N_15276,N_15020,N_14967);
or U15277 (N_15277,N_14715,N_15117);
nand U15278 (N_15278,N_15002,N_14466);
nor U15279 (N_15279,N_15148,N_14833);
or U15280 (N_15280,N_14894,N_15098);
xnor U15281 (N_15281,N_15115,N_14447);
xnor U15282 (N_15282,N_14804,N_14810);
xnor U15283 (N_15283,N_14537,N_15024);
nand U15284 (N_15284,N_15193,N_14774);
nand U15285 (N_15285,N_14608,N_14816);
nand U15286 (N_15286,N_15137,N_15022);
or U15287 (N_15287,N_14959,N_14946);
nand U15288 (N_15288,N_14637,N_14766);
or U15289 (N_15289,N_14941,N_14878);
and U15290 (N_15290,N_14873,N_15109);
nor U15291 (N_15291,N_14827,N_14875);
nand U15292 (N_15292,N_14588,N_14525);
and U15293 (N_15293,N_15017,N_14699);
or U15294 (N_15294,N_15045,N_14678);
or U15295 (N_15295,N_14891,N_14596);
or U15296 (N_15296,N_14644,N_14949);
or U15297 (N_15297,N_14755,N_14653);
or U15298 (N_15298,N_14921,N_15090);
and U15299 (N_15299,N_14552,N_15144);
nand U15300 (N_15300,N_14761,N_15027);
nand U15301 (N_15301,N_14506,N_14970);
and U15302 (N_15302,N_14533,N_15032);
and U15303 (N_15303,N_14798,N_14559);
or U15304 (N_15304,N_14713,N_14937);
and U15305 (N_15305,N_14915,N_14829);
xnor U15306 (N_15306,N_14416,N_14847);
and U15307 (N_15307,N_15036,N_14789);
nor U15308 (N_15308,N_14853,N_14705);
nand U15309 (N_15309,N_14609,N_14410);
nand U15310 (N_15310,N_14725,N_14613);
nand U15311 (N_15311,N_14759,N_14790);
and U15312 (N_15312,N_14871,N_14752);
and U15313 (N_15313,N_14729,N_14425);
nor U15314 (N_15314,N_15142,N_14467);
nor U15315 (N_15315,N_14695,N_14586);
xor U15316 (N_15316,N_14627,N_14992);
or U15317 (N_15317,N_14401,N_14488);
or U15318 (N_15318,N_14923,N_14538);
xor U15319 (N_15319,N_15031,N_14697);
nand U15320 (N_15320,N_15030,N_14408);
or U15321 (N_15321,N_15107,N_15092);
xnor U15322 (N_15322,N_14777,N_15106);
xnor U15323 (N_15323,N_14996,N_15043);
xor U15324 (N_15324,N_14420,N_14452);
or U15325 (N_15325,N_15188,N_14960);
xnor U15326 (N_15326,N_14978,N_15055);
xnor U15327 (N_15327,N_14579,N_14628);
xnor U15328 (N_15328,N_14592,N_14989);
nand U15329 (N_15329,N_14995,N_14824);
xor U15330 (N_15330,N_15035,N_14578);
nand U15331 (N_15331,N_14661,N_14445);
xor U15332 (N_15332,N_14856,N_14965);
or U15333 (N_15333,N_14511,N_15169);
xnor U15334 (N_15334,N_14522,N_15140);
nand U15335 (N_15335,N_15118,N_14957);
nand U15336 (N_15336,N_15029,N_14534);
or U15337 (N_15337,N_14544,N_14706);
and U15338 (N_15338,N_14916,N_14884);
nand U15339 (N_15339,N_14432,N_14745);
and U15340 (N_15340,N_14964,N_14822);
and U15341 (N_15341,N_14739,N_15180);
or U15342 (N_15342,N_14550,N_14618);
nand U15343 (N_15343,N_14412,N_15156);
nand U15344 (N_15344,N_14730,N_14616);
nand U15345 (N_15345,N_14625,N_14993);
xnor U15346 (N_15346,N_14951,N_14717);
nand U15347 (N_15347,N_14581,N_14712);
and U15348 (N_15348,N_14422,N_15175);
or U15349 (N_15349,N_14589,N_15044);
or U15350 (N_15350,N_15141,N_14404);
and U15351 (N_15351,N_14998,N_15010);
or U15352 (N_15352,N_14832,N_14863);
xor U15353 (N_15353,N_14955,N_14530);
or U15354 (N_15354,N_14457,N_14835);
nor U15355 (N_15355,N_14411,N_14859);
nor U15356 (N_15356,N_14966,N_14564);
nand U15357 (N_15357,N_15096,N_14944);
xnor U15358 (N_15358,N_14775,N_14834);
nand U15359 (N_15359,N_14561,N_14433);
or U15360 (N_15360,N_14744,N_14840);
nand U15361 (N_15361,N_14762,N_14990);
or U15362 (N_15362,N_14830,N_14418);
nand U15363 (N_15363,N_15056,N_14436);
and U15364 (N_15364,N_15102,N_14855);
or U15365 (N_15365,N_14801,N_15086);
nor U15366 (N_15366,N_15018,N_14907);
xnor U15367 (N_15367,N_14818,N_15127);
or U15368 (N_15368,N_14691,N_14465);
nor U15369 (N_15369,N_14570,N_15155);
nor U15370 (N_15370,N_14956,N_15139);
nor U15371 (N_15371,N_15136,N_15033);
nand U15372 (N_15372,N_15194,N_14431);
and U15373 (N_15373,N_14876,N_14649);
nand U15374 (N_15374,N_14647,N_14783);
nor U15375 (N_15375,N_14841,N_14831);
nand U15376 (N_15376,N_14672,N_14553);
nand U15377 (N_15377,N_14486,N_15150);
nand U15378 (N_15378,N_14554,N_14562);
or U15379 (N_15379,N_14626,N_14743);
nand U15380 (N_15380,N_14597,N_15146);
or U15381 (N_15381,N_15120,N_14604);
nand U15382 (N_15382,N_14987,N_14444);
and U15383 (N_15383,N_15057,N_14805);
nor U15384 (N_15384,N_14443,N_15165);
or U15385 (N_15385,N_14489,N_14899);
xnor U15386 (N_15386,N_15023,N_14454);
nor U15387 (N_15387,N_14720,N_14567);
xor U15388 (N_15388,N_14696,N_14531);
nand U15389 (N_15389,N_14499,N_15046);
nand U15390 (N_15390,N_14880,N_15012);
xor U15391 (N_15391,N_14557,N_14472);
nor U15392 (N_15392,N_14666,N_14476);
nor U15393 (N_15393,N_14800,N_14500);
or U15394 (N_15394,N_14931,N_14714);
nor U15395 (N_15395,N_14958,N_15171);
and U15396 (N_15396,N_15186,N_14814);
and U15397 (N_15397,N_14969,N_14947);
xor U15398 (N_15398,N_15112,N_14787);
xor U15399 (N_15399,N_14490,N_14797);
nand U15400 (N_15400,N_15129,N_14638);
nor U15401 (N_15401,N_14686,N_15050);
xor U15402 (N_15402,N_14435,N_15088);
xnor U15403 (N_15403,N_15091,N_15162);
xnor U15404 (N_15404,N_14983,N_14971);
nand U15405 (N_15405,N_14642,N_15093);
and U15406 (N_15406,N_15074,N_14828);
xnor U15407 (N_15407,N_15038,N_14895);
or U15408 (N_15408,N_14668,N_15181);
nor U15409 (N_15409,N_15048,N_14904);
or U15410 (N_15410,N_14942,N_14684);
nor U15411 (N_15411,N_14519,N_15051);
nand U15412 (N_15412,N_14903,N_14400);
nor U15413 (N_15413,N_14722,N_14930);
nor U15414 (N_15414,N_14607,N_14536);
nor U15415 (N_15415,N_14723,N_15158);
or U15416 (N_15416,N_14807,N_14979);
xor U15417 (N_15417,N_14667,N_14428);
xnor U15418 (N_15418,N_14975,N_14498);
nor U15419 (N_15419,N_14865,N_14708);
and U15420 (N_15420,N_15177,N_14929);
nand U15421 (N_15421,N_15099,N_15066);
and U15422 (N_15422,N_14605,N_14494);
nor U15423 (N_15423,N_14767,N_14496);
nor U15424 (N_15424,N_14529,N_14509);
or U15425 (N_15425,N_14540,N_14483);
and U15426 (N_15426,N_14690,N_14424);
nor U15427 (N_15427,N_15039,N_14430);
nand U15428 (N_15428,N_14776,N_15094);
xor U15429 (N_15429,N_14442,N_14663);
or U15430 (N_15430,N_14693,N_14909);
nand U15431 (N_15431,N_15133,N_15196);
and U15432 (N_15432,N_14603,N_14439);
xnor U15433 (N_15433,N_15011,N_15138);
nor U15434 (N_15434,N_14640,N_14634);
and U15435 (N_15435,N_15182,N_15015);
nor U15436 (N_15436,N_14702,N_14460);
nor U15437 (N_15437,N_14858,N_14513);
and U15438 (N_15438,N_14948,N_14643);
nand U15439 (N_15439,N_14786,N_15082);
or U15440 (N_15440,N_15166,N_14721);
and U15441 (N_15441,N_14670,N_14870);
nor U15442 (N_15442,N_14980,N_15134);
xor U15443 (N_15443,N_15034,N_14694);
nand U15444 (N_15444,N_14994,N_15110);
nor U15445 (N_15445,N_15163,N_14484);
nor U15446 (N_15446,N_14718,N_14808);
and U15447 (N_15447,N_14414,N_14913);
nor U15448 (N_15448,N_15184,N_14646);
and U15449 (N_15449,N_14481,N_15062);
nor U15450 (N_15450,N_14902,N_15068);
or U15451 (N_15451,N_14584,N_14461);
xor U15452 (N_15452,N_15195,N_14687);
nor U15453 (N_15453,N_14886,N_14520);
nor U15454 (N_15454,N_14815,N_14747);
xor U15455 (N_15455,N_15073,N_14523);
nor U15456 (N_15456,N_14857,N_14655);
xnor U15457 (N_15457,N_14785,N_14754);
nor U15458 (N_15458,N_14510,N_14429);
xnor U15459 (N_15459,N_14826,N_15172);
xor U15460 (N_15460,N_14836,N_14505);
xnor U15461 (N_15461,N_14517,N_14772);
or U15462 (N_15462,N_14573,N_14526);
nand U15463 (N_15463,N_14560,N_14571);
xnor U15464 (N_15464,N_14842,N_14763);
or U15465 (N_15465,N_14771,N_14662);
or U15466 (N_15466,N_15168,N_14676);
nand U15467 (N_15467,N_14753,N_14514);
and U15468 (N_15468,N_15135,N_15079);
or U15469 (N_15469,N_15132,N_14939);
and U15470 (N_15470,N_14485,N_15143);
xnor U15471 (N_15471,N_14438,N_14732);
and U15472 (N_15472,N_14539,N_15147);
nor U15473 (N_15473,N_14984,N_15100);
nand U15474 (N_15474,N_14576,N_14405);
and U15475 (N_15475,N_14555,N_15058);
and U15476 (N_15476,N_14898,N_14610);
and U15477 (N_15477,N_15192,N_14867);
or U15478 (N_15478,N_14469,N_14654);
or U15479 (N_15479,N_14569,N_14547);
nor U15480 (N_15480,N_14707,N_15111);
nor U15481 (N_15481,N_14908,N_14617);
nor U15482 (N_15482,N_14650,N_14426);
and U15483 (N_15483,N_14577,N_14535);
and U15484 (N_15484,N_14621,N_14925);
or U15485 (N_15485,N_15007,N_14748);
and U15486 (N_15486,N_14587,N_14599);
and U15487 (N_15487,N_14749,N_14950);
nor U15488 (N_15488,N_15063,N_14402);
nand U15489 (N_15489,N_14583,N_15085);
and U15490 (N_15490,N_14688,N_14985);
xnor U15491 (N_15491,N_14988,N_14905);
nor U15492 (N_15492,N_14524,N_14594);
xnor U15493 (N_15493,N_14981,N_14883);
nand U15494 (N_15494,N_15089,N_14677);
nand U15495 (N_15495,N_15167,N_15178);
nor U15496 (N_15496,N_14468,N_15081);
nand U15497 (N_15497,N_14735,N_14409);
nand U15498 (N_15498,N_14492,N_14882);
nand U15499 (N_15499,N_14532,N_14651);
nand U15500 (N_15500,N_14516,N_14972);
nand U15501 (N_15501,N_14779,N_15189);
xnor U15502 (N_15502,N_14817,N_14582);
and U15503 (N_15503,N_14624,N_14421);
nand U15504 (N_15504,N_14645,N_14887);
nor U15505 (N_15505,N_15087,N_14665);
xnor U15506 (N_15506,N_15037,N_14795);
xnor U15507 (N_15507,N_14778,N_14441);
nand U15508 (N_15508,N_14659,N_14977);
and U15509 (N_15509,N_15126,N_14656);
or U15510 (N_15510,N_14664,N_15187);
xnor U15511 (N_15511,N_14632,N_14591);
or U15512 (N_15512,N_14475,N_14423);
or U15513 (N_15513,N_14657,N_14741);
and U15514 (N_15514,N_14751,N_14812);
and U15515 (N_15515,N_14719,N_15113);
and U15516 (N_15516,N_14580,N_14874);
or U15517 (N_15517,N_14548,N_14997);
nand U15518 (N_15518,N_14737,N_15105);
nor U15519 (N_15519,N_14927,N_15000);
nor U15520 (N_15520,N_14542,N_14727);
xnor U15521 (N_15521,N_14926,N_15161);
nor U15522 (N_15522,N_14954,N_14961);
and U15523 (N_15523,N_14528,N_14945);
and U15524 (N_15524,N_14417,N_14615);
and U15525 (N_15525,N_14518,N_14669);
nor U15526 (N_15526,N_14837,N_14809);
and U15527 (N_15527,N_14478,N_14549);
nand U15528 (N_15528,N_15065,N_14917);
or U15529 (N_15529,N_14700,N_14704);
nor U15530 (N_15530,N_14565,N_15199);
or U15531 (N_15531,N_14403,N_14792);
nor U15532 (N_15532,N_15069,N_14862);
nand U15533 (N_15533,N_14890,N_15185);
xor U15534 (N_15534,N_14773,N_15076);
or U15535 (N_15535,N_14845,N_15019);
and U15536 (N_15536,N_14726,N_15159);
and U15537 (N_15537,N_14631,N_14943);
xor U15538 (N_15538,N_14860,N_14869);
nor U15539 (N_15539,N_14742,N_14673);
or U15540 (N_15540,N_14455,N_14462);
nor U15541 (N_15541,N_14864,N_14541);
or U15542 (N_15542,N_14660,N_14456);
nand U15543 (N_15543,N_14558,N_14440);
xor U15544 (N_15544,N_14734,N_14574);
nand U15545 (N_15545,N_14813,N_14434);
or U15546 (N_15546,N_14780,N_14629);
xnor U15547 (N_15547,N_14709,N_15130);
nor U15548 (N_15548,N_14612,N_14991);
nand U15549 (N_15549,N_14844,N_14623);
xnor U15550 (N_15550,N_14620,N_15064);
and U15551 (N_15551,N_14639,N_15054);
nand U15552 (N_15552,N_14760,N_14746);
nand U15553 (N_15553,N_14852,N_14710);
and U15554 (N_15554,N_14934,N_14448);
xor U15555 (N_15555,N_14611,N_15114);
xnor U15556 (N_15556,N_15041,N_15191);
xnor U15557 (N_15557,N_14464,N_14585);
nor U15558 (N_15558,N_14652,N_14940);
nor U15559 (N_15559,N_14764,N_15067);
nand U15560 (N_15560,N_15080,N_15047);
xnor U15561 (N_15561,N_14449,N_15152);
or U15562 (N_15562,N_14799,N_14590);
or U15563 (N_15563,N_14796,N_14453);
or U15564 (N_15564,N_14563,N_14986);
xor U15565 (N_15565,N_14508,N_15028);
xnor U15566 (N_15566,N_14872,N_14619);
xor U15567 (N_15567,N_14846,N_14733);
and U15568 (N_15568,N_15131,N_14982);
nand U15569 (N_15569,N_14861,N_14973);
and U15570 (N_15570,N_15078,N_15176);
nand U15571 (N_15571,N_15083,N_14963);
or U15572 (N_15572,N_14556,N_14630);
and U15573 (N_15573,N_14593,N_14784);
and U15574 (N_15574,N_14843,N_14888);
nand U15575 (N_15575,N_14768,N_14848);
nand U15576 (N_15576,N_14692,N_14595);
nand U15577 (N_15577,N_14839,N_14962);
xnor U15578 (N_15578,N_14914,N_14912);
nand U15579 (N_15579,N_15190,N_14546);
nand U15580 (N_15580,N_15049,N_14782);
or U15581 (N_15581,N_15040,N_14658);
or U15582 (N_15582,N_14738,N_14470);
nand U15583 (N_15583,N_15014,N_14999);
xor U15584 (N_15584,N_14918,N_14451);
xor U15585 (N_15585,N_14838,N_14689);
or U15586 (N_15586,N_15077,N_14504);
xor U15587 (N_15587,N_14819,N_15116);
and U15588 (N_15588,N_15183,N_14892);
nand U15589 (N_15589,N_14674,N_15075);
xor U15590 (N_15590,N_15095,N_14901);
or U15591 (N_15591,N_14769,N_14793);
nand U15592 (N_15592,N_14911,N_14473);
or U15593 (N_15593,N_14724,N_14575);
nor U15594 (N_15594,N_14924,N_14825);
nor U15595 (N_15595,N_14680,N_14897);
xor U15596 (N_15596,N_15072,N_14413);
nor U15597 (N_15597,N_14479,N_14459);
nor U15598 (N_15598,N_15016,N_15121);
nor U15599 (N_15599,N_14491,N_15149);
and U15600 (N_15600,N_15129,N_15155);
and U15601 (N_15601,N_14863,N_14587);
nor U15602 (N_15602,N_14933,N_14990);
and U15603 (N_15603,N_14870,N_14962);
nand U15604 (N_15604,N_14757,N_14768);
or U15605 (N_15605,N_14859,N_14503);
or U15606 (N_15606,N_14678,N_14439);
xnor U15607 (N_15607,N_14542,N_14812);
nand U15608 (N_15608,N_15149,N_14407);
or U15609 (N_15609,N_14525,N_14920);
and U15610 (N_15610,N_14846,N_14884);
nor U15611 (N_15611,N_15116,N_14678);
nand U15612 (N_15612,N_15108,N_14440);
nor U15613 (N_15613,N_14689,N_14516);
nor U15614 (N_15614,N_14641,N_15026);
nor U15615 (N_15615,N_14794,N_14464);
and U15616 (N_15616,N_14675,N_14518);
xor U15617 (N_15617,N_14485,N_14533);
nor U15618 (N_15618,N_14495,N_14549);
xnor U15619 (N_15619,N_14734,N_14530);
xor U15620 (N_15620,N_14739,N_15106);
xnor U15621 (N_15621,N_15066,N_14498);
xor U15622 (N_15622,N_14752,N_14771);
and U15623 (N_15623,N_14986,N_15121);
or U15624 (N_15624,N_14871,N_14663);
xor U15625 (N_15625,N_15002,N_14585);
xor U15626 (N_15626,N_14886,N_14681);
and U15627 (N_15627,N_14787,N_14451);
nor U15628 (N_15628,N_15138,N_14417);
nand U15629 (N_15629,N_14758,N_14558);
xnor U15630 (N_15630,N_15093,N_14428);
nand U15631 (N_15631,N_14971,N_14668);
and U15632 (N_15632,N_14502,N_14658);
and U15633 (N_15633,N_14761,N_14916);
and U15634 (N_15634,N_14733,N_14837);
nor U15635 (N_15635,N_14453,N_15064);
nand U15636 (N_15636,N_14715,N_14730);
nand U15637 (N_15637,N_14916,N_14817);
nand U15638 (N_15638,N_15010,N_14684);
xnor U15639 (N_15639,N_14622,N_14493);
nor U15640 (N_15640,N_15023,N_14612);
nor U15641 (N_15641,N_15040,N_15131);
xor U15642 (N_15642,N_14909,N_15072);
nand U15643 (N_15643,N_14526,N_15073);
nand U15644 (N_15644,N_14687,N_14598);
nand U15645 (N_15645,N_14716,N_14949);
xor U15646 (N_15646,N_14505,N_14610);
nand U15647 (N_15647,N_15152,N_14664);
nand U15648 (N_15648,N_14670,N_14557);
or U15649 (N_15649,N_14756,N_15150);
and U15650 (N_15650,N_14579,N_14523);
xnor U15651 (N_15651,N_15074,N_14421);
nand U15652 (N_15652,N_14472,N_14583);
and U15653 (N_15653,N_14762,N_14919);
or U15654 (N_15654,N_14803,N_14994);
and U15655 (N_15655,N_14588,N_15087);
or U15656 (N_15656,N_14988,N_14910);
nand U15657 (N_15657,N_14560,N_14899);
and U15658 (N_15658,N_15109,N_14541);
nand U15659 (N_15659,N_14806,N_15051);
or U15660 (N_15660,N_14428,N_15044);
xnor U15661 (N_15661,N_14793,N_15189);
or U15662 (N_15662,N_14422,N_15188);
nand U15663 (N_15663,N_14710,N_14488);
xnor U15664 (N_15664,N_14429,N_14632);
or U15665 (N_15665,N_14647,N_14938);
nand U15666 (N_15666,N_14901,N_14826);
nand U15667 (N_15667,N_14440,N_14842);
and U15668 (N_15668,N_14407,N_14533);
or U15669 (N_15669,N_14721,N_14915);
nor U15670 (N_15670,N_15092,N_14793);
or U15671 (N_15671,N_14952,N_14851);
nor U15672 (N_15672,N_14842,N_14660);
or U15673 (N_15673,N_14883,N_14757);
and U15674 (N_15674,N_14865,N_14845);
xor U15675 (N_15675,N_14519,N_14819);
xnor U15676 (N_15676,N_15115,N_15156);
and U15677 (N_15677,N_14718,N_14431);
nor U15678 (N_15678,N_14926,N_14553);
xor U15679 (N_15679,N_14918,N_14535);
nand U15680 (N_15680,N_14419,N_14741);
xor U15681 (N_15681,N_14587,N_14463);
xor U15682 (N_15682,N_14955,N_15098);
or U15683 (N_15683,N_15095,N_14448);
and U15684 (N_15684,N_14949,N_15052);
xnor U15685 (N_15685,N_14885,N_15156);
or U15686 (N_15686,N_15106,N_15199);
or U15687 (N_15687,N_14698,N_15085);
and U15688 (N_15688,N_14565,N_15064);
nand U15689 (N_15689,N_14591,N_14660);
nand U15690 (N_15690,N_14904,N_14447);
nand U15691 (N_15691,N_14822,N_15177);
nor U15692 (N_15692,N_14559,N_14445);
xor U15693 (N_15693,N_14802,N_14429);
and U15694 (N_15694,N_14912,N_14502);
or U15695 (N_15695,N_14460,N_14815);
xor U15696 (N_15696,N_14777,N_14822);
nand U15697 (N_15697,N_15137,N_14561);
and U15698 (N_15698,N_14515,N_14708);
nand U15699 (N_15699,N_14743,N_15088);
nor U15700 (N_15700,N_14928,N_15062);
nand U15701 (N_15701,N_15092,N_14577);
or U15702 (N_15702,N_14654,N_15051);
xnor U15703 (N_15703,N_14429,N_14705);
nor U15704 (N_15704,N_14735,N_14498);
nor U15705 (N_15705,N_14655,N_14788);
and U15706 (N_15706,N_14726,N_14559);
nand U15707 (N_15707,N_14904,N_14918);
nand U15708 (N_15708,N_14955,N_14887);
xor U15709 (N_15709,N_14897,N_14792);
xnor U15710 (N_15710,N_14647,N_15002);
and U15711 (N_15711,N_14511,N_14433);
and U15712 (N_15712,N_15051,N_15094);
xnor U15713 (N_15713,N_15198,N_14683);
nand U15714 (N_15714,N_14562,N_14813);
or U15715 (N_15715,N_14656,N_15100);
xor U15716 (N_15716,N_15006,N_14453);
xor U15717 (N_15717,N_14433,N_14715);
xor U15718 (N_15718,N_14629,N_14705);
xor U15719 (N_15719,N_14585,N_14552);
nor U15720 (N_15720,N_15031,N_14595);
and U15721 (N_15721,N_15022,N_15047);
nor U15722 (N_15722,N_14750,N_14498);
and U15723 (N_15723,N_14720,N_14445);
nor U15724 (N_15724,N_14507,N_15193);
or U15725 (N_15725,N_14682,N_14542);
nand U15726 (N_15726,N_14854,N_14781);
xnor U15727 (N_15727,N_15119,N_14460);
nand U15728 (N_15728,N_15127,N_14473);
or U15729 (N_15729,N_14646,N_14450);
xnor U15730 (N_15730,N_14691,N_15061);
and U15731 (N_15731,N_14422,N_14975);
or U15732 (N_15732,N_15025,N_14724);
or U15733 (N_15733,N_14973,N_14911);
xnor U15734 (N_15734,N_14951,N_15191);
nor U15735 (N_15735,N_15006,N_15048);
or U15736 (N_15736,N_14479,N_15176);
xnor U15737 (N_15737,N_14919,N_14797);
xor U15738 (N_15738,N_14456,N_14509);
or U15739 (N_15739,N_14773,N_14817);
or U15740 (N_15740,N_14490,N_14494);
nor U15741 (N_15741,N_15157,N_14931);
nor U15742 (N_15742,N_14674,N_14952);
and U15743 (N_15743,N_15198,N_14891);
nand U15744 (N_15744,N_14483,N_15119);
or U15745 (N_15745,N_15117,N_14700);
xor U15746 (N_15746,N_14450,N_14527);
nor U15747 (N_15747,N_14439,N_14892);
xor U15748 (N_15748,N_14539,N_14529);
and U15749 (N_15749,N_14753,N_14944);
nand U15750 (N_15750,N_15136,N_14401);
nand U15751 (N_15751,N_14857,N_14796);
xor U15752 (N_15752,N_14599,N_15169);
nor U15753 (N_15753,N_14491,N_15071);
nand U15754 (N_15754,N_14685,N_15019);
xor U15755 (N_15755,N_14897,N_14893);
or U15756 (N_15756,N_15087,N_14944);
nor U15757 (N_15757,N_14811,N_14481);
nor U15758 (N_15758,N_14523,N_14692);
or U15759 (N_15759,N_14592,N_14840);
nor U15760 (N_15760,N_14834,N_14522);
or U15761 (N_15761,N_14774,N_14811);
xnor U15762 (N_15762,N_15024,N_15116);
and U15763 (N_15763,N_14896,N_14632);
or U15764 (N_15764,N_14474,N_15197);
nor U15765 (N_15765,N_15162,N_14616);
nor U15766 (N_15766,N_15070,N_14859);
and U15767 (N_15767,N_14903,N_14983);
or U15768 (N_15768,N_14412,N_14454);
xnor U15769 (N_15769,N_15093,N_14939);
xor U15770 (N_15770,N_14940,N_14435);
and U15771 (N_15771,N_14564,N_14948);
nand U15772 (N_15772,N_14699,N_14443);
nor U15773 (N_15773,N_14592,N_14496);
and U15774 (N_15774,N_14737,N_14720);
nor U15775 (N_15775,N_14610,N_15162);
nand U15776 (N_15776,N_14933,N_14430);
and U15777 (N_15777,N_15192,N_14728);
and U15778 (N_15778,N_15026,N_14745);
xnor U15779 (N_15779,N_14605,N_14423);
or U15780 (N_15780,N_14909,N_14850);
and U15781 (N_15781,N_14838,N_15195);
nor U15782 (N_15782,N_14570,N_14653);
and U15783 (N_15783,N_14680,N_14721);
nand U15784 (N_15784,N_14952,N_14676);
xnor U15785 (N_15785,N_14570,N_14713);
xor U15786 (N_15786,N_14855,N_14943);
xor U15787 (N_15787,N_14764,N_15170);
and U15788 (N_15788,N_14943,N_14622);
xor U15789 (N_15789,N_14714,N_14999);
and U15790 (N_15790,N_14947,N_14693);
xor U15791 (N_15791,N_14760,N_14910);
xor U15792 (N_15792,N_15009,N_14701);
nand U15793 (N_15793,N_14747,N_14664);
or U15794 (N_15794,N_14657,N_15035);
nand U15795 (N_15795,N_14933,N_14984);
or U15796 (N_15796,N_15175,N_14649);
nor U15797 (N_15797,N_15095,N_15098);
nor U15798 (N_15798,N_15155,N_14588);
nand U15799 (N_15799,N_14816,N_14677);
or U15800 (N_15800,N_14864,N_14551);
nand U15801 (N_15801,N_14768,N_15138);
and U15802 (N_15802,N_14624,N_14680);
nand U15803 (N_15803,N_15023,N_14618);
nor U15804 (N_15804,N_15108,N_14555);
xnor U15805 (N_15805,N_15013,N_14613);
nand U15806 (N_15806,N_15162,N_14501);
nor U15807 (N_15807,N_15176,N_14660);
and U15808 (N_15808,N_14527,N_14778);
nor U15809 (N_15809,N_14528,N_14839);
nor U15810 (N_15810,N_14905,N_14544);
nand U15811 (N_15811,N_14961,N_15174);
xnor U15812 (N_15812,N_14918,N_14468);
nor U15813 (N_15813,N_14670,N_15082);
nand U15814 (N_15814,N_14514,N_14652);
xor U15815 (N_15815,N_14473,N_15146);
nor U15816 (N_15816,N_14490,N_14943);
or U15817 (N_15817,N_14711,N_14487);
nand U15818 (N_15818,N_15186,N_14759);
and U15819 (N_15819,N_14875,N_14729);
nand U15820 (N_15820,N_14952,N_14629);
xnor U15821 (N_15821,N_14562,N_15016);
or U15822 (N_15822,N_14610,N_14627);
or U15823 (N_15823,N_14959,N_14856);
nand U15824 (N_15824,N_14775,N_14955);
and U15825 (N_15825,N_14507,N_15149);
nor U15826 (N_15826,N_15110,N_14987);
nand U15827 (N_15827,N_14665,N_14869);
nor U15828 (N_15828,N_14515,N_14517);
and U15829 (N_15829,N_14819,N_14562);
xnor U15830 (N_15830,N_14926,N_15189);
nor U15831 (N_15831,N_14998,N_14915);
nand U15832 (N_15832,N_14592,N_15081);
xor U15833 (N_15833,N_14758,N_14404);
or U15834 (N_15834,N_14418,N_14977);
and U15835 (N_15835,N_14915,N_15011);
xnor U15836 (N_15836,N_14994,N_14515);
and U15837 (N_15837,N_14660,N_14759);
nand U15838 (N_15838,N_14519,N_14441);
and U15839 (N_15839,N_14939,N_14555);
xor U15840 (N_15840,N_14995,N_14652);
xnor U15841 (N_15841,N_14730,N_14631);
or U15842 (N_15842,N_14956,N_15077);
nor U15843 (N_15843,N_14955,N_14604);
or U15844 (N_15844,N_14925,N_14514);
and U15845 (N_15845,N_14681,N_14611);
or U15846 (N_15846,N_14534,N_15189);
xor U15847 (N_15847,N_14672,N_14407);
or U15848 (N_15848,N_15034,N_14800);
and U15849 (N_15849,N_14631,N_14767);
xor U15850 (N_15850,N_15159,N_14850);
or U15851 (N_15851,N_15083,N_15131);
xor U15852 (N_15852,N_15009,N_15192);
and U15853 (N_15853,N_14965,N_14500);
nand U15854 (N_15854,N_14805,N_14416);
nand U15855 (N_15855,N_15170,N_15075);
nand U15856 (N_15856,N_15076,N_14544);
nor U15857 (N_15857,N_15050,N_14956);
xnor U15858 (N_15858,N_14703,N_14494);
nand U15859 (N_15859,N_15198,N_14782);
and U15860 (N_15860,N_14460,N_14911);
nor U15861 (N_15861,N_15109,N_15139);
or U15862 (N_15862,N_14638,N_14586);
nand U15863 (N_15863,N_15016,N_14508);
and U15864 (N_15864,N_14623,N_14989);
or U15865 (N_15865,N_14754,N_14529);
nand U15866 (N_15866,N_14566,N_14776);
nor U15867 (N_15867,N_14468,N_14981);
nor U15868 (N_15868,N_15064,N_14474);
and U15869 (N_15869,N_14594,N_14607);
and U15870 (N_15870,N_14476,N_14855);
xor U15871 (N_15871,N_15131,N_14847);
or U15872 (N_15872,N_14496,N_14558);
nand U15873 (N_15873,N_15110,N_14556);
or U15874 (N_15874,N_15187,N_14915);
nor U15875 (N_15875,N_14803,N_14632);
nor U15876 (N_15876,N_14821,N_14855);
nor U15877 (N_15877,N_14771,N_14678);
nor U15878 (N_15878,N_14637,N_15140);
nor U15879 (N_15879,N_14827,N_14572);
and U15880 (N_15880,N_15069,N_14730);
nor U15881 (N_15881,N_15069,N_14437);
nand U15882 (N_15882,N_14842,N_14714);
nand U15883 (N_15883,N_14673,N_14444);
nand U15884 (N_15884,N_14840,N_14963);
and U15885 (N_15885,N_14577,N_15161);
nor U15886 (N_15886,N_14616,N_14525);
nor U15887 (N_15887,N_14703,N_14882);
nand U15888 (N_15888,N_14856,N_14467);
xor U15889 (N_15889,N_14665,N_14825);
xor U15890 (N_15890,N_15174,N_14426);
or U15891 (N_15891,N_14533,N_15169);
nor U15892 (N_15892,N_14787,N_14438);
nand U15893 (N_15893,N_14718,N_14745);
nand U15894 (N_15894,N_15174,N_14837);
xnor U15895 (N_15895,N_14453,N_14657);
nand U15896 (N_15896,N_14438,N_14922);
or U15897 (N_15897,N_14797,N_14714);
nor U15898 (N_15898,N_14633,N_15100);
or U15899 (N_15899,N_14574,N_15022);
and U15900 (N_15900,N_14512,N_14536);
xor U15901 (N_15901,N_14994,N_14742);
nand U15902 (N_15902,N_14557,N_14805);
and U15903 (N_15903,N_15153,N_15069);
or U15904 (N_15904,N_14773,N_15111);
and U15905 (N_15905,N_14905,N_14799);
xnor U15906 (N_15906,N_14738,N_14627);
xnor U15907 (N_15907,N_15047,N_15019);
nand U15908 (N_15908,N_14820,N_14482);
nand U15909 (N_15909,N_15071,N_15019);
xnor U15910 (N_15910,N_14775,N_15064);
and U15911 (N_15911,N_14891,N_14852);
xor U15912 (N_15912,N_15096,N_14803);
nor U15913 (N_15913,N_14439,N_14613);
nand U15914 (N_15914,N_14879,N_14966);
and U15915 (N_15915,N_14652,N_15150);
and U15916 (N_15916,N_15170,N_14784);
and U15917 (N_15917,N_14520,N_15018);
or U15918 (N_15918,N_15011,N_14835);
xor U15919 (N_15919,N_15036,N_14579);
or U15920 (N_15920,N_14868,N_14738);
nand U15921 (N_15921,N_14704,N_14865);
xor U15922 (N_15922,N_14634,N_14492);
nor U15923 (N_15923,N_14648,N_14836);
nor U15924 (N_15924,N_14504,N_15031);
nor U15925 (N_15925,N_14919,N_15095);
or U15926 (N_15926,N_14458,N_14930);
or U15927 (N_15927,N_14411,N_15016);
or U15928 (N_15928,N_14550,N_14978);
xnor U15929 (N_15929,N_14782,N_14631);
nand U15930 (N_15930,N_14612,N_15167);
and U15931 (N_15931,N_14810,N_14805);
nand U15932 (N_15932,N_14600,N_14870);
xor U15933 (N_15933,N_14680,N_14410);
xor U15934 (N_15934,N_14864,N_14618);
nor U15935 (N_15935,N_14664,N_14835);
xnor U15936 (N_15936,N_14416,N_14866);
and U15937 (N_15937,N_14987,N_14651);
nand U15938 (N_15938,N_14851,N_14506);
nand U15939 (N_15939,N_14826,N_15196);
and U15940 (N_15940,N_14588,N_14459);
nor U15941 (N_15941,N_14490,N_14910);
nor U15942 (N_15942,N_15182,N_14897);
and U15943 (N_15943,N_14906,N_14843);
and U15944 (N_15944,N_15130,N_15074);
and U15945 (N_15945,N_14564,N_14592);
nand U15946 (N_15946,N_15156,N_14785);
xnor U15947 (N_15947,N_14667,N_15065);
or U15948 (N_15948,N_14664,N_14869);
nand U15949 (N_15949,N_14921,N_14516);
and U15950 (N_15950,N_15170,N_14813);
nor U15951 (N_15951,N_14848,N_14759);
and U15952 (N_15952,N_14734,N_15060);
or U15953 (N_15953,N_14681,N_14418);
nor U15954 (N_15954,N_14822,N_14935);
and U15955 (N_15955,N_15032,N_14858);
and U15956 (N_15956,N_14420,N_14937);
xnor U15957 (N_15957,N_14698,N_14475);
nand U15958 (N_15958,N_14594,N_15039);
xor U15959 (N_15959,N_14463,N_14431);
nor U15960 (N_15960,N_15154,N_14857);
nand U15961 (N_15961,N_14622,N_15112);
xor U15962 (N_15962,N_15145,N_14901);
xor U15963 (N_15963,N_14437,N_15090);
or U15964 (N_15964,N_14593,N_15049);
xnor U15965 (N_15965,N_14872,N_14444);
or U15966 (N_15966,N_14602,N_15067);
nor U15967 (N_15967,N_14850,N_14841);
and U15968 (N_15968,N_15186,N_14670);
or U15969 (N_15969,N_15007,N_14734);
xnor U15970 (N_15970,N_14867,N_15173);
nand U15971 (N_15971,N_14867,N_14785);
and U15972 (N_15972,N_14876,N_14630);
and U15973 (N_15973,N_14762,N_14804);
and U15974 (N_15974,N_15112,N_14880);
nor U15975 (N_15975,N_15098,N_14528);
nor U15976 (N_15976,N_14966,N_14510);
nor U15977 (N_15977,N_15112,N_14569);
xor U15978 (N_15978,N_14439,N_15154);
and U15979 (N_15979,N_15007,N_14893);
and U15980 (N_15980,N_14858,N_14843);
or U15981 (N_15981,N_14680,N_15115);
xnor U15982 (N_15982,N_14973,N_15148);
nor U15983 (N_15983,N_15008,N_14536);
or U15984 (N_15984,N_14412,N_14820);
nor U15985 (N_15985,N_14494,N_15047);
nor U15986 (N_15986,N_14998,N_14500);
nor U15987 (N_15987,N_14961,N_14670);
and U15988 (N_15988,N_14457,N_15069);
and U15989 (N_15989,N_14905,N_14698);
xor U15990 (N_15990,N_14618,N_15137);
xnor U15991 (N_15991,N_14412,N_15053);
xor U15992 (N_15992,N_14684,N_15016);
or U15993 (N_15993,N_14932,N_15091);
nor U15994 (N_15994,N_15026,N_14773);
xor U15995 (N_15995,N_14920,N_15007);
xor U15996 (N_15996,N_14457,N_14800);
xor U15997 (N_15997,N_15056,N_15148);
or U15998 (N_15998,N_14695,N_14897);
xnor U15999 (N_15999,N_14957,N_14674);
nor U16000 (N_16000,N_15490,N_15434);
and U16001 (N_16001,N_15921,N_15429);
nor U16002 (N_16002,N_15536,N_15478);
nor U16003 (N_16003,N_15769,N_15849);
nor U16004 (N_16004,N_15621,N_15427);
and U16005 (N_16005,N_15602,N_15263);
nand U16006 (N_16006,N_15311,N_15458);
xor U16007 (N_16007,N_15312,N_15895);
or U16008 (N_16008,N_15467,N_15858);
xnor U16009 (N_16009,N_15278,N_15357);
nand U16010 (N_16010,N_15564,N_15724);
nand U16011 (N_16011,N_15876,N_15615);
nor U16012 (N_16012,N_15364,N_15674);
or U16013 (N_16013,N_15843,N_15552);
or U16014 (N_16014,N_15409,N_15725);
or U16015 (N_16015,N_15595,N_15786);
nand U16016 (N_16016,N_15599,N_15760);
or U16017 (N_16017,N_15874,N_15879);
and U16018 (N_16018,N_15231,N_15282);
nor U16019 (N_16019,N_15672,N_15625);
xnor U16020 (N_16020,N_15320,N_15776);
nand U16021 (N_16021,N_15562,N_15783);
xnor U16022 (N_16022,N_15986,N_15648);
xor U16023 (N_16023,N_15697,N_15577);
or U16024 (N_16024,N_15811,N_15711);
and U16025 (N_16025,N_15442,N_15293);
xnor U16026 (N_16026,N_15779,N_15670);
xor U16027 (N_16027,N_15369,N_15271);
or U16028 (N_16028,N_15499,N_15385);
or U16029 (N_16029,N_15937,N_15634);
xor U16030 (N_16030,N_15780,N_15756);
or U16031 (N_16031,N_15754,N_15448);
or U16032 (N_16032,N_15775,N_15923);
and U16033 (N_16033,N_15790,N_15755);
and U16034 (N_16034,N_15911,N_15534);
nor U16035 (N_16035,N_15353,N_15864);
nor U16036 (N_16036,N_15208,N_15985);
nand U16037 (N_16037,N_15390,N_15688);
or U16038 (N_16038,N_15306,N_15463);
nor U16039 (N_16039,N_15245,N_15881);
or U16040 (N_16040,N_15363,N_15408);
nand U16041 (N_16041,N_15421,N_15276);
and U16042 (N_16042,N_15514,N_15383);
and U16043 (N_16043,N_15547,N_15909);
xor U16044 (N_16044,N_15557,N_15594);
nand U16045 (N_16045,N_15791,N_15492);
nand U16046 (N_16046,N_15651,N_15638);
or U16047 (N_16047,N_15800,N_15927);
nor U16048 (N_16048,N_15804,N_15329);
nand U16049 (N_16049,N_15834,N_15546);
nand U16050 (N_16050,N_15907,N_15298);
nor U16051 (N_16051,N_15323,N_15220);
and U16052 (N_16052,N_15686,N_15246);
nand U16053 (N_16053,N_15657,N_15758);
nor U16054 (N_16054,N_15314,N_15336);
nand U16055 (N_16055,N_15677,N_15331);
xor U16056 (N_16056,N_15974,N_15232);
xor U16057 (N_16057,N_15846,N_15238);
and U16058 (N_16058,N_15867,N_15799);
xnor U16059 (N_16059,N_15721,N_15788);
and U16060 (N_16060,N_15713,N_15432);
and U16061 (N_16061,N_15468,N_15452);
and U16062 (N_16062,N_15344,N_15793);
and U16063 (N_16063,N_15837,N_15877);
nand U16064 (N_16064,N_15759,N_15588);
and U16065 (N_16065,N_15341,N_15700);
xnor U16066 (N_16066,N_15257,N_15701);
xor U16067 (N_16067,N_15568,N_15705);
xnor U16068 (N_16068,N_15582,N_15764);
nor U16069 (N_16069,N_15498,N_15723);
nor U16070 (N_16070,N_15941,N_15641);
nor U16071 (N_16071,N_15515,N_15862);
and U16072 (N_16072,N_15838,N_15805);
nand U16073 (N_16073,N_15847,N_15614);
nor U16074 (N_16074,N_15503,N_15976);
nand U16075 (N_16075,N_15887,N_15461);
nor U16076 (N_16076,N_15603,N_15506);
xnor U16077 (N_16077,N_15241,N_15367);
xnor U16078 (N_16078,N_15339,N_15980);
nor U16079 (N_16079,N_15437,N_15494);
xnor U16080 (N_16080,N_15496,N_15617);
nand U16081 (N_16081,N_15281,N_15845);
or U16082 (N_16082,N_15944,N_15646);
nand U16083 (N_16083,N_15317,N_15857);
nand U16084 (N_16084,N_15354,N_15925);
nor U16085 (N_16085,N_15290,N_15253);
nor U16086 (N_16086,N_15806,N_15850);
nand U16087 (N_16087,N_15528,N_15213);
and U16088 (N_16088,N_15508,N_15237);
xor U16089 (N_16089,N_15728,N_15678);
or U16090 (N_16090,N_15495,N_15510);
nor U16091 (N_16091,N_15493,N_15532);
nand U16092 (N_16092,N_15280,N_15897);
nand U16093 (N_16093,N_15939,N_15908);
or U16094 (N_16094,N_15295,N_15457);
and U16095 (N_16095,N_15446,N_15596);
and U16096 (N_16096,N_15481,N_15613);
and U16097 (N_16097,N_15797,N_15265);
nor U16098 (N_16098,N_15914,N_15450);
xor U16099 (N_16099,N_15900,N_15635);
nor U16100 (N_16100,N_15992,N_15853);
nand U16101 (N_16101,N_15420,N_15441);
and U16102 (N_16102,N_15894,N_15299);
or U16103 (N_16103,N_15979,N_15398);
and U16104 (N_16104,N_15233,N_15440);
nand U16105 (N_16105,N_15655,N_15752);
and U16106 (N_16106,N_15476,N_15663);
xnor U16107 (N_16107,N_15844,N_15541);
nand U16108 (N_16108,N_15659,N_15491);
nor U16109 (N_16109,N_15501,N_15951);
nand U16110 (N_16110,N_15570,N_15839);
xor U16111 (N_16111,N_15465,N_15773);
nand U16112 (N_16112,N_15535,N_15611);
xnor U16113 (N_16113,N_15928,N_15487);
nand U16114 (N_16114,N_15789,N_15716);
nor U16115 (N_16115,N_15229,N_15886);
nand U16116 (N_16116,N_15328,N_15763);
nand U16117 (N_16117,N_15652,N_15955);
and U16118 (N_16118,N_15903,N_15256);
nor U16119 (N_16119,N_15419,N_15227);
and U16120 (N_16120,N_15393,N_15627);
nand U16121 (N_16121,N_15386,N_15466);
xnor U16122 (N_16122,N_15718,N_15737);
nand U16123 (N_16123,N_15968,N_15203);
and U16124 (N_16124,N_15435,N_15949);
nand U16125 (N_16125,N_15661,N_15702);
nor U16126 (N_16126,N_15272,N_15214);
nand U16127 (N_16127,N_15527,N_15379);
nand U16128 (N_16128,N_15916,N_15860);
xor U16129 (N_16129,N_15294,N_15943);
or U16130 (N_16130,N_15489,N_15308);
and U16131 (N_16131,N_15606,N_15592);
nand U16132 (N_16132,N_15973,N_15774);
or U16133 (N_16133,N_15848,N_15926);
and U16134 (N_16134,N_15544,N_15802);
nand U16135 (N_16135,N_15956,N_15778);
nor U16136 (N_16136,N_15445,N_15486);
xor U16137 (N_16137,N_15946,N_15745);
or U16138 (N_16138,N_15566,N_15443);
nor U16139 (N_16139,N_15283,N_15572);
nor U16140 (N_16140,N_15488,N_15972);
nand U16141 (N_16141,N_15731,N_15313);
and U16142 (N_16142,N_15275,N_15706);
nand U16143 (N_16143,N_15977,N_15746);
and U16144 (N_16144,N_15223,N_15736);
nor U16145 (N_16145,N_15694,N_15975);
or U16146 (N_16146,N_15219,N_15819);
nor U16147 (N_16147,N_15719,N_15551);
nand U16148 (N_16148,N_15966,N_15247);
and U16149 (N_16149,N_15243,N_15822);
xor U16150 (N_16150,N_15264,N_15391);
or U16151 (N_16151,N_15593,N_15342);
nor U16152 (N_16152,N_15349,N_15416);
and U16153 (N_16153,N_15631,N_15988);
or U16154 (N_16154,N_15689,N_15206);
or U16155 (N_16155,N_15423,N_15337);
xnor U16156 (N_16156,N_15543,N_15201);
and U16157 (N_16157,N_15970,N_15259);
and U16158 (N_16158,N_15809,N_15549);
xor U16159 (N_16159,N_15865,N_15675);
xnor U16160 (N_16160,N_15965,N_15827);
or U16161 (N_16161,N_15803,N_15270);
and U16162 (N_16162,N_15384,N_15394);
xnor U16163 (N_16163,N_15859,N_15696);
or U16164 (N_16164,N_15401,N_15642);
nand U16165 (N_16165,N_15600,N_15296);
nor U16166 (N_16166,N_15581,N_15338);
nor U16167 (N_16167,N_15679,N_15509);
or U16168 (N_16168,N_15669,N_15738);
xor U16169 (N_16169,N_15643,N_15917);
and U16170 (N_16170,N_15332,N_15340);
and U16171 (N_16171,N_15953,N_15878);
nand U16172 (N_16172,N_15998,N_15691);
nor U16173 (N_16173,N_15832,N_15812);
xnor U16174 (N_16174,N_15473,N_15560);
nor U16175 (N_16175,N_15469,N_15934);
nand U16176 (N_16176,N_15919,N_15649);
or U16177 (N_16177,N_15483,N_15211);
nor U16178 (N_16178,N_15396,N_15781);
nor U16179 (N_16179,N_15359,N_15708);
or U16180 (N_16180,N_15471,N_15334);
and U16181 (N_16181,N_15958,N_15905);
or U16182 (N_16182,N_15815,N_15870);
nand U16183 (N_16183,N_15930,N_15413);
and U16184 (N_16184,N_15288,N_15795);
xor U16185 (N_16185,N_15831,N_15727);
nor U16186 (N_16186,N_15439,N_15428);
nor U16187 (N_16187,N_15890,N_15348);
nor U16188 (N_16188,N_15584,N_15964);
nand U16189 (N_16189,N_15565,N_15714);
or U16190 (N_16190,N_15747,N_15880);
xnor U16191 (N_16191,N_15202,N_15963);
xnor U16192 (N_16192,N_15768,N_15215);
nor U16193 (N_16193,N_15355,N_15269);
nand U16194 (N_16194,N_15325,N_15404);
xor U16195 (N_16195,N_15816,N_15381);
xor U16196 (N_16196,N_15589,N_15371);
nor U16197 (N_16197,N_15410,N_15852);
xor U16198 (N_16198,N_15531,N_15580);
and U16199 (N_16199,N_15388,N_15889);
or U16200 (N_16200,N_15695,N_15268);
nand U16201 (N_16201,N_15931,N_15239);
and U16202 (N_16202,N_15961,N_15733);
or U16203 (N_16203,N_15628,N_15835);
and U16204 (N_16204,N_15550,N_15912);
and U16205 (N_16205,N_15633,N_15578);
nand U16206 (N_16206,N_15885,N_15533);
or U16207 (N_16207,N_15472,N_15922);
and U16208 (N_16208,N_15662,N_15983);
and U16209 (N_16209,N_15374,N_15569);
nor U16210 (N_16210,N_15632,N_15740);
nand U16211 (N_16211,N_15684,N_15365);
nand U16212 (N_16212,N_15540,N_15345);
or U16213 (N_16213,N_15598,N_15400);
or U16214 (N_16214,N_15671,N_15757);
and U16215 (N_16215,N_15654,N_15292);
nand U16216 (N_16216,N_15967,N_15414);
xnor U16217 (N_16217,N_15475,N_15525);
nand U16218 (N_16218,N_15729,N_15987);
or U16219 (N_16219,N_15235,N_15782);
or U16220 (N_16220,N_15717,N_15297);
and U16221 (N_16221,N_15884,N_15431);
and U16222 (N_16222,N_15346,N_15573);
nor U16223 (N_16223,N_15751,N_15563);
nand U16224 (N_16224,N_15530,N_15990);
nand U16225 (N_16225,N_15392,N_15318);
nor U16226 (N_16226,N_15521,N_15861);
or U16227 (N_16227,N_15637,N_15750);
nand U16228 (N_16228,N_15277,N_15918);
or U16229 (N_16229,N_15796,N_15403);
or U16230 (N_16230,N_15542,N_15397);
xor U16231 (N_16231,N_15376,N_15366);
or U16232 (N_16232,N_15553,N_15712);
nor U16233 (N_16233,N_15624,N_15230);
xor U16234 (N_16234,N_15667,N_15330);
or U16235 (N_16235,N_15869,N_15555);
xnor U16236 (N_16236,N_15749,N_15996);
nor U16237 (N_16237,N_15537,N_15315);
and U16238 (N_16238,N_15629,N_15682);
or U16239 (N_16239,N_15842,N_15971);
nand U16240 (N_16240,N_15978,N_15303);
nor U16241 (N_16241,N_15673,N_15698);
or U16242 (N_16242,N_15484,N_15607);
or U16243 (N_16243,N_15828,N_15244);
xor U16244 (N_16244,N_15212,N_15952);
and U16245 (N_16245,N_15326,N_15455);
xor U16246 (N_16246,N_15482,N_15236);
xnor U16247 (N_16247,N_15902,N_15856);
or U16248 (N_16248,N_15609,N_15507);
xor U16249 (N_16249,N_15561,N_15430);
nand U16250 (N_16250,N_15658,N_15873);
and U16251 (N_16251,N_15204,N_15205);
or U16252 (N_16252,N_15449,N_15304);
xnor U16253 (N_16253,N_15833,N_15300);
or U16254 (N_16254,N_15875,N_15447);
or U16255 (N_16255,N_15222,N_15456);
nand U16256 (N_16256,N_15305,N_15411);
xor U16257 (N_16257,N_15480,N_15929);
and U16258 (N_16258,N_15785,N_15993);
nor U16259 (N_16259,N_15765,N_15310);
nand U16260 (N_16260,N_15444,N_15517);
xor U16261 (N_16261,N_15368,N_15459);
xnor U16262 (N_16262,N_15512,N_15734);
and U16263 (N_16263,N_15210,N_15591);
nand U16264 (N_16264,N_15732,N_15286);
or U16265 (N_16265,N_15520,N_15370);
and U16266 (N_16266,N_15777,N_15935);
and U16267 (N_16267,N_15302,N_15529);
or U16268 (N_16268,N_15739,N_15741);
or U16269 (N_16269,N_15947,N_15618);
nor U16270 (N_16270,N_15335,N_15377);
nand U16271 (N_16271,N_15619,N_15343);
nand U16272 (N_16272,N_15722,N_15415);
and U16273 (N_16273,N_15539,N_15575);
or U16274 (N_16274,N_15989,N_15771);
nand U16275 (N_16275,N_15920,N_15319);
and U16276 (N_16276,N_15378,N_15735);
and U16277 (N_16277,N_15685,N_15620);
nor U16278 (N_16278,N_15524,N_15321);
nand U16279 (N_16279,N_15226,N_15882);
and U16280 (N_16280,N_15267,N_15587);
or U16281 (N_16281,N_15893,N_15585);
xnor U16282 (N_16282,N_15801,N_15762);
and U16283 (N_16283,N_15942,N_15358);
nor U16284 (N_16284,N_15502,N_15548);
or U16285 (N_16285,N_15823,N_15709);
or U16286 (N_16286,N_15406,N_15207);
or U16287 (N_16287,N_15352,N_15266);
nor U16288 (N_16288,N_15422,N_15938);
xnor U16289 (N_16289,N_15761,N_15924);
nand U16290 (N_16290,N_15913,N_15704);
nand U16291 (N_16291,N_15854,N_15960);
and U16292 (N_16292,N_15579,N_15676);
and U16293 (N_16293,N_15307,N_15453);
and U16294 (N_16294,N_15950,N_15571);
and U16295 (N_16295,N_15871,N_15687);
nand U16296 (N_16296,N_15683,N_15558);
and U16297 (N_16297,N_15242,N_15792);
xor U16298 (N_16298,N_15821,N_15898);
or U16299 (N_16299,N_15418,N_15770);
xor U16300 (N_16300,N_15690,N_15892);
xor U16301 (N_16301,N_15840,N_15720);
nand U16302 (N_16302,N_15896,N_15604);
xnor U16303 (N_16303,N_15753,N_15258);
or U16304 (N_16304,N_15991,N_15824);
nand U16305 (N_16305,N_15522,N_15375);
or U16306 (N_16306,N_15647,N_15818);
nand U16307 (N_16307,N_15820,N_15608);
nor U16308 (N_16308,N_15807,N_15436);
nand U16309 (N_16309,N_15622,N_15464);
or U16310 (N_16310,N_15645,N_15954);
xor U16311 (N_16311,N_15680,N_15863);
nor U16312 (N_16312,N_15224,N_15526);
nor U16313 (N_16313,N_15590,N_15324);
nor U16314 (N_16314,N_15945,N_15399);
or U16315 (N_16315,N_15612,N_15250);
nor U16316 (N_16316,N_15656,N_15743);
and U16317 (N_16317,N_15730,N_15855);
or U16318 (N_16318,N_15322,N_15511);
and U16319 (N_16319,N_15969,N_15836);
xnor U16320 (N_16320,N_15451,N_15699);
or U16321 (N_16321,N_15668,N_15813);
nor U16322 (N_16322,N_15999,N_15382);
nor U16323 (N_16323,N_15829,N_15910);
or U16324 (N_16324,N_15940,N_15915);
xnor U16325 (N_16325,N_15742,N_15426);
xnor U16326 (N_16326,N_15601,N_15538);
xor U16327 (N_16327,N_15218,N_15362);
nand U16328 (N_16328,N_15356,N_15200);
and U16329 (N_16329,N_15479,N_15767);
and U16330 (N_16330,N_15518,N_15660);
nand U16331 (N_16331,N_15994,N_15744);
nor U16332 (N_16332,N_15545,N_15361);
and U16333 (N_16333,N_15650,N_15932);
nand U16334 (N_16334,N_15957,N_15872);
xnor U16335 (N_16335,N_15309,N_15389);
xnor U16336 (N_16336,N_15639,N_15891);
and U16337 (N_16337,N_15485,N_15395);
nand U16338 (N_16338,N_15273,N_15424);
and U16339 (N_16339,N_15826,N_15327);
xor U16340 (N_16340,N_15692,N_15640);
xnor U16341 (N_16341,N_15787,N_15347);
xnor U16342 (N_16342,N_15351,N_15810);
and U16343 (N_16343,N_15981,N_15523);
and U16344 (N_16344,N_15626,N_15438);
or U16345 (N_16345,N_15715,N_15221);
xnor U16346 (N_16346,N_15681,N_15653);
or U16347 (N_16347,N_15262,N_15372);
or U16348 (N_16348,N_15405,N_15301);
nor U16349 (N_16349,N_15610,N_15567);
nand U16350 (N_16350,N_15784,N_15707);
or U16351 (N_16351,N_15808,N_15576);
nor U16352 (N_16352,N_15556,N_15462);
nand U16353 (N_16353,N_15425,N_15516);
or U16354 (N_16354,N_15586,N_15583);
and U16355 (N_16355,N_15825,N_15841);
or U16356 (N_16356,N_15228,N_15623);
xnor U16357 (N_16357,N_15817,N_15666);
and U16358 (N_16358,N_15962,N_15559);
nand U16359 (N_16359,N_15664,N_15255);
xor U16360 (N_16360,N_15693,N_15497);
nand U16361 (N_16361,N_15251,N_15794);
xnor U16362 (N_16362,N_15748,N_15387);
nor U16363 (N_16363,N_15261,N_15726);
nor U16364 (N_16364,N_15830,N_15616);
nor U16365 (N_16365,N_15407,N_15982);
xor U16366 (N_16366,N_15316,N_15703);
nand U16367 (N_16367,N_15630,N_15766);
nor U16368 (N_16368,N_15460,N_15225);
or U16369 (N_16369,N_15901,N_15995);
nor U16370 (N_16370,N_15883,N_15254);
nor U16371 (N_16371,N_15868,N_15710);
xnor U16372 (N_16372,N_15904,N_15933);
nand U16373 (N_16373,N_15888,N_15997);
nand U16374 (N_16374,N_15216,N_15513);
nand U16375 (N_16375,N_15500,N_15380);
or U16376 (N_16376,N_15412,N_15289);
or U16377 (N_16377,N_15984,N_15249);
or U16378 (N_16378,N_15454,N_15798);
nor U16379 (N_16379,N_15285,N_15252);
xnor U16380 (N_16380,N_15279,N_15284);
and U16381 (N_16381,N_15665,N_15209);
and U16382 (N_16382,N_15240,N_15899);
xor U16383 (N_16383,N_15360,N_15866);
or U16384 (N_16384,N_15636,N_15519);
or U16385 (N_16385,N_15948,N_15959);
nand U16386 (N_16386,N_15851,N_15287);
nand U16387 (N_16387,N_15477,N_15260);
nand U16388 (N_16388,N_15417,N_15936);
nor U16389 (N_16389,N_15217,N_15574);
and U16390 (N_16390,N_15597,N_15505);
or U16391 (N_16391,N_15474,N_15333);
nand U16392 (N_16392,N_15644,N_15605);
nand U16393 (N_16393,N_15373,N_15274);
nor U16394 (N_16394,N_15433,N_15504);
nor U16395 (N_16395,N_15248,N_15470);
and U16396 (N_16396,N_15350,N_15291);
nand U16397 (N_16397,N_15814,N_15402);
xnor U16398 (N_16398,N_15234,N_15554);
or U16399 (N_16399,N_15772,N_15906);
nor U16400 (N_16400,N_15870,N_15267);
nand U16401 (N_16401,N_15653,N_15582);
nor U16402 (N_16402,N_15247,N_15239);
nor U16403 (N_16403,N_15826,N_15296);
nand U16404 (N_16404,N_15621,N_15223);
xnor U16405 (N_16405,N_15227,N_15706);
nor U16406 (N_16406,N_15789,N_15719);
nand U16407 (N_16407,N_15462,N_15975);
and U16408 (N_16408,N_15864,N_15711);
and U16409 (N_16409,N_15342,N_15389);
nor U16410 (N_16410,N_15392,N_15577);
or U16411 (N_16411,N_15634,N_15695);
nor U16412 (N_16412,N_15449,N_15232);
nand U16413 (N_16413,N_15416,N_15783);
nor U16414 (N_16414,N_15326,N_15424);
nor U16415 (N_16415,N_15488,N_15573);
and U16416 (N_16416,N_15506,N_15358);
nand U16417 (N_16417,N_15637,N_15685);
nor U16418 (N_16418,N_15581,N_15232);
and U16419 (N_16419,N_15463,N_15885);
or U16420 (N_16420,N_15236,N_15226);
nand U16421 (N_16421,N_15655,N_15606);
and U16422 (N_16422,N_15740,N_15589);
xor U16423 (N_16423,N_15999,N_15433);
and U16424 (N_16424,N_15285,N_15971);
xnor U16425 (N_16425,N_15246,N_15454);
nand U16426 (N_16426,N_15658,N_15989);
xnor U16427 (N_16427,N_15299,N_15308);
or U16428 (N_16428,N_15236,N_15749);
nor U16429 (N_16429,N_15816,N_15497);
xor U16430 (N_16430,N_15916,N_15333);
nor U16431 (N_16431,N_15669,N_15330);
and U16432 (N_16432,N_15664,N_15485);
or U16433 (N_16433,N_15534,N_15593);
nand U16434 (N_16434,N_15323,N_15719);
nor U16435 (N_16435,N_15840,N_15302);
nand U16436 (N_16436,N_15857,N_15593);
xnor U16437 (N_16437,N_15206,N_15344);
nand U16438 (N_16438,N_15739,N_15489);
nand U16439 (N_16439,N_15495,N_15743);
xnor U16440 (N_16440,N_15938,N_15580);
nand U16441 (N_16441,N_15251,N_15493);
or U16442 (N_16442,N_15243,N_15294);
nand U16443 (N_16443,N_15859,N_15620);
nor U16444 (N_16444,N_15693,N_15954);
or U16445 (N_16445,N_15399,N_15230);
or U16446 (N_16446,N_15907,N_15658);
and U16447 (N_16447,N_15701,N_15377);
xor U16448 (N_16448,N_15959,N_15424);
nand U16449 (N_16449,N_15892,N_15920);
and U16450 (N_16450,N_15267,N_15687);
xor U16451 (N_16451,N_15251,N_15376);
xor U16452 (N_16452,N_15940,N_15936);
xnor U16453 (N_16453,N_15932,N_15894);
and U16454 (N_16454,N_15552,N_15404);
nand U16455 (N_16455,N_15301,N_15816);
nand U16456 (N_16456,N_15667,N_15293);
xnor U16457 (N_16457,N_15384,N_15454);
nor U16458 (N_16458,N_15899,N_15610);
xor U16459 (N_16459,N_15341,N_15442);
nor U16460 (N_16460,N_15906,N_15872);
and U16461 (N_16461,N_15332,N_15603);
nand U16462 (N_16462,N_15708,N_15580);
nand U16463 (N_16463,N_15733,N_15992);
nand U16464 (N_16464,N_15557,N_15930);
xor U16465 (N_16465,N_15475,N_15496);
nand U16466 (N_16466,N_15708,N_15805);
and U16467 (N_16467,N_15828,N_15747);
xor U16468 (N_16468,N_15205,N_15547);
and U16469 (N_16469,N_15606,N_15304);
nor U16470 (N_16470,N_15935,N_15420);
xnor U16471 (N_16471,N_15597,N_15744);
nand U16472 (N_16472,N_15467,N_15826);
or U16473 (N_16473,N_15737,N_15860);
and U16474 (N_16474,N_15623,N_15535);
or U16475 (N_16475,N_15371,N_15767);
nor U16476 (N_16476,N_15273,N_15737);
and U16477 (N_16477,N_15380,N_15483);
nor U16478 (N_16478,N_15722,N_15395);
or U16479 (N_16479,N_15730,N_15504);
and U16480 (N_16480,N_15327,N_15246);
nand U16481 (N_16481,N_15591,N_15213);
xnor U16482 (N_16482,N_15339,N_15321);
xnor U16483 (N_16483,N_15946,N_15802);
or U16484 (N_16484,N_15255,N_15332);
nand U16485 (N_16485,N_15642,N_15282);
or U16486 (N_16486,N_15365,N_15988);
nor U16487 (N_16487,N_15635,N_15545);
nor U16488 (N_16488,N_15569,N_15329);
and U16489 (N_16489,N_15253,N_15791);
and U16490 (N_16490,N_15848,N_15551);
and U16491 (N_16491,N_15272,N_15488);
and U16492 (N_16492,N_15569,N_15764);
and U16493 (N_16493,N_15844,N_15498);
nand U16494 (N_16494,N_15530,N_15446);
or U16495 (N_16495,N_15769,N_15938);
and U16496 (N_16496,N_15639,N_15520);
or U16497 (N_16497,N_15491,N_15886);
nor U16498 (N_16498,N_15442,N_15995);
nor U16499 (N_16499,N_15217,N_15311);
or U16500 (N_16500,N_15264,N_15325);
xnor U16501 (N_16501,N_15863,N_15990);
nand U16502 (N_16502,N_15505,N_15315);
nor U16503 (N_16503,N_15684,N_15560);
xnor U16504 (N_16504,N_15962,N_15589);
nor U16505 (N_16505,N_15762,N_15396);
or U16506 (N_16506,N_15368,N_15694);
nand U16507 (N_16507,N_15481,N_15928);
xnor U16508 (N_16508,N_15711,N_15446);
xnor U16509 (N_16509,N_15807,N_15875);
or U16510 (N_16510,N_15914,N_15746);
or U16511 (N_16511,N_15401,N_15971);
xnor U16512 (N_16512,N_15342,N_15425);
nand U16513 (N_16513,N_15497,N_15907);
or U16514 (N_16514,N_15632,N_15244);
and U16515 (N_16515,N_15838,N_15430);
and U16516 (N_16516,N_15321,N_15724);
nand U16517 (N_16517,N_15819,N_15644);
xor U16518 (N_16518,N_15654,N_15718);
nor U16519 (N_16519,N_15594,N_15746);
nand U16520 (N_16520,N_15202,N_15978);
or U16521 (N_16521,N_15227,N_15255);
or U16522 (N_16522,N_15638,N_15664);
and U16523 (N_16523,N_15976,N_15934);
or U16524 (N_16524,N_15796,N_15528);
or U16525 (N_16525,N_15450,N_15540);
or U16526 (N_16526,N_15637,N_15456);
or U16527 (N_16527,N_15952,N_15705);
xor U16528 (N_16528,N_15423,N_15305);
nand U16529 (N_16529,N_15715,N_15763);
xor U16530 (N_16530,N_15405,N_15695);
and U16531 (N_16531,N_15479,N_15317);
nand U16532 (N_16532,N_15938,N_15202);
nor U16533 (N_16533,N_15205,N_15434);
nand U16534 (N_16534,N_15969,N_15415);
and U16535 (N_16535,N_15933,N_15881);
nand U16536 (N_16536,N_15861,N_15776);
and U16537 (N_16537,N_15583,N_15756);
xor U16538 (N_16538,N_15931,N_15785);
and U16539 (N_16539,N_15352,N_15970);
nand U16540 (N_16540,N_15887,N_15300);
or U16541 (N_16541,N_15675,N_15289);
nor U16542 (N_16542,N_15628,N_15251);
and U16543 (N_16543,N_15410,N_15445);
nand U16544 (N_16544,N_15883,N_15786);
xor U16545 (N_16545,N_15818,N_15239);
or U16546 (N_16546,N_15781,N_15412);
or U16547 (N_16547,N_15717,N_15933);
and U16548 (N_16548,N_15711,N_15674);
or U16549 (N_16549,N_15272,N_15812);
nor U16550 (N_16550,N_15792,N_15473);
nand U16551 (N_16551,N_15920,N_15568);
nand U16552 (N_16552,N_15421,N_15924);
or U16553 (N_16553,N_15955,N_15530);
xor U16554 (N_16554,N_15628,N_15503);
xnor U16555 (N_16555,N_15470,N_15899);
and U16556 (N_16556,N_15464,N_15627);
xor U16557 (N_16557,N_15970,N_15832);
nor U16558 (N_16558,N_15393,N_15908);
and U16559 (N_16559,N_15665,N_15563);
nor U16560 (N_16560,N_15886,N_15665);
nor U16561 (N_16561,N_15439,N_15317);
and U16562 (N_16562,N_15594,N_15914);
nand U16563 (N_16563,N_15200,N_15401);
or U16564 (N_16564,N_15303,N_15890);
or U16565 (N_16565,N_15649,N_15797);
xor U16566 (N_16566,N_15423,N_15263);
and U16567 (N_16567,N_15900,N_15666);
and U16568 (N_16568,N_15567,N_15988);
or U16569 (N_16569,N_15892,N_15418);
or U16570 (N_16570,N_15368,N_15219);
and U16571 (N_16571,N_15875,N_15968);
and U16572 (N_16572,N_15368,N_15960);
nor U16573 (N_16573,N_15281,N_15618);
xor U16574 (N_16574,N_15628,N_15305);
or U16575 (N_16575,N_15729,N_15429);
and U16576 (N_16576,N_15554,N_15872);
xnor U16577 (N_16577,N_15614,N_15415);
and U16578 (N_16578,N_15216,N_15690);
or U16579 (N_16579,N_15274,N_15386);
or U16580 (N_16580,N_15969,N_15864);
nor U16581 (N_16581,N_15699,N_15672);
and U16582 (N_16582,N_15790,N_15301);
xor U16583 (N_16583,N_15975,N_15277);
nand U16584 (N_16584,N_15358,N_15343);
or U16585 (N_16585,N_15213,N_15261);
and U16586 (N_16586,N_15692,N_15613);
nor U16587 (N_16587,N_15830,N_15498);
xnor U16588 (N_16588,N_15379,N_15861);
nor U16589 (N_16589,N_15266,N_15793);
or U16590 (N_16590,N_15880,N_15229);
xnor U16591 (N_16591,N_15725,N_15327);
and U16592 (N_16592,N_15279,N_15761);
or U16593 (N_16593,N_15745,N_15523);
nor U16594 (N_16594,N_15454,N_15308);
and U16595 (N_16595,N_15550,N_15747);
xor U16596 (N_16596,N_15499,N_15510);
or U16597 (N_16597,N_15581,N_15446);
xnor U16598 (N_16598,N_15927,N_15813);
or U16599 (N_16599,N_15777,N_15559);
xnor U16600 (N_16600,N_15555,N_15714);
and U16601 (N_16601,N_15821,N_15255);
nand U16602 (N_16602,N_15878,N_15457);
nor U16603 (N_16603,N_15613,N_15870);
or U16604 (N_16604,N_15972,N_15858);
and U16605 (N_16605,N_15545,N_15307);
or U16606 (N_16606,N_15905,N_15419);
and U16607 (N_16607,N_15237,N_15554);
nand U16608 (N_16608,N_15740,N_15727);
and U16609 (N_16609,N_15422,N_15355);
or U16610 (N_16610,N_15898,N_15709);
and U16611 (N_16611,N_15307,N_15585);
or U16612 (N_16612,N_15393,N_15336);
nand U16613 (N_16613,N_15890,N_15248);
and U16614 (N_16614,N_15452,N_15216);
nand U16615 (N_16615,N_15590,N_15370);
nor U16616 (N_16616,N_15870,N_15441);
or U16617 (N_16617,N_15430,N_15717);
xor U16618 (N_16618,N_15599,N_15433);
xnor U16619 (N_16619,N_15364,N_15216);
nor U16620 (N_16620,N_15710,N_15920);
and U16621 (N_16621,N_15360,N_15724);
nor U16622 (N_16622,N_15296,N_15808);
nand U16623 (N_16623,N_15787,N_15391);
nand U16624 (N_16624,N_15605,N_15424);
and U16625 (N_16625,N_15383,N_15827);
and U16626 (N_16626,N_15205,N_15611);
nand U16627 (N_16627,N_15926,N_15706);
and U16628 (N_16628,N_15916,N_15547);
nor U16629 (N_16629,N_15440,N_15671);
nor U16630 (N_16630,N_15857,N_15262);
nand U16631 (N_16631,N_15940,N_15298);
xor U16632 (N_16632,N_15580,N_15461);
xnor U16633 (N_16633,N_15516,N_15304);
xnor U16634 (N_16634,N_15860,N_15811);
nor U16635 (N_16635,N_15674,N_15355);
and U16636 (N_16636,N_15255,N_15617);
nand U16637 (N_16637,N_15815,N_15440);
nor U16638 (N_16638,N_15944,N_15706);
or U16639 (N_16639,N_15444,N_15450);
nor U16640 (N_16640,N_15325,N_15556);
or U16641 (N_16641,N_15430,N_15307);
nor U16642 (N_16642,N_15844,N_15615);
xor U16643 (N_16643,N_15981,N_15351);
nor U16644 (N_16644,N_15516,N_15534);
and U16645 (N_16645,N_15257,N_15543);
or U16646 (N_16646,N_15654,N_15834);
xor U16647 (N_16647,N_15517,N_15648);
and U16648 (N_16648,N_15946,N_15952);
or U16649 (N_16649,N_15648,N_15568);
xor U16650 (N_16650,N_15391,N_15832);
and U16651 (N_16651,N_15349,N_15496);
or U16652 (N_16652,N_15853,N_15395);
or U16653 (N_16653,N_15286,N_15885);
and U16654 (N_16654,N_15576,N_15800);
nor U16655 (N_16655,N_15550,N_15824);
nor U16656 (N_16656,N_15871,N_15339);
and U16657 (N_16657,N_15892,N_15229);
xnor U16658 (N_16658,N_15201,N_15902);
and U16659 (N_16659,N_15456,N_15653);
and U16660 (N_16660,N_15934,N_15722);
or U16661 (N_16661,N_15818,N_15398);
xnor U16662 (N_16662,N_15423,N_15408);
and U16663 (N_16663,N_15608,N_15261);
nand U16664 (N_16664,N_15567,N_15440);
nor U16665 (N_16665,N_15580,N_15610);
and U16666 (N_16666,N_15729,N_15328);
nand U16667 (N_16667,N_15275,N_15328);
nor U16668 (N_16668,N_15849,N_15278);
nor U16669 (N_16669,N_15987,N_15899);
nor U16670 (N_16670,N_15675,N_15597);
xnor U16671 (N_16671,N_15678,N_15606);
and U16672 (N_16672,N_15890,N_15807);
xor U16673 (N_16673,N_15696,N_15352);
or U16674 (N_16674,N_15564,N_15740);
or U16675 (N_16675,N_15567,N_15950);
and U16676 (N_16676,N_15301,N_15738);
xnor U16677 (N_16677,N_15373,N_15247);
or U16678 (N_16678,N_15552,N_15756);
or U16679 (N_16679,N_15235,N_15800);
and U16680 (N_16680,N_15273,N_15915);
or U16681 (N_16681,N_15716,N_15533);
or U16682 (N_16682,N_15564,N_15961);
nand U16683 (N_16683,N_15887,N_15315);
nor U16684 (N_16684,N_15817,N_15864);
nand U16685 (N_16685,N_15201,N_15819);
nor U16686 (N_16686,N_15744,N_15862);
and U16687 (N_16687,N_15272,N_15451);
and U16688 (N_16688,N_15697,N_15761);
and U16689 (N_16689,N_15303,N_15630);
xnor U16690 (N_16690,N_15360,N_15855);
xnor U16691 (N_16691,N_15276,N_15320);
or U16692 (N_16692,N_15979,N_15783);
or U16693 (N_16693,N_15888,N_15959);
xnor U16694 (N_16694,N_15504,N_15303);
nor U16695 (N_16695,N_15949,N_15764);
nor U16696 (N_16696,N_15999,N_15250);
nor U16697 (N_16697,N_15429,N_15289);
or U16698 (N_16698,N_15670,N_15309);
and U16699 (N_16699,N_15379,N_15953);
or U16700 (N_16700,N_15845,N_15883);
or U16701 (N_16701,N_15924,N_15707);
nand U16702 (N_16702,N_15825,N_15974);
nand U16703 (N_16703,N_15275,N_15603);
xor U16704 (N_16704,N_15937,N_15895);
and U16705 (N_16705,N_15213,N_15842);
or U16706 (N_16706,N_15262,N_15764);
nand U16707 (N_16707,N_15446,N_15666);
and U16708 (N_16708,N_15916,N_15429);
xor U16709 (N_16709,N_15322,N_15450);
or U16710 (N_16710,N_15854,N_15972);
nor U16711 (N_16711,N_15253,N_15357);
and U16712 (N_16712,N_15542,N_15473);
or U16713 (N_16713,N_15484,N_15968);
nor U16714 (N_16714,N_15733,N_15984);
and U16715 (N_16715,N_15527,N_15231);
nand U16716 (N_16716,N_15237,N_15269);
xnor U16717 (N_16717,N_15567,N_15304);
nand U16718 (N_16718,N_15707,N_15899);
and U16719 (N_16719,N_15353,N_15457);
xor U16720 (N_16720,N_15622,N_15695);
xnor U16721 (N_16721,N_15295,N_15210);
and U16722 (N_16722,N_15463,N_15800);
or U16723 (N_16723,N_15659,N_15762);
xor U16724 (N_16724,N_15215,N_15957);
or U16725 (N_16725,N_15491,N_15831);
or U16726 (N_16726,N_15867,N_15507);
nor U16727 (N_16727,N_15647,N_15563);
xnor U16728 (N_16728,N_15281,N_15951);
or U16729 (N_16729,N_15461,N_15330);
nand U16730 (N_16730,N_15592,N_15976);
nor U16731 (N_16731,N_15361,N_15513);
and U16732 (N_16732,N_15772,N_15752);
and U16733 (N_16733,N_15600,N_15276);
xnor U16734 (N_16734,N_15974,N_15966);
nor U16735 (N_16735,N_15765,N_15857);
nand U16736 (N_16736,N_15255,N_15743);
xnor U16737 (N_16737,N_15534,N_15678);
xnor U16738 (N_16738,N_15576,N_15250);
nand U16739 (N_16739,N_15205,N_15258);
nor U16740 (N_16740,N_15245,N_15228);
nand U16741 (N_16741,N_15856,N_15331);
nand U16742 (N_16742,N_15675,N_15682);
and U16743 (N_16743,N_15854,N_15662);
or U16744 (N_16744,N_15253,N_15545);
nand U16745 (N_16745,N_15622,N_15540);
and U16746 (N_16746,N_15992,N_15868);
and U16747 (N_16747,N_15767,N_15320);
xnor U16748 (N_16748,N_15965,N_15746);
nand U16749 (N_16749,N_15599,N_15465);
nand U16750 (N_16750,N_15489,N_15444);
and U16751 (N_16751,N_15829,N_15604);
nand U16752 (N_16752,N_15210,N_15784);
xnor U16753 (N_16753,N_15728,N_15716);
or U16754 (N_16754,N_15290,N_15517);
and U16755 (N_16755,N_15488,N_15618);
xnor U16756 (N_16756,N_15500,N_15508);
nor U16757 (N_16757,N_15973,N_15218);
xnor U16758 (N_16758,N_15272,N_15359);
nor U16759 (N_16759,N_15589,N_15485);
nand U16760 (N_16760,N_15933,N_15793);
nand U16761 (N_16761,N_15538,N_15421);
and U16762 (N_16762,N_15320,N_15578);
nor U16763 (N_16763,N_15705,N_15652);
xnor U16764 (N_16764,N_15495,N_15657);
xor U16765 (N_16765,N_15952,N_15793);
nand U16766 (N_16766,N_15941,N_15419);
nand U16767 (N_16767,N_15519,N_15360);
or U16768 (N_16768,N_15265,N_15874);
and U16769 (N_16769,N_15217,N_15910);
or U16770 (N_16770,N_15774,N_15486);
xor U16771 (N_16771,N_15631,N_15757);
xor U16772 (N_16772,N_15683,N_15561);
or U16773 (N_16773,N_15639,N_15695);
nor U16774 (N_16774,N_15658,N_15609);
nor U16775 (N_16775,N_15998,N_15594);
xor U16776 (N_16776,N_15520,N_15995);
xnor U16777 (N_16777,N_15985,N_15653);
nor U16778 (N_16778,N_15895,N_15997);
nand U16779 (N_16779,N_15933,N_15240);
nor U16780 (N_16780,N_15626,N_15468);
and U16781 (N_16781,N_15361,N_15607);
nor U16782 (N_16782,N_15609,N_15282);
xor U16783 (N_16783,N_15519,N_15694);
or U16784 (N_16784,N_15273,N_15372);
xor U16785 (N_16785,N_15897,N_15863);
or U16786 (N_16786,N_15882,N_15246);
xor U16787 (N_16787,N_15466,N_15564);
and U16788 (N_16788,N_15790,N_15948);
nand U16789 (N_16789,N_15945,N_15563);
nor U16790 (N_16790,N_15654,N_15692);
or U16791 (N_16791,N_15610,N_15285);
xor U16792 (N_16792,N_15968,N_15291);
or U16793 (N_16793,N_15204,N_15580);
and U16794 (N_16794,N_15204,N_15806);
nor U16795 (N_16795,N_15801,N_15655);
and U16796 (N_16796,N_15936,N_15609);
and U16797 (N_16797,N_15496,N_15827);
xor U16798 (N_16798,N_15738,N_15218);
or U16799 (N_16799,N_15913,N_15998);
nor U16800 (N_16800,N_16298,N_16148);
nor U16801 (N_16801,N_16137,N_16061);
nand U16802 (N_16802,N_16026,N_16668);
or U16803 (N_16803,N_16636,N_16005);
nand U16804 (N_16804,N_16373,N_16192);
or U16805 (N_16805,N_16627,N_16696);
nand U16806 (N_16806,N_16799,N_16057);
xnor U16807 (N_16807,N_16366,N_16112);
nor U16808 (N_16808,N_16055,N_16170);
nor U16809 (N_16809,N_16455,N_16491);
or U16810 (N_16810,N_16609,N_16033);
and U16811 (N_16811,N_16637,N_16706);
nand U16812 (N_16812,N_16386,N_16722);
xnor U16813 (N_16813,N_16710,N_16405);
nor U16814 (N_16814,N_16506,N_16252);
and U16815 (N_16815,N_16716,N_16259);
xnor U16816 (N_16816,N_16437,N_16363);
xnor U16817 (N_16817,N_16034,N_16218);
nor U16818 (N_16818,N_16253,N_16368);
and U16819 (N_16819,N_16633,N_16798);
nand U16820 (N_16820,N_16233,N_16529);
nand U16821 (N_16821,N_16447,N_16182);
and U16822 (N_16822,N_16143,N_16275);
nor U16823 (N_16823,N_16757,N_16231);
nor U16824 (N_16824,N_16283,N_16793);
and U16825 (N_16825,N_16770,N_16240);
xor U16826 (N_16826,N_16665,N_16213);
nand U16827 (N_16827,N_16356,N_16600);
nor U16828 (N_16828,N_16224,N_16206);
or U16829 (N_16829,N_16084,N_16277);
or U16830 (N_16830,N_16530,N_16689);
or U16831 (N_16831,N_16395,N_16272);
or U16832 (N_16832,N_16513,N_16420);
or U16833 (N_16833,N_16255,N_16642);
nand U16834 (N_16834,N_16071,N_16569);
or U16835 (N_16835,N_16583,N_16700);
and U16836 (N_16836,N_16563,N_16495);
nor U16837 (N_16837,N_16508,N_16621);
nor U16838 (N_16838,N_16557,N_16021);
nor U16839 (N_16839,N_16701,N_16264);
and U16840 (N_16840,N_16527,N_16296);
nand U16841 (N_16841,N_16337,N_16760);
nand U16842 (N_16842,N_16573,N_16490);
nand U16843 (N_16843,N_16762,N_16379);
and U16844 (N_16844,N_16528,N_16538);
xnor U16845 (N_16845,N_16531,N_16287);
xnor U16846 (N_16846,N_16592,N_16352);
or U16847 (N_16847,N_16324,N_16375);
xnor U16848 (N_16848,N_16485,N_16736);
and U16849 (N_16849,N_16318,N_16691);
nor U16850 (N_16850,N_16299,N_16791);
or U16851 (N_16851,N_16499,N_16606);
xnor U16852 (N_16852,N_16131,N_16388);
nand U16853 (N_16853,N_16501,N_16780);
nor U16854 (N_16854,N_16079,N_16176);
or U16855 (N_16855,N_16778,N_16484);
nand U16856 (N_16856,N_16288,N_16759);
or U16857 (N_16857,N_16291,N_16751);
xor U16858 (N_16858,N_16140,N_16579);
nor U16859 (N_16859,N_16322,N_16436);
nand U16860 (N_16860,N_16685,N_16384);
and U16861 (N_16861,N_16221,N_16747);
nor U16862 (N_16862,N_16173,N_16243);
nor U16863 (N_16863,N_16695,N_16043);
xor U16864 (N_16864,N_16456,N_16237);
xnor U16865 (N_16865,N_16086,N_16385);
xnor U16866 (N_16866,N_16185,N_16096);
nor U16867 (N_16867,N_16149,N_16461);
xnor U16868 (N_16868,N_16274,N_16300);
nor U16869 (N_16869,N_16425,N_16784);
and U16870 (N_16870,N_16415,N_16066);
nor U16871 (N_16871,N_16153,N_16678);
or U16872 (N_16872,N_16400,N_16768);
and U16873 (N_16873,N_16587,N_16301);
or U16874 (N_16874,N_16248,N_16167);
nor U16875 (N_16875,N_16432,N_16006);
or U16876 (N_16876,N_16207,N_16397);
and U16877 (N_16877,N_16596,N_16630);
and U16878 (N_16878,N_16074,N_16645);
or U16879 (N_16879,N_16104,N_16335);
nor U16880 (N_16880,N_16660,N_16315);
nand U16881 (N_16881,N_16601,N_16174);
or U16882 (N_16882,N_16681,N_16486);
or U16883 (N_16883,N_16551,N_16466);
nor U16884 (N_16884,N_16163,N_16354);
nor U16885 (N_16885,N_16577,N_16441);
nand U16886 (N_16886,N_16469,N_16521);
nor U16887 (N_16887,N_16687,N_16216);
nand U16888 (N_16888,N_16171,N_16746);
nor U16889 (N_16889,N_16719,N_16686);
or U16890 (N_16890,N_16404,N_16795);
or U16891 (N_16891,N_16351,N_16323);
xnor U16892 (N_16892,N_16305,N_16520);
nor U16893 (N_16893,N_16113,N_16347);
or U16894 (N_16894,N_16052,N_16554);
xor U16895 (N_16895,N_16050,N_16503);
nand U16896 (N_16896,N_16348,N_16027);
and U16897 (N_16897,N_16230,N_16572);
nand U16898 (N_16898,N_16403,N_16412);
or U16899 (N_16899,N_16064,N_16378);
or U16900 (N_16900,N_16256,N_16444);
nor U16901 (N_16901,N_16029,N_16732);
nor U16902 (N_16902,N_16735,N_16342);
or U16903 (N_16903,N_16109,N_16576);
nand U16904 (N_16904,N_16279,N_16377);
nor U16905 (N_16905,N_16196,N_16344);
nor U16906 (N_16906,N_16445,N_16118);
nand U16907 (N_16907,N_16741,N_16376);
or U16908 (N_16908,N_16451,N_16470);
or U16909 (N_16909,N_16629,N_16419);
nand U16910 (N_16910,N_16399,N_16136);
nor U16911 (N_16911,N_16797,N_16225);
nor U16912 (N_16912,N_16281,N_16201);
nor U16913 (N_16913,N_16615,N_16350);
xnor U16914 (N_16914,N_16028,N_16565);
and U16915 (N_16915,N_16115,N_16449);
or U16916 (N_16916,N_16493,N_16679);
nand U16917 (N_16917,N_16250,N_16160);
nand U16918 (N_16918,N_16263,N_16193);
and U16919 (N_16919,N_16720,N_16197);
and U16920 (N_16920,N_16144,N_16316);
and U16921 (N_16921,N_16122,N_16478);
nand U16922 (N_16922,N_16737,N_16650);
xor U16923 (N_16923,N_16589,N_16699);
xnor U16924 (N_16924,N_16777,N_16523);
or U16925 (N_16925,N_16640,N_16708);
nand U16926 (N_16926,N_16638,N_16219);
nor U16927 (N_16927,N_16093,N_16675);
xor U16928 (N_16928,N_16236,N_16653);
or U16929 (N_16929,N_16763,N_16001);
and U16930 (N_16930,N_16724,N_16663);
nand U16931 (N_16931,N_16391,N_16526);
xor U16932 (N_16932,N_16308,N_16254);
and U16933 (N_16933,N_16138,N_16035);
and U16934 (N_16934,N_16556,N_16726);
or U16935 (N_16935,N_16246,N_16048);
and U16936 (N_16936,N_16059,N_16776);
or U16937 (N_16937,N_16519,N_16326);
xnor U16938 (N_16938,N_16032,N_16658);
or U16939 (N_16939,N_16178,N_16772);
nor U16940 (N_16940,N_16383,N_16133);
and U16941 (N_16941,N_16030,N_16620);
xor U16942 (N_16942,N_16234,N_16533);
or U16943 (N_16943,N_16209,N_16756);
and U16944 (N_16944,N_16690,N_16704);
and U16945 (N_16945,N_16771,N_16319);
xor U16946 (N_16946,N_16677,N_16282);
nor U16947 (N_16947,N_16090,N_16217);
nand U16948 (N_16948,N_16588,N_16498);
or U16949 (N_16949,N_16198,N_16458);
nor U16950 (N_16950,N_16428,N_16155);
nor U16951 (N_16951,N_16078,N_16649);
xor U16952 (N_16952,N_16743,N_16166);
or U16953 (N_16953,N_16085,N_16302);
nand U16954 (N_16954,N_16159,N_16013);
nor U16955 (N_16955,N_16179,N_16730);
and U16956 (N_16956,N_16471,N_16421);
nand U16957 (N_16957,N_16157,N_16709);
xnor U16958 (N_16958,N_16295,N_16715);
xor U16959 (N_16959,N_16742,N_16416);
nor U16960 (N_16960,N_16422,N_16102);
or U16961 (N_16961,N_16036,N_16473);
and U16962 (N_16962,N_16651,N_16580);
or U16963 (N_16963,N_16489,N_16492);
and U16964 (N_16964,N_16602,N_16229);
nor U16965 (N_16965,N_16518,N_16380);
or U16966 (N_16966,N_16512,N_16619);
nand U16967 (N_16967,N_16270,N_16666);
xnor U16968 (N_16968,N_16475,N_16189);
nor U16969 (N_16969,N_16524,N_16023);
or U16970 (N_16970,N_16744,N_16188);
nand U16971 (N_16971,N_16442,N_16543);
or U16972 (N_16972,N_16306,N_16164);
nand U16973 (N_16973,N_16063,N_16483);
nand U16974 (N_16974,N_16123,N_16697);
nand U16975 (N_16975,N_16494,N_16725);
xnor U16976 (N_16976,N_16703,N_16345);
nand U16977 (N_16977,N_16408,N_16394);
or U16978 (N_16978,N_16424,N_16152);
and U16979 (N_16979,N_16532,N_16657);
nand U16980 (N_16980,N_16738,N_16003);
nor U16981 (N_16981,N_16245,N_16370);
xnor U16982 (N_16982,N_16010,N_16570);
nor U16983 (N_16983,N_16783,N_16477);
xor U16984 (N_16984,N_16076,N_16124);
nand U16985 (N_16985,N_16616,N_16022);
nand U16986 (N_16986,N_16232,N_16622);
and U16987 (N_16987,N_16500,N_16154);
nor U16988 (N_16988,N_16625,N_16349);
xor U16989 (N_16989,N_16567,N_16177);
and U16990 (N_16990,N_16460,N_16313);
or U16991 (N_16991,N_16586,N_16119);
xor U16992 (N_16992,N_16247,N_16314);
and U16993 (N_16993,N_16514,N_16381);
or U16994 (N_16994,N_16094,N_16355);
nor U16995 (N_16995,N_16748,N_16121);
or U16996 (N_16996,N_16558,N_16099);
nor U16997 (N_16997,N_16562,N_16434);
xor U16998 (N_16998,N_16517,N_16639);
nand U16999 (N_16999,N_16509,N_16410);
nor U17000 (N_17000,N_16362,N_16135);
nor U17001 (N_17001,N_16750,N_16430);
xor U17002 (N_17002,N_16360,N_16566);
xor U17003 (N_17003,N_16037,N_16018);
or U17004 (N_17004,N_16480,N_16393);
xnor U17005 (N_17005,N_16550,N_16194);
nand U17006 (N_17006,N_16238,N_16794);
and U17007 (N_17007,N_16260,N_16559);
and U17008 (N_17008,N_16753,N_16025);
and U17009 (N_17009,N_16435,N_16235);
nor U17010 (N_17010,N_16398,N_16593);
or U17011 (N_17011,N_16151,N_16479);
and U17012 (N_17012,N_16082,N_16116);
or U17013 (N_17013,N_16648,N_16613);
nand U17014 (N_17014,N_16330,N_16773);
and U17015 (N_17015,N_16017,N_16634);
nor U17016 (N_17016,N_16534,N_16605);
xor U17017 (N_17017,N_16284,N_16000);
xnor U17018 (N_17018,N_16100,N_16474);
or U17019 (N_17019,N_16598,N_16031);
nand U17020 (N_17020,N_16340,N_16423);
xor U17021 (N_17021,N_16597,N_16611);
or U17022 (N_17022,N_16047,N_16754);
nor U17023 (N_17023,N_16227,N_16226);
xor U17024 (N_17024,N_16038,N_16712);
nand U17025 (N_17025,N_16016,N_16214);
or U17026 (N_17026,N_16454,N_16095);
xor U17027 (N_17027,N_16183,N_16108);
or U17028 (N_17028,N_16367,N_16088);
or U17029 (N_17029,N_16548,N_16204);
nand U17030 (N_17030,N_16536,N_16591);
xor U17031 (N_17031,N_16464,N_16012);
and U17032 (N_17032,N_16443,N_16303);
or U17033 (N_17033,N_16585,N_16786);
xor U17034 (N_17034,N_16147,N_16073);
or U17035 (N_17035,N_16267,N_16120);
nand U17036 (N_17036,N_16242,N_16212);
nand U17037 (N_17037,N_16325,N_16705);
xnor U17038 (N_17038,N_16535,N_16610);
or U17039 (N_17039,N_16150,N_16262);
xnor U17040 (N_17040,N_16504,N_16056);
xnor U17041 (N_17041,N_16614,N_16781);
nand U17042 (N_17042,N_16788,N_16215);
or U17043 (N_17043,N_16683,N_16041);
xor U17044 (N_17044,N_16406,N_16244);
xor U17045 (N_17045,N_16292,N_16560);
or U17046 (N_17046,N_16612,N_16594);
nand U17047 (N_17047,N_16792,N_16643);
xor U17048 (N_17048,N_16293,N_16522);
or U17049 (N_17049,N_16785,N_16603);
nor U17050 (N_17050,N_16007,N_16662);
and U17051 (N_17051,N_16427,N_16769);
and U17052 (N_17052,N_16286,N_16546);
nand U17053 (N_17053,N_16008,N_16542);
and U17054 (N_17054,N_16659,N_16733);
and U17055 (N_17055,N_16269,N_16114);
xor U17056 (N_17056,N_16317,N_16265);
nor U17057 (N_17057,N_16667,N_16321);
or U17058 (N_17058,N_16544,N_16654);
or U17059 (N_17059,N_16239,N_16482);
or U17060 (N_17060,N_16172,N_16635);
and U17061 (N_17061,N_16652,N_16463);
xor U17062 (N_17062,N_16223,N_16693);
or U17063 (N_17063,N_16014,N_16186);
nor U17064 (N_17064,N_16540,N_16617);
nor U17065 (N_17065,N_16202,N_16343);
xnor U17066 (N_17066,N_16555,N_16672);
nand U17067 (N_17067,N_16561,N_16191);
and U17068 (N_17068,N_16407,N_16258);
or U17069 (N_17069,N_16053,N_16448);
xor U17070 (N_17070,N_16162,N_16049);
or U17071 (N_17071,N_16068,N_16009);
and U17072 (N_17072,N_16790,N_16595);
nor U17073 (N_17073,N_16765,N_16714);
and U17074 (N_17074,N_16329,N_16488);
nand U17075 (N_17075,N_16257,N_16702);
or U17076 (N_17076,N_16020,N_16101);
and U17077 (N_17077,N_16389,N_16045);
and U17078 (N_17078,N_16042,N_16199);
nor U17079 (N_17079,N_16452,N_16180);
and U17080 (N_17080,N_16761,N_16111);
and U17081 (N_17081,N_16766,N_16467);
or U17082 (N_17082,N_16307,N_16070);
and U17083 (N_17083,N_16626,N_16132);
and U17084 (N_17084,N_16142,N_16497);
nor U17085 (N_17085,N_16103,N_16165);
nand U17086 (N_17086,N_16549,N_16433);
xor U17087 (N_17087,N_16062,N_16450);
nor U17088 (N_17088,N_16208,N_16628);
and U17089 (N_17089,N_16106,N_16752);
nor U17090 (N_17090,N_16789,N_16655);
or U17091 (N_17091,N_16039,N_16599);
and U17092 (N_17092,N_16401,N_16320);
nor U17093 (N_17093,N_16065,N_16117);
and U17094 (N_17094,N_16713,N_16089);
nand U17095 (N_17095,N_16740,N_16080);
nand U17096 (N_17096,N_16688,N_16525);
and U17097 (N_17097,N_16092,N_16333);
or U17098 (N_17098,N_16755,N_16767);
nor U17099 (N_17099,N_16656,N_16134);
and U17100 (N_17100,N_16098,N_16564);
xor U17101 (N_17101,N_16220,N_16072);
nor U17102 (N_17102,N_16129,N_16146);
and U17103 (N_17103,N_16728,N_16141);
xnor U17104 (N_17104,N_16075,N_16673);
nand U17105 (N_17105,N_16083,N_16717);
nor U17106 (N_17106,N_16453,N_16414);
and U17107 (N_17107,N_16545,N_16390);
nand U17108 (N_17108,N_16511,N_16758);
and U17109 (N_17109,N_16462,N_16327);
and U17110 (N_17110,N_16409,N_16357);
and U17111 (N_17111,N_16251,N_16341);
and U17112 (N_17112,N_16294,N_16507);
xnor U17113 (N_17113,N_16331,N_16004);
nor U17114 (N_17114,N_16446,N_16418);
nor U17115 (N_17115,N_16684,N_16727);
nor U17116 (N_17116,N_16261,N_16547);
xor U17117 (N_17117,N_16002,N_16130);
nand U17118 (N_17118,N_16110,N_16280);
or U17119 (N_17119,N_16145,N_16734);
nand U17120 (N_17120,N_16336,N_16431);
xor U17121 (N_17121,N_16019,N_16775);
xor U17122 (N_17122,N_16024,N_16161);
or U17123 (N_17123,N_16632,N_16782);
xnor U17124 (N_17124,N_16505,N_16011);
nand U17125 (N_17125,N_16387,N_16481);
xor U17126 (N_17126,N_16175,N_16077);
nor U17127 (N_17127,N_16676,N_16015);
nor U17128 (N_17128,N_16158,N_16210);
nor U17129 (N_17129,N_16359,N_16107);
xor U17130 (N_17130,N_16718,N_16631);
xnor U17131 (N_17131,N_16510,N_16181);
xnor U17132 (N_17132,N_16670,N_16439);
or U17133 (N_17133,N_16374,N_16440);
nand U17134 (N_17134,N_16698,N_16273);
nand U17135 (N_17135,N_16516,N_16312);
nor U17136 (N_17136,N_16334,N_16457);
and U17137 (N_17137,N_16607,N_16353);
xnor U17138 (N_17138,N_16338,N_16097);
or U17139 (N_17139,N_16618,N_16044);
xnor U17140 (N_17140,N_16241,N_16417);
and U17141 (N_17141,N_16156,N_16332);
xor U17142 (N_17142,N_16276,N_16623);
nand U17143 (N_17143,N_16578,N_16304);
xor U17144 (N_17144,N_16680,N_16311);
nand U17145 (N_17145,N_16465,N_16552);
nor U17146 (N_17146,N_16515,N_16184);
and U17147 (N_17147,N_16694,N_16139);
xor U17148 (N_17148,N_16127,N_16669);
xnor U17149 (N_17149,N_16711,N_16268);
nor U17150 (N_17150,N_16200,N_16372);
xor U17151 (N_17151,N_16721,N_16060);
nand U17152 (N_17152,N_16476,N_16438);
xnor U17153 (N_17153,N_16249,N_16346);
nor U17154 (N_17154,N_16553,N_16087);
xnor U17155 (N_17155,N_16169,N_16644);
and U17156 (N_17156,N_16289,N_16537);
and U17157 (N_17157,N_16723,N_16222);
or U17158 (N_17158,N_16392,N_16128);
nand U17159 (N_17159,N_16040,N_16682);
nand U17160 (N_17160,N_16496,N_16468);
xor U17161 (N_17161,N_16067,N_16729);
or U17162 (N_17162,N_16647,N_16285);
or U17163 (N_17163,N_16787,N_16774);
and U17164 (N_17164,N_16369,N_16069);
and U17165 (N_17165,N_16168,N_16271);
nand U17166 (N_17166,N_16571,N_16297);
and U17167 (N_17167,N_16081,N_16541);
xor U17168 (N_17168,N_16402,N_16364);
nand U17169 (N_17169,N_16054,N_16487);
and U17170 (N_17170,N_16779,N_16105);
or U17171 (N_17171,N_16584,N_16371);
nor U17172 (N_17172,N_16358,N_16731);
nand U17173 (N_17173,N_16661,N_16575);
or U17174 (N_17174,N_16574,N_16365);
xnor U17175 (N_17175,N_16581,N_16707);
or U17176 (N_17176,N_16382,N_16502);
nand U17177 (N_17177,N_16459,N_16278);
and U17178 (N_17178,N_16211,N_16413);
or U17179 (N_17179,N_16472,N_16604);
xnor U17180 (N_17180,N_16739,N_16091);
and U17181 (N_17181,N_16539,N_16187);
nor U17182 (N_17182,N_16582,N_16749);
nand U17183 (N_17183,N_16692,N_16396);
and U17184 (N_17184,N_16745,N_16126);
nand U17185 (N_17185,N_16568,N_16058);
or U17186 (N_17186,N_16125,N_16328);
xnor U17187 (N_17187,N_16361,N_16590);
or U17188 (N_17188,N_16671,N_16796);
nor U17189 (N_17189,N_16309,N_16429);
xor U17190 (N_17190,N_16046,N_16339);
xor U17191 (N_17191,N_16051,N_16426);
nor U17192 (N_17192,N_16641,N_16624);
nor U17193 (N_17193,N_16203,N_16608);
xor U17194 (N_17194,N_16195,N_16190);
nor U17195 (N_17195,N_16228,N_16290);
nand U17196 (N_17196,N_16646,N_16266);
nand U17197 (N_17197,N_16205,N_16664);
and U17198 (N_17198,N_16674,N_16310);
nor U17199 (N_17199,N_16764,N_16411);
nor U17200 (N_17200,N_16760,N_16714);
nor U17201 (N_17201,N_16747,N_16186);
nand U17202 (N_17202,N_16682,N_16621);
nand U17203 (N_17203,N_16104,N_16782);
and U17204 (N_17204,N_16419,N_16627);
and U17205 (N_17205,N_16362,N_16723);
and U17206 (N_17206,N_16668,N_16408);
nand U17207 (N_17207,N_16328,N_16681);
or U17208 (N_17208,N_16794,N_16518);
xor U17209 (N_17209,N_16386,N_16363);
or U17210 (N_17210,N_16613,N_16783);
nand U17211 (N_17211,N_16025,N_16784);
or U17212 (N_17212,N_16660,N_16691);
and U17213 (N_17213,N_16139,N_16536);
or U17214 (N_17214,N_16460,N_16287);
nor U17215 (N_17215,N_16560,N_16622);
xor U17216 (N_17216,N_16757,N_16210);
or U17217 (N_17217,N_16270,N_16585);
nor U17218 (N_17218,N_16251,N_16105);
nor U17219 (N_17219,N_16013,N_16745);
nand U17220 (N_17220,N_16407,N_16693);
xor U17221 (N_17221,N_16028,N_16393);
nor U17222 (N_17222,N_16211,N_16459);
xor U17223 (N_17223,N_16769,N_16771);
and U17224 (N_17224,N_16158,N_16332);
or U17225 (N_17225,N_16515,N_16297);
nor U17226 (N_17226,N_16264,N_16545);
nor U17227 (N_17227,N_16415,N_16020);
nor U17228 (N_17228,N_16421,N_16146);
nand U17229 (N_17229,N_16261,N_16623);
or U17230 (N_17230,N_16495,N_16549);
nor U17231 (N_17231,N_16576,N_16168);
nand U17232 (N_17232,N_16286,N_16110);
nand U17233 (N_17233,N_16495,N_16698);
or U17234 (N_17234,N_16514,N_16246);
nor U17235 (N_17235,N_16461,N_16752);
and U17236 (N_17236,N_16768,N_16231);
or U17237 (N_17237,N_16684,N_16649);
or U17238 (N_17238,N_16388,N_16776);
and U17239 (N_17239,N_16694,N_16123);
xnor U17240 (N_17240,N_16365,N_16315);
xnor U17241 (N_17241,N_16493,N_16688);
xor U17242 (N_17242,N_16263,N_16359);
nand U17243 (N_17243,N_16562,N_16334);
or U17244 (N_17244,N_16593,N_16131);
xnor U17245 (N_17245,N_16315,N_16482);
or U17246 (N_17246,N_16076,N_16577);
nand U17247 (N_17247,N_16195,N_16662);
nor U17248 (N_17248,N_16046,N_16607);
nand U17249 (N_17249,N_16490,N_16375);
nand U17250 (N_17250,N_16282,N_16469);
nand U17251 (N_17251,N_16696,N_16384);
nor U17252 (N_17252,N_16738,N_16531);
nor U17253 (N_17253,N_16497,N_16593);
or U17254 (N_17254,N_16771,N_16784);
and U17255 (N_17255,N_16431,N_16335);
nand U17256 (N_17256,N_16352,N_16575);
or U17257 (N_17257,N_16217,N_16422);
xor U17258 (N_17258,N_16247,N_16395);
nor U17259 (N_17259,N_16620,N_16745);
or U17260 (N_17260,N_16578,N_16711);
or U17261 (N_17261,N_16722,N_16010);
and U17262 (N_17262,N_16646,N_16230);
xnor U17263 (N_17263,N_16150,N_16319);
nor U17264 (N_17264,N_16044,N_16732);
nor U17265 (N_17265,N_16246,N_16631);
or U17266 (N_17266,N_16268,N_16052);
nand U17267 (N_17267,N_16369,N_16009);
nor U17268 (N_17268,N_16476,N_16647);
nand U17269 (N_17269,N_16281,N_16023);
xnor U17270 (N_17270,N_16621,N_16714);
nand U17271 (N_17271,N_16584,N_16471);
nor U17272 (N_17272,N_16241,N_16531);
and U17273 (N_17273,N_16783,N_16286);
and U17274 (N_17274,N_16041,N_16063);
xnor U17275 (N_17275,N_16214,N_16186);
nor U17276 (N_17276,N_16119,N_16471);
or U17277 (N_17277,N_16180,N_16339);
nor U17278 (N_17278,N_16020,N_16644);
nor U17279 (N_17279,N_16013,N_16702);
or U17280 (N_17280,N_16062,N_16379);
nand U17281 (N_17281,N_16218,N_16385);
xor U17282 (N_17282,N_16499,N_16089);
or U17283 (N_17283,N_16749,N_16474);
or U17284 (N_17284,N_16676,N_16561);
and U17285 (N_17285,N_16520,N_16644);
nor U17286 (N_17286,N_16477,N_16218);
nor U17287 (N_17287,N_16780,N_16272);
or U17288 (N_17288,N_16743,N_16732);
xnor U17289 (N_17289,N_16332,N_16221);
nand U17290 (N_17290,N_16470,N_16123);
and U17291 (N_17291,N_16123,N_16640);
nand U17292 (N_17292,N_16781,N_16578);
or U17293 (N_17293,N_16372,N_16554);
nand U17294 (N_17294,N_16482,N_16419);
xnor U17295 (N_17295,N_16207,N_16707);
or U17296 (N_17296,N_16435,N_16795);
or U17297 (N_17297,N_16613,N_16484);
nor U17298 (N_17298,N_16749,N_16432);
xnor U17299 (N_17299,N_16247,N_16079);
xnor U17300 (N_17300,N_16536,N_16289);
xor U17301 (N_17301,N_16768,N_16323);
and U17302 (N_17302,N_16675,N_16581);
xor U17303 (N_17303,N_16680,N_16078);
nand U17304 (N_17304,N_16534,N_16514);
or U17305 (N_17305,N_16170,N_16740);
nand U17306 (N_17306,N_16164,N_16249);
xnor U17307 (N_17307,N_16063,N_16261);
and U17308 (N_17308,N_16683,N_16136);
and U17309 (N_17309,N_16017,N_16651);
nand U17310 (N_17310,N_16251,N_16092);
and U17311 (N_17311,N_16115,N_16366);
and U17312 (N_17312,N_16279,N_16729);
nor U17313 (N_17313,N_16609,N_16255);
nor U17314 (N_17314,N_16505,N_16347);
nor U17315 (N_17315,N_16692,N_16476);
and U17316 (N_17316,N_16370,N_16176);
xnor U17317 (N_17317,N_16626,N_16248);
nand U17318 (N_17318,N_16406,N_16676);
nand U17319 (N_17319,N_16589,N_16530);
and U17320 (N_17320,N_16585,N_16232);
nor U17321 (N_17321,N_16205,N_16175);
xnor U17322 (N_17322,N_16194,N_16710);
or U17323 (N_17323,N_16000,N_16294);
and U17324 (N_17324,N_16342,N_16629);
xor U17325 (N_17325,N_16058,N_16792);
and U17326 (N_17326,N_16445,N_16090);
or U17327 (N_17327,N_16112,N_16223);
nand U17328 (N_17328,N_16184,N_16239);
xor U17329 (N_17329,N_16598,N_16770);
xnor U17330 (N_17330,N_16459,N_16677);
xnor U17331 (N_17331,N_16783,N_16636);
xnor U17332 (N_17332,N_16631,N_16103);
and U17333 (N_17333,N_16447,N_16573);
nand U17334 (N_17334,N_16457,N_16185);
nand U17335 (N_17335,N_16787,N_16546);
nor U17336 (N_17336,N_16306,N_16034);
and U17337 (N_17337,N_16031,N_16245);
nand U17338 (N_17338,N_16498,N_16510);
nor U17339 (N_17339,N_16170,N_16748);
xor U17340 (N_17340,N_16441,N_16727);
nand U17341 (N_17341,N_16666,N_16041);
xor U17342 (N_17342,N_16631,N_16081);
and U17343 (N_17343,N_16466,N_16450);
nand U17344 (N_17344,N_16456,N_16025);
or U17345 (N_17345,N_16390,N_16167);
nor U17346 (N_17346,N_16041,N_16307);
or U17347 (N_17347,N_16217,N_16124);
or U17348 (N_17348,N_16454,N_16012);
xor U17349 (N_17349,N_16660,N_16740);
and U17350 (N_17350,N_16153,N_16383);
xnor U17351 (N_17351,N_16764,N_16280);
nand U17352 (N_17352,N_16302,N_16687);
or U17353 (N_17353,N_16112,N_16768);
nand U17354 (N_17354,N_16231,N_16026);
nand U17355 (N_17355,N_16269,N_16177);
nor U17356 (N_17356,N_16456,N_16131);
nand U17357 (N_17357,N_16000,N_16245);
xnor U17358 (N_17358,N_16286,N_16171);
and U17359 (N_17359,N_16596,N_16511);
and U17360 (N_17360,N_16303,N_16319);
and U17361 (N_17361,N_16336,N_16471);
nor U17362 (N_17362,N_16402,N_16425);
or U17363 (N_17363,N_16145,N_16700);
or U17364 (N_17364,N_16154,N_16687);
and U17365 (N_17365,N_16575,N_16401);
or U17366 (N_17366,N_16338,N_16008);
xnor U17367 (N_17367,N_16492,N_16000);
nand U17368 (N_17368,N_16640,N_16772);
xor U17369 (N_17369,N_16629,N_16728);
xor U17370 (N_17370,N_16040,N_16007);
nand U17371 (N_17371,N_16440,N_16760);
nor U17372 (N_17372,N_16505,N_16707);
nand U17373 (N_17373,N_16576,N_16251);
nor U17374 (N_17374,N_16726,N_16689);
or U17375 (N_17375,N_16083,N_16473);
or U17376 (N_17376,N_16680,N_16007);
nand U17377 (N_17377,N_16687,N_16399);
or U17378 (N_17378,N_16413,N_16439);
nor U17379 (N_17379,N_16161,N_16093);
nor U17380 (N_17380,N_16002,N_16498);
xor U17381 (N_17381,N_16109,N_16537);
and U17382 (N_17382,N_16119,N_16016);
and U17383 (N_17383,N_16049,N_16034);
and U17384 (N_17384,N_16497,N_16337);
and U17385 (N_17385,N_16360,N_16510);
or U17386 (N_17386,N_16179,N_16079);
or U17387 (N_17387,N_16417,N_16688);
nand U17388 (N_17388,N_16673,N_16385);
nand U17389 (N_17389,N_16152,N_16263);
xor U17390 (N_17390,N_16246,N_16499);
nand U17391 (N_17391,N_16643,N_16472);
xor U17392 (N_17392,N_16592,N_16057);
xnor U17393 (N_17393,N_16284,N_16057);
nor U17394 (N_17394,N_16005,N_16482);
and U17395 (N_17395,N_16474,N_16061);
nand U17396 (N_17396,N_16557,N_16631);
or U17397 (N_17397,N_16237,N_16398);
or U17398 (N_17398,N_16044,N_16439);
nand U17399 (N_17399,N_16186,N_16343);
nand U17400 (N_17400,N_16774,N_16022);
and U17401 (N_17401,N_16144,N_16574);
and U17402 (N_17402,N_16077,N_16176);
nand U17403 (N_17403,N_16542,N_16035);
and U17404 (N_17404,N_16414,N_16202);
xor U17405 (N_17405,N_16599,N_16336);
and U17406 (N_17406,N_16279,N_16181);
or U17407 (N_17407,N_16768,N_16227);
nor U17408 (N_17408,N_16137,N_16019);
nand U17409 (N_17409,N_16030,N_16581);
nand U17410 (N_17410,N_16369,N_16227);
xnor U17411 (N_17411,N_16313,N_16238);
and U17412 (N_17412,N_16723,N_16308);
nor U17413 (N_17413,N_16708,N_16587);
or U17414 (N_17414,N_16182,N_16730);
and U17415 (N_17415,N_16796,N_16133);
or U17416 (N_17416,N_16631,N_16179);
nor U17417 (N_17417,N_16450,N_16089);
nand U17418 (N_17418,N_16699,N_16663);
nor U17419 (N_17419,N_16267,N_16573);
xor U17420 (N_17420,N_16350,N_16492);
or U17421 (N_17421,N_16418,N_16559);
nand U17422 (N_17422,N_16742,N_16492);
and U17423 (N_17423,N_16190,N_16581);
xnor U17424 (N_17424,N_16570,N_16549);
and U17425 (N_17425,N_16193,N_16536);
nand U17426 (N_17426,N_16184,N_16379);
nand U17427 (N_17427,N_16726,N_16491);
xnor U17428 (N_17428,N_16259,N_16762);
and U17429 (N_17429,N_16011,N_16065);
xnor U17430 (N_17430,N_16180,N_16230);
nor U17431 (N_17431,N_16344,N_16696);
nor U17432 (N_17432,N_16038,N_16048);
xnor U17433 (N_17433,N_16632,N_16585);
and U17434 (N_17434,N_16696,N_16658);
and U17435 (N_17435,N_16711,N_16568);
nor U17436 (N_17436,N_16632,N_16144);
nor U17437 (N_17437,N_16738,N_16119);
and U17438 (N_17438,N_16287,N_16789);
and U17439 (N_17439,N_16058,N_16355);
or U17440 (N_17440,N_16730,N_16311);
xor U17441 (N_17441,N_16109,N_16056);
nand U17442 (N_17442,N_16679,N_16759);
and U17443 (N_17443,N_16618,N_16524);
nor U17444 (N_17444,N_16246,N_16037);
nand U17445 (N_17445,N_16698,N_16358);
and U17446 (N_17446,N_16049,N_16437);
nor U17447 (N_17447,N_16490,N_16799);
nand U17448 (N_17448,N_16649,N_16199);
and U17449 (N_17449,N_16346,N_16262);
or U17450 (N_17450,N_16047,N_16638);
and U17451 (N_17451,N_16046,N_16458);
nor U17452 (N_17452,N_16488,N_16674);
nand U17453 (N_17453,N_16265,N_16756);
or U17454 (N_17454,N_16111,N_16230);
or U17455 (N_17455,N_16520,N_16238);
nand U17456 (N_17456,N_16725,N_16574);
nor U17457 (N_17457,N_16369,N_16020);
nand U17458 (N_17458,N_16250,N_16549);
xor U17459 (N_17459,N_16194,N_16481);
nand U17460 (N_17460,N_16342,N_16276);
and U17461 (N_17461,N_16338,N_16437);
nor U17462 (N_17462,N_16402,N_16270);
nor U17463 (N_17463,N_16287,N_16219);
and U17464 (N_17464,N_16067,N_16768);
nor U17465 (N_17465,N_16515,N_16542);
nand U17466 (N_17466,N_16106,N_16107);
nor U17467 (N_17467,N_16575,N_16471);
nand U17468 (N_17468,N_16156,N_16183);
nor U17469 (N_17469,N_16496,N_16642);
nor U17470 (N_17470,N_16353,N_16715);
xnor U17471 (N_17471,N_16729,N_16769);
and U17472 (N_17472,N_16369,N_16716);
or U17473 (N_17473,N_16591,N_16325);
nand U17474 (N_17474,N_16474,N_16773);
nand U17475 (N_17475,N_16082,N_16721);
xor U17476 (N_17476,N_16449,N_16732);
xnor U17477 (N_17477,N_16197,N_16774);
or U17478 (N_17478,N_16126,N_16076);
nand U17479 (N_17479,N_16631,N_16578);
xnor U17480 (N_17480,N_16440,N_16204);
nor U17481 (N_17481,N_16552,N_16775);
nand U17482 (N_17482,N_16603,N_16197);
or U17483 (N_17483,N_16518,N_16467);
or U17484 (N_17484,N_16579,N_16674);
nand U17485 (N_17485,N_16109,N_16336);
and U17486 (N_17486,N_16071,N_16337);
xor U17487 (N_17487,N_16353,N_16199);
or U17488 (N_17488,N_16785,N_16046);
and U17489 (N_17489,N_16208,N_16301);
nor U17490 (N_17490,N_16423,N_16428);
xor U17491 (N_17491,N_16723,N_16304);
and U17492 (N_17492,N_16792,N_16149);
and U17493 (N_17493,N_16007,N_16643);
nor U17494 (N_17494,N_16404,N_16414);
or U17495 (N_17495,N_16409,N_16070);
and U17496 (N_17496,N_16624,N_16002);
xor U17497 (N_17497,N_16131,N_16635);
xor U17498 (N_17498,N_16208,N_16372);
or U17499 (N_17499,N_16380,N_16342);
and U17500 (N_17500,N_16269,N_16553);
xnor U17501 (N_17501,N_16184,N_16712);
and U17502 (N_17502,N_16623,N_16123);
and U17503 (N_17503,N_16246,N_16400);
or U17504 (N_17504,N_16571,N_16057);
nor U17505 (N_17505,N_16588,N_16149);
nand U17506 (N_17506,N_16490,N_16014);
xnor U17507 (N_17507,N_16105,N_16148);
nor U17508 (N_17508,N_16695,N_16058);
or U17509 (N_17509,N_16100,N_16504);
nor U17510 (N_17510,N_16068,N_16321);
nand U17511 (N_17511,N_16171,N_16734);
and U17512 (N_17512,N_16279,N_16735);
xor U17513 (N_17513,N_16092,N_16623);
nand U17514 (N_17514,N_16081,N_16682);
nand U17515 (N_17515,N_16180,N_16532);
nand U17516 (N_17516,N_16183,N_16169);
nand U17517 (N_17517,N_16254,N_16761);
nand U17518 (N_17518,N_16646,N_16396);
and U17519 (N_17519,N_16101,N_16405);
nand U17520 (N_17520,N_16260,N_16028);
nand U17521 (N_17521,N_16371,N_16067);
nand U17522 (N_17522,N_16328,N_16131);
xor U17523 (N_17523,N_16750,N_16406);
xor U17524 (N_17524,N_16229,N_16754);
nor U17525 (N_17525,N_16017,N_16792);
and U17526 (N_17526,N_16277,N_16541);
nand U17527 (N_17527,N_16056,N_16573);
and U17528 (N_17528,N_16181,N_16560);
nor U17529 (N_17529,N_16029,N_16460);
xnor U17530 (N_17530,N_16756,N_16420);
or U17531 (N_17531,N_16363,N_16039);
or U17532 (N_17532,N_16654,N_16773);
or U17533 (N_17533,N_16431,N_16651);
or U17534 (N_17534,N_16100,N_16073);
xor U17535 (N_17535,N_16069,N_16078);
and U17536 (N_17536,N_16732,N_16358);
nand U17537 (N_17537,N_16300,N_16295);
or U17538 (N_17538,N_16381,N_16445);
nand U17539 (N_17539,N_16668,N_16395);
and U17540 (N_17540,N_16650,N_16594);
nand U17541 (N_17541,N_16219,N_16185);
nor U17542 (N_17542,N_16189,N_16059);
xor U17543 (N_17543,N_16188,N_16493);
or U17544 (N_17544,N_16050,N_16305);
and U17545 (N_17545,N_16172,N_16240);
and U17546 (N_17546,N_16059,N_16473);
nor U17547 (N_17547,N_16674,N_16471);
nand U17548 (N_17548,N_16052,N_16501);
nor U17549 (N_17549,N_16250,N_16239);
xnor U17550 (N_17550,N_16620,N_16577);
nor U17551 (N_17551,N_16023,N_16558);
nor U17552 (N_17552,N_16284,N_16054);
xnor U17553 (N_17553,N_16645,N_16307);
nor U17554 (N_17554,N_16404,N_16525);
nand U17555 (N_17555,N_16010,N_16177);
or U17556 (N_17556,N_16461,N_16609);
xor U17557 (N_17557,N_16588,N_16391);
nand U17558 (N_17558,N_16183,N_16678);
or U17559 (N_17559,N_16384,N_16057);
or U17560 (N_17560,N_16176,N_16627);
nor U17561 (N_17561,N_16744,N_16451);
or U17562 (N_17562,N_16268,N_16385);
nand U17563 (N_17563,N_16592,N_16227);
nor U17564 (N_17564,N_16394,N_16287);
or U17565 (N_17565,N_16737,N_16047);
nand U17566 (N_17566,N_16229,N_16650);
nand U17567 (N_17567,N_16268,N_16570);
xnor U17568 (N_17568,N_16349,N_16298);
nor U17569 (N_17569,N_16669,N_16516);
nand U17570 (N_17570,N_16050,N_16115);
nand U17571 (N_17571,N_16421,N_16406);
nor U17572 (N_17572,N_16751,N_16270);
and U17573 (N_17573,N_16049,N_16417);
or U17574 (N_17574,N_16354,N_16177);
and U17575 (N_17575,N_16391,N_16002);
xnor U17576 (N_17576,N_16285,N_16256);
or U17577 (N_17577,N_16022,N_16389);
nor U17578 (N_17578,N_16473,N_16205);
nand U17579 (N_17579,N_16566,N_16415);
or U17580 (N_17580,N_16473,N_16351);
xor U17581 (N_17581,N_16706,N_16152);
nor U17582 (N_17582,N_16100,N_16576);
nor U17583 (N_17583,N_16117,N_16142);
or U17584 (N_17584,N_16526,N_16288);
and U17585 (N_17585,N_16487,N_16129);
or U17586 (N_17586,N_16317,N_16381);
xnor U17587 (N_17587,N_16410,N_16080);
or U17588 (N_17588,N_16382,N_16675);
or U17589 (N_17589,N_16520,N_16744);
nand U17590 (N_17590,N_16617,N_16303);
and U17591 (N_17591,N_16048,N_16640);
nand U17592 (N_17592,N_16531,N_16491);
or U17593 (N_17593,N_16057,N_16254);
nor U17594 (N_17594,N_16233,N_16191);
nand U17595 (N_17595,N_16779,N_16375);
nand U17596 (N_17596,N_16354,N_16044);
and U17597 (N_17597,N_16303,N_16015);
and U17598 (N_17598,N_16049,N_16353);
nor U17599 (N_17599,N_16339,N_16648);
xnor U17600 (N_17600,N_16852,N_17525);
xor U17601 (N_17601,N_17571,N_17488);
and U17602 (N_17602,N_17458,N_17090);
and U17603 (N_17603,N_17174,N_17251);
and U17604 (N_17604,N_16969,N_17221);
nand U17605 (N_17605,N_16924,N_17404);
or U17606 (N_17606,N_17370,N_17348);
and U17607 (N_17607,N_17580,N_17529);
nor U17608 (N_17608,N_17298,N_16865);
or U17609 (N_17609,N_17585,N_16932);
nor U17610 (N_17610,N_16911,N_17475);
xor U17611 (N_17611,N_17112,N_17169);
or U17612 (N_17612,N_17422,N_17255);
nand U17613 (N_17613,N_17012,N_17390);
xor U17614 (N_17614,N_17568,N_17031);
xor U17615 (N_17615,N_17599,N_16925);
xnor U17616 (N_17616,N_17321,N_17130);
and U17617 (N_17617,N_16869,N_17444);
nor U17618 (N_17618,N_16950,N_17335);
xnor U17619 (N_17619,N_17233,N_17108);
xnor U17620 (N_17620,N_17282,N_16824);
xnor U17621 (N_17621,N_17076,N_17201);
nand U17622 (N_17622,N_17360,N_17164);
or U17623 (N_17623,N_17092,N_17582);
nor U17624 (N_17624,N_17492,N_17111);
or U17625 (N_17625,N_17554,N_17392);
or U17626 (N_17626,N_17426,N_17096);
nor U17627 (N_17627,N_16981,N_17354);
and U17628 (N_17628,N_17350,N_17095);
nor U17629 (N_17629,N_17474,N_16933);
and U17630 (N_17630,N_16971,N_17218);
and U17631 (N_17631,N_17119,N_16816);
nand U17632 (N_17632,N_17516,N_17094);
nand U17633 (N_17633,N_17132,N_17099);
xnor U17634 (N_17634,N_16917,N_17195);
nor U17635 (N_17635,N_16850,N_17377);
nand U17636 (N_17636,N_16980,N_17100);
nor U17637 (N_17637,N_17328,N_16835);
xnor U17638 (N_17638,N_16934,N_17334);
nand U17639 (N_17639,N_16944,N_16918);
xor U17640 (N_17640,N_16817,N_16949);
or U17641 (N_17641,N_16825,N_16939);
or U17642 (N_17642,N_17534,N_17331);
nor U17643 (N_17643,N_16879,N_17441);
nor U17644 (N_17644,N_17013,N_17170);
xnor U17645 (N_17645,N_16913,N_17546);
and U17646 (N_17646,N_17409,N_17081);
nand U17647 (N_17647,N_17087,N_17461);
xor U17648 (N_17648,N_16901,N_17540);
nor U17649 (N_17649,N_17155,N_17439);
nand U17650 (N_17650,N_17598,N_16912);
nand U17651 (N_17651,N_16866,N_17402);
or U17652 (N_17652,N_16800,N_16877);
or U17653 (N_17653,N_17583,N_17339);
nand U17654 (N_17654,N_16900,N_16998);
nor U17655 (N_17655,N_17269,N_17501);
xnor U17656 (N_17656,N_17210,N_17032);
and U17657 (N_17657,N_17594,N_17188);
or U17658 (N_17658,N_17535,N_17347);
nor U17659 (N_17659,N_17427,N_17121);
or U17660 (N_17660,N_17225,N_17105);
xnor U17661 (N_17661,N_17468,N_17091);
or U17662 (N_17662,N_17143,N_17485);
xnor U17663 (N_17663,N_16831,N_17460);
and U17664 (N_17664,N_16953,N_17406);
or U17665 (N_17665,N_17234,N_17035);
nand U17666 (N_17666,N_17093,N_17122);
nor U17667 (N_17667,N_17559,N_17489);
xor U17668 (N_17668,N_17504,N_17002);
or U17669 (N_17669,N_16826,N_17068);
and U17670 (N_17670,N_17048,N_17053);
nand U17671 (N_17671,N_16996,N_17576);
xor U17672 (N_17672,N_17246,N_17072);
and U17673 (N_17673,N_17301,N_16887);
xnor U17674 (N_17674,N_17189,N_17033);
nor U17675 (N_17675,N_17472,N_16837);
xor U17676 (N_17676,N_17179,N_16952);
nand U17677 (N_17677,N_17393,N_17565);
and U17678 (N_17678,N_17456,N_17366);
nand U17679 (N_17679,N_17553,N_17476);
nand U17680 (N_17680,N_17268,N_17413);
and U17681 (N_17681,N_16848,N_17544);
nor U17682 (N_17682,N_17541,N_17587);
or U17683 (N_17683,N_17500,N_17300);
nor U17684 (N_17684,N_17001,N_17308);
nor U17685 (N_17685,N_17363,N_16903);
nand U17686 (N_17686,N_17004,N_17141);
and U17687 (N_17687,N_17177,N_16937);
and U17688 (N_17688,N_16841,N_17327);
nor U17689 (N_17689,N_16859,N_17579);
nor U17690 (N_17690,N_17262,N_17223);
nor U17691 (N_17691,N_17447,N_16878);
or U17692 (N_17692,N_17584,N_17482);
nor U17693 (N_17693,N_17523,N_17103);
xor U17694 (N_17694,N_17396,N_16814);
xnor U17695 (N_17695,N_17556,N_16987);
nor U17696 (N_17696,N_17333,N_17527);
and U17697 (N_17697,N_17136,N_17232);
and U17698 (N_17698,N_17054,N_16983);
xor U17699 (N_17699,N_17542,N_17397);
nor U17700 (N_17700,N_16965,N_17137);
nand U17701 (N_17701,N_17416,N_17520);
nand U17702 (N_17702,N_16957,N_17345);
nand U17703 (N_17703,N_17290,N_17168);
nand U17704 (N_17704,N_17320,N_17277);
nand U17705 (N_17705,N_17346,N_16893);
or U17706 (N_17706,N_17185,N_17182);
nor U17707 (N_17707,N_17293,N_17196);
nand U17708 (N_17708,N_17212,N_17593);
nor U17709 (N_17709,N_17551,N_16976);
xnor U17710 (N_17710,N_17569,N_17371);
nand U17711 (N_17711,N_16858,N_16875);
and U17712 (N_17712,N_17278,N_17515);
and U17713 (N_17713,N_17537,N_16884);
nor U17714 (N_17714,N_17194,N_17059);
nor U17715 (N_17715,N_16919,N_16802);
or U17716 (N_17716,N_16829,N_17432);
xor U17717 (N_17717,N_17040,N_17131);
nor U17718 (N_17718,N_17307,N_17052);
and U17719 (N_17719,N_17419,N_17249);
nand U17720 (N_17720,N_17027,N_17271);
xor U17721 (N_17721,N_17358,N_17330);
and U17722 (N_17722,N_17086,N_16982);
nand U17723 (N_17723,N_17424,N_17592);
or U17724 (N_17724,N_17317,N_16871);
nand U17725 (N_17725,N_17502,N_16992);
nand U17726 (N_17726,N_17057,N_17299);
and U17727 (N_17727,N_17442,N_16991);
xnor U17728 (N_17728,N_17467,N_17231);
nand U17729 (N_17729,N_17288,N_16897);
xor U17730 (N_17730,N_17499,N_17379);
nor U17731 (N_17731,N_17250,N_17047);
and U17732 (N_17732,N_16986,N_17563);
xor U17733 (N_17733,N_16895,N_16896);
nand U17734 (N_17734,N_17267,N_17236);
or U17735 (N_17735,N_17016,N_17158);
nor U17736 (N_17736,N_17566,N_17311);
and U17737 (N_17737,N_17483,N_17226);
xor U17738 (N_17738,N_17386,N_17443);
xor U17739 (N_17739,N_17437,N_16885);
or U17740 (N_17740,N_17157,N_17058);
nor U17741 (N_17741,N_16938,N_17110);
xnor U17742 (N_17742,N_17166,N_17552);
nor U17743 (N_17743,N_17506,N_16929);
xnor U17744 (N_17744,N_17147,N_16993);
and U17745 (N_17745,N_17149,N_17503);
nor U17746 (N_17746,N_17391,N_17146);
nor U17747 (N_17747,N_17340,N_17211);
xnor U17748 (N_17748,N_17056,N_16973);
xnor U17749 (N_17749,N_17558,N_17316);
and U17750 (N_17750,N_17193,N_17264);
nor U17751 (N_17751,N_16943,N_17043);
or U17752 (N_17752,N_17548,N_17509);
nand U17753 (N_17753,N_16836,N_17285);
or U17754 (N_17754,N_17570,N_17038);
nand U17755 (N_17755,N_17434,N_17309);
nor U17756 (N_17756,N_17270,N_17303);
nor U17757 (N_17757,N_17517,N_17577);
nor U17758 (N_17758,N_17549,N_17042);
nand U17759 (N_17759,N_17411,N_17152);
or U17760 (N_17760,N_17009,N_16898);
or U17761 (N_17761,N_17524,N_17050);
nand U17762 (N_17762,N_16926,N_16923);
nor U17763 (N_17763,N_17011,N_17315);
nor U17764 (N_17764,N_17313,N_17597);
nand U17765 (N_17765,N_16935,N_16979);
and U17766 (N_17766,N_17238,N_17245);
nand U17767 (N_17767,N_16974,N_17590);
nor U17768 (N_17768,N_16988,N_17470);
nor U17769 (N_17769,N_17428,N_17162);
xor U17770 (N_17770,N_17254,N_17528);
xnor U17771 (N_17771,N_17046,N_17202);
and U17772 (N_17772,N_17248,N_17319);
nand U17773 (N_17773,N_17414,N_17055);
and U17774 (N_17774,N_17167,N_17505);
and U17775 (N_17775,N_17260,N_16851);
or U17776 (N_17776,N_17003,N_17224);
or U17777 (N_17777,N_17464,N_17065);
and U17778 (N_17778,N_16854,N_16855);
and U17779 (N_17779,N_17265,N_16927);
nor U17780 (N_17780,N_17097,N_17425);
and U17781 (N_17781,N_17532,N_16963);
or U17782 (N_17782,N_16872,N_16922);
xnor U17783 (N_17783,N_16916,N_16806);
and U17784 (N_17784,N_17395,N_17030);
xnor U17785 (N_17785,N_16815,N_17436);
nor U17786 (N_17786,N_17399,N_16968);
or U17787 (N_17787,N_17586,N_16847);
nor U17788 (N_17788,N_17230,N_17306);
or U17789 (N_17789,N_17186,N_17508);
and U17790 (N_17790,N_17036,N_17114);
or U17791 (N_17791,N_17173,N_17385);
nor U17792 (N_17792,N_17102,N_17061);
xor U17793 (N_17793,N_16906,N_17295);
nand U17794 (N_17794,N_16890,N_16962);
nand U17795 (N_17795,N_16989,N_17589);
xnor U17796 (N_17796,N_16834,N_16830);
nand U17797 (N_17797,N_17337,N_17024);
and U17798 (N_17798,N_17291,N_17420);
or U17799 (N_17799,N_16945,N_17342);
xor U17800 (N_17800,N_17326,N_17417);
and U17801 (N_17801,N_16964,N_17204);
nor U17802 (N_17802,N_16818,N_17244);
nor U17803 (N_17803,N_17010,N_17338);
or U17804 (N_17804,N_17187,N_17486);
xnor U17805 (N_17805,N_17477,N_17365);
nor U17806 (N_17806,N_17261,N_16921);
nor U17807 (N_17807,N_16857,N_16819);
nand U17808 (N_17808,N_17478,N_17324);
nand U17809 (N_17809,N_17421,N_17165);
and U17810 (N_17810,N_17150,N_17567);
nor U17811 (N_17811,N_17557,N_17418);
and U17812 (N_17812,N_16881,N_16880);
nand U17813 (N_17813,N_16864,N_17560);
xnor U17814 (N_17814,N_17355,N_17382);
nand U17815 (N_17815,N_17550,N_17521);
xor U17816 (N_17816,N_17466,N_17106);
and U17817 (N_17817,N_17332,N_17219);
and U17818 (N_17818,N_17180,N_17148);
nor U17819 (N_17819,N_17286,N_17533);
xnor U17820 (N_17820,N_17575,N_17343);
nor U17821 (N_17821,N_17394,N_17435);
nor U17822 (N_17822,N_16889,N_17116);
xor U17823 (N_17823,N_16842,N_17017);
nor U17824 (N_17824,N_17401,N_16808);
xor U17825 (N_17825,N_17539,N_17075);
nor U17826 (N_17826,N_17430,N_17257);
or U17827 (N_17827,N_17138,N_17198);
nand U17828 (N_17828,N_17304,N_17274);
nor U17829 (N_17829,N_16977,N_17214);
and U17830 (N_17830,N_17019,N_17127);
and U17831 (N_17831,N_17083,N_17514);
or U17832 (N_17832,N_17595,N_16801);
nand U17833 (N_17833,N_17135,N_17453);
or U17834 (N_17834,N_17410,N_17247);
nor U17835 (N_17835,N_16955,N_17438);
nand U17836 (N_17836,N_17465,N_17373);
or U17837 (N_17837,N_17353,N_17028);
nor U17838 (N_17838,N_17263,N_17536);
xor U17839 (N_17839,N_17071,N_17215);
xor U17840 (N_17840,N_16905,N_16860);
nand U17841 (N_17841,N_17006,N_17118);
xnor U17842 (N_17842,N_17126,N_17491);
or U17843 (N_17843,N_17125,N_17082);
nand U17844 (N_17844,N_17000,N_17412);
and U17845 (N_17845,N_17423,N_17120);
or U17846 (N_17846,N_17449,N_17151);
nand U17847 (N_17847,N_17085,N_17561);
or U17848 (N_17848,N_17243,N_17213);
xnor U17849 (N_17849,N_17511,N_17596);
nor U17850 (N_17850,N_17279,N_17239);
nand U17851 (N_17851,N_16915,N_17258);
xor U17852 (N_17852,N_17044,N_17415);
nand U17853 (N_17853,N_17176,N_17161);
or U17854 (N_17854,N_17578,N_17266);
nor U17855 (N_17855,N_16894,N_16822);
or U17856 (N_17856,N_17113,N_17369);
and U17857 (N_17857,N_17495,N_17172);
xor U17858 (N_17858,N_17220,N_17440);
xor U17859 (N_17859,N_17314,N_17356);
xor U17860 (N_17860,N_17387,N_17153);
nand U17861 (N_17861,N_16812,N_17216);
and U17862 (N_17862,N_16823,N_17341);
xor U17863 (N_17863,N_16868,N_17513);
xnor U17864 (N_17864,N_17374,N_16930);
nand U17865 (N_17865,N_16967,N_17088);
nand U17866 (N_17866,N_17252,N_17007);
xnor U17867 (N_17867,N_17455,N_17389);
and U17868 (N_17868,N_16804,N_17322);
xnor U17869 (N_17869,N_16892,N_17140);
and U17870 (N_17870,N_17543,N_17496);
or U17871 (N_17871,N_17256,N_16863);
nand U17872 (N_17872,N_17227,N_17450);
nor U17873 (N_17873,N_16948,N_16886);
or U17874 (N_17874,N_16839,N_17429);
or U17875 (N_17875,N_17545,N_17318);
and U17876 (N_17876,N_17296,N_17124);
nand U17877 (N_17877,N_17005,N_16909);
nand U17878 (N_17878,N_17388,N_17175);
or U17879 (N_17879,N_17273,N_17519);
or U17880 (N_17880,N_17206,N_16994);
and U17881 (N_17881,N_17408,N_17357);
or U17882 (N_17882,N_16845,N_17183);
nor U17883 (N_17883,N_17159,N_17015);
nand U17884 (N_17884,N_16972,N_17446);
nor U17885 (N_17885,N_17208,N_17361);
nand U17886 (N_17886,N_17115,N_17041);
nor U17887 (N_17887,N_17139,N_17284);
and U17888 (N_17888,N_17021,N_17574);
or U17889 (N_17889,N_17022,N_17289);
and U17890 (N_17890,N_17479,N_17134);
and U17891 (N_17891,N_17078,N_17084);
and U17892 (N_17892,N_17351,N_17445);
nand U17893 (N_17893,N_17480,N_17008);
nor U17894 (N_17894,N_16960,N_16861);
nand U17895 (N_17895,N_17462,N_17171);
or U17896 (N_17896,N_17481,N_17302);
nand U17897 (N_17897,N_17512,N_17229);
or U17898 (N_17898,N_16947,N_17433);
nand U17899 (N_17899,N_16844,N_16999);
xnor U17900 (N_17900,N_17259,N_16961);
nor U17901 (N_17901,N_17184,N_16920);
nor U17902 (N_17902,N_16853,N_17142);
nor U17903 (N_17903,N_17497,N_16820);
and U17904 (N_17904,N_17240,N_16902);
and U17905 (N_17905,N_17192,N_16941);
nor U17906 (N_17906,N_16928,N_17060);
or U17907 (N_17907,N_16870,N_17469);
or U17908 (N_17908,N_17372,N_17063);
xor U17909 (N_17909,N_17381,N_17080);
nor U17910 (N_17910,N_16908,N_17237);
nor U17911 (N_17911,N_17484,N_17473);
or U17912 (N_17912,N_17518,N_17283);
nand U17913 (N_17913,N_17564,N_17375);
xor U17914 (N_17914,N_17026,N_17209);
nor U17915 (N_17915,N_17181,N_17281);
nor U17916 (N_17916,N_17359,N_17384);
xor U17917 (N_17917,N_17066,N_17522);
xnor U17918 (N_17918,N_16984,N_17197);
xor U17919 (N_17919,N_17029,N_17378);
nor U17920 (N_17920,N_17051,N_17275);
or U17921 (N_17921,N_17368,N_17156);
nand U17922 (N_17922,N_17217,N_16813);
xor U17923 (N_17923,N_17272,N_17325);
xnor U17924 (N_17924,N_17154,N_16946);
or U17925 (N_17925,N_17023,N_17448);
and U17926 (N_17926,N_16810,N_16832);
and U17927 (N_17927,N_17045,N_17538);
nor U17928 (N_17928,N_16856,N_16931);
xor U17929 (N_17929,N_16914,N_17352);
nor U17930 (N_17930,N_16975,N_17280);
nand U17931 (N_17931,N_17487,N_17064);
xnor U17932 (N_17932,N_16849,N_16838);
nor U17933 (N_17933,N_17200,N_17588);
nand U17934 (N_17934,N_17203,N_16828);
xor U17935 (N_17935,N_17025,N_17376);
or U17936 (N_17936,N_16990,N_16891);
or U17937 (N_17937,N_16840,N_17109);
or U17938 (N_17938,N_16958,N_16956);
nand U17939 (N_17939,N_17190,N_17494);
or U17940 (N_17940,N_17160,N_16809);
xor U17941 (N_17941,N_17241,N_17312);
nand U17942 (N_17942,N_16873,N_16985);
nand U17943 (N_17943,N_17128,N_16833);
nor U17944 (N_17944,N_16959,N_16995);
and U17945 (N_17945,N_17510,N_17098);
nand U17946 (N_17946,N_17431,N_17457);
or U17947 (N_17947,N_16876,N_17530);
nand U17948 (N_17948,N_17362,N_16940);
and U17949 (N_17949,N_17133,N_16997);
xnor U17950 (N_17950,N_17235,N_16807);
or U17951 (N_17951,N_17400,N_17531);
and U17952 (N_17952,N_17039,N_17049);
xor U17953 (N_17953,N_17207,N_17073);
nor U17954 (N_17954,N_16951,N_17079);
nand U17955 (N_17955,N_17367,N_17129);
nand U17956 (N_17956,N_17305,N_16811);
and U17957 (N_17957,N_17323,N_16936);
nor U17958 (N_17958,N_17222,N_17364);
and U17959 (N_17959,N_16907,N_17242);
xnor U17960 (N_17960,N_16805,N_17507);
xor U17961 (N_17961,N_17077,N_17178);
or U17962 (N_17962,N_16843,N_16910);
xnor U17963 (N_17963,N_16867,N_17020);
and U17964 (N_17964,N_17037,N_17526);
or U17965 (N_17965,N_17069,N_17228);
nand U17966 (N_17966,N_17463,N_17349);
nand U17967 (N_17967,N_17451,N_17070);
and U17968 (N_17968,N_17034,N_17336);
nand U17969 (N_17969,N_17581,N_17383);
nand U17970 (N_17970,N_17205,N_17555);
nor U17971 (N_17971,N_17403,N_17573);
nand U17972 (N_17972,N_16882,N_17107);
nand U17973 (N_17973,N_16874,N_17329);
nor U17974 (N_17974,N_17067,N_17498);
and U17975 (N_17975,N_16883,N_17253);
xor U17976 (N_17976,N_17089,N_17380);
and U17977 (N_17977,N_17591,N_17310);
xor U17978 (N_17978,N_17344,N_17287);
nand U17979 (N_17979,N_16904,N_17547);
or U17980 (N_17980,N_16899,N_16970);
or U17981 (N_17981,N_16954,N_17276);
xnor U17982 (N_17982,N_17062,N_16827);
nand U17983 (N_17983,N_16888,N_17018);
nand U17984 (N_17984,N_17297,N_16966);
or U17985 (N_17985,N_17572,N_17471);
and U17986 (N_17986,N_17493,N_17294);
nor U17987 (N_17987,N_16821,N_16942);
or U17988 (N_17988,N_17014,N_16862);
and U17989 (N_17989,N_17452,N_17163);
and U17990 (N_17990,N_17398,N_17117);
and U17991 (N_17991,N_17145,N_17459);
nand U17992 (N_17992,N_17407,N_17123);
or U17993 (N_17993,N_17562,N_17104);
xnor U17994 (N_17994,N_17490,N_17454);
and U17995 (N_17995,N_16846,N_17101);
xor U17996 (N_17996,N_17074,N_17144);
nand U17997 (N_17997,N_16803,N_17199);
nor U17998 (N_17998,N_17405,N_16978);
or U17999 (N_17999,N_17292,N_17191);
nor U18000 (N_18000,N_17390,N_17089);
nor U18001 (N_18001,N_17348,N_17563);
nor U18002 (N_18002,N_17414,N_17186);
xnor U18003 (N_18003,N_17222,N_17085);
nor U18004 (N_18004,N_16970,N_17298);
nor U18005 (N_18005,N_17176,N_17480);
nor U18006 (N_18006,N_17416,N_17567);
nor U18007 (N_18007,N_17585,N_16943);
nand U18008 (N_18008,N_17349,N_16804);
or U18009 (N_18009,N_17586,N_16918);
nor U18010 (N_18010,N_16928,N_16929);
nand U18011 (N_18011,N_17127,N_17436);
nand U18012 (N_18012,N_16889,N_17112);
xor U18013 (N_18013,N_17060,N_17023);
xnor U18014 (N_18014,N_17416,N_17082);
nand U18015 (N_18015,N_17287,N_17398);
nand U18016 (N_18016,N_16974,N_17500);
and U18017 (N_18017,N_16849,N_16830);
or U18018 (N_18018,N_16977,N_17122);
nand U18019 (N_18019,N_16816,N_17462);
and U18020 (N_18020,N_16824,N_16843);
nor U18021 (N_18021,N_16837,N_16830);
and U18022 (N_18022,N_17473,N_17576);
or U18023 (N_18023,N_17546,N_17464);
and U18024 (N_18024,N_16846,N_16960);
nand U18025 (N_18025,N_16879,N_17404);
nor U18026 (N_18026,N_17191,N_17039);
or U18027 (N_18027,N_16976,N_17188);
and U18028 (N_18028,N_17267,N_17424);
and U18029 (N_18029,N_17287,N_16928);
or U18030 (N_18030,N_17060,N_17355);
or U18031 (N_18031,N_17405,N_17170);
nand U18032 (N_18032,N_16824,N_17155);
and U18033 (N_18033,N_17209,N_17132);
or U18034 (N_18034,N_17152,N_17056);
xor U18035 (N_18035,N_17390,N_17315);
nor U18036 (N_18036,N_16881,N_17220);
or U18037 (N_18037,N_17299,N_17240);
nand U18038 (N_18038,N_16993,N_17519);
and U18039 (N_18039,N_17455,N_17230);
nand U18040 (N_18040,N_17206,N_17293);
nand U18041 (N_18041,N_16993,N_17407);
nor U18042 (N_18042,N_17294,N_17202);
and U18043 (N_18043,N_16920,N_17185);
or U18044 (N_18044,N_16991,N_17061);
or U18045 (N_18045,N_16915,N_17043);
or U18046 (N_18046,N_16994,N_17339);
nand U18047 (N_18047,N_17286,N_17037);
nor U18048 (N_18048,N_17597,N_17570);
nor U18049 (N_18049,N_17165,N_17128);
nor U18050 (N_18050,N_17165,N_17313);
nand U18051 (N_18051,N_17469,N_17244);
or U18052 (N_18052,N_16890,N_17111);
or U18053 (N_18053,N_17531,N_17184);
or U18054 (N_18054,N_16960,N_17369);
nand U18055 (N_18055,N_17123,N_16807);
and U18056 (N_18056,N_16961,N_16857);
nand U18057 (N_18057,N_17224,N_17458);
nand U18058 (N_18058,N_17516,N_17014);
nand U18059 (N_18059,N_16873,N_17369);
nand U18060 (N_18060,N_16967,N_16988);
or U18061 (N_18061,N_16971,N_17131);
xnor U18062 (N_18062,N_17134,N_16867);
nand U18063 (N_18063,N_16867,N_17493);
nand U18064 (N_18064,N_16871,N_17048);
nand U18065 (N_18065,N_17210,N_17562);
nand U18066 (N_18066,N_17286,N_17433);
or U18067 (N_18067,N_17034,N_17296);
or U18068 (N_18068,N_17510,N_17085);
or U18069 (N_18069,N_17128,N_17433);
and U18070 (N_18070,N_17397,N_17439);
nor U18071 (N_18071,N_17429,N_17572);
nor U18072 (N_18072,N_17165,N_17571);
nor U18073 (N_18073,N_17049,N_17500);
or U18074 (N_18074,N_17298,N_17556);
and U18075 (N_18075,N_17009,N_16968);
nor U18076 (N_18076,N_17339,N_17076);
and U18077 (N_18077,N_17318,N_17205);
nand U18078 (N_18078,N_17090,N_17569);
nand U18079 (N_18079,N_17384,N_17564);
and U18080 (N_18080,N_17535,N_17331);
nor U18081 (N_18081,N_17099,N_17326);
xnor U18082 (N_18082,N_17203,N_17429);
nand U18083 (N_18083,N_17318,N_17157);
or U18084 (N_18084,N_16888,N_17528);
and U18085 (N_18085,N_17367,N_17332);
or U18086 (N_18086,N_17138,N_17305);
nor U18087 (N_18087,N_17395,N_17187);
nor U18088 (N_18088,N_17332,N_16947);
nor U18089 (N_18089,N_17398,N_16987);
nor U18090 (N_18090,N_17025,N_16803);
nor U18091 (N_18091,N_17168,N_17169);
or U18092 (N_18092,N_17096,N_17136);
nor U18093 (N_18093,N_17121,N_17273);
and U18094 (N_18094,N_17381,N_17254);
xor U18095 (N_18095,N_17239,N_17465);
nand U18096 (N_18096,N_17213,N_17473);
nand U18097 (N_18097,N_17448,N_17450);
xnor U18098 (N_18098,N_17220,N_16813);
or U18099 (N_18099,N_17571,N_17205);
nor U18100 (N_18100,N_17221,N_17328);
nor U18101 (N_18101,N_17368,N_17080);
xnor U18102 (N_18102,N_17061,N_16904);
or U18103 (N_18103,N_17126,N_17208);
nand U18104 (N_18104,N_17599,N_17124);
nand U18105 (N_18105,N_17541,N_17422);
nor U18106 (N_18106,N_17187,N_17421);
and U18107 (N_18107,N_16836,N_17024);
and U18108 (N_18108,N_17498,N_17564);
nor U18109 (N_18109,N_17310,N_17459);
xor U18110 (N_18110,N_17414,N_17023);
or U18111 (N_18111,N_17325,N_17249);
xnor U18112 (N_18112,N_17517,N_17433);
or U18113 (N_18113,N_17053,N_17062);
nand U18114 (N_18114,N_17076,N_17597);
and U18115 (N_18115,N_17029,N_17597);
nand U18116 (N_18116,N_16958,N_17521);
and U18117 (N_18117,N_17000,N_17052);
and U18118 (N_18118,N_17287,N_17595);
and U18119 (N_18119,N_17097,N_17421);
xnor U18120 (N_18120,N_17053,N_16908);
xnor U18121 (N_18121,N_17299,N_16861);
nor U18122 (N_18122,N_17210,N_17413);
xor U18123 (N_18123,N_17219,N_17595);
or U18124 (N_18124,N_17331,N_17171);
nor U18125 (N_18125,N_17190,N_17411);
and U18126 (N_18126,N_17217,N_17136);
nand U18127 (N_18127,N_17345,N_16815);
nor U18128 (N_18128,N_17522,N_17339);
or U18129 (N_18129,N_17328,N_17468);
nor U18130 (N_18130,N_16886,N_17030);
xor U18131 (N_18131,N_17363,N_17421);
nor U18132 (N_18132,N_17420,N_17158);
nor U18133 (N_18133,N_17355,N_17465);
and U18134 (N_18134,N_17286,N_17301);
nand U18135 (N_18135,N_17298,N_17591);
nor U18136 (N_18136,N_16814,N_16836);
or U18137 (N_18137,N_16887,N_16881);
nand U18138 (N_18138,N_17541,N_17548);
xnor U18139 (N_18139,N_17308,N_16993);
nand U18140 (N_18140,N_17276,N_17252);
nand U18141 (N_18141,N_17506,N_17490);
and U18142 (N_18142,N_17090,N_17396);
nor U18143 (N_18143,N_17227,N_17306);
nor U18144 (N_18144,N_16869,N_17142);
xor U18145 (N_18145,N_17055,N_17464);
xnor U18146 (N_18146,N_16902,N_16887);
and U18147 (N_18147,N_16894,N_16881);
xor U18148 (N_18148,N_17577,N_17555);
and U18149 (N_18149,N_17186,N_17209);
xnor U18150 (N_18150,N_17548,N_17127);
or U18151 (N_18151,N_17583,N_17514);
or U18152 (N_18152,N_17515,N_17192);
or U18153 (N_18153,N_17588,N_17234);
xor U18154 (N_18154,N_17348,N_17111);
and U18155 (N_18155,N_17090,N_16936);
and U18156 (N_18156,N_17132,N_17363);
or U18157 (N_18157,N_16982,N_16889);
and U18158 (N_18158,N_17132,N_17245);
or U18159 (N_18159,N_17593,N_17247);
nor U18160 (N_18160,N_17411,N_17287);
xnor U18161 (N_18161,N_17586,N_17173);
nand U18162 (N_18162,N_16846,N_17102);
nor U18163 (N_18163,N_17379,N_16890);
or U18164 (N_18164,N_17456,N_17527);
xor U18165 (N_18165,N_16881,N_16842);
nand U18166 (N_18166,N_16864,N_17537);
nor U18167 (N_18167,N_16831,N_17543);
and U18168 (N_18168,N_16927,N_16948);
and U18169 (N_18169,N_17586,N_17156);
nand U18170 (N_18170,N_17400,N_16949);
nand U18171 (N_18171,N_17547,N_17131);
or U18172 (N_18172,N_16852,N_17010);
nor U18173 (N_18173,N_17467,N_16930);
nand U18174 (N_18174,N_17316,N_16939);
xor U18175 (N_18175,N_17009,N_17003);
xnor U18176 (N_18176,N_17528,N_17585);
xor U18177 (N_18177,N_17313,N_17178);
or U18178 (N_18178,N_17586,N_16903);
or U18179 (N_18179,N_17263,N_16987);
xor U18180 (N_18180,N_17295,N_16939);
or U18181 (N_18181,N_17228,N_17293);
and U18182 (N_18182,N_16907,N_17071);
xor U18183 (N_18183,N_17546,N_17592);
nand U18184 (N_18184,N_17039,N_17260);
nor U18185 (N_18185,N_17444,N_17473);
and U18186 (N_18186,N_17478,N_17402);
or U18187 (N_18187,N_17540,N_17035);
or U18188 (N_18188,N_16854,N_16961);
xor U18189 (N_18189,N_17479,N_17491);
nor U18190 (N_18190,N_17295,N_17129);
nor U18191 (N_18191,N_16993,N_17376);
and U18192 (N_18192,N_17297,N_17585);
and U18193 (N_18193,N_17413,N_17013);
nor U18194 (N_18194,N_17059,N_17130);
or U18195 (N_18195,N_16915,N_17388);
xor U18196 (N_18196,N_17322,N_17312);
and U18197 (N_18197,N_16902,N_17132);
and U18198 (N_18198,N_16838,N_16856);
nand U18199 (N_18199,N_17406,N_17301);
nand U18200 (N_18200,N_17489,N_17302);
nor U18201 (N_18201,N_16814,N_17034);
xnor U18202 (N_18202,N_17437,N_17263);
nor U18203 (N_18203,N_17330,N_17250);
xnor U18204 (N_18204,N_17194,N_17271);
xnor U18205 (N_18205,N_16834,N_16840);
nand U18206 (N_18206,N_17486,N_17324);
or U18207 (N_18207,N_17557,N_17042);
and U18208 (N_18208,N_17507,N_17042);
or U18209 (N_18209,N_16804,N_17365);
nand U18210 (N_18210,N_17426,N_17441);
or U18211 (N_18211,N_17242,N_17139);
or U18212 (N_18212,N_17388,N_16899);
nor U18213 (N_18213,N_17221,N_16921);
nor U18214 (N_18214,N_16942,N_16827);
and U18215 (N_18215,N_16856,N_17598);
and U18216 (N_18216,N_17485,N_17238);
nand U18217 (N_18217,N_16990,N_16868);
nor U18218 (N_18218,N_16807,N_17328);
and U18219 (N_18219,N_17076,N_17131);
nor U18220 (N_18220,N_17002,N_17362);
nor U18221 (N_18221,N_17518,N_17089);
or U18222 (N_18222,N_16846,N_16938);
xor U18223 (N_18223,N_17325,N_17075);
xor U18224 (N_18224,N_16810,N_17233);
nand U18225 (N_18225,N_17246,N_16923);
nand U18226 (N_18226,N_16841,N_17395);
xor U18227 (N_18227,N_17330,N_17272);
xnor U18228 (N_18228,N_17532,N_17133);
and U18229 (N_18229,N_16872,N_17056);
and U18230 (N_18230,N_16891,N_17368);
nor U18231 (N_18231,N_17421,N_17194);
nor U18232 (N_18232,N_16815,N_17264);
and U18233 (N_18233,N_16915,N_16831);
and U18234 (N_18234,N_16810,N_17064);
and U18235 (N_18235,N_17188,N_17143);
and U18236 (N_18236,N_17170,N_16897);
nand U18237 (N_18237,N_17090,N_17500);
xor U18238 (N_18238,N_17468,N_17523);
nand U18239 (N_18239,N_17045,N_17244);
or U18240 (N_18240,N_17415,N_17450);
or U18241 (N_18241,N_16973,N_17518);
nand U18242 (N_18242,N_17197,N_17366);
or U18243 (N_18243,N_17340,N_16827);
and U18244 (N_18244,N_16966,N_17394);
or U18245 (N_18245,N_17581,N_17488);
or U18246 (N_18246,N_17184,N_17578);
nor U18247 (N_18247,N_17204,N_17066);
nor U18248 (N_18248,N_17004,N_17080);
nand U18249 (N_18249,N_17056,N_17016);
or U18250 (N_18250,N_17463,N_17277);
xor U18251 (N_18251,N_17380,N_17064);
or U18252 (N_18252,N_17388,N_17503);
and U18253 (N_18253,N_17454,N_17233);
xnor U18254 (N_18254,N_17441,N_17477);
xnor U18255 (N_18255,N_17266,N_17403);
xnor U18256 (N_18256,N_17114,N_16993);
nand U18257 (N_18257,N_16843,N_17489);
and U18258 (N_18258,N_16902,N_17259);
or U18259 (N_18259,N_17303,N_17469);
and U18260 (N_18260,N_16865,N_17099);
nand U18261 (N_18261,N_17266,N_17307);
or U18262 (N_18262,N_16950,N_17029);
or U18263 (N_18263,N_16853,N_17291);
xnor U18264 (N_18264,N_17223,N_16897);
xor U18265 (N_18265,N_16930,N_17249);
nand U18266 (N_18266,N_17536,N_17245);
nor U18267 (N_18267,N_17431,N_17160);
nor U18268 (N_18268,N_17565,N_17476);
nor U18269 (N_18269,N_16940,N_17599);
xnor U18270 (N_18270,N_17120,N_17191);
xnor U18271 (N_18271,N_17185,N_17313);
nor U18272 (N_18272,N_17201,N_17333);
and U18273 (N_18273,N_17109,N_17392);
nand U18274 (N_18274,N_16956,N_17238);
or U18275 (N_18275,N_17046,N_17023);
nand U18276 (N_18276,N_17157,N_17151);
and U18277 (N_18277,N_17414,N_17233);
xor U18278 (N_18278,N_17537,N_17244);
and U18279 (N_18279,N_16904,N_17077);
xnor U18280 (N_18280,N_17031,N_17412);
xor U18281 (N_18281,N_16852,N_17469);
nor U18282 (N_18282,N_17513,N_17544);
nor U18283 (N_18283,N_17284,N_17478);
xor U18284 (N_18284,N_17118,N_17507);
nand U18285 (N_18285,N_17471,N_16936);
or U18286 (N_18286,N_17035,N_17499);
xor U18287 (N_18287,N_17260,N_17267);
and U18288 (N_18288,N_17129,N_16859);
nand U18289 (N_18289,N_17421,N_17106);
xor U18290 (N_18290,N_17128,N_17402);
or U18291 (N_18291,N_17192,N_17013);
nor U18292 (N_18292,N_17170,N_17025);
xor U18293 (N_18293,N_17588,N_17371);
nor U18294 (N_18294,N_17473,N_17142);
nor U18295 (N_18295,N_17055,N_17435);
nor U18296 (N_18296,N_17248,N_17573);
nor U18297 (N_18297,N_17319,N_16848);
or U18298 (N_18298,N_17243,N_17545);
xor U18299 (N_18299,N_17532,N_17519);
or U18300 (N_18300,N_17235,N_17093);
nand U18301 (N_18301,N_16925,N_17059);
or U18302 (N_18302,N_16921,N_16989);
nand U18303 (N_18303,N_17421,N_17425);
and U18304 (N_18304,N_16806,N_17055);
xnor U18305 (N_18305,N_17521,N_16944);
xor U18306 (N_18306,N_17561,N_16800);
nand U18307 (N_18307,N_17375,N_17577);
xor U18308 (N_18308,N_17240,N_17599);
nor U18309 (N_18309,N_16946,N_17311);
xor U18310 (N_18310,N_16999,N_16957);
xnor U18311 (N_18311,N_17134,N_16914);
and U18312 (N_18312,N_17072,N_17442);
nor U18313 (N_18313,N_17219,N_17542);
or U18314 (N_18314,N_17078,N_17011);
and U18315 (N_18315,N_17425,N_17110);
nand U18316 (N_18316,N_17138,N_17590);
and U18317 (N_18317,N_17430,N_16975);
nor U18318 (N_18318,N_17528,N_17577);
nor U18319 (N_18319,N_16842,N_17587);
nand U18320 (N_18320,N_16958,N_17335);
xnor U18321 (N_18321,N_17108,N_17430);
or U18322 (N_18322,N_17374,N_16885);
nor U18323 (N_18323,N_16832,N_17392);
nand U18324 (N_18324,N_17541,N_17387);
nor U18325 (N_18325,N_17244,N_17304);
and U18326 (N_18326,N_17299,N_17143);
or U18327 (N_18327,N_17366,N_17208);
xor U18328 (N_18328,N_16838,N_17116);
nor U18329 (N_18329,N_17070,N_17389);
nor U18330 (N_18330,N_17466,N_16956);
nand U18331 (N_18331,N_17002,N_17428);
xor U18332 (N_18332,N_17542,N_17210);
xnor U18333 (N_18333,N_17246,N_17130);
or U18334 (N_18334,N_17505,N_17150);
or U18335 (N_18335,N_17533,N_17248);
xor U18336 (N_18336,N_17492,N_17108);
and U18337 (N_18337,N_16997,N_17177);
and U18338 (N_18338,N_17055,N_17513);
nor U18339 (N_18339,N_16815,N_17228);
and U18340 (N_18340,N_17003,N_16935);
or U18341 (N_18341,N_17164,N_17144);
xor U18342 (N_18342,N_17266,N_17211);
xnor U18343 (N_18343,N_16822,N_17283);
or U18344 (N_18344,N_17063,N_16904);
or U18345 (N_18345,N_17325,N_17432);
xnor U18346 (N_18346,N_17488,N_17311);
or U18347 (N_18347,N_17505,N_17195);
nand U18348 (N_18348,N_16856,N_16824);
or U18349 (N_18349,N_17180,N_17141);
nor U18350 (N_18350,N_16874,N_17147);
or U18351 (N_18351,N_17560,N_17212);
and U18352 (N_18352,N_17599,N_17069);
or U18353 (N_18353,N_17321,N_16853);
or U18354 (N_18354,N_16939,N_17509);
nor U18355 (N_18355,N_17326,N_17394);
or U18356 (N_18356,N_17113,N_16901);
and U18357 (N_18357,N_17462,N_17021);
nor U18358 (N_18358,N_17157,N_17049);
nor U18359 (N_18359,N_17591,N_17260);
nor U18360 (N_18360,N_17397,N_17205);
and U18361 (N_18361,N_17443,N_17321);
and U18362 (N_18362,N_17140,N_17160);
nand U18363 (N_18363,N_17009,N_17103);
and U18364 (N_18364,N_16864,N_17118);
nand U18365 (N_18365,N_17474,N_17370);
nor U18366 (N_18366,N_16854,N_17076);
xnor U18367 (N_18367,N_16865,N_16985);
nand U18368 (N_18368,N_17009,N_17465);
and U18369 (N_18369,N_17554,N_17176);
nor U18370 (N_18370,N_16862,N_17429);
xor U18371 (N_18371,N_17014,N_17153);
xnor U18372 (N_18372,N_17053,N_17118);
nand U18373 (N_18373,N_17590,N_16812);
xor U18374 (N_18374,N_17324,N_16991);
and U18375 (N_18375,N_16870,N_17346);
nand U18376 (N_18376,N_16844,N_17580);
nor U18377 (N_18377,N_17005,N_16876);
xnor U18378 (N_18378,N_16911,N_17442);
nand U18379 (N_18379,N_16928,N_17337);
nor U18380 (N_18380,N_16989,N_17210);
and U18381 (N_18381,N_17556,N_16864);
nand U18382 (N_18382,N_17049,N_17230);
nor U18383 (N_18383,N_17460,N_16803);
nor U18384 (N_18384,N_17428,N_17298);
nor U18385 (N_18385,N_17050,N_17146);
xor U18386 (N_18386,N_17017,N_17123);
nor U18387 (N_18387,N_17425,N_17270);
nor U18388 (N_18388,N_16806,N_16945);
or U18389 (N_18389,N_17176,N_17507);
or U18390 (N_18390,N_17139,N_17291);
nor U18391 (N_18391,N_17135,N_17256);
nand U18392 (N_18392,N_17022,N_16910);
and U18393 (N_18393,N_17409,N_17546);
and U18394 (N_18394,N_16948,N_16915);
and U18395 (N_18395,N_17153,N_17463);
nand U18396 (N_18396,N_17554,N_17455);
nor U18397 (N_18397,N_16898,N_17027);
xnor U18398 (N_18398,N_17460,N_17303);
xor U18399 (N_18399,N_17077,N_17267);
and U18400 (N_18400,N_18086,N_17823);
xor U18401 (N_18401,N_18274,N_18043);
nand U18402 (N_18402,N_17670,N_17644);
xor U18403 (N_18403,N_17680,N_18275);
nor U18404 (N_18404,N_18161,N_18369);
nor U18405 (N_18405,N_17972,N_17933);
xor U18406 (N_18406,N_18368,N_18357);
or U18407 (N_18407,N_17960,N_18197);
or U18408 (N_18408,N_17982,N_18067);
nand U18409 (N_18409,N_17978,N_18070);
or U18410 (N_18410,N_17946,N_18032);
or U18411 (N_18411,N_17973,N_18269);
xnor U18412 (N_18412,N_18149,N_18062);
nand U18413 (N_18413,N_17937,N_18088);
and U18414 (N_18414,N_18261,N_17854);
and U18415 (N_18415,N_18291,N_18205);
nor U18416 (N_18416,N_17601,N_17781);
xnor U18417 (N_18417,N_17749,N_17906);
xor U18418 (N_18418,N_17888,N_18359);
nand U18419 (N_18419,N_18074,N_17721);
and U18420 (N_18420,N_17650,N_18083);
xor U18421 (N_18421,N_17782,N_17943);
nand U18422 (N_18422,N_18103,N_18133);
xnor U18423 (N_18423,N_18356,N_18372);
xnor U18424 (N_18424,N_17815,N_18021);
and U18425 (N_18425,N_18000,N_17712);
and U18426 (N_18426,N_18178,N_17754);
nor U18427 (N_18427,N_18039,N_17738);
nor U18428 (N_18428,N_18075,N_18255);
nor U18429 (N_18429,N_17614,N_18335);
xor U18430 (N_18430,N_18251,N_18189);
nand U18431 (N_18431,N_17914,N_17934);
nand U18432 (N_18432,N_18122,N_18293);
and U18433 (N_18433,N_17818,N_18366);
nand U18434 (N_18434,N_17735,N_17967);
or U18435 (N_18435,N_17968,N_18210);
nand U18436 (N_18436,N_17775,N_17811);
xor U18437 (N_18437,N_18303,N_18329);
nor U18438 (N_18438,N_17665,N_18365);
xor U18439 (N_18439,N_18202,N_17727);
or U18440 (N_18440,N_18132,N_18333);
xnor U18441 (N_18441,N_18337,N_18102);
or U18442 (N_18442,N_17926,N_17662);
nand U18443 (N_18443,N_18124,N_18342);
xnor U18444 (N_18444,N_18272,N_18127);
nor U18445 (N_18445,N_17851,N_18037);
xnor U18446 (N_18446,N_17897,N_17828);
nand U18447 (N_18447,N_17750,N_17990);
or U18448 (N_18448,N_17890,N_17959);
nand U18449 (N_18449,N_17718,N_17915);
or U18450 (N_18450,N_18131,N_17814);
and U18451 (N_18451,N_17841,N_17645);
and U18452 (N_18452,N_18284,N_17923);
nor U18453 (N_18453,N_17675,N_17954);
nor U18454 (N_18454,N_18384,N_17808);
nand U18455 (N_18455,N_18173,N_17955);
or U18456 (N_18456,N_17772,N_17704);
nand U18457 (N_18457,N_18136,N_17711);
nor U18458 (N_18458,N_18256,N_17682);
nand U18459 (N_18459,N_17637,N_18171);
nor U18460 (N_18460,N_18388,N_18162);
and U18461 (N_18461,N_18073,N_18362);
or U18462 (N_18462,N_17622,N_17824);
or U18463 (N_18463,N_17974,N_17862);
or U18464 (N_18464,N_18006,N_18024);
or U18465 (N_18465,N_18154,N_17907);
nor U18466 (N_18466,N_18240,N_18081);
xor U18467 (N_18467,N_17669,N_17916);
nand U18468 (N_18468,N_17836,N_18265);
nand U18469 (N_18469,N_18168,N_18228);
or U18470 (N_18470,N_17930,N_17663);
xor U18471 (N_18471,N_17701,N_18207);
xor U18472 (N_18472,N_17667,N_18307);
nor U18473 (N_18473,N_17809,N_17760);
nor U18474 (N_18474,N_17758,N_18018);
nor U18475 (N_18475,N_17941,N_18239);
xor U18476 (N_18476,N_18104,N_18276);
nor U18477 (N_18477,N_17661,N_17668);
xnor U18478 (N_18478,N_17742,N_17776);
nand U18479 (N_18479,N_17688,N_18244);
xor U18480 (N_18480,N_17694,N_17654);
nand U18481 (N_18481,N_18271,N_17684);
and U18482 (N_18482,N_17903,N_17692);
nand U18483 (N_18483,N_18213,N_18302);
nor U18484 (N_18484,N_18097,N_17655);
nand U18485 (N_18485,N_17857,N_17917);
or U18486 (N_18486,N_17633,N_18076);
nor U18487 (N_18487,N_18105,N_17612);
and U18488 (N_18488,N_18186,N_18332);
nor U18489 (N_18489,N_18395,N_17608);
xor U18490 (N_18490,N_18094,N_17947);
and U18491 (N_18491,N_18257,N_17709);
nand U18492 (N_18492,N_18031,N_17865);
nand U18493 (N_18493,N_17904,N_18393);
nor U18494 (N_18494,N_17602,N_18059);
or U18495 (N_18495,N_18108,N_18001);
nor U18496 (N_18496,N_17853,N_18254);
nor U18497 (N_18497,N_17869,N_18199);
and U18498 (N_18498,N_18340,N_17896);
and U18499 (N_18499,N_17696,N_17993);
nor U18500 (N_18500,N_18208,N_18113);
and U18501 (N_18501,N_17698,N_18223);
xor U18502 (N_18502,N_18128,N_18106);
xor U18503 (N_18503,N_18301,N_17658);
xnor U18504 (N_18504,N_18048,N_17646);
and U18505 (N_18505,N_18373,N_18236);
and U18506 (N_18506,N_18014,N_18294);
or U18507 (N_18507,N_18180,N_17998);
or U18508 (N_18508,N_17855,N_18153);
and U18509 (N_18509,N_18306,N_17892);
xor U18510 (N_18510,N_18308,N_17731);
xor U18511 (N_18511,N_18049,N_17653);
and U18512 (N_18512,N_18166,N_18015);
or U18513 (N_18513,N_17970,N_17902);
nand U18514 (N_18514,N_18379,N_18297);
and U18515 (N_18515,N_18025,N_17878);
or U18516 (N_18516,N_18027,N_17879);
or U18517 (N_18517,N_18120,N_17691);
or U18518 (N_18518,N_18175,N_18305);
or U18519 (N_18519,N_17813,N_17605);
xor U18520 (N_18520,N_17844,N_18169);
xor U18521 (N_18521,N_18397,N_17991);
nand U18522 (N_18522,N_18142,N_18188);
nor U18523 (N_18523,N_18320,N_18350);
nand U18524 (N_18524,N_18389,N_18220);
or U18525 (N_18525,N_18182,N_18063);
or U18526 (N_18526,N_18098,N_18065);
or U18527 (N_18527,N_17866,N_17859);
and U18528 (N_18528,N_17631,N_17726);
nand U18529 (N_18529,N_17635,N_18252);
nor U18530 (N_18530,N_17791,N_17801);
nor U18531 (N_18531,N_18242,N_18194);
nand U18532 (N_18532,N_17796,N_17618);
nor U18533 (N_18533,N_18217,N_17604);
nand U18534 (N_18534,N_17626,N_17699);
or U18535 (N_18535,N_18177,N_18058);
or U18536 (N_18536,N_18147,N_17697);
xor U18537 (N_18537,N_18110,N_18211);
xor U18538 (N_18538,N_17804,N_17861);
or U18539 (N_18539,N_17679,N_18262);
and U18540 (N_18540,N_17985,N_17921);
xnor U18541 (N_18541,N_18116,N_17807);
nor U18542 (N_18542,N_18351,N_18247);
and U18543 (N_18543,N_18117,N_18367);
and U18544 (N_18544,N_18078,N_18278);
and U18545 (N_18545,N_18172,N_17621);
or U18546 (N_18546,N_18055,N_17913);
nor U18547 (N_18547,N_17910,N_18341);
and U18548 (N_18548,N_17932,N_18057);
nand U18549 (N_18549,N_17880,N_17900);
nor U18550 (N_18550,N_18030,N_18250);
nor U18551 (N_18551,N_18299,N_18390);
nand U18552 (N_18552,N_17634,N_17950);
and U18553 (N_18553,N_17924,N_18327);
nor U18554 (N_18554,N_18371,N_17838);
nor U18555 (N_18555,N_18158,N_18363);
and U18556 (N_18556,N_18093,N_17827);
and U18557 (N_18557,N_18347,N_17953);
xnor U18558 (N_18558,N_18045,N_18036);
xnor U18559 (N_18559,N_17632,N_17690);
nand U18560 (N_18560,N_18010,N_18259);
or U18561 (N_18561,N_17651,N_17920);
nand U18562 (N_18562,N_17969,N_18016);
nor U18563 (N_18563,N_18085,N_17639);
nand U18564 (N_18564,N_17964,N_17952);
and U18565 (N_18565,N_18192,N_17895);
nor U18566 (N_18566,N_17822,N_18003);
or U18567 (N_18567,N_17929,N_17774);
and U18568 (N_18568,N_18077,N_18007);
or U18569 (N_18569,N_18290,N_17852);
and U18570 (N_18570,N_17683,N_18383);
and U18571 (N_18571,N_18090,N_17871);
or U18572 (N_18572,N_18193,N_17966);
nand U18573 (N_18573,N_17840,N_17716);
nand U18574 (N_18574,N_18135,N_17999);
nor U18575 (N_18575,N_18280,N_17977);
and U18576 (N_18576,N_18052,N_18061);
or U18577 (N_18577,N_17835,N_17961);
nand U18578 (N_18578,N_17842,N_17905);
nand U18579 (N_18579,N_17778,N_17648);
or U18580 (N_18580,N_17764,N_17997);
nand U18581 (N_18581,N_17785,N_18165);
and U18582 (N_18582,N_18398,N_17962);
and U18583 (N_18583,N_18109,N_17886);
and U18584 (N_18584,N_17868,N_18300);
or U18585 (N_18585,N_18391,N_18355);
xor U18586 (N_18586,N_18143,N_17988);
and U18587 (N_18587,N_18319,N_17613);
or U18588 (N_18588,N_17700,N_17723);
and U18589 (N_18589,N_18394,N_17800);
and U18590 (N_18590,N_18241,N_18163);
and U18591 (N_18591,N_17640,N_18151);
or U18592 (N_18592,N_17761,N_17673);
or U18593 (N_18593,N_18339,N_17805);
nor U18594 (N_18594,N_18126,N_17743);
nand U18595 (N_18595,N_17765,N_17752);
nand U18596 (N_18596,N_18164,N_17912);
nor U18597 (N_18597,N_18377,N_17976);
nor U18598 (N_18598,N_18185,N_17714);
nand U18599 (N_18599,N_18328,N_18376);
nand U18600 (N_18600,N_18231,N_17919);
or U18601 (N_18601,N_17705,N_18237);
and U18602 (N_18602,N_18079,N_17734);
nor U18603 (N_18603,N_17736,N_18321);
nor U18604 (N_18604,N_18206,N_18283);
nor U18605 (N_18605,N_17918,N_18227);
and U18606 (N_18606,N_18249,N_17770);
or U18607 (N_18607,N_18386,N_17681);
or U18608 (N_18608,N_17627,N_17739);
nor U18609 (N_18609,N_18222,N_17908);
and U18610 (N_18610,N_17725,N_18204);
or U18611 (N_18611,N_17769,N_17792);
nand U18612 (N_18612,N_18080,N_17837);
nor U18613 (N_18613,N_17607,N_17810);
nand U18614 (N_18614,N_17887,N_18047);
nor U18615 (N_18615,N_18179,N_18101);
xor U18616 (N_18616,N_18196,N_17942);
and U18617 (N_18617,N_18130,N_17717);
or U18618 (N_18618,N_18226,N_18009);
nand U18619 (N_18619,N_18289,N_17816);
xor U18620 (N_18620,N_18100,N_17773);
nand U18621 (N_18621,N_17659,N_18029);
xor U18622 (N_18622,N_18344,N_17703);
nor U18623 (N_18623,N_18349,N_18091);
xnor U18624 (N_18624,N_17883,N_18295);
or U18625 (N_18625,N_17636,N_17802);
and U18626 (N_18626,N_18381,N_17893);
nor U18627 (N_18627,N_17643,N_17821);
or U18628 (N_18628,N_18148,N_18121);
nand U18629 (N_18629,N_17812,N_17931);
xnor U18630 (N_18630,N_18155,N_17945);
xor U18631 (N_18631,N_18345,N_17702);
nand U18632 (N_18632,N_18087,N_18160);
nor U18633 (N_18633,N_18107,N_18174);
nor U18634 (N_18634,N_17877,N_17656);
or U18635 (N_18635,N_18114,N_17984);
nand U18636 (N_18636,N_18243,N_17986);
and U18637 (N_18637,N_18396,N_17641);
nor U18638 (N_18638,N_17677,N_18159);
nor U18639 (N_18639,N_18380,N_18071);
and U18640 (N_18640,N_17676,N_18312);
xor U18641 (N_18641,N_18129,N_17797);
nand U18642 (N_18642,N_17882,N_17664);
xnor U18643 (N_18643,N_18286,N_18035);
or U18644 (N_18644,N_17979,N_18184);
and U18645 (N_18645,N_17720,N_17863);
xor U18646 (N_18646,N_18387,N_17678);
or U18647 (N_18647,N_17831,N_18214);
nor U18648 (N_18648,N_17755,N_18298);
nor U18649 (N_18649,N_18013,N_17820);
nand U18650 (N_18650,N_18044,N_18361);
nor U18651 (N_18651,N_17777,N_18358);
xor U18652 (N_18652,N_17898,N_18137);
nor U18653 (N_18653,N_17759,N_18331);
and U18654 (N_18654,N_18364,N_17671);
nor U18655 (N_18655,N_17944,N_18068);
nand U18656 (N_18656,N_17713,N_18040);
or U18657 (N_18657,N_17995,N_18144);
or U18658 (N_18658,N_17666,N_17687);
nand U18659 (N_18659,N_18092,N_17767);
and U18660 (N_18660,N_17826,N_18285);
nor U18661 (N_18661,N_17845,N_18141);
and U18662 (N_18662,N_18118,N_17956);
nor U18663 (N_18663,N_18183,N_18195);
nand U18664 (N_18664,N_18336,N_17600);
xor U18665 (N_18665,N_17981,N_18370);
nor U18666 (N_18666,N_18156,N_18323);
xnor U18667 (N_18667,N_17695,N_17874);
or U18668 (N_18668,N_17891,N_17829);
or U18669 (N_18669,N_18146,N_18281);
nor U18670 (N_18670,N_18054,N_17722);
and U18671 (N_18671,N_18046,N_17860);
or U18672 (N_18672,N_17783,N_18317);
and U18673 (N_18673,N_18212,N_17751);
nor U18674 (N_18674,N_18082,N_18224);
nor U18675 (N_18675,N_17748,N_17787);
or U18676 (N_18676,N_18176,N_17992);
xnor U18677 (N_18677,N_17948,N_17747);
or U18678 (N_18678,N_18209,N_18002);
and U18679 (N_18679,N_18330,N_18115);
or U18680 (N_18680,N_17935,N_17872);
or U18681 (N_18681,N_18248,N_17963);
nand U18682 (N_18682,N_17615,N_17980);
and U18683 (N_18683,N_17672,N_17839);
or U18684 (N_18684,N_17647,N_18019);
or U18685 (N_18685,N_18041,N_17843);
and U18686 (N_18686,N_17762,N_18221);
or U18687 (N_18687,N_17957,N_18277);
nor U18688 (N_18688,N_18119,N_18038);
nand U18689 (N_18689,N_18215,N_18099);
nand U18690 (N_18690,N_18318,N_18051);
nand U18691 (N_18691,N_18287,N_18198);
or U18692 (N_18692,N_17707,N_17958);
and U18693 (N_18693,N_18399,N_18216);
nand U18694 (N_18694,N_17911,N_18263);
nand U18695 (N_18695,N_17833,N_18382);
nor U18696 (N_18696,N_18053,N_18234);
nand U18697 (N_18697,N_18203,N_18028);
xor U18698 (N_18698,N_17779,N_17889);
or U18699 (N_18699,N_17951,N_18012);
or U18700 (N_18700,N_17850,N_17719);
or U18701 (N_18701,N_17847,N_17885);
xnor U18702 (N_18702,N_17975,N_17971);
xnor U18703 (N_18703,N_17925,N_17740);
xnor U18704 (N_18704,N_17795,N_18279);
or U18705 (N_18705,N_17674,N_17724);
nor U18706 (N_18706,N_18201,N_18020);
and U18707 (N_18707,N_18313,N_17649);
and U18708 (N_18708,N_18112,N_17884);
nand U18709 (N_18709,N_18170,N_18246);
or U18710 (N_18710,N_17628,N_17710);
nand U18711 (N_18711,N_18056,N_17730);
and U18712 (N_18712,N_17803,N_17901);
xor U18713 (N_18713,N_18140,N_17771);
and U18714 (N_18714,N_17638,N_18258);
and U18715 (N_18715,N_18343,N_17728);
and U18716 (N_18716,N_18060,N_17806);
nand U18717 (N_18717,N_17881,N_18334);
nand U18718 (N_18718,N_18392,N_18353);
nor U18719 (N_18719,N_18245,N_17620);
nand U18720 (N_18720,N_17625,N_18253);
nand U18721 (N_18721,N_17819,N_18152);
and U18722 (N_18722,N_17788,N_18023);
xor U18723 (N_18723,N_17642,N_18325);
or U18724 (N_18724,N_18233,N_18123);
and U18725 (N_18725,N_18374,N_17603);
or U18726 (N_18726,N_17623,N_18292);
xnor U18727 (N_18727,N_17753,N_18125);
nand U18728 (N_18728,N_18360,N_18026);
xor U18729 (N_18729,N_18084,N_17825);
xnor U18730 (N_18730,N_18314,N_18311);
nand U18731 (N_18731,N_18266,N_17793);
or U18732 (N_18732,N_17657,N_17830);
or U18733 (N_18733,N_18264,N_17732);
and U18734 (N_18734,N_17799,N_17611);
nor U18735 (N_18735,N_18011,N_17832);
or U18736 (N_18736,N_18230,N_17790);
nor U18737 (N_18737,N_18378,N_17876);
nand U18738 (N_18738,N_17744,N_17909);
or U18739 (N_18739,N_18235,N_18069);
xor U18740 (N_18740,N_18187,N_18096);
nand U18741 (N_18741,N_17846,N_17606);
or U18742 (N_18742,N_17619,N_17817);
nor U18743 (N_18743,N_18326,N_17756);
nor U18744 (N_18744,N_18066,N_18157);
or U18745 (N_18745,N_17927,N_18050);
nand U18746 (N_18746,N_17936,N_18273);
nand U18747 (N_18747,N_18034,N_17780);
xor U18748 (N_18748,N_18095,N_18072);
nor U18749 (N_18749,N_17928,N_18138);
nor U18750 (N_18750,N_18134,N_17987);
or U18751 (N_18751,N_18229,N_17894);
nand U18752 (N_18752,N_18008,N_18346);
and U18753 (N_18753,N_18270,N_17875);
nor U18754 (N_18754,N_18348,N_18005);
or U18755 (N_18755,N_17630,N_17737);
xnor U18756 (N_18756,N_18042,N_18260);
xnor U18757 (N_18757,N_18225,N_18111);
or U18758 (N_18758,N_17685,N_18338);
xor U18759 (N_18759,N_17786,N_17660);
xor U18760 (N_18760,N_18268,N_18200);
nor U18761 (N_18761,N_18167,N_17870);
and U18762 (N_18762,N_18385,N_17849);
nand U18763 (N_18763,N_17864,N_18238);
and U18764 (N_18764,N_17624,N_17938);
nor U18765 (N_18765,N_17746,N_17745);
nand U18766 (N_18766,N_17609,N_18288);
nand U18767 (N_18767,N_18033,N_18352);
xor U18768 (N_18768,N_18324,N_17616);
and U18769 (N_18769,N_18296,N_17922);
nand U18770 (N_18770,N_18139,N_18304);
and U18771 (N_18771,N_17996,N_17939);
nand U18772 (N_18772,N_17789,N_17706);
nor U18773 (N_18773,N_17686,N_17708);
xnor U18774 (N_18774,N_17834,N_18375);
nor U18775 (N_18775,N_17741,N_17858);
or U18776 (N_18776,N_18145,N_18267);
nand U18777 (N_18777,N_17629,N_17766);
xor U18778 (N_18778,N_17733,N_18150);
nor U18779 (N_18779,N_17715,N_17768);
nand U18780 (N_18780,N_17610,N_17784);
or U18781 (N_18781,N_17867,N_18022);
xor U18782 (N_18782,N_18232,N_17983);
and U18783 (N_18783,N_17856,N_17873);
and U18784 (N_18784,N_18004,N_18064);
nand U18785 (N_18785,N_17940,N_18190);
or U18786 (N_18786,N_18218,N_17899);
nand U18787 (N_18787,N_17763,N_18354);
or U18788 (N_18788,N_17729,N_17965);
nand U18789 (N_18789,N_17994,N_18282);
xor U18790 (N_18790,N_18089,N_17757);
or U18791 (N_18791,N_17693,N_17689);
or U18792 (N_18792,N_18315,N_17794);
nor U18793 (N_18793,N_18017,N_18310);
xnor U18794 (N_18794,N_18219,N_18181);
and U18795 (N_18795,N_17652,N_18316);
or U18796 (N_18796,N_18191,N_18322);
xnor U18797 (N_18797,N_17848,N_17798);
nor U18798 (N_18798,N_17989,N_18309);
xor U18799 (N_18799,N_17617,N_17949);
xor U18800 (N_18800,N_17731,N_17834);
nand U18801 (N_18801,N_18113,N_17871);
and U18802 (N_18802,N_18111,N_17720);
nor U18803 (N_18803,N_17919,N_18208);
and U18804 (N_18804,N_18163,N_17740);
or U18805 (N_18805,N_17633,N_18095);
nor U18806 (N_18806,N_18274,N_17884);
and U18807 (N_18807,N_17740,N_17818);
nand U18808 (N_18808,N_18316,N_18241);
nor U18809 (N_18809,N_18027,N_18055);
and U18810 (N_18810,N_18257,N_17772);
nand U18811 (N_18811,N_17849,N_18355);
or U18812 (N_18812,N_17642,N_17729);
xnor U18813 (N_18813,N_17929,N_17700);
or U18814 (N_18814,N_18041,N_18330);
xnor U18815 (N_18815,N_17794,N_17839);
nor U18816 (N_18816,N_17634,N_17603);
nand U18817 (N_18817,N_17797,N_18349);
and U18818 (N_18818,N_17631,N_17771);
nand U18819 (N_18819,N_17679,N_17985);
and U18820 (N_18820,N_17954,N_17687);
nand U18821 (N_18821,N_17965,N_17675);
nor U18822 (N_18822,N_17988,N_18318);
nor U18823 (N_18823,N_18174,N_17824);
or U18824 (N_18824,N_18238,N_17716);
nor U18825 (N_18825,N_18226,N_18309);
nor U18826 (N_18826,N_18261,N_18116);
and U18827 (N_18827,N_17878,N_17710);
or U18828 (N_18828,N_17741,N_17767);
or U18829 (N_18829,N_17693,N_17976);
nand U18830 (N_18830,N_18008,N_18120);
nand U18831 (N_18831,N_17928,N_18275);
xnor U18832 (N_18832,N_18037,N_18307);
xor U18833 (N_18833,N_18164,N_18054);
or U18834 (N_18834,N_17671,N_18174);
nand U18835 (N_18835,N_17636,N_18100);
and U18836 (N_18836,N_18182,N_18317);
nor U18837 (N_18837,N_17903,N_17608);
xnor U18838 (N_18838,N_17854,N_17631);
nand U18839 (N_18839,N_18235,N_18142);
nor U18840 (N_18840,N_17864,N_18222);
nor U18841 (N_18841,N_18340,N_18167);
or U18842 (N_18842,N_18203,N_17856);
nand U18843 (N_18843,N_18270,N_18300);
xnor U18844 (N_18844,N_17658,N_18291);
xnor U18845 (N_18845,N_18209,N_17832);
or U18846 (N_18846,N_18222,N_17724);
nand U18847 (N_18847,N_17977,N_18226);
or U18848 (N_18848,N_18025,N_17728);
xor U18849 (N_18849,N_18314,N_18030);
nor U18850 (N_18850,N_18277,N_18046);
xnor U18851 (N_18851,N_17645,N_18171);
nor U18852 (N_18852,N_18202,N_17983);
or U18853 (N_18853,N_17842,N_17776);
and U18854 (N_18854,N_17874,N_17750);
or U18855 (N_18855,N_18272,N_17891);
nor U18856 (N_18856,N_18105,N_18030);
or U18857 (N_18857,N_17826,N_17792);
or U18858 (N_18858,N_17781,N_18296);
nor U18859 (N_18859,N_17646,N_18210);
nand U18860 (N_18860,N_18215,N_17867);
nor U18861 (N_18861,N_17778,N_17600);
nand U18862 (N_18862,N_17865,N_17778);
or U18863 (N_18863,N_17670,N_18182);
and U18864 (N_18864,N_17957,N_18255);
or U18865 (N_18865,N_17646,N_18127);
nand U18866 (N_18866,N_18247,N_17963);
nand U18867 (N_18867,N_18146,N_17653);
nor U18868 (N_18868,N_18213,N_18148);
and U18869 (N_18869,N_17762,N_18368);
or U18870 (N_18870,N_17691,N_17937);
or U18871 (N_18871,N_17998,N_17700);
nor U18872 (N_18872,N_18356,N_17927);
and U18873 (N_18873,N_18013,N_18025);
nor U18874 (N_18874,N_18219,N_18163);
nor U18875 (N_18875,N_17966,N_17706);
or U18876 (N_18876,N_18206,N_17603);
nand U18877 (N_18877,N_17829,N_17972);
and U18878 (N_18878,N_17877,N_17968);
and U18879 (N_18879,N_17627,N_18173);
or U18880 (N_18880,N_17761,N_17946);
xnor U18881 (N_18881,N_18184,N_17712);
and U18882 (N_18882,N_17676,N_17626);
xor U18883 (N_18883,N_18077,N_18373);
nor U18884 (N_18884,N_18036,N_18165);
or U18885 (N_18885,N_18094,N_17766);
nor U18886 (N_18886,N_18334,N_17756);
nand U18887 (N_18887,N_18105,N_17828);
and U18888 (N_18888,N_18067,N_17791);
xor U18889 (N_18889,N_17986,N_18172);
nand U18890 (N_18890,N_17759,N_18116);
or U18891 (N_18891,N_18264,N_18040);
and U18892 (N_18892,N_17663,N_18344);
nand U18893 (N_18893,N_18105,N_17779);
nand U18894 (N_18894,N_17795,N_18238);
or U18895 (N_18895,N_18049,N_18105);
nor U18896 (N_18896,N_18231,N_17943);
or U18897 (N_18897,N_17970,N_18232);
or U18898 (N_18898,N_17796,N_17812);
nand U18899 (N_18899,N_17979,N_17877);
nand U18900 (N_18900,N_18265,N_18391);
and U18901 (N_18901,N_18129,N_17737);
nand U18902 (N_18902,N_18282,N_17966);
nor U18903 (N_18903,N_17810,N_18242);
and U18904 (N_18904,N_17758,N_17874);
nor U18905 (N_18905,N_17942,N_17750);
nand U18906 (N_18906,N_18112,N_17911);
nand U18907 (N_18907,N_17642,N_18302);
nand U18908 (N_18908,N_17791,N_18000);
xnor U18909 (N_18909,N_18376,N_17972);
or U18910 (N_18910,N_18238,N_17941);
nand U18911 (N_18911,N_17976,N_17704);
or U18912 (N_18912,N_17691,N_17704);
nand U18913 (N_18913,N_18261,N_18136);
nor U18914 (N_18914,N_17993,N_18321);
nand U18915 (N_18915,N_17986,N_17714);
xor U18916 (N_18916,N_18385,N_17700);
and U18917 (N_18917,N_18368,N_18111);
xnor U18918 (N_18918,N_17690,N_17871);
or U18919 (N_18919,N_17899,N_17798);
nor U18920 (N_18920,N_18324,N_18176);
and U18921 (N_18921,N_17944,N_17762);
nand U18922 (N_18922,N_17686,N_17804);
xnor U18923 (N_18923,N_17957,N_17849);
or U18924 (N_18924,N_18273,N_18229);
nor U18925 (N_18925,N_17619,N_17673);
xnor U18926 (N_18926,N_17887,N_18286);
xor U18927 (N_18927,N_17775,N_17667);
and U18928 (N_18928,N_18105,N_17968);
nor U18929 (N_18929,N_18312,N_17836);
and U18930 (N_18930,N_18380,N_17911);
xor U18931 (N_18931,N_17785,N_17792);
nand U18932 (N_18932,N_17867,N_18315);
nor U18933 (N_18933,N_18030,N_18203);
nor U18934 (N_18934,N_17943,N_17621);
xor U18935 (N_18935,N_18135,N_17868);
and U18936 (N_18936,N_17835,N_18277);
or U18937 (N_18937,N_17906,N_17627);
nor U18938 (N_18938,N_18010,N_17779);
nand U18939 (N_18939,N_17831,N_17761);
or U18940 (N_18940,N_17703,N_17916);
and U18941 (N_18941,N_17733,N_18104);
xnor U18942 (N_18942,N_17984,N_17793);
and U18943 (N_18943,N_17838,N_18241);
nand U18944 (N_18944,N_17688,N_18209);
or U18945 (N_18945,N_18174,N_17742);
xor U18946 (N_18946,N_17961,N_18086);
nand U18947 (N_18947,N_18093,N_17982);
or U18948 (N_18948,N_17700,N_17674);
xor U18949 (N_18949,N_17777,N_18055);
and U18950 (N_18950,N_18144,N_17886);
and U18951 (N_18951,N_17774,N_17968);
or U18952 (N_18952,N_17783,N_18152);
or U18953 (N_18953,N_17922,N_18019);
nand U18954 (N_18954,N_17887,N_17603);
nand U18955 (N_18955,N_17779,N_18204);
xor U18956 (N_18956,N_17831,N_18209);
nand U18957 (N_18957,N_17960,N_17746);
or U18958 (N_18958,N_18385,N_17722);
nand U18959 (N_18959,N_18077,N_18289);
nor U18960 (N_18960,N_17880,N_18259);
nor U18961 (N_18961,N_18041,N_18029);
or U18962 (N_18962,N_17671,N_17745);
nand U18963 (N_18963,N_17931,N_18105);
xnor U18964 (N_18964,N_17977,N_18350);
and U18965 (N_18965,N_17957,N_18373);
nor U18966 (N_18966,N_18292,N_18102);
xor U18967 (N_18967,N_18269,N_17860);
xnor U18968 (N_18968,N_18240,N_18143);
nand U18969 (N_18969,N_17691,N_18345);
xnor U18970 (N_18970,N_17705,N_17780);
xnor U18971 (N_18971,N_17620,N_18150);
nand U18972 (N_18972,N_17965,N_18096);
and U18973 (N_18973,N_17728,N_17922);
or U18974 (N_18974,N_17764,N_18057);
or U18975 (N_18975,N_17893,N_18299);
or U18976 (N_18976,N_18200,N_17616);
or U18977 (N_18977,N_18362,N_17978);
and U18978 (N_18978,N_17934,N_17811);
nand U18979 (N_18979,N_17936,N_17633);
nor U18980 (N_18980,N_17987,N_18108);
nand U18981 (N_18981,N_17636,N_17838);
nand U18982 (N_18982,N_18396,N_18006);
nor U18983 (N_18983,N_17653,N_18162);
and U18984 (N_18984,N_17605,N_18093);
and U18985 (N_18985,N_18290,N_17724);
nand U18986 (N_18986,N_17601,N_17946);
xor U18987 (N_18987,N_18193,N_18075);
xor U18988 (N_18988,N_18248,N_17792);
xor U18989 (N_18989,N_17681,N_17777);
xnor U18990 (N_18990,N_18379,N_18243);
nor U18991 (N_18991,N_18113,N_18347);
xnor U18992 (N_18992,N_17758,N_17821);
nand U18993 (N_18993,N_18164,N_18212);
or U18994 (N_18994,N_18332,N_17604);
nand U18995 (N_18995,N_17713,N_17734);
and U18996 (N_18996,N_18087,N_18198);
nor U18997 (N_18997,N_17670,N_18398);
xnor U18998 (N_18998,N_18043,N_18132);
and U18999 (N_18999,N_17865,N_18215);
nor U19000 (N_19000,N_18302,N_17922);
nor U19001 (N_19001,N_18229,N_18014);
or U19002 (N_19002,N_18348,N_18016);
nor U19003 (N_19003,N_18315,N_17994);
nor U19004 (N_19004,N_17642,N_18089);
or U19005 (N_19005,N_17629,N_18142);
xnor U19006 (N_19006,N_17977,N_18396);
nand U19007 (N_19007,N_18189,N_17854);
and U19008 (N_19008,N_18313,N_17901);
nand U19009 (N_19009,N_17713,N_18045);
and U19010 (N_19010,N_18055,N_18106);
nor U19011 (N_19011,N_18089,N_18383);
nand U19012 (N_19012,N_18085,N_18379);
or U19013 (N_19013,N_17893,N_17983);
nand U19014 (N_19014,N_17783,N_18275);
nor U19015 (N_19015,N_17767,N_18248);
xor U19016 (N_19016,N_17654,N_17621);
or U19017 (N_19017,N_17814,N_18196);
nor U19018 (N_19018,N_17759,N_18263);
nor U19019 (N_19019,N_18272,N_17621);
or U19020 (N_19020,N_17760,N_18017);
and U19021 (N_19021,N_18329,N_18382);
or U19022 (N_19022,N_18315,N_17883);
nand U19023 (N_19023,N_18333,N_17715);
xor U19024 (N_19024,N_17876,N_18376);
xor U19025 (N_19025,N_17699,N_18396);
nand U19026 (N_19026,N_18388,N_18348);
nor U19027 (N_19027,N_17697,N_18303);
nand U19028 (N_19028,N_18163,N_18261);
nor U19029 (N_19029,N_17837,N_17825);
nor U19030 (N_19030,N_17960,N_18263);
nand U19031 (N_19031,N_17861,N_18079);
nor U19032 (N_19032,N_18131,N_18132);
xor U19033 (N_19033,N_18392,N_17768);
xnor U19034 (N_19034,N_17885,N_17790);
or U19035 (N_19035,N_18336,N_17898);
and U19036 (N_19036,N_17644,N_18012);
or U19037 (N_19037,N_17790,N_18022);
or U19038 (N_19038,N_17646,N_17783);
or U19039 (N_19039,N_17600,N_18208);
and U19040 (N_19040,N_17653,N_17664);
or U19041 (N_19041,N_18228,N_18381);
xnor U19042 (N_19042,N_18028,N_17853);
xor U19043 (N_19043,N_17900,N_17906);
nand U19044 (N_19044,N_17725,N_17779);
and U19045 (N_19045,N_17645,N_18176);
or U19046 (N_19046,N_18036,N_17985);
or U19047 (N_19047,N_18389,N_18149);
nand U19048 (N_19048,N_18359,N_18096);
nand U19049 (N_19049,N_18356,N_18157);
or U19050 (N_19050,N_17662,N_18275);
nor U19051 (N_19051,N_18368,N_18098);
or U19052 (N_19052,N_18059,N_18215);
xnor U19053 (N_19053,N_18083,N_18080);
nand U19054 (N_19054,N_18074,N_18238);
or U19055 (N_19055,N_17721,N_17628);
xnor U19056 (N_19056,N_18040,N_17974);
or U19057 (N_19057,N_17903,N_18199);
nor U19058 (N_19058,N_18097,N_17993);
nand U19059 (N_19059,N_18048,N_18067);
nand U19060 (N_19060,N_17775,N_17651);
and U19061 (N_19061,N_17703,N_17959);
nand U19062 (N_19062,N_18195,N_18048);
and U19063 (N_19063,N_18001,N_17937);
xnor U19064 (N_19064,N_17925,N_17726);
nor U19065 (N_19065,N_17623,N_17741);
or U19066 (N_19066,N_17784,N_18228);
nand U19067 (N_19067,N_18277,N_17608);
nand U19068 (N_19068,N_18345,N_18121);
nor U19069 (N_19069,N_17684,N_17885);
nor U19070 (N_19070,N_18144,N_18138);
xnor U19071 (N_19071,N_18282,N_17804);
nor U19072 (N_19072,N_18090,N_18271);
nor U19073 (N_19073,N_17885,N_18225);
or U19074 (N_19074,N_17937,N_18153);
nor U19075 (N_19075,N_18022,N_17715);
nand U19076 (N_19076,N_17954,N_17650);
xnor U19077 (N_19077,N_18090,N_17700);
or U19078 (N_19078,N_17833,N_17654);
nor U19079 (N_19079,N_17885,N_17755);
xor U19080 (N_19080,N_17932,N_18228);
or U19081 (N_19081,N_17898,N_17789);
xnor U19082 (N_19082,N_18358,N_18334);
or U19083 (N_19083,N_17671,N_18083);
nor U19084 (N_19084,N_17916,N_18242);
xnor U19085 (N_19085,N_18256,N_17675);
or U19086 (N_19086,N_18223,N_17613);
xor U19087 (N_19087,N_18245,N_17925);
xnor U19088 (N_19088,N_18145,N_18313);
nor U19089 (N_19089,N_18385,N_18370);
nor U19090 (N_19090,N_18200,N_18250);
nand U19091 (N_19091,N_17682,N_18353);
nor U19092 (N_19092,N_17713,N_17683);
nand U19093 (N_19093,N_17943,N_17918);
and U19094 (N_19094,N_17713,N_18220);
xor U19095 (N_19095,N_18062,N_18078);
nand U19096 (N_19096,N_17772,N_17614);
and U19097 (N_19097,N_18225,N_17872);
and U19098 (N_19098,N_18239,N_18328);
xor U19099 (N_19099,N_17661,N_17934);
nand U19100 (N_19100,N_17771,N_18169);
nor U19101 (N_19101,N_18214,N_17661);
nor U19102 (N_19102,N_18160,N_18101);
nor U19103 (N_19103,N_18238,N_17763);
or U19104 (N_19104,N_18053,N_18362);
nor U19105 (N_19105,N_17727,N_18331);
and U19106 (N_19106,N_18345,N_17661);
or U19107 (N_19107,N_18192,N_17600);
and U19108 (N_19108,N_18215,N_18054);
and U19109 (N_19109,N_18148,N_18046);
or U19110 (N_19110,N_17841,N_18306);
nor U19111 (N_19111,N_18295,N_17933);
xor U19112 (N_19112,N_18090,N_17642);
and U19113 (N_19113,N_17968,N_17851);
nor U19114 (N_19114,N_18264,N_17646);
or U19115 (N_19115,N_18368,N_17705);
or U19116 (N_19116,N_18281,N_18094);
nor U19117 (N_19117,N_18073,N_18340);
and U19118 (N_19118,N_17620,N_18100);
nor U19119 (N_19119,N_18161,N_18057);
nand U19120 (N_19120,N_17611,N_18200);
or U19121 (N_19121,N_18362,N_18371);
and U19122 (N_19122,N_17884,N_18154);
xnor U19123 (N_19123,N_18308,N_18145);
or U19124 (N_19124,N_17845,N_18322);
nand U19125 (N_19125,N_18344,N_17649);
xnor U19126 (N_19126,N_17691,N_17618);
and U19127 (N_19127,N_17754,N_18220);
or U19128 (N_19128,N_17895,N_17843);
nand U19129 (N_19129,N_18031,N_17669);
nor U19130 (N_19130,N_17842,N_18273);
xor U19131 (N_19131,N_17698,N_17721);
or U19132 (N_19132,N_18112,N_18005);
xnor U19133 (N_19133,N_18198,N_17636);
xor U19134 (N_19134,N_17906,N_17667);
and U19135 (N_19135,N_17843,N_18123);
nand U19136 (N_19136,N_18077,N_17982);
nand U19137 (N_19137,N_18194,N_17985);
xnor U19138 (N_19138,N_18202,N_17745);
nand U19139 (N_19139,N_17723,N_18380);
or U19140 (N_19140,N_18287,N_17942);
nand U19141 (N_19141,N_18013,N_17947);
or U19142 (N_19142,N_18189,N_17903);
or U19143 (N_19143,N_17797,N_18068);
nor U19144 (N_19144,N_17608,N_18385);
xnor U19145 (N_19145,N_17640,N_17711);
xor U19146 (N_19146,N_18116,N_18145);
and U19147 (N_19147,N_18223,N_17859);
nand U19148 (N_19148,N_17704,N_17747);
or U19149 (N_19149,N_17633,N_17722);
and U19150 (N_19150,N_18305,N_18268);
or U19151 (N_19151,N_18239,N_18254);
xor U19152 (N_19152,N_18236,N_18276);
and U19153 (N_19153,N_18102,N_17720);
xnor U19154 (N_19154,N_17780,N_18285);
or U19155 (N_19155,N_17876,N_18068);
and U19156 (N_19156,N_17890,N_17947);
or U19157 (N_19157,N_18150,N_17859);
and U19158 (N_19158,N_18112,N_17950);
and U19159 (N_19159,N_17819,N_18364);
and U19160 (N_19160,N_18038,N_17759);
and U19161 (N_19161,N_18273,N_17944);
xnor U19162 (N_19162,N_17703,N_18237);
and U19163 (N_19163,N_17700,N_17706);
nand U19164 (N_19164,N_18325,N_17957);
nand U19165 (N_19165,N_18222,N_17666);
or U19166 (N_19166,N_17697,N_18323);
and U19167 (N_19167,N_18364,N_18206);
xnor U19168 (N_19168,N_17748,N_17955);
nand U19169 (N_19169,N_18268,N_18294);
and U19170 (N_19170,N_17655,N_18014);
or U19171 (N_19171,N_17838,N_18267);
nand U19172 (N_19172,N_17860,N_17686);
nand U19173 (N_19173,N_17719,N_17948);
and U19174 (N_19174,N_18238,N_17869);
nand U19175 (N_19175,N_18341,N_18330);
nand U19176 (N_19176,N_17602,N_18190);
nor U19177 (N_19177,N_17816,N_17977);
nand U19178 (N_19178,N_18340,N_18123);
and U19179 (N_19179,N_17941,N_18094);
or U19180 (N_19180,N_17872,N_18310);
xor U19181 (N_19181,N_18114,N_17723);
nor U19182 (N_19182,N_17819,N_18146);
and U19183 (N_19183,N_18267,N_18002);
or U19184 (N_19184,N_18136,N_17790);
or U19185 (N_19185,N_18293,N_17751);
and U19186 (N_19186,N_18154,N_17933);
nand U19187 (N_19187,N_17728,N_18389);
and U19188 (N_19188,N_17830,N_17920);
nor U19189 (N_19189,N_17897,N_17809);
xor U19190 (N_19190,N_18151,N_17887);
nor U19191 (N_19191,N_18256,N_17980);
or U19192 (N_19192,N_17789,N_18206);
xnor U19193 (N_19193,N_17913,N_18111);
nor U19194 (N_19194,N_18348,N_17749);
and U19195 (N_19195,N_17785,N_18170);
or U19196 (N_19196,N_18390,N_18009);
or U19197 (N_19197,N_18207,N_17947);
or U19198 (N_19198,N_18078,N_18142);
and U19199 (N_19199,N_17704,N_17900);
nor U19200 (N_19200,N_18594,N_18601);
or U19201 (N_19201,N_19097,N_18839);
or U19202 (N_19202,N_18935,N_18825);
nand U19203 (N_19203,N_18520,N_18497);
xnor U19204 (N_19204,N_18879,N_19092);
or U19205 (N_19205,N_19091,N_18857);
nand U19206 (N_19206,N_18755,N_19129);
and U19207 (N_19207,N_18807,N_19064);
or U19208 (N_19208,N_19143,N_18609);
or U19209 (N_19209,N_19073,N_18760);
xor U19210 (N_19210,N_18990,N_18424);
or U19211 (N_19211,N_18584,N_18853);
or U19212 (N_19212,N_18618,N_18585);
or U19213 (N_19213,N_18648,N_18923);
or U19214 (N_19214,N_18692,N_18626);
nand U19215 (N_19215,N_18826,N_19106);
nor U19216 (N_19216,N_18819,N_18462);
and U19217 (N_19217,N_18629,N_18421);
nand U19218 (N_19218,N_18414,N_18632);
and U19219 (N_19219,N_18754,N_18565);
and U19220 (N_19220,N_19116,N_19036);
nand U19221 (N_19221,N_18509,N_18737);
nor U19222 (N_19222,N_18578,N_18989);
and U19223 (N_19223,N_18722,N_19068);
or U19224 (N_19224,N_18920,N_18443);
xnor U19225 (N_19225,N_18426,N_19152);
xor U19226 (N_19226,N_18457,N_18590);
xor U19227 (N_19227,N_18720,N_18716);
nand U19228 (N_19228,N_18587,N_18882);
and U19229 (N_19229,N_18476,N_18725);
nand U19230 (N_19230,N_18795,N_19090);
and U19231 (N_19231,N_19004,N_19085);
nor U19232 (N_19232,N_19126,N_18740);
xor U19233 (N_19233,N_18417,N_19155);
xor U19234 (N_19234,N_19055,N_19124);
nor U19235 (N_19235,N_18714,N_19066);
and U19236 (N_19236,N_18663,N_18928);
nor U19237 (N_19237,N_18723,N_18447);
or U19238 (N_19238,N_18786,N_19191);
or U19239 (N_19239,N_18903,N_18436);
and U19240 (N_19240,N_18611,N_18619);
or U19241 (N_19241,N_19083,N_18892);
and U19242 (N_19242,N_18486,N_18652);
nand U19243 (N_19243,N_18470,N_18769);
or U19244 (N_19244,N_18844,N_18772);
or U19245 (N_19245,N_18583,N_19169);
nor U19246 (N_19246,N_18883,N_18501);
xnor U19247 (N_19247,N_18739,N_18442);
or U19248 (N_19248,N_18938,N_19054);
nand U19249 (N_19249,N_19132,N_18773);
nor U19250 (N_19250,N_19110,N_19029);
nand U19251 (N_19251,N_18849,N_19135);
and U19252 (N_19252,N_19179,N_18876);
or U19253 (N_19253,N_18752,N_18451);
xnor U19254 (N_19254,N_18530,N_18402);
nor U19255 (N_19255,N_18809,N_18915);
xnor U19256 (N_19256,N_18834,N_18449);
or U19257 (N_19257,N_18841,N_18662);
nand U19258 (N_19258,N_18728,N_19077);
or U19259 (N_19259,N_19125,N_18867);
xnor U19260 (N_19260,N_18660,N_19052);
xnor U19261 (N_19261,N_18868,N_18713);
or U19262 (N_19262,N_19112,N_18902);
xor U19263 (N_19263,N_18502,N_18899);
or U19264 (N_19264,N_18524,N_18461);
nor U19265 (N_19265,N_18638,N_19161);
xor U19266 (N_19266,N_18790,N_18789);
and U19267 (N_19267,N_18690,N_18753);
nand U19268 (N_19268,N_18535,N_18710);
nand U19269 (N_19269,N_18976,N_18408);
or U19270 (N_19270,N_18680,N_18434);
nor U19271 (N_19271,N_19149,N_18797);
xnor U19272 (N_19272,N_19153,N_18614);
and U19273 (N_19273,N_19021,N_18897);
and U19274 (N_19274,N_19127,N_18569);
nor U19275 (N_19275,N_18644,N_19034);
nand U19276 (N_19276,N_19166,N_18829);
or U19277 (N_19277,N_18922,N_18610);
nand U19278 (N_19278,N_18788,N_19070);
and U19279 (N_19279,N_19115,N_18653);
nand U19280 (N_19280,N_18956,N_18598);
and U19281 (N_19281,N_18541,N_18794);
xnor U19282 (N_19282,N_18507,N_18553);
nand U19283 (N_19283,N_18670,N_18729);
nand U19284 (N_19284,N_18848,N_19067);
xnor U19285 (N_19285,N_18946,N_18767);
and U19286 (N_19286,N_18700,N_19030);
xor U19287 (N_19287,N_18912,N_18743);
xor U19288 (N_19288,N_18908,N_19145);
xnor U19289 (N_19289,N_18593,N_19053);
nand U19290 (N_19290,N_18727,N_18850);
or U19291 (N_19291,N_18861,N_19185);
nand U19292 (N_19292,N_18953,N_18699);
or U19293 (N_19293,N_18961,N_18822);
or U19294 (N_19294,N_18924,N_18955);
xnor U19295 (N_19295,N_19105,N_18950);
or U19296 (N_19296,N_18437,N_18523);
nand U19297 (N_19297,N_18532,N_18419);
or U19298 (N_19298,N_19048,N_18613);
nor U19299 (N_19299,N_19078,N_18589);
nand U19300 (N_19300,N_18639,N_18537);
nand U19301 (N_19301,N_19009,N_19136);
nor U19302 (N_19302,N_18534,N_18745);
xnor U19303 (N_19303,N_18811,N_18905);
xor U19304 (N_19304,N_18561,N_18664);
or U19305 (N_19305,N_19069,N_19050);
or U19306 (N_19306,N_18456,N_18431);
and U19307 (N_19307,N_18941,N_18854);
xor U19308 (N_19308,N_18813,N_18832);
and U19309 (N_19309,N_18872,N_18793);
or U19310 (N_19310,N_18792,N_18758);
xnor U19311 (N_19311,N_18525,N_18642);
and U19312 (N_19312,N_18916,N_19177);
nor U19313 (N_19313,N_18545,N_18816);
nand U19314 (N_19314,N_18407,N_19001);
or U19315 (N_19315,N_18459,N_18776);
and U19316 (N_19316,N_18641,N_18563);
xnor U19317 (N_19317,N_19180,N_18546);
nand U19318 (N_19318,N_18576,N_18891);
xnor U19319 (N_19319,N_18453,N_18901);
or U19320 (N_19320,N_19074,N_18499);
xor U19321 (N_19321,N_18762,N_19003);
and U19322 (N_19322,N_18668,N_18513);
nor U19323 (N_19323,N_19103,N_19075);
xnor U19324 (N_19324,N_18791,N_18873);
xnor U19325 (N_19325,N_19139,N_19170);
and U19326 (N_19326,N_18615,N_18870);
and U19327 (N_19327,N_19163,N_18746);
nor U19328 (N_19328,N_19174,N_18931);
xnor U19329 (N_19329,N_19089,N_18706);
nor U19330 (N_19330,N_19108,N_19111);
or U19331 (N_19331,N_18591,N_18770);
nand U19332 (N_19332,N_18866,N_19164);
nor U19333 (N_19333,N_18688,N_19141);
nand U19334 (N_19334,N_18603,N_18784);
or U19335 (N_19335,N_19150,N_18573);
nand U19336 (N_19336,N_18625,N_18675);
or U19337 (N_19337,N_18798,N_19168);
xnor U19338 (N_19338,N_18577,N_18435);
and U19339 (N_19339,N_18705,N_19013);
nor U19340 (N_19340,N_18588,N_18702);
or U19341 (N_19341,N_19040,N_18712);
and U19342 (N_19342,N_19035,N_19061);
nand U19343 (N_19343,N_18674,N_18572);
nand U19344 (N_19344,N_18778,N_19140);
and U19345 (N_19345,N_19042,N_19080);
and U19346 (N_19346,N_18503,N_18781);
nand U19347 (N_19347,N_18930,N_19015);
or U19348 (N_19348,N_19095,N_19165);
nor U19349 (N_19349,N_18659,N_18815);
and U19350 (N_19350,N_18889,N_18880);
or U19351 (N_19351,N_18810,N_18682);
and U19352 (N_19352,N_18683,N_19008);
xor U19353 (N_19353,N_18708,N_18818);
xnor U19354 (N_19354,N_19192,N_18646);
and U19355 (N_19355,N_18616,N_19197);
and U19356 (N_19356,N_18557,N_19046);
nor U19357 (N_19357,N_18496,N_19184);
or U19358 (N_19358,N_18742,N_18858);
or U19359 (N_19359,N_18914,N_18978);
and U19360 (N_19360,N_19100,N_18721);
nor U19361 (N_19361,N_18544,N_18604);
or U19362 (N_19362,N_19007,N_18697);
nor U19363 (N_19363,N_19117,N_18959);
nor U19364 (N_19364,N_18952,N_18869);
xnor U19365 (N_19365,N_18804,N_18526);
or U19366 (N_19366,N_18846,N_18962);
nand U19367 (N_19367,N_19157,N_18785);
or U19368 (N_19368,N_19199,N_18831);
or U19369 (N_19369,N_18475,N_18988);
or U19370 (N_19370,N_18748,N_19109);
nand U19371 (N_19371,N_18860,N_18987);
and U19372 (N_19372,N_18695,N_18766);
or U19373 (N_19373,N_18726,N_18763);
nand U19374 (N_19374,N_18562,N_18432);
or U19375 (N_19375,N_18884,N_18677);
or U19376 (N_19376,N_18932,N_19119);
or U19377 (N_19377,N_19156,N_19084);
xnor U19378 (N_19378,N_18636,N_18518);
xnor U19379 (N_19379,N_19181,N_18581);
and U19380 (N_19380,N_18717,N_19006);
nor U19381 (N_19381,N_18471,N_18968);
xor U19382 (N_19382,N_19058,N_19183);
xnor U19383 (N_19383,N_18898,N_19138);
and U19384 (N_19384,N_18511,N_19028);
and U19385 (N_19385,N_18489,N_18627);
or U19386 (N_19386,N_18761,N_18970);
nor U19387 (N_19387,N_19059,N_18516);
nor U19388 (N_19388,N_18744,N_18780);
nand U19389 (N_19389,N_19014,N_19167);
and U19390 (N_19390,N_18993,N_18802);
xnor U19391 (N_19391,N_18691,N_18567);
xor U19392 (N_19392,N_19194,N_18528);
xnor U19393 (N_19393,N_18540,N_18881);
and U19394 (N_19394,N_18856,N_19189);
nand U19395 (N_19395,N_19151,N_18894);
xor U19396 (N_19396,N_18775,N_19056);
nand U19397 (N_19397,N_19137,N_18492);
nand U19398 (N_19398,N_18482,N_19107);
nor U19399 (N_19399,N_18508,N_18862);
nand U19400 (N_19400,N_18505,N_18694);
or U19401 (N_19401,N_18582,N_19027);
and U19402 (N_19402,N_18756,N_18676);
or U19403 (N_19403,N_18665,N_18607);
and U19404 (N_19404,N_18689,N_19144);
xor U19405 (N_19405,N_18579,N_19079);
nand U19406 (N_19406,N_18733,N_18983);
nand U19407 (N_19407,N_18494,N_18531);
nor U19408 (N_19408,N_18661,N_19128);
nor U19409 (N_19409,N_18715,N_18425);
and U19410 (N_19410,N_18416,N_19016);
nand U19411 (N_19411,N_19032,N_18801);
xor U19412 (N_19412,N_18647,N_18900);
or U19413 (N_19413,N_18430,N_18568);
nor U19414 (N_19414,N_18735,N_19195);
xnor U19415 (N_19415,N_18612,N_18851);
nand U19416 (N_19416,N_18823,N_19047);
xnor U19417 (N_19417,N_18560,N_18467);
or U19418 (N_19418,N_18672,N_18977);
nor U19419 (N_19419,N_18491,N_18921);
and U19420 (N_19420,N_18599,N_18472);
nor U19421 (N_19421,N_19057,N_18799);
xnor U19422 (N_19422,N_19175,N_18440);
and U19423 (N_19423,N_18515,N_18913);
nand U19424 (N_19424,N_18574,N_18965);
xor U19425 (N_19425,N_18777,N_18498);
xor U19426 (N_19426,N_19099,N_18824);
or U19427 (N_19427,N_18969,N_18877);
or U19428 (N_19428,N_18842,N_18468);
nand U19429 (N_19429,N_18973,N_18975);
or U19430 (N_19430,N_18926,N_18904);
nand U19431 (N_19431,N_18787,N_18687);
nand U19432 (N_19432,N_18982,N_18991);
nand U19433 (N_19433,N_18997,N_18620);
and U19434 (N_19434,N_19019,N_19018);
nor U19435 (N_19435,N_18463,N_18586);
nor U19436 (N_19436,N_18413,N_19041);
and U19437 (N_19437,N_18711,N_19060);
nor U19438 (N_19438,N_18759,N_18566);
or U19439 (N_19439,N_19065,N_18893);
xnor U19440 (N_19440,N_19026,N_19198);
or U19441 (N_19441,N_18685,N_18643);
and U19442 (N_19442,N_18446,N_18992);
nor U19443 (N_19443,N_19037,N_18645);
xnor U19444 (N_19444,N_19002,N_18985);
or U19445 (N_19445,N_18478,N_18655);
nor U19446 (N_19446,N_19159,N_18600);
xor U19447 (N_19447,N_19102,N_18656);
xnor U19448 (N_19448,N_19012,N_18843);
nand U19449 (N_19449,N_18479,N_18465);
xnor U19450 (N_19450,N_18444,N_18731);
nand U19451 (N_19451,N_18483,N_18814);
and U19452 (N_19452,N_19130,N_19134);
nor U19453 (N_19453,N_18657,N_18450);
nor U19454 (N_19454,N_18830,N_18782);
nor U19455 (N_19455,N_18634,N_18596);
or U19456 (N_19456,N_18623,N_18597);
and U19457 (N_19457,N_18986,N_19000);
or U19458 (N_19458,N_18438,N_18765);
or U19459 (N_19459,N_19114,N_19154);
nand U19460 (N_19460,N_18995,N_18847);
and U19461 (N_19461,N_18400,N_18865);
nor U19462 (N_19462,N_19176,N_19096);
xor U19463 (N_19463,N_18556,N_18418);
nand U19464 (N_19464,N_18836,N_18490);
and U19465 (N_19465,N_18917,N_18741);
nor U19466 (N_19466,N_19148,N_19045);
nor U19467 (N_19467,N_19005,N_19082);
xnor U19468 (N_19468,N_18564,N_18747);
or U19469 (N_19469,N_18999,N_18821);
nor U19470 (N_19470,N_18441,N_18484);
and U19471 (N_19471,N_18533,N_18673);
nand U19472 (N_19472,N_18547,N_19121);
xnor U19473 (N_19473,N_18919,N_18863);
or U19474 (N_19474,N_19088,N_18696);
nor U19475 (N_19475,N_18828,N_18718);
xor U19476 (N_19476,N_19044,N_18548);
and U19477 (N_19477,N_19022,N_18666);
or U19478 (N_19478,N_18888,N_18401);
nand U19479 (N_19479,N_18543,N_19011);
nor U19480 (N_19480,N_18979,N_19147);
or U19481 (N_19481,N_18409,N_18940);
or U19482 (N_19482,N_18403,N_18488);
and U19483 (N_19483,N_19173,N_19023);
and U19484 (N_19484,N_18838,N_18466);
and U19485 (N_19485,N_18495,N_18907);
nor U19486 (N_19486,N_18994,N_19188);
or U19487 (N_19487,N_18671,N_18805);
and U19488 (N_19488,N_18605,N_18944);
xnor U19489 (N_19489,N_18684,N_18948);
and U19490 (N_19490,N_19193,N_18833);
and U19491 (N_19491,N_18551,N_18817);
nand U19492 (N_19492,N_19017,N_18529);
nand U19493 (N_19493,N_19087,N_18972);
and U19494 (N_19494,N_18527,N_18939);
xnor U19495 (N_19495,N_18906,N_18649);
xor U19496 (N_19496,N_18945,N_19076);
nand U19497 (N_19497,N_19024,N_18730);
or U19498 (N_19498,N_18942,N_18640);
or U19499 (N_19499,N_18493,N_18933);
nand U19500 (N_19500,N_19093,N_18943);
or U19501 (N_19501,N_19146,N_18559);
or U19502 (N_19502,N_19072,N_18925);
nand U19503 (N_19503,N_19094,N_19039);
nor U19504 (N_19504,N_18783,N_18423);
nand U19505 (N_19505,N_18473,N_18658);
or U19506 (N_19506,N_18521,N_18996);
or U19507 (N_19507,N_18411,N_18885);
xor U19508 (N_19508,N_18448,N_18796);
xnor U19509 (N_19509,N_18764,N_18552);
or U19510 (N_19510,N_18859,N_18410);
and U19511 (N_19511,N_18779,N_18592);
and U19512 (N_19512,N_19081,N_18454);
xnor U19513 (N_19513,N_18927,N_18558);
nor U19514 (N_19514,N_18510,N_18654);
nand U19515 (N_19515,N_18433,N_18678);
nand U19516 (N_19516,N_19172,N_18837);
and U19517 (N_19517,N_18637,N_18420);
nor U19518 (N_19518,N_18845,N_19038);
nor U19519 (N_19519,N_19122,N_18538);
nor U19520 (N_19520,N_19162,N_18422);
nand U19521 (N_19521,N_19118,N_18774);
nor U19522 (N_19522,N_18506,N_19071);
or U19523 (N_19523,N_18957,N_18622);
or U19524 (N_19524,N_18624,N_18840);
or U19525 (N_19525,N_18487,N_18406);
and U19526 (N_19526,N_18517,N_18910);
or U19527 (N_19527,N_18549,N_19120);
or U19528 (N_19528,N_18981,N_18542);
and U19529 (N_19529,N_18911,N_18539);
and U19530 (N_19530,N_18878,N_18669);
or U19531 (N_19531,N_18428,N_18896);
xnor U19532 (N_19532,N_18575,N_18522);
or U19533 (N_19533,N_18724,N_19171);
nor U19534 (N_19534,N_18820,N_18980);
xnor U19535 (N_19535,N_18404,N_19133);
and U19536 (N_19536,N_19033,N_18890);
xnor U19537 (N_19537,N_18936,N_18460);
and U19538 (N_19538,N_18966,N_18963);
nand U19539 (N_19539,N_18806,N_18635);
nor U19540 (N_19540,N_18679,N_18681);
and U19541 (N_19541,N_18949,N_19186);
nor U19542 (N_19542,N_18958,N_18550);
nand U19543 (N_19543,N_18855,N_18909);
or U19544 (N_19544,N_18480,N_18571);
or U19545 (N_19545,N_18427,N_18631);
and U19546 (N_19546,N_18701,N_19101);
and U19547 (N_19547,N_18749,N_19178);
xnor U19548 (N_19548,N_18474,N_18536);
and U19549 (N_19549,N_19010,N_19113);
nor U19550 (N_19550,N_18452,N_18808);
nand U19551 (N_19551,N_18458,N_18469);
or U19552 (N_19552,N_18934,N_18512);
xnor U19553 (N_19553,N_18971,N_18628);
nor U19554 (N_19554,N_18736,N_18595);
nor U19555 (N_19555,N_19104,N_18415);
or U19556 (N_19556,N_19190,N_18703);
nor U19557 (N_19557,N_18709,N_18606);
and U19558 (N_19558,N_19062,N_18738);
nand U19559 (N_19559,N_18998,N_19020);
nor U19560 (N_19560,N_18960,N_18871);
xor U19561 (N_19561,N_19142,N_18602);
or U19562 (N_19562,N_18608,N_18751);
nand U19563 (N_19563,N_19160,N_18750);
xnor U19564 (N_19564,N_19063,N_18617);
nand U19565 (N_19565,N_18918,N_18481);
and U19566 (N_19566,N_19123,N_18554);
or U19567 (N_19567,N_18734,N_18514);
and U19568 (N_19568,N_18947,N_18651);
nor U19569 (N_19569,N_18771,N_18929);
or U19570 (N_19570,N_18800,N_19031);
and U19571 (N_19571,N_18732,N_18964);
and U19572 (N_19572,N_19025,N_18768);
and U19573 (N_19573,N_18698,N_18827);
or U19574 (N_19574,N_18874,N_18650);
nor U19575 (N_19575,N_18429,N_18951);
nor U19576 (N_19576,N_18500,N_18954);
and U19577 (N_19577,N_18519,N_19051);
nand U19578 (N_19578,N_19098,N_19043);
nor U19579 (N_19579,N_18570,N_18803);
or U19580 (N_19580,N_19086,N_18412);
nor U19581 (N_19581,N_18895,N_18937);
nand U19582 (N_19582,N_19187,N_18852);
or U19583 (N_19583,N_18864,N_19158);
and U19584 (N_19584,N_18967,N_18455);
nor U19585 (N_19585,N_18704,N_18633);
xnor U19586 (N_19586,N_18984,N_18812);
nor U19587 (N_19587,N_18405,N_18580);
nor U19588 (N_19588,N_18464,N_18555);
xor U19589 (N_19589,N_18477,N_18667);
or U19590 (N_19590,N_18887,N_18504);
or U19591 (N_19591,N_18439,N_18693);
nor U19592 (N_19592,N_18719,N_18974);
or U19593 (N_19593,N_18707,N_18485);
nor U19594 (N_19594,N_18630,N_18875);
nor U19595 (N_19595,N_19131,N_18886);
and U19596 (N_19596,N_19049,N_18757);
nor U19597 (N_19597,N_18835,N_18445);
or U19598 (N_19598,N_18686,N_19182);
or U19599 (N_19599,N_18621,N_19196);
nand U19600 (N_19600,N_19012,N_18792);
xnor U19601 (N_19601,N_18915,N_18714);
or U19602 (N_19602,N_18669,N_18424);
nor U19603 (N_19603,N_18857,N_18746);
and U19604 (N_19604,N_19162,N_18494);
or U19605 (N_19605,N_18946,N_18917);
nor U19606 (N_19606,N_18999,N_19099);
nand U19607 (N_19607,N_18868,N_19018);
or U19608 (N_19608,N_18897,N_19154);
or U19609 (N_19609,N_18486,N_19137);
nand U19610 (N_19610,N_19157,N_19142);
or U19611 (N_19611,N_18510,N_18584);
xnor U19612 (N_19612,N_18745,N_19191);
and U19613 (N_19613,N_18822,N_18963);
nand U19614 (N_19614,N_18902,N_18668);
and U19615 (N_19615,N_18886,N_18744);
or U19616 (N_19616,N_18966,N_18567);
xor U19617 (N_19617,N_18994,N_18507);
xor U19618 (N_19618,N_18711,N_18543);
nand U19619 (N_19619,N_18811,N_18660);
and U19620 (N_19620,N_18631,N_18480);
nand U19621 (N_19621,N_18600,N_18575);
nor U19622 (N_19622,N_19157,N_18680);
xor U19623 (N_19623,N_19186,N_19195);
and U19624 (N_19624,N_18901,N_19008);
xor U19625 (N_19625,N_18551,N_18478);
and U19626 (N_19626,N_18778,N_18855);
xnor U19627 (N_19627,N_18899,N_19180);
or U19628 (N_19628,N_18477,N_18420);
or U19629 (N_19629,N_19028,N_18548);
or U19630 (N_19630,N_18803,N_18974);
xnor U19631 (N_19631,N_18751,N_19183);
and U19632 (N_19632,N_19156,N_18440);
or U19633 (N_19633,N_19197,N_18423);
and U19634 (N_19634,N_19096,N_19004);
xnor U19635 (N_19635,N_18445,N_18523);
nor U19636 (N_19636,N_19068,N_18511);
xnor U19637 (N_19637,N_18782,N_18925);
or U19638 (N_19638,N_18924,N_18935);
xnor U19639 (N_19639,N_18459,N_19182);
or U19640 (N_19640,N_18556,N_18452);
and U19641 (N_19641,N_18493,N_18714);
nor U19642 (N_19642,N_19088,N_18702);
nand U19643 (N_19643,N_18598,N_19091);
nand U19644 (N_19644,N_18664,N_18834);
or U19645 (N_19645,N_18456,N_19122);
nand U19646 (N_19646,N_18543,N_18908);
or U19647 (N_19647,N_19163,N_18503);
or U19648 (N_19648,N_19035,N_18865);
nand U19649 (N_19649,N_18850,N_18916);
xor U19650 (N_19650,N_19092,N_18563);
or U19651 (N_19651,N_19083,N_18486);
and U19652 (N_19652,N_19158,N_18965);
or U19653 (N_19653,N_19103,N_18994);
nor U19654 (N_19654,N_18943,N_18471);
nor U19655 (N_19655,N_18861,N_18784);
nor U19656 (N_19656,N_19086,N_19079);
xor U19657 (N_19657,N_19128,N_18940);
and U19658 (N_19658,N_19153,N_18888);
and U19659 (N_19659,N_18464,N_18829);
or U19660 (N_19660,N_19065,N_18503);
xor U19661 (N_19661,N_18961,N_18449);
and U19662 (N_19662,N_18999,N_18877);
or U19663 (N_19663,N_19048,N_18913);
and U19664 (N_19664,N_18815,N_18485);
and U19665 (N_19665,N_19019,N_18901);
or U19666 (N_19666,N_19144,N_19163);
xnor U19667 (N_19667,N_18570,N_19119);
nand U19668 (N_19668,N_18676,N_19178);
and U19669 (N_19669,N_19090,N_19150);
or U19670 (N_19670,N_19072,N_18882);
and U19671 (N_19671,N_18729,N_18639);
xor U19672 (N_19672,N_18773,N_18406);
xor U19673 (N_19673,N_18432,N_18434);
nand U19674 (N_19674,N_18942,N_18743);
xnor U19675 (N_19675,N_18911,N_18457);
and U19676 (N_19676,N_18633,N_18750);
and U19677 (N_19677,N_18568,N_18504);
or U19678 (N_19678,N_19165,N_18650);
nand U19679 (N_19679,N_18979,N_18899);
xor U19680 (N_19680,N_18648,N_18538);
or U19681 (N_19681,N_18700,N_18920);
and U19682 (N_19682,N_19069,N_19127);
or U19683 (N_19683,N_19004,N_18975);
nor U19684 (N_19684,N_18857,N_19042);
nor U19685 (N_19685,N_19194,N_18462);
nor U19686 (N_19686,N_18993,N_18895);
nand U19687 (N_19687,N_18489,N_18997);
and U19688 (N_19688,N_18967,N_18958);
or U19689 (N_19689,N_18907,N_18791);
xor U19690 (N_19690,N_18742,N_18992);
and U19691 (N_19691,N_19011,N_18990);
and U19692 (N_19692,N_18527,N_18558);
nor U19693 (N_19693,N_19191,N_18623);
or U19694 (N_19694,N_19018,N_18931);
xnor U19695 (N_19695,N_18441,N_18865);
and U19696 (N_19696,N_18593,N_18963);
xnor U19697 (N_19697,N_18953,N_18542);
nor U19698 (N_19698,N_19122,N_18681);
nor U19699 (N_19699,N_18638,N_19128);
nand U19700 (N_19700,N_18550,N_19198);
nor U19701 (N_19701,N_18602,N_18947);
and U19702 (N_19702,N_18565,N_19064);
and U19703 (N_19703,N_18413,N_18796);
or U19704 (N_19704,N_18420,N_19131);
nand U19705 (N_19705,N_18784,N_18642);
xor U19706 (N_19706,N_18956,N_18632);
and U19707 (N_19707,N_19099,N_18902);
xor U19708 (N_19708,N_18699,N_19180);
xor U19709 (N_19709,N_19196,N_18842);
xor U19710 (N_19710,N_18732,N_18518);
nor U19711 (N_19711,N_18457,N_18420);
xor U19712 (N_19712,N_18863,N_18769);
nor U19713 (N_19713,N_18664,N_18859);
nand U19714 (N_19714,N_19046,N_18440);
nor U19715 (N_19715,N_18407,N_18735);
nand U19716 (N_19716,N_19007,N_18852);
nor U19717 (N_19717,N_18419,N_18514);
and U19718 (N_19718,N_18996,N_18705);
nand U19719 (N_19719,N_18508,N_19073);
xor U19720 (N_19720,N_18476,N_18424);
and U19721 (N_19721,N_18827,N_18655);
xor U19722 (N_19722,N_18804,N_18462);
nand U19723 (N_19723,N_19146,N_18922);
and U19724 (N_19724,N_18692,N_18405);
xor U19725 (N_19725,N_18826,N_18987);
nand U19726 (N_19726,N_18845,N_18959);
nand U19727 (N_19727,N_18462,N_18787);
and U19728 (N_19728,N_18442,N_18777);
nand U19729 (N_19729,N_18870,N_18623);
xor U19730 (N_19730,N_18985,N_18797);
xor U19731 (N_19731,N_18796,N_19035);
and U19732 (N_19732,N_18582,N_19130);
xnor U19733 (N_19733,N_18478,N_18781);
or U19734 (N_19734,N_18777,N_18408);
and U19735 (N_19735,N_18982,N_19193);
or U19736 (N_19736,N_18513,N_18616);
or U19737 (N_19737,N_18809,N_18626);
xnor U19738 (N_19738,N_19044,N_18932);
xor U19739 (N_19739,N_19152,N_18834);
or U19740 (N_19740,N_18777,N_18464);
xnor U19741 (N_19741,N_18742,N_19164);
xor U19742 (N_19742,N_19044,N_19144);
nand U19743 (N_19743,N_18737,N_19092);
nor U19744 (N_19744,N_19137,N_18804);
nand U19745 (N_19745,N_18501,N_18432);
nand U19746 (N_19746,N_18653,N_18722);
and U19747 (N_19747,N_18947,N_19001);
or U19748 (N_19748,N_18710,N_19108);
or U19749 (N_19749,N_18823,N_18501);
nand U19750 (N_19750,N_19100,N_19033);
and U19751 (N_19751,N_18534,N_19133);
nor U19752 (N_19752,N_18467,N_19154);
and U19753 (N_19753,N_19023,N_19120);
xor U19754 (N_19754,N_18833,N_18476);
xor U19755 (N_19755,N_18574,N_19034);
or U19756 (N_19756,N_18943,N_18705);
nor U19757 (N_19757,N_18432,N_18466);
nor U19758 (N_19758,N_19171,N_18734);
xnor U19759 (N_19759,N_19016,N_18454);
or U19760 (N_19760,N_18434,N_18600);
xnor U19761 (N_19761,N_18562,N_19023);
or U19762 (N_19762,N_18403,N_18983);
or U19763 (N_19763,N_18871,N_18722);
or U19764 (N_19764,N_19031,N_18933);
and U19765 (N_19765,N_18797,N_18749);
nand U19766 (N_19766,N_19129,N_19137);
and U19767 (N_19767,N_18774,N_18534);
nor U19768 (N_19768,N_18473,N_18956);
nand U19769 (N_19769,N_18555,N_19193);
or U19770 (N_19770,N_18681,N_19184);
and U19771 (N_19771,N_18819,N_18568);
and U19772 (N_19772,N_19170,N_18474);
or U19773 (N_19773,N_19076,N_19104);
or U19774 (N_19774,N_18451,N_18815);
nor U19775 (N_19775,N_19064,N_18538);
nor U19776 (N_19776,N_18654,N_19173);
nor U19777 (N_19777,N_18700,N_18417);
and U19778 (N_19778,N_18655,N_19035);
and U19779 (N_19779,N_18818,N_18569);
nor U19780 (N_19780,N_18607,N_18634);
xor U19781 (N_19781,N_18528,N_18642);
nand U19782 (N_19782,N_19019,N_18666);
or U19783 (N_19783,N_19185,N_19147);
nand U19784 (N_19784,N_18714,N_18529);
xor U19785 (N_19785,N_18963,N_18820);
or U19786 (N_19786,N_18464,N_18654);
or U19787 (N_19787,N_18733,N_18651);
or U19788 (N_19788,N_19190,N_19064);
and U19789 (N_19789,N_18593,N_18561);
xnor U19790 (N_19790,N_19176,N_18750);
xnor U19791 (N_19791,N_18878,N_18546);
xor U19792 (N_19792,N_19103,N_18615);
nor U19793 (N_19793,N_19081,N_18481);
nand U19794 (N_19794,N_19049,N_18511);
and U19795 (N_19795,N_18619,N_18650);
and U19796 (N_19796,N_18931,N_19117);
and U19797 (N_19797,N_19194,N_18507);
and U19798 (N_19798,N_18666,N_18753);
and U19799 (N_19799,N_18752,N_19067);
nand U19800 (N_19800,N_18903,N_19048);
xnor U19801 (N_19801,N_18463,N_18743);
or U19802 (N_19802,N_18753,N_18577);
xnor U19803 (N_19803,N_18687,N_18959);
nand U19804 (N_19804,N_18806,N_18587);
or U19805 (N_19805,N_19148,N_18971);
or U19806 (N_19806,N_18932,N_18581);
and U19807 (N_19807,N_19035,N_18421);
xor U19808 (N_19808,N_18542,N_18492);
or U19809 (N_19809,N_18845,N_19103);
nand U19810 (N_19810,N_18882,N_18532);
xnor U19811 (N_19811,N_18711,N_18892);
xor U19812 (N_19812,N_18625,N_18421);
nand U19813 (N_19813,N_18627,N_18930);
xor U19814 (N_19814,N_18806,N_18470);
or U19815 (N_19815,N_18568,N_18563);
xor U19816 (N_19816,N_18466,N_18971);
or U19817 (N_19817,N_18602,N_18897);
xnor U19818 (N_19818,N_18550,N_19136);
or U19819 (N_19819,N_19028,N_19088);
and U19820 (N_19820,N_18947,N_18523);
and U19821 (N_19821,N_18739,N_18769);
nand U19822 (N_19822,N_18821,N_18458);
or U19823 (N_19823,N_18768,N_18734);
nand U19824 (N_19824,N_18571,N_18424);
nor U19825 (N_19825,N_18691,N_19098);
or U19826 (N_19826,N_18809,N_18869);
and U19827 (N_19827,N_19177,N_18918);
nand U19828 (N_19828,N_18814,N_19086);
nor U19829 (N_19829,N_18864,N_18832);
and U19830 (N_19830,N_18853,N_18823);
and U19831 (N_19831,N_19043,N_18674);
xor U19832 (N_19832,N_18441,N_18801);
and U19833 (N_19833,N_19039,N_18672);
and U19834 (N_19834,N_18789,N_18480);
nor U19835 (N_19835,N_18630,N_18658);
nor U19836 (N_19836,N_18973,N_18423);
xnor U19837 (N_19837,N_18811,N_18697);
nor U19838 (N_19838,N_18870,N_18453);
xnor U19839 (N_19839,N_18652,N_18519);
nor U19840 (N_19840,N_18807,N_18813);
or U19841 (N_19841,N_18746,N_18506);
nor U19842 (N_19842,N_18409,N_18959);
nor U19843 (N_19843,N_19096,N_18665);
xor U19844 (N_19844,N_19083,N_18765);
nand U19845 (N_19845,N_18835,N_18751);
and U19846 (N_19846,N_18992,N_19016);
and U19847 (N_19847,N_18515,N_19037);
or U19848 (N_19848,N_18481,N_18759);
nand U19849 (N_19849,N_19149,N_18969);
or U19850 (N_19850,N_18478,N_18839);
nand U19851 (N_19851,N_19166,N_19140);
nand U19852 (N_19852,N_18427,N_18589);
or U19853 (N_19853,N_18484,N_18964);
nor U19854 (N_19854,N_18606,N_18736);
xor U19855 (N_19855,N_19098,N_18508);
nand U19856 (N_19856,N_18981,N_18829);
or U19857 (N_19857,N_18443,N_18863);
and U19858 (N_19858,N_18471,N_18421);
or U19859 (N_19859,N_18773,N_18873);
nand U19860 (N_19860,N_18525,N_18847);
and U19861 (N_19861,N_18747,N_18629);
and U19862 (N_19862,N_18707,N_19125);
or U19863 (N_19863,N_19183,N_18667);
and U19864 (N_19864,N_18718,N_19016);
and U19865 (N_19865,N_19145,N_18621);
nand U19866 (N_19866,N_19076,N_18896);
xnor U19867 (N_19867,N_18578,N_19019);
xnor U19868 (N_19868,N_19196,N_18777);
xnor U19869 (N_19869,N_18449,N_18947);
xnor U19870 (N_19870,N_18505,N_18651);
and U19871 (N_19871,N_19106,N_18775);
xor U19872 (N_19872,N_19007,N_18872);
nand U19873 (N_19873,N_18892,N_18588);
or U19874 (N_19874,N_18785,N_18524);
and U19875 (N_19875,N_18755,N_18846);
and U19876 (N_19876,N_19015,N_19030);
and U19877 (N_19877,N_18859,N_19116);
nor U19878 (N_19878,N_18728,N_18961);
or U19879 (N_19879,N_18961,N_18899);
or U19880 (N_19880,N_18928,N_18960);
nand U19881 (N_19881,N_18707,N_18843);
nor U19882 (N_19882,N_19058,N_18516);
or U19883 (N_19883,N_18609,N_18881);
or U19884 (N_19884,N_19142,N_18425);
nor U19885 (N_19885,N_18545,N_18940);
nand U19886 (N_19886,N_18444,N_18576);
and U19887 (N_19887,N_18714,N_18903);
and U19888 (N_19888,N_18874,N_18450);
and U19889 (N_19889,N_18594,N_18795);
and U19890 (N_19890,N_18967,N_18848);
nand U19891 (N_19891,N_18492,N_19111);
nand U19892 (N_19892,N_19146,N_18461);
xnor U19893 (N_19893,N_18458,N_18714);
or U19894 (N_19894,N_18524,N_19044);
and U19895 (N_19895,N_19024,N_18624);
xnor U19896 (N_19896,N_18531,N_19147);
nand U19897 (N_19897,N_18627,N_18538);
nand U19898 (N_19898,N_18498,N_18832);
or U19899 (N_19899,N_18566,N_18860);
and U19900 (N_19900,N_18510,N_18848);
nand U19901 (N_19901,N_18736,N_18964);
nand U19902 (N_19902,N_18737,N_19008);
nor U19903 (N_19903,N_19075,N_18602);
and U19904 (N_19904,N_18890,N_19003);
nor U19905 (N_19905,N_18653,N_18774);
nor U19906 (N_19906,N_18495,N_19072);
and U19907 (N_19907,N_18791,N_18976);
or U19908 (N_19908,N_18990,N_18885);
nor U19909 (N_19909,N_18401,N_18575);
and U19910 (N_19910,N_18906,N_19075);
nand U19911 (N_19911,N_18593,N_18749);
xnor U19912 (N_19912,N_19007,N_19022);
nor U19913 (N_19913,N_18577,N_18442);
xor U19914 (N_19914,N_18818,N_18835);
or U19915 (N_19915,N_19059,N_18745);
nand U19916 (N_19916,N_19100,N_19131);
nand U19917 (N_19917,N_18476,N_19088);
xor U19918 (N_19918,N_18907,N_18951);
and U19919 (N_19919,N_18533,N_18843);
nand U19920 (N_19920,N_18451,N_18404);
or U19921 (N_19921,N_18706,N_18650);
nand U19922 (N_19922,N_18906,N_18643);
xor U19923 (N_19923,N_19163,N_19019);
and U19924 (N_19924,N_18585,N_19148);
xnor U19925 (N_19925,N_18676,N_18850);
nand U19926 (N_19926,N_18888,N_18876);
or U19927 (N_19927,N_19127,N_18805);
nor U19928 (N_19928,N_18566,N_18869);
and U19929 (N_19929,N_18620,N_19147);
nand U19930 (N_19930,N_18584,N_18756);
or U19931 (N_19931,N_18932,N_19011);
nand U19932 (N_19932,N_18760,N_18574);
xnor U19933 (N_19933,N_18931,N_19185);
nor U19934 (N_19934,N_18830,N_18547);
nor U19935 (N_19935,N_18595,N_18891);
nor U19936 (N_19936,N_18513,N_18874);
xnor U19937 (N_19937,N_18539,N_18693);
and U19938 (N_19938,N_18412,N_19069);
or U19939 (N_19939,N_18823,N_18807);
xnor U19940 (N_19940,N_18462,N_18760);
xor U19941 (N_19941,N_18783,N_18734);
xnor U19942 (N_19942,N_18530,N_18625);
nand U19943 (N_19943,N_18938,N_19030);
xnor U19944 (N_19944,N_18869,N_19193);
xor U19945 (N_19945,N_18825,N_19170);
xor U19946 (N_19946,N_18792,N_18644);
and U19947 (N_19947,N_18833,N_19186);
xnor U19948 (N_19948,N_18796,N_19057);
and U19949 (N_19949,N_18620,N_19010);
nand U19950 (N_19950,N_18917,N_19076);
or U19951 (N_19951,N_18550,N_19013);
nand U19952 (N_19952,N_19183,N_18725);
or U19953 (N_19953,N_18525,N_19116);
xnor U19954 (N_19954,N_18929,N_18974);
xnor U19955 (N_19955,N_18510,N_18650);
nor U19956 (N_19956,N_18979,N_19018);
and U19957 (N_19957,N_18494,N_18658);
nand U19958 (N_19958,N_19181,N_18436);
nor U19959 (N_19959,N_18407,N_18853);
and U19960 (N_19960,N_18492,N_18640);
xor U19961 (N_19961,N_18741,N_19079);
or U19962 (N_19962,N_18704,N_18985);
xnor U19963 (N_19963,N_18956,N_18677);
nor U19964 (N_19964,N_18992,N_18652);
nor U19965 (N_19965,N_18750,N_18588);
xnor U19966 (N_19966,N_18855,N_18930);
and U19967 (N_19967,N_19157,N_18489);
xor U19968 (N_19968,N_18463,N_19160);
and U19969 (N_19969,N_18941,N_18424);
nor U19970 (N_19970,N_19066,N_18961);
or U19971 (N_19971,N_18845,N_19154);
or U19972 (N_19972,N_19079,N_18711);
or U19973 (N_19973,N_19114,N_18411);
and U19974 (N_19974,N_18805,N_18807);
or U19975 (N_19975,N_18973,N_18565);
xnor U19976 (N_19976,N_18765,N_18636);
or U19977 (N_19977,N_19111,N_18611);
or U19978 (N_19978,N_18510,N_18628);
nor U19979 (N_19979,N_18455,N_18676);
and U19980 (N_19980,N_18442,N_18718);
and U19981 (N_19981,N_18750,N_19167);
or U19982 (N_19982,N_18536,N_19161);
xor U19983 (N_19983,N_18638,N_19094);
and U19984 (N_19984,N_18998,N_18668);
nor U19985 (N_19985,N_18972,N_19049);
and U19986 (N_19986,N_18466,N_18950);
nand U19987 (N_19987,N_18599,N_19191);
xnor U19988 (N_19988,N_19087,N_18883);
xor U19989 (N_19989,N_18782,N_19191);
xnor U19990 (N_19990,N_18858,N_18642);
and U19991 (N_19991,N_18671,N_18626);
and U19992 (N_19992,N_18744,N_18558);
or U19993 (N_19993,N_18874,N_18721);
nor U19994 (N_19994,N_18657,N_18609);
nor U19995 (N_19995,N_18736,N_19158);
or U19996 (N_19996,N_19129,N_18707);
and U19997 (N_19997,N_18896,N_18585);
xnor U19998 (N_19998,N_18806,N_19018);
nor U19999 (N_19999,N_18554,N_18643);
nand UO_0 (O_0,N_19228,N_19525);
nor UO_1 (O_1,N_19892,N_19596);
nand UO_2 (O_2,N_19867,N_19311);
nand UO_3 (O_3,N_19509,N_19550);
nand UO_4 (O_4,N_19471,N_19413);
or UO_5 (O_5,N_19869,N_19487);
xnor UO_6 (O_6,N_19896,N_19830);
nor UO_7 (O_7,N_19322,N_19443);
xor UO_8 (O_8,N_19782,N_19607);
nor UO_9 (O_9,N_19784,N_19383);
nand UO_10 (O_10,N_19408,N_19964);
nor UO_11 (O_11,N_19420,N_19912);
nand UO_12 (O_12,N_19865,N_19366);
xnor UO_13 (O_13,N_19367,N_19635);
xnor UO_14 (O_14,N_19465,N_19579);
nand UO_15 (O_15,N_19794,N_19988);
or UO_16 (O_16,N_19209,N_19762);
or UO_17 (O_17,N_19280,N_19642);
and UO_18 (O_18,N_19645,N_19445);
nand UO_19 (O_19,N_19557,N_19499);
or UO_20 (O_20,N_19619,N_19270);
nand UO_21 (O_21,N_19974,N_19944);
or UO_22 (O_22,N_19205,N_19775);
nand UO_23 (O_23,N_19336,N_19301);
and UO_24 (O_24,N_19754,N_19340);
nand UO_25 (O_25,N_19513,N_19318);
or UO_26 (O_26,N_19661,N_19781);
nand UO_27 (O_27,N_19751,N_19600);
nand UO_28 (O_28,N_19660,N_19750);
nor UO_29 (O_29,N_19686,N_19658);
or UO_30 (O_30,N_19657,N_19516);
xnor UO_31 (O_31,N_19728,N_19272);
or UO_32 (O_32,N_19877,N_19970);
nor UO_33 (O_33,N_19588,N_19310);
nor UO_34 (O_34,N_19584,N_19925);
or UO_35 (O_35,N_19883,N_19552);
or UO_36 (O_36,N_19558,N_19911);
xnor UO_37 (O_37,N_19479,N_19456);
nor UO_38 (O_38,N_19563,N_19293);
and UO_39 (O_39,N_19214,N_19822);
and UO_40 (O_40,N_19341,N_19795);
xnor UO_41 (O_41,N_19387,N_19868);
nor UO_42 (O_42,N_19723,N_19705);
and UO_43 (O_43,N_19326,N_19717);
nand UO_44 (O_44,N_19647,N_19519);
nand UO_45 (O_45,N_19609,N_19874);
nor UO_46 (O_46,N_19587,N_19601);
or UO_47 (O_47,N_19483,N_19960);
nor UO_48 (O_48,N_19540,N_19440);
nor UO_49 (O_49,N_19947,N_19521);
nand UO_50 (O_50,N_19790,N_19282);
xnor UO_51 (O_51,N_19767,N_19941);
nor UO_52 (O_52,N_19783,N_19304);
or UO_53 (O_53,N_19757,N_19298);
nand UO_54 (O_54,N_19539,N_19332);
or UO_55 (O_55,N_19543,N_19756);
nand UO_56 (O_56,N_19325,N_19360);
nor UO_57 (O_57,N_19294,N_19888);
and UO_58 (O_58,N_19247,N_19889);
nor UO_59 (O_59,N_19855,N_19991);
and UO_60 (O_60,N_19396,N_19204);
and UO_61 (O_61,N_19417,N_19859);
and UO_62 (O_62,N_19863,N_19286);
and UO_63 (O_63,N_19873,N_19504);
or UO_64 (O_64,N_19410,N_19449);
or UO_65 (O_65,N_19772,N_19544);
xor UO_66 (O_66,N_19371,N_19350);
xnor UO_67 (O_67,N_19671,N_19624);
nand UO_68 (O_68,N_19524,N_19740);
xor UO_69 (O_69,N_19996,N_19844);
and UO_70 (O_70,N_19778,N_19501);
or UO_71 (O_71,N_19345,N_19429);
xor UO_72 (O_72,N_19560,N_19886);
nand UO_73 (O_73,N_19743,N_19320);
xor UO_74 (O_74,N_19989,N_19983);
and UO_75 (O_75,N_19779,N_19735);
or UO_76 (O_76,N_19695,N_19853);
and UO_77 (O_77,N_19585,N_19678);
or UO_78 (O_78,N_19771,N_19526);
xnor UO_79 (O_79,N_19799,N_19528);
and UO_80 (O_80,N_19264,N_19680);
xor UO_81 (O_81,N_19724,N_19399);
nor UO_82 (O_82,N_19871,N_19495);
or UO_83 (O_83,N_19901,N_19463);
nor UO_84 (O_84,N_19916,N_19712);
or UO_85 (O_85,N_19802,N_19218);
xor UO_86 (O_86,N_19927,N_19358);
and UO_87 (O_87,N_19200,N_19651);
or UO_88 (O_88,N_19774,N_19237);
xor UO_89 (O_89,N_19469,N_19250);
nand UO_90 (O_90,N_19694,N_19577);
nand UO_91 (O_91,N_19667,N_19404);
nor UO_92 (O_92,N_19634,N_19826);
or UO_93 (O_93,N_19485,N_19663);
nand UO_94 (O_94,N_19720,N_19477);
xor UO_95 (O_95,N_19679,N_19491);
or UO_96 (O_96,N_19818,N_19226);
or UO_97 (O_97,N_19673,N_19805);
and UO_98 (O_98,N_19520,N_19628);
nor UO_99 (O_99,N_19356,N_19212);
nor UO_100 (O_100,N_19776,N_19913);
xnor UO_101 (O_101,N_19536,N_19255);
nand UO_102 (O_102,N_19254,N_19407);
or UO_103 (O_103,N_19419,N_19581);
nor UO_104 (O_104,N_19820,N_19578);
xnor UO_105 (O_105,N_19765,N_19347);
or UO_106 (O_106,N_19738,N_19953);
xor UO_107 (O_107,N_19403,N_19241);
xnor UO_108 (O_108,N_19676,N_19530);
nor UO_109 (O_109,N_19814,N_19801);
nand UO_110 (O_110,N_19849,N_19342);
xor UO_111 (O_111,N_19299,N_19380);
xor UO_112 (O_112,N_19880,N_19458);
and UO_113 (O_113,N_19936,N_19637);
or UO_114 (O_114,N_19897,N_19636);
nand UO_115 (O_115,N_19986,N_19269);
or UO_116 (O_116,N_19426,N_19923);
xnor UO_117 (O_117,N_19773,N_19887);
and UO_118 (O_118,N_19608,N_19289);
nand UO_119 (O_119,N_19278,N_19405);
nor UO_120 (O_120,N_19786,N_19502);
xor UO_121 (O_121,N_19593,N_19732);
or UO_122 (O_122,N_19955,N_19571);
nor UO_123 (O_123,N_19677,N_19210);
xor UO_124 (O_124,N_19514,N_19486);
nor UO_125 (O_125,N_19351,N_19933);
xnor UO_126 (O_126,N_19703,N_19438);
nand UO_127 (O_127,N_19261,N_19850);
or UO_128 (O_128,N_19731,N_19721);
nor UO_129 (O_129,N_19696,N_19373);
nor UO_130 (O_130,N_19249,N_19576);
or UO_131 (O_131,N_19534,N_19494);
nand UO_132 (O_132,N_19812,N_19498);
nand UO_133 (O_133,N_19496,N_19545);
xnor UO_134 (O_134,N_19851,N_19630);
xnor UO_135 (O_135,N_19856,N_19924);
or UO_136 (O_136,N_19234,N_19872);
nor UO_137 (O_137,N_19833,N_19353);
xor UO_138 (O_138,N_19309,N_19674);
xnor UO_139 (O_139,N_19616,N_19908);
nor UO_140 (O_140,N_19764,N_19281);
nand UO_141 (O_141,N_19948,N_19837);
and UO_142 (O_142,N_19659,N_19905);
nand UO_143 (O_143,N_19727,N_19461);
or UO_144 (O_144,N_19468,N_19422);
nand UO_145 (O_145,N_19506,N_19357);
and UO_146 (O_146,N_19453,N_19533);
nor UO_147 (O_147,N_19719,N_19981);
or UO_148 (O_148,N_19917,N_19315);
nor UO_149 (O_149,N_19308,N_19839);
and UO_150 (O_150,N_19497,N_19233);
xnor UO_151 (O_151,N_19243,N_19537);
or UO_152 (O_152,N_19825,N_19484);
and UO_153 (O_153,N_19423,N_19388);
xnor UO_154 (O_154,N_19610,N_19971);
nand UO_155 (O_155,N_19303,N_19758);
xor UO_156 (O_156,N_19527,N_19605);
and UO_157 (O_157,N_19736,N_19492);
nand UO_158 (O_158,N_19231,N_19523);
nand UO_159 (O_159,N_19878,N_19565);
nor UO_160 (O_160,N_19421,N_19207);
and UO_161 (O_161,N_19554,N_19796);
nor UO_162 (O_162,N_19666,N_19392);
nand UO_163 (O_163,N_19531,N_19699);
nor UO_164 (O_164,N_19515,N_19920);
xor UO_165 (O_165,N_19361,N_19391);
nor UO_166 (O_166,N_19760,N_19306);
xnor UO_167 (O_167,N_19507,N_19295);
or UO_168 (O_168,N_19283,N_19427);
and UO_169 (O_169,N_19276,N_19447);
nor UO_170 (O_170,N_19561,N_19314);
nand UO_171 (O_171,N_19646,N_19446);
and UO_172 (O_172,N_19797,N_19791);
nor UO_173 (O_173,N_19393,N_19572);
and UO_174 (O_174,N_19542,N_19535);
nor UO_175 (O_175,N_19442,N_19595);
or UO_176 (O_176,N_19745,N_19586);
nor UO_177 (O_177,N_19846,N_19599);
nand UO_178 (O_178,N_19291,N_19631);
or UO_179 (O_179,N_19945,N_19473);
or UO_180 (O_180,N_19662,N_19928);
nor UO_181 (O_181,N_19547,N_19777);
nand UO_182 (O_182,N_19838,N_19653);
and UO_183 (O_183,N_19211,N_19302);
or UO_184 (O_184,N_19379,N_19954);
nor UO_185 (O_185,N_19275,N_19604);
and UO_186 (O_186,N_19994,N_19847);
and UO_187 (O_187,N_19843,N_19223);
xor UO_188 (O_188,N_19919,N_19359);
nor UO_189 (O_189,N_19733,N_19685);
or UO_190 (O_190,N_19215,N_19329);
nand UO_191 (O_191,N_19459,N_19553);
or UO_192 (O_192,N_19323,N_19793);
or UO_193 (O_193,N_19397,N_19489);
nand UO_194 (O_194,N_19956,N_19297);
xnor UO_195 (O_195,N_19979,N_19242);
nor UO_196 (O_196,N_19821,N_19382);
nand UO_197 (O_197,N_19759,N_19993);
xnor UO_198 (O_198,N_19984,N_19934);
or UO_199 (O_199,N_19222,N_19747);
nor UO_200 (O_200,N_19603,N_19374);
nor UO_201 (O_201,N_19997,N_19834);
xnor UO_202 (O_202,N_19963,N_19655);
xnor UO_203 (O_203,N_19879,N_19672);
nor UO_204 (O_204,N_19618,N_19448);
or UO_205 (O_205,N_19355,N_19292);
xor UO_206 (O_206,N_19225,N_19935);
nor UO_207 (O_207,N_19706,N_19615);
nor UO_208 (O_208,N_19472,N_19606);
or UO_209 (O_209,N_19835,N_19707);
nand UO_210 (O_210,N_19462,N_19556);
nor UO_211 (O_211,N_19395,N_19832);
nor UO_212 (O_212,N_19348,N_19860);
and UO_213 (O_213,N_19726,N_19766);
or UO_214 (O_214,N_19288,N_19650);
nor UO_215 (O_215,N_19918,N_19828);
nand UO_216 (O_216,N_19335,N_19900);
and UO_217 (O_217,N_19914,N_19962);
nand UO_218 (O_218,N_19389,N_19381);
or UO_219 (O_219,N_19433,N_19296);
or UO_220 (O_220,N_19891,N_19598);
and UO_221 (O_221,N_19253,N_19493);
or UO_222 (O_222,N_19475,N_19803);
or UO_223 (O_223,N_19575,N_19780);
nor UO_224 (O_224,N_19273,N_19592);
nand UO_225 (O_225,N_19546,N_19852);
xor UO_226 (O_226,N_19375,N_19248);
and UO_227 (O_227,N_19246,N_19614);
nor UO_228 (O_228,N_19861,N_19890);
or UO_229 (O_229,N_19952,N_19836);
and UO_230 (O_230,N_19922,N_19701);
nand UO_231 (O_231,N_19252,N_19641);
nor UO_232 (O_232,N_19875,N_19319);
xor UO_233 (O_233,N_19439,N_19627);
nor UO_234 (O_234,N_19260,N_19508);
and UO_235 (O_235,N_19338,N_19415);
and UO_236 (O_236,N_19700,N_19206);
and UO_237 (O_237,N_19398,N_19966);
or UO_238 (O_238,N_19684,N_19203);
nand UO_239 (O_239,N_19245,N_19969);
nand UO_240 (O_240,N_19792,N_19620);
nand UO_241 (O_241,N_19416,N_19798);
nor UO_242 (O_242,N_19227,N_19364);
or UO_243 (O_243,N_19734,N_19749);
nor UO_244 (O_244,N_19467,N_19470);
nor UO_245 (O_245,N_19744,N_19845);
and UO_246 (O_246,N_19590,N_19510);
xnor UO_247 (O_247,N_19815,N_19999);
nor UO_248 (O_248,N_19414,N_19321);
and UO_249 (O_249,N_19580,N_19394);
nor UO_250 (O_250,N_19939,N_19343);
xor UO_251 (O_251,N_19808,N_19800);
or UO_252 (O_252,N_19406,N_19597);
and UO_253 (O_253,N_19946,N_19995);
xnor UO_254 (O_254,N_19482,N_19229);
nand UO_255 (O_255,N_19625,N_19428);
xnor UO_256 (O_256,N_19682,N_19817);
nand UO_257 (O_257,N_19583,N_19788);
nor UO_258 (O_258,N_19266,N_19412);
or UO_259 (O_259,N_19307,N_19804);
or UO_260 (O_260,N_19591,N_19431);
and UO_261 (O_261,N_19327,N_19372);
or UO_262 (O_262,N_19626,N_19702);
and UO_263 (O_263,N_19787,N_19377);
or UO_264 (O_264,N_19967,N_19538);
nor UO_265 (O_265,N_19259,N_19907);
or UO_266 (O_266,N_19904,N_19263);
nor UO_267 (O_267,N_19725,N_19555);
xor UO_268 (O_268,N_19882,N_19384);
nand UO_269 (O_269,N_19457,N_19434);
or UO_270 (O_270,N_19612,N_19741);
or UO_271 (O_271,N_19769,N_19938);
and UO_272 (O_272,N_19737,N_19568);
or UO_273 (O_273,N_19349,N_19648);
and UO_274 (O_274,N_19687,N_19770);
nand UO_275 (O_275,N_19268,N_19668);
xor UO_276 (O_276,N_19220,N_19236);
nor UO_277 (O_277,N_19279,N_19257);
and UO_278 (O_278,N_19567,N_19602);
nand UO_279 (O_279,N_19213,N_19709);
xnor UO_280 (O_280,N_19208,N_19884);
and UO_281 (O_281,N_19354,N_19858);
nor UO_282 (O_282,N_19722,N_19277);
and UO_283 (O_283,N_19569,N_19240);
xor UO_284 (O_284,N_19930,N_19730);
xor UO_285 (O_285,N_19481,N_19511);
or UO_286 (O_286,N_19235,N_19566);
xor UO_287 (O_287,N_19573,N_19441);
and UO_288 (O_288,N_19866,N_19224);
or UO_289 (O_289,N_19450,N_19337);
nor UO_290 (O_290,N_19386,N_19763);
or UO_291 (O_291,N_19681,N_19937);
nor UO_292 (O_292,N_19632,N_19940);
or UO_293 (O_293,N_19895,N_19665);
nand UO_294 (O_294,N_19430,N_19339);
nand UO_295 (O_295,N_19957,N_19488);
nor UO_296 (O_296,N_19522,N_19312);
nand UO_297 (O_297,N_19840,N_19638);
nor UO_298 (O_298,N_19400,N_19857);
xnor UO_299 (O_299,N_19714,N_19718);
and UO_300 (O_300,N_19819,N_19894);
or UO_301 (O_301,N_19965,N_19987);
and UO_302 (O_302,N_19480,N_19490);
nor UO_303 (O_303,N_19972,N_19915);
or UO_304 (O_304,N_19689,N_19369);
xor UO_305 (O_305,N_19958,N_19378);
or UO_306 (O_306,N_19451,N_19929);
nor UO_307 (O_307,N_19401,N_19752);
nand UO_308 (O_308,N_19985,N_19729);
or UO_309 (O_309,N_19761,N_19902);
and UO_310 (O_310,N_19432,N_19824);
or UO_311 (O_311,N_19324,N_19809);
nor UO_312 (O_312,N_19711,N_19697);
nand UO_313 (O_313,N_19640,N_19316);
and UO_314 (O_314,N_19466,N_19633);
nand UO_315 (O_315,N_19217,N_19742);
nand UO_316 (O_316,N_19644,N_19346);
or UO_317 (O_317,N_19444,N_19334);
xor UO_318 (O_318,N_19256,N_19518);
xor UO_319 (O_319,N_19950,N_19232);
nand UO_320 (O_320,N_19436,N_19500);
and UO_321 (O_321,N_19219,N_19768);
and UO_322 (O_322,N_19976,N_19649);
and UO_323 (O_323,N_19810,N_19921);
and UO_324 (O_324,N_19715,N_19906);
nor UO_325 (O_325,N_19376,N_19949);
nor UO_326 (O_326,N_19704,N_19271);
xor UO_327 (O_327,N_19411,N_19532);
xnor UO_328 (O_328,N_19909,N_19221);
xnor UO_329 (O_329,N_19594,N_19331);
xor UO_330 (O_330,N_19710,N_19474);
and UO_331 (O_331,N_19746,N_19362);
xor UO_332 (O_332,N_19691,N_19239);
nor UO_333 (O_333,N_19352,N_19425);
nand UO_334 (O_334,N_19476,N_19437);
and UO_335 (O_335,N_19899,N_19574);
nand UO_336 (O_336,N_19238,N_19409);
xnor UO_337 (O_337,N_19675,N_19258);
xor UO_338 (O_338,N_19452,N_19670);
nor UO_339 (O_339,N_19885,N_19693);
xor UO_340 (O_340,N_19716,N_19622);
or UO_341 (O_341,N_19910,N_19823);
and UO_342 (O_342,N_19202,N_19541);
nor UO_343 (O_343,N_19284,N_19942);
and UO_344 (O_344,N_19455,N_19621);
or UO_345 (O_345,N_19652,N_19785);
xor UO_346 (O_346,N_19683,N_19251);
xnor UO_347 (O_347,N_19931,N_19643);
xor UO_348 (O_348,N_19424,N_19402);
nor UO_349 (O_349,N_19980,N_19300);
or UO_350 (O_350,N_19998,N_19903);
xor UO_351 (O_351,N_19317,N_19570);
xnor UO_352 (O_352,N_19265,N_19517);
nor UO_353 (O_353,N_19639,N_19201);
nand UO_354 (O_354,N_19244,N_19713);
and UO_355 (O_355,N_19503,N_19418);
xor UO_356 (O_356,N_19330,N_19992);
nor UO_357 (O_357,N_19978,N_19664);
nor UO_358 (O_358,N_19739,N_19274);
or UO_359 (O_359,N_19559,N_19529);
xnor UO_360 (O_360,N_19629,N_19842);
xor UO_361 (O_361,N_19582,N_19562);
and UO_362 (O_362,N_19977,N_19611);
or UO_363 (O_363,N_19959,N_19898);
nor UO_364 (O_364,N_19753,N_19982);
and UO_365 (O_365,N_19973,N_19287);
xor UO_366 (O_366,N_19816,N_19454);
or UO_367 (O_367,N_19654,N_19831);
nand UO_368 (O_368,N_19813,N_19698);
nor UO_369 (O_369,N_19267,N_19656);
xor UO_370 (O_370,N_19841,N_19990);
or UO_371 (O_371,N_19623,N_19881);
xor UO_372 (O_372,N_19893,N_19564);
or UO_373 (O_373,N_19313,N_19807);
nor UO_374 (O_374,N_19333,N_19549);
and UO_375 (O_375,N_19806,N_19435);
nand UO_376 (O_376,N_19951,N_19328);
xnor UO_377 (O_377,N_19368,N_19617);
and UO_378 (O_378,N_19864,N_19363);
xnor UO_379 (O_379,N_19262,N_19505);
xnor UO_380 (O_380,N_19755,N_19344);
nand UO_381 (O_381,N_19370,N_19876);
and UO_382 (O_382,N_19551,N_19968);
xor UO_383 (O_383,N_19365,N_19926);
nand UO_384 (O_384,N_19870,N_19748);
xor UO_385 (O_385,N_19811,N_19789);
and UO_386 (O_386,N_19613,N_19548);
or UO_387 (O_387,N_19305,N_19512);
xnor UO_388 (O_388,N_19589,N_19464);
nand UO_389 (O_389,N_19961,N_19478);
nand UO_390 (O_390,N_19290,N_19943);
and UO_391 (O_391,N_19690,N_19708);
nand UO_392 (O_392,N_19862,N_19692);
and UO_393 (O_393,N_19975,N_19932);
xor UO_394 (O_394,N_19854,N_19230);
nor UO_395 (O_395,N_19829,N_19669);
and UO_396 (O_396,N_19848,N_19460);
nand UO_397 (O_397,N_19390,N_19688);
xor UO_398 (O_398,N_19216,N_19285);
xnor UO_399 (O_399,N_19827,N_19385);
and UO_400 (O_400,N_19821,N_19734);
nand UO_401 (O_401,N_19329,N_19295);
nor UO_402 (O_402,N_19656,N_19290);
nand UO_403 (O_403,N_19853,N_19906);
nand UO_404 (O_404,N_19705,N_19879);
nor UO_405 (O_405,N_19450,N_19604);
or UO_406 (O_406,N_19522,N_19570);
nand UO_407 (O_407,N_19957,N_19988);
nor UO_408 (O_408,N_19566,N_19348);
xnor UO_409 (O_409,N_19709,N_19761);
or UO_410 (O_410,N_19220,N_19405);
nor UO_411 (O_411,N_19732,N_19969);
or UO_412 (O_412,N_19742,N_19730);
or UO_413 (O_413,N_19719,N_19286);
or UO_414 (O_414,N_19422,N_19967);
or UO_415 (O_415,N_19400,N_19411);
xnor UO_416 (O_416,N_19223,N_19869);
nor UO_417 (O_417,N_19847,N_19644);
xor UO_418 (O_418,N_19806,N_19831);
or UO_419 (O_419,N_19970,N_19352);
xor UO_420 (O_420,N_19964,N_19854);
or UO_421 (O_421,N_19525,N_19823);
and UO_422 (O_422,N_19856,N_19378);
nor UO_423 (O_423,N_19799,N_19403);
or UO_424 (O_424,N_19811,N_19508);
nand UO_425 (O_425,N_19974,N_19566);
nor UO_426 (O_426,N_19354,N_19425);
nand UO_427 (O_427,N_19265,N_19499);
or UO_428 (O_428,N_19288,N_19292);
nand UO_429 (O_429,N_19301,N_19732);
and UO_430 (O_430,N_19921,N_19918);
nor UO_431 (O_431,N_19738,N_19982);
and UO_432 (O_432,N_19887,N_19470);
nor UO_433 (O_433,N_19392,N_19783);
xor UO_434 (O_434,N_19918,N_19896);
nor UO_435 (O_435,N_19388,N_19513);
or UO_436 (O_436,N_19681,N_19543);
nand UO_437 (O_437,N_19320,N_19976);
and UO_438 (O_438,N_19615,N_19453);
or UO_439 (O_439,N_19480,N_19744);
nor UO_440 (O_440,N_19342,N_19471);
or UO_441 (O_441,N_19584,N_19835);
or UO_442 (O_442,N_19749,N_19979);
xor UO_443 (O_443,N_19525,N_19750);
nor UO_444 (O_444,N_19359,N_19367);
and UO_445 (O_445,N_19697,N_19370);
xnor UO_446 (O_446,N_19637,N_19836);
or UO_447 (O_447,N_19575,N_19266);
xor UO_448 (O_448,N_19334,N_19341);
nand UO_449 (O_449,N_19749,N_19620);
and UO_450 (O_450,N_19660,N_19617);
nor UO_451 (O_451,N_19783,N_19951);
nand UO_452 (O_452,N_19983,N_19315);
xor UO_453 (O_453,N_19628,N_19733);
nor UO_454 (O_454,N_19602,N_19308);
xor UO_455 (O_455,N_19512,N_19922);
and UO_456 (O_456,N_19298,N_19583);
nor UO_457 (O_457,N_19801,N_19586);
xor UO_458 (O_458,N_19399,N_19910);
xnor UO_459 (O_459,N_19501,N_19441);
xor UO_460 (O_460,N_19644,N_19371);
nand UO_461 (O_461,N_19810,N_19479);
or UO_462 (O_462,N_19836,N_19898);
nand UO_463 (O_463,N_19301,N_19203);
or UO_464 (O_464,N_19309,N_19769);
or UO_465 (O_465,N_19914,N_19605);
xnor UO_466 (O_466,N_19718,N_19311);
and UO_467 (O_467,N_19577,N_19468);
or UO_468 (O_468,N_19239,N_19491);
nor UO_469 (O_469,N_19790,N_19423);
and UO_470 (O_470,N_19246,N_19322);
and UO_471 (O_471,N_19256,N_19587);
or UO_472 (O_472,N_19299,N_19724);
xnor UO_473 (O_473,N_19700,N_19931);
xnor UO_474 (O_474,N_19705,N_19808);
and UO_475 (O_475,N_19214,N_19281);
and UO_476 (O_476,N_19822,N_19651);
and UO_477 (O_477,N_19786,N_19492);
nand UO_478 (O_478,N_19761,N_19931);
nor UO_479 (O_479,N_19855,N_19851);
xor UO_480 (O_480,N_19265,N_19796);
and UO_481 (O_481,N_19284,N_19887);
or UO_482 (O_482,N_19880,N_19691);
nand UO_483 (O_483,N_19978,N_19840);
and UO_484 (O_484,N_19273,N_19320);
and UO_485 (O_485,N_19600,N_19369);
nor UO_486 (O_486,N_19345,N_19821);
xnor UO_487 (O_487,N_19661,N_19690);
or UO_488 (O_488,N_19443,N_19864);
and UO_489 (O_489,N_19770,N_19566);
and UO_490 (O_490,N_19893,N_19735);
nor UO_491 (O_491,N_19477,N_19703);
nand UO_492 (O_492,N_19836,N_19429);
or UO_493 (O_493,N_19259,N_19721);
nand UO_494 (O_494,N_19856,N_19269);
nor UO_495 (O_495,N_19487,N_19579);
xor UO_496 (O_496,N_19352,N_19608);
or UO_497 (O_497,N_19577,N_19650);
nor UO_498 (O_498,N_19715,N_19229);
and UO_499 (O_499,N_19332,N_19723);
and UO_500 (O_500,N_19380,N_19514);
nor UO_501 (O_501,N_19564,N_19905);
xnor UO_502 (O_502,N_19974,N_19919);
and UO_503 (O_503,N_19783,N_19451);
xor UO_504 (O_504,N_19517,N_19464);
xor UO_505 (O_505,N_19213,N_19592);
nor UO_506 (O_506,N_19656,N_19801);
or UO_507 (O_507,N_19592,N_19925);
or UO_508 (O_508,N_19451,N_19245);
nand UO_509 (O_509,N_19497,N_19321);
or UO_510 (O_510,N_19404,N_19400);
nor UO_511 (O_511,N_19736,N_19287);
or UO_512 (O_512,N_19999,N_19753);
nor UO_513 (O_513,N_19443,N_19690);
nor UO_514 (O_514,N_19228,N_19309);
xor UO_515 (O_515,N_19664,N_19412);
xnor UO_516 (O_516,N_19879,N_19459);
xnor UO_517 (O_517,N_19683,N_19423);
nand UO_518 (O_518,N_19801,N_19477);
nand UO_519 (O_519,N_19975,N_19985);
xnor UO_520 (O_520,N_19978,N_19628);
or UO_521 (O_521,N_19311,N_19241);
xor UO_522 (O_522,N_19312,N_19473);
nand UO_523 (O_523,N_19469,N_19311);
and UO_524 (O_524,N_19360,N_19897);
or UO_525 (O_525,N_19726,N_19413);
and UO_526 (O_526,N_19738,N_19894);
and UO_527 (O_527,N_19477,N_19795);
nor UO_528 (O_528,N_19511,N_19682);
nand UO_529 (O_529,N_19393,N_19566);
or UO_530 (O_530,N_19258,N_19844);
xor UO_531 (O_531,N_19613,N_19867);
nor UO_532 (O_532,N_19573,N_19728);
xor UO_533 (O_533,N_19652,N_19362);
or UO_534 (O_534,N_19960,N_19227);
nor UO_535 (O_535,N_19664,N_19801);
nand UO_536 (O_536,N_19667,N_19556);
xnor UO_537 (O_537,N_19352,N_19952);
xor UO_538 (O_538,N_19595,N_19653);
and UO_539 (O_539,N_19805,N_19229);
and UO_540 (O_540,N_19711,N_19419);
nor UO_541 (O_541,N_19976,N_19837);
or UO_542 (O_542,N_19545,N_19387);
xor UO_543 (O_543,N_19257,N_19583);
nor UO_544 (O_544,N_19388,N_19667);
and UO_545 (O_545,N_19748,N_19745);
or UO_546 (O_546,N_19445,N_19441);
and UO_547 (O_547,N_19470,N_19366);
nand UO_548 (O_548,N_19457,N_19948);
nor UO_549 (O_549,N_19589,N_19521);
nand UO_550 (O_550,N_19356,N_19388);
and UO_551 (O_551,N_19705,N_19234);
or UO_552 (O_552,N_19374,N_19567);
and UO_553 (O_553,N_19450,N_19852);
nand UO_554 (O_554,N_19226,N_19854);
or UO_555 (O_555,N_19696,N_19433);
nor UO_556 (O_556,N_19417,N_19394);
nor UO_557 (O_557,N_19575,N_19298);
nand UO_558 (O_558,N_19658,N_19435);
xor UO_559 (O_559,N_19709,N_19873);
or UO_560 (O_560,N_19579,N_19362);
and UO_561 (O_561,N_19680,N_19837);
nand UO_562 (O_562,N_19828,N_19454);
nor UO_563 (O_563,N_19625,N_19703);
and UO_564 (O_564,N_19721,N_19232);
xnor UO_565 (O_565,N_19749,N_19841);
xnor UO_566 (O_566,N_19971,N_19643);
and UO_567 (O_567,N_19261,N_19929);
xnor UO_568 (O_568,N_19884,N_19290);
xnor UO_569 (O_569,N_19714,N_19268);
nor UO_570 (O_570,N_19766,N_19426);
nand UO_571 (O_571,N_19441,N_19747);
or UO_572 (O_572,N_19373,N_19968);
or UO_573 (O_573,N_19881,N_19934);
and UO_574 (O_574,N_19532,N_19947);
and UO_575 (O_575,N_19745,N_19603);
nand UO_576 (O_576,N_19348,N_19555);
xnor UO_577 (O_577,N_19703,N_19533);
or UO_578 (O_578,N_19777,N_19662);
and UO_579 (O_579,N_19216,N_19998);
and UO_580 (O_580,N_19503,N_19800);
xnor UO_581 (O_581,N_19410,N_19711);
or UO_582 (O_582,N_19846,N_19855);
nor UO_583 (O_583,N_19797,N_19288);
and UO_584 (O_584,N_19839,N_19590);
or UO_585 (O_585,N_19544,N_19438);
xor UO_586 (O_586,N_19213,N_19770);
or UO_587 (O_587,N_19538,N_19547);
nand UO_588 (O_588,N_19314,N_19270);
nor UO_589 (O_589,N_19967,N_19741);
xnor UO_590 (O_590,N_19257,N_19896);
or UO_591 (O_591,N_19834,N_19697);
or UO_592 (O_592,N_19839,N_19507);
nor UO_593 (O_593,N_19381,N_19270);
and UO_594 (O_594,N_19678,N_19483);
nand UO_595 (O_595,N_19226,N_19379);
or UO_596 (O_596,N_19977,N_19231);
or UO_597 (O_597,N_19328,N_19758);
nor UO_598 (O_598,N_19435,N_19520);
and UO_599 (O_599,N_19731,N_19631);
nand UO_600 (O_600,N_19617,N_19684);
or UO_601 (O_601,N_19951,N_19723);
xnor UO_602 (O_602,N_19715,N_19773);
or UO_603 (O_603,N_19434,N_19541);
and UO_604 (O_604,N_19721,N_19379);
or UO_605 (O_605,N_19657,N_19226);
or UO_606 (O_606,N_19233,N_19514);
and UO_607 (O_607,N_19431,N_19874);
and UO_608 (O_608,N_19628,N_19213);
nand UO_609 (O_609,N_19943,N_19673);
nor UO_610 (O_610,N_19899,N_19516);
or UO_611 (O_611,N_19918,N_19797);
xnor UO_612 (O_612,N_19829,N_19989);
and UO_613 (O_613,N_19888,N_19636);
nand UO_614 (O_614,N_19364,N_19541);
or UO_615 (O_615,N_19815,N_19564);
nor UO_616 (O_616,N_19597,N_19745);
and UO_617 (O_617,N_19690,N_19232);
nand UO_618 (O_618,N_19483,N_19836);
xnor UO_619 (O_619,N_19289,N_19979);
and UO_620 (O_620,N_19808,N_19884);
or UO_621 (O_621,N_19366,N_19978);
nor UO_622 (O_622,N_19412,N_19892);
or UO_623 (O_623,N_19649,N_19229);
and UO_624 (O_624,N_19217,N_19556);
or UO_625 (O_625,N_19480,N_19518);
nand UO_626 (O_626,N_19315,N_19469);
nor UO_627 (O_627,N_19365,N_19909);
xnor UO_628 (O_628,N_19880,N_19972);
nor UO_629 (O_629,N_19868,N_19873);
nand UO_630 (O_630,N_19783,N_19611);
and UO_631 (O_631,N_19419,N_19921);
or UO_632 (O_632,N_19516,N_19957);
nor UO_633 (O_633,N_19248,N_19996);
and UO_634 (O_634,N_19657,N_19671);
nand UO_635 (O_635,N_19963,N_19907);
or UO_636 (O_636,N_19850,N_19515);
nor UO_637 (O_637,N_19278,N_19806);
or UO_638 (O_638,N_19639,N_19891);
nor UO_639 (O_639,N_19838,N_19667);
nand UO_640 (O_640,N_19528,N_19386);
xor UO_641 (O_641,N_19909,N_19408);
or UO_642 (O_642,N_19961,N_19344);
nor UO_643 (O_643,N_19574,N_19670);
xnor UO_644 (O_644,N_19852,N_19996);
nand UO_645 (O_645,N_19204,N_19333);
and UO_646 (O_646,N_19518,N_19606);
xor UO_647 (O_647,N_19240,N_19303);
or UO_648 (O_648,N_19498,N_19326);
nand UO_649 (O_649,N_19379,N_19448);
nand UO_650 (O_650,N_19412,N_19670);
nor UO_651 (O_651,N_19400,N_19882);
or UO_652 (O_652,N_19420,N_19246);
xnor UO_653 (O_653,N_19467,N_19627);
and UO_654 (O_654,N_19318,N_19660);
nor UO_655 (O_655,N_19592,N_19807);
nand UO_656 (O_656,N_19483,N_19260);
nand UO_657 (O_657,N_19683,N_19865);
xnor UO_658 (O_658,N_19469,N_19878);
nand UO_659 (O_659,N_19672,N_19302);
xnor UO_660 (O_660,N_19309,N_19740);
nand UO_661 (O_661,N_19522,N_19519);
and UO_662 (O_662,N_19891,N_19325);
nor UO_663 (O_663,N_19596,N_19559);
nor UO_664 (O_664,N_19568,N_19578);
xor UO_665 (O_665,N_19578,N_19838);
nand UO_666 (O_666,N_19642,N_19786);
nor UO_667 (O_667,N_19883,N_19442);
nor UO_668 (O_668,N_19574,N_19960);
nand UO_669 (O_669,N_19449,N_19660);
xor UO_670 (O_670,N_19419,N_19331);
nor UO_671 (O_671,N_19706,N_19296);
xor UO_672 (O_672,N_19420,N_19827);
or UO_673 (O_673,N_19289,N_19452);
nand UO_674 (O_674,N_19584,N_19487);
xor UO_675 (O_675,N_19555,N_19593);
nor UO_676 (O_676,N_19664,N_19409);
and UO_677 (O_677,N_19999,N_19872);
nor UO_678 (O_678,N_19400,N_19551);
xnor UO_679 (O_679,N_19798,N_19579);
nor UO_680 (O_680,N_19368,N_19310);
and UO_681 (O_681,N_19932,N_19293);
and UO_682 (O_682,N_19781,N_19575);
or UO_683 (O_683,N_19239,N_19760);
nor UO_684 (O_684,N_19729,N_19404);
nor UO_685 (O_685,N_19952,N_19954);
and UO_686 (O_686,N_19632,N_19586);
nand UO_687 (O_687,N_19941,N_19374);
and UO_688 (O_688,N_19630,N_19846);
and UO_689 (O_689,N_19229,N_19849);
and UO_690 (O_690,N_19722,N_19937);
and UO_691 (O_691,N_19810,N_19531);
nor UO_692 (O_692,N_19278,N_19625);
xnor UO_693 (O_693,N_19250,N_19398);
nand UO_694 (O_694,N_19950,N_19816);
nand UO_695 (O_695,N_19907,N_19807);
xnor UO_696 (O_696,N_19420,N_19890);
and UO_697 (O_697,N_19810,N_19626);
xor UO_698 (O_698,N_19924,N_19779);
and UO_699 (O_699,N_19307,N_19570);
or UO_700 (O_700,N_19305,N_19452);
nand UO_701 (O_701,N_19611,N_19443);
nand UO_702 (O_702,N_19424,N_19939);
nand UO_703 (O_703,N_19550,N_19451);
xor UO_704 (O_704,N_19864,N_19715);
xnor UO_705 (O_705,N_19458,N_19829);
xor UO_706 (O_706,N_19342,N_19399);
nor UO_707 (O_707,N_19774,N_19985);
xor UO_708 (O_708,N_19776,N_19458);
and UO_709 (O_709,N_19637,N_19967);
or UO_710 (O_710,N_19550,N_19887);
or UO_711 (O_711,N_19883,N_19612);
xor UO_712 (O_712,N_19395,N_19901);
and UO_713 (O_713,N_19631,N_19449);
or UO_714 (O_714,N_19527,N_19431);
xnor UO_715 (O_715,N_19343,N_19684);
or UO_716 (O_716,N_19655,N_19503);
nand UO_717 (O_717,N_19280,N_19703);
and UO_718 (O_718,N_19939,N_19742);
nor UO_719 (O_719,N_19750,N_19786);
nor UO_720 (O_720,N_19351,N_19813);
or UO_721 (O_721,N_19979,N_19661);
nor UO_722 (O_722,N_19271,N_19597);
or UO_723 (O_723,N_19804,N_19473);
or UO_724 (O_724,N_19671,N_19464);
or UO_725 (O_725,N_19791,N_19743);
nand UO_726 (O_726,N_19740,N_19311);
nand UO_727 (O_727,N_19249,N_19232);
or UO_728 (O_728,N_19583,N_19415);
and UO_729 (O_729,N_19214,N_19271);
xor UO_730 (O_730,N_19612,N_19521);
nand UO_731 (O_731,N_19824,N_19424);
xnor UO_732 (O_732,N_19473,N_19812);
nor UO_733 (O_733,N_19844,N_19999);
or UO_734 (O_734,N_19636,N_19405);
and UO_735 (O_735,N_19559,N_19511);
xor UO_736 (O_736,N_19751,N_19542);
and UO_737 (O_737,N_19579,N_19727);
and UO_738 (O_738,N_19582,N_19629);
and UO_739 (O_739,N_19528,N_19247);
and UO_740 (O_740,N_19520,N_19405);
nor UO_741 (O_741,N_19504,N_19764);
nor UO_742 (O_742,N_19449,N_19299);
or UO_743 (O_743,N_19543,N_19403);
nor UO_744 (O_744,N_19836,N_19228);
xor UO_745 (O_745,N_19283,N_19609);
and UO_746 (O_746,N_19237,N_19805);
or UO_747 (O_747,N_19772,N_19528);
xnor UO_748 (O_748,N_19702,N_19411);
and UO_749 (O_749,N_19582,N_19392);
or UO_750 (O_750,N_19352,N_19572);
xor UO_751 (O_751,N_19317,N_19228);
nand UO_752 (O_752,N_19385,N_19455);
or UO_753 (O_753,N_19627,N_19816);
or UO_754 (O_754,N_19407,N_19204);
nor UO_755 (O_755,N_19489,N_19543);
nor UO_756 (O_756,N_19874,N_19365);
and UO_757 (O_757,N_19418,N_19296);
nor UO_758 (O_758,N_19803,N_19544);
and UO_759 (O_759,N_19254,N_19696);
xnor UO_760 (O_760,N_19764,N_19599);
or UO_761 (O_761,N_19847,N_19404);
nand UO_762 (O_762,N_19232,N_19945);
nand UO_763 (O_763,N_19407,N_19637);
xnor UO_764 (O_764,N_19654,N_19276);
and UO_765 (O_765,N_19457,N_19863);
nor UO_766 (O_766,N_19641,N_19812);
nor UO_767 (O_767,N_19658,N_19375);
and UO_768 (O_768,N_19236,N_19745);
nand UO_769 (O_769,N_19369,N_19680);
nand UO_770 (O_770,N_19217,N_19518);
and UO_771 (O_771,N_19753,N_19722);
xnor UO_772 (O_772,N_19396,N_19291);
or UO_773 (O_773,N_19464,N_19489);
and UO_774 (O_774,N_19461,N_19731);
xnor UO_775 (O_775,N_19748,N_19507);
or UO_776 (O_776,N_19437,N_19501);
nand UO_777 (O_777,N_19720,N_19393);
or UO_778 (O_778,N_19958,N_19632);
xnor UO_779 (O_779,N_19523,N_19837);
nand UO_780 (O_780,N_19885,N_19406);
nand UO_781 (O_781,N_19258,N_19310);
xor UO_782 (O_782,N_19922,N_19975);
nor UO_783 (O_783,N_19456,N_19462);
nand UO_784 (O_784,N_19377,N_19460);
and UO_785 (O_785,N_19816,N_19250);
xnor UO_786 (O_786,N_19404,N_19651);
or UO_787 (O_787,N_19202,N_19646);
nor UO_788 (O_788,N_19673,N_19819);
xor UO_789 (O_789,N_19358,N_19738);
and UO_790 (O_790,N_19986,N_19983);
nor UO_791 (O_791,N_19732,N_19432);
nor UO_792 (O_792,N_19855,N_19356);
nand UO_793 (O_793,N_19540,N_19237);
nor UO_794 (O_794,N_19976,N_19366);
nand UO_795 (O_795,N_19558,N_19944);
nand UO_796 (O_796,N_19665,N_19630);
xnor UO_797 (O_797,N_19382,N_19572);
or UO_798 (O_798,N_19861,N_19924);
nand UO_799 (O_799,N_19955,N_19697);
nor UO_800 (O_800,N_19739,N_19270);
and UO_801 (O_801,N_19530,N_19573);
xnor UO_802 (O_802,N_19297,N_19451);
xor UO_803 (O_803,N_19715,N_19946);
nand UO_804 (O_804,N_19764,N_19277);
nor UO_805 (O_805,N_19442,N_19793);
nor UO_806 (O_806,N_19808,N_19445);
nor UO_807 (O_807,N_19219,N_19239);
nand UO_808 (O_808,N_19553,N_19470);
or UO_809 (O_809,N_19390,N_19318);
and UO_810 (O_810,N_19469,N_19760);
xnor UO_811 (O_811,N_19274,N_19230);
nor UO_812 (O_812,N_19872,N_19556);
nor UO_813 (O_813,N_19282,N_19824);
nor UO_814 (O_814,N_19858,N_19814);
nor UO_815 (O_815,N_19711,N_19406);
nor UO_816 (O_816,N_19678,N_19204);
or UO_817 (O_817,N_19795,N_19768);
nand UO_818 (O_818,N_19707,N_19605);
xnor UO_819 (O_819,N_19687,N_19714);
nand UO_820 (O_820,N_19892,N_19331);
xnor UO_821 (O_821,N_19822,N_19329);
nand UO_822 (O_822,N_19249,N_19620);
nand UO_823 (O_823,N_19466,N_19947);
nand UO_824 (O_824,N_19776,N_19259);
nor UO_825 (O_825,N_19602,N_19970);
nand UO_826 (O_826,N_19603,N_19970);
and UO_827 (O_827,N_19324,N_19432);
and UO_828 (O_828,N_19295,N_19926);
xor UO_829 (O_829,N_19791,N_19521);
nor UO_830 (O_830,N_19654,N_19675);
or UO_831 (O_831,N_19339,N_19885);
or UO_832 (O_832,N_19410,N_19279);
nand UO_833 (O_833,N_19762,N_19788);
nor UO_834 (O_834,N_19509,N_19894);
nand UO_835 (O_835,N_19847,N_19205);
xor UO_836 (O_836,N_19336,N_19561);
nand UO_837 (O_837,N_19884,N_19623);
and UO_838 (O_838,N_19598,N_19829);
nand UO_839 (O_839,N_19439,N_19912);
nand UO_840 (O_840,N_19597,N_19432);
xnor UO_841 (O_841,N_19871,N_19863);
or UO_842 (O_842,N_19931,N_19984);
xnor UO_843 (O_843,N_19687,N_19539);
and UO_844 (O_844,N_19898,N_19309);
and UO_845 (O_845,N_19252,N_19721);
nor UO_846 (O_846,N_19348,N_19683);
nor UO_847 (O_847,N_19647,N_19842);
nor UO_848 (O_848,N_19535,N_19775);
nor UO_849 (O_849,N_19545,N_19379);
nand UO_850 (O_850,N_19340,N_19619);
and UO_851 (O_851,N_19484,N_19550);
or UO_852 (O_852,N_19430,N_19671);
nor UO_853 (O_853,N_19987,N_19669);
or UO_854 (O_854,N_19362,N_19892);
xor UO_855 (O_855,N_19552,N_19983);
or UO_856 (O_856,N_19897,N_19670);
and UO_857 (O_857,N_19950,N_19982);
xnor UO_858 (O_858,N_19625,N_19552);
nor UO_859 (O_859,N_19439,N_19312);
nor UO_860 (O_860,N_19491,N_19574);
xnor UO_861 (O_861,N_19632,N_19773);
and UO_862 (O_862,N_19226,N_19323);
and UO_863 (O_863,N_19702,N_19965);
xnor UO_864 (O_864,N_19680,N_19928);
xor UO_865 (O_865,N_19204,N_19954);
and UO_866 (O_866,N_19761,N_19260);
nand UO_867 (O_867,N_19967,N_19235);
nor UO_868 (O_868,N_19372,N_19334);
nor UO_869 (O_869,N_19244,N_19990);
nand UO_870 (O_870,N_19931,N_19538);
nand UO_871 (O_871,N_19999,N_19691);
xnor UO_872 (O_872,N_19945,N_19555);
or UO_873 (O_873,N_19430,N_19260);
and UO_874 (O_874,N_19508,N_19457);
and UO_875 (O_875,N_19719,N_19616);
and UO_876 (O_876,N_19551,N_19931);
nand UO_877 (O_877,N_19332,N_19822);
nor UO_878 (O_878,N_19328,N_19811);
xnor UO_879 (O_879,N_19368,N_19594);
nand UO_880 (O_880,N_19875,N_19439);
and UO_881 (O_881,N_19440,N_19780);
and UO_882 (O_882,N_19982,N_19861);
nand UO_883 (O_883,N_19319,N_19675);
nor UO_884 (O_884,N_19576,N_19411);
nand UO_885 (O_885,N_19452,N_19567);
nand UO_886 (O_886,N_19552,N_19300);
xnor UO_887 (O_887,N_19989,N_19544);
and UO_888 (O_888,N_19777,N_19703);
and UO_889 (O_889,N_19303,N_19746);
or UO_890 (O_890,N_19821,N_19425);
nand UO_891 (O_891,N_19505,N_19841);
and UO_892 (O_892,N_19357,N_19583);
and UO_893 (O_893,N_19232,N_19914);
and UO_894 (O_894,N_19262,N_19252);
nand UO_895 (O_895,N_19867,N_19786);
or UO_896 (O_896,N_19767,N_19723);
and UO_897 (O_897,N_19210,N_19420);
xor UO_898 (O_898,N_19262,N_19336);
and UO_899 (O_899,N_19902,N_19765);
xor UO_900 (O_900,N_19411,N_19361);
nor UO_901 (O_901,N_19499,N_19687);
or UO_902 (O_902,N_19526,N_19400);
xor UO_903 (O_903,N_19788,N_19370);
or UO_904 (O_904,N_19661,N_19992);
xor UO_905 (O_905,N_19344,N_19257);
nor UO_906 (O_906,N_19513,N_19423);
or UO_907 (O_907,N_19481,N_19714);
nand UO_908 (O_908,N_19909,N_19774);
and UO_909 (O_909,N_19326,N_19933);
xnor UO_910 (O_910,N_19764,N_19286);
nand UO_911 (O_911,N_19432,N_19717);
nor UO_912 (O_912,N_19531,N_19977);
or UO_913 (O_913,N_19539,N_19818);
nand UO_914 (O_914,N_19337,N_19761);
or UO_915 (O_915,N_19616,N_19685);
nor UO_916 (O_916,N_19320,N_19834);
nand UO_917 (O_917,N_19857,N_19413);
nor UO_918 (O_918,N_19542,N_19883);
nor UO_919 (O_919,N_19624,N_19556);
and UO_920 (O_920,N_19635,N_19701);
and UO_921 (O_921,N_19831,N_19552);
and UO_922 (O_922,N_19488,N_19552);
and UO_923 (O_923,N_19675,N_19935);
xor UO_924 (O_924,N_19970,N_19228);
xor UO_925 (O_925,N_19826,N_19667);
and UO_926 (O_926,N_19837,N_19420);
or UO_927 (O_927,N_19954,N_19284);
or UO_928 (O_928,N_19292,N_19470);
nand UO_929 (O_929,N_19490,N_19218);
nand UO_930 (O_930,N_19650,N_19634);
nor UO_931 (O_931,N_19736,N_19787);
and UO_932 (O_932,N_19561,N_19430);
xnor UO_933 (O_933,N_19335,N_19259);
xor UO_934 (O_934,N_19484,N_19313);
xnor UO_935 (O_935,N_19653,N_19787);
or UO_936 (O_936,N_19702,N_19432);
and UO_937 (O_937,N_19505,N_19806);
nor UO_938 (O_938,N_19208,N_19450);
xor UO_939 (O_939,N_19858,N_19394);
nor UO_940 (O_940,N_19256,N_19555);
nand UO_941 (O_941,N_19780,N_19322);
xnor UO_942 (O_942,N_19268,N_19517);
or UO_943 (O_943,N_19781,N_19701);
and UO_944 (O_944,N_19710,N_19790);
and UO_945 (O_945,N_19984,N_19983);
nor UO_946 (O_946,N_19697,N_19264);
nor UO_947 (O_947,N_19832,N_19839);
nand UO_948 (O_948,N_19856,N_19368);
nand UO_949 (O_949,N_19806,N_19217);
and UO_950 (O_950,N_19482,N_19538);
and UO_951 (O_951,N_19533,N_19259);
nor UO_952 (O_952,N_19845,N_19519);
xor UO_953 (O_953,N_19633,N_19276);
and UO_954 (O_954,N_19226,N_19465);
xnor UO_955 (O_955,N_19517,N_19500);
or UO_956 (O_956,N_19549,N_19695);
nand UO_957 (O_957,N_19913,N_19629);
nor UO_958 (O_958,N_19369,N_19206);
nor UO_959 (O_959,N_19849,N_19809);
nand UO_960 (O_960,N_19398,N_19446);
nor UO_961 (O_961,N_19504,N_19689);
or UO_962 (O_962,N_19381,N_19781);
nand UO_963 (O_963,N_19878,N_19675);
or UO_964 (O_964,N_19592,N_19762);
xor UO_965 (O_965,N_19378,N_19715);
or UO_966 (O_966,N_19759,N_19596);
and UO_967 (O_967,N_19935,N_19888);
nor UO_968 (O_968,N_19278,N_19729);
nor UO_969 (O_969,N_19968,N_19890);
nand UO_970 (O_970,N_19206,N_19493);
or UO_971 (O_971,N_19714,N_19783);
or UO_972 (O_972,N_19936,N_19833);
and UO_973 (O_973,N_19452,N_19599);
nand UO_974 (O_974,N_19651,N_19679);
or UO_975 (O_975,N_19833,N_19942);
or UO_976 (O_976,N_19259,N_19995);
or UO_977 (O_977,N_19865,N_19503);
or UO_978 (O_978,N_19909,N_19563);
xnor UO_979 (O_979,N_19214,N_19940);
nand UO_980 (O_980,N_19338,N_19706);
or UO_981 (O_981,N_19638,N_19574);
nor UO_982 (O_982,N_19823,N_19386);
and UO_983 (O_983,N_19891,N_19502);
nor UO_984 (O_984,N_19417,N_19364);
nor UO_985 (O_985,N_19698,N_19219);
and UO_986 (O_986,N_19568,N_19708);
nor UO_987 (O_987,N_19901,N_19885);
xor UO_988 (O_988,N_19643,N_19964);
and UO_989 (O_989,N_19365,N_19388);
or UO_990 (O_990,N_19878,N_19697);
or UO_991 (O_991,N_19388,N_19793);
xnor UO_992 (O_992,N_19722,N_19263);
and UO_993 (O_993,N_19253,N_19283);
xor UO_994 (O_994,N_19316,N_19512);
nor UO_995 (O_995,N_19934,N_19432);
and UO_996 (O_996,N_19647,N_19674);
nand UO_997 (O_997,N_19703,N_19262);
nand UO_998 (O_998,N_19747,N_19371);
or UO_999 (O_999,N_19606,N_19383);
nand UO_1000 (O_1000,N_19827,N_19363);
or UO_1001 (O_1001,N_19974,N_19519);
nand UO_1002 (O_1002,N_19512,N_19553);
nand UO_1003 (O_1003,N_19238,N_19420);
nand UO_1004 (O_1004,N_19478,N_19249);
nand UO_1005 (O_1005,N_19738,N_19717);
and UO_1006 (O_1006,N_19700,N_19689);
or UO_1007 (O_1007,N_19491,N_19920);
nor UO_1008 (O_1008,N_19838,N_19964);
nor UO_1009 (O_1009,N_19761,N_19553);
xnor UO_1010 (O_1010,N_19255,N_19256);
xnor UO_1011 (O_1011,N_19936,N_19712);
or UO_1012 (O_1012,N_19227,N_19779);
or UO_1013 (O_1013,N_19256,N_19721);
nor UO_1014 (O_1014,N_19894,N_19678);
nor UO_1015 (O_1015,N_19348,N_19922);
or UO_1016 (O_1016,N_19395,N_19983);
or UO_1017 (O_1017,N_19974,N_19657);
nor UO_1018 (O_1018,N_19483,N_19745);
nor UO_1019 (O_1019,N_19451,N_19898);
xor UO_1020 (O_1020,N_19424,N_19861);
and UO_1021 (O_1021,N_19321,N_19714);
and UO_1022 (O_1022,N_19441,N_19666);
or UO_1023 (O_1023,N_19868,N_19871);
and UO_1024 (O_1024,N_19379,N_19843);
nor UO_1025 (O_1025,N_19676,N_19791);
xor UO_1026 (O_1026,N_19297,N_19440);
nor UO_1027 (O_1027,N_19728,N_19203);
and UO_1028 (O_1028,N_19491,N_19926);
nor UO_1029 (O_1029,N_19487,N_19208);
nand UO_1030 (O_1030,N_19531,N_19214);
nand UO_1031 (O_1031,N_19905,N_19618);
nand UO_1032 (O_1032,N_19721,N_19315);
xor UO_1033 (O_1033,N_19607,N_19608);
xnor UO_1034 (O_1034,N_19644,N_19810);
or UO_1035 (O_1035,N_19997,N_19336);
and UO_1036 (O_1036,N_19738,N_19294);
or UO_1037 (O_1037,N_19372,N_19401);
xnor UO_1038 (O_1038,N_19849,N_19733);
xnor UO_1039 (O_1039,N_19307,N_19694);
and UO_1040 (O_1040,N_19492,N_19995);
nor UO_1041 (O_1041,N_19870,N_19540);
or UO_1042 (O_1042,N_19978,N_19868);
nor UO_1043 (O_1043,N_19539,N_19667);
xnor UO_1044 (O_1044,N_19642,N_19365);
xor UO_1045 (O_1045,N_19272,N_19484);
and UO_1046 (O_1046,N_19298,N_19205);
nor UO_1047 (O_1047,N_19302,N_19854);
and UO_1048 (O_1048,N_19254,N_19310);
nor UO_1049 (O_1049,N_19753,N_19778);
nand UO_1050 (O_1050,N_19832,N_19399);
xnor UO_1051 (O_1051,N_19440,N_19533);
nor UO_1052 (O_1052,N_19692,N_19360);
nand UO_1053 (O_1053,N_19992,N_19780);
xnor UO_1054 (O_1054,N_19951,N_19990);
nor UO_1055 (O_1055,N_19606,N_19784);
nand UO_1056 (O_1056,N_19400,N_19980);
or UO_1057 (O_1057,N_19215,N_19647);
or UO_1058 (O_1058,N_19919,N_19780);
xor UO_1059 (O_1059,N_19896,N_19600);
nand UO_1060 (O_1060,N_19650,N_19490);
and UO_1061 (O_1061,N_19548,N_19850);
nand UO_1062 (O_1062,N_19923,N_19284);
and UO_1063 (O_1063,N_19213,N_19952);
or UO_1064 (O_1064,N_19531,N_19974);
nor UO_1065 (O_1065,N_19993,N_19516);
and UO_1066 (O_1066,N_19417,N_19851);
nor UO_1067 (O_1067,N_19919,N_19737);
nor UO_1068 (O_1068,N_19612,N_19570);
nand UO_1069 (O_1069,N_19912,N_19552);
or UO_1070 (O_1070,N_19840,N_19738);
nand UO_1071 (O_1071,N_19908,N_19376);
and UO_1072 (O_1072,N_19724,N_19855);
or UO_1073 (O_1073,N_19995,N_19288);
nand UO_1074 (O_1074,N_19704,N_19733);
nand UO_1075 (O_1075,N_19619,N_19286);
xor UO_1076 (O_1076,N_19689,N_19283);
xor UO_1077 (O_1077,N_19591,N_19426);
nor UO_1078 (O_1078,N_19271,N_19299);
and UO_1079 (O_1079,N_19599,N_19254);
or UO_1080 (O_1080,N_19778,N_19703);
xor UO_1081 (O_1081,N_19571,N_19643);
xnor UO_1082 (O_1082,N_19764,N_19830);
nor UO_1083 (O_1083,N_19697,N_19397);
nor UO_1084 (O_1084,N_19477,N_19332);
or UO_1085 (O_1085,N_19914,N_19676);
nor UO_1086 (O_1086,N_19817,N_19588);
and UO_1087 (O_1087,N_19272,N_19482);
nor UO_1088 (O_1088,N_19460,N_19492);
xor UO_1089 (O_1089,N_19923,N_19770);
nand UO_1090 (O_1090,N_19340,N_19890);
or UO_1091 (O_1091,N_19865,N_19334);
nand UO_1092 (O_1092,N_19916,N_19338);
nand UO_1093 (O_1093,N_19463,N_19908);
and UO_1094 (O_1094,N_19690,N_19307);
and UO_1095 (O_1095,N_19552,N_19774);
xor UO_1096 (O_1096,N_19352,N_19448);
nand UO_1097 (O_1097,N_19953,N_19731);
or UO_1098 (O_1098,N_19891,N_19214);
xor UO_1099 (O_1099,N_19497,N_19676);
nand UO_1100 (O_1100,N_19273,N_19524);
nand UO_1101 (O_1101,N_19726,N_19992);
nor UO_1102 (O_1102,N_19630,N_19272);
xnor UO_1103 (O_1103,N_19540,N_19963);
xor UO_1104 (O_1104,N_19852,N_19505);
xor UO_1105 (O_1105,N_19804,N_19990);
or UO_1106 (O_1106,N_19235,N_19453);
nor UO_1107 (O_1107,N_19939,N_19724);
and UO_1108 (O_1108,N_19221,N_19343);
nand UO_1109 (O_1109,N_19997,N_19831);
xor UO_1110 (O_1110,N_19799,N_19493);
or UO_1111 (O_1111,N_19941,N_19502);
xor UO_1112 (O_1112,N_19352,N_19769);
or UO_1113 (O_1113,N_19452,N_19250);
nand UO_1114 (O_1114,N_19629,N_19523);
nor UO_1115 (O_1115,N_19789,N_19464);
nor UO_1116 (O_1116,N_19393,N_19826);
and UO_1117 (O_1117,N_19242,N_19550);
xnor UO_1118 (O_1118,N_19926,N_19414);
xor UO_1119 (O_1119,N_19320,N_19499);
or UO_1120 (O_1120,N_19861,N_19845);
and UO_1121 (O_1121,N_19696,N_19722);
nand UO_1122 (O_1122,N_19891,N_19771);
xnor UO_1123 (O_1123,N_19931,N_19333);
and UO_1124 (O_1124,N_19991,N_19211);
nand UO_1125 (O_1125,N_19402,N_19706);
nor UO_1126 (O_1126,N_19499,N_19671);
or UO_1127 (O_1127,N_19852,N_19468);
nor UO_1128 (O_1128,N_19753,N_19490);
and UO_1129 (O_1129,N_19549,N_19926);
nand UO_1130 (O_1130,N_19688,N_19821);
or UO_1131 (O_1131,N_19607,N_19304);
and UO_1132 (O_1132,N_19383,N_19437);
or UO_1133 (O_1133,N_19398,N_19467);
xor UO_1134 (O_1134,N_19769,N_19303);
and UO_1135 (O_1135,N_19723,N_19853);
and UO_1136 (O_1136,N_19375,N_19743);
nor UO_1137 (O_1137,N_19403,N_19616);
or UO_1138 (O_1138,N_19982,N_19664);
nand UO_1139 (O_1139,N_19942,N_19629);
and UO_1140 (O_1140,N_19340,N_19856);
or UO_1141 (O_1141,N_19643,N_19435);
xnor UO_1142 (O_1142,N_19548,N_19213);
nand UO_1143 (O_1143,N_19624,N_19965);
nand UO_1144 (O_1144,N_19495,N_19596);
xnor UO_1145 (O_1145,N_19821,N_19479);
nor UO_1146 (O_1146,N_19976,N_19509);
nor UO_1147 (O_1147,N_19850,N_19546);
xor UO_1148 (O_1148,N_19429,N_19787);
or UO_1149 (O_1149,N_19503,N_19263);
or UO_1150 (O_1150,N_19441,N_19873);
nor UO_1151 (O_1151,N_19692,N_19725);
xnor UO_1152 (O_1152,N_19989,N_19786);
and UO_1153 (O_1153,N_19801,N_19683);
and UO_1154 (O_1154,N_19818,N_19214);
nand UO_1155 (O_1155,N_19630,N_19950);
or UO_1156 (O_1156,N_19655,N_19904);
nor UO_1157 (O_1157,N_19336,N_19828);
and UO_1158 (O_1158,N_19536,N_19323);
xnor UO_1159 (O_1159,N_19554,N_19660);
and UO_1160 (O_1160,N_19830,N_19617);
and UO_1161 (O_1161,N_19894,N_19416);
or UO_1162 (O_1162,N_19200,N_19539);
or UO_1163 (O_1163,N_19559,N_19563);
nand UO_1164 (O_1164,N_19286,N_19945);
nor UO_1165 (O_1165,N_19486,N_19492);
nor UO_1166 (O_1166,N_19579,N_19516);
nor UO_1167 (O_1167,N_19945,N_19431);
nand UO_1168 (O_1168,N_19844,N_19708);
or UO_1169 (O_1169,N_19381,N_19924);
or UO_1170 (O_1170,N_19750,N_19437);
nand UO_1171 (O_1171,N_19486,N_19659);
and UO_1172 (O_1172,N_19638,N_19790);
xnor UO_1173 (O_1173,N_19654,N_19318);
or UO_1174 (O_1174,N_19744,N_19407);
or UO_1175 (O_1175,N_19816,N_19706);
or UO_1176 (O_1176,N_19570,N_19281);
and UO_1177 (O_1177,N_19516,N_19694);
xor UO_1178 (O_1178,N_19624,N_19683);
and UO_1179 (O_1179,N_19369,N_19338);
nand UO_1180 (O_1180,N_19890,N_19225);
nand UO_1181 (O_1181,N_19987,N_19613);
and UO_1182 (O_1182,N_19656,N_19662);
xor UO_1183 (O_1183,N_19411,N_19663);
nor UO_1184 (O_1184,N_19564,N_19242);
or UO_1185 (O_1185,N_19859,N_19789);
nand UO_1186 (O_1186,N_19917,N_19796);
nand UO_1187 (O_1187,N_19887,N_19840);
or UO_1188 (O_1188,N_19663,N_19799);
or UO_1189 (O_1189,N_19471,N_19732);
or UO_1190 (O_1190,N_19658,N_19647);
nor UO_1191 (O_1191,N_19876,N_19516);
or UO_1192 (O_1192,N_19669,N_19551);
and UO_1193 (O_1193,N_19525,N_19526);
or UO_1194 (O_1194,N_19864,N_19233);
nand UO_1195 (O_1195,N_19437,N_19742);
nand UO_1196 (O_1196,N_19600,N_19532);
xor UO_1197 (O_1197,N_19932,N_19308);
nand UO_1198 (O_1198,N_19803,N_19502);
nand UO_1199 (O_1199,N_19618,N_19565);
or UO_1200 (O_1200,N_19809,N_19975);
nand UO_1201 (O_1201,N_19871,N_19818);
xor UO_1202 (O_1202,N_19474,N_19681);
nor UO_1203 (O_1203,N_19741,N_19737);
or UO_1204 (O_1204,N_19525,N_19541);
nand UO_1205 (O_1205,N_19799,N_19286);
xnor UO_1206 (O_1206,N_19248,N_19719);
and UO_1207 (O_1207,N_19756,N_19889);
xnor UO_1208 (O_1208,N_19446,N_19502);
nor UO_1209 (O_1209,N_19644,N_19342);
nand UO_1210 (O_1210,N_19740,N_19254);
nor UO_1211 (O_1211,N_19398,N_19629);
or UO_1212 (O_1212,N_19755,N_19481);
nor UO_1213 (O_1213,N_19218,N_19638);
nand UO_1214 (O_1214,N_19255,N_19384);
and UO_1215 (O_1215,N_19689,N_19722);
nor UO_1216 (O_1216,N_19975,N_19741);
and UO_1217 (O_1217,N_19773,N_19583);
or UO_1218 (O_1218,N_19778,N_19942);
and UO_1219 (O_1219,N_19443,N_19341);
and UO_1220 (O_1220,N_19588,N_19713);
nand UO_1221 (O_1221,N_19519,N_19207);
and UO_1222 (O_1222,N_19683,N_19301);
nand UO_1223 (O_1223,N_19251,N_19381);
nor UO_1224 (O_1224,N_19218,N_19991);
and UO_1225 (O_1225,N_19640,N_19406);
nand UO_1226 (O_1226,N_19919,N_19819);
nor UO_1227 (O_1227,N_19450,N_19813);
xnor UO_1228 (O_1228,N_19432,N_19788);
nand UO_1229 (O_1229,N_19389,N_19554);
xnor UO_1230 (O_1230,N_19669,N_19316);
xnor UO_1231 (O_1231,N_19641,N_19351);
xnor UO_1232 (O_1232,N_19432,N_19562);
xor UO_1233 (O_1233,N_19966,N_19557);
nand UO_1234 (O_1234,N_19962,N_19267);
or UO_1235 (O_1235,N_19718,N_19548);
or UO_1236 (O_1236,N_19903,N_19820);
or UO_1237 (O_1237,N_19888,N_19695);
nor UO_1238 (O_1238,N_19819,N_19390);
nor UO_1239 (O_1239,N_19971,N_19505);
and UO_1240 (O_1240,N_19859,N_19496);
nor UO_1241 (O_1241,N_19428,N_19976);
nand UO_1242 (O_1242,N_19914,N_19248);
xnor UO_1243 (O_1243,N_19515,N_19779);
xnor UO_1244 (O_1244,N_19206,N_19519);
xor UO_1245 (O_1245,N_19259,N_19891);
nor UO_1246 (O_1246,N_19805,N_19257);
or UO_1247 (O_1247,N_19604,N_19914);
nor UO_1248 (O_1248,N_19537,N_19940);
and UO_1249 (O_1249,N_19379,N_19642);
nand UO_1250 (O_1250,N_19299,N_19441);
nand UO_1251 (O_1251,N_19255,N_19582);
nor UO_1252 (O_1252,N_19674,N_19321);
nand UO_1253 (O_1253,N_19844,N_19780);
nand UO_1254 (O_1254,N_19585,N_19365);
xnor UO_1255 (O_1255,N_19944,N_19480);
nand UO_1256 (O_1256,N_19759,N_19669);
xor UO_1257 (O_1257,N_19895,N_19992);
xor UO_1258 (O_1258,N_19270,N_19303);
xnor UO_1259 (O_1259,N_19976,N_19406);
or UO_1260 (O_1260,N_19454,N_19536);
or UO_1261 (O_1261,N_19416,N_19301);
or UO_1262 (O_1262,N_19294,N_19600);
nor UO_1263 (O_1263,N_19575,N_19304);
nor UO_1264 (O_1264,N_19987,N_19681);
nand UO_1265 (O_1265,N_19792,N_19324);
nand UO_1266 (O_1266,N_19457,N_19941);
and UO_1267 (O_1267,N_19714,N_19934);
and UO_1268 (O_1268,N_19550,N_19256);
xor UO_1269 (O_1269,N_19774,N_19841);
and UO_1270 (O_1270,N_19212,N_19661);
and UO_1271 (O_1271,N_19569,N_19527);
xnor UO_1272 (O_1272,N_19409,N_19760);
or UO_1273 (O_1273,N_19934,N_19520);
or UO_1274 (O_1274,N_19310,N_19865);
and UO_1275 (O_1275,N_19860,N_19444);
nand UO_1276 (O_1276,N_19734,N_19865);
nor UO_1277 (O_1277,N_19694,N_19618);
or UO_1278 (O_1278,N_19231,N_19831);
or UO_1279 (O_1279,N_19583,N_19690);
nand UO_1280 (O_1280,N_19756,N_19818);
and UO_1281 (O_1281,N_19610,N_19501);
xor UO_1282 (O_1282,N_19294,N_19610);
or UO_1283 (O_1283,N_19504,N_19400);
nor UO_1284 (O_1284,N_19404,N_19451);
xnor UO_1285 (O_1285,N_19592,N_19445);
xnor UO_1286 (O_1286,N_19807,N_19979);
xor UO_1287 (O_1287,N_19874,N_19676);
xor UO_1288 (O_1288,N_19295,N_19851);
xnor UO_1289 (O_1289,N_19816,N_19595);
and UO_1290 (O_1290,N_19555,N_19280);
nor UO_1291 (O_1291,N_19814,N_19673);
nand UO_1292 (O_1292,N_19564,N_19206);
and UO_1293 (O_1293,N_19759,N_19522);
nor UO_1294 (O_1294,N_19766,N_19317);
nor UO_1295 (O_1295,N_19904,N_19245);
nor UO_1296 (O_1296,N_19320,N_19537);
nand UO_1297 (O_1297,N_19222,N_19939);
nor UO_1298 (O_1298,N_19437,N_19752);
nor UO_1299 (O_1299,N_19307,N_19477);
or UO_1300 (O_1300,N_19960,N_19410);
xor UO_1301 (O_1301,N_19804,N_19915);
and UO_1302 (O_1302,N_19721,N_19537);
nor UO_1303 (O_1303,N_19381,N_19797);
nand UO_1304 (O_1304,N_19250,N_19322);
and UO_1305 (O_1305,N_19315,N_19403);
or UO_1306 (O_1306,N_19312,N_19995);
and UO_1307 (O_1307,N_19720,N_19217);
and UO_1308 (O_1308,N_19440,N_19821);
nor UO_1309 (O_1309,N_19411,N_19343);
nand UO_1310 (O_1310,N_19473,N_19340);
nand UO_1311 (O_1311,N_19355,N_19784);
xor UO_1312 (O_1312,N_19362,N_19955);
nand UO_1313 (O_1313,N_19610,N_19975);
or UO_1314 (O_1314,N_19835,N_19404);
xor UO_1315 (O_1315,N_19294,N_19316);
or UO_1316 (O_1316,N_19496,N_19697);
and UO_1317 (O_1317,N_19882,N_19229);
nor UO_1318 (O_1318,N_19289,N_19935);
xnor UO_1319 (O_1319,N_19213,N_19586);
nand UO_1320 (O_1320,N_19888,N_19794);
and UO_1321 (O_1321,N_19492,N_19359);
or UO_1322 (O_1322,N_19619,N_19769);
and UO_1323 (O_1323,N_19476,N_19264);
nor UO_1324 (O_1324,N_19832,N_19715);
nand UO_1325 (O_1325,N_19864,N_19214);
or UO_1326 (O_1326,N_19316,N_19791);
xnor UO_1327 (O_1327,N_19527,N_19835);
or UO_1328 (O_1328,N_19559,N_19907);
nand UO_1329 (O_1329,N_19958,N_19625);
xor UO_1330 (O_1330,N_19653,N_19741);
nand UO_1331 (O_1331,N_19898,N_19871);
and UO_1332 (O_1332,N_19758,N_19807);
nand UO_1333 (O_1333,N_19552,N_19551);
xor UO_1334 (O_1334,N_19944,N_19240);
xor UO_1335 (O_1335,N_19801,N_19680);
or UO_1336 (O_1336,N_19270,N_19758);
nor UO_1337 (O_1337,N_19229,N_19711);
nor UO_1338 (O_1338,N_19751,N_19348);
nand UO_1339 (O_1339,N_19637,N_19509);
xor UO_1340 (O_1340,N_19763,N_19638);
and UO_1341 (O_1341,N_19334,N_19590);
or UO_1342 (O_1342,N_19505,N_19357);
or UO_1343 (O_1343,N_19263,N_19694);
nand UO_1344 (O_1344,N_19699,N_19944);
nand UO_1345 (O_1345,N_19204,N_19891);
and UO_1346 (O_1346,N_19383,N_19219);
nand UO_1347 (O_1347,N_19611,N_19568);
nand UO_1348 (O_1348,N_19383,N_19986);
nor UO_1349 (O_1349,N_19512,N_19540);
or UO_1350 (O_1350,N_19323,N_19670);
nor UO_1351 (O_1351,N_19568,N_19711);
xor UO_1352 (O_1352,N_19782,N_19702);
or UO_1353 (O_1353,N_19315,N_19718);
or UO_1354 (O_1354,N_19956,N_19773);
or UO_1355 (O_1355,N_19480,N_19687);
or UO_1356 (O_1356,N_19657,N_19882);
xnor UO_1357 (O_1357,N_19687,N_19720);
xor UO_1358 (O_1358,N_19923,N_19449);
nand UO_1359 (O_1359,N_19237,N_19890);
xor UO_1360 (O_1360,N_19355,N_19970);
nor UO_1361 (O_1361,N_19829,N_19909);
xor UO_1362 (O_1362,N_19849,N_19460);
and UO_1363 (O_1363,N_19414,N_19526);
or UO_1364 (O_1364,N_19359,N_19627);
nor UO_1365 (O_1365,N_19228,N_19355);
or UO_1366 (O_1366,N_19641,N_19285);
nand UO_1367 (O_1367,N_19734,N_19283);
and UO_1368 (O_1368,N_19838,N_19457);
nand UO_1369 (O_1369,N_19338,N_19832);
nand UO_1370 (O_1370,N_19475,N_19776);
xnor UO_1371 (O_1371,N_19439,N_19595);
nor UO_1372 (O_1372,N_19573,N_19433);
or UO_1373 (O_1373,N_19935,N_19660);
nor UO_1374 (O_1374,N_19542,N_19821);
xnor UO_1375 (O_1375,N_19952,N_19808);
and UO_1376 (O_1376,N_19766,N_19557);
and UO_1377 (O_1377,N_19525,N_19775);
or UO_1378 (O_1378,N_19330,N_19628);
and UO_1379 (O_1379,N_19306,N_19841);
nor UO_1380 (O_1380,N_19493,N_19264);
nor UO_1381 (O_1381,N_19934,N_19595);
xor UO_1382 (O_1382,N_19828,N_19343);
nor UO_1383 (O_1383,N_19464,N_19225);
nand UO_1384 (O_1384,N_19822,N_19483);
or UO_1385 (O_1385,N_19734,N_19281);
nor UO_1386 (O_1386,N_19621,N_19908);
or UO_1387 (O_1387,N_19417,N_19825);
xnor UO_1388 (O_1388,N_19360,N_19954);
xnor UO_1389 (O_1389,N_19629,N_19477);
or UO_1390 (O_1390,N_19838,N_19291);
xor UO_1391 (O_1391,N_19238,N_19280);
nor UO_1392 (O_1392,N_19889,N_19637);
or UO_1393 (O_1393,N_19949,N_19742);
xor UO_1394 (O_1394,N_19712,N_19686);
or UO_1395 (O_1395,N_19842,N_19820);
or UO_1396 (O_1396,N_19876,N_19589);
or UO_1397 (O_1397,N_19758,N_19442);
and UO_1398 (O_1398,N_19361,N_19472);
and UO_1399 (O_1399,N_19975,N_19587);
nand UO_1400 (O_1400,N_19321,N_19907);
and UO_1401 (O_1401,N_19989,N_19222);
nor UO_1402 (O_1402,N_19644,N_19274);
nand UO_1403 (O_1403,N_19415,N_19810);
nand UO_1404 (O_1404,N_19858,N_19681);
xnor UO_1405 (O_1405,N_19945,N_19309);
or UO_1406 (O_1406,N_19897,N_19722);
nor UO_1407 (O_1407,N_19883,N_19937);
nor UO_1408 (O_1408,N_19209,N_19219);
nor UO_1409 (O_1409,N_19570,N_19306);
nor UO_1410 (O_1410,N_19948,N_19775);
nor UO_1411 (O_1411,N_19228,N_19265);
and UO_1412 (O_1412,N_19358,N_19596);
and UO_1413 (O_1413,N_19633,N_19526);
xnor UO_1414 (O_1414,N_19433,N_19689);
and UO_1415 (O_1415,N_19447,N_19995);
nand UO_1416 (O_1416,N_19814,N_19232);
and UO_1417 (O_1417,N_19267,N_19640);
or UO_1418 (O_1418,N_19747,N_19631);
or UO_1419 (O_1419,N_19204,N_19325);
and UO_1420 (O_1420,N_19701,N_19473);
or UO_1421 (O_1421,N_19830,N_19354);
xnor UO_1422 (O_1422,N_19922,N_19819);
and UO_1423 (O_1423,N_19430,N_19584);
nand UO_1424 (O_1424,N_19759,N_19791);
and UO_1425 (O_1425,N_19747,N_19356);
nor UO_1426 (O_1426,N_19348,N_19996);
or UO_1427 (O_1427,N_19805,N_19789);
or UO_1428 (O_1428,N_19431,N_19323);
nand UO_1429 (O_1429,N_19769,N_19438);
or UO_1430 (O_1430,N_19948,N_19498);
nand UO_1431 (O_1431,N_19776,N_19465);
and UO_1432 (O_1432,N_19795,N_19889);
and UO_1433 (O_1433,N_19877,N_19467);
nand UO_1434 (O_1434,N_19752,N_19654);
nor UO_1435 (O_1435,N_19800,N_19400);
xnor UO_1436 (O_1436,N_19980,N_19857);
xor UO_1437 (O_1437,N_19462,N_19213);
or UO_1438 (O_1438,N_19314,N_19974);
or UO_1439 (O_1439,N_19906,N_19658);
nand UO_1440 (O_1440,N_19574,N_19209);
xor UO_1441 (O_1441,N_19262,N_19263);
xor UO_1442 (O_1442,N_19591,N_19867);
nor UO_1443 (O_1443,N_19544,N_19949);
nor UO_1444 (O_1444,N_19909,N_19719);
nor UO_1445 (O_1445,N_19553,N_19530);
nand UO_1446 (O_1446,N_19636,N_19651);
or UO_1447 (O_1447,N_19572,N_19962);
xor UO_1448 (O_1448,N_19531,N_19434);
nand UO_1449 (O_1449,N_19683,N_19448);
and UO_1450 (O_1450,N_19648,N_19818);
xor UO_1451 (O_1451,N_19810,N_19309);
xnor UO_1452 (O_1452,N_19867,N_19737);
nand UO_1453 (O_1453,N_19289,N_19565);
or UO_1454 (O_1454,N_19325,N_19660);
and UO_1455 (O_1455,N_19927,N_19518);
xor UO_1456 (O_1456,N_19306,N_19299);
or UO_1457 (O_1457,N_19350,N_19802);
nand UO_1458 (O_1458,N_19642,N_19876);
xnor UO_1459 (O_1459,N_19388,N_19313);
and UO_1460 (O_1460,N_19658,N_19948);
xor UO_1461 (O_1461,N_19782,N_19384);
nand UO_1462 (O_1462,N_19645,N_19894);
and UO_1463 (O_1463,N_19592,N_19365);
xor UO_1464 (O_1464,N_19415,N_19766);
nor UO_1465 (O_1465,N_19485,N_19468);
and UO_1466 (O_1466,N_19317,N_19513);
xnor UO_1467 (O_1467,N_19947,N_19346);
nand UO_1468 (O_1468,N_19457,N_19225);
and UO_1469 (O_1469,N_19242,N_19420);
nand UO_1470 (O_1470,N_19406,N_19593);
nand UO_1471 (O_1471,N_19846,N_19272);
xor UO_1472 (O_1472,N_19470,N_19690);
or UO_1473 (O_1473,N_19633,N_19398);
xnor UO_1474 (O_1474,N_19753,N_19587);
or UO_1475 (O_1475,N_19954,N_19813);
nor UO_1476 (O_1476,N_19265,N_19813);
nand UO_1477 (O_1477,N_19439,N_19645);
nand UO_1478 (O_1478,N_19944,N_19792);
and UO_1479 (O_1479,N_19463,N_19948);
and UO_1480 (O_1480,N_19574,N_19825);
xor UO_1481 (O_1481,N_19278,N_19734);
nand UO_1482 (O_1482,N_19526,N_19748);
nand UO_1483 (O_1483,N_19680,N_19861);
nand UO_1484 (O_1484,N_19746,N_19494);
nor UO_1485 (O_1485,N_19322,N_19663);
and UO_1486 (O_1486,N_19394,N_19937);
nor UO_1487 (O_1487,N_19507,N_19319);
nor UO_1488 (O_1488,N_19666,N_19625);
or UO_1489 (O_1489,N_19936,N_19217);
xor UO_1490 (O_1490,N_19380,N_19906);
or UO_1491 (O_1491,N_19318,N_19224);
nor UO_1492 (O_1492,N_19743,N_19333);
and UO_1493 (O_1493,N_19881,N_19931);
or UO_1494 (O_1494,N_19575,N_19682);
and UO_1495 (O_1495,N_19787,N_19251);
nand UO_1496 (O_1496,N_19265,N_19216);
nand UO_1497 (O_1497,N_19973,N_19553);
nor UO_1498 (O_1498,N_19540,N_19914);
or UO_1499 (O_1499,N_19887,N_19229);
nand UO_1500 (O_1500,N_19892,N_19919);
nor UO_1501 (O_1501,N_19687,N_19440);
and UO_1502 (O_1502,N_19221,N_19389);
xnor UO_1503 (O_1503,N_19763,N_19857);
nor UO_1504 (O_1504,N_19420,N_19390);
or UO_1505 (O_1505,N_19668,N_19354);
nor UO_1506 (O_1506,N_19203,N_19654);
nand UO_1507 (O_1507,N_19212,N_19955);
or UO_1508 (O_1508,N_19808,N_19987);
nor UO_1509 (O_1509,N_19761,N_19692);
nand UO_1510 (O_1510,N_19381,N_19713);
nor UO_1511 (O_1511,N_19821,N_19212);
xor UO_1512 (O_1512,N_19218,N_19622);
or UO_1513 (O_1513,N_19892,N_19206);
nand UO_1514 (O_1514,N_19737,N_19717);
or UO_1515 (O_1515,N_19984,N_19828);
nand UO_1516 (O_1516,N_19962,N_19797);
or UO_1517 (O_1517,N_19927,N_19359);
and UO_1518 (O_1518,N_19524,N_19506);
or UO_1519 (O_1519,N_19469,N_19514);
nor UO_1520 (O_1520,N_19863,N_19580);
nand UO_1521 (O_1521,N_19586,N_19825);
nand UO_1522 (O_1522,N_19354,N_19602);
and UO_1523 (O_1523,N_19260,N_19446);
or UO_1524 (O_1524,N_19868,N_19796);
and UO_1525 (O_1525,N_19712,N_19245);
nor UO_1526 (O_1526,N_19220,N_19394);
nor UO_1527 (O_1527,N_19641,N_19472);
or UO_1528 (O_1528,N_19352,N_19482);
or UO_1529 (O_1529,N_19612,N_19458);
xnor UO_1530 (O_1530,N_19999,N_19206);
xnor UO_1531 (O_1531,N_19544,N_19334);
nor UO_1532 (O_1532,N_19246,N_19947);
nand UO_1533 (O_1533,N_19567,N_19914);
xor UO_1534 (O_1534,N_19975,N_19660);
nor UO_1535 (O_1535,N_19952,N_19310);
and UO_1536 (O_1536,N_19529,N_19628);
nor UO_1537 (O_1537,N_19291,N_19356);
and UO_1538 (O_1538,N_19359,N_19355);
or UO_1539 (O_1539,N_19452,N_19489);
nand UO_1540 (O_1540,N_19943,N_19441);
nor UO_1541 (O_1541,N_19713,N_19614);
nor UO_1542 (O_1542,N_19632,N_19665);
nor UO_1543 (O_1543,N_19694,N_19870);
xor UO_1544 (O_1544,N_19654,N_19213);
xnor UO_1545 (O_1545,N_19320,N_19519);
xor UO_1546 (O_1546,N_19448,N_19960);
nand UO_1547 (O_1547,N_19749,N_19597);
and UO_1548 (O_1548,N_19595,N_19807);
and UO_1549 (O_1549,N_19881,N_19648);
nand UO_1550 (O_1550,N_19670,N_19229);
and UO_1551 (O_1551,N_19790,N_19717);
nor UO_1552 (O_1552,N_19757,N_19432);
and UO_1553 (O_1553,N_19630,N_19845);
or UO_1554 (O_1554,N_19688,N_19787);
nand UO_1555 (O_1555,N_19375,N_19294);
or UO_1556 (O_1556,N_19595,N_19279);
and UO_1557 (O_1557,N_19550,N_19870);
or UO_1558 (O_1558,N_19673,N_19396);
xnor UO_1559 (O_1559,N_19361,N_19489);
nor UO_1560 (O_1560,N_19592,N_19232);
and UO_1561 (O_1561,N_19951,N_19447);
and UO_1562 (O_1562,N_19748,N_19717);
or UO_1563 (O_1563,N_19856,N_19864);
or UO_1564 (O_1564,N_19592,N_19722);
and UO_1565 (O_1565,N_19432,N_19758);
xor UO_1566 (O_1566,N_19993,N_19742);
nor UO_1567 (O_1567,N_19700,N_19848);
and UO_1568 (O_1568,N_19938,N_19792);
xor UO_1569 (O_1569,N_19846,N_19677);
nand UO_1570 (O_1570,N_19501,N_19278);
or UO_1571 (O_1571,N_19908,N_19980);
xnor UO_1572 (O_1572,N_19302,N_19603);
or UO_1573 (O_1573,N_19868,N_19598);
nand UO_1574 (O_1574,N_19799,N_19398);
nor UO_1575 (O_1575,N_19865,N_19562);
xnor UO_1576 (O_1576,N_19881,N_19993);
or UO_1577 (O_1577,N_19666,N_19305);
nand UO_1578 (O_1578,N_19660,N_19918);
or UO_1579 (O_1579,N_19489,N_19632);
or UO_1580 (O_1580,N_19975,N_19500);
or UO_1581 (O_1581,N_19425,N_19717);
and UO_1582 (O_1582,N_19577,N_19868);
nor UO_1583 (O_1583,N_19527,N_19546);
nand UO_1584 (O_1584,N_19424,N_19726);
nor UO_1585 (O_1585,N_19804,N_19410);
xor UO_1586 (O_1586,N_19233,N_19894);
and UO_1587 (O_1587,N_19994,N_19672);
nand UO_1588 (O_1588,N_19976,N_19827);
or UO_1589 (O_1589,N_19379,N_19462);
or UO_1590 (O_1590,N_19977,N_19441);
xor UO_1591 (O_1591,N_19306,N_19372);
nand UO_1592 (O_1592,N_19213,N_19604);
xnor UO_1593 (O_1593,N_19403,N_19474);
xnor UO_1594 (O_1594,N_19468,N_19709);
or UO_1595 (O_1595,N_19306,N_19216);
nand UO_1596 (O_1596,N_19250,N_19868);
and UO_1597 (O_1597,N_19480,N_19344);
xnor UO_1598 (O_1598,N_19980,N_19389);
and UO_1599 (O_1599,N_19777,N_19566);
nand UO_1600 (O_1600,N_19826,N_19492);
xnor UO_1601 (O_1601,N_19682,N_19490);
or UO_1602 (O_1602,N_19795,N_19552);
nand UO_1603 (O_1603,N_19818,N_19319);
and UO_1604 (O_1604,N_19546,N_19653);
or UO_1605 (O_1605,N_19370,N_19325);
or UO_1606 (O_1606,N_19381,N_19538);
and UO_1607 (O_1607,N_19307,N_19312);
nand UO_1608 (O_1608,N_19274,N_19725);
nand UO_1609 (O_1609,N_19521,N_19641);
or UO_1610 (O_1610,N_19201,N_19843);
nor UO_1611 (O_1611,N_19279,N_19470);
nand UO_1612 (O_1612,N_19312,N_19936);
nand UO_1613 (O_1613,N_19671,N_19427);
and UO_1614 (O_1614,N_19625,N_19561);
nor UO_1615 (O_1615,N_19694,N_19439);
nand UO_1616 (O_1616,N_19960,N_19824);
xor UO_1617 (O_1617,N_19703,N_19988);
nand UO_1618 (O_1618,N_19584,N_19628);
or UO_1619 (O_1619,N_19256,N_19605);
and UO_1620 (O_1620,N_19273,N_19297);
nor UO_1621 (O_1621,N_19933,N_19892);
or UO_1622 (O_1622,N_19799,N_19301);
nand UO_1623 (O_1623,N_19457,N_19891);
or UO_1624 (O_1624,N_19307,N_19677);
xor UO_1625 (O_1625,N_19585,N_19703);
xnor UO_1626 (O_1626,N_19816,N_19965);
and UO_1627 (O_1627,N_19556,N_19791);
xnor UO_1628 (O_1628,N_19850,N_19499);
nor UO_1629 (O_1629,N_19677,N_19544);
xor UO_1630 (O_1630,N_19533,N_19365);
xor UO_1631 (O_1631,N_19808,N_19803);
xnor UO_1632 (O_1632,N_19793,N_19585);
nor UO_1633 (O_1633,N_19908,N_19792);
nor UO_1634 (O_1634,N_19215,N_19233);
or UO_1635 (O_1635,N_19876,N_19925);
and UO_1636 (O_1636,N_19204,N_19476);
xor UO_1637 (O_1637,N_19597,N_19860);
or UO_1638 (O_1638,N_19230,N_19409);
xnor UO_1639 (O_1639,N_19638,N_19698);
xor UO_1640 (O_1640,N_19568,N_19664);
and UO_1641 (O_1641,N_19705,N_19516);
nand UO_1642 (O_1642,N_19555,N_19731);
or UO_1643 (O_1643,N_19747,N_19485);
or UO_1644 (O_1644,N_19483,N_19707);
nor UO_1645 (O_1645,N_19731,N_19260);
xnor UO_1646 (O_1646,N_19402,N_19888);
xnor UO_1647 (O_1647,N_19646,N_19700);
or UO_1648 (O_1648,N_19520,N_19762);
nand UO_1649 (O_1649,N_19488,N_19386);
and UO_1650 (O_1650,N_19881,N_19863);
nor UO_1651 (O_1651,N_19715,N_19538);
nor UO_1652 (O_1652,N_19515,N_19523);
nand UO_1653 (O_1653,N_19477,N_19323);
nor UO_1654 (O_1654,N_19402,N_19365);
xnor UO_1655 (O_1655,N_19548,N_19829);
xnor UO_1656 (O_1656,N_19400,N_19314);
nand UO_1657 (O_1657,N_19942,N_19884);
and UO_1658 (O_1658,N_19950,N_19611);
nor UO_1659 (O_1659,N_19686,N_19543);
or UO_1660 (O_1660,N_19341,N_19610);
nor UO_1661 (O_1661,N_19487,N_19953);
and UO_1662 (O_1662,N_19646,N_19790);
nand UO_1663 (O_1663,N_19633,N_19219);
xnor UO_1664 (O_1664,N_19274,N_19802);
nor UO_1665 (O_1665,N_19282,N_19740);
nor UO_1666 (O_1666,N_19703,N_19385);
xor UO_1667 (O_1667,N_19549,N_19821);
xor UO_1668 (O_1668,N_19279,N_19482);
nand UO_1669 (O_1669,N_19908,N_19610);
or UO_1670 (O_1670,N_19498,N_19679);
nor UO_1671 (O_1671,N_19275,N_19594);
and UO_1672 (O_1672,N_19344,N_19461);
and UO_1673 (O_1673,N_19855,N_19841);
nand UO_1674 (O_1674,N_19455,N_19460);
xnor UO_1675 (O_1675,N_19752,N_19541);
xnor UO_1676 (O_1676,N_19852,N_19406);
xor UO_1677 (O_1677,N_19756,N_19445);
nand UO_1678 (O_1678,N_19371,N_19236);
xor UO_1679 (O_1679,N_19409,N_19614);
or UO_1680 (O_1680,N_19657,N_19417);
nor UO_1681 (O_1681,N_19585,N_19677);
nor UO_1682 (O_1682,N_19541,N_19764);
nand UO_1683 (O_1683,N_19451,N_19251);
and UO_1684 (O_1684,N_19350,N_19907);
nor UO_1685 (O_1685,N_19999,N_19876);
or UO_1686 (O_1686,N_19411,N_19472);
nand UO_1687 (O_1687,N_19532,N_19390);
nand UO_1688 (O_1688,N_19845,N_19273);
and UO_1689 (O_1689,N_19584,N_19311);
nand UO_1690 (O_1690,N_19908,N_19525);
or UO_1691 (O_1691,N_19559,N_19339);
and UO_1692 (O_1692,N_19482,N_19829);
nor UO_1693 (O_1693,N_19936,N_19778);
xnor UO_1694 (O_1694,N_19390,N_19615);
or UO_1695 (O_1695,N_19394,N_19467);
nor UO_1696 (O_1696,N_19206,N_19907);
xor UO_1697 (O_1697,N_19972,N_19298);
nand UO_1698 (O_1698,N_19378,N_19869);
nor UO_1699 (O_1699,N_19462,N_19243);
or UO_1700 (O_1700,N_19668,N_19556);
or UO_1701 (O_1701,N_19888,N_19376);
or UO_1702 (O_1702,N_19542,N_19409);
nor UO_1703 (O_1703,N_19676,N_19579);
xnor UO_1704 (O_1704,N_19456,N_19426);
or UO_1705 (O_1705,N_19441,N_19672);
nor UO_1706 (O_1706,N_19804,N_19355);
and UO_1707 (O_1707,N_19635,N_19830);
xor UO_1708 (O_1708,N_19404,N_19887);
nand UO_1709 (O_1709,N_19399,N_19569);
nor UO_1710 (O_1710,N_19392,N_19744);
and UO_1711 (O_1711,N_19851,N_19286);
xor UO_1712 (O_1712,N_19555,N_19766);
nand UO_1713 (O_1713,N_19992,N_19675);
or UO_1714 (O_1714,N_19940,N_19457);
or UO_1715 (O_1715,N_19694,N_19286);
xor UO_1716 (O_1716,N_19771,N_19490);
xor UO_1717 (O_1717,N_19480,N_19503);
or UO_1718 (O_1718,N_19496,N_19655);
and UO_1719 (O_1719,N_19832,N_19255);
and UO_1720 (O_1720,N_19263,N_19683);
or UO_1721 (O_1721,N_19763,N_19510);
xor UO_1722 (O_1722,N_19620,N_19290);
xor UO_1723 (O_1723,N_19225,N_19294);
nand UO_1724 (O_1724,N_19954,N_19850);
and UO_1725 (O_1725,N_19535,N_19730);
nor UO_1726 (O_1726,N_19233,N_19481);
nand UO_1727 (O_1727,N_19958,N_19863);
nor UO_1728 (O_1728,N_19682,N_19571);
xor UO_1729 (O_1729,N_19786,N_19778);
xnor UO_1730 (O_1730,N_19974,N_19517);
xor UO_1731 (O_1731,N_19244,N_19344);
nor UO_1732 (O_1732,N_19277,N_19358);
xor UO_1733 (O_1733,N_19247,N_19855);
xor UO_1734 (O_1734,N_19604,N_19257);
and UO_1735 (O_1735,N_19387,N_19434);
nand UO_1736 (O_1736,N_19985,N_19296);
and UO_1737 (O_1737,N_19810,N_19930);
and UO_1738 (O_1738,N_19491,N_19621);
nor UO_1739 (O_1739,N_19580,N_19374);
nand UO_1740 (O_1740,N_19898,N_19727);
and UO_1741 (O_1741,N_19747,N_19983);
or UO_1742 (O_1742,N_19478,N_19862);
and UO_1743 (O_1743,N_19332,N_19805);
nor UO_1744 (O_1744,N_19527,N_19345);
and UO_1745 (O_1745,N_19237,N_19620);
or UO_1746 (O_1746,N_19315,N_19705);
and UO_1747 (O_1747,N_19757,N_19833);
xor UO_1748 (O_1748,N_19260,N_19263);
xnor UO_1749 (O_1749,N_19474,N_19654);
or UO_1750 (O_1750,N_19861,N_19732);
or UO_1751 (O_1751,N_19586,N_19532);
xor UO_1752 (O_1752,N_19262,N_19763);
nor UO_1753 (O_1753,N_19916,N_19684);
nand UO_1754 (O_1754,N_19758,N_19936);
and UO_1755 (O_1755,N_19242,N_19447);
nor UO_1756 (O_1756,N_19487,N_19875);
and UO_1757 (O_1757,N_19423,N_19835);
nor UO_1758 (O_1758,N_19448,N_19416);
nor UO_1759 (O_1759,N_19597,N_19262);
and UO_1760 (O_1760,N_19996,N_19973);
or UO_1761 (O_1761,N_19944,N_19894);
nor UO_1762 (O_1762,N_19271,N_19357);
nor UO_1763 (O_1763,N_19579,N_19699);
and UO_1764 (O_1764,N_19901,N_19401);
and UO_1765 (O_1765,N_19271,N_19966);
nand UO_1766 (O_1766,N_19379,N_19926);
or UO_1767 (O_1767,N_19782,N_19568);
or UO_1768 (O_1768,N_19621,N_19794);
xnor UO_1769 (O_1769,N_19580,N_19246);
nor UO_1770 (O_1770,N_19555,N_19786);
nand UO_1771 (O_1771,N_19426,N_19364);
nor UO_1772 (O_1772,N_19837,N_19843);
or UO_1773 (O_1773,N_19424,N_19614);
nand UO_1774 (O_1774,N_19330,N_19612);
or UO_1775 (O_1775,N_19919,N_19978);
nand UO_1776 (O_1776,N_19419,N_19230);
xor UO_1777 (O_1777,N_19961,N_19832);
xor UO_1778 (O_1778,N_19910,N_19718);
or UO_1779 (O_1779,N_19555,N_19432);
nor UO_1780 (O_1780,N_19229,N_19444);
or UO_1781 (O_1781,N_19995,N_19701);
or UO_1782 (O_1782,N_19231,N_19379);
xnor UO_1783 (O_1783,N_19910,N_19515);
xnor UO_1784 (O_1784,N_19624,N_19708);
and UO_1785 (O_1785,N_19370,N_19484);
and UO_1786 (O_1786,N_19210,N_19553);
and UO_1787 (O_1787,N_19955,N_19924);
xnor UO_1788 (O_1788,N_19889,N_19451);
xnor UO_1789 (O_1789,N_19657,N_19467);
xnor UO_1790 (O_1790,N_19249,N_19213);
or UO_1791 (O_1791,N_19563,N_19599);
or UO_1792 (O_1792,N_19822,N_19354);
nor UO_1793 (O_1793,N_19436,N_19569);
or UO_1794 (O_1794,N_19219,N_19218);
nand UO_1795 (O_1795,N_19245,N_19776);
or UO_1796 (O_1796,N_19640,N_19215);
xor UO_1797 (O_1797,N_19846,N_19570);
nor UO_1798 (O_1798,N_19331,N_19451);
xnor UO_1799 (O_1799,N_19578,N_19749);
and UO_1800 (O_1800,N_19375,N_19865);
nor UO_1801 (O_1801,N_19951,N_19344);
or UO_1802 (O_1802,N_19334,N_19765);
xnor UO_1803 (O_1803,N_19695,N_19351);
xnor UO_1804 (O_1804,N_19230,N_19250);
xor UO_1805 (O_1805,N_19368,N_19795);
or UO_1806 (O_1806,N_19486,N_19452);
nand UO_1807 (O_1807,N_19663,N_19563);
and UO_1808 (O_1808,N_19402,N_19652);
xor UO_1809 (O_1809,N_19380,N_19462);
and UO_1810 (O_1810,N_19618,N_19850);
or UO_1811 (O_1811,N_19862,N_19287);
nor UO_1812 (O_1812,N_19863,N_19310);
nand UO_1813 (O_1813,N_19890,N_19316);
or UO_1814 (O_1814,N_19877,N_19213);
or UO_1815 (O_1815,N_19239,N_19444);
nor UO_1816 (O_1816,N_19826,N_19850);
nand UO_1817 (O_1817,N_19894,N_19913);
nand UO_1818 (O_1818,N_19372,N_19626);
nor UO_1819 (O_1819,N_19685,N_19451);
and UO_1820 (O_1820,N_19973,N_19412);
nand UO_1821 (O_1821,N_19924,N_19376);
nand UO_1822 (O_1822,N_19697,N_19968);
and UO_1823 (O_1823,N_19991,N_19713);
nor UO_1824 (O_1824,N_19626,N_19224);
or UO_1825 (O_1825,N_19763,N_19606);
nand UO_1826 (O_1826,N_19735,N_19302);
or UO_1827 (O_1827,N_19980,N_19248);
xnor UO_1828 (O_1828,N_19321,N_19380);
nor UO_1829 (O_1829,N_19247,N_19913);
xnor UO_1830 (O_1830,N_19562,N_19684);
xnor UO_1831 (O_1831,N_19756,N_19880);
nor UO_1832 (O_1832,N_19574,N_19739);
nand UO_1833 (O_1833,N_19738,N_19838);
or UO_1834 (O_1834,N_19889,N_19701);
xnor UO_1835 (O_1835,N_19997,N_19311);
or UO_1836 (O_1836,N_19302,N_19357);
and UO_1837 (O_1837,N_19317,N_19597);
or UO_1838 (O_1838,N_19667,N_19800);
nor UO_1839 (O_1839,N_19976,N_19367);
xnor UO_1840 (O_1840,N_19850,N_19770);
nand UO_1841 (O_1841,N_19471,N_19585);
xor UO_1842 (O_1842,N_19900,N_19730);
and UO_1843 (O_1843,N_19276,N_19718);
xor UO_1844 (O_1844,N_19233,N_19484);
nand UO_1845 (O_1845,N_19669,N_19293);
xor UO_1846 (O_1846,N_19351,N_19479);
xnor UO_1847 (O_1847,N_19481,N_19805);
xnor UO_1848 (O_1848,N_19428,N_19479);
nand UO_1849 (O_1849,N_19309,N_19625);
nand UO_1850 (O_1850,N_19909,N_19793);
or UO_1851 (O_1851,N_19492,N_19814);
xnor UO_1852 (O_1852,N_19736,N_19537);
or UO_1853 (O_1853,N_19205,N_19251);
nor UO_1854 (O_1854,N_19859,N_19822);
nand UO_1855 (O_1855,N_19737,N_19340);
nand UO_1856 (O_1856,N_19283,N_19920);
or UO_1857 (O_1857,N_19453,N_19513);
and UO_1858 (O_1858,N_19702,N_19286);
nand UO_1859 (O_1859,N_19656,N_19246);
or UO_1860 (O_1860,N_19605,N_19890);
xnor UO_1861 (O_1861,N_19286,N_19527);
or UO_1862 (O_1862,N_19821,N_19927);
or UO_1863 (O_1863,N_19751,N_19269);
or UO_1864 (O_1864,N_19486,N_19215);
or UO_1865 (O_1865,N_19397,N_19592);
or UO_1866 (O_1866,N_19504,N_19561);
nand UO_1867 (O_1867,N_19956,N_19300);
nor UO_1868 (O_1868,N_19879,N_19494);
nor UO_1869 (O_1869,N_19264,N_19468);
xnor UO_1870 (O_1870,N_19905,N_19577);
nor UO_1871 (O_1871,N_19551,N_19408);
or UO_1872 (O_1872,N_19663,N_19706);
xnor UO_1873 (O_1873,N_19461,N_19320);
nand UO_1874 (O_1874,N_19325,N_19914);
xnor UO_1875 (O_1875,N_19221,N_19869);
nor UO_1876 (O_1876,N_19839,N_19846);
xnor UO_1877 (O_1877,N_19475,N_19730);
or UO_1878 (O_1878,N_19516,N_19204);
or UO_1879 (O_1879,N_19700,N_19866);
xor UO_1880 (O_1880,N_19889,N_19621);
nand UO_1881 (O_1881,N_19948,N_19861);
or UO_1882 (O_1882,N_19935,N_19801);
nand UO_1883 (O_1883,N_19597,N_19877);
nor UO_1884 (O_1884,N_19355,N_19512);
xnor UO_1885 (O_1885,N_19707,N_19540);
or UO_1886 (O_1886,N_19732,N_19812);
nand UO_1887 (O_1887,N_19975,N_19904);
xor UO_1888 (O_1888,N_19622,N_19595);
nor UO_1889 (O_1889,N_19351,N_19419);
nand UO_1890 (O_1890,N_19912,N_19216);
xor UO_1891 (O_1891,N_19236,N_19914);
and UO_1892 (O_1892,N_19537,N_19569);
xnor UO_1893 (O_1893,N_19903,N_19686);
xnor UO_1894 (O_1894,N_19234,N_19808);
xor UO_1895 (O_1895,N_19566,N_19737);
or UO_1896 (O_1896,N_19794,N_19859);
nand UO_1897 (O_1897,N_19685,N_19396);
nand UO_1898 (O_1898,N_19749,N_19629);
nand UO_1899 (O_1899,N_19647,N_19287);
nand UO_1900 (O_1900,N_19717,N_19744);
and UO_1901 (O_1901,N_19462,N_19581);
nand UO_1902 (O_1902,N_19405,N_19900);
nor UO_1903 (O_1903,N_19998,N_19504);
and UO_1904 (O_1904,N_19924,N_19931);
and UO_1905 (O_1905,N_19333,N_19797);
nand UO_1906 (O_1906,N_19703,N_19969);
or UO_1907 (O_1907,N_19770,N_19587);
and UO_1908 (O_1908,N_19207,N_19213);
nand UO_1909 (O_1909,N_19426,N_19769);
nor UO_1910 (O_1910,N_19672,N_19839);
or UO_1911 (O_1911,N_19454,N_19824);
and UO_1912 (O_1912,N_19571,N_19991);
nand UO_1913 (O_1913,N_19799,N_19372);
nand UO_1914 (O_1914,N_19955,N_19953);
nand UO_1915 (O_1915,N_19800,N_19802);
nor UO_1916 (O_1916,N_19945,N_19416);
or UO_1917 (O_1917,N_19950,N_19793);
and UO_1918 (O_1918,N_19984,N_19520);
xnor UO_1919 (O_1919,N_19403,N_19545);
xor UO_1920 (O_1920,N_19565,N_19896);
or UO_1921 (O_1921,N_19293,N_19750);
nor UO_1922 (O_1922,N_19716,N_19689);
nand UO_1923 (O_1923,N_19451,N_19730);
or UO_1924 (O_1924,N_19489,N_19701);
or UO_1925 (O_1925,N_19960,N_19765);
xnor UO_1926 (O_1926,N_19865,N_19478);
and UO_1927 (O_1927,N_19865,N_19639);
or UO_1928 (O_1928,N_19442,N_19232);
and UO_1929 (O_1929,N_19882,N_19999);
xnor UO_1930 (O_1930,N_19972,N_19471);
nor UO_1931 (O_1931,N_19787,N_19940);
nor UO_1932 (O_1932,N_19212,N_19556);
xor UO_1933 (O_1933,N_19694,N_19778);
xnor UO_1934 (O_1934,N_19672,N_19862);
nor UO_1935 (O_1935,N_19376,N_19955);
xor UO_1936 (O_1936,N_19392,N_19773);
nand UO_1937 (O_1937,N_19905,N_19289);
nor UO_1938 (O_1938,N_19464,N_19828);
and UO_1939 (O_1939,N_19523,N_19476);
and UO_1940 (O_1940,N_19332,N_19509);
or UO_1941 (O_1941,N_19726,N_19446);
nand UO_1942 (O_1942,N_19321,N_19255);
nor UO_1943 (O_1943,N_19853,N_19843);
nand UO_1944 (O_1944,N_19240,N_19767);
xor UO_1945 (O_1945,N_19364,N_19495);
nor UO_1946 (O_1946,N_19723,N_19885);
xnor UO_1947 (O_1947,N_19207,N_19399);
nand UO_1948 (O_1948,N_19556,N_19860);
nor UO_1949 (O_1949,N_19739,N_19854);
nand UO_1950 (O_1950,N_19777,N_19576);
and UO_1951 (O_1951,N_19324,N_19975);
or UO_1952 (O_1952,N_19589,N_19741);
xnor UO_1953 (O_1953,N_19680,N_19694);
nand UO_1954 (O_1954,N_19681,N_19774);
and UO_1955 (O_1955,N_19217,N_19274);
nor UO_1956 (O_1956,N_19287,N_19505);
or UO_1957 (O_1957,N_19449,N_19358);
nor UO_1958 (O_1958,N_19517,N_19629);
nor UO_1959 (O_1959,N_19490,N_19785);
nand UO_1960 (O_1960,N_19761,N_19436);
nor UO_1961 (O_1961,N_19720,N_19411);
or UO_1962 (O_1962,N_19895,N_19257);
xor UO_1963 (O_1963,N_19454,N_19749);
or UO_1964 (O_1964,N_19825,N_19957);
xor UO_1965 (O_1965,N_19952,N_19828);
or UO_1966 (O_1966,N_19527,N_19414);
or UO_1967 (O_1967,N_19335,N_19617);
nor UO_1968 (O_1968,N_19286,N_19242);
and UO_1969 (O_1969,N_19516,N_19850);
xnor UO_1970 (O_1970,N_19293,N_19304);
xnor UO_1971 (O_1971,N_19628,N_19700);
xnor UO_1972 (O_1972,N_19359,N_19467);
or UO_1973 (O_1973,N_19992,N_19728);
nor UO_1974 (O_1974,N_19256,N_19497);
nand UO_1975 (O_1975,N_19849,N_19930);
nand UO_1976 (O_1976,N_19639,N_19242);
and UO_1977 (O_1977,N_19505,N_19990);
nor UO_1978 (O_1978,N_19390,N_19990);
nor UO_1979 (O_1979,N_19244,N_19218);
nand UO_1980 (O_1980,N_19274,N_19776);
nand UO_1981 (O_1981,N_19552,N_19732);
xor UO_1982 (O_1982,N_19878,N_19823);
and UO_1983 (O_1983,N_19925,N_19345);
or UO_1984 (O_1984,N_19419,N_19200);
and UO_1985 (O_1985,N_19473,N_19789);
and UO_1986 (O_1986,N_19611,N_19956);
and UO_1987 (O_1987,N_19718,N_19463);
and UO_1988 (O_1988,N_19636,N_19262);
nand UO_1989 (O_1989,N_19230,N_19481);
nor UO_1990 (O_1990,N_19661,N_19596);
or UO_1991 (O_1991,N_19968,N_19203);
nand UO_1992 (O_1992,N_19724,N_19621);
and UO_1993 (O_1993,N_19555,N_19732);
nand UO_1994 (O_1994,N_19833,N_19997);
xor UO_1995 (O_1995,N_19857,N_19235);
and UO_1996 (O_1996,N_19488,N_19510);
nand UO_1997 (O_1997,N_19739,N_19763);
nand UO_1998 (O_1998,N_19204,N_19381);
and UO_1999 (O_1999,N_19474,N_19257);
nor UO_2000 (O_2000,N_19670,N_19932);
nand UO_2001 (O_2001,N_19200,N_19659);
and UO_2002 (O_2002,N_19745,N_19814);
nor UO_2003 (O_2003,N_19809,N_19448);
nand UO_2004 (O_2004,N_19331,N_19896);
nand UO_2005 (O_2005,N_19444,N_19602);
nor UO_2006 (O_2006,N_19220,N_19408);
xnor UO_2007 (O_2007,N_19470,N_19815);
or UO_2008 (O_2008,N_19747,N_19213);
and UO_2009 (O_2009,N_19803,N_19689);
and UO_2010 (O_2010,N_19312,N_19524);
nor UO_2011 (O_2011,N_19580,N_19871);
nand UO_2012 (O_2012,N_19433,N_19679);
or UO_2013 (O_2013,N_19501,N_19448);
nand UO_2014 (O_2014,N_19652,N_19881);
or UO_2015 (O_2015,N_19202,N_19265);
nand UO_2016 (O_2016,N_19856,N_19780);
or UO_2017 (O_2017,N_19513,N_19407);
nand UO_2018 (O_2018,N_19528,N_19829);
and UO_2019 (O_2019,N_19331,N_19498);
nand UO_2020 (O_2020,N_19278,N_19870);
xor UO_2021 (O_2021,N_19814,N_19555);
and UO_2022 (O_2022,N_19779,N_19642);
xor UO_2023 (O_2023,N_19944,N_19249);
and UO_2024 (O_2024,N_19971,N_19234);
nor UO_2025 (O_2025,N_19718,N_19365);
or UO_2026 (O_2026,N_19220,N_19252);
xnor UO_2027 (O_2027,N_19201,N_19637);
or UO_2028 (O_2028,N_19863,N_19378);
nand UO_2029 (O_2029,N_19436,N_19783);
nand UO_2030 (O_2030,N_19600,N_19710);
and UO_2031 (O_2031,N_19582,N_19402);
and UO_2032 (O_2032,N_19865,N_19724);
or UO_2033 (O_2033,N_19555,N_19618);
nor UO_2034 (O_2034,N_19485,N_19327);
or UO_2035 (O_2035,N_19636,N_19747);
and UO_2036 (O_2036,N_19528,N_19898);
xnor UO_2037 (O_2037,N_19813,N_19840);
xor UO_2038 (O_2038,N_19663,N_19269);
xor UO_2039 (O_2039,N_19679,N_19994);
and UO_2040 (O_2040,N_19869,N_19220);
nor UO_2041 (O_2041,N_19907,N_19223);
or UO_2042 (O_2042,N_19637,N_19268);
nor UO_2043 (O_2043,N_19718,N_19904);
nor UO_2044 (O_2044,N_19388,N_19233);
or UO_2045 (O_2045,N_19405,N_19258);
nor UO_2046 (O_2046,N_19469,N_19562);
nor UO_2047 (O_2047,N_19435,N_19791);
xor UO_2048 (O_2048,N_19899,N_19695);
xor UO_2049 (O_2049,N_19420,N_19261);
xor UO_2050 (O_2050,N_19249,N_19994);
and UO_2051 (O_2051,N_19416,N_19948);
or UO_2052 (O_2052,N_19803,N_19902);
or UO_2053 (O_2053,N_19425,N_19535);
or UO_2054 (O_2054,N_19582,N_19494);
nand UO_2055 (O_2055,N_19327,N_19601);
nand UO_2056 (O_2056,N_19216,N_19390);
and UO_2057 (O_2057,N_19531,N_19408);
and UO_2058 (O_2058,N_19904,N_19389);
xor UO_2059 (O_2059,N_19896,N_19871);
and UO_2060 (O_2060,N_19349,N_19655);
and UO_2061 (O_2061,N_19528,N_19498);
nand UO_2062 (O_2062,N_19725,N_19530);
nand UO_2063 (O_2063,N_19271,N_19658);
and UO_2064 (O_2064,N_19498,N_19729);
nor UO_2065 (O_2065,N_19977,N_19695);
and UO_2066 (O_2066,N_19729,N_19548);
and UO_2067 (O_2067,N_19940,N_19380);
and UO_2068 (O_2068,N_19627,N_19649);
nand UO_2069 (O_2069,N_19830,N_19820);
nand UO_2070 (O_2070,N_19806,N_19326);
nor UO_2071 (O_2071,N_19387,N_19326);
nor UO_2072 (O_2072,N_19893,N_19438);
nand UO_2073 (O_2073,N_19544,N_19205);
nand UO_2074 (O_2074,N_19317,N_19258);
nor UO_2075 (O_2075,N_19507,N_19656);
nor UO_2076 (O_2076,N_19922,N_19973);
xor UO_2077 (O_2077,N_19630,N_19924);
and UO_2078 (O_2078,N_19635,N_19417);
nor UO_2079 (O_2079,N_19580,N_19428);
and UO_2080 (O_2080,N_19663,N_19902);
nand UO_2081 (O_2081,N_19964,N_19200);
nand UO_2082 (O_2082,N_19756,N_19412);
nor UO_2083 (O_2083,N_19679,N_19353);
or UO_2084 (O_2084,N_19874,N_19530);
and UO_2085 (O_2085,N_19915,N_19760);
or UO_2086 (O_2086,N_19658,N_19515);
xor UO_2087 (O_2087,N_19205,N_19593);
and UO_2088 (O_2088,N_19710,N_19925);
nand UO_2089 (O_2089,N_19353,N_19237);
or UO_2090 (O_2090,N_19873,N_19340);
and UO_2091 (O_2091,N_19779,N_19439);
nand UO_2092 (O_2092,N_19539,N_19614);
nand UO_2093 (O_2093,N_19535,N_19445);
nor UO_2094 (O_2094,N_19633,N_19692);
nor UO_2095 (O_2095,N_19985,N_19300);
nand UO_2096 (O_2096,N_19267,N_19501);
xor UO_2097 (O_2097,N_19598,N_19680);
xnor UO_2098 (O_2098,N_19667,N_19451);
nand UO_2099 (O_2099,N_19579,N_19294);
nor UO_2100 (O_2100,N_19475,N_19910);
nor UO_2101 (O_2101,N_19515,N_19826);
nand UO_2102 (O_2102,N_19773,N_19883);
or UO_2103 (O_2103,N_19921,N_19247);
and UO_2104 (O_2104,N_19300,N_19421);
xor UO_2105 (O_2105,N_19790,N_19704);
xor UO_2106 (O_2106,N_19591,N_19252);
xnor UO_2107 (O_2107,N_19635,N_19685);
nor UO_2108 (O_2108,N_19733,N_19313);
nand UO_2109 (O_2109,N_19744,N_19257);
nand UO_2110 (O_2110,N_19283,N_19580);
nor UO_2111 (O_2111,N_19692,N_19718);
nand UO_2112 (O_2112,N_19351,N_19417);
xnor UO_2113 (O_2113,N_19489,N_19893);
xnor UO_2114 (O_2114,N_19391,N_19408);
and UO_2115 (O_2115,N_19770,N_19697);
nand UO_2116 (O_2116,N_19396,N_19243);
or UO_2117 (O_2117,N_19447,N_19822);
nor UO_2118 (O_2118,N_19386,N_19352);
nand UO_2119 (O_2119,N_19433,N_19515);
xor UO_2120 (O_2120,N_19298,N_19386);
and UO_2121 (O_2121,N_19255,N_19864);
xnor UO_2122 (O_2122,N_19717,N_19798);
xnor UO_2123 (O_2123,N_19974,N_19557);
nor UO_2124 (O_2124,N_19770,N_19392);
nand UO_2125 (O_2125,N_19863,N_19488);
xnor UO_2126 (O_2126,N_19480,N_19488);
nand UO_2127 (O_2127,N_19859,N_19534);
xor UO_2128 (O_2128,N_19941,N_19917);
or UO_2129 (O_2129,N_19972,N_19636);
xnor UO_2130 (O_2130,N_19274,N_19745);
nor UO_2131 (O_2131,N_19743,N_19705);
nor UO_2132 (O_2132,N_19602,N_19225);
xnor UO_2133 (O_2133,N_19859,N_19388);
nor UO_2134 (O_2134,N_19642,N_19533);
xor UO_2135 (O_2135,N_19704,N_19658);
or UO_2136 (O_2136,N_19226,N_19445);
xor UO_2137 (O_2137,N_19730,N_19249);
xnor UO_2138 (O_2138,N_19712,N_19983);
nand UO_2139 (O_2139,N_19970,N_19828);
or UO_2140 (O_2140,N_19386,N_19225);
xnor UO_2141 (O_2141,N_19756,N_19619);
nor UO_2142 (O_2142,N_19980,N_19347);
and UO_2143 (O_2143,N_19448,N_19863);
nor UO_2144 (O_2144,N_19580,N_19363);
xor UO_2145 (O_2145,N_19544,N_19757);
and UO_2146 (O_2146,N_19690,N_19848);
nand UO_2147 (O_2147,N_19923,N_19330);
nand UO_2148 (O_2148,N_19320,N_19314);
or UO_2149 (O_2149,N_19306,N_19619);
nand UO_2150 (O_2150,N_19456,N_19599);
nor UO_2151 (O_2151,N_19215,N_19976);
and UO_2152 (O_2152,N_19422,N_19595);
or UO_2153 (O_2153,N_19844,N_19611);
nand UO_2154 (O_2154,N_19608,N_19247);
xor UO_2155 (O_2155,N_19349,N_19205);
nor UO_2156 (O_2156,N_19854,N_19545);
nor UO_2157 (O_2157,N_19391,N_19385);
and UO_2158 (O_2158,N_19890,N_19924);
nand UO_2159 (O_2159,N_19753,N_19494);
or UO_2160 (O_2160,N_19997,N_19688);
nand UO_2161 (O_2161,N_19882,N_19755);
nand UO_2162 (O_2162,N_19426,N_19654);
xor UO_2163 (O_2163,N_19844,N_19837);
xnor UO_2164 (O_2164,N_19482,N_19562);
and UO_2165 (O_2165,N_19288,N_19483);
xnor UO_2166 (O_2166,N_19556,N_19572);
and UO_2167 (O_2167,N_19726,N_19632);
or UO_2168 (O_2168,N_19703,N_19859);
xnor UO_2169 (O_2169,N_19499,N_19973);
and UO_2170 (O_2170,N_19516,N_19820);
nor UO_2171 (O_2171,N_19556,N_19307);
or UO_2172 (O_2172,N_19681,N_19993);
nor UO_2173 (O_2173,N_19850,N_19598);
nor UO_2174 (O_2174,N_19621,N_19203);
and UO_2175 (O_2175,N_19836,N_19820);
or UO_2176 (O_2176,N_19375,N_19913);
nand UO_2177 (O_2177,N_19594,N_19892);
xnor UO_2178 (O_2178,N_19931,N_19799);
or UO_2179 (O_2179,N_19442,N_19814);
xor UO_2180 (O_2180,N_19235,N_19977);
xnor UO_2181 (O_2181,N_19502,N_19595);
and UO_2182 (O_2182,N_19552,N_19859);
or UO_2183 (O_2183,N_19960,N_19217);
and UO_2184 (O_2184,N_19823,N_19447);
and UO_2185 (O_2185,N_19642,N_19668);
or UO_2186 (O_2186,N_19540,N_19534);
and UO_2187 (O_2187,N_19409,N_19307);
nand UO_2188 (O_2188,N_19373,N_19896);
nor UO_2189 (O_2189,N_19773,N_19962);
nand UO_2190 (O_2190,N_19882,N_19707);
and UO_2191 (O_2191,N_19759,N_19474);
nand UO_2192 (O_2192,N_19251,N_19482);
nand UO_2193 (O_2193,N_19274,N_19439);
and UO_2194 (O_2194,N_19928,N_19478);
nand UO_2195 (O_2195,N_19584,N_19523);
or UO_2196 (O_2196,N_19807,N_19636);
nor UO_2197 (O_2197,N_19334,N_19396);
nand UO_2198 (O_2198,N_19204,N_19757);
nor UO_2199 (O_2199,N_19799,N_19999);
xnor UO_2200 (O_2200,N_19210,N_19762);
xnor UO_2201 (O_2201,N_19509,N_19969);
nor UO_2202 (O_2202,N_19910,N_19882);
and UO_2203 (O_2203,N_19533,N_19513);
nor UO_2204 (O_2204,N_19477,N_19909);
or UO_2205 (O_2205,N_19731,N_19548);
or UO_2206 (O_2206,N_19954,N_19754);
nor UO_2207 (O_2207,N_19594,N_19701);
nand UO_2208 (O_2208,N_19416,N_19451);
and UO_2209 (O_2209,N_19429,N_19258);
nand UO_2210 (O_2210,N_19820,N_19915);
and UO_2211 (O_2211,N_19704,N_19742);
nor UO_2212 (O_2212,N_19937,N_19953);
xnor UO_2213 (O_2213,N_19456,N_19654);
and UO_2214 (O_2214,N_19720,N_19458);
xnor UO_2215 (O_2215,N_19223,N_19438);
xnor UO_2216 (O_2216,N_19317,N_19869);
nand UO_2217 (O_2217,N_19991,N_19786);
or UO_2218 (O_2218,N_19608,N_19964);
nor UO_2219 (O_2219,N_19799,N_19324);
and UO_2220 (O_2220,N_19579,N_19499);
xor UO_2221 (O_2221,N_19979,N_19383);
and UO_2222 (O_2222,N_19559,N_19473);
and UO_2223 (O_2223,N_19352,N_19730);
xor UO_2224 (O_2224,N_19306,N_19264);
nor UO_2225 (O_2225,N_19623,N_19819);
xnor UO_2226 (O_2226,N_19414,N_19573);
or UO_2227 (O_2227,N_19427,N_19865);
nand UO_2228 (O_2228,N_19615,N_19928);
nor UO_2229 (O_2229,N_19861,N_19742);
and UO_2230 (O_2230,N_19895,N_19463);
or UO_2231 (O_2231,N_19207,N_19701);
nand UO_2232 (O_2232,N_19353,N_19219);
nand UO_2233 (O_2233,N_19438,N_19594);
xor UO_2234 (O_2234,N_19456,N_19607);
nor UO_2235 (O_2235,N_19317,N_19443);
and UO_2236 (O_2236,N_19693,N_19773);
nand UO_2237 (O_2237,N_19494,N_19689);
and UO_2238 (O_2238,N_19939,N_19903);
and UO_2239 (O_2239,N_19502,N_19616);
xnor UO_2240 (O_2240,N_19424,N_19578);
and UO_2241 (O_2241,N_19332,N_19445);
xor UO_2242 (O_2242,N_19782,N_19721);
nand UO_2243 (O_2243,N_19495,N_19784);
or UO_2244 (O_2244,N_19918,N_19207);
nand UO_2245 (O_2245,N_19591,N_19574);
or UO_2246 (O_2246,N_19585,N_19447);
and UO_2247 (O_2247,N_19480,N_19543);
nand UO_2248 (O_2248,N_19665,N_19910);
or UO_2249 (O_2249,N_19316,N_19670);
xnor UO_2250 (O_2250,N_19850,N_19486);
xor UO_2251 (O_2251,N_19412,N_19989);
and UO_2252 (O_2252,N_19248,N_19482);
and UO_2253 (O_2253,N_19742,N_19482);
and UO_2254 (O_2254,N_19566,N_19922);
or UO_2255 (O_2255,N_19364,N_19479);
xor UO_2256 (O_2256,N_19666,N_19633);
xor UO_2257 (O_2257,N_19741,N_19781);
xor UO_2258 (O_2258,N_19386,N_19879);
and UO_2259 (O_2259,N_19491,N_19676);
nand UO_2260 (O_2260,N_19471,N_19805);
xor UO_2261 (O_2261,N_19319,N_19687);
nand UO_2262 (O_2262,N_19243,N_19275);
or UO_2263 (O_2263,N_19824,N_19539);
xor UO_2264 (O_2264,N_19871,N_19922);
xnor UO_2265 (O_2265,N_19443,N_19874);
xnor UO_2266 (O_2266,N_19443,N_19471);
nor UO_2267 (O_2267,N_19593,N_19488);
xnor UO_2268 (O_2268,N_19230,N_19661);
nand UO_2269 (O_2269,N_19340,N_19445);
and UO_2270 (O_2270,N_19507,N_19634);
or UO_2271 (O_2271,N_19226,N_19947);
xnor UO_2272 (O_2272,N_19570,N_19859);
nand UO_2273 (O_2273,N_19339,N_19360);
or UO_2274 (O_2274,N_19834,N_19841);
or UO_2275 (O_2275,N_19811,N_19236);
nand UO_2276 (O_2276,N_19776,N_19393);
nor UO_2277 (O_2277,N_19523,N_19686);
nand UO_2278 (O_2278,N_19757,N_19480);
and UO_2279 (O_2279,N_19294,N_19979);
xnor UO_2280 (O_2280,N_19493,N_19355);
nor UO_2281 (O_2281,N_19933,N_19964);
nor UO_2282 (O_2282,N_19692,N_19568);
nor UO_2283 (O_2283,N_19590,N_19354);
xnor UO_2284 (O_2284,N_19295,N_19517);
and UO_2285 (O_2285,N_19658,N_19238);
and UO_2286 (O_2286,N_19233,N_19648);
xnor UO_2287 (O_2287,N_19963,N_19456);
or UO_2288 (O_2288,N_19816,N_19531);
or UO_2289 (O_2289,N_19982,N_19612);
xor UO_2290 (O_2290,N_19738,N_19285);
or UO_2291 (O_2291,N_19979,N_19893);
or UO_2292 (O_2292,N_19664,N_19549);
xnor UO_2293 (O_2293,N_19962,N_19756);
xor UO_2294 (O_2294,N_19644,N_19309);
or UO_2295 (O_2295,N_19652,N_19277);
or UO_2296 (O_2296,N_19284,N_19374);
nor UO_2297 (O_2297,N_19404,N_19221);
and UO_2298 (O_2298,N_19243,N_19803);
and UO_2299 (O_2299,N_19703,N_19207);
nand UO_2300 (O_2300,N_19965,N_19204);
nor UO_2301 (O_2301,N_19254,N_19906);
and UO_2302 (O_2302,N_19558,N_19211);
xnor UO_2303 (O_2303,N_19951,N_19766);
xnor UO_2304 (O_2304,N_19435,N_19842);
xnor UO_2305 (O_2305,N_19625,N_19581);
nand UO_2306 (O_2306,N_19602,N_19228);
xnor UO_2307 (O_2307,N_19632,N_19463);
nand UO_2308 (O_2308,N_19798,N_19969);
nor UO_2309 (O_2309,N_19553,N_19223);
and UO_2310 (O_2310,N_19818,N_19479);
xnor UO_2311 (O_2311,N_19544,N_19704);
nand UO_2312 (O_2312,N_19362,N_19487);
nand UO_2313 (O_2313,N_19258,N_19368);
nor UO_2314 (O_2314,N_19382,N_19989);
xor UO_2315 (O_2315,N_19772,N_19765);
nor UO_2316 (O_2316,N_19741,N_19359);
nor UO_2317 (O_2317,N_19472,N_19407);
or UO_2318 (O_2318,N_19692,N_19485);
nor UO_2319 (O_2319,N_19438,N_19943);
xnor UO_2320 (O_2320,N_19900,N_19961);
and UO_2321 (O_2321,N_19506,N_19574);
or UO_2322 (O_2322,N_19624,N_19469);
nor UO_2323 (O_2323,N_19340,N_19605);
nor UO_2324 (O_2324,N_19672,N_19835);
nand UO_2325 (O_2325,N_19443,N_19403);
nand UO_2326 (O_2326,N_19808,N_19785);
or UO_2327 (O_2327,N_19354,N_19748);
and UO_2328 (O_2328,N_19945,N_19202);
or UO_2329 (O_2329,N_19546,N_19469);
nor UO_2330 (O_2330,N_19443,N_19589);
nor UO_2331 (O_2331,N_19664,N_19628);
and UO_2332 (O_2332,N_19592,N_19334);
xor UO_2333 (O_2333,N_19820,N_19221);
nor UO_2334 (O_2334,N_19293,N_19978);
nand UO_2335 (O_2335,N_19612,N_19911);
xor UO_2336 (O_2336,N_19344,N_19610);
nor UO_2337 (O_2337,N_19826,N_19711);
nor UO_2338 (O_2338,N_19773,N_19367);
xor UO_2339 (O_2339,N_19506,N_19877);
xor UO_2340 (O_2340,N_19278,N_19446);
nand UO_2341 (O_2341,N_19386,N_19654);
xnor UO_2342 (O_2342,N_19607,N_19870);
nor UO_2343 (O_2343,N_19849,N_19876);
nand UO_2344 (O_2344,N_19924,N_19677);
and UO_2345 (O_2345,N_19905,N_19548);
or UO_2346 (O_2346,N_19350,N_19983);
nor UO_2347 (O_2347,N_19341,N_19497);
nor UO_2348 (O_2348,N_19309,N_19885);
and UO_2349 (O_2349,N_19678,N_19595);
nor UO_2350 (O_2350,N_19472,N_19307);
nor UO_2351 (O_2351,N_19575,N_19852);
or UO_2352 (O_2352,N_19387,N_19569);
and UO_2353 (O_2353,N_19555,N_19305);
and UO_2354 (O_2354,N_19784,N_19948);
or UO_2355 (O_2355,N_19799,N_19609);
nand UO_2356 (O_2356,N_19343,N_19630);
xnor UO_2357 (O_2357,N_19309,N_19450);
xnor UO_2358 (O_2358,N_19257,N_19626);
nand UO_2359 (O_2359,N_19240,N_19812);
or UO_2360 (O_2360,N_19698,N_19250);
nand UO_2361 (O_2361,N_19451,N_19590);
nor UO_2362 (O_2362,N_19668,N_19465);
xnor UO_2363 (O_2363,N_19646,N_19542);
nand UO_2364 (O_2364,N_19367,N_19268);
or UO_2365 (O_2365,N_19412,N_19909);
and UO_2366 (O_2366,N_19257,N_19476);
nor UO_2367 (O_2367,N_19508,N_19238);
and UO_2368 (O_2368,N_19922,N_19964);
nand UO_2369 (O_2369,N_19561,N_19294);
xnor UO_2370 (O_2370,N_19706,N_19824);
or UO_2371 (O_2371,N_19368,N_19850);
xnor UO_2372 (O_2372,N_19816,N_19932);
nand UO_2373 (O_2373,N_19226,N_19413);
or UO_2374 (O_2374,N_19756,N_19827);
xor UO_2375 (O_2375,N_19285,N_19920);
nor UO_2376 (O_2376,N_19492,N_19673);
and UO_2377 (O_2377,N_19906,N_19809);
nor UO_2378 (O_2378,N_19886,N_19744);
or UO_2379 (O_2379,N_19809,N_19284);
nor UO_2380 (O_2380,N_19326,N_19377);
or UO_2381 (O_2381,N_19338,N_19951);
nand UO_2382 (O_2382,N_19646,N_19798);
nand UO_2383 (O_2383,N_19603,N_19301);
or UO_2384 (O_2384,N_19878,N_19465);
xor UO_2385 (O_2385,N_19423,N_19719);
xor UO_2386 (O_2386,N_19878,N_19688);
or UO_2387 (O_2387,N_19879,N_19552);
nand UO_2388 (O_2388,N_19282,N_19239);
xnor UO_2389 (O_2389,N_19360,N_19485);
and UO_2390 (O_2390,N_19627,N_19745);
nor UO_2391 (O_2391,N_19972,N_19530);
nor UO_2392 (O_2392,N_19815,N_19958);
and UO_2393 (O_2393,N_19322,N_19608);
xor UO_2394 (O_2394,N_19264,N_19922);
nor UO_2395 (O_2395,N_19443,N_19817);
or UO_2396 (O_2396,N_19665,N_19392);
and UO_2397 (O_2397,N_19461,N_19819);
nand UO_2398 (O_2398,N_19287,N_19499);
xor UO_2399 (O_2399,N_19964,N_19360);
xor UO_2400 (O_2400,N_19985,N_19979);
and UO_2401 (O_2401,N_19865,N_19575);
or UO_2402 (O_2402,N_19723,N_19997);
or UO_2403 (O_2403,N_19991,N_19288);
nor UO_2404 (O_2404,N_19285,N_19841);
nand UO_2405 (O_2405,N_19854,N_19731);
nor UO_2406 (O_2406,N_19547,N_19499);
or UO_2407 (O_2407,N_19999,N_19440);
and UO_2408 (O_2408,N_19674,N_19247);
nor UO_2409 (O_2409,N_19232,N_19629);
nand UO_2410 (O_2410,N_19824,N_19336);
and UO_2411 (O_2411,N_19673,N_19816);
and UO_2412 (O_2412,N_19631,N_19771);
nor UO_2413 (O_2413,N_19533,N_19946);
nand UO_2414 (O_2414,N_19885,N_19705);
nor UO_2415 (O_2415,N_19573,N_19757);
nand UO_2416 (O_2416,N_19872,N_19976);
xor UO_2417 (O_2417,N_19356,N_19774);
xnor UO_2418 (O_2418,N_19453,N_19247);
nand UO_2419 (O_2419,N_19289,N_19260);
xnor UO_2420 (O_2420,N_19298,N_19483);
xor UO_2421 (O_2421,N_19377,N_19363);
or UO_2422 (O_2422,N_19961,N_19938);
or UO_2423 (O_2423,N_19717,N_19378);
or UO_2424 (O_2424,N_19601,N_19408);
and UO_2425 (O_2425,N_19719,N_19927);
or UO_2426 (O_2426,N_19206,N_19535);
xnor UO_2427 (O_2427,N_19347,N_19981);
xnor UO_2428 (O_2428,N_19762,N_19316);
or UO_2429 (O_2429,N_19445,N_19583);
nand UO_2430 (O_2430,N_19593,N_19982);
nand UO_2431 (O_2431,N_19441,N_19377);
nand UO_2432 (O_2432,N_19813,N_19754);
nand UO_2433 (O_2433,N_19736,N_19235);
nand UO_2434 (O_2434,N_19850,N_19691);
or UO_2435 (O_2435,N_19227,N_19336);
xnor UO_2436 (O_2436,N_19681,N_19992);
nor UO_2437 (O_2437,N_19499,N_19225);
nand UO_2438 (O_2438,N_19394,N_19398);
and UO_2439 (O_2439,N_19719,N_19636);
or UO_2440 (O_2440,N_19643,N_19576);
nor UO_2441 (O_2441,N_19436,N_19518);
or UO_2442 (O_2442,N_19934,N_19403);
and UO_2443 (O_2443,N_19613,N_19675);
and UO_2444 (O_2444,N_19512,N_19615);
xnor UO_2445 (O_2445,N_19426,N_19436);
xor UO_2446 (O_2446,N_19783,N_19979);
and UO_2447 (O_2447,N_19505,N_19937);
nand UO_2448 (O_2448,N_19783,N_19809);
nand UO_2449 (O_2449,N_19776,N_19481);
nor UO_2450 (O_2450,N_19966,N_19527);
nor UO_2451 (O_2451,N_19372,N_19634);
and UO_2452 (O_2452,N_19998,N_19371);
nor UO_2453 (O_2453,N_19496,N_19590);
xor UO_2454 (O_2454,N_19751,N_19825);
and UO_2455 (O_2455,N_19520,N_19292);
or UO_2456 (O_2456,N_19255,N_19998);
xnor UO_2457 (O_2457,N_19706,N_19379);
and UO_2458 (O_2458,N_19364,N_19213);
nor UO_2459 (O_2459,N_19749,N_19890);
xnor UO_2460 (O_2460,N_19730,N_19546);
nor UO_2461 (O_2461,N_19846,N_19745);
nor UO_2462 (O_2462,N_19782,N_19906);
and UO_2463 (O_2463,N_19827,N_19856);
xor UO_2464 (O_2464,N_19974,N_19582);
and UO_2465 (O_2465,N_19424,N_19546);
nand UO_2466 (O_2466,N_19606,N_19824);
or UO_2467 (O_2467,N_19858,N_19827);
and UO_2468 (O_2468,N_19600,N_19735);
and UO_2469 (O_2469,N_19943,N_19517);
or UO_2470 (O_2470,N_19212,N_19810);
xor UO_2471 (O_2471,N_19602,N_19209);
nor UO_2472 (O_2472,N_19703,N_19323);
nand UO_2473 (O_2473,N_19210,N_19860);
and UO_2474 (O_2474,N_19934,N_19364);
or UO_2475 (O_2475,N_19623,N_19288);
nor UO_2476 (O_2476,N_19376,N_19453);
and UO_2477 (O_2477,N_19214,N_19588);
nand UO_2478 (O_2478,N_19576,N_19926);
xnor UO_2479 (O_2479,N_19876,N_19871);
nand UO_2480 (O_2480,N_19972,N_19576);
or UO_2481 (O_2481,N_19344,N_19698);
nor UO_2482 (O_2482,N_19247,N_19531);
and UO_2483 (O_2483,N_19875,N_19689);
nand UO_2484 (O_2484,N_19829,N_19905);
and UO_2485 (O_2485,N_19642,N_19318);
nand UO_2486 (O_2486,N_19821,N_19265);
and UO_2487 (O_2487,N_19481,N_19661);
nand UO_2488 (O_2488,N_19770,N_19759);
nand UO_2489 (O_2489,N_19624,N_19537);
nand UO_2490 (O_2490,N_19483,N_19352);
nor UO_2491 (O_2491,N_19825,N_19245);
xor UO_2492 (O_2492,N_19704,N_19987);
or UO_2493 (O_2493,N_19778,N_19682);
or UO_2494 (O_2494,N_19654,N_19885);
xor UO_2495 (O_2495,N_19954,N_19571);
nor UO_2496 (O_2496,N_19998,N_19740);
or UO_2497 (O_2497,N_19235,N_19535);
or UO_2498 (O_2498,N_19938,N_19864);
or UO_2499 (O_2499,N_19909,N_19485);
endmodule