module basic_500_3000_500_6_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_481,In_444);
nor U1 (N_1,In_25,In_119);
or U2 (N_2,In_190,In_46);
nand U3 (N_3,In_62,In_290);
nor U4 (N_4,In_122,In_333);
xor U5 (N_5,In_467,In_446);
nand U6 (N_6,In_71,In_200);
and U7 (N_7,In_284,In_322);
and U8 (N_8,In_246,In_282);
nand U9 (N_9,In_330,In_240);
nor U10 (N_10,In_9,In_139);
or U11 (N_11,In_472,In_499);
nand U12 (N_12,In_430,In_41);
or U13 (N_13,In_453,In_85);
or U14 (N_14,In_188,In_103);
or U15 (N_15,In_293,In_329);
or U16 (N_16,In_59,In_133);
xnor U17 (N_17,In_64,In_318);
nand U18 (N_18,In_118,In_101);
nor U19 (N_19,In_38,In_3);
nor U20 (N_20,In_301,In_313);
or U21 (N_21,In_392,In_332);
and U22 (N_22,In_275,In_426);
xor U23 (N_23,In_482,In_311);
nand U24 (N_24,In_255,In_74);
nor U25 (N_25,In_107,In_160);
nor U26 (N_26,In_123,In_184);
nand U27 (N_27,In_115,In_137);
and U28 (N_28,In_490,In_89);
and U29 (N_29,In_324,In_36);
and U30 (N_30,In_341,In_323);
nand U31 (N_31,In_68,In_460);
nor U32 (N_32,In_13,In_286);
and U33 (N_33,In_479,In_358);
and U34 (N_34,In_28,In_164);
nor U35 (N_35,In_335,In_17);
and U36 (N_36,In_11,In_440);
and U37 (N_37,In_260,In_40);
or U38 (N_38,In_245,In_43);
xnor U39 (N_39,In_203,In_56);
and U40 (N_40,In_256,In_192);
or U41 (N_41,In_242,In_497);
nor U42 (N_42,In_304,In_182);
and U43 (N_43,In_208,In_54);
nor U44 (N_44,In_220,In_194);
and U45 (N_45,In_196,In_369);
and U46 (N_46,In_69,In_129);
nor U47 (N_47,In_469,In_209);
or U48 (N_48,In_436,In_462);
nand U49 (N_49,In_211,In_90);
nand U50 (N_50,In_361,In_346);
nand U51 (N_51,In_165,In_105);
xnor U52 (N_52,In_20,In_163);
and U53 (N_53,In_47,In_368);
nand U54 (N_54,In_404,In_77);
nor U55 (N_55,In_87,In_224);
and U56 (N_56,In_433,In_14);
or U57 (N_57,In_178,In_191);
nor U58 (N_58,In_32,In_314);
and U59 (N_59,In_398,In_104);
xor U60 (N_60,In_340,In_316);
nand U61 (N_61,In_420,In_63);
nor U62 (N_62,In_276,In_2);
xor U63 (N_63,In_488,In_266);
nand U64 (N_64,In_130,In_249);
nand U65 (N_65,In_327,In_253);
nor U66 (N_66,In_379,In_179);
or U67 (N_67,In_8,In_274);
and U68 (N_68,In_371,In_149);
nand U69 (N_69,In_380,In_342);
nor U70 (N_70,In_31,In_365);
or U71 (N_71,In_385,In_394);
or U72 (N_72,In_432,In_108);
or U73 (N_73,In_66,In_378);
nor U74 (N_74,In_262,In_395);
or U75 (N_75,In_4,In_70);
or U76 (N_76,In_307,In_281);
or U77 (N_77,In_35,In_489);
and U78 (N_78,In_474,In_429);
or U79 (N_79,In_278,In_338);
and U80 (N_80,In_265,In_228);
nor U81 (N_81,In_112,In_232);
nor U82 (N_82,In_351,In_187);
nand U83 (N_83,In_494,In_498);
and U84 (N_84,In_419,In_10);
and U85 (N_85,In_331,In_78);
and U86 (N_86,In_389,In_128);
nor U87 (N_87,In_248,In_213);
nand U88 (N_88,In_388,In_458);
xor U89 (N_89,In_243,In_370);
and U90 (N_90,In_470,In_212);
nor U91 (N_91,In_382,In_7);
nor U92 (N_92,In_259,In_124);
nand U93 (N_93,In_1,In_496);
nor U94 (N_94,In_390,In_95);
and U95 (N_95,In_448,In_493);
or U96 (N_96,In_227,In_268);
nand U97 (N_97,In_152,In_310);
or U98 (N_98,In_263,In_306);
nand U99 (N_99,In_159,In_477);
or U100 (N_100,In_218,In_174);
or U101 (N_101,In_29,In_162);
and U102 (N_102,In_277,In_72);
nand U103 (N_103,In_297,In_219);
nand U104 (N_104,In_229,In_261);
nor U105 (N_105,In_45,In_201);
nor U106 (N_106,In_173,In_347);
or U107 (N_107,In_121,In_237);
nor U108 (N_108,In_391,In_126);
and U109 (N_109,In_355,In_403);
or U110 (N_110,In_143,In_483);
and U111 (N_111,In_199,In_473);
and U112 (N_112,In_65,In_442);
and U113 (N_113,In_405,In_186);
or U114 (N_114,In_250,In_37);
or U115 (N_115,In_450,In_67);
nand U116 (N_116,In_337,In_258);
and U117 (N_117,In_106,In_454);
nor U118 (N_118,In_315,In_157);
nand U119 (N_119,In_295,In_50);
nor U120 (N_120,In_471,In_94);
nand U121 (N_121,In_434,In_6);
or U122 (N_122,In_366,In_49);
xor U123 (N_123,In_58,In_110);
xnor U124 (N_124,In_197,In_23);
nor U125 (N_125,In_92,In_222);
nand U126 (N_126,In_456,In_424);
nor U127 (N_127,In_257,In_406);
nor U128 (N_128,In_421,In_233);
or U129 (N_129,In_99,In_81);
and U130 (N_130,In_21,In_189);
nand U131 (N_131,In_384,In_397);
nand U132 (N_132,In_180,In_113);
and U133 (N_133,In_270,In_480);
or U134 (N_134,In_412,In_158);
nor U135 (N_135,In_252,In_308);
and U136 (N_136,In_125,In_296);
nand U137 (N_137,In_217,In_247);
or U138 (N_138,In_451,In_349);
and U139 (N_139,In_417,In_215);
and U140 (N_140,In_207,In_98);
nor U141 (N_141,In_326,In_16);
and U142 (N_142,In_53,In_413);
and U143 (N_143,In_445,In_334);
or U144 (N_144,In_84,In_373);
xnor U145 (N_145,In_466,In_39);
or U146 (N_146,In_485,In_280);
nand U147 (N_147,In_343,In_377);
and U148 (N_148,In_131,In_264);
and U149 (N_149,In_150,In_367);
or U150 (N_150,In_435,In_291);
nor U151 (N_151,In_399,In_336);
xnor U152 (N_152,In_177,In_96);
or U153 (N_153,In_487,In_18);
nand U154 (N_154,In_210,In_411);
and U155 (N_155,In_86,In_302);
and U156 (N_156,In_309,In_166);
nand U157 (N_157,In_205,In_319);
nand U158 (N_158,In_231,In_492);
nor U159 (N_159,In_476,In_431);
nand U160 (N_160,In_27,In_52);
nor U161 (N_161,In_26,In_285);
nor U162 (N_162,In_386,In_321);
xor U163 (N_163,In_34,In_5);
nor U164 (N_164,In_48,In_147);
or U165 (N_165,In_272,In_168);
or U166 (N_166,In_475,In_292);
or U167 (N_167,In_57,In_100);
or U168 (N_168,In_51,In_19);
and U169 (N_169,In_61,In_279);
nor U170 (N_170,In_452,In_195);
nor U171 (N_171,In_269,In_423);
or U172 (N_172,In_97,In_238);
nor U173 (N_173,In_114,In_93);
or U174 (N_174,In_364,In_409);
or U175 (N_175,In_127,In_156);
and U176 (N_176,In_437,In_354);
nor U177 (N_177,In_294,In_396);
xor U178 (N_178,In_486,In_142);
nand U179 (N_179,In_387,In_225);
and U180 (N_180,In_353,In_161);
and U181 (N_181,In_441,In_414);
nor U182 (N_182,In_339,In_464);
nand U183 (N_183,In_136,In_241);
and U184 (N_184,In_167,In_172);
xor U185 (N_185,In_300,In_244);
nor U186 (N_186,In_181,In_221);
xor U187 (N_187,In_465,In_216);
or U188 (N_188,In_102,In_468);
or U189 (N_189,In_317,In_75);
or U190 (N_190,In_374,In_138);
or U191 (N_191,In_185,In_357);
nand U192 (N_192,In_155,In_42);
or U193 (N_193,In_345,In_193);
nand U194 (N_194,In_134,In_350);
xnor U195 (N_195,In_44,In_55);
nand U196 (N_196,In_375,In_202);
and U197 (N_197,In_271,In_145);
nor U198 (N_198,In_132,In_60);
and U199 (N_199,In_383,In_363);
and U200 (N_200,In_267,In_116);
nor U201 (N_201,In_325,In_381);
and U202 (N_202,In_24,In_299);
and U203 (N_203,In_356,In_457);
and U204 (N_204,In_204,In_15);
nand U205 (N_205,In_273,In_30);
nand U206 (N_206,In_140,In_352);
or U207 (N_207,In_214,In_88);
xor U208 (N_208,In_117,In_425);
nand U209 (N_209,In_459,In_234);
nand U210 (N_210,In_175,In_236);
or U211 (N_211,In_120,In_415);
and U212 (N_212,In_410,In_455);
or U213 (N_213,In_359,In_146);
nand U214 (N_214,In_289,In_298);
and U215 (N_215,In_461,In_428);
or U216 (N_216,In_495,In_491);
nor U217 (N_217,In_449,In_109);
nand U218 (N_218,In_484,In_206);
and U219 (N_219,In_376,In_401);
nand U220 (N_220,In_416,In_312);
xor U221 (N_221,In_223,In_239);
or U222 (N_222,In_151,In_80);
and U223 (N_223,In_393,In_226);
nor U224 (N_224,In_183,In_303);
and U225 (N_225,In_344,In_283);
nor U226 (N_226,In_22,In_141);
or U227 (N_227,In_73,In_443);
nor U228 (N_228,In_320,In_362);
nand U229 (N_229,In_407,In_402);
nand U230 (N_230,In_12,In_360);
and U231 (N_231,In_76,In_328);
or U232 (N_232,In_230,In_478);
or U233 (N_233,In_372,In_169);
and U234 (N_234,In_400,In_408);
xnor U235 (N_235,In_235,In_135);
or U236 (N_236,In_148,In_170);
nor U237 (N_237,In_288,In_0);
or U238 (N_238,In_254,In_287);
xnor U239 (N_239,In_251,In_176);
xnor U240 (N_240,In_154,In_463);
or U241 (N_241,In_447,In_83);
nand U242 (N_242,In_427,In_348);
nand U243 (N_243,In_305,In_111);
nand U244 (N_244,In_439,In_422);
nand U245 (N_245,In_33,In_153);
or U246 (N_246,In_144,In_171);
or U247 (N_247,In_198,In_79);
or U248 (N_248,In_91,In_82);
nand U249 (N_249,In_418,In_438);
nand U250 (N_250,In_105,In_18);
or U251 (N_251,In_251,In_481);
or U252 (N_252,In_301,In_338);
or U253 (N_253,In_63,In_380);
and U254 (N_254,In_454,In_128);
and U255 (N_255,In_357,In_232);
and U256 (N_256,In_438,In_2);
or U257 (N_257,In_453,In_182);
and U258 (N_258,In_89,In_419);
nor U259 (N_259,In_254,In_316);
and U260 (N_260,In_117,In_68);
nor U261 (N_261,In_124,In_425);
nor U262 (N_262,In_165,In_493);
and U263 (N_263,In_93,In_419);
and U264 (N_264,In_417,In_332);
nor U265 (N_265,In_232,In_46);
nor U266 (N_266,In_371,In_295);
nand U267 (N_267,In_383,In_410);
or U268 (N_268,In_177,In_28);
and U269 (N_269,In_24,In_31);
nand U270 (N_270,In_59,In_127);
nor U271 (N_271,In_398,In_388);
nand U272 (N_272,In_398,In_399);
or U273 (N_273,In_233,In_462);
nor U274 (N_274,In_493,In_457);
nor U275 (N_275,In_48,In_230);
xor U276 (N_276,In_337,In_245);
or U277 (N_277,In_493,In_446);
or U278 (N_278,In_186,In_465);
or U279 (N_279,In_218,In_231);
nand U280 (N_280,In_478,In_95);
xor U281 (N_281,In_243,In_497);
nor U282 (N_282,In_2,In_440);
nand U283 (N_283,In_1,In_99);
or U284 (N_284,In_471,In_371);
nor U285 (N_285,In_438,In_451);
nand U286 (N_286,In_22,In_24);
or U287 (N_287,In_389,In_70);
nor U288 (N_288,In_199,In_412);
or U289 (N_289,In_313,In_55);
nor U290 (N_290,In_155,In_68);
nor U291 (N_291,In_420,In_361);
xor U292 (N_292,In_204,In_200);
nand U293 (N_293,In_437,In_171);
nor U294 (N_294,In_373,In_323);
nand U295 (N_295,In_54,In_314);
or U296 (N_296,In_90,In_325);
and U297 (N_297,In_166,In_89);
or U298 (N_298,In_138,In_238);
or U299 (N_299,In_306,In_495);
nor U300 (N_300,In_0,In_131);
and U301 (N_301,In_393,In_450);
xnor U302 (N_302,In_157,In_407);
nand U303 (N_303,In_437,In_102);
nor U304 (N_304,In_185,In_304);
or U305 (N_305,In_473,In_12);
and U306 (N_306,In_261,In_11);
nor U307 (N_307,In_130,In_5);
nand U308 (N_308,In_253,In_78);
nor U309 (N_309,In_148,In_298);
nand U310 (N_310,In_308,In_359);
nor U311 (N_311,In_35,In_231);
nand U312 (N_312,In_353,In_411);
or U313 (N_313,In_3,In_8);
or U314 (N_314,In_479,In_487);
and U315 (N_315,In_248,In_269);
nand U316 (N_316,In_420,In_159);
xnor U317 (N_317,In_305,In_82);
nand U318 (N_318,In_38,In_458);
nor U319 (N_319,In_454,In_148);
xor U320 (N_320,In_236,In_66);
nor U321 (N_321,In_97,In_17);
xor U322 (N_322,In_145,In_273);
and U323 (N_323,In_259,In_316);
nand U324 (N_324,In_406,In_428);
xor U325 (N_325,In_469,In_459);
and U326 (N_326,In_275,In_320);
nand U327 (N_327,In_210,In_450);
nor U328 (N_328,In_390,In_429);
nor U329 (N_329,In_5,In_212);
and U330 (N_330,In_264,In_54);
and U331 (N_331,In_178,In_265);
xnor U332 (N_332,In_93,In_14);
nor U333 (N_333,In_83,In_320);
nand U334 (N_334,In_475,In_436);
and U335 (N_335,In_19,In_143);
nor U336 (N_336,In_206,In_387);
or U337 (N_337,In_44,In_304);
nand U338 (N_338,In_382,In_85);
nor U339 (N_339,In_39,In_438);
or U340 (N_340,In_377,In_280);
or U341 (N_341,In_74,In_21);
or U342 (N_342,In_492,In_153);
xor U343 (N_343,In_493,In_324);
nor U344 (N_344,In_240,In_26);
nand U345 (N_345,In_418,In_88);
nor U346 (N_346,In_331,In_234);
or U347 (N_347,In_404,In_342);
nor U348 (N_348,In_354,In_371);
nand U349 (N_349,In_318,In_450);
and U350 (N_350,In_92,In_342);
or U351 (N_351,In_281,In_21);
nand U352 (N_352,In_35,In_459);
and U353 (N_353,In_403,In_201);
xor U354 (N_354,In_454,In_295);
and U355 (N_355,In_356,In_94);
or U356 (N_356,In_491,In_391);
xnor U357 (N_357,In_144,In_270);
and U358 (N_358,In_398,In_310);
nand U359 (N_359,In_277,In_86);
nor U360 (N_360,In_172,In_493);
nand U361 (N_361,In_286,In_380);
nor U362 (N_362,In_35,In_115);
nor U363 (N_363,In_315,In_458);
and U364 (N_364,In_136,In_255);
and U365 (N_365,In_297,In_138);
or U366 (N_366,In_380,In_108);
and U367 (N_367,In_175,In_126);
nand U368 (N_368,In_67,In_218);
nor U369 (N_369,In_131,In_21);
or U370 (N_370,In_178,In_359);
nand U371 (N_371,In_305,In_362);
and U372 (N_372,In_448,In_70);
nand U373 (N_373,In_37,In_358);
and U374 (N_374,In_269,In_70);
nor U375 (N_375,In_462,In_102);
nand U376 (N_376,In_338,In_40);
and U377 (N_377,In_381,In_309);
nand U378 (N_378,In_364,In_61);
nor U379 (N_379,In_229,In_421);
nand U380 (N_380,In_296,In_123);
nor U381 (N_381,In_416,In_64);
nor U382 (N_382,In_88,In_244);
nor U383 (N_383,In_18,In_52);
or U384 (N_384,In_488,In_335);
and U385 (N_385,In_275,In_47);
nor U386 (N_386,In_486,In_230);
nand U387 (N_387,In_411,In_92);
nor U388 (N_388,In_205,In_264);
nor U389 (N_389,In_286,In_275);
nand U390 (N_390,In_269,In_128);
and U391 (N_391,In_124,In_452);
nand U392 (N_392,In_439,In_257);
nor U393 (N_393,In_19,In_388);
or U394 (N_394,In_39,In_445);
nor U395 (N_395,In_230,In_130);
or U396 (N_396,In_399,In_29);
nor U397 (N_397,In_498,In_412);
nand U398 (N_398,In_394,In_23);
xnor U399 (N_399,In_141,In_146);
nor U400 (N_400,In_308,In_213);
and U401 (N_401,In_167,In_254);
or U402 (N_402,In_310,In_256);
nor U403 (N_403,In_376,In_453);
nor U404 (N_404,In_410,In_319);
nor U405 (N_405,In_280,In_417);
or U406 (N_406,In_175,In_25);
nand U407 (N_407,In_115,In_418);
or U408 (N_408,In_126,In_316);
or U409 (N_409,In_428,In_239);
and U410 (N_410,In_280,In_324);
or U411 (N_411,In_195,In_448);
or U412 (N_412,In_99,In_195);
and U413 (N_413,In_234,In_28);
nor U414 (N_414,In_331,In_145);
or U415 (N_415,In_22,In_328);
nand U416 (N_416,In_351,In_375);
nand U417 (N_417,In_293,In_315);
or U418 (N_418,In_64,In_441);
nand U419 (N_419,In_207,In_143);
or U420 (N_420,In_213,In_380);
nor U421 (N_421,In_176,In_451);
nor U422 (N_422,In_256,In_377);
and U423 (N_423,In_100,In_73);
nand U424 (N_424,In_479,In_363);
nand U425 (N_425,In_22,In_441);
nor U426 (N_426,In_59,In_331);
nand U427 (N_427,In_439,In_228);
xor U428 (N_428,In_434,In_306);
or U429 (N_429,In_422,In_458);
nor U430 (N_430,In_170,In_68);
or U431 (N_431,In_255,In_110);
or U432 (N_432,In_386,In_329);
and U433 (N_433,In_330,In_229);
and U434 (N_434,In_179,In_144);
or U435 (N_435,In_150,In_189);
nand U436 (N_436,In_283,In_203);
and U437 (N_437,In_337,In_496);
or U438 (N_438,In_386,In_390);
xor U439 (N_439,In_42,In_287);
or U440 (N_440,In_216,In_469);
nor U441 (N_441,In_203,In_427);
nor U442 (N_442,In_250,In_436);
nand U443 (N_443,In_135,In_207);
xnor U444 (N_444,In_123,In_498);
nor U445 (N_445,In_381,In_42);
nor U446 (N_446,In_21,In_351);
nand U447 (N_447,In_346,In_236);
or U448 (N_448,In_103,In_431);
and U449 (N_449,In_430,In_243);
and U450 (N_450,In_457,In_376);
nand U451 (N_451,In_125,In_321);
or U452 (N_452,In_330,In_255);
nor U453 (N_453,In_417,In_297);
nor U454 (N_454,In_203,In_431);
xor U455 (N_455,In_173,In_4);
or U456 (N_456,In_293,In_85);
and U457 (N_457,In_258,In_307);
and U458 (N_458,In_162,In_30);
or U459 (N_459,In_333,In_65);
nor U460 (N_460,In_69,In_404);
and U461 (N_461,In_278,In_400);
or U462 (N_462,In_386,In_135);
nor U463 (N_463,In_324,In_67);
nor U464 (N_464,In_449,In_126);
xor U465 (N_465,In_152,In_400);
and U466 (N_466,In_195,In_96);
nor U467 (N_467,In_465,In_2);
and U468 (N_468,In_109,In_467);
nor U469 (N_469,In_462,In_2);
nor U470 (N_470,In_294,In_68);
nand U471 (N_471,In_384,In_163);
xnor U472 (N_472,In_276,In_294);
and U473 (N_473,In_90,In_465);
and U474 (N_474,In_300,In_265);
nand U475 (N_475,In_156,In_401);
nor U476 (N_476,In_459,In_89);
and U477 (N_477,In_448,In_444);
nand U478 (N_478,In_126,In_154);
and U479 (N_479,In_157,In_68);
and U480 (N_480,In_399,In_194);
xnor U481 (N_481,In_284,In_183);
or U482 (N_482,In_260,In_32);
nand U483 (N_483,In_388,In_384);
nand U484 (N_484,In_101,In_469);
nor U485 (N_485,In_152,In_47);
or U486 (N_486,In_427,In_59);
and U487 (N_487,In_187,In_190);
and U488 (N_488,In_220,In_159);
nand U489 (N_489,In_465,In_185);
xor U490 (N_490,In_234,In_143);
and U491 (N_491,In_435,In_281);
and U492 (N_492,In_313,In_388);
or U493 (N_493,In_131,In_449);
and U494 (N_494,In_346,In_219);
and U495 (N_495,In_163,In_494);
nor U496 (N_496,In_409,In_13);
or U497 (N_497,In_480,In_155);
nand U498 (N_498,In_407,In_63);
nor U499 (N_499,In_487,In_275);
nand U500 (N_500,N_219,N_38);
and U501 (N_501,N_37,N_132);
nor U502 (N_502,N_251,N_53);
and U503 (N_503,N_294,N_307);
xor U504 (N_504,N_310,N_372);
and U505 (N_505,N_325,N_94);
or U506 (N_506,N_292,N_123);
xor U507 (N_507,N_249,N_150);
or U508 (N_508,N_342,N_341);
or U509 (N_509,N_92,N_468);
and U510 (N_510,N_184,N_74);
and U511 (N_511,N_466,N_269);
nand U512 (N_512,N_234,N_409);
nand U513 (N_513,N_240,N_474);
nand U514 (N_514,N_424,N_289);
nor U515 (N_515,N_161,N_496);
or U516 (N_516,N_298,N_222);
and U517 (N_517,N_323,N_336);
and U518 (N_518,N_112,N_202);
or U519 (N_519,N_290,N_483);
or U520 (N_520,N_41,N_369);
nor U521 (N_521,N_394,N_319);
and U522 (N_522,N_238,N_439);
nand U523 (N_523,N_295,N_475);
and U524 (N_524,N_371,N_355);
and U525 (N_525,N_0,N_271);
or U526 (N_526,N_177,N_126);
nor U527 (N_527,N_199,N_429);
nor U528 (N_528,N_340,N_125);
and U529 (N_529,N_55,N_183);
xnor U530 (N_530,N_337,N_284);
nand U531 (N_531,N_406,N_430);
nor U532 (N_532,N_343,N_314);
nand U533 (N_533,N_34,N_418);
or U534 (N_534,N_90,N_257);
nand U535 (N_535,N_487,N_435);
xnor U536 (N_536,N_356,N_423);
and U537 (N_537,N_347,N_27);
and U538 (N_538,N_171,N_130);
and U539 (N_539,N_272,N_277);
nor U540 (N_540,N_111,N_331);
and U541 (N_541,N_84,N_388);
nor U542 (N_542,N_247,N_65);
or U543 (N_543,N_172,N_66);
and U544 (N_544,N_89,N_116);
nand U545 (N_545,N_207,N_100);
and U546 (N_546,N_281,N_450);
nand U547 (N_547,N_252,N_210);
xor U548 (N_548,N_73,N_72);
nor U549 (N_549,N_164,N_11);
nand U550 (N_550,N_114,N_485);
nor U551 (N_551,N_478,N_137);
or U552 (N_552,N_245,N_267);
nor U553 (N_553,N_157,N_415);
nand U554 (N_554,N_278,N_120);
and U555 (N_555,N_254,N_127);
nand U556 (N_556,N_235,N_302);
or U557 (N_557,N_448,N_459);
xnor U558 (N_558,N_462,N_358);
and U559 (N_559,N_231,N_160);
nor U560 (N_560,N_316,N_133);
or U561 (N_561,N_64,N_403);
and U562 (N_562,N_486,N_497);
and U563 (N_563,N_33,N_259);
or U564 (N_564,N_70,N_43);
and U565 (N_565,N_383,N_451);
nand U566 (N_566,N_62,N_276);
nand U567 (N_567,N_168,N_54);
nand U568 (N_568,N_421,N_155);
and U569 (N_569,N_106,N_83);
and U570 (N_570,N_149,N_320);
nand U571 (N_571,N_283,N_365);
or U572 (N_572,N_442,N_56);
or U573 (N_573,N_99,N_140);
nand U574 (N_574,N_334,N_373);
nand U575 (N_575,N_456,N_328);
nor U576 (N_576,N_274,N_102);
and U577 (N_577,N_344,N_351);
nand U578 (N_578,N_236,N_44);
nand U579 (N_579,N_174,N_194);
nand U580 (N_580,N_255,N_443);
nor U581 (N_581,N_198,N_395);
nor U582 (N_582,N_285,N_22);
and U583 (N_583,N_4,N_10);
nor U584 (N_584,N_154,N_213);
and U585 (N_585,N_63,N_107);
or U586 (N_586,N_303,N_218);
or U587 (N_587,N_364,N_482);
or U588 (N_588,N_384,N_189);
or U589 (N_589,N_117,N_408);
and U590 (N_590,N_7,N_472);
xnor U591 (N_591,N_441,N_42);
nand U592 (N_592,N_329,N_492);
and U593 (N_593,N_119,N_413);
nor U594 (N_594,N_146,N_346);
and U595 (N_595,N_363,N_221);
nand U596 (N_596,N_477,N_412);
and U597 (N_597,N_118,N_368);
and U598 (N_598,N_258,N_246);
nor U599 (N_599,N_81,N_124);
or U600 (N_600,N_353,N_170);
or U601 (N_601,N_498,N_152);
and U602 (N_602,N_345,N_77);
nor U603 (N_603,N_489,N_359);
nor U604 (N_604,N_85,N_61);
and U605 (N_605,N_280,N_2);
nand U606 (N_606,N_244,N_312);
nor U607 (N_607,N_349,N_232);
or U608 (N_608,N_265,N_82);
nand U609 (N_609,N_391,N_392);
or U610 (N_610,N_287,N_301);
nor U611 (N_611,N_420,N_299);
nor U612 (N_612,N_321,N_432);
nor U613 (N_613,N_217,N_490);
and U614 (N_614,N_187,N_122);
nand U615 (N_615,N_262,N_227);
or U616 (N_616,N_402,N_93);
nand U617 (N_617,N_317,N_288);
and U618 (N_618,N_370,N_204);
or U619 (N_619,N_291,N_398);
nand U620 (N_620,N_458,N_109);
nor U621 (N_621,N_19,N_333);
and U622 (N_622,N_181,N_438);
nor U623 (N_623,N_239,N_385);
and U624 (N_624,N_98,N_326);
nor U625 (N_625,N_382,N_476);
nor U626 (N_626,N_223,N_248);
xor U627 (N_627,N_226,N_79);
nand U628 (N_628,N_381,N_87);
or U629 (N_629,N_159,N_444);
nand U630 (N_630,N_49,N_148);
nand U631 (N_631,N_129,N_454);
or U632 (N_632,N_266,N_484);
or U633 (N_633,N_179,N_209);
nor U634 (N_634,N_455,N_163);
or U635 (N_635,N_305,N_36);
xnor U636 (N_636,N_12,N_110);
or U637 (N_637,N_339,N_216);
nor U638 (N_638,N_224,N_225);
and U639 (N_639,N_135,N_88);
nand U640 (N_640,N_243,N_479);
nand U641 (N_641,N_354,N_367);
nand U642 (N_642,N_52,N_306);
nor U643 (N_643,N_16,N_230);
and U644 (N_644,N_495,N_350);
or U645 (N_645,N_68,N_147);
and U646 (N_646,N_101,N_446);
and U647 (N_647,N_39,N_440);
nor U648 (N_648,N_193,N_237);
nand U649 (N_649,N_215,N_461);
and U650 (N_650,N_3,N_15);
and U651 (N_651,N_208,N_115);
nor U652 (N_652,N_390,N_95);
nor U653 (N_653,N_268,N_396);
nor U654 (N_654,N_315,N_96);
and U655 (N_655,N_410,N_141);
nor U656 (N_656,N_182,N_51);
and U657 (N_657,N_58,N_180);
or U658 (N_658,N_48,N_309);
or U659 (N_659,N_104,N_434);
nand U660 (N_660,N_414,N_300);
xor U661 (N_661,N_40,N_436);
and U662 (N_662,N_233,N_205);
or U663 (N_663,N_499,N_293);
xor U664 (N_664,N_488,N_286);
nor U665 (N_665,N_206,N_6);
nand U666 (N_666,N_360,N_151);
or U667 (N_667,N_464,N_50);
nand U668 (N_668,N_5,N_375);
or U669 (N_669,N_256,N_433);
and U670 (N_670,N_361,N_178);
nand U671 (N_671,N_393,N_9);
nand U672 (N_672,N_47,N_428);
nor U673 (N_673,N_203,N_445);
or U674 (N_674,N_453,N_228);
and U675 (N_675,N_18,N_437);
and U676 (N_676,N_380,N_404);
and U677 (N_677,N_220,N_481);
nor U678 (N_678,N_308,N_399);
nor U679 (N_679,N_400,N_91);
and U680 (N_680,N_175,N_211);
and U681 (N_681,N_447,N_405);
nor U682 (N_682,N_145,N_327);
nor U683 (N_683,N_431,N_452);
nand U684 (N_684,N_214,N_416);
xor U685 (N_685,N_57,N_457);
and U686 (N_686,N_425,N_78);
and U687 (N_687,N_261,N_167);
nor U688 (N_688,N_318,N_142);
or U689 (N_689,N_279,N_23);
and U690 (N_690,N_494,N_35);
nand U691 (N_691,N_80,N_465);
and U692 (N_692,N_196,N_176);
and U693 (N_693,N_463,N_190);
or U694 (N_694,N_469,N_378);
nand U695 (N_695,N_185,N_24);
xnor U696 (N_696,N_426,N_26);
and U697 (N_697,N_297,N_67);
xor U698 (N_698,N_97,N_21);
and U699 (N_699,N_379,N_173);
and U700 (N_700,N_60,N_470);
or U701 (N_701,N_338,N_275);
nor U702 (N_702,N_330,N_45);
nor U703 (N_703,N_491,N_69);
nand U704 (N_704,N_144,N_14);
or U705 (N_705,N_260,N_270);
and U706 (N_706,N_407,N_195);
and U707 (N_707,N_422,N_108);
and U708 (N_708,N_139,N_471);
xor U709 (N_709,N_138,N_1);
nand U710 (N_710,N_201,N_158);
nand U711 (N_711,N_17,N_480);
xor U712 (N_712,N_493,N_313);
or U713 (N_713,N_162,N_20);
or U714 (N_714,N_186,N_212);
and U715 (N_715,N_30,N_401);
or U716 (N_716,N_25,N_31);
or U717 (N_717,N_322,N_417);
and U718 (N_718,N_153,N_134);
or U719 (N_719,N_13,N_348);
nor U720 (N_720,N_143,N_131);
and U721 (N_721,N_86,N_188);
nand U722 (N_722,N_169,N_282);
and U723 (N_723,N_387,N_229);
nand U724 (N_724,N_264,N_165);
nor U725 (N_725,N_166,N_377);
xor U726 (N_726,N_427,N_263);
nand U727 (N_727,N_8,N_376);
and U728 (N_728,N_473,N_156);
and U729 (N_729,N_352,N_128);
nor U730 (N_730,N_103,N_191);
nor U731 (N_731,N_335,N_242);
and U732 (N_732,N_374,N_273);
nor U733 (N_733,N_366,N_311);
and U734 (N_734,N_332,N_357);
nand U735 (N_735,N_253,N_449);
nor U736 (N_736,N_411,N_241);
and U737 (N_737,N_75,N_467);
nor U738 (N_738,N_29,N_121);
or U739 (N_739,N_397,N_460);
or U740 (N_740,N_386,N_200);
nand U741 (N_741,N_113,N_59);
nand U742 (N_742,N_32,N_250);
nor U743 (N_743,N_46,N_76);
nand U744 (N_744,N_389,N_197);
nor U745 (N_745,N_362,N_304);
or U746 (N_746,N_296,N_105);
nand U747 (N_747,N_324,N_28);
or U748 (N_748,N_136,N_419);
and U749 (N_749,N_192,N_71);
xnor U750 (N_750,N_421,N_146);
or U751 (N_751,N_337,N_392);
and U752 (N_752,N_153,N_135);
nand U753 (N_753,N_443,N_379);
and U754 (N_754,N_445,N_462);
nor U755 (N_755,N_240,N_46);
or U756 (N_756,N_37,N_155);
or U757 (N_757,N_15,N_7);
nor U758 (N_758,N_265,N_239);
and U759 (N_759,N_341,N_370);
and U760 (N_760,N_15,N_4);
nor U761 (N_761,N_118,N_418);
nand U762 (N_762,N_41,N_155);
nor U763 (N_763,N_88,N_38);
xor U764 (N_764,N_146,N_163);
nand U765 (N_765,N_45,N_253);
nand U766 (N_766,N_365,N_96);
nand U767 (N_767,N_299,N_383);
nand U768 (N_768,N_306,N_443);
nand U769 (N_769,N_81,N_375);
nand U770 (N_770,N_14,N_324);
xnor U771 (N_771,N_285,N_106);
nor U772 (N_772,N_458,N_407);
and U773 (N_773,N_149,N_29);
nand U774 (N_774,N_356,N_251);
and U775 (N_775,N_460,N_58);
and U776 (N_776,N_178,N_68);
nor U777 (N_777,N_345,N_346);
and U778 (N_778,N_481,N_476);
or U779 (N_779,N_190,N_363);
nand U780 (N_780,N_393,N_357);
and U781 (N_781,N_53,N_361);
and U782 (N_782,N_222,N_179);
nor U783 (N_783,N_356,N_11);
or U784 (N_784,N_357,N_414);
and U785 (N_785,N_314,N_497);
and U786 (N_786,N_149,N_194);
or U787 (N_787,N_232,N_353);
or U788 (N_788,N_332,N_408);
xnor U789 (N_789,N_89,N_190);
or U790 (N_790,N_9,N_165);
nand U791 (N_791,N_202,N_123);
xnor U792 (N_792,N_373,N_325);
nor U793 (N_793,N_451,N_319);
nand U794 (N_794,N_257,N_490);
nand U795 (N_795,N_320,N_499);
nand U796 (N_796,N_156,N_179);
and U797 (N_797,N_449,N_435);
nor U798 (N_798,N_3,N_236);
or U799 (N_799,N_378,N_451);
or U800 (N_800,N_313,N_331);
nor U801 (N_801,N_314,N_67);
and U802 (N_802,N_458,N_16);
or U803 (N_803,N_452,N_124);
and U804 (N_804,N_429,N_417);
and U805 (N_805,N_237,N_121);
nor U806 (N_806,N_61,N_192);
or U807 (N_807,N_175,N_404);
nor U808 (N_808,N_458,N_262);
and U809 (N_809,N_229,N_126);
nor U810 (N_810,N_169,N_255);
or U811 (N_811,N_290,N_115);
nor U812 (N_812,N_149,N_424);
xnor U813 (N_813,N_87,N_424);
nor U814 (N_814,N_257,N_121);
nand U815 (N_815,N_351,N_65);
and U816 (N_816,N_407,N_275);
nor U817 (N_817,N_45,N_148);
or U818 (N_818,N_384,N_469);
and U819 (N_819,N_101,N_200);
nand U820 (N_820,N_268,N_93);
and U821 (N_821,N_495,N_10);
nor U822 (N_822,N_285,N_134);
and U823 (N_823,N_211,N_389);
and U824 (N_824,N_410,N_264);
nand U825 (N_825,N_215,N_336);
nor U826 (N_826,N_246,N_75);
xor U827 (N_827,N_253,N_148);
nor U828 (N_828,N_381,N_138);
xor U829 (N_829,N_185,N_67);
nand U830 (N_830,N_202,N_151);
nand U831 (N_831,N_94,N_393);
and U832 (N_832,N_293,N_67);
nor U833 (N_833,N_495,N_20);
xnor U834 (N_834,N_39,N_378);
nor U835 (N_835,N_317,N_155);
or U836 (N_836,N_166,N_314);
nand U837 (N_837,N_453,N_182);
nor U838 (N_838,N_135,N_99);
and U839 (N_839,N_244,N_133);
nand U840 (N_840,N_50,N_54);
nor U841 (N_841,N_68,N_34);
nand U842 (N_842,N_219,N_231);
and U843 (N_843,N_68,N_51);
or U844 (N_844,N_99,N_479);
nor U845 (N_845,N_195,N_498);
or U846 (N_846,N_341,N_486);
or U847 (N_847,N_209,N_108);
nand U848 (N_848,N_416,N_11);
and U849 (N_849,N_268,N_204);
nor U850 (N_850,N_454,N_327);
and U851 (N_851,N_262,N_382);
or U852 (N_852,N_272,N_72);
xor U853 (N_853,N_479,N_95);
nor U854 (N_854,N_498,N_11);
nor U855 (N_855,N_450,N_284);
nand U856 (N_856,N_341,N_464);
nand U857 (N_857,N_197,N_401);
nor U858 (N_858,N_365,N_487);
xnor U859 (N_859,N_311,N_264);
and U860 (N_860,N_15,N_207);
xor U861 (N_861,N_107,N_305);
and U862 (N_862,N_6,N_411);
nand U863 (N_863,N_154,N_374);
nor U864 (N_864,N_338,N_244);
or U865 (N_865,N_403,N_336);
nand U866 (N_866,N_36,N_168);
and U867 (N_867,N_91,N_411);
nor U868 (N_868,N_43,N_133);
nand U869 (N_869,N_67,N_154);
and U870 (N_870,N_8,N_317);
nand U871 (N_871,N_484,N_311);
xor U872 (N_872,N_165,N_20);
and U873 (N_873,N_163,N_195);
or U874 (N_874,N_475,N_456);
nor U875 (N_875,N_156,N_248);
nand U876 (N_876,N_46,N_439);
nand U877 (N_877,N_57,N_232);
nor U878 (N_878,N_189,N_40);
and U879 (N_879,N_220,N_163);
nand U880 (N_880,N_354,N_175);
and U881 (N_881,N_97,N_70);
nor U882 (N_882,N_240,N_35);
nand U883 (N_883,N_257,N_115);
and U884 (N_884,N_170,N_157);
nand U885 (N_885,N_405,N_414);
nor U886 (N_886,N_140,N_341);
and U887 (N_887,N_354,N_302);
or U888 (N_888,N_396,N_378);
nand U889 (N_889,N_45,N_355);
xnor U890 (N_890,N_23,N_426);
and U891 (N_891,N_292,N_213);
nor U892 (N_892,N_424,N_483);
or U893 (N_893,N_465,N_129);
nand U894 (N_894,N_108,N_311);
nor U895 (N_895,N_286,N_44);
and U896 (N_896,N_282,N_217);
and U897 (N_897,N_493,N_404);
or U898 (N_898,N_386,N_158);
and U899 (N_899,N_18,N_101);
nor U900 (N_900,N_14,N_308);
or U901 (N_901,N_145,N_277);
or U902 (N_902,N_473,N_208);
nand U903 (N_903,N_232,N_66);
and U904 (N_904,N_456,N_193);
nor U905 (N_905,N_422,N_391);
nor U906 (N_906,N_59,N_215);
or U907 (N_907,N_484,N_102);
xnor U908 (N_908,N_443,N_295);
or U909 (N_909,N_6,N_217);
or U910 (N_910,N_237,N_153);
xor U911 (N_911,N_68,N_405);
nand U912 (N_912,N_363,N_256);
and U913 (N_913,N_217,N_487);
and U914 (N_914,N_302,N_43);
nand U915 (N_915,N_304,N_431);
nand U916 (N_916,N_378,N_348);
and U917 (N_917,N_214,N_301);
nor U918 (N_918,N_171,N_380);
or U919 (N_919,N_92,N_401);
nand U920 (N_920,N_155,N_328);
or U921 (N_921,N_61,N_129);
nand U922 (N_922,N_71,N_261);
nand U923 (N_923,N_54,N_370);
nor U924 (N_924,N_337,N_76);
nor U925 (N_925,N_320,N_387);
and U926 (N_926,N_172,N_147);
or U927 (N_927,N_61,N_496);
and U928 (N_928,N_114,N_52);
nor U929 (N_929,N_261,N_66);
nand U930 (N_930,N_414,N_412);
nand U931 (N_931,N_77,N_93);
or U932 (N_932,N_347,N_320);
and U933 (N_933,N_232,N_9);
nand U934 (N_934,N_444,N_450);
or U935 (N_935,N_284,N_262);
nand U936 (N_936,N_305,N_139);
or U937 (N_937,N_135,N_326);
nor U938 (N_938,N_376,N_159);
nand U939 (N_939,N_250,N_142);
and U940 (N_940,N_90,N_335);
or U941 (N_941,N_140,N_86);
nor U942 (N_942,N_127,N_245);
or U943 (N_943,N_154,N_113);
nor U944 (N_944,N_393,N_38);
or U945 (N_945,N_281,N_262);
xor U946 (N_946,N_196,N_44);
nor U947 (N_947,N_497,N_177);
nand U948 (N_948,N_498,N_104);
xor U949 (N_949,N_245,N_201);
and U950 (N_950,N_396,N_214);
and U951 (N_951,N_250,N_327);
nor U952 (N_952,N_263,N_264);
or U953 (N_953,N_341,N_442);
nand U954 (N_954,N_168,N_405);
nor U955 (N_955,N_112,N_192);
and U956 (N_956,N_120,N_97);
nor U957 (N_957,N_448,N_23);
or U958 (N_958,N_465,N_381);
and U959 (N_959,N_59,N_62);
nor U960 (N_960,N_34,N_142);
nor U961 (N_961,N_346,N_213);
nand U962 (N_962,N_437,N_290);
nor U963 (N_963,N_34,N_277);
and U964 (N_964,N_162,N_238);
and U965 (N_965,N_401,N_461);
nand U966 (N_966,N_459,N_98);
or U967 (N_967,N_65,N_436);
or U968 (N_968,N_39,N_468);
nor U969 (N_969,N_382,N_172);
or U970 (N_970,N_260,N_117);
xnor U971 (N_971,N_51,N_168);
nand U972 (N_972,N_445,N_439);
nor U973 (N_973,N_493,N_220);
and U974 (N_974,N_402,N_128);
nand U975 (N_975,N_392,N_377);
nor U976 (N_976,N_166,N_34);
nand U977 (N_977,N_89,N_12);
nand U978 (N_978,N_377,N_347);
xnor U979 (N_979,N_59,N_347);
nor U980 (N_980,N_364,N_80);
and U981 (N_981,N_60,N_140);
or U982 (N_982,N_256,N_132);
nor U983 (N_983,N_378,N_444);
xnor U984 (N_984,N_318,N_149);
nand U985 (N_985,N_350,N_431);
xor U986 (N_986,N_145,N_499);
and U987 (N_987,N_354,N_319);
and U988 (N_988,N_20,N_410);
and U989 (N_989,N_457,N_361);
nand U990 (N_990,N_42,N_322);
nor U991 (N_991,N_378,N_236);
nor U992 (N_992,N_419,N_113);
nor U993 (N_993,N_93,N_432);
nor U994 (N_994,N_0,N_256);
nand U995 (N_995,N_38,N_239);
and U996 (N_996,N_229,N_285);
or U997 (N_997,N_181,N_450);
and U998 (N_998,N_259,N_184);
and U999 (N_999,N_13,N_110);
xnor U1000 (N_1000,N_591,N_722);
and U1001 (N_1001,N_980,N_706);
nor U1002 (N_1002,N_903,N_547);
and U1003 (N_1003,N_877,N_901);
nand U1004 (N_1004,N_569,N_508);
nor U1005 (N_1005,N_866,N_767);
nand U1006 (N_1006,N_509,N_935);
nand U1007 (N_1007,N_904,N_926);
xnor U1008 (N_1008,N_671,N_654);
nor U1009 (N_1009,N_518,N_691);
nand U1010 (N_1010,N_517,N_515);
or U1011 (N_1011,N_557,N_962);
nor U1012 (N_1012,N_886,N_910);
or U1013 (N_1013,N_727,N_735);
nand U1014 (N_1014,N_564,N_530);
nand U1015 (N_1015,N_775,N_837);
nor U1016 (N_1016,N_666,N_682);
nand U1017 (N_1017,N_617,N_719);
nor U1018 (N_1018,N_818,N_835);
or U1019 (N_1019,N_634,N_716);
nand U1020 (N_1020,N_810,N_754);
or U1021 (N_1021,N_848,N_705);
nand U1022 (N_1022,N_804,N_858);
nor U1023 (N_1023,N_713,N_536);
or U1024 (N_1024,N_884,N_918);
nand U1025 (N_1025,N_825,N_867);
and U1026 (N_1026,N_865,N_681);
nand U1027 (N_1027,N_768,N_791);
or U1028 (N_1028,N_966,N_795);
nor U1029 (N_1029,N_685,N_802);
or U1030 (N_1030,N_813,N_953);
and U1031 (N_1031,N_940,N_951);
and U1032 (N_1032,N_743,N_650);
nand U1033 (N_1033,N_830,N_657);
or U1034 (N_1034,N_834,N_897);
and U1035 (N_1035,N_733,N_533);
nor U1036 (N_1036,N_799,N_624);
nand U1037 (N_1037,N_637,N_573);
and U1038 (N_1038,N_552,N_783);
or U1039 (N_1039,N_970,N_581);
nor U1040 (N_1040,N_724,N_506);
and U1041 (N_1041,N_781,N_700);
nor U1042 (N_1042,N_527,N_586);
or U1043 (N_1043,N_758,N_572);
nand U1044 (N_1044,N_669,N_869);
nor U1045 (N_1045,N_973,N_680);
nor U1046 (N_1046,N_687,N_971);
or U1047 (N_1047,N_765,N_964);
nand U1048 (N_1048,N_792,N_568);
or U1049 (N_1049,N_729,N_675);
nor U1050 (N_1050,N_892,N_651);
nor U1051 (N_1051,N_546,N_839);
and U1052 (N_1052,N_954,N_645);
and U1053 (N_1053,N_526,N_927);
nand U1054 (N_1054,N_598,N_847);
nand U1055 (N_1055,N_542,N_749);
or U1056 (N_1056,N_993,N_959);
nand U1057 (N_1057,N_592,N_896);
or U1058 (N_1058,N_872,N_704);
and U1059 (N_1059,N_678,N_823);
nand U1060 (N_1060,N_524,N_965);
and U1061 (N_1061,N_659,N_602);
nand U1062 (N_1062,N_882,N_701);
and U1063 (N_1063,N_836,N_832);
nand U1064 (N_1064,N_922,N_957);
or U1065 (N_1065,N_528,N_694);
nor U1066 (N_1066,N_764,N_779);
xnor U1067 (N_1067,N_516,N_871);
and U1068 (N_1068,N_730,N_788);
nor U1069 (N_1069,N_560,N_899);
or U1070 (N_1070,N_519,N_614);
or U1071 (N_1071,N_889,N_909);
nor U1072 (N_1072,N_511,N_874);
xnor U1073 (N_1073,N_587,N_797);
and U1074 (N_1074,N_679,N_913);
or U1075 (N_1075,N_851,N_961);
nand U1076 (N_1076,N_597,N_761);
and U1077 (N_1077,N_611,N_539);
or U1078 (N_1078,N_820,N_950);
or U1079 (N_1079,N_814,N_708);
or U1080 (N_1080,N_649,N_714);
and U1081 (N_1081,N_610,N_693);
nor U1082 (N_1082,N_898,N_696);
or U1083 (N_1083,N_990,N_766);
nor U1084 (N_1084,N_929,N_646);
nor U1085 (N_1085,N_987,N_821);
xor U1086 (N_1086,N_686,N_751);
and U1087 (N_1087,N_933,N_510);
and U1088 (N_1088,N_500,N_626);
nand U1089 (N_1089,N_878,N_692);
or U1090 (N_1090,N_908,N_969);
nor U1091 (N_1091,N_502,N_535);
nor U1092 (N_1092,N_930,N_842);
nand U1093 (N_1093,N_523,N_702);
nor U1094 (N_1094,N_759,N_576);
and U1095 (N_1095,N_653,N_777);
or U1096 (N_1096,N_603,N_566);
or U1097 (N_1097,N_589,N_710);
xor U1098 (N_1098,N_997,N_999);
nor U1099 (N_1099,N_737,N_948);
and U1100 (N_1100,N_796,N_844);
or U1101 (N_1101,N_621,N_859);
or U1102 (N_1102,N_963,N_739);
and U1103 (N_1103,N_556,N_752);
xor U1104 (N_1104,N_697,N_928);
xnor U1105 (N_1105,N_638,N_606);
nor U1106 (N_1106,N_667,N_811);
nand U1107 (N_1107,N_647,N_974);
nand U1108 (N_1108,N_562,N_563);
or U1109 (N_1109,N_545,N_805);
nor U1110 (N_1110,N_575,N_815);
xnor U1111 (N_1111,N_937,N_984);
or U1112 (N_1112,N_849,N_652);
or U1113 (N_1113,N_541,N_543);
nand U1114 (N_1114,N_828,N_833);
nand U1115 (N_1115,N_622,N_656);
nand U1116 (N_1116,N_934,N_852);
or U1117 (N_1117,N_763,N_731);
nor U1118 (N_1118,N_695,N_888);
nor U1119 (N_1119,N_967,N_944);
and U1120 (N_1120,N_827,N_721);
nand U1121 (N_1121,N_520,N_537);
or U1122 (N_1122,N_570,N_583);
or U1123 (N_1123,N_982,N_664);
nor U1124 (N_1124,N_949,N_590);
nand U1125 (N_1125,N_907,N_760);
and U1126 (N_1126,N_817,N_919);
nand U1127 (N_1127,N_931,N_941);
or U1128 (N_1128,N_529,N_550);
nor U1129 (N_1129,N_985,N_785);
xnor U1130 (N_1130,N_994,N_932);
or U1131 (N_1131,N_640,N_718);
xnor U1132 (N_1132,N_880,N_881);
and U1133 (N_1133,N_635,N_513);
or U1134 (N_1134,N_861,N_579);
nand U1135 (N_1135,N_822,N_891);
xnor U1136 (N_1136,N_643,N_553);
nand U1137 (N_1137,N_612,N_672);
and U1138 (N_1138,N_840,N_798);
nand U1139 (N_1139,N_639,N_620);
nand U1140 (N_1140,N_769,N_856);
nand U1141 (N_1141,N_806,N_846);
or U1142 (N_1142,N_914,N_829);
nand U1143 (N_1143,N_600,N_793);
nor U1144 (N_1144,N_741,N_728);
and U1145 (N_1145,N_608,N_744);
nand U1146 (N_1146,N_843,N_942);
nand U1147 (N_1147,N_633,N_831);
and U1148 (N_1148,N_561,N_955);
nor U1149 (N_1149,N_644,N_824);
nand U1150 (N_1150,N_816,N_902);
and U1151 (N_1151,N_915,N_551);
nor U1152 (N_1152,N_663,N_594);
nand U1153 (N_1153,N_558,N_544);
nor U1154 (N_1154,N_601,N_996);
nand U1155 (N_1155,N_631,N_522);
nor U1156 (N_1156,N_862,N_740);
or U1157 (N_1157,N_503,N_578);
nand U1158 (N_1158,N_890,N_947);
and U1159 (N_1159,N_770,N_660);
nand U1160 (N_1160,N_986,N_658);
nand U1161 (N_1161,N_923,N_699);
nor U1162 (N_1162,N_916,N_850);
and U1163 (N_1163,N_845,N_642);
or U1164 (N_1164,N_636,N_958);
nand U1165 (N_1165,N_812,N_826);
xor U1166 (N_1166,N_905,N_596);
and U1167 (N_1167,N_809,N_900);
and U1168 (N_1168,N_703,N_956);
or U1169 (N_1169,N_819,N_968);
or U1170 (N_1170,N_943,N_975);
nor U1171 (N_1171,N_599,N_565);
and U1172 (N_1172,N_559,N_734);
or U1173 (N_1173,N_683,N_723);
xnor U1174 (N_1174,N_738,N_906);
nand U1175 (N_1175,N_748,N_774);
xnor U1176 (N_1176,N_725,N_717);
nor U1177 (N_1177,N_661,N_938);
nand U1178 (N_1178,N_841,N_534);
and U1179 (N_1179,N_887,N_674);
xnor U1180 (N_1180,N_567,N_665);
xnor U1181 (N_1181,N_540,N_757);
xnor U1182 (N_1182,N_801,N_525);
and U1183 (N_1183,N_504,N_607);
and U1184 (N_1184,N_613,N_588);
xnor U1185 (N_1185,N_776,N_782);
nand U1186 (N_1186,N_616,N_808);
xor U1187 (N_1187,N_979,N_921);
nor U1188 (N_1188,N_641,N_689);
or U1189 (N_1189,N_627,N_623);
xor U1190 (N_1190,N_756,N_873);
and U1191 (N_1191,N_521,N_605);
nor U1192 (N_1192,N_514,N_772);
or U1193 (N_1193,N_755,N_936);
nor U1194 (N_1194,N_619,N_615);
nand U1195 (N_1195,N_800,N_911);
nor U1196 (N_1196,N_549,N_711);
nor U1197 (N_1197,N_707,N_747);
nand U1198 (N_1198,N_625,N_629);
or U1199 (N_1199,N_609,N_712);
nand U1200 (N_1200,N_585,N_628);
and U1201 (N_1201,N_532,N_574);
nand U1202 (N_1202,N_555,N_582);
nand U1203 (N_1203,N_771,N_946);
nand U1204 (N_1204,N_976,N_736);
and U1205 (N_1205,N_875,N_655);
and U1206 (N_1206,N_593,N_690);
nand U1207 (N_1207,N_732,N_720);
or U1208 (N_1208,N_981,N_577);
and U1209 (N_1209,N_726,N_854);
or U1210 (N_1210,N_920,N_879);
or U1211 (N_1211,N_715,N_784);
nand U1212 (N_1212,N_632,N_883);
nand U1213 (N_1213,N_787,N_863);
nor U1214 (N_1214,N_807,N_917);
or U1215 (N_1215,N_960,N_512);
or U1216 (N_1216,N_548,N_584);
and U1217 (N_1217,N_789,N_618);
or U1218 (N_1218,N_794,N_945);
nand U1219 (N_1219,N_885,N_668);
and U1220 (N_1220,N_753,N_648);
nand U1221 (N_1221,N_745,N_876);
nor U1222 (N_1222,N_972,N_604);
xor U1223 (N_1223,N_989,N_998);
and U1224 (N_1224,N_670,N_742);
or U1225 (N_1225,N_992,N_554);
and U1226 (N_1226,N_912,N_630);
xnor U1227 (N_1227,N_790,N_750);
nor U1228 (N_1228,N_698,N_853);
and U1229 (N_1229,N_988,N_924);
or U1230 (N_1230,N_688,N_580);
and U1231 (N_1231,N_894,N_925);
nor U1232 (N_1232,N_673,N_786);
or U1233 (N_1233,N_709,N_995);
nor U1234 (N_1234,N_952,N_864);
nand U1235 (N_1235,N_505,N_746);
and U1236 (N_1236,N_780,N_838);
nand U1237 (N_1237,N_531,N_893);
and U1238 (N_1238,N_538,N_803);
nand U1239 (N_1239,N_870,N_571);
and U1240 (N_1240,N_507,N_978);
nand U1241 (N_1241,N_778,N_857);
or U1242 (N_1242,N_501,N_662);
or U1243 (N_1243,N_762,N_895);
and U1244 (N_1244,N_677,N_684);
or U1245 (N_1245,N_977,N_595);
nor U1246 (N_1246,N_860,N_855);
nor U1247 (N_1247,N_939,N_773);
nor U1248 (N_1248,N_676,N_868);
nor U1249 (N_1249,N_983,N_991);
nand U1250 (N_1250,N_926,N_506);
nor U1251 (N_1251,N_701,N_899);
and U1252 (N_1252,N_629,N_666);
and U1253 (N_1253,N_737,N_955);
or U1254 (N_1254,N_708,N_709);
nor U1255 (N_1255,N_684,N_726);
nor U1256 (N_1256,N_522,N_936);
or U1257 (N_1257,N_763,N_559);
nor U1258 (N_1258,N_693,N_555);
or U1259 (N_1259,N_629,N_601);
or U1260 (N_1260,N_879,N_892);
nor U1261 (N_1261,N_822,N_640);
or U1262 (N_1262,N_974,N_909);
or U1263 (N_1263,N_532,N_945);
xnor U1264 (N_1264,N_595,N_957);
or U1265 (N_1265,N_750,N_869);
nor U1266 (N_1266,N_665,N_758);
and U1267 (N_1267,N_660,N_996);
nand U1268 (N_1268,N_635,N_824);
nor U1269 (N_1269,N_745,N_762);
or U1270 (N_1270,N_502,N_991);
nor U1271 (N_1271,N_788,N_710);
nand U1272 (N_1272,N_547,N_981);
nor U1273 (N_1273,N_591,N_686);
or U1274 (N_1274,N_923,N_644);
nor U1275 (N_1275,N_671,N_629);
and U1276 (N_1276,N_739,N_959);
nand U1277 (N_1277,N_833,N_880);
nor U1278 (N_1278,N_986,N_634);
or U1279 (N_1279,N_853,N_735);
nand U1280 (N_1280,N_643,N_540);
nor U1281 (N_1281,N_705,N_831);
nor U1282 (N_1282,N_518,N_631);
or U1283 (N_1283,N_730,N_627);
nand U1284 (N_1284,N_780,N_644);
nor U1285 (N_1285,N_723,N_759);
or U1286 (N_1286,N_899,N_696);
xnor U1287 (N_1287,N_804,N_672);
nor U1288 (N_1288,N_941,N_999);
or U1289 (N_1289,N_573,N_870);
and U1290 (N_1290,N_674,N_620);
and U1291 (N_1291,N_994,N_760);
and U1292 (N_1292,N_912,N_755);
nand U1293 (N_1293,N_921,N_561);
and U1294 (N_1294,N_871,N_863);
or U1295 (N_1295,N_749,N_726);
nand U1296 (N_1296,N_808,N_842);
nand U1297 (N_1297,N_514,N_920);
nand U1298 (N_1298,N_928,N_599);
nand U1299 (N_1299,N_747,N_828);
nand U1300 (N_1300,N_959,N_899);
nand U1301 (N_1301,N_733,N_612);
nor U1302 (N_1302,N_500,N_513);
or U1303 (N_1303,N_847,N_552);
or U1304 (N_1304,N_771,N_581);
nor U1305 (N_1305,N_925,N_519);
and U1306 (N_1306,N_949,N_818);
nor U1307 (N_1307,N_908,N_994);
and U1308 (N_1308,N_777,N_572);
nand U1309 (N_1309,N_523,N_559);
and U1310 (N_1310,N_557,N_591);
xor U1311 (N_1311,N_979,N_861);
or U1312 (N_1312,N_961,N_889);
nor U1313 (N_1313,N_762,N_728);
and U1314 (N_1314,N_797,N_702);
xnor U1315 (N_1315,N_805,N_660);
and U1316 (N_1316,N_922,N_644);
and U1317 (N_1317,N_796,N_780);
or U1318 (N_1318,N_852,N_773);
nor U1319 (N_1319,N_919,N_632);
nor U1320 (N_1320,N_771,N_739);
nor U1321 (N_1321,N_882,N_593);
and U1322 (N_1322,N_802,N_694);
nand U1323 (N_1323,N_781,N_620);
nand U1324 (N_1324,N_643,N_587);
nor U1325 (N_1325,N_503,N_728);
and U1326 (N_1326,N_747,N_736);
nor U1327 (N_1327,N_644,N_814);
or U1328 (N_1328,N_686,N_612);
xor U1329 (N_1329,N_768,N_613);
and U1330 (N_1330,N_788,N_554);
xnor U1331 (N_1331,N_744,N_696);
and U1332 (N_1332,N_504,N_932);
or U1333 (N_1333,N_979,N_577);
or U1334 (N_1334,N_536,N_874);
nor U1335 (N_1335,N_756,N_730);
and U1336 (N_1336,N_638,N_934);
nand U1337 (N_1337,N_856,N_660);
nand U1338 (N_1338,N_562,N_793);
nor U1339 (N_1339,N_663,N_742);
and U1340 (N_1340,N_764,N_686);
and U1341 (N_1341,N_698,N_984);
nand U1342 (N_1342,N_531,N_562);
and U1343 (N_1343,N_951,N_851);
and U1344 (N_1344,N_912,N_829);
and U1345 (N_1345,N_743,N_883);
nor U1346 (N_1346,N_829,N_669);
nand U1347 (N_1347,N_520,N_959);
nor U1348 (N_1348,N_760,N_671);
nand U1349 (N_1349,N_550,N_950);
and U1350 (N_1350,N_823,N_980);
and U1351 (N_1351,N_716,N_913);
and U1352 (N_1352,N_612,N_809);
or U1353 (N_1353,N_617,N_608);
nor U1354 (N_1354,N_546,N_611);
and U1355 (N_1355,N_684,N_600);
nor U1356 (N_1356,N_582,N_988);
or U1357 (N_1357,N_562,N_757);
nand U1358 (N_1358,N_988,N_952);
nand U1359 (N_1359,N_539,N_834);
nor U1360 (N_1360,N_664,N_960);
nand U1361 (N_1361,N_656,N_523);
and U1362 (N_1362,N_545,N_846);
or U1363 (N_1363,N_655,N_794);
and U1364 (N_1364,N_973,N_824);
xnor U1365 (N_1365,N_805,N_579);
and U1366 (N_1366,N_770,N_537);
nand U1367 (N_1367,N_593,N_770);
or U1368 (N_1368,N_546,N_903);
and U1369 (N_1369,N_944,N_837);
and U1370 (N_1370,N_529,N_952);
and U1371 (N_1371,N_975,N_901);
or U1372 (N_1372,N_874,N_678);
or U1373 (N_1373,N_627,N_927);
nand U1374 (N_1374,N_850,N_935);
xor U1375 (N_1375,N_704,N_814);
xnor U1376 (N_1376,N_628,N_519);
or U1377 (N_1377,N_864,N_623);
xnor U1378 (N_1378,N_807,N_520);
nand U1379 (N_1379,N_923,N_885);
or U1380 (N_1380,N_853,N_640);
and U1381 (N_1381,N_734,N_894);
nor U1382 (N_1382,N_855,N_808);
nor U1383 (N_1383,N_874,N_846);
xnor U1384 (N_1384,N_953,N_520);
nand U1385 (N_1385,N_927,N_909);
or U1386 (N_1386,N_817,N_573);
nor U1387 (N_1387,N_548,N_634);
xor U1388 (N_1388,N_753,N_684);
nand U1389 (N_1389,N_804,N_719);
nor U1390 (N_1390,N_680,N_831);
and U1391 (N_1391,N_982,N_626);
and U1392 (N_1392,N_751,N_991);
or U1393 (N_1393,N_777,N_716);
nand U1394 (N_1394,N_919,N_967);
nand U1395 (N_1395,N_653,N_759);
nand U1396 (N_1396,N_573,N_828);
nand U1397 (N_1397,N_881,N_816);
and U1398 (N_1398,N_662,N_805);
and U1399 (N_1399,N_603,N_761);
or U1400 (N_1400,N_819,N_906);
or U1401 (N_1401,N_906,N_715);
and U1402 (N_1402,N_851,N_764);
nor U1403 (N_1403,N_618,N_792);
or U1404 (N_1404,N_698,N_538);
nor U1405 (N_1405,N_631,N_761);
nand U1406 (N_1406,N_624,N_577);
or U1407 (N_1407,N_658,N_905);
or U1408 (N_1408,N_985,N_800);
and U1409 (N_1409,N_653,N_790);
nand U1410 (N_1410,N_622,N_922);
or U1411 (N_1411,N_781,N_931);
xor U1412 (N_1412,N_725,N_547);
nand U1413 (N_1413,N_997,N_797);
nand U1414 (N_1414,N_990,N_897);
nor U1415 (N_1415,N_737,N_682);
or U1416 (N_1416,N_696,N_560);
or U1417 (N_1417,N_721,N_898);
nand U1418 (N_1418,N_532,N_717);
and U1419 (N_1419,N_618,N_868);
and U1420 (N_1420,N_531,N_901);
nand U1421 (N_1421,N_573,N_708);
and U1422 (N_1422,N_795,N_653);
xnor U1423 (N_1423,N_870,N_634);
nand U1424 (N_1424,N_736,N_808);
nand U1425 (N_1425,N_657,N_524);
or U1426 (N_1426,N_636,N_803);
or U1427 (N_1427,N_504,N_723);
xor U1428 (N_1428,N_987,N_561);
or U1429 (N_1429,N_604,N_548);
nand U1430 (N_1430,N_818,N_595);
nor U1431 (N_1431,N_597,N_863);
and U1432 (N_1432,N_872,N_890);
and U1433 (N_1433,N_946,N_919);
or U1434 (N_1434,N_532,N_760);
and U1435 (N_1435,N_762,N_637);
nand U1436 (N_1436,N_690,N_871);
nor U1437 (N_1437,N_784,N_656);
and U1438 (N_1438,N_747,N_712);
or U1439 (N_1439,N_961,N_860);
nor U1440 (N_1440,N_755,N_831);
nor U1441 (N_1441,N_758,N_603);
nand U1442 (N_1442,N_809,N_568);
and U1443 (N_1443,N_862,N_824);
and U1444 (N_1444,N_954,N_765);
nand U1445 (N_1445,N_954,N_933);
nand U1446 (N_1446,N_617,N_811);
or U1447 (N_1447,N_657,N_928);
nand U1448 (N_1448,N_821,N_936);
or U1449 (N_1449,N_660,N_614);
nand U1450 (N_1450,N_684,N_512);
xnor U1451 (N_1451,N_838,N_584);
or U1452 (N_1452,N_634,N_938);
or U1453 (N_1453,N_526,N_664);
nor U1454 (N_1454,N_506,N_612);
or U1455 (N_1455,N_626,N_520);
xnor U1456 (N_1456,N_862,N_596);
or U1457 (N_1457,N_753,N_824);
nand U1458 (N_1458,N_936,N_919);
or U1459 (N_1459,N_529,N_744);
xnor U1460 (N_1460,N_871,N_524);
nor U1461 (N_1461,N_904,N_856);
nor U1462 (N_1462,N_884,N_510);
xnor U1463 (N_1463,N_507,N_688);
and U1464 (N_1464,N_695,N_796);
or U1465 (N_1465,N_676,N_817);
and U1466 (N_1466,N_546,N_710);
nand U1467 (N_1467,N_623,N_724);
nor U1468 (N_1468,N_925,N_702);
and U1469 (N_1469,N_919,N_952);
xor U1470 (N_1470,N_587,N_634);
nand U1471 (N_1471,N_764,N_955);
xor U1472 (N_1472,N_898,N_532);
nor U1473 (N_1473,N_893,N_526);
and U1474 (N_1474,N_781,N_782);
nand U1475 (N_1475,N_513,N_762);
nand U1476 (N_1476,N_918,N_734);
and U1477 (N_1477,N_902,N_665);
and U1478 (N_1478,N_736,N_706);
nand U1479 (N_1479,N_760,N_985);
and U1480 (N_1480,N_952,N_711);
nand U1481 (N_1481,N_943,N_543);
nand U1482 (N_1482,N_854,N_658);
and U1483 (N_1483,N_589,N_528);
nor U1484 (N_1484,N_787,N_533);
xor U1485 (N_1485,N_769,N_828);
or U1486 (N_1486,N_903,N_662);
and U1487 (N_1487,N_504,N_824);
or U1488 (N_1488,N_849,N_978);
or U1489 (N_1489,N_778,N_790);
xor U1490 (N_1490,N_786,N_903);
xnor U1491 (N_1491,N_842,N_747);
nor U1492 (N_1492,N_879,N_902);
or U1493 (N_1493,N_765,N_646);
nor U1494 (N_1494,N_819,N_738);
and U1495 (N_1495,N_792,N_887);
xor U1496 (N_1496,N_964,N_714);
nand U1497 (N_1497,N_619,N_523);
or U1498 (N_1498,N_964,N_579);
nand U1499 (N_1499,N_877,N_703);
and U1500 (N_1500,N_1081,N_1225);
and U1501 (N_1501,N_1441,N_1235);
or U1502 (N_1502,N_1119,N_1268);
xor U1503 (N_1503,N_1052,N_1229);
nor U1504 (N_1504,N_1038,N_1070);
or U1505 (N_1505,N_1005,N_1158);
xor U1506 (N_1506,N_1347,N_1267);
xnor U1507 (N_1507,N_1170,N_1438);
or U1508 (N_1508,N_1204,N_1228);
nand U1509 (N_1509,N_1405,N_1142);
nand U1510 (N_1510,N_1205,N_1289);
or U1511 (N_1511,N_1084,N_1395);
and U1512 (N_1512,N_1303,N_1226);
or U1513 (N_1513,N_1244,N_1296);
xor U1514 (N_1514,N_1026,N_1360);
nor U1515 (N_1515,N_1050,N_1497);
xnor U1516 (N_1516,N_1416,N_1449);
xnor U1517 (N_1517,N_1234,N_1265);
and U1518 (N_1518,N_1271,N_1138);
nor U1519 (N_1519,N_1317,N_1136);
and U1520 (N_1520,N_1112,N_1091);
nand U1521 (N_1521,N_1067,N_1080);
nor U1522 (N_1522,N_1049,N_1340);
nand U1523 (N_1523,N_1428,N_1288);
and U1524 (N_1524,N_1351,N_1315);
nand U1525 (N_1525,N_1383,N_1321);
nand U1526 (N_1526,N_1373,N_1043);
nand U1527 (N_1527,N_1398,N_1261);
nor U1528 (N_1528,N_1217,N_1314);
nand U1529 (N_1529,N_1237,N_1069);
and U1530 (N_1530,N_1446,N_1251);
nand U1531 (N_1531,N_1272,N_1174);
xnor U1532 (N_1532,N_1248,N_1019);
and U1533 (N_1533,N_1392,N_1483);
nand U1534 (N_1534,N_1278,N_1144);
nand U1535 (N_1535,N_1320,N_1364);
nand U1536 (N_1536,N_1419,N_1117);
and U1537 (N_1537,N_1254,N_1245);
nand U1538 (N_1538,N_1150,N_1089);
and U1539 (N_1539,N_1216,N_1285);
nand U1540 (N_1540,N_1143,N_1442);
and U1541 (N_1541,N_1368,N_1280);
or U1542 (N_1542,N_1433,N_1088);
nor U1543 (N_1543,N_1236,N_1424);
and U1544 (N_1544,N_1182,N_1023);
and U1545 (N_1545,N_1013,N_1313);
or U1546 (N_1546,N_1279,N_1128);
nand U1547 (N_1547,N_1400,N_1057);
nor U1548 (N_1548,N_1467,N_1202);
xnor U1549 (N_1549,N_1412,N_1406);
nand U1550 (N_1550,N_1463,N_1105);
and U1551 (N_1551,N_1075,N_1430);
or U1552 (N_1552,N_1127,N_1427);
and U1553 (N_1553,N_1155,N_1309);
nand U1554 (N_1554,N_1354,N_1218);
and U1555 (N_1555,N_1344,N_1482);
or U1556 (N_1556,N_1121,N_1055);
nor U1557 (N_1557,N_1472,N_1357);
or U1558 (N_1558,N_1066,N_1030);
nand U1559 (N_1559,N_1471,N_1387);
or U1560 (N_1560,N_1450,N_1118);
nand U1561 (N_1561,N_1042,N_1290);
nand U1562 (N_1562,N_1311,N_1012);
or U1563 (N_1563,N_1431,N_1444);
nor U1564 (N_1564,N_1407,N_1281);
or U1565 (N_1565,N_1453,N_1132);
and U1566 (N_1566,N_1458,N_1270);
nor U1567 (N_1567,N_1097,N_1141);
or U1568 (N_1568,N_1410,N_1096);
nor U1569 (N_1569,N_1255,N_1054);
and U1570 (N_1570,N_1061,N_1260);
nand U1571 (N_1571,N_1157,N_1399);
xor U1572 (N_1572,N_1106,N_1420);
or U1573 (N_1573,N_1196,N_1102);
xor U1574 (N_1574,N_1445,N_1099);
nor U1575 (N_1575,N_1083,N_1086);
or U1576 (N_1576,N_1448,N_1153);
xor U1577 (N_1577,N_1263,N_1133);
nor U1578 (N_1578,N_1404,N_1116);
nor U1579 (N_1579,N_1486,N_1488);
or U1580 (N_1580,N_1169,N_1499);
nor U1581 (N_1581,N_1479,N_1293);
nor U1582 (N_1582,N_1362,N_1429);
nor U1583 (N_1583,N_1455,N_1485);
nor U1584 (N_1584,N_1258,N_1187);
nand U1585 (N_1585,N_1198,N_1037);
nor U1586 (N_1586,N_1292,N_1257);
or U1587 (N_1587,N_1440,N_1101);
and U1588 (N_1588,N_1126,N_1186);
nand U1589 (N_1589,N_1266,N_1179);
and U1590 (N_1590,N_1165,N_1490);
nand U1591 (N_1591,N_1298,N_1018);
and U1592 (N_1592,N_1008,N_1327);
nand U1593 (N_1593,N_1339,N_1131);
nor U1594 (N_1594,N_1149,N_1011);
nor U1595 (N_1595,N_1495,N_1418);
or U1596 (N_1596,N_1283,N_1353);
or U1597 (N_1597,N_1171,N_1252);
nand U1598 (N_1598,N_1286,N_1434);
nor U1599 (N_1599,N_1491,N_1063);
nor U1600 (N_1600,N_1206,N_1231);
nor U1601 (N_1601,N_1468,N_1284);
or U1602 (N_1602,N_1194,N_1243);
and U1603 (N_1603,N_1496,N_1297);
and U1604 (N_1604,N_1466,N_1178);
or U1605 (N_1605,N_1017,N_1164);
or U1606 (N_1606,N_1181,N_1432);
nand U1607 (N_1607,N_1048,N_1422);
xnor U1608 (N_1608,N_1197,N_1145);
xor U1609 (N_1609,N_1060,N_1001);
nand U1610 (N_1610,N_1058,N_1010);
or U1611 (N_1611,N_1457,N_1123);
and U1612 (N_1612,N_1389,N_1473);
and U1613 (N_1613,N_1276,N_1113);
nand U1614 (N_1614,N_1319,N_1299);
and U1615 (N_1615,N_1213,N_1190);
nand U1616 (N_1616,N_1221,N_1476);
nor U1617 (N_1617,N_1016,N_1435);
and U1618 (N_1618,N_1401,N_1377);
and U1619 (N_1619,N_1059,N_1437);
or U1620 (N_1620,N_1129,N_1343);
or U1621 (N_1621,N_1064,N_1318);
nor U1622 (N_1622,N_1072,N_1305);
or U1623 (N_1623,N_1200,N_1277);
nand U1624 (N_1624,N_1421,N_1274);
nand U1625 (N_1625,N_1210,N_1323);
or U1626 (N_1626,N_1220,N_1162);
nand U1627 (N_1627,N_1139,N_1291);
xnor U1628 (N_1628,N_1163,N_1029);
and U1629 (N_1629,N_1349,N_1372);
nand U1630 (N_1630,N_1459,N_1413);
and U1631 (N_1631,N_1079,N_1098);
and U1632 (N_1632,N_1385,N_1125);
nor U1633 (N_1633,N_1045,N_1047);
and U1634 (N_1634,N_1262,N_1199);
or U1635 (N_1635,N_1253,N_1002);
nor U1636 (N_1636,N_1341,N_1247);
nand U1637 (N_1637,N_1146,N_1452);
nor U1638 (N_1638,N_1095,N_1172);
or U1639 (N_1639,N_1073,N_1183);
xnor U1640 (N_1640,N_1487,N_1122);
nor U1641 (N_1641,N_1300,N_1051);
or U1642 (N_1642,N_1147,N_1022);
and U1643 (N_1643,N_1068,N_1369);
nand U1644 (N_1644,N_1214,N_1361);
or U1645 (N_1645,N_1111,N_1185);
nand U1646 (N_1646,N_1065,N_1304);
nand U1647 (N_1647,N_1159,N_1464);
and U1648 (N_1648,N_1148,N_1242);
and U1649 (N_1649,N_1396,N_1379);
nor U1650 (N_1650,N_1191,N_1484);
and U1651 (N_1651,N_1233,N_1462);
and U1652 (N_1652,N_1036,N_1366);
nand U1653 (N_1653,N_1256,N_1295);
nand U1654 (N_1654,N_1020,N_1166);
or U1655 (N_1655,N_1024,N_1219);
and U1656 (N_1656,N_1409,N_1180);
or U1657 (N_1657,N_1140,N_1135);
nand U1658 (N_1658,N_1308,N_1201);
or U1659 (N_1659,N_1077,N_1408);
or U1660 (N_1660,N_1367,N_1041);
nand U1661 (N_1661,N_1474,N_1439);
or U1662 (N_1662,N_1134,N_1325);
nand U1663 (N_1663,N_1227,N_1469);
or U1664 (N_1664,N_1436,N_1342);
or U1665 (N_1665,N_1397,N_1239);
nor U1666 (N_1666,N_1212,N_1447);
xnor U1667 (N_1667,N_1371,N_1222);
and U1668 (N_1668,N_1302,N_1329);
and U1669 (N_1669,N_1374,N_1346);
and U1670 (N_1670,N_1259,N_1100);
nand U1671 (N_1671,N_1451,N_1076);
and U1672 (N_1672,N_1335,N_1411);
nand U1673 (N_1673,N_1137,N_1332);
or U1674 (N_1674,N_1004,N_1287);
or U1675 (N_1675,N_1224,N_1350);
and U1676 (N_1676,N_1039,N_1376);
or U1677 (N_1677,N_1326,N_1306);
xor U1678 (N_1678,N_1173,N_1282);
nand U1679 (N_1679,N_1114,N_1027);
nor U1680 (N_1680,N_1082,N_1230);
nand U1681 (N_1681,N_1322,N_1324);
and U1682 (N_1682,N_1209,N_1380);
nor U1683 (N_1683,N_1167,N_1124);
or U1684 (N_1684,N_1078,N_1208);
xnor U1685 (N_1685,N_1470,N_1307);
and U1686 (N_1686,N_1269,N_1034);
nor U1687 (N_1687,N_1152,N_1093);
nor U1688 (N_1688,N_1168,N_1333);
or U1689 (N_1689,N_1378,N_1035);
xor U1690 (N_1690,N_1195,N_1414);
nor U1691 (N_1691,N_1193,N_1090);
and U1692 (N_1692,N_1381,N_1087);
and U1693 (N_1693,N_1189,N_1074);
or U1694 (N_1694,N_1071,N_1365);
and U1695 (N_1695,N_1211,N_1188);
xnor U1696 (N_1696,N_1423,N_1358);
or U1697 (N_1697,N_1443,N_1130);
xnor U1698 (N_1698,N_1330,N_1337);
nor U1699 (N_1699,N_1477,N_1000);
nor U1700 (N_1700,N_1316,N_1031);
or U1701 (N_1701,N_1103,N_1348);
nand U1702 (N_1702,N_1223,N_1033);
or U1703 (N_1703,N_1240,N_1352);
or U1704 (N_1704,N_1192,N_1046);
or U1705 (N_1705,N_1454,N_1456);
nor U1706 (N_1706,N_1402,N_1294);
xnor U1707 (N_1707,N_1085,N_1154);
nand U1708 (N_1708,N_1151,N_1184);
nand U1709 (N_1709,N_1215,N_1492);
nand U1710 (N_1710,N_1044,N_1336);
nand U1711 (N_1711,N_1177,N_1104);
or U1712 (N_1712,N_1207,N_1370);
nor U1713 (N_1713,N_1460,N_1246);
nor U1714 (N_1714,N_1040,N_1249);
nand U1715 (N_1715,N_1375,N_1015);
or U1716 (N_1716,N_1062,N_1475);
and U1717 (N_1717,N_1388,N_1417);
nor U1718 (N_1718,N_1107,N_1489);
or U1719 (N_1719,N_1310,N_1498);
nand U1720 (N_1720,N_1056,N_1390);
nor U1721 (N_1721,N_1156,N_1108);
xnor U1722 (N_1722,N_1250,N_1160);
nor U1723 (N_1723,N_1312,N_1110);
xnor U1724 (N_1724,N_1355,N_1403);
nor U1725 (N_1725,N_1394,N_1032);
or U1726 (N_1726,N_1120,N_1391);
nor U1727 (N_1727,N_1175,N_1264);
nand U1728 (N_1728,N_1053,N_1275);
nor U1729 (N_1729,N_1334,N_1363);
and U1730 (N_1730,N_1480,N_1345);
xor U1731 (N_1731,N_1494,N_1384);
and U1732 (N_1732,N_1426,N_1094);
xnor U1733 (N_1733,N_1241,N_1161);
xor U1734 (N_1734,N_1425,N_1478);
or U1735 (N_1735,N_1176,N_1232);
nand U1736 (N_1736,N_1481,N_1493);
and U1737 (N_1737,N_1007,N_1338);
or U1738 (N_1738,N_1415,N_1203);
and U1739 (N_1739,N_1003,N_1238);
nor U1740 (N_1740,N_1115,N_1359);
and U1741 (N_1741,N_1006,N_1393);
nor U1742 (N_1742,N_1331,N_1014);
nor U1743 (N_1743,N_1465,N_1021);
or U1744 (N_1744,N_1382,N_1386);
xor U1745 (N_1745,N_1301,N_1009);
or U1746 (N_1746,N_1328,N_1092);
nand U1747 (N_1747,N_1109,N_1028);
nor U1748 (N_1748,N_1025,N_1461);
and U1749 (N_1749,N_1273,N_1356);
or U1750 (N_1750,N_1235,N_1364);
and U1751 (N_1751,N_1399,N_1236);
nor U1752 (N_1752,N_1084,N_1146);
nor U1753 (N_1753,N_1012,N_1003);
and U1754 (N_1754,N_1350,N_1243);
and U1755 (N_1755,N_1186,N_1272);
xnor U1756 (N_1756,N_1269,N_1429);
nor U1757 (N_1757,N_1088,N_1375);
or U1758 (N_1758,N_1077,N_1211);
nor U1759 (N_1759,N_1046,N_1391);
nand U1760 (N_1760,N_1330,N_1010);
or U1761 (N_1761,N_1000,N_1313);
or U1762 (N_1762,N_1058,N_1143);
and U1763 (N_1763,N_1284,N_1067);
and U1764 (N_1764,N_1259,N_1350);
and U1765 (N_1765,N_1172,N_1021);
or U1766 (N_1766,N_1469,N_1025);
xnor U1767 (N_1767,N_1415,N_1191);
nand U1768 (N_1768,N_1291,N_1395);
nand U1769 (N_1769,N_1249,N_1160);
nand U1770 (N_1770,N_1020,N_1490);
or U1771 (N_1771,N_1187,N_1316);
nor U1772 (N_1772,N_1478,N_1491);
nand U1773 (N_1773,N_1093,N_1365);
nor U1774 (N_1774,N_1007,N_1498);
nand U1775 (N_1775,N_1146,N_1209);
or U1776 (N_1776,N_1174,N_1181);
xor U1777 (N_1777,N_1332,N_1129);
nand U1778 (N_1778,N_1116,N_1007);
nand U1779 (N_1779,N_1392,N_1399);
and U1780 (N_1780,N_1320,N_1052);
nor U1781 (N_1781,N_1076,N_1005);
nand U1782 (N_1782,N_1043,N_1036);
and U1783 (N_1783,N_1088,N_1066);
or U1784 (N_1784,N_1294,N_1191);
nor U1785 (N_1785,N_1150,N_1046);
and U1786 (N_1786,N_1070,N_1159);
and U1787 (N_1787,N_1158,N_1438);
and U1788 (N_1788,N_1012,N_1397);
and U1789 (N_1789,N_1382,N_1473);
xor U1790 (N_1790,N_1126,N_1071);
nor U1791 (N_1791,N_1370,N_1461);
and U1792 (N_1792,N_1435,N_1074);
nand U1793 (N_1793,N_1072,N_1213);
and U1794 (N_1794,N_1125,N_1208);
or U1795 (N_1795,N_1254,N_1000);
nor U1796 (N_1796,N_1139,N_1475);
and U1797 (N_1797,N_1224,N_1448);
and U1798 (N_1798,N_1368,N_1058);
and U1799 (N_1799,N_1254,N_1422);
nand U1800 (N_1800,N_1465,N_1229);
or U1801 (N_1801,N_1263,N_1189);
xor U1802 (N_1802,N_1280,N_1224);
xnor U1803 (N_1803,N_1119,N_1322);
or U1804 (N_1804,N_1290,N_1316);
and U1805 (N_1805,N_1345,N_1496);
nand U1806 (N_1806,N_1140,N_1235);
nor U1807 (N_1807,N_1146,N_1303);
nand U1808 (N_1808,N_1442,N_1280);
nand U1809 (N_1809,N_1389,N_1262);
and U1810 (N_1810,N_1325,N_1126);
nor U1811 (N_1811,N_1052,N_1221);
xor U1812 (N_1812,N_1461,N_1289);
and U1813 (N_1813,N_1483,N_1165);
nand U1814 (N_1814,N_1249,N_1412);
nor U1815 (N_1815,N_1245,N_1216);
and U1816 (N_1816,N_1008,N_1139);
nor U1817 (N_1817,N_1312,N_1320);
and U1818 (N_1818,N_1009,N_1384);
nor U1819 (N_1819,N_1243,N_1364);
or U1820 (N_1820,N_1428,N_1037);
nand U1821 (N_1821,N_1403,N_1155);
or U1822 (N_1822,N_1256,N_1492);
and U1823 (N_1823,N_1021,N_1234);
or U1824 (N_1824,N_1176,N_1413);
nand U1825 (N_1825,N_1004,N_1345);
or U1826 (N_1826,N_1041,N_1000);
nand U1827 (N_1827,N_1114,N_1205);
or U1828 (N_1828,N_1106,N_1424);
xnor U1829 (N_1829,N_1324,N_1218);
and U1830 (N_1830,N_1139,N_1227);
and U1831 (N_1831,N_1043,N_1240);
nand U1832 (N_1832,N_1224,N_1218);
and U1833 (N_1833,N_1356,N_1031);
nor U1834 (N_1834,N_1354,N_1103);
and U1835 (N_1835,N_1138,N_1220);
nand U1836 (N_1836,N_1251,N_1003);
or U1837 (N_1837,N_1366,N_1340);
nand U1838 (N_1838,N_1409,N_1276);
nor U1839 (N_1839,N_1406,N_1067);
or U1840 (N_1840,N_1496,N_1072);
xnor U1841 (N_1841,N_1105,N_1047);
nor U1842 (N_1842,N_1259,N_1486);
or U1843 (N_1843,N_1101,N_1382);
and U1844 (N_1844,N_1465,N_1158);
nand U1845 (N_1845,N_1452,N_1453);
nand U1846 (N_1846,N_1107,N_1449);
nand U1847 (N_1847,N_1008,N_1031);
nand U1848 (N_1848,N_1085,N_1267);
xor U1849 (N_1849,N_1486,N_1119);
nor U1850 (N_1850,N_1433,N_1335);
and U1851 (N_1851,N_1400,N_1053);
and U1852 (N_1852,N_1445,N_1079);
or U1853 (N_1853,N_1373,N_1410);
and U1854 (N_1854,N_1369,N_1001);
xnor U1855 (N_1855,N_1069,N_1410);
or U1856 (N_1856,N_1199,N_1043);
nand U1857 (N_1857,N_1435,N_1216);
nand U1858 (N_1858,N_1299,N_1488);
xor U1859 (N_1859,N_1159,N_1295);
or U1860 (N_1860,N_1380,N_1123);
nor U1861 (N_1861,N_1262,N_1333);
or U1862 (N_1862,N_1498,N_1302);
nand U1863 (N_1863,N_1412,N_1025);
nor U1864 (N_1864,N_1285,N_1012);
or U1865 (N_1865,N_1453,N_1428);
or U1866 (N_1866,N_1465,N_1061);
xor U1867 (N_1867,N_1080,N_1034);
or U1868 (N_1868,N_1119,N_1236);
or U1869 (N_1869,N_1467,N_1354);
and U1870 (N_1870,N_1342,N_1083);
and U1871 (N_1871,N_1007,N_1480);
xor U1872 (N_1872,N_1171,N_1189);
and U1873 (N_1873,N_1399,N_1050);
nor U1874 (N_1874,N_1444,N_1220);
nor U1875 (N_1875,N_1165,N_1401);
xnor U1876 (N_1876,N_1038,N_1189);
xor U1877 (N_1877,N_1030,N_1027);
or U1878 (N_1878,N_1215,N_1491);
and U1879 (N_1879,N_1496,N_1300);
nor U1880 (N_1880,N_1121,N_1200);
nor U1881 (N_1881,N_1423,N_1062);
nor U1882 (N_1882,N_1080,N_1050);
and U1883 (N_1883,N_1403,N_1340);
nand U1884 (N_1884,N_1178,N_1199);
nor U1885 (N_1885,N_1268,N_1338);
nor U1886 (N_1886,N_1078,N_1281);
or U1887 (N_1887,N_1061,N_1296);
and U1888 (N_1888,N_1078,N_1226);
nor U1889 (N_1889,N_1023,N_1209);
or U1890 (N_1890,N_1137,N_1377);
nor U1891 (N_1891,N_1482,N_1325);
nor U1892 (N_1892,N_1391,N_1276);
xor U1893 (N_1893,N_1299,N_1010);
or U1894 (N_1894,N_1475,N_1270);
nand U1895 (N_1895,N_1202,N_1167);
or U1896 (N_1896,N_1386,N_1268);
nor U1897 (N_1897,N_1202,N_1452);
xnor U1898 (N_1898,N_1275,N_1391);
and U1899 (N_1899,N_1408,N_1325);
nor U1900 (N_1900,N_1070,N_1482);
and U1901 (N_1901,N_1208,N_1029);
xnor U1902 (N_1902,N_1358,N_1262);
or U1903 (N_1903,N_1360,N_1217);
nand U1904 (N_1904,N_1361,N_1177);
nor U1905 (N_1905,N_1172,N_1379);
nor U1906 (N_1906,N_1440,N_1186);
nand U1907 (N_1907,N_1459,N_1308);
xor U1908 (N_1908,N_1103,N_1232);
and U1909 (N_1909,N_1491,N_1125);
and U1910 (N_1910,N_1133,N_1187);
or U1911 (N_1911,N_1467,N_1209);
nor U1912 (N_1912,N_1080,N_1114);
nor U1913 (N_1913,N_1236,N_1353);
or U1914 (N_1914,N_1401,N_1309);
nand U1915 (N_1915,N_1095,N_1188);
nor U1916 (N_1916,N_1017,N_1122);
xnor U1917 (N_1917,N_1017,N_1055);
or U1918 (N_1918,N_1485,N_1330);
nand U1919 (N_1919,N_1427,N_1032);
nand U1920 (N_1920,N_1262,N_1263);
or U1921 (N_1921,N_1006,N_1132);
or U1922 (N_1922,N_1000,N_1413);
nand U1923 (N_1923,N_1434,N_1492);
and U1924 (N_1924,N_1253,N_1282);
or U1925 (N_1925,N_1071,N_1015);
nor U1926 (N_1926,N_1111,N_1212);
or U1927 (N_1927,N_1441,N_1335);
nor U1928 (N_1928,N_1431,N_1270);
nor U1929 (N_1929,N_1192,N_1119);
or U1930 (N_1930,N_1485,N_1499);
nor U1931 (N_1931,N_1004,N_1402);
nor U1932 (N_1932,N_1382,N_1027);
nor U1933 (N_1933,N_1218,N_1016);
nor U1934 (N_1934,N_1310,N_1007);
xnor U1935 (N_1935,N_1051,N_1377);
and U1936 (N_1936,N_1097,N_1297);
nor U1937 (N_1937,N_1442,N_1026);
and U1938 (N_1938,N_1123,N_1215);
xor U1939 (N_1939,N_1209,N_1084);
and U1940 (N_1940,N_1212,N_1096);
nor U1941 (N_1941,N_1179,N_1453);
nor U1942 (N_1942,N_1077,N_1104);
or U1943 (N_1943,N_1137,N_1433);
nand U1944 (N_1944,N_1056,N_1030);
or U1945 (N_1945,N_1441,N_1385);
nor U1946 (N_1946,N_1179,N_1041);
nand U1947 (N_1947,N_1026,N_1410);
xnor U1948 (N_1948,N_1485,N_1109);
or U1949 (N_1949,N_1319,N_1483);
nand U1950 (N_1950,N_1174,N_1290);
and U1951 (N_1951,N_1273,N_1474);
nand U1952 (N_1952,N_1242,N_1351);
and U1953 (N_1953,N_1244,N_1038);
nor U1954 (N_1954,N_1060,N_1175);
or U1955 (N_1955,N_1088,N_1242);
and U1956 (N_1956,N_1309,N_1209);
xnor U1957 (N_1957,N_1169,N_1370);
and U1958 (N_1958,N_1232,N_1343);
and U1959 (N_1959,N_1356,N_1292);
and U1960 (N_1960,N_1492,N_1080);
or U1961 (N_1961,N_1198,N_1400);
nand U1962 (N_1962,N_1131,N_1176);
nand U1963 (N_1963,N_1348,N_1281);
xnor U1964 (N_1964,N_1119,N_1421);
and U1965 (N_1965,N_1044,N_1135);
nand U1966 (N_1966,N_1118,N_1084);
nor U1967 (N_1967,N_1153,N_1156);
nor U1968 (N_1968,N_1244,N_1062);
or U1969 (N_1969,N_1003,N_1415);
nand U1970 (N_1970,N_1172,N_1404);
or U1971 (N_1971,N_1334,N_1212);
nor U1972 (N_1972,N_1349,N_1299);
nand U1973 (N_1973,N_1232,N_1449);
nor U1974 (N_1974,N_1498,N_1316);
and U1975 (N_1975,N_1096,N_1136);
and U1976 (N_1976,N_1436,N_1404);
and U1977 (N_1977,N_1127,N_1357);
nor U1978 (N_1978,N_1219,N_1402);
nand U1979 (N_1979,N_1036,N_1333);
xor U1980 (N_1980,N_1241,N_1065);
or U1981 (N_1981,N_1116,N_1121);
nand U1982 (N_1982,N_1446,N_1387);
nand U1983 (N_1983,N_1041,N_1185);
or U1984 (N_1984,N_1483,N_1432);
nor U1985 (N_1985,N_1444,N_1032);
nor U1986 (N_1986,N_1286,N_1124);
nor U1987 (N_1987,N_1048,N_1338);
nor U1988 (N_1988,N_1418,N_1322);
nand U1989 (N_1989,N_1468,N_1110);
and U1990 (N_1990,N_1399,N_1409);
nand U1991 (N_1991,N_1058,N_1480);
or U1992 (N_1992,N_1393,N_1363);
or U1993 (N_1993,N_1496,N_1295);
or U1994 (N_1994,N_1328,N_1151);
nand U1995 (N_1995,N_1115,N_1192);
nand U1996 (N_1996,N_1031,N_1113);
or U1997 (N_1997,N_1288,N_1265);
or U1998 (N_1998,N_1493,N_1142);
and U1999 (N_1999,N_1258,N_1302);
or U2000 (N_2000,N_1583,N_1554);
or U2001 (N_2001,N_1979,N_1515);
nor U2002 (N_2002,N_1881,N_1910);
or U2003 (N_2003,N_1586,N_1607);
and U2004 (N_2004,N_1955,N_1510);
xor U2005 (N_2005,N_1538,N_1502);
nand U2006 (N_2006,N_1895,N_1900);
nand U2007 (N_2007,N_1858,N_1570);
and U2008 (N_2008,N_1822,N_1621);
nand U2009 (N_2009,N_1928,N_1521);
nor U2010 (N_2010,N_1985,N_1546);
nand U2011 (N_2011,N_1509,N_1736);
or U2012 (N_2012,N_1735,N_1567);
and U2013 (N_2013,N_1639,N_1615);
nand U2014 (N_2014,N_1804,N_1951);
nor U2015 (N_2015,N_1786,N_1633);
nor U2016 (N_2016,N_1749,N_1721);
or U2017 (N_2017,N_1645,N_1933);
nor U2018 (N_2018,N_1726,N_1924);
nor U2019 (N_2019,N_1823,N_1661);
and U2020 (N_2020,N_1730,N_1802);
xnor U2021 (N_2021,N_1988,N_1803);
nand U2022 (N_2022,N_1576,N_1571);
nor U2023 (N_2023,N_1609,N_1624);
nor U2024 (N_2024,N_1818,N_1580);
nand U2025 (N_2025,N_1534,N_1631);
xnor U2026 (N_2026,N_1968,N_1632);
or U2027 (N_2027,N_1666,N_1612);
and U2028 (N_2028,N_1608,N_1662);
or U2029 (N_2029,N_1716,N_1693);
or U2030 (N_2030,N_1634,N_1992);
and U2031 (N_2031,N_1519,N_1854);
and U2032 (N_2032,N_1866,N_1750);
and U2033 (N_2033,N_1815,N_1941);
or U2034 (N_2034,N_1880,N_1691);
nor U2035 (N_2035,N_1766,N_1655);
nor U2036 (N_2036,N_1562,N_1522);
nand U2037 (N_2037,N_1500,N_1986);
and U2038 (N_2038,N_1757,N_1848);
xnor U2039 (N_2039,N_1764,N_1877);
and U2040 (N_2040,N_1630,N_1511);
or U2041 (N_2041,N_1518,N_1808);
nand U2042 (N_2042,N_1626,N_1718);
nor U2043 (N_2043,N_1821,N_1715);
and U2044 (N_2044,N_1589,N_1679);
xor U2045 (N_2045,N_1878,N_1660);
nand U2046 (N_2046,N_1953,N_1669);
and U2047 (N_2047,N_1779,N_1654);
nand U2048 (N_2048,N_1755,N_1969);
nand U2049 (N_2049,N_1742,N_1667);
nand U2050 (N_2050,N_1962,N_1973);
nand U2051 (N_2051,N_1672,N_1991);
nor U2052 (N_2052,N_1835,N_1945);
nor U2053 (N_2053,N_1839,N_1532);
nor U2054 (N_2054,N_1801,N_1996);
nand U2055 (N_2055,N_1588,N_1575);
nor U2056 (N_2056,N_1677,N_1700);
and U2057 (N_2057,N_1787,N_1710);
or U2058 (N_2058,N_1772,N_1850);
nor U2059 (N_2059,N_1717,N_1694);
xor U2060 (N_2060,N_1705,N_1875);
nand U2061 (N_2061,N_1657,N_1563);
xor U2062 (N_2062,N_1731,N_1874);
and U2063 (N_2063,N_1957,N_1796);
or U2064 (N_2064,N_1926,N_1758);
nand U2065 (N_2065,N_1959,N_1884);
and U2066 (N_2066,N_1919,N_1865);
nor U2067 (N_2067,N_1635,N_1975);
or U2068 (N_2068,N_1762,N_1552);
nor U2069 (N_2069,N_1771,N_1596);
nor U2070 (N_2070,N_1743,N_1964);
xnor U2071 (N_2071,N_1756,N_1685);
and U2072 (N_2072,N_1847,N_1864);
nand U2073 (N_2073,N_1961,N_1703);
nand U2074 (N_2074,N_1564,N_1838);
and U2075 (N_2075,N_1820,N_1551);
nand U2076 (N_2076,N_1828,N_1870);
xor U2077 (N_2077,N_1826,N_1656);
and U2078 (N_2078,N_1722,N_1976);
nor U2079 (N_2079,N_1760,N_1605);
nor U2080 (N_2080,N_1747,N_1692);
or U2081 (N_2081,N_1610,N_1582);
or U2082 (N_2082,N_1876,N_1739);
and U2083 (N_2083,N_1573,N_1812);
nor U2084 (N_2084,N_1636,N_1934);
xor U2085 (N_2085,N_1545,N_1768);
and U2086 (N_2086,N_1713,N_1687);
or U2087 (N_2087,N_1763,N_1673);
or U2088 (N_2088,N_1723,N_1547);
nand U2089 (N_2089,N_1653,N_1983);
or U2090 (N_2090,N_1784,N_1907);
nor U2091 (N_2091,N_1912,N_1528);
nand U2092 (N_2092,N_1972,N_1819);
or U2093 (N_2093,N_1593,N_1618);
nand U2094 (N_2094,N_1863,N_1602);
or U2095 (N_2095,N_1861,N_1652);
or U2096 (N_2096,N_1872,N_1981);
and U2097 (N_2097,N_1627,N_1642);
nor U2098 (N_2098,N_1777,N_1670);
nor U2099 (N_2099,N_1845,N_1792);
or U2100 (N_2100,N_1684,N_1711);
nand U2101 (N_2101,N_1560,N_1892);
or U2102 (N_2102,N_1680,N_1949);
or U2103 (N_2103,N_1943,N_1782);
and U2104 (N_2104,N_1543,N_1753);
or U2105 (N_2105,N_1944,N_1851);
xor U2106 (N_2106,N_1927,N_1879);
nor U2107 (N_2107,N_1888,N_1550);
xor U2108 (N_2108,N_1971,N_1585);
or U2109 (N_2109,N_1688,N_1650);
xor U2110 (N_2110,N_1849,N_1520);
nor U2111 (N_2111,N_1725,N_1530);
nand U2112 (N_2112,N_1794,N_1728);
and U2113 (N_2113,N_1614,N_1590);
nor U2114 (N_2114,N_1891,N_1556);
and U2115 (N_2115,N_1512,N_1997);
or U2116 (N_2116,N_1906,N_1526);
nor U2117 (N_2117,N_1911,N_1974);
or U2118 (N_2118,N_1681,N_1938);
or U2119 (N_2119,N_1853,N_1899);
nor U2120 (N_2120,N_1523,N_1896);
or U2121 (N_2121,N_1600,N_1886);
nand U2122 (N_2122,N_1824,N_1995);
or U2123 (N_2123,N_1952,N_1869);
or U2124 (N_2124,N_1531,N_1574);
nor U2125 (N_2125,N_1651,N_1587);
nand U2126 (N_2126,N_1929,N_1540);
and U2127 (N_2127,N_1727,N_1914);
nor U2128 (N_2128,N_1533,N_1595);
and U2129 (N_2129,N_1620,N_1836);
and U2130 (N_2130,N_1769,N_1606);
and U2131 (N_2131,N_1675,N_1601);
nand U2132 (N_2132,N_1561,N_1708);
and U2133 (N_2133,N_1935,N_1733);
or U2134 (N_2134,N_1579,N_1581);
and U2135 (N_2135,N_1852,N_1553);
nor U2136 (N_2136,N_1682,N_1873);
and U2137 (N_2137,N_1844,N_1846);
or U2138 (N_2138,N_1748,N_1829);
or U2139 (N_2139,N_1781,N_1699);
nand U2140 (N_2140,N_1536,N_1701);
xnor U2141 (N_2141,N_1984,N_1734);
and U2142 (N_2142,N_1939,N_1702);
nor U2143 (N_2143,N_1738,N_1663);
or U2144 (N_2144,N_1999,N_1640);
and U2145 (N_2145,N_1559,N_1506);
xor U2146 (N_2146,N_1629,N_1931);
or U2147 (N_2147,N_1987,N_1737);
and U2148 (N_2148,N_1752,N_1658);
or U2149 (N_2149,N_1720,N_1555);
or U2150 (N_2150,N_1584,N_1857);
and U2151 (N_2151,N_1767,N_1568);
nand U2152 (N_2152,N_1572,N_1901);
nand U2153 (N_2153,N_1619,N_1665);
nand U2154 (N_2154,N_1746,N_1825);
or U2155 (N_2155,N_1980,N_1548);
or U2156 (N_2156,N_1709,N_1916);
nand U2157 (N_2157,N_1732,N_1505);
nor U2158 (N_2158,N_1978,N_1990);
nor U2159 (N_2159,N_1729,N_1946);
xnor U2160 (N_2160,N_1960,N_1867);
nand U2161 (N_2161,N_1807,N_1542);
or U2162 (N_2162,N_1887,N_1625);
and U2163 (N_2163,N_1811,N_1517);
nand U2164 (N_2164,N_1800,N_1789);
nor U2165 (N_2165,N_1628,N_1671);
xor U2166 (N_2166,N_1503,N_1741);
and U2167 (N_2167,N_1967,N_1837);
and U2168 (N_2168,N_1578,N_1833);
and U2169 (N_2169,N_1780,N_1791);
nand U2170 (N_2170,N_1604,N_1740);
xnor U2171 (N_2171,N_1659,N_1898);
or U2172 (N_2172,N_1908,N_1966);
nor U2173 (N_2173,N_1504,N_1797);
xnor U2174 (N_2174,N_1759,N_1539);
or U2175 (N_2175,N_1501,N_1641);
nor U2176 (N_2176,N_1603,N_1599);
or U2177 (N_2177,N_1695,N_1566);
and U2178 (N_2178,N_1617,N_1788);
and U2179 (N_2179,N_1790,N_1765);
nor U2180 (N_2180,N_1597,N_1936);
nand U2181 (N_2181,N_1909,N_1882);
nor U2182 (N_2182,N_1649,N_1842);
or U2183 (N_2183,N_1817,N_1834);
nand U2184 (N_2184,N_1982,N_1754);
or U2185 (N_2185,N_1527,N_1883);
and U2186 (N_2186,N_1577,N_1696);
and U2187 (N_2187,N_1954,N_1776);
or U2188 (N_2188,N_1594,N_1745);
and U2189 (N_2189,N_1668,N_1647);
or U2190 (N_2190,N_1557,N_1831);
or U2191 (N_2191,N_1989,N_1816);
nor U2192 (N_2192,N_1686,N_1591);
nand U2193 (N_2193,N_1813,N_1856);
nor U2194 (N_2194,N_1902,N_1915);
nor U2195 (N_2195,N_1947,N_1956);
or U2196 (N_2196,N_1507,N_1994);
nand U2197 (N_2197,N_1970,N_1643);
nand U2198 (N_2198,N_1644,N_1958);
or U2199 (N_2199,N_1932,N_1917);
or U2200 (N_2200,N_1761,N_1508);
or U2201 (N_2201,N_1683,N_1707);
nor U2202 (N_2202,N_1950,N_1798);
xnor U2203 (N_2203,N_1697,N_1751);
nand U2204 (N_2204,N_1814,N_1859);
and U2205 (N_2205,N_1637,N_1773);
nor U2206 (N_2206,N_1623,N_1930);
xor U2207 (N_2207,N_1993,N_1525);
and U2208 (N_2208,N_1775,N_1558);
nand U2209 (N_2209,N_1862,N_1674);
or U2210 (N_2210,N_1598,N_1616);
nor U2211 (N_2211,N_1793,N_1940);
or U2212 (N_2212,N_1913,N_1925);
xnor U2213 (N_2213,N_1805,N_1611);
or U2214 (N_2214,N_1690,N_1885);
xor U2215 (N_2215,N_1855,N_1860);
or U2216 (N_2216,N_1706,N_1638);
or U2217 (N_2217,N_1799,N_1689);
xnor U2218 (N_2218,N_1774,N_1537);
and U2219 (N_2219,N_1920,N_1942);
or U2220 (N_2220,N_1905,N_1806);
and U2221 (N_2221,N_1809,N_1785);
or U2222 (N_2222,N_1843,N_1921);
or U2223 (N_2223,N_1937,N_1963);
and U2224 (N_2224,N_1516,N_1524);
and U2225 (N_2225,N_1678,N_1513);
and U2226 (N_2226,N_1676,N_1889);
xor U2227 (N_2227,N_1698,N_1744);
nor U2228 (N_2228,N_1646,N_1549);
or U2229 (N_2229,N_1923,N_1569);
or U2230 (N_2230,N_1778,N_1918);
nand U2231 (N_2231,N_1894,N_1893);
and U2232 (N_2232,N_1903,N_1830);
nor U2233 (N_2233,N_1904,N_1622);
and U2234 (N_2234,N_1565,N_1704);
xnor U2235 (N_2235,N_1890,N_1795);
and U2236 (N_2236,N_1827,N_1770);
or U2237 (N_2237,N_1832,N_1719);
and U2238 (N_2238,N_1998,N_1810);
xnor U2239 (N_2239,N_1613,N_1514);
nor U2240 (N_2240,N_1529,N_1922);
nand U2241 (N_2241,N_1724,N_1535);
nor U2242 (N_2242,N_1840,N_1712);
nand U2243 (N_2243,N_1544,N_1948);
and U2244 (N_2244,N_1648,N_1871);
and U2245 (N_2245,N_1868,N_1714);
xnor U2246 (N_2246,N_1783,N_1977);
and U2247 (N_2247,N_1965,N_1841);
xnor U2248 (N_2248,N_1541,N_1897);
xor U2249 (N_2249,N_1592,N_1664);
xor U2250 (N_2250,N_1695,N_1896);
nor U2251 (N_2251,N_1771,N_1662);
or U2252 (N_2252,N_1834,N_1623);
xor U2253 (N_2253,N_1878,N_1812);
nand U2254 (N_2254,N_1827,N_1852);
or U2255 (N_2255,N_1518,N_1573);
or U2256 (N_2256,N_1904,N_1619);
nor U2257 (N_2257,N_1974,N_1871);
xor U2258 (N_2258,N_1589,N_1631);
and U2259 (N_2259,N_1524,N_1679);
and U2260 (N_2260,N_1826,N_1794);
nor U2261 (N_2261,N_1549,N_1502);
and U2262 (N_2262,N_1570,N_1629);
xor U2263 (N_2263,N_1803,N_1833);
nor U2264 (N_2264,N_1921,N_1735);
and U2265 (N_2265,N_1683,N_1845);
nor U2266 (N_2266,N_1599,N_1554);
nand U2267 (N_2267,N_1506,N_1665);
or U2268 (N_2268,N_1656,N_1762);
nor U2269 (N_2269,N_1731,N_1586);
or U2270 (N_2270,N_1974,N_1888);
or U2271 (N_2271,N_1701,N_1848);
or U2272 (N_2272,N_1735,N_1552);
xor U2273 (N_2273,N_1964,N_1752);
and U2274 (N_2274,N_1781,N_1833);
nand U2275 (N_2275,N_1596,N_1518);
and U2276 (N_2276,N_1552,N_1722);
or U2277 (N_2277,N_1599,N_1715);
or U2278 (N_2278,N_1683,N_1798);
nand U2279 (N_2279,N_1512,N_1621);
nor U2280 (N_2280,N_1937,N_1755);
or U2281 (N_2281,N_1679,N_1644);
or U2282 (N_2282,N_1503,N_1645);
and U2283 (N_2283,N_1932,N_1605);
and U2284 (N_2284,N_1514,N_1969);
and U2285 (N_2285,N_1674,N_1795);
and U2286 (N_2286,N_1892,N_1816);
and U2287 (N_2287,N_1935,N_1727);
and U2288 (N_2288,N_1757,N_1505);
nor U2289 (N_2289,N_1942,N_1753);
nor U2290 (N_2290,N_1708,N_1749);
nand U2291 (N_2291,N_1518,N_1629);
and U2292 (N_2292,N_1638,N_1972);
nand U2293 (N_2293,N_1843,N_1608);
nor U2294 (N_2294,N_1781,N_1913);
nand U2295 (N_2295,N_1812,N_1888);
xnor U2296 (N_2296,N_1512,N_1704);
or U2297 (N_2297,N_1946,N_1959);
nor U2298 (N_2298,N_1723,N_1511);
or U2299 (N_2299,N_1660,N_1730);
nor U2300 (N_2300,N_1963,N_1654);
nor U2301 (N_2301,N_1742,N_1642);
nand U2302 (N_2302,N_1906,N_1846);
or U2303 (N_2303,N_1886,N_1960);
nor U2304 (N_2304,N_1775,N_1760);
or U2305 (N_2305,N_1534,N_1506);
xor U2306 (N_2306,N_1657,N_1746);
nor U2307 (N_2307,N_1889,N_1613);
xor U2308 (N_2308,N_1526,N_1563);
nand U2309 (N_2309,N_1833,N_1527);
xor U2310 (N_2310,N_1960,N_1724);
nor U2311 (N_2311,N_1729,N_1664);
nor U2312 (N_2312,N_1867,N_1851);
nand U2313 (N_2313,N_1823,N_1585);
or U2314 (N_2314,N_1909,N_1527);
or U2315 (N_2315,N_1898,N_1734);
nor U2316 (N_2316,N_1632,N_1737);
nand U2317 (N_2317,N_1775,N_1951);
nor U2318 (N_2318,N_1798,N_1779);
or U2319 (N_2319,N_1563,N_1938);
nor U2320 (N_2320,N_1944,N_1766);
nand U2321 (N_2321,N_1858,N_1808);
nor U2322 (N_2322,N_1946,N_1634);
xnor U2323 (N_2323,N_1508,N_1635);
or U2324 (N_2324,N_1540,N_1906);
nand U2325 (N_2325,N_1689,N_1744);
nor U2326 (N_2326,N_1595,N_1646);
and U2327 (N_2327,N_1906,N_1531);
and U2328 (N_2328,N_1548,N_1733);
or U2329 (N_2329,N_1520,N_1689);
nor U2330 (N_2330,N_1987,N_1699);
nor U2331 (N_2331,N_1525,N_1930);
and U2332 (N_2332,N_1933,N_1590);
nand U2333 (N_2333,N_1914,N_1600);
and U2334 (N_2334,N_1825,N_1687);
nor U2335 (N_2335,N_1726,N_1979);
nand U2336 (N_2336,N_1566,N_1749);
nor U2337 (N_2337,N_1784,N_1534);
nand U2338 (N_2338,N_1704,N_1756);
nand U2339 (N_2339,N_1948,N_1745);
and U2340 (N_2340,N_1589,N_1962);
or U2341 (N_2341,N_1883,N_1844);
or U2342 (N_2342,N_1782,N_1553);
or U2343 (N_2343,N_1743,N_1806);
or U2344 (N_2344,N_1745,N_1952);
and U2345 (N_2345,N_1914,N_1610);
nor U2346 (N_2346,N_1893,N_1900);
nor U2347 (N_2347,N_1839,N_1934);
nor U2348 (N_2348,N_1664,N_1807);
nand U2349 (N_2349,N_1754,N_1778);
nand U2350 (N_2350,N_1954,N_1773);
and U2351 (N_2351,N_1843,N_1658);
nor U2352 (N_2352,N_1511,N_1861);
or U2353 (N_2353,N_1869,N_1908);
and U2354 (N_2354,N_1912,N_1868);
or U2355 (N_2355,N_1890,N_1781);
or U2356 (N_2356,N_1559,N_1630);
nor U2357 (N_2357,N_1536,N_1610);
and U2358 (N_2358,N_1633,N_1936);
xnor U2359 (N_2359,N_1694,N_1807);
nand U2360 (N_2360,N_1658,N_1730);
nor U2361 (N_2361,N_1602,N_1727);
xnor U2362 (N_2362,N_1872,N_1615);
nand U2363 (N_2363,N_1803,N_1895);
or U2364 (N_2364,N_1809,N_1601);
or U2365 (N_2365,N_1508,N_1974);
nand U2366 (N_2366,N_1636,N_1982);
nor U2367 (N_2367,N_1853,N_1963);
xor U2368 (N_2368,N_1909,N_1964);
and U2369 (N_2369,N_1575,N_1893);
nand U2370 (N_2370,N_1942,N_1991);
and U2371 (N_2371,N_1783,N_1651);
or U2372 (N_2372,N_1797,N_1573);
or U2373 (N_2373,N_1774,N_1689);
nor U2374 (N_2374,N_1668,N_1515);
and U2375 (N_2375,N_1538,N_1620);
and U2376 (N_2376,N_1976,N_1539);
nor U2377 (N_2377,N_1684,N_1999);
and U2378 (N_2378,N_1899,N_1512);
nor U2379 (N_2379,N_1888,N_1703);
nor U2380 (N_2380,N_1836,N_1876);
nand U2381 (N_2381,N_1621,N_1523);
nand U2382 (N_2382,N_1811,N_1698);
nor U2383 (N_2383,N_1735,N_1612);
and U2384 (N_2384,N_1928,N_1583);
or U2385 (N_2385,N_1643,N_1532);
nor U2386 (N_2386,N_1905,N_1677);
and U2387 (N_2387,N_1898,N_1736);
nor U2388 (N_2388,N_1876,N_1793);
xor U2389 (N_2389,N_1642,N_1508);
nor U2390 (N_2390,N_1848,N_1759);
and U2391 (N_2391,N_1690,N_1586);
or U2392 (N_2392,N_1587,N_1560);
nand U2393 (N_2393,N_1906,N_1678);
xor U2394 (N_2394,N_1507,N_1744);
and U2395 (N_2395,N_1936,N_1631);
and U2396 (N_2396,N_1919,N_1756);
nor U2397 (N_2397,N_1692,N_1639);
or U2398 (N_2398,N_1641,N_1808);
nor U2399 (N_2399,N_1950,N_1743);
or U2400 (N_2400,N_1729,N_1804);
or U2401 (N_2401,N_1807,N_1867);
xor U2402 (N_2402,N_1851,N_1673);
nand U2403 (N_2403,N_1501,N_1698);
nand U2404 (N_2404,N_1537,N_1930);
or U2405 (N_2405,N_1983,N_1562);
or U2406 (N_2406,N_1734,N_1995);
or U2407 (N_2407,N_1903,N_1805);
nor U2408 (N_2408,N_1646,N_1584);
nor U2409 (N_2409,N_1565,N_1771);
nand U2410 (N_2410,N_1961,N_1734);
and U2411 (N_2411,N_1523,N_1700);
nor U2412 (N_2412,N_1992,N_1799);
nor U2413 (N_2413,N_1910,N_1679);
or U2414 (N_2414,N_1972,N_1563);
nand U2415 (N_2415,N_1541,N_1576);
xnor U2416 (N_2416,N_1937,N_1561);
and U2417 (N_2417,N_1915,N_1689);
nand U2418 (N_2418,N_1838,N_1912);
xnor U2419 (N_2419,N_1914,N_1738);
nor U2420 (N_2420,N_1577,N_1706);
or U2421 (N_2421,N_1820,N_1831);
nor U2422 (N_2422,N_1568,N_1723);
or U2423 (N_2423,N_1791,N_1631);
nor U2424 (N_2424,N_1511,N_1502);
nand U2425 (N_2425,N_1685,N_1637);
or U2426 (N_2426,N_1645,N_1852);
or U2427 (N_2427,N_1823,N_1828);
or U2428 (N_2428,N_1974,N_1717);
xor U2429 (N_2429,N_1564,N_1839);
and U2430 (N_2430,N_1769,N_1763);
and U2431 (N_2431,N_1702,N_1942);
nor U2432 (N_2432,N_1955,N_1977);
nand U2433 (N_2433,N_1663,N_1675);
nor U2434 (N_2434,N_1874,N_1578);
nor U2435 (N_2435,N_1842,N_1602);
and U2436 (N_2436,N_1980,N_1558);
or U2437 (N_2437,N_1962,N_1646);
nand U2438 (N_2438,N_1742,N_1849);
and U2439 (N_2439,N_1843,N_1743);
nand U2440 (N_2440,N_1894,N_1942);
nor U2441 (N_2441,N_1764,N_1993);
or U2442 (N_2442,N_1653,N_1796);
nand U2443 (N_2443,N_1686,N_1840);
nand U2444 (N_2444,N_1849,N_1559);
or U2445 (N_2445,N_1963,N_1706);
nand U2446 (N_2446,N_1791,N_1601);
or U2447 (N_2447,N_1765,N_1586);
nor U2448 (N_2448,N_1903,N_1889);
nor U2449 (N_2449,N_1680,N_1846);
nand U2450 (N_2450,N_1827,N_1800);
or U2451 (N_2451,N_1773,N_1561);
xnor U2452 (N_2452,N_1913,N_1651);
or U2453 (N_2453,N_1925,N_1617);
and U2454 (N_2454,N_1959,N_1758);
and U2455 (N_2455,N_1848,N_1753);
nand U2456 (N_2456,N_1753,N_1896);
and U2457 (N_2457,N_1965,N_1904);
or U2458 (N_2458,N_1656,N_1742);
xor U2459 (N_2459,N_1589,N_1956);
or U2460 (N_2460,N_1700,N_1886);
or U2461 (N_2461,N_1544,N_1864);
nand U2462 (N_2462,N_1807,N_1916);
nor U2463 (N_2463,N_1585,N_1883);
nor U2464 (N_2464,N_1587,N_1958);
nor U2465 (N_2465,N_1808,N_1735);
nand U2466 (N_2466,N_1854,N_1884);
or U2467 (N_2467,N_1680,N_1886);
and U2468 (N_2468,N_1735,N_1983);
nand U2469 (N_2469,N_1559,N_1936);
nor U2470 (N_2470,N_1860,N_1950);
xnor U2471 (N_2471,N_1571,N_1733);
and U2472 (N_2472,N_1921,N_1577);
xor U2473 (N_2473,N_1848,N_1532);
nor U2474 (N_2474,N_1856,N_1985);
or U2475 (N_2475,N_1658,N_1589);
or U2476 (N_2476,N_1897,N_1734);
nor U2477 (N_2477,N_1631,N_1573);
and U2478 (N_2478,N_1897,N_1710);
xor U2479 (N_2479,N_1544,N_1514);
nand U2480 (N_2480,N_1605,N_1603);
and U2481 (N_2481,N_1803,N_1996);
nand U2482 (N_2482,N_1503,N_1500);
or U2483 (N_2483,N_1715,N_1585);
nand U2484 (N_2484,N_1700,N_1947);
xor U2485 (N_2485,N_1539,N_1661);
nor U2486 (N_2486,N_1927,N_1946);
nor U2487 (N_2487,N_1832,N_1574);
or U2488 (N_2488,N_1633,N_1954);
nand U2489 (N_2489,N_1872,N_1717);
nand U2490 (N_2490,N_1955,N_1990);
or U2491 (N_2491,N_1751,N_1673);
nand U2492 (N_2492,N_1662,N_1680);
nand U2493 (N_2493,N_1649,N_1550);
nand U2494 (N_2494,N_1536,N_1724);
nor U2495 (N_2495,N_1861,N_1544);
or U2496 (N_2496,N_1721,N_1618);
or U2497 (N_2497,N_1527,N_1856);
xor U2498 (N_2498,N_1959,N_1546);
and U2499 (N_2499,N_1671,N_1615);
nor U2500 (N_2500,N_2014,N_2073);
or U2501 (N_2501,N_2460,N_2354);
and U2502 (N_2502,N_2126,N_2383);
or U2503 (N_2503,N_2470,N_2416);
nand U2504 (N_2504,N_2472,N_2045);
nor U2505 (N_2505,N_2150,N_2272);
nand U2506 (N_2506,N_2418,N_2101);
and U2507 (N_2507,N_2125,N_2321);
or U2508 (N_2508,N_2459,N_2095);
nand U2509 (N_2509,N_2113,N_2395);
xnor U2510 (N_2510,N_2443,N_2121);
nand U2511 (N_2511,N_2074,N_2001);
nand U2512 (N_2512,N_2000,N_2270);
nand U2513 (N_2513,N_2240,N_2377);
xor U2514 (N_2514,N_2365,N_2067);
or U2515 (N_2515,N_2286,N_2071);
nor U2516 (N_2516,N_2363,N_2037);
and U2517 (N_2517,N_2489,N_2437);
nand U2518 (N_2518,N_2168,N_2124);
nor U2519 (N_2519,N_2066,N_2090);
nand U2520 (N_2520,N_2083,N_2183);
nand U2521 (N_2521,N_2043,N_2211);
xnor U2522 (N_2522,N_2372,N_2431);
or U2523 (N_2523,N_2213,N_2140);
and U2524 (N_2524,N_2376,N_2017);
or U2525 (N_2525,N_2084,N_2026);
and U2526 (N_2526,N_2430,N_2208);
nand U2527 (N_2527,N_2441,N_2166);
or U2528 (N_2528,N_2191,N_2495);
nand U2529 (N_2529,N_2050,N_2297);
or U2530 (N_2530,N_2072,N_2147);
nand U2531 (N_2531,N_2223,N_2389);
nor U2532 (N_2532,N_2417,N_2467);
and U2533 (N_2533,N_2406,N_2359);
or U2534 (N_2534,N_2302,N_2410);
nor U2535 (N_2535,N_2362,N_2224);
nor U2536 (N_2536,N_2241,N_2231);
nor U2537 (N_2537,N_2347,N_2261);
or U2538 (N_2538,N_2475,N_2190);
nand U2539 (N_2539,N_2453,N_2051);
nor U2540 (N_2540,N_2222,N_2141);
nand U2541 (N_2541,N_2341,N_2420);
or U2542 (N_2542,N_2474,N_2275);
or U2543 (N_2543,N_2257,N_2122);
xor U2544 (N_2544,N_2198,N_2271);
or U2545 (N_2545,N_2137,N_2465);
nand U2546 (N_2546,N_2314,N_2016);
nand U2547 (N_2547,N_2234,N_2295);
xor U2548 (N_2548,N_2278,N_2352);
and U2549 (N_2549,N_2119,N_2434);
nor U2550 (N_2550,N_2149,N_2024);
or U2551 (N_2551,N_2139,N_2323);
and U2552 (N_2552,N_2447,N_2205);
and U2553 (N_2553,N_2276,N_2233);
nand U2554 (N_2554,N_2326,N_2367);
or U2555 (N_2555,N_2053,N_2446);
nor U2556 (N_2556,N_2209,N_2401);
and U2557 (N_2557,N_2157,N_2151);
or U2558 (N_2558,N_2288,N_2044);
and U2559 (N_2559,N_2282,N_2337);
nor U2560 (N_2560,N_2007,N_2138);
nor U2561 (N_2561,N_2109,N_2445);
or U2562 (N_2562,N_2184,N_2468);
nand U2563 (N_2563,N_2329,N_2306);
nor U2564 (N_2564,N_2448,N_2207);
or U2565 (N_2565,N_2079,N_2128);
nor U2566 (N_2566,N_2309,N_2332);
nor U2567 (N_2567,N_2269,N_2415);
and U2568 (N_2568,N_2159,N_2035);
and U2569 (N_2569,N_2313,N_2496);
nor U2570 (N_2570,N_2498,N_2186);
and U2571 (N_2571,N_2433,N_2093);
or U2572 (N_2572,N_2330,N_2200);
and U2573 (N_2573,N_2478,N_2492);
and U2574 (N_2574,N_2413,N_2350);
nand U2575 (N_2575,N_2015,N_2065);
nor U2576 (N_2576,N_2246,N_2253);
and U2577 (N_2577,N_2387,N_2252);
nand U2578 (N_2578,N_2038,N_2206);
and U2579 (N_2579,N_2245,N_2345);
and U2580 (N_2580,N_2167,N_2268);
nor U2581 (N_2581,N_2366,N_2423);
nor U2582 (N_2582,N_2098,N_2155);
nand U2583 (N_2583,N_2199,N_2236);
or U2584 (N_2584,N_2439,N_2456);
nand U2585 (N_2585,N_2108,N_2123);
or U2586 (N_2586,N_2412,N_2349);
xnor U2587 (N_2587,N_2392,N_2148);
and U2588 (N_2588,N_2449,N_2325);
nor U2589 (N_2589,N_2266,N_2114);
nand U2590 (N_2590,N_2006,N_2409);
and U2591 (N_2591,N_2146,N_2384);
nand U2592 (N_2592,N_2432,N_2440);
nand U2593 (N_2593,N_2466,N_2444);
and U2594 (N_2594,N_2331,N_2228);
xnor U2595 (N_2595,N_2361,N_2092);
nor U2596 (N_2596,N_2005,N_2283);
nand U2597 (N_2597,N_2391,N_2086);
or U2598 (N_2598,N_2277,N_2102);
and U2599 (N_2599,N_2394,N_2379);
nor U2600 (N_2600,N_2303,N_2356);
nand U2601 (N_2601,N_2239,N_2103);
and U2602 (N_2602,N_2235,N_2442);
xnor U2603 (N_2603,N_2076,N_2009);
nand U2604 (N_2604,N_2134,N_2068);
xor U2605 (N_2605,N_2197,N_2457);
nand U2606 (N_2606,N_2491,N_2061);
nor U2607 (N_2607,N_2482,N_2486);
or U2608 (N_2608,N_2304,N_2059);
nor U2609 (N_2609,N_2497,N_2493);
or U2610 (N_2610,N_2192,N_2471);
nor U2611 (N_2611,N_2202,N_2133);
nor U2612 (N_2612,N_2402,N_2374);
nor U2613 (N_2613,N_2256,N_2262);
nand U2614 (N_2614,N_2291,N_2225);
nor U2615 (N_2615,N_2057,N_2487);
or U2616 (N_2616,N_2088,N_2120);
nor U2617 (N_2617,N_2311,N_2230);
nor U2618 (N_2618,N_2294,N_2336);
xnor U2619 (N_2619,N_2034,N_2382);
xnor U2620 (N_2620,N_2244,N_2408);
nor U2621 (N_2621,N_2259,N_2381);
nand U2622 (N_2622,N_2054,N_2210);
nand U2623 (N_2623,N_2369,N_2110);
nand U2624 (N_2624,N_2390,N_2477);
nand U2625 (N_2625,N_2055,N_2081);
and U2626 (N_2626,N_2307,N_2364);
xor U2627 (N_2627,N_2082,N_2116);
or U2628 (N_2628,N_2339,N_2499);
nand U2629 (N_2629,N_2025,N_2154);
xnor U2630 (N_2630,N_2135,N_2164);
and U2631 (N_2631,N_2106,N_2263);
xor U2632 (N_2632,N_2033,N_2293);
xnor U2633 (N_2633,N_2020,N_2435);
nand U2634 (N_2634,N_2046,N_2237);
nand U2635 (N_2635,N_2274,N_2127);
nor U2636 (N_2636,N_2204,N_2075);
nor U2637 (N_2637,N_2370,N_2187);
nand U2638 (N_2638,N_2115,N_2042);
nand U2639 (N_2639,N_2426,N_2170);
nor U2640 (N_2640,N_2194,N_2319);
nor U2641 (N_2641,N_2112,N_2255);
and U2642 (N_2642,N_2094,N_2156);
or U2643 (N_2643,N_2188,N_2398);
and U2644 (N_2644,N_2182,N_2411);
or U2645 (N_2645,N_2162,N_2250);
xnor U2646 (N_2646,N_2405,N_2480);
or U2647 (N_2647,N_2279,N_2320);
and U2648 (N_2648,N_2342,N_2327);
and U2649 (N_2649,N_2039,N_2056);
and U2650 (N_2650,N_2344,N_2158);
xnor U2651 (N_2651,N_2028,N_2021);
or U2652 (N_2652,N_2479,N_2403);
nand U2653 (N_2653,N_2064,N_2041);
nor U2654 (N_2654,N_2196,N_2011);
nor U2655 (N_2655,N_2258,N_2380);
nand U2656 (N_2656,N_2425,N_2142);
and U2657 (N_2657,N_2008,N_2060);
and U2658 (N_2658,N_2203,N_2179);
nand U2659 (N_2659,N_2218,N_2251);
nor U2660 (N_2660,N_2216,N_2399);
or U2661 (N_2661,N_2227,N_2130);
and U2662 (N_2662,N_2414,N_2049);
nor U2663 (N_2663,N_2284,N_2385);
nor U2664 (N_2664,N_2404,N_2273);
nor U2665 (N_2665,N_2328,N_2305);
nor U2666 (N_2666,N_2464,N_2317);
nand U2667 (N_2667,N_2058,N_2104);
or U2668 (N_2668,N_2287,N_2285);
and U2669 (N_2669,N_2221,N_2312);
and U2670 (N_2670,N_2040,N_2338);
nand U2671 (N_2671,N_2238,N_2476);
nor U2672 (N_2672,N_2032,N_2107);
nand U2673 (N_2673,N_2243,N_2152);
and U2674 (N_2674,N_2018,N_2462);
and U2675 (N_2675,N_2163,N_2185);
nor U2676 (N_2676,N_2036,N_2219);
nor U2677 (N_2677,N_2248,N_2217);
nor U2678 (N_2678,N_2173,N_2111);
or U2679 (N_2679,N_2407,N_2171);
nor U2680 (N_2680,N_2085,N_2469);
and U2681 (N_2681,N_2396,N_2281);
nand U2682 (N_2682,N_2193,N_2069);
or U2683 (N_2683,N_2355,N_2165);
nand U2684 (N_2684,N_2176,N_2299);
xor U2685 (N_2685,N_2454,N_2030);
nor U2686 (N_2686,N_2220,N_2343);
nand U2687 (N_2687,N_2129,N_2091);
or U2688 (N_2688,N_2484,N_2031);
and U2689 (N_2689,N_2153,N_2027);
or U2690 (N_2690,N_2428,N_2333);
nand U2691 (N_2691,N_2419,N_2136);
xor U2692 (N_2692,N_2013,N_2292);
and U2693 (N_2693,N_2003,N_2161);
nor U2694 (N_2694,N_2375,N_2178);
nor U2695 (N_2695,N_2451,N_2436);
or U2696 (N_2696,N_2145,N_2169);
or U2697 (N_2697,N_2463,N_2290);
or U2698 (N_2698,N_2265,N_2310);
or U2699 (N_2699,N_2080,N_2022);
and U2700 (N_2700,N_2247,N_2023);
nand U2701 (N_2701,N_2483,N_2229);
and U2702 (N_2702,N_2180,N_2117);
nand U2703 (N_2703,N_2455,N_2019);
or U2704 (N_2704,N_2400,N_2070);
nand U2705 (N_2705,N_2450,N_2490);
or U2706 (N_2706,N_2316,N_2485);
nor U2707 (N_2707,N_2357,N_2063);
xor U2708 (N_2708,N_2010,N_2105);
nand U2709 (N_2709,N_2368,N_2301);
nand U2710 (N_2710,N_2346,N_2334);
or U2711 (N_2711,N_2300,N_2089);
and U2712 (N_2712,N_2232,N_2077);
and U2713 (N_2713,N_2048,N_2118);
nand U2714 (N_2714,N_2260,N_2289);
nor U2715 (N_2715,N_2249,N_2393);
or U2716 (N_2716,N_2308,N_2264);
nand U2717 (N_2717,N_2452,N_2473);
and U2718 (N_2718,N_2358,N_2378);
or U2719 (N_2719,N_2132,N_2189);
nand U2720 (N_2720,N_2422,N_2386);
or U2721 (N_2721,N_2087,N_2096);
nor U2722 (N_2722,N_2315,N_2296);
and U2723 (N_2723,N_2160,N_2004);
nand U2724 (N_2724,N_2078,N_2052);
or U2725 (N_2725,N_2143,N_2298);
nor U2726 (N_2726,N_2012,N_2100);
xor U2727 (N_2727,N_2360,N_2172);
and U2728 (N_2728,N_2174,N_2373);
nor U2729 (N_2729,N_2429,N_2371);
xnor U2730 (N_2730,N_2215,N_2340);
or U2731 (N_2731,N_2181,N_2318);
nor U2732 (N_2732,N_2195,N_2280);
or U2733 (N_2733,N_2397,N_2214);
and U2734 (N_2734,N_2421,N_2458);
and U2735 (N_2735,N_2062,N_2461);
nand U2736 (N_2736,N_2175,N_2348);
or U2737 (N_2737,N_2177,N_2322);
nand U2738 (N_2738,N_2267,N_2481);
and U2739 (N_2739,N_2254,N_2029);
xnor U2740 (N_2740,N_2242,N_2201);
nor U2741 (N_2741,N_2097,N_2488);
nand U2742 (N_2742,N_2353,N_2099);
nand U2743 (N_2743,N_2335,N_2438);
nand U2744 (N_2744,N_2427,N_2144);
or U2745 (N_2745,N_2424,N_2212);
nor U2746 (N_2746,N_2351,N_2047);
or U2747 (N_2747,N_2494,N_2131);
and U2748 (N_2748,N_2226,N_2388);
xnor U2749 (N_2749,N_2002,N_2324);
nor U2750 (N_2750,N_2057,N_2044);
nor U2751 (N_2751,N_2461,N_2418);
or U2752 (N_2752,N_2066,N_2050);
or U2753 (N_2753,N_2367,N_2198);
nand U2754 (N_2754,N_2416,N_2358);
nand U2755 (N_2755,N_2269,N_2480);
or U2756 (N_2756,N_2285,N_2300);
nor U2757 (N_2757,N_2415,N_2410);
nand U2758 (N_2758,N_2009,N_2360);
nand U2759 (N_2759,N_2393,N_2361);
or U2760 (N_2760,N_2263,N_2450);
nor U2761 (N_2761,N_2406,N_2166);
or U2762 (N_2762,N_2453,N_2034);
or U2763 (N_2763,N_2251,N_2288);
xnor U2764 (N_2764,N_2151,N_2422);
or U2765 (N_2765,N_2272,N_2125);
nor U2766 (N_2766,N_2258,N_2279);
xnor U2767 (N_2767,N_2448,N_2264);
and U2768 (N_2768,N_2429,N_2417);
xor U2769 (N_2769,N_2484,N_2417);
or U2770 (N_2770,N_2159,N_2395);
or U2771 (N_2771,N_2449,N_2053);
and U2772 (N_2772,N_2310,N_2206);
xnor U2773 (N_2773,N_2353,N_2351);
nand U2774 (N_2774,N_2191,N_2275);
nor U2775 (N_2775,N_2271,N_2320);
xnor U2776 (N_2776,N_2414,N_2263);
nor U2777 (N_2777,N_2054,N_2052);
and U2778 (N_2778,N_2487,N_2222);
or U2779 (N_2779,N_2071,N_2199);
or U2780 (N_2780,N_2121,N_2068);
nand U2781 (N_2781,N_2017,N_2358);
or U2782 (N_2782,N_2342,N_2128);
nor U2783 (N_2783,N_2269,N_2291);
nand U2784 (N_2784,N_2314,N_2181);
or U2785 (N_2785,N_2400,N_2214);
and U2786 (N_2786,N_2035,N_2382);
nand U2787 (N_2787,N_2135,N_2086);
nor U2788 (N_2788,N_2086,N_2399);
nor U2789 (N_2789,N_2030,N_2429);
and U2790 (N_2790,N_2317,N_2349);
xnor U2791 (N_2791,N_2223,N_2112);
nor U2792 (N_2792,N_2499,N_2099);
or U2793 (N_2793,N_2311,N_2474);
or U2794 (N_2794,N_2078,N_2252);
or U2795 (N_2795,N_2281,N_2095);
or U2796 (N_2796,N_2485,N_2094);
or U2797 (N_2797,N_2333,N_2038);
nor U2798 (N_2798,N_2194,N_2071);
nand U2799 (N_2799,N_2024,N_2300);
or U2800 (N_2800,N_2132,N_2016);
nor U2801 (N_2801,N_2497,N_2052);
nor U2802 (N_2802,N_2182,N_2194);
nand U2803 (N_2803,N_2229,N_2054);
nor U2804 (N_2804,N_2386,N_2431);
and U2805 (N_2805,N_2134,N_2433);
or U2806 (N_2806,N_2169,N_2097);
or U2807 (N_2807,N_2380,N_2059);
and U2808 (N_2808,N_2003,N_2475);
and U2809 (N_2809,N_2033,N_2113);
nand U2810 (N_2810,N_2318,N_2371);
and U2811 (N_2811,N_2001,N_2496);
nor U2812 (N_2812,N_2065,N_2259);
or U2813 (N_2813,N_2088,N_2300);
and U2814 (N_2814,N_2023,N_2443);
and U2815 (N_2815,N_2374,N_2138);
and U2816 (N_2816,N_2023,N_2169);
and U2817 (N_2817,N_2215,N_2188);
and U2818 (N_2818,N_2112,N_2235);
xor U2819 (N_2819,N_2111,N_2148);
nor U2820 (N_2820,N_2374,N_2083);
nand U2821 (N_2821,N_2306,N_2356);
nor U2822 (N_2822,N_2401,N_2412);
and U2823 (N_2823,N_2081,N_2414);
nand U2824 (N_2824,N_2159,N_2194);
nand U2825 (N_2825,N_2416,N_2226);
and U2826 (N_2826,N_2272,N_2048);
nor U2827 (N_2827,N_2260,N_2016);
and U2828 (N_2828,N_2003,N_2354);
nor U2829 (N_2829,N_2201,N_2341);
nor U2830 (N_2830,N_2221,N_2227);
nor U2831 (N_2831,N_2200,N_2263);
and U2832 (N_2832,N_2421,N_2225);
nor U2833 (N_2833,N_2437,N_2114);
xnor U2834 (N_2834,N_2385,N_2099);
and U2835 (N_2835,N_2273,N_2191);
nor U2836 (N_2836,N_2385,N_2123);
and U2837 (N_2837,N_2011,N_2359);
and U2838 (N_2838,N_2472,N_2100);
nand U2839 (N_2839,N_2087,N_2227);
nor U2840 (N_2840,N_2494,N_2336);
or U2841 (N_2841,N_2191,N_2416);
xnor U2842 (N_2842,N_2378,N_2382);
xor U2843 (N_2843,N_2133,N_2296);
nor U2844 (N_2844,N_2417,N_2243);
nand U2845 (N_2845,N_2328,N_2050);
or U2846 (N_2846,N_2394,N_2031);
nand U2847 (N_2847,N_2267,N_2260);
or U2848 (N_2848,N_2385,N_2143);
nor U2849 (N_2849,N_2304,N_2204);
nor U2850 (N_2850,N_2454,N_2202);
and U2851 (N_2851,N_2278,N_2012);
xor U2852 (N_2852,N_2071,N_2478);
or U2853 (N_2853,N_2134,N_2450);
nor U2854 (N_2854,N_2126,N_2087);
nor U2855 (N_2855,N_2082,N_2074);
nand U2856 (N_2856,N_2284,N_2157);
and U2857 (N_2857,N_2408,N_2155);
and U2858 (N_2858,N_2007,N_2457);
nand U2859 (N_2859,N_2216,N_2224);
or U2860 (N_2860,N_2195,N_2453);
nor U2861 (N_2861,N_2049,N_2011);
or U2862 (N_2862,N_2245,N_2182);
and U2863 (N_2863,N_2402,N_2338);
and U2864 (N_2864,N_2379,N_2033);
nor U2865 (N_2865,N_2462,N_2086);
nand U2866 (N_2866,N_2411,N_2303);
or U2867 (N_2867,N_2282,N_2286);
and U2868 (N_2868,N_2218,N_2088);
nand U2869 (N_2869,N_2022,N_2269);
nand U2870 (N_2870,N_2079,N_2368);
xnor U2871 (N_2871,N_2217,N_2486);
or U2872 (N_2872,N_2321,N_2040);
nand U2873 (N_2873,N_2343,N_2122);
nor U2874 (N_2874,N_2402,N_2315);
and U2875 (N_2875,N_2270,N_2444);
nand U2876 (N_2876,N_2346,N_2225);
nand U2877 (N_2877,N_2457,N_2383);
xnor U2878 (N_2878,N_2438,N_2012);
nand U2879 (N_2879,N_2275,N_2220);
nor U2880 (N_2880,N_2135,N_2344);
xor U2881 (N_2881,N_2059,N_2470);
or U2882 (N_2882,N_2267,N_2468);
nand U2883 (N_2883,N_2145,N_2459);
or U2884 (N_2884,N_2371,N_2354);
nor U2885 (N_2885,N_2199,N_2421);
nand U2886 (N_2886,N_2061,N_2317);
nand U2887 (N_2887,N_2451,N_2076);
or U2888 (N_2888,N_2136,N_2139);
nand U2889 (N_2889,N_2243,N_2443);
nor U2890 (N_2890,N_2376,N_2405);
xor U2891 (N_2891,N_2042,N_2002);
or U2892 (N_2892,N_2318,N_2321);
nand U2893 (N_2893,N_2302,N_2345);
xnor U2894 (N_2894,N_2104,N_2087);
or U2895 (N_2895,N_2387,N_2243);
nor U2896 (N_2896,N_2238,N_2256);
nand U2897 (N_2897,N_2455,N_2136);
or U2898 (N_2898,N_2421,N_2481);
or U2899 (N_2899,N_2461,N_2008);
nor U2900 (N_2900,N_2403,N_2379);
and U2901 (N_2901,N_2135,N_2210);
and U2902 (N_2902,N_2088,N_2208);
xor U2903 (N_2903,N_2451,N_2478);
nand U2904 (N_2904,N_2204,N_2202);
or U2905 (N_2905,N_2375,N_2097);
nand U2906 (N_2906,N_2321,N_2469);
or U2907 (N_2907,N_2198,N_2409);
nand U2908 (N_2908,N_2030,N_2348);
and U2909 (N_2909,N_2473,N_2466);
and U2910 (N_2910,N_2115,N_2421);
xnor U2911 (N_2911,N_2176,N_2052);
nor U2912 (N_2912,N_2021,N_2241);
nand U2913 (N_2913,N_2227,N_2038);
xor U2914 (N_2914,N_2262,N_2299);
nand U2915 (N_2915,N_2053,N_2097);
nand U2916 (N_2916,N_2105,N_2197);
nand U2917 (N_2917,N_2118,N_2250);
or U2918 (N_2918,N_2338,N_2240);
nor U2919 (N_2919,N_2396,N_2435);
and U2920 (N_2920,N_2193,N_2424);
nor U2921 (N_2921,N_2456,N_2352);
or U2922 (N_2922,N_2366,N_2329);
or U2923 (N_2923,N_2229,N_2232);
or U2924 (N_2924,N_2436,N_2407);
or U2925 (N_2925,N_2168,N_2073);
or U2926 (N_2926,N_2030,N_2289);
nor U2927 (N_2927,N_2114,N_2301);
nor U2928 (N_2928,N_2300,N_2052);
or U2929 (N_2929,N_2266,N_2231);
nor U2930 (N_2930,N_2217,N_2084);
or U2931 (N_2931,N_2424,N_2425);
or U2932 (N_2932,N_2458,N_2006);
nor U2933 (N_2933,N_2464,N_2035);
xor U2934 (N_2934,N_2428,N_2490);
nor U2935 (N_2935,N_2456,N_2375);
nand U2936 (N_2936,N_2309,N_2163);
xnor U2937 (N_2937,N_2363,N_2105);
and U2938 (N_2938,N_2338,N_2323);
nor U2939 (N_2939,N_2016,N_2226);
or U2940 (N_2940,N_2255,N_2009);
xnor U2941 (N_2941,N_2465,N_2045);
and U2942 (N_2942,N_2198,N_2417);
and U2943 (N_2943,N_2110,N_2202);
and U2944 (N_2944,N_2019,N_2199);
and U2945 (N_2945,N_2068,N_2333);
nor U2946 (N_2946,N_2482,N_2084);
nor U2947 (N_2947,N_2031,N_2236);
nor U2948 (N_2948,N_2361,N_2201);
or U2949 (N_2949,N_2286,N_2382);
and U2950 (N_2950,N_2368,N_2256);
nand U2951 (N_2951,N_2357,N_2204);
nor U2952 (N_2952,N_2480,N_2006);
or U2953 (N_2953,N_2447,N_2339);
or U2954 (N_2954,N_2392,N_2427);
xnor U2955 (N_2955,N_2114,N_2310);
nand U2956 (N_2956,N_2469,N_2170);
nand U2957 (N_2957,N_2132,N_2105);
and U2958 (N_2958,N_2160,N_2081);
or U2959 (N_2959,N_2055,N_2360);
and U2960 (N_2960,N_2190,N_2292);
nand U2961 (N_2961,N_2039,N_2404);
or U2962 (N_2962,N_2200,N_2248);
and U2963 (N_2963,N_2290,N_2040);
xnor U2964 (N_2964,N_2466,N_2088);
nor U2965 (N_2965,N_2303,N_2024);
nand U2966 (N_2966,N_2121,N_2210);
nand U2967 (N_2967,N_2328,N_2194);
and U2968 (N_2968,N_2218,N_2188);
xor U2969 (N_2969,N_2399,N_2304);
nor U2970 (N_2970,N_2014,N_2036);
xor U2971 (N_2971,N_2053,N_2241);
nor U2972 (N_2972,N_2058,N_2303);
and U2973 (N_2973,N_2071,N_2122);
or U2974 (N_2974,N_2230,N_2277);
and U2975 (N_2975,N_2427,N_2256);
xnor U2976 (N_2976,N_2471,N_2362);
nor U2977 (N_2977,N_2042,N_2075);
or U2978 (N_2978,N_2202,N_2125);
nor U2979 (N_2979,N_2022,N_2381);
nor U2980 (N_2980,N_2097,N_2478);
nand U2981 (N_2981,N_2336,N_2366);
nor U2982 (N_2982,N_2136,N_2454);
nor U2983 (N_2983,N_2268,N_2239);
xnor U2984 (N_2984,N_2128,N_2333);
and U2985 (N_2985,N_2160,N_2391);
and U2986 (N_2986,N_2277,N_2119);
or U2987 (N_2987,N_2359,N_2211);
nand U2988 (N_2988,N_2167,N_2118);
or U2989 (N_2989,N_2007,N_2489);
and U2990 (N_2990,N_2233,N_2234);
nor U2991 (N_2991,N_2239,N_2151);
nor U2992 (N_2992,N_2120,N_2069);
nor U2993 (N_2993,N_2197,N_2026);
and U2994 (N_2994,N_2188,N_2052);
or U2995 (N_2995,N_2140,N_2353);
nand U2996 (N_2996,N_2329,N_2260);
nand U2997 (N_2997,N_2418,N_2296);
nand U2998 (N_2998,N_2070,N_2006);
nor U2999 (N_2999,N_2426,N_2241);
and UO_0 (O_0,N_2541,N_2919);
and UO_1 (O_1,N_2904,N_2589);
or UO_2 (O_2,N_2552,N_2730);
nor UO_3 (O_3,N_2618,N_2538);
nand UO_4 (O_4,N_2952,N_2984);
or UO_5 (O_5,N_2850,N_2505);
and UO_6 (O_6,N_2802,N_2683);
and UO_7 (O_7,N_2985,N_2709);
nand UO_8 (O_8,N_2908,N_2955);
or UO_9 (O_9,N_2918,N_2767);
or UO_10 (O_10,N_2871,N_2579);
and UO_11 (O_11,N_2640,N_2670);
and UO_12 (O_12,N_2556,N_2916);
nand UO_13 (O_13,N_2615,N_2788);
or UO_14 (O_14,N_2858,N_2956);
nand UO_15 (O_15,N_2811,N_2612);
nor UO_16 (O_16,N_2831,N_2666);
nor UO_17 (O_17,N_2634,N_2769);
nor UO_18 (O_18,N_2617,N_2868);
nand UO_19 (O_19,N_2862,N_2905);
nand UO_20 (O_20,N_2652,N_2583);
and UO_21 (O_21,N_2582,N_2795);
and UO_22 (O_22,N_2942,N_2914);
and UO_23 (O_23,N_2792,N_2524);
xor UO_24 (O_24,N_2658,N_2772);
or UO_25 (O_25,N_2863,N_2633);
or UO_26 (O_26,N_2890,N_2716);
xor UO_27 (O_27,N_2570,N_2969);
or UO_28 (O_28,N_2963,N_2768);
nor UO_29 (O_29,N_2878,N_2674);
nor UO_30 (O_30,N_2735,N_2819);
or UO_31 (O_31,N_2758,N_2915);
or UO_32 (O_32,N_2751,N_2564);
or UO_33 (O_33,N_2877,N_2760);
or UO_34 (O_34,N_2539,N_2650);
nand UO_35 (O_35,N_2886,N_2827);
nand UO_36 (O_36,N_2693,N_2746);
nand UO_37 (O_37,N_2752,N_2742);
nor UO_38 (O_38,N_2600,N_2630);
and UO_39 (O_39,N_2697,N_2978);
and UO_40 (O_40,N_2959,N_2880);
or UO_41 (O_41,N_2786,N_2704);
nor UO_42 (O_42,N_2747,N_2722);
and UO_43 (O_43,N_2660,N_2764);
and UO_44 (O_44,N_2983,N_2950);
or UO_45 (O_45,N_2972,N_2558);
nand UO_46 (O_46,N_2691,N_2990);
or UO_47 (O_47,N_2531,N_2812);
nand UO_48 (O_48,N_2869,N_2563);
nor UO_49 (O_49,N_2585,N_2551);
nor UO_50 (O_50,N_2514,N_2519);
or UO_51 (O_51,N_2961,N_2870);
or UO_52 (O_52,N_2997,N_2866);
nor UO_53 (O_53,N_2999,N_2835);
nand UO_54 (O_54,N_2912,N_2989);
nor UO_55 (O_55,N_2938,N_2940);
nand UO_56 (O_56,N_2976,N_2561);
or UO_57 (O_57,N_2794,N_2529);
or UO_58 (O_58,N_2718,N_2549);
and UO_59 (O_59,N_2909,N_2766);
xor UO_60 (O_60,N_2613,N_2619);
and UO_61 (O_61,N_2554,N_2864);
nor UO_62 (O_62,N_2667,N_2995);
xnor UO_63 (O_63,N_2713,N_2951);
and UO_64 (O_64,N_2726,N_2793);
xor UO_65 (O_65,N_2857,N_2837);
and UO_66 (O_66,N_2702,N_2671);
nor UO_67 (O_67,N_2939,N_2875);
nand UO_68 (O_68,N_2987,N_2818);
or UO_69 (O_69,N_2889,N_2700);
nor UO_70 (O_70,N_2892,N_2816);
nand UO_71 (O_71,N_2848,N_2879);
and UO_72 (O_72,N_2991,N_2679);
xnor UO_73 (O_73,N_2616,N_2611);
nor UO_74 (O_74,N_2913,N_2993);
nor UO_75 (O_75,N_2572,N_2902);
nand UO_76 (O_76,N_2946,N_2609);
nor UO_77 (O_77,N_2928,N_2607);
xnor UO_78 (O_78,N_2631,N_2703);
or UO_79 (O_79,N_2724,N_2966);
xnor UO_80 (O_80,N_2810,N_2622);
nand UO_81 (O_81,N_2753,N_2729);
or UO_82 (O_82,N_2555,N_2646);
nor UO_83 (O_83,N_2967,N_2673);
and UO_84 (O_84,N_2771,N_2936);
and UO_85 (O_85,N_2744,N_2834);
or UO_86 (O_86,N_2645,N_2559);
nand UO_87 (O_87,N_2755,N_2822);
nand UO_88 (O_88,N_2521,N_2533);
or UO_89 (O_89,N_2506,N_2575);
or UO_90 (O_90,N_2856,N_2924);
nor UO_91 (O_91,N_2553,N_2785);
nor UO_92 (O_92,N_2605,N_2637);
nor UO_93 (O_93,N_2720,N_2860);
nor UO_94 (O_94,N_2784,N_2896);
and UO_95 (O_95,N_2900,N_2820);
nand UO_96 (O_96,N_2632,N_2728);
nand UO_97 (O_97,N_2895,N_2920);
and UO_98 (O_98,N_2690,N_2849);
and UO_99 (O_99,N_2845,N_2664);
nand UO_100 (O_100,N_2933,N_2780);
or UO_101 (O_101,N_2762,N_2901);
nor UO_102 (O_102,N_2872,N_2705);
or UO_103 (O_103,N_2659,N_2948);
nand UO_104 (O_104,N_2765,N_2750);
nand UO_105 (O_105,N_2839,N_2584);
and UO_106 (O_106,N_2960,N_2921);
or UO_107 (O_107,N_2844,N_2814);
and UO_108 (O_108,N_2687,N_2782);
or UO_109 (O_109,N_2642,N_2894);
and UO_110 (O_110,N_2668,N_2715);
and UO_111 (O_111,N_2958,N_2757);
nor UO_112 (O_112,N_2635,N_2681);
nor UO_113 (O_113,N_2798,N_2843);
and UO_114 (O_114,N_2534,N_2931);
and UO_115 (O_115,N_2624,N_2712);
nand UO_116 (O_116,N_2917,N_2677);
nand UO_117 (O_117,N_2692,N_2675);
nor UO_118 (O_118,N_2754,N_2801);
nand UO_119 (O_119,N_2628,N_2927);
xnor UO_120 (O_120,N_2592,N_2580);
or UO_121 (O_121,N_2520,N_2898);
or UO_122 (O_122,N_2906,N_2593);
or UO_123 (O_123,N_2610,N_2682);
or UO_124 (O_124,N_2595,N_2560);
or UO_125 (O_125,N_2644,N_2779);
and UO_126 (O_126,N_2964,N_2528);
nor UO_127 (O_127,N_2789,N_2817);
and UO_128 (O_128,N_2523,N_2803);
or UO_129 (O_129,N_2513,N_2945);
xnor UO_130 (O_130,N_2832,N_2508);
nor UO_131 (O_131,N_2708,N_2680);
xnor UO_132 (O_132,N_2926,N_2694);
or UO_133 (O_133,N_2651,N_2525);
and UO_134 (O_134,N_2623,N_2606);
xnor UO_135 (O_135,N_2778,N_2587);
nand UO_136 (O_136,N_2851,N_2594);
and UO_137 (O_137,N_2581,N_2970);
nor UO_138 (O_138,N_2689,N_2669);
and UO_139 (O_139,N_2865,N_2907);
xnor UO_140 (O_140,N_2806,N_2661);
and UO_141 (O_141,N_2500,N_2929);
nor UO_142 (O_142,N_2867,N_2602);
nand UO_143 (O_143,N_2711,N_2821);
nor UO_144 (O_144,N_2740,N_2852);
or UO_145 (O_145,N_2887,N_2725);
and UO_146 (O_146,N_2504,N_2608);
nor UO_147 (O_147,N_2992,N_2597);
and UO_148 (O_148,N_2947,N_2885);
and UO_149 (O_149,N_2808,N_2629);
nor UO_150 (O_150,N_2599,N_2626);
nor UO_151 (O_151,N_2957,N_2676);
or UO_152 (O_152,N_2973,N_2698);
nand UO_153 (O_153,N_2734,N_2743);
nand UO_154 (O_154,N_2568,N_2535);
and UO_155 (O_155,N_2893,N_2853);
xnor UO_156 (O_156,N_2546,N_2965);
or UO_157 (O_157,N_2761,N_2986);
and UO_158 (O_158,N_2790,N_2620);
and UO_159 (O_159,N_2515,N_2897);
nand UO_160 (O_160,N_2737,N_2756);
nor UO_161 (O_161,N_2799,N_2569);
or UO_162 (O_162,N_2807,N_2510);
nand UO_163 (O_163,N_2684,N_2688);
nor UO_164 (O_164,N_2748,N_2596);
and UO_165 (O_165,N_2815,N_2565);
nor UO_166 (O_166,N_2826,N_2621);
or UO_167 (O_167,N_2643,N_2547);
nand UO_168 (O_168,N_2836,N_2502);
xnor UO_169 (O_169,N_2935,N_2923);
nor UO_170 (O_170,N_2598,N_2977);
nand UO_171 (O_171,N_2943,N_2962);
and UO_172 (O_172,N_2882,N_2516);
nand UO_173 (O_173,N_2578,N_2603);
nand UO_174 (O_174,N_2557,N_2823);
nor UO_175 (O_175,N_2988,N_2588);
nor UO_176 (O_176,N_2562,N_2522);
xnor UO_177 (O_177,N_2614,N_2566);
nor UO_178 (O_178,N_2574,N_2625);
nand UO_179 (O_179,N_2861,N_2544);
nand UO_180 (O_180,N_2517,N_2731);
or UO_181 (O_181,N_2974,N_2774);
xor UO_182 (O_182,N_2672,N_2749);
or UO_183 (O_183,N_2888,N_2759);
nor UO_184 (O_184,N_2571,N_2797);
and UO_185 (O_185,N_2873,N_2706);
nand UO_186 (O_186,N_2655,N_2639);
or UO_187 (O_187,N_2507,N_2859);
or UO_188 (O_188,N_2663,N_2512);
and UO_189 (O_189,N_2841,N_2548);
nor UO_190 (O_190,N_2738,N_2719);
and UO_191 (O_191,N_2590,N_2922);
xor UO_192 (O_192,N_2805,N_2739);
nor UO_193 (O_193,N_2911,N_2653);
nand UO_194 (O_194,N_2994,N_2604);
and UO_195 (O_195,N_2511,N_2770);
and UO_196 (O_196,N_2833,N_2696);
and UO_197 (O_197,N_2874,N_2733);
nand UO_198 (O_198,N_2601,N_2787);
nand UO_199 (O_199,N_2781,N_2540);
and UO_200 (O_200,N_2884,N_2775);
or UO_201 (O_201,N_2981,N_2518);
nand UO_202 (O_202,N_2876,N_2550);
and UO_203 (O_203,N_2649,N_2745);
nand UO_204 (O_204,N_2654,N_2537);
and UO_205 (O_205,N_2526,N_2883);
and UO_206 (O_206,N_2838,N_2910);
or UO_207 (O_207,N_2527,N_2809);
xnor UO_208 (O_208,N_2727,N_2846);
nand UO_209 (O_209,N_2800,N_2699);
nor UO_210 (O_210,N_2944,N_2627);
and UO_211 (O_211,N_2847,N_2891);
xor UO_212 (O_212,N_2545,N_2685);
nor UO_213 (O_213,N_2825,N_2854);
or UO_214 (O_214,N_2828,N_2543);
xnor UO_215 (O_215,N_2968,N_2773);
and UO_216 (O_216,N_2736,N_2695);
nand UO_217 (O_217,N_2542,N_2586);
or UO_218 (O_218,N_2641,N_2855);
xor UO_219 (O_219,N_2707,N_2953);
and UO_220 (O_220,N_2656,N_2723);
and UO_221 (O_221,N_2842,N_2949);
and UO_222 (O_222,N_2934,N_2783);
or UO_223 (O_223,N_2573,N_2567);
nor UO_224 (O_224,N_2930,N_2647);
and UO_225 (O_225,N_2721,N_2982);
or UO_226 (O_226,N_2813,N_2975);
and UO_227 (O_227,N_2648,N_2678);
or UO_228 (O_228,N_2638,N_2941);
nor UO_229 (O_229,N_2530,N_2777);
nor UO_230 (O_230,N_2503,N_2717);
and UO_231 (O_231,N_2732,N_2881);
and UO_232 (O_232,N_2830,N_2577);
nor UO_233 (O_233,N_2971,N_2932);
xnor UO_234 (O_234,N_2501,N_2954);
nand UO_235 (O_235,N_2665,N_2980);
xor UO_236 (O_236,N_2576,N_2996);
nor UO_237 (O_237,N_2509,N_2796);
nor UO_238 (O_238,N_2532,N_2824);
or UO_239 (O_239,N_2925,N_2829);
nor UO_240 (O_240,N_2657,N_2536);
or UO_241 (O_241,N_2701,N_2591);
nand UO_242 (O_242,N_2791,N_2776);
and UO_243 (O_243,N_2979,N_2937);
and UO_244 (O_244,N_2686,N_2714);
and UO_245 (O_245,N_2899,N_2998);
or UO_246 (O_246,N_2804,N_2903);
nand UO_247 (O_247,N_2636,N_2763);
or UO_248 (O_248,N_2741,N_2710);
nand UO_249 (O_249,N_2840,N_2662);
xor UO_250 (O_250,N_2638,N_2712);
and UO_251 (O_251,N_2874,N_2742);
nand UO_252 (O_252,N_2856,N_2658);
xnor UO_253 (O_253,N_2675,N_2562);
nor UO_254 (O_254,N_2868,N_2699);
and UO_255 (O_255,N_2741,N_2683);
nor UO_256 (O_256,N_2805,N_2913);
or UO_257 (O_257,N_2994,N_2651);
nand UO_258 (O_258,N_2570,N_2953);
nor UO_259 (O_259,N_2908,N_2756);
nand UO_260 (O_260,N_2613,N_2737);
or UO_261 (O_261,N_2928,N_2877);
nand UO_262 (O_262,N_2547,N_2960);
nand UO_263 (O_263,N_2575,N_2553);
or UO_264 (O_264,N_2723,N_2737);
or UO_265 (O_265,N_2830,N_2530);
nand UO_266 (O_266,N_2589,N_2523);
or UO_267 (O_267,N_2807,N_2696);
or UO_268 (O_268,N_2808,N_2931);
or UO_269 (O_269,N_2507,N_2846);
xor UO_270 (O_270,N_2912,N_2760);
nor UO_271 (O_271,N_2871,N_2724);
or UO_272 (O_272,N_2811,N_2738);
or UO_273 (O_273,N_2963,N_2846);
nand UO_274 (O_274,N_2550,N_2655);
nand UO_275 (O_275,N_2638,N_2943);
nand UO_276 (O_276,N_2695,N_2605);
nor UO_277 (O_277,N_2887,N_2993);
nor UO_278 (O_278,N_2583,N_2719);
and UO_279 (O_279,N_2676,N_2545);
nor UO_280 (O_280,N_2905,N_2752);
or UO_281 (O_281,N_2888,N_2915);
and UO_282 (O_282,N_2904,N_2977);
and UO_283 (O_283,N_2558,N_2820);
nor UO_284 (O_284,N_2781,N_2868);
xnor UO_285 (O_285,N_2969,N_2573);
nand UO_286 (O_286,N_2785,N_2591);
or UO_287 (O_287,N_2837,N_2540);
nand UO_288 (O_288,N_2684,N_2565);
and UO_289 (O_289,N_2621,N_2680);
nand UO_290 (O_290,N_2890,N_2846);
nor UO_291 (O_291,N_2500,N_2587);
and UO_292 (O_292,N_2909,N_2578);
nor UO_293 (O_293,N_2685,N_2710);
nand UO_294 (O_294,N_2851,N_2604);
and UO_295 (O_295,N_2974,N_2841);
or UO_296 (O_296,N_2655,N_2668);
and UO_297 (O_297,N_2953,N_2871);
nor UO_298 (O_298,N_2606,N_2930);
nand UO_299 (O_299,N_2801,N_2987);
or UO_300 (O_300,N_2890,N_2560);
and UO_301 (O_301,N_2972,N_2857);
and UO_302 (O_302,N_2954,N_2826);
nand UO_303 (O_303,N_2741,N_2858);
nand UO_304 (O_304,N_2990,N_2606);
nor UO_305 (O_305,N_2727,N_2773);
and UO_306 (O_306,N_2679,N_2538);
nand UO_307 (O_307,N_2669,N_2612);
nand UO_308 (O_308,N_2866,N_2755);
or UO_309 (O_309,N_2895,N_2745);
nor UO_310 (O_310,N_2690,N_2904);
nand UO_311 (O_311,N_2544,N_2841);
or UO_312 (O_312,N_2699,N_2952);
nor UO_313 (O_313,N_2768,N_2664);
nor UO_314 (O_314,N_2779,N_2840);
or UO_315 (O_315,N_2531,N_2769);
or UO_316 (O_316,N_2520,N_2756);
or UO_317 (O_317,N_2974,N_2929);
or UO_318 (O_318,N_2639,N_2718);
or UO_319 (O_319,N_2854,N_2863);
nor UO_320 (O_320,N_2699,N_2608);
or UO_321 (O_321,N_2700,N_2625);
and UO_322 (O_322,N_2783,N_2906);
or UO_323 (O_323,N_2693,N_2985);
and UO_324 (O_324,N_2905,N_2515);
nand UO_325 (O_325,N_2614,N_2848);
nor UO_326 (O_326,N_2701,N_2768);
nor UO_327 (O_327,N_2559,N_2945);
and UO_328 (O_328,N_2528,N_2989);
and UO_329 (O_329,N_2967,N_2864);
xnor UO_330 (O_330,N_2794,N_2843);
nand UO_331 (O_331,N_2717,N_2599);
and UO_332 (O_332,N_2623,N_2721);
xor UO_333 (O_333,N_2515,N_2507);
or UO_334 (O_334,N_2705,N_2879);
nor UO_335 (O_335,N_2771,N_2648);
and UO_336 (O_336,N_2857,N_2532);
and UO_337 (O_337,N_2878,N_2864);
nor UO_338 (O_338,N_2875,N_2991);
nor UO_339 (O_339,N_2980,N_2831);
and UO_340 (O_340,N_2560,N_2981);
nand UO_341 (O_341,N_2661,N_2840);
xnor UO_342 (O_342,N_2977,N_2664);
nand UO_343 (O_343,N_2723,N_2516);
and UO_344 (O_344,N_2887,N_2808);
nand UO_345 (O_345,N_2655,N_2749);
nor UO_346 (O_346,N_2717,N_2879);
nand UO_347 (O_347,N_2786,N_2904);
or UO_348 (O_348,N_2931,N_2990);
nor UO_349 (O_349,N_2941,N_2789);
nand UO_350 (O_350,N_2840,N_2516);
and UO_351 (O_351,N_2774,N_2562);
and UO_352 (O_352,N_2992,N_2827);
nand UO_353 (O_353,N_2656,N_2517);
nand UO_354 (O_354,N_2511,N_2672);
nor UO_355 (O_355,N_2749,N_2877);
or UO_356 (O_356,N_2986,N_2994);
and UO_357 (O_357,N_2747,N_2850);
nand UO_358 (O_358,N_2995,N_2789);
nor UO_359 (O_359,N_2652,N_2875);
or UO_360 (O_360,N_2714,N_2544);
and UO_361 (O_361,N_2731,N_2914);
nand UO_362 (O_362,N_2511,N_2831);
and UO_363 (O_363,N_2977,N_2981);
or UO_364 (O_364,N_2518,N_2735);
or UO_365 (O_365,N_2820,N_2746);
nor UO_366 (O_366,N_2570,N_2917);
nor UO_367 (O_367,N_2736,N_2754);
nand UO_368 (O_368,N_2870,N_2812);
nor UO_369 (O_369,N_2993,N_2659);
or UO_370 (O_370,N_2519,N_2602);
nor UO_371 (O_371,N_2794,N_2953);
and UO_372 (O_372,N_2607,N_2978);
or UO_373 (O_373,N_2753,N_2549);
nand UO_374 (O_374,N_2716,N_2961);
or UO_375 (O_375,N_2798,N_2519);
or UO_376 (O_376,N_2583,N_2655);
or UO_377 (O_377,N_2513,N_2962);
nand UO_378 (O_378,N_2825,N_2652);
and UO_379 (O_379,N_2612,N_2516);
or UO_380 (O_380,N_2745,N_2653);
nor UO_381 (O_381,N_2747,N_2783);
nand UO_382 (O_382,N_2908,N_2605);
and UO_383 (O_383,N_2885,N_2533);
nand UO_384 (O_384,N_2824,N_2731);
and UO_385 (O_385,N_2885,N_2871);
and UO_386 (O_386,N_2615,N_2782);
nand UO_387 (O_387,N_2620,N_2991);
and UO_388 (O_388,N_2728,N_2888);
or UO_389 (O_389,N_2718,N_2781);
xnor UO_390 (O_390,N_2769,N_2589);
nand UO_391 (O_391,N_2980,N_2705);
or UO_392 (O_392,N_2924,N_2559);
and UO_393 (O_393,N_2640,N_2591);
nand UO_394 (O_394,N_2819,N_2617);
nor UO_395 (O_395,N_2795,N_2641);
nand UO_396 (O_396,N_2984,N_2514);
xnor UO_397 (O_397,N_2884,N_2755);
xnor UO_398 (O_398,N_2600,N_2968);
nor UO_399 (O_399,N_2975,N_2771);
and UO_400 (O_400,N_2568,N_2534);
nor UO_401 (O_401,N_2705,N_2964);
nand UO_402 (O_402,N_2928,N_2639);
xnor UO_403 (O_403,N_2852,N_2733);
nand UO_404 (O_404,N_2984,N_2688);
or UO_405 (O_405,N_2753,N_2536);
or UO_406 (O_406,N_2989,N_2947);
and UO_407 (O_407,N_2961,N_2526);
or UO_408 (O_408,N_2596,N_2747);
xnor UO_409 (O_409,N_2586,N_2621);
nor UO_410 (O_410,N_2554,N_2697);
nand UO_411 (O_411,N_2888,N_2761);
and UO_412 (O_412,N_2529,N_2876);
nand UO_413 (O_413,N_2767,N_2828);
nor UO_414 (O_414,N_2657,N_2798);
nand UO_415 (O_415,N_2929,N_2973);
xnor UO_416 (O_416,N_2720,N_2699);
nor UO_417 (O_417,N_2945,N_2618);
nand UO_418 (O_418,N_2556,N_2600);
and UO_419 (O_419,N_2508,N_2723);
nor UO_420 (O_420,N_2980,N_2578);
nand UO_421 (O_421,N_2769,N_2920);
and UO_422 (O_422,N_2756,N_2888);
nand UO_423 (O_423,N_2822,N_2969);
or UO_424 (O_424,N_2875,N_2817);
or UO_425 (O_425,N_2514,N_2805);
nor UO_426 (O_426,N_2799,N_2987);
or UO_427 (O_427,N_2919,N_2590);
nor UO_428 (O_428,N_2521,N_2920);
nor UO_429 (O_429,N_2524,N_2943);
nand UO_430 (O_430,N_2980,N_2911);
nor UO_431 (O_431,N_2939,N_2984);
or UO_432 (O_432,N_2797,N_2523);
or UO_433 (O_433,N_2794,N_2702);
nor UO_434 (O_434,N_2669,N_2701);
nand UO_435 (O_435,N_2670,N_2934);
or UO_436 (O_436,N_2926,N_2516);
nor UO_437 (O_437,N_2730,N_2644);
xnor UO_438 (O_438,N_2561,N_2673);
and UO_439 (O_439,N_2815,N_2679);
xor UO_440 (O_440,N_2912,N_2843);
and UO_441 (O_441,N_2606,N_2641);
nor UO_442 (O_442,N_2607,N_2871);
or UO_443 (O_443,N_2523,N_2682);
or UO_444 (O_444,N_2918,N_2544);
or UO_445 (O_445,N_2712,N_2823);
nand UO_446 (O_446,N_2593,N_2939);
xor UO_447 (O_447,N_2582,N_2770);
and UO_448 (O_448,N_2878,N_2949);
and UO_449 (O_449,N_2906,N_2875);
nor UO_450 (O_450,N_2567,N_2896);
nand UO_451 (O_451,N_2666,N_2609);
nor UO_452 (O_452,N_2512,N_2597);
nor UO_453 (O_453,N_2668,N_2551);
nor UO_454 (O_454,N_2594,N_2970);
or UO_455 (O_455,N_2630,N_2504);
and UO_456 (O_456,N_2578,N_2676);
nor UO_457 (O_457,N_2545,N_2576);
nand UO_458 (O_458,N_2715,N_2914);
and UO_459 (O_459,N_2763,N_2618);
or UO_460 (O_460,N_2826,N_2821);
nand UO_461 (O_461,N_2978,N_2541);
nor UO_462 (O_462,N_2805,N_2906);
nand UO_463 (O_463,N_2752,N_2681);
nor UO_464 (O_464,N_2755,N_2911);
nor UO_465 (O_465,N_2970,N_2682);
or UO_466 (O_466,N_2607,N_2938);
or UO_467 (O_467,N_2880,N_2708);
and UO_468 (O_468,N_2703,N_2777);
nand UO_469 (O_469,N_2849,N_2575);
nand UO_470 (O_470,N_2524,N_2781);
nand UO_471 (O_471,N_2573,N_2695);
and UO_472 (O_472,N_2872,N_2881);
and UO_473 (O_473,N_2637,N_2944);
and UO_474 (O_474,N_2623,N_2779);
nor UO_475 (O_475,N_2744,N_2778);
and UO_476 (O_476,N_2854,N_2504);
nand UO_477 (O_477,N_2575,N_2683);
nor UO_478 (O_478,N_2745,N_2769);
or UO_479 (O_479,N_2525,N_2719);
nand UO_480 (O_480,N_2707,N_2869);
nor UO_481 (O_481,N_2651,N_2558);
xor UO_482 (O_482,N_2622,N_2803);
and UO_483 (O_483,N_2533,N_2841);
and UO_484 (O_484,N_2735,N_2660);
and UO_485 (O_485,N_2767,N_2824);
nor UO_486 (O_486,N_2778,N_2560);
nand UO_487 (O_487,N_2990,N_2573);
and UO_488 (O_488,N_2512,N_2835);
or UO_489 (O_489,N_2731,N_2883);
nor UO_490 (O_490,N_2502,N_2847);
or UO_491 (O_491,N_2950,N_2792);
or UO_492 (O_492,N_2815,N_2783);
nand UO_493 (O_493,N_2648,N_2653);
and UO_494 (O_494,N_2890,N_2575);
xnor UO_495 (O_495,N_2993,N_2721);
or UO_496 (O_496,N_2522,N_2609);
or UO_497 (O_497,N_2999,N_2754);
or UO_498 (O_498,N_2947,N_2756);
nor UO_499 (O_499,N_2880,N_2585);
endmodule