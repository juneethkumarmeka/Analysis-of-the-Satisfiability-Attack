module basic_3000_30000_3500_15_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_718,In_2657);
xnor U1 (N_1,In_224,In_2191);
or U2 (N_2,In_252,In_896);
xor U3 (N_3,In_209,In_2552);
or U4 (N_4,In_11,In_1266);
or U5 (N_5,In_393,In_2634);
xor U6 (N_6,In_1654,In_2611);
nand U7 (N_7,In_2619,In_1234);
or U8 (N_8,In_320,In_423);
nor U9 (N_9,In_2969,In_507);
nor U10 (N_10,In_1496,In_175);
nand U11 (N_11,In_2118,In_2779);
nor U12 (N_12,In_1066,In_1252);
or U13 (N_13,In_2012,In_1959);
or U14 (N_14,In_2823,In_2160);
or U15 (N_15,In_2062,In_923);
and U16 (N_16,In_2028,In_1396);
nand U17 (N_17,In_2682,In_993);
nand U18 (N_18,In_678,In_1624);
nand U19 (N_19,In_309,In_1514);
and U20 (N_20,In_2744,In_1732);
or U21 (N_21,In_970,In_2255);
xnor U22 (N_22,In_2957,In_1416);
and U23 (N_23,In_2145,In_949);
or U24 (N_24,In_2425,In_1344);
nand U25 (N_25,In_515,In_1681);
or U26 (N_26,In_345,In_2275);
nand U27 (N_27,In_675,In_1801);
or U28 (N_28,In_1841,In_1071);
nand U29 (N_29,In_2207,In_1237);
or U30 (N_30,In_1986,In_91);
nor U31 (N_31,In_350,In_490);
xor U32 (N_32,In_259,In_2888);
xnor U33 (N_33,In_2679,In_34);
nand U34 (N_34,In_546,In_2607);
xnor U35 (N_35,In_396,In_2785);
xor U36 (N_36,In_2767,In_2471);
nor U37 (N_37,In_2421,In_426);
or U38 (N_38,In_2579,In_762);
or U39 (N_39,In_2623,In_2499);
and U40 (N_40,In_2448,In_2513);
and U41 (N_41,In_860,In_30);
and U42 (N_42,In_2060,In_2429);
nor U43 (N_43,In_461,In_2998);
and U44 (N_44,In_1610,In_402);
nor U45 (N_45,In_2587,In_1035);
nor U46 (N_46,In_1847,In_639);
xnor U47 (N_47,In_1797,In_682);
or U48 (N_48,In_2363,In_253);
nand U49 (N_49,In_316,In_198);
and U50 (N_50,In_1937,In_2885);
xnor U51 (N_51,In_2949,In_963);
xnor U52 (N_52,In_1985,In_2535);
xnor U53 (N_53,In_1042,In_1615);
or U54 (N_54,In_2104,In_2913);
nor U55 (N_55,In_1440,In_2635);
nor U56 (N_56,In_400,In_1486);
nor U57 (N_57,In_2299,In_1189);
nor U58 (N_58,In_744,In_1968);
and U59 (N_59,In_1991,In_185);
or U60 (N_60,In_2642,In_2443);
nand U61 (N_61,In_2397,In_2939);
and U62 (N_62,In_105,In_1914);
xnor U63 (N_63,In_73,In_1291);
and U64 (N_64,In_2346,In_1334);
xor U65 (N_65,In_1069,In_971);
or U66 (N_66,In_741,In_2662);
nor U67 (N_67,In_1152,In_1784);
or U68 (N_68,In_1782,In_1738);
and U69 (N_69,In_1211,In_805);
nand U70 (N_70,In_2307,In_766);
nand U71 (N_71,In_2797,In_2088);
nand U72 (N_72,In_903,In_2940);
or U73 (N_73,In_1169,In_2517);
and U74 (N_74,In_1418,In_14);
xnor U75 (N_75,In_726,In_2142);
and U76 (N_76,In_2031,In_257);
or U77 (N_77,In_2869,In_2985);
nand U78 (N_78,In_761,In_592);
nand U79 (N_79,In_2659,In_2864);
and U80 (N_80,In_1825,In_568);
or U81 (N_81,In_887,In_647);
nor U82 (N_82,In_1747,In_702);
or U83 (N_83,In_1730,In_1756);
or U84 (N_84,In_2732,In_2391);
and U85 (N_85,In_996,In_1114);
or U86 (N_86,In_1607,In_235);
nand U87 (N_87,In_2813,In_1412);
and U88 (N_88,In_1371,In_116);
xnor U89 (N_89,In_2417,In_677);
nand U90 (N_90,In_2598,In_1917);
nand U91 (N_91,In_2324,In_504);
nand U92 (N_92,In_1193,In_1158);
or U93 (N_93,In_167,In_1030);
and U94 (N_94,In_140,In_1491);
xor U95 (N_95,In_2043,In_1928);
xor U96 (N_96,In_2321,In_2845);
nand U97 (N_97,In_2546,In_403);
or U98 (N_98,In_1240,In_1389);
and U99 (N_99,In_583,In_1168);
xnor U100 (N_100,In_1280,In_551);
or U101 (N_101,In_2020,In_2734);
or U102 (N_102,In_434,In_244);
nor U103 (N_103,In_570,In_727);
xnor U104 (N_104,In_1346,In_1787);
nand U105 (N_105,In_2064,In_1668);
nor U106 (N_106,In_2234,In_1564);
nor U107 (N_107,In_35,In_219);
nor U108 (N_108,In_2412,In_848);
or U109 (N_109,In_1839,In_139);
nand U110 (N_110,In_2373,In_1622);
xnor U111 (N_111,In_1734,In_796);
nand U112 (N_112,In_894,In_2592);
nand U113 (N_113,In_1587,In_1859);
nor U114 (N_114,In_468,In_2441);
xnor U115 (N_115,In_2304,In_1325);
xor U116 (N_116,In_2453,In_1699);
nor U117 (N_117,In_531,In_918);
or U118 (N_118,In_260,In_1214);
xnor U119 (N_119,In_2449,In_2730);
nand U120 (N_120,In_453,In_1829);
or U121 (N_121,In_2035,In_2388);
nor U122 (N_122,In_2537,In_128);
nand U123 (N_123,In_2084,In_2896);
xnor U124 (N_124,In_2863,In_847);
or U125 (N_125,In_1369,In_1261);
or U126 (N_126,In_1101,In_1268);
nor U127 (N_127,In_2955,In_2743);
or U128 (N_128,In_1692,In_489);
nand U129 (N_129,In_287,In_26);
xor U130 (N_130,In_1414,In_2001);
and U131 (N_131,In_2868,In_1037);
or U132 (N_132,In_2567,In_2383);
and U133 (N_133,In_1964,In_954);
or U134 (N_134,In_496,In_829);
nand U135 (N_135,In_2105,In_2435);
xor U136 (N_136,In_1499,In_2288);
and U137 (N_137,In_2401,In_389);
and U138 (N_138,In_1793,In_588);
or U139 (N_139,In_2678,In_2958);
or U140 (N_140,In_2572,In_2353);
or U141 (N_141,In_992,In_1843);
xor U142 (N_142,In_638,In_150);
and U143 (N_143,In_1674,In_1115);
xnor U144 (N_144,In_2519,In_440);
or U145 (N_145,In_2037,In_1238);
xnor U146 (N_146,In_2811,In_513);
xor U147 (N_147,In_2948,In_2691);
nor U148 (N_148,In_1980,In_2695);
and U149 (N_149,In_2800,In_2741);
xnor U150 (N_150,In_1625,In_437);
nor U151 (N_151,In_2706,In_842);
nor U152 (N_152,In_2524,In_2230);
or U153 (N_153,In_1867,In_1804);
nand U154 (N_154,In_170,In_325);
nor U155 (N_155,In_2201,In_286);
xnor U156 (N_156,In_1792,In_2500);
nor U157 (N_157,In_876,In_2268);
and U158 (N_158,In_1011,In_79);
and U159 (N_159,In_417,In_1139);
nor U160 (N_160,In_2652,In_637);
nor U161 (N_161,In_1818,In_1285);
xor U162 (N_162,In_1679,In_2971);
or U163 (N_163,In_2256,In_240);
xnor U164 (N_164,In_545,In_2919);
and U165 (N_165,In_2338,In_1871);
nor U166 (N_166,In_977,In_1195);
or U167 (N_167,In_1576,In_1061);
xor U168 (N_168,In_1929,In_1126);
nor U169 (N_169,In_280,In_1733);
xor U170 (N_170,In_2886,In_1006);
nor U171 (N_171,In_1306,In_817);
and U172 (N_172,In_1120,In_473);
nor U173 (N_173,In_1145,In_1254);
nand U174 (N_174,In_2830,In_1803);
xor U175 (N_175,In_2467,In_2171);
xnor U176 (N_176,In_331,In_2218);
nand U177 (N_177,In_2664,In_2177);
xnor U178 (N_178,In_2228,In_2150);
nand U179 (N_179,In_2025,In_2458);
xor U180 (N_180,In_1310,In_1833);
or U181 (N_181,In_142,In_2935);
nand U182 (N_182,In_982,In_1997);
nor U183 (N_183,In_1753,In_311);
nor U184 (N_184,In_1762,In_46);
and U185 (N_185,In_905,In_1510);
xnor U186 (N_186,In_1390,In_2720);
and U187 (N_187,In_1323,In_1076);
or U188 (N_188,In_2224,In_382);
nand U189 (N_189,In_1180,In_2481);
or U190 (N_190,In_673,In_2477);
nor U191 (N_191,In_2543,In_2115);
nand U192 (N_192,In_376,In_45);
or U193 (N_193,In_1495,In_2464);
and U194 (N_194,In_522,In_2451);
and U195 (N_195,In_2596,In_874);
and U196 (N_196,In_337,In_733);
xor U197 (N_197,In_1581,In_1335);
xor U198 (N_198,In_2106,In_1439);
nor U199 (N_199,In_2157,In_2525);
and U200 (N_200,In_1933,In_1863);
and U201 (N_201,In_2496,In_2468);
or U202 (N_202,In_1994,In_2747);
or U203 (N_203,In_1527,In_1500);
and U204 (N_204,In_221,In_869);
nand U205 (N_205,In_1611,In_843);
nand U206 (N_206,In_1451,In_2236);
or U207 (N_207,In_467,In_870);
and U208 (N_208,In_2643,In_2908);
nand U209 (N_209,In_2030,In_2409);
nor U210 (N_210,In_2289,In_121);
xor U211 (N_211,In_1218,In_1653);
xor U212 (N_212,In_288,In_1813);
nor U213 (N_213,In_1472,In_505);
or U214 (N_214,In_880,In_296);
nor U215 (N_215,In_1893,In_2112);
nor U216 (N_216,In_332,In_1164);
nor U217 (N_217,In_607,In_1821);
or U218 (N_218,In_218,In_430);
xor U219 (N_219,In_2962,In_342);
or U220 (N_220,In_2238,In_2053);
xor U221 (N_221,In_940,In_2462);
nor U222 (N_222,In_657,In_2272);
and U223 (N_223,In_38,In_2193);
nand U224 (N_224,In_1864,In_2252);
nor U225 (N_225,In_1532,In_1106);
or U226 (N_226,In_854,In_2100);
nand U227 (N_227,In_196,In_1039);
or U228 (N_228,In_1050,In_2198);
nand U229 (N_229,In_2384,In_1176);
nand U230 (N_230,In_1525,In_1410);
nor U231 (N_231,In_1819,In_1952);
nor U232 (N_232,In_2622,In_614);
xor U233 (N_233,In_338,In_1122);
nand U234 (N_234,In_1689,In_2337);
nand U235 (N_235,In_2295,In_1918);
and U236 (N_236,In_1236,In_2941);
nand U237 (N_237,In_594,In_945);
nand U238 (N_238,In_1200,In_2683);
and U239 (N_239,In_1562,In_267);
and U240 (N_240,In_2707,In_1312);
xnor U241 (N_241,In_539,In_2394);
nand U242 (N_242,In_1031,In_1675);
and U243 (N_243,In_1719,In_1590);
nor U244 (N_244,In_1912,In_2648);
or U245 (N_245,In_2128,In_2347);
and U246 (N_246,In_106,In_2424);
xnor U247 (N_247,In_1661,In_1317);
and U248 (N_248,In_962,In_1380);
nand U249 (N_249,In_1349,In_1638);
or U250 (N_250,In_2372,In_133);
and U251 (N_251,In_1274,In_519);
nor U252 (N_252,In_1569,In_1503);
and U253 (N_253,In_778,In_2442);
and U254 (N_254,In_2008,In_439);
or U255 (N_255,In_104,In_1393);
nor U256 (N_256,In_1573,In_2219);
xor U257 (N_257,In_575,In_781);
xor U258 (N_258,In_2536,In_1057);
xor U259 (N_259,In_2640,In_823);
nor U260 (N_260,In_1981,In_96);
and U261 (N_261,In_1476,In_1328);
or U262 (N_262,In_1953,In_1685);
nor U263 (N_263,In_2312,In_2526);
nor U264 (N_264,In_3,In_2821);
xnor U265 (N_265,In_2984,In_112);
nand U266 (N_266,In_486,In_2170);
and U267 (N_267,In_2563,In_1643);
xnor U268 (N_268,In_1333,In_2716);
xnor U269 (N_269,In_107,In_1515);
nor U270 (N_270,In_284,In_1);
nand U271 (N_271,In_242,In_1999);
xor U272 (N_272,In_1769,In_1359);
nand U273 (N_273,In_2831,In_1905);
nor U274 (N_274,In_708,In_2260);
nor U275 (N_275,In_51,In_2791);
and U276 (N_276,In_573,In_1277);
nor U277 (N_277,In_2459,In_16);
and U278 (N_278,In_1591,In_703);
nand U279 (N_279,In_730,In_194);
or U280 (N_280,In_2922,In_1342);
or U281 (N_281,In_2848,In_208);
xnor U282 (N_282,In_1882,In_743);
nand U283 (N_283,In_1174,In_2124);
nor U284 (N_284,In_1568,In_1276);
or U285 (N_285,In_1233,In_2748);
or U286 (N_286,In_1074,In_472);
nand U287 (N_287,In_408,In_1924);
xor U288 (N_288,In_862,In_2223);
nor U289 (N_289,In_1094,In_1623);
xor U290 (N_290,In_557,In_1113);
nand U291 (N_291,In_995,In_1022);
nor U292 (N_292,In_2091,In_318);
and U293 (N_293,In_146,In_404);
and U294 (N_294,In_2708,In_956);
and U295 (N_295,In_793,In_736);
and U296 (N_296,In_523,In_2736);
nor U297 (N_297,In_2604,In_2923);
xnor U298 (N_298,In_1155,In_446);
xnor U299 (N_299,In_1130,In_563);
xnor U300 (N_300,In_2445,In_2993);
nand U301 (N_301,In_1029,In_2093);
or U302 (N_302,In_1855,In_1300);
nand U303 (N_303,In_173,In_1466);
xnor U304 (N_304,In_968,In_910);
nand U305 (N_305,In_2858,In_1243);
or U306 (N_306,In_1353,In_425);
and U307 (N_307,In_2095,In_119);
or U308 (N_308,In_143,In_1951);
and U309 (N_309,In_2309,In_2203);
nand U310 (N_310,In_81,In_2929);
or U311 (N_311,In_2614,In_2280);
nand U312 (N_312,In_1060,In_1226);
xnor U313 (N_313,In_558,In_601);
nand U314 (N_314,In_44,In_1198);
nand U315 (N_315,In_344,In_725);
nand U316 (N_316,In_2013,In_2290);
xor U317 (N_317,In_1976,In_2192);
nand U318 (N_318,In_413,In_827);
xor U319 (N_319,In_77,In_2887);
xnor U320 (N_320,In_1194,In_1707);
and U321 (N_321,In_2501,In_202);
xor U322 (N_322,In_2396,In_2658);
and U323 (N_323,In_729,In_873);
nor U324 (N_324,In_1429,In_585);
nor U325 (N_325,In_828,In_2656);
xor U326 (N_326,In_2808,In_2239);
or U327 (N_327,In_1383,In_2882);
xor U328 (N_328,In_1460,In_1776);
xor U329 (N_329,In_2773,In_749);
nor U330 (N_330,In_2788,In_1121);
xor U331 (N_331,In_1441,In_1448);
nand U332 (N_332,In_2423,In_1916);
or U333 (N_333,In_1931,In_2931);
or U334 (N_334,In_1081,In_1866);
nand U335 (N_335,In_1960,In_29);
xor U336 (N_336,In_2340,In_217);
nand U337 (N_337,In_1468,In_2076);
or U338 (N_338,In_1696,In_2943);
and U339 (N_339,In_695,In_1461);
and U340 (N_340,In_2972,In_989);
nor U341 (N_341,In_1260,In_1603);
nand U342 (N_342,In_1090,In_2533);
xor U343 (N_343,In_1606,In_1567);
nor U344 (N_344,In_1979,In_2731);
xor U345 (N_345,In_1477,In_1305);
nor U346 (N_346,In_1572,In_908);
nand U347 (N_347,In_70,In_365);
or U348 (N_348,In_2389,In_1682);
nand U349 (N_349,In_2070,In_2566);
nor U350 (N_350,In_998,In_1178);
nand U351 (N_351,In_2143,In_1505);
nand U352 (N_352,In_1432,In_1583);
and U353 (N_353,In_2475,In_39);
and U354 (N_354,In_1850,In_751);
nand U355 (N_355,In_2126,In_2291);
or U356 (N_356,In_1788,In_1352);
or U357 (N_357,In_1786,In_2505);
nor U358 (N_358,In_734,In_1593);
and U359 (N_359,In_388,In_1805);
nor U360 (N_360,In_2778,In_2410);
and U361 (N_361,In_1494,In_2632);
xnor U362 (N_362,In_1906,In_1435);
or U363 (N_363,In_1513,In_2905);
nor U364 (N_364,In_635,In_1815);
xor U365 (N_365,In_1336,In_1025);
nor U366 (N_366,In_1700,In_902);
or U367 (N_367,In_1868,In_1549);
and U368 (N_368,In_2367,In_2541);
and U369 (N_369,In_2478,In_2564);
nand U370 (N_370,In_213,In_2975);
nand U371 (N_371,In_1713,In_69);
nor U372 (N_372,In_2277,In_1190);
xor U373 (N_373,In_1018,In_470);
and U374 (N_374,In_258,In_1517);
or U375 (N_375,In_836,In_1823);
nor U376 (N_376,In_2544,In_2153);
nor U377 (N_377,In_99,In_1442);
xnor U378 (N_378,In_1473,In_2195);
nand U379 (N_379,In_2527,In_777);
or U380 (N_380,In_2322,In_1507);
nand U381 (N_381,In_2495,In_1127);
nand U382 (N_382,In_871,In_2819);
and U383 (N_383,In_2803,In_1519);
xnor U384 (N_384,In_1457,In_1015);
nor U385 (N_385,In_1487,In_891);
and U386 (N_386,In_1338,In_2586);
nor U387 (N_387,In_438,In_1715);
or U388 (N_388,In_135,In_1783);
nor U389 (N_389,In_679,In_2359);
nor U390 (N_390,In_2251,In_2220);
nand U391 (N_391,In_2974,In_609);
nand U392 (N_392,In_877,In_2173);
nand U393 (N_393,In_2063,In_436);
nand U394 (N_394,In_972,In_1571);
nand U395 (N_395,In_2103,In_2189);
or U396 (N_396,In_1563,In_1141);
nand U397 (N_397,In_1327,In_1154);
xor U398 (N_398,In_1907,In_236);
xor U399 (N_399,In_2318,In_690);
nor U400 (N_400,In_745,In_1512);
or U401 (N_401,In_394,In_172);
or U402 (N_402,In_149,In_705);
nor U403 (N_403,In_186,In_1827);
xnor U404 (N_404,In_1664,In_463);
or U405 (N_405,In_1246,In_2601);
nand U406 (N_406,In_203,In_2225);
or U407 (N_407,In_1004,In_1256);
nor U408 (N_408,In_2422,In_1750);
nand U409 (N_409,In_328,In_1550);
xor U410 (N_410,In_1215,In_2071);
nor U411 (N_411,In_549,In_562);
xnor U412 (N_412,In_844,In_986);
nand U413 (N_413,In_1904,In_444);
or U414 (N_414,In_624,In_1975);
or U415 (N_415,In_1191,In_78);
and U416 (N_416,In_1806,In_49);
or U417 (N_417,In_1329,In_2085);
and U418 (N_418,In_2825,In_2686);
or U419 (N_419,In_2240,In_1136);
xnor U420 (N_420,In_2986,In_2616);
nor U421 (N_421,In_2655,In_1752);
xnor U422 (N_422,In_676,In_2287);
nor U423 (N_423,In_450,In_861);
nor U424 (N_424,In_2867,In_1923);
xor U425 (N_425,In_2556,In_530);
nor U426 (N_426,In_1438,In_1040);
xor U427 (N_427,In_2828,In_1777);
or U428 (N_428,In_2096,In_2694);
and U429 (N_429,In_924,In_2456);
nand U430 (N_430,In_1911,In_1854);
nand U431 (N_431,In_62,In_2069);
or U432 (N_432,In_1279,In_1162);
nor U433 (N_433,In_1686,In_2283);
and U434 (N_434,In_1922,In_590);
nor U435 (N_435,In_2861,In_380);
or U436 (N_436,In_1227,In_458);
nor U437 (N_437,In_270,In_1641);
nor U438 (N_438,In_1208,In_990);
and U439 (N_439,In_1027,In_1411);
and U440 (N_440,In_520,In_837);
or U441 (N_441,In_636,In_2521);
xor U442 (N_442,In_2875,In_1857);
or U443 (N_443,In_2787,In_2711);
xor U444 (N_444,In_2420,In_2405);
nor U445 (N_445,In_2320,In_528);
or U446 (N_446,In_2558,In_2710);
nor U447 (N_447,In_1767,In_275);
xor U448 (N_448,In_2625,In_2631);
nor U449 (N_449,In_2434,In_2621);
nor U450 (N_450,In_643,In_2554);
and U451 (N_451,In_697,In_2690);
xnor U452 (N_452,In_857,In_1067);
nor U453 (N_453,In_1524,In_1087);
and U454 (N_454,In_1452,In_1125);
nor U455 (N_455,In_1566,In_2376);
and U456 (N_456,In_2319,In_656);
and U457 (N_457,In_1171,In_699);
xor U458 (N_458,In_1002,In_2480);
nor U459 (N_459,In_2206,In_2768);
nand U460 (N_460,In_1766,In_2483);
xor U461 (N_461,In_1824,In_1000);
xnor U462 (N_462,In_2874,In_2727);
nor U463 (N_463,In_1651,In_2578);
nand U464 (N_464,In_2452,In_321);
or U465 (N_465,In_1666,In_8);
xnor U466 (N_466,In_2641,In_580);
nand U467 (N_467,In_1271,In_1892);
or U468 (N_468,In_299,In_359);
and U469 (N_469,In_651,In_1987);
or U470 (N_470,In_2046,In_2990);
nor U471 (N_471,In_2645,In_340);
or U472 (N_472,In_988,In_1594);
xnor U473 (N_473,In_826,In_542);
nor U474 (N_474,In_1541,In_1913);
nand U475 (N_475,In_168,In_2583);
nand U476 (N_476,In_2865,In_881);
nor U477 (N_477,In_653,In_2661);
nand U478 (N_478,In_2786,In_2034);
xnor U479 (N_479,In_1112,In_448);
nand U480 (N_480,In_460,In_1727);
or U481 (N_481,In_750,In_83);
xnor U482 (N_482,In_180,In_576);
and U483 (N_483,In_1354,In_334);
xnor U484 (N_484,In_2506,In_1597);
and U485 (N_485,In_1490,In_1872);
xor U486 (N_486,In_1258,In_1462);
and U487 (N_487,In_455,In_629);
nand U488 (N_488,In_2348,In_1989);
nor U489 (N_489,In_1433,In_731);
nor U490 (N_490,In_1034,In_432);
nor U491 (N_491,In_1209,In_1357);
xnor U492 (N_492,In_2488,In_190);
nand U493 (N_493,In_2925,In_1062);
nor U494 (N_494,In_2044,In_882);
nand U495 (N_495,In_1151,In_1710);
xor U496 (N_496,In_2589,In_1384);
xnor U497 (N_497,In_1528,In_1721);
nor U498 (N_498,In_1637,In_947);
xnor U499 (N_499,In_1420,In_1299);
xnor U500 (N_500,In_2113,In_2790);
xor U501 (N_501,In_958,In_2212);
or U502 (N_502,In_1676,In_2158);
nand U503 (N_503,In_2894,In_849);
nand U504 (N_504,In_374,In_2573);
or U505 (N_505,In_1504,In_1533);
nor U506 (N_506,In_710,In_1751);
nor U507 (N_507,In_2980,In_1984);
and U508 (N_508,In_1372,In_985);
nor U509 (N_509,In_1092,In_757);
nand U510 (N_510,In_498,In_2784);
or U511 (N_511,In_1469,In_192);
xor U512 (N_512,In_1848,In_2244);
and U513 (N_513,In_2833,In_2726);
xnor U514 (N_514,In_2983,In_951);
nor U515 (N_515,In_825,In_2147);
nand U516 (N_516,In_1941,In_1326);
xnor U517 (N_517,In_2676,In_113);
xnor U518 (N_518,In_2279,In_808);
nand U519 (N_519,In_2700,In_2651);
xor U520 (N_520,In_1146,In_2061);
nand U521 (N_521,In_1657,In_907);
and U522 (N_522,In_1636,In_1307);
and U523 (N_523,In_1417,In_794);
and U524 (N_524,In_1016,In_2469);
nand U525 (N_525,In_1013,In_2973);
xor U526 (N_526,In_2427,In_2792);
or U527 (N_527,In_2109,In_2810);
nand U528 (N_528,In_2756,In_231);
nand U529 (N_529,In_1118,In_713);
xnor U530 (N_530,In_2350,In_2293);
nor U531 (N_531,In_572,In_851);
nor U532 (N_532,In_1635,In_147);
xor U533 (N_533,In_1345,In_707);
xnor U534 (N_534,In_1883,In_2847);
nand U535 (N_535,In_1413,In_2737);
nor U536 (N_536,In_1160,In_481);
and U537 (N_537,In_1645,In_109);
and U538 (N_538,In_790,In_277);
xnor U539 (N_539,In_567,In_2841);
or U540 (N_540,In_784,In_2814);
nor U541 (N_541,In_2418,In_921);
nor U542 (N_542,In_1406,In_2159);
xnor U543 (N_543,In_474,In_760);
nand U544 (N_544,In_1614,In_2738);
or U545 (N_545,In_1639,In_606);
xnor U546 (N_546,In_571,In_72);
xnor U547 (N_547,In_2038,In_1851);
xor U548 (N_548,In_1055,In_2516);
nand U549 (N_549,In_2644,In_1124);
xor U550 (N_550,In_630,In_2129);
nor U551 (N_551,In_991,In_2630);
xnor U552 (N_552,In_1073,In_1836);
and U553 (N_553,In_1835,In_1842);
xnor U554 (N_554,In_1840,In_2551);
nor U555 (N_555,In_2560,In_2548);
or U556 (N_556,In_2715,In_521);
and U557 (N_557,In_997,In_2430);
or U558 (N_558,In_2411,In_1758);
or U559 (N_559,In_2542,In_2981);
xor U560 (N_560,In_2221,In_2301);
nor U561 (N_561,In_1706,In_952);
or U562 (N_562,In_2123,In_846);
nand U563 (N_563,In_371,In_2392);
nor U564 (N_564,In_1838,In_1579);
or U565 (N_565,In_2050,In_2450);
nand U566 (N_566,In_2102,In_2826);
nand U567 (N_567,In_2245,In_1880);
and U568 (N_568,In_1370,In_941);
nand U569 (N_569,In_511,In_552);
nand U570 (N_570,In_1773,In_901);
nor U571 (N_571,In_2089,In_2026);
and U572 (N_572,In_2215,In_1509);
nor U573 (N_573,In_2794,In_307);
nor U574 (N_574,In_171,In_1041);
xor U575 (N_575,In_2599,In_2247);
and U576 (N_576,In_1012,In_852);
or U577 (N_577,In_2989,In_1763);
nand U578 (N_578,In_1596,In_333);
or U579 (N_579,In_158,In_375);
or U580 (N_580,In_1790,In_1014);
nand U581 (N_581,In_780,In_1063);
or U582 (N_582,In_2681,In_223);
nor U583 (N_583,In_264,In_2994);
nand U584 (N_584,In_2457,In_1478);
and U585 (N_585,In_2265,In_2358);
xor U586 (N_586,In_292,In_2746);
nor U587 (N_587,In_1249,In_1578);
nor U588 (N_588,In_1634,In_302);
nand U589 (N_589,In_618,In_1398);
nand U590 (N_590,In_2895,In_60);
xnor U591 (N_591,In_1592,In_503);
xor U592 (N_592,In_864,In_1314);
and U593 (N_593,In_205,In_765);
nand U594 (N_594,In_548,In_2436);
xnor U595 (N_595,In_608,In_412);
or U596 (N_596,In_2242,In_2565);
nor U597 (N_597,In_271,In_1257);
or U598 (N_598,In_850,In_1995);
nor U599 (N_599,In_2125,In_2618);
nand U600 (N_600,In_206,In_2511);
nor U601 (N_601,In_2374,In_502);
and U602 (N_602,In_999,In_2021);
nand U603 (N_603,In_2036,In_2615);
nand U604 (N_604,In_2675,In_885);
or U605 (N_605,In_652,In_268);
nand U606 (N_606,In_2624,In_482);
and U607 (N_607,In_2065,In_1147);
nand U608 (N_608,In_2883,In_50);
and U609 (N_609,In_976,In_84);
nor U610 (N_610,In_2761,In_210);
nand U611 (N_611,In_163,In_1373);
xor U612 (N_612,In_111,In_824);
xor U613 (N_613,In_1068,In_1482);
nor U614 (N_614,In_930,In_1172);
xnor U615 (N_615,In_1315,In_465);
nand U616 (N_616,In_2493,In_893);
xnor U617 (N_617,In_251,In_2666);
nor U618 (N_618,In_603,In_322);
nand U619 (N_619,In_2961,In_904);
or U620 (N_620,In_1678,In_418);
nand U621 (N_621,In_818,In_1729);
or U622 (N_622,In_174,In_1244);
xor U623 (N_623,In_2211,In_2938);
and U624 (N_624,In_1971,In_1267);
nor U625 (N_625,In_795,In_2812);
or U626 (N_626,In_1023,In_582);
nand U627 (N_627,In_838,In_1128);
and U628 (N_628,In_1708,In_364);
and U629 (N_629,In_604,In_1650);
or U630 (N_630,In_1956,In_2257);
nor U631 (N_631,In_922,In_555);
xnor U632 (N_632,In_1506,In_2361);
and U633 (N_633,In_680,In_2626);
or U634 (N_634,In_1895,In_1456);
nand U635 (N_635,In_955,In_2671);
or U636 (N_636,In_1116,In_36);
nor U637 (N_637,In_303,In_2952);
xnor U638 (N_638,In_1731,In_1311);
and U639 (N_639,In_626,In_2856);
nand U640 (N_640,In_1633,In_1405);
and U641 (N_641,In_1365,In_1695);
and U642 (N_642,In_889,In_2944);
xnor U643 (N_643,In_125,In_1740);
nor U644 (N_644,In_890,In_1133);
and U645 (N_645,In_2132,In_1546);
and U646 (N_646,In_2907,In_2491);
xnor U647 (N_647,In_2668,In_1202);
and U648 (N_648,In_1351,In_1337);
xor U649 (N_649,In_942,In_724);
nand U650 (N_650,In_533,In_1192);
and U651 (N_651,In_2764,In_1612);
nor U652 (N_652,In_2512,In_2003);
xor U653 (N_653,In_2742,In_768);
xor U654 (N_654,In_385,In_456);
or U655 (N_655,In_97,In_2054);
nand U656 (N_656,In_1775,In_87);
xnor U657 (N_657,In_1800,In_2698);
and U658 (N_658,In_715,In_654);
nand U659 (N_659,In_1038,In_1467);
xor U660 (N_660,In_801,In_201);
and U661 (N_661,In_2723,In_1630);
and U662 (N_662,In_1347,In_819);
xnor U663 (N_663,In_88,In_2568);
nand U664 (N_664,In_2571,In_2303);
nand U665 (N_665,In_310,In_1049);
or U666 (N_666,In_2920,In_2771);
nor U667 (N_667,In_2688,In_2344);
or U668 (N_668,In_1245,In_879);
or U669 (N_669,In_1409,In_1425);
nand U670 (N_670,In_1107,In_1701);
or U671 (N_671,In_1134,In_2646);
nand U672 (N_672,In_1089,In_2824);
nor U673 (N_673,In_1086,In_525);
xor U674 (N_674,In_1974,In_2140);
xor U675 (N_675,In_2292,In_354);
or U676 (N_676,In_276,In_1771);
or U677 (N_677,In_925,In_2357);
and U678 (N_678,In_599,In_612);
nor U679 (N_679,In_2862,In_500);
xor U680 (N_680,In_2278,In_159);
and U681 (N_681,In_2210,In_1966);
nand U682 (N_682,In_2775,In_685);
and U683 (N_683,In_2183,In_1470);
xnor U684 (N_684,In_1156,In_506);
or U685 (N_685,In_1621,In_428);
xnor U686 (N_686,In_518,In_2432);
nor U687 (N_687,In_162,In_646);
nand U688 (N_688,In_464,In_1620);
nor U689 (N_689,In_2182,In_1972);
or U690 (N_690,In_1455,In_1899);
or U691 (N_691,In_2162,In_295);
xnor U692 (N_692,In_686,In_2000);
or U693 (N_693,In_1749,In_2014);
and U694 (N_694,In_1748,In_2758);
or U695 (N_695,In_591,In_758);
nor U696 (N_696,In_117,In_1230);
xnor U697 (N_697,In_2375,In_1132);
nor U698 (N_698,In_2360,In_2002);
or U699 (N_699,In_1047,In_538);
or U700 (N_700,In_304,In_2890);
nor U701 (N_701,In_1698,In_1796);
xnor U702 (N_702,In_1648,In_145);
nor U703 (N_703,In_1744,In_1672);
and U704 (N_704,In_1765,In_2249);
nor U705 (N_705,In_1554,In_2254);
nand U706 (N_706,In_800,In_1761);
and U707 (N_707,In_2629,In_1556);
or U708 (N_708,In_1565,In_1946);
nor U709 (N_709,In_1694,In_2446);
and U710 (N_710,In_1225,In_20);
xnor U711 (N_711,In_2722,In_2264);
nand U712 (N_712,In_2712,In_704);
or U713 (N_713,In_152,In_360);
or U714 (N_714,In_2705,In_2335);
and U715 (N_715,In_683,In_1526);
and U716 (N_716,In_256,In_625);
xnor U717 (N_717,In_2068,In_1489);
or U718 (N_718,In_2721,In_536);
or U719 (N_719,In_1760,In_2364);
xor U720 (N_720,In_177,In_2860);
nand U721 (N_721,In_363,In_1900);
or U722 (N_722,In_1811,In_1117);
nor U723 (N_723,In_2217,In_462);
nand U724 (N_724,In_1222,In_2739);
nand U725 (N_725,In_2345,In_740);
xnor U726 (N_726,In_2006,In_2932);
or U727 (N_727,In_18,In_2793);
xor U728 (N_728,In_1426,In_1096);
nand U729 (N_729,In_1703,In_1403);
nor U730 (N_730,In_1909,In_2950);
and U731 (N_731,In_1497,In_329);
or U732 (N_732,In_82,In_220);
nand U733 (N_733,In_1862,In_1350);
nand U734 (N_734,In_1264,In_2074);
nand U735 (N_735,In_742,In_2492);
nor U736 (N_736,In_1772,In_2151);
or U737 (N_737,In_1876,In_2839);
or U738 (N_738,In_2593,In_841);
nand U739 (N_739,In_1397,In_1363);
and U740 (N_740,In_1822,In_1229);
nor U741 (N_741,In_917,In_2332);
or U742 (N_742,In_1536,In_2300);
nand U743 (N_743,In_1535,In_1053);
and U744 (N_744,In_913,In_47);
xor U745 (N_745,In_339,In_2968);
and U746 (N_746,In_1781,In_1599);
nand U747 (N_747,In_2976,In_973);
or U748 (N_748,In_1757,In_978);
and U749 (N_749,In_2233,In_2083);
nand U750 (N_750,In_2266,In_720);
xnor U751 (N_751,In_2127,In_2763);
xor U752 (N_752,In_927,In_2719);
xor U753 (N_753,In_1100,In_1618);
xor U754 (N_754,In_421,In_2197);
xnor U755 (N_755,In_323,In_687);
nand U756 (N_756,In_2628,In_2087);
or U757 (N_757,In_1054,In_2996);
and U758 (N_758,In_670,In_1736);
or U759 (N_759,In_2378,In_2482);
nand U760 (N_760,In_2612,In_534);
xnor U761 (N_761,In_2437,In_746);
nand U762 (N_762,In_2509,In_2032);
nand U763 (N_763,In_706,In_1436);
xnor U764 (N_764,In_2582,In_2194);
xor U765 (N_765,In_716,In_2702);
and U766 (N_766,In_2273,In_1430);
and U767 (N_767,In_2101,In_1877);
xnor U768 (N_768,In_449,In_64);
and U769 (N_769,In_1241,In_2978);
nor U770 (N_770,In_1865,In_1137);
xor U771 (N_771,In_22,In_2130);
xor U772 (N_772,In_888,In_2796);
and U773 (N_773,In_265,In_274);
and U774 (N_774,In_2687,In_2015);
and U775 (N_775,In_2759,In_1213);
and U776 (N_776,In_1270,In_1498);
or U777 (N_777,In_2470,In_948);
nand U778 (N_778,In_2930,In_2782);
nor U779 (N_779,In_1212,In_915);
and U780 (N_780,In_642,In_1802);
nand U781 (N_781,In_2352,In_1609);
nor U782 (N_782,In_2766,In_200);
nand U783 (N_783,In_232,In_2334);
nor U784 (N_784,In_445,In_1794);
xnor U785 (N_785,In_2997,In_2966);
nand U786 (N_786,In_532,In_1884);
nand U787 (N_787,In_960,In_1021);
xor U788 (N_788,In_1182,In_856);
nor U789 (N_789,In_967,In_1962);
or U790 (N_790,In_1091,In_1673);
or U791 (N_791,In_484,In_859);
nor U792 (N_792,In_2979,In_1167);
nand U793 (N_793,In_2042,In_2406);
or U794 (N_794,In_610,In_1600);
or U795 (N_795,In_1891,In_1095);
nand U796 (N_796,In_830,In_92);
nand U797 (N_797,In_797,In_415);
nor U798 (N_798,In_1020,In_1157);
xnor U799 (N_799,In_1224,In_1272);
xnor U800 (N_800,In_187,In_1944);
xnor U801 (N_801,In_865,In_2161);
and U802 (N_802,In_2382,In_1930);
or U803 (N_803,In_2528,In_2179);
and U804 (N_804,In_246,In_2880);
or U805 (N_805,In_2263,In_2588);
nand U806 (N_806,In_2078,In_1078);
and U807 (N_807,In_1366,In_2802);
xor U808 (N_808,In_1295,In_898);
xor U809 (N_809,In_2199,In_906);
nor U810 (N_810,In_2185,In_804);
nand U811 (N_811,In_2704,In_477);
or U812 (N_812,In_1103,In_1934);
nand U813 (N_813,In_2148,In_2853);
xnor U814 (N_814,In_2740,In_2377);
nand U815 (N_815,In_2822,In_1471);
nand U816 (N_816,In_2461,In_2945);
and U817 (N_817,In_693,In_2580);
or U818 (N_818,In_554,In_979);
or U819 (N_819,In_357,In_747);
and U820 (N_820,In_1024,In_739);
xor U821 (N_821,In_665,In_1860);
nor U822 (N_822,In_1647,In_294);
nand U823 (N_823,In_2872,In_2801);
and U824 (N_824,In_493,In_293);
nor U825 (N_825,In_2877,In_2540);
nor U826 (N_826,In_2214,In_475);
nand U827 (N_827,In_547,In_2696);
nor U828 (N_828,In_1795,In_1628);
or U829 (N_829,In_1714,In_565);
nor U830 (N_830,In_641,In_2933);
and U831 (N_831,In_2386,In_1464);
nor U832 (N_832,In_2851,In_1341);
or U833 (N_833,In_688,In_247);
nor U834 (N_834,In_7,In_2444);
and U835 (N_835,In_2765,In_2575);
xor U836 (N_836,In_1321,In_634);
nand U837 (N_837,In_1175,In_1149);
or U838 (N_838,In_2817,In_2341);
nor U839 (N_839,In_517,In_2597);
nand U840 (N_840,In_207,In_619);
and U841 (N_841,In_2018,In_1950);
xnor U842 (N_842,In_1990,In_214);
xor U843 (N_843,In_347,In_884);
and U844 (N_844,In_764,In_1723);
or U845 (N_845,In_692,In_2753);
xnor U846 (N_846,In_269,In_2146);
or U847 (N_847,In_1570,In_2270);
or U848 (N_848,In_420,In_1640);
or U849 (N_849,In_2581,In_1320);
nand U850 (N_850,In_272,In_1742);
nand U851 (N_851,In_2520,In_919);
xor U852 (N_852,In_182,In_578);
nand U853 (N_853,In_422,In_2951);
and U854 (N_854,In_944,In_2889);
xnor U855 (N_855,In_1520,In_226);
or U856 (N_856,In_2016,In_1123);
nor U857 (N_857,In_1377,In_1481);
xnor U858 (N_858,In_1688,In_37);
nor U859 (N_859,In_1205,In_2281);
nand U860 (N_860,In_110,In_2898);
or U861 (N_861,In_24,In_1206);
nor U862 (N_862,In_2549,In_204);
and U863 (N_863,In_1262,In_1896);
nor U864 (N_864,In_2010,In_1910);
xnor U865 (N_865,In_2440,In_1450);
nor U866 (N_866,In_1954,In_598);
and U867 (N_867,In_1890,In_1529);
or U868 (N_868,In_2172,In_12);
nor U869 (N_869,In_811,In_1908);
nand U870 (N_870,In_914,In_1831);
nor U871 (N_871,In_807,In_1998);
and U872 (N_872,In_0,In_2305);
nor U873 (N_873,In_492,In_234);
nand U874 (N_874,In_2909,In_2180);
xor U875 (N_875,In_1575,In_1627);
xnor U876 (N_876,In_2404,In_2912);
or U877 (N_877,In_2884,In_254);
or U878 (N_878,In_1454,In_752);
xor U879 (N_879,In_1873,In_863);
xnor U880 (N_880,In_2489,In_1809);
nor U881 (N_881,In_1743,In_2916);
xor U882 (N_882,In_1474,In_2058);
nand U883 (N_883,In_2439,In_2815);
xnor U884 (N_884,In_2937,In_663);
and U885 (N_885,In_566,In_2138);
or U886 (N_886,In_1273,In_263);
nand U887 (N_887,In_356,In_13);
xnor U888 (N_888,In_1309,In_5);
or U889 (N_889,In_2362,In_2647);
and U890 (N_890,In_2041,In_694);
and U891 (N_891,In_2045,In_2590);
xor U892 (N_892,In_1577,In_21);
and U893 (N_893,In_381,In_2605);
and U894 (N_894,In_2460,In_2529);
nand U895 (N_895,In_33,In_2798);
nand U896 (N_896,In_10,In_593);
nand U897 (N_897,In_397,In_243);
nand U898 (N_898,In_165,In_2379);
xor U899 (N_899,In_2455,In_1728);
nor U900 (N_900,In_717,In_414);
nand U901 (N_901,In_2208,In_621);
xnor U902 (N_902,In_1545,In_80);
xor U903 (N_903,In_153,In_410);
or U904 (N_904,In_2286,In_883);
or U905 (N_905,In_1088,In_2235);
xor U906 (N_906,In_378,In_2977);
xnor U907 (N_907,In_1667,In_892);
nor U908 (N_908,In_379,In_1492);
and U909 (N_909,In_1358,In_1702);
or U910 (N_910,In_1032,In_306);
nand U911 (N_911,In_497,In_2385);
and U912 (N_912,In_297,In_1415);
nor U913 (N_913,In_2004,In_2413);
or U914 (N_914,In_1791,In_627);
xor U915 (N_915,In_1662,In_315);
or U916 (N_916,In_1186,In_649);
nand U917 (N_917,In_85,In_2395);
nor U918 (N_918,In_2594,In_1083);
and U919 (N_919,In_1082,In_931);
nand U920 (N_920,In_789,In_2547);
or U921 (N_921,In_2964,In_1391);
nand U922 (N_922,In_2987,In_1138);
nand U923 (N_923,In_1109,In_1009);
xor U924 (N_924,In_1308,In_42);
nor U925 (N_925,In_1967,In_141);
and U926 (N_926,In_1297,In_2317);
xnor U927 (N_927,In_2472,In_2693);
and U928 (N_928,In_1902,In_2190);
or U929 (N_929,In_975,In_395);
xor U930 (N_930,In_386,In_454);
nor U931 (N_931,In_2390,In_788);
xnor U932 (N_932,In_289,In_791);
nand U933 (N_933,In_1834,In_431);
xnor U934 (N_934,In_136,In_2673);
xnor U935 (N_935,In_108,In_723);
nor U936 (N_936,In_2703,In_2750);
or U937 (N_937,In_1453,In_510);
and U938 (N_938,In_2510,In_2473);
nor U939 (N_939,In_1632,In_806);
nand U940 (N_940,In_2900,In_1379);
nor U941 (N_941,In_1290,In_2842);
and U942 (N_942,In_834,In_1445);
and U943 (N_943,In_595,In_1217);
xor U944 (N_944,In_459,In_1626);
nand U945 (N_945,In_2557,In_2855);
and U946 (N_946,In_89,In_1522);
nor U947 (N_947,In_2871,In_2999);
nand U948 (N_948,In_469,In_1724);
and U949 (N_949,In_346,In_405);
xor U950 (N_950,In_581,In_55);
or U951 (N_951,In_770,In_774);
or U952 (N_952,In_164,In_946);
xnor U953 (N_953,In_1385,In_2677);
and U954 (N_954,In_1356,In_138);
nor U955 (N_955,In_2302,In_361);
or U956 (N_956,In_2067,In_2072);
nand U957 (N_957,In_2834,In_2426);
nand U958 (N_958,In_2947,In_65);
xnor U959 (N_959,In_1830,In_1926);
nand U960 (N_960,In_124,In_471);
nor U961 (N_961,In_1530,In_1973);
nand U962 (N_962,In_1881,In_559);
nor U963 (N_963,In_2774,In_1001);
nor U964 (N_964,In_2486,In_2620);
nand U965 (N_965,In_840,In_2209);
or U966 (N_966,In_2371,In_1875);
nor U967 (N_967,In_1816,In_809);
or U968 (N_968,In_1861,In_181);
xor U969 (N_969,In_2804,In_424);
xor U970 (N_970,In_1458,In_2107);
and U971 (N_971,In_86,In_2899);
and U972 (N_972,In_391,In_1817);
nor U973 (N_973,In_230,In_645);
or U974 (N_974,In_27,In_1434);
nor U975 (N_975,In_383,In_786);
and U976 (N_976,In_667,In_2248);
nor U977 (N_977,In_362,In_2893);
nor U978 (N_978,In_1242,In_2166);
nor U979 (N_979,In_2953,In_661);
or U980 (N_980,In_1879,In_1281);
xor U981 (N_981,In_2328,In_1148);
and U982 (N_982,In_1339,In_2027);
and U983 (N_983,In_427,In_366);
nand U984 (N_984,In_1142,In_701);
or U985 (N_985,In_868,In_541);
xor U986 (N_986,In_537,In_1915);
nor U987 (N_987,In_308,In_1659);
xnor U988 (N_988,In_238,In_1446);
or U989 (N_989,In_1722,In_526);
nor U990 (N_990,In_1343,In_2733);
nand U991 (N_991,In_2370,In_406);
or U992 (N_992,In_2892,In_2398);
xor U993 (N_993,In_1718,In_858);
nor U994 (N_994,In_2174,In_1887);
or U995 (N_995,In_735,In_821);
and U996 (N_996,In_615,In_1932);
xor U997 (N_997,In_250,In_1376);
and U998 (N_998,In_1364,In_1203);
xor U999 (N_999,In_193,In_1983);
xor U1000 (N_1000,In_2415,In_1228);
or U1001 (N_1001,In_2165,In_2075);
xor U1002 (N_1002,In_509,In_1197);
xor U1003 (N_1003,In_916,In_353);
and U1004 (N_1004,In_2507,In_2323);
nor U1005 (N_1005,In_1844,In_1144);
or U1006 (N_1006,In_313,In_2117);
and U1007 (N_1007,In_225,In_2246);
or U1008 (N_1008,In_816,In_1521);
and U1009 (N_1009,In_2827,In_1542);
xnor U1010 (N_1010,In_1010,In_2136);
and U1011 (N_1011,In_798,In_1404);
xor U1012 (N_1012,In_348,In_775);
and U1013 (N_1013,In_2820,In_1077);
nor U1014 (N_1014,In_126,In_1259);
or U1015 (N_1015,In_684,In_2354);
or U1016 (N_1016,In_2366,In_237);
nand U1017 (N_1017,In_54,In_872);
nor U1018 (N_1018,In_2,In_1283);
nand U1019 (N_1019,In_1303,In_1140);
or U1020 (N_1020,In_1812,In_1296);
nand U1021 (N_1021,In_1745,In_1316);
nor U1022 (N_1022,In_419,In_25);
or U1023 (N_1023,In_282,In_2674);
and U1024 (N_1024,In_1340,In_2267);
nand U1025 (N_1025,In_2701,In_964);
and U1026 (N_1026,In_1709,In_773);
or U1027 (N_1027,In_1945,In_1552);
xor U1028 (N_1028,In_2667,In_957);
and U1029 (N_1029,In_1993,In_1419);
nor U1030 (N_1030,In_1553,In_2613);
nor U1031 (N_1031,In_1755,In_127);
xnor U1032 (N_1032,In_156,In_1026);
nor U1033 (N_1033,In_933,In_980);
xor U1034 (N_1034,In_1459,In_2325);
xnor U1035 (N_1035,In_2805,In_41);
xor U1036 (N_1036,In_2514,In_512);
xor U1037 (N_1037,In_544,In_1282);
nor U1038 (N_1038,In_1483,In_2186);
or U1039 (N_1039,In_779,In_211);
xnor U1040 (N_1040,In_1302,In_867);
nand U1041 (N_1041,In_833,In_748);
or U1042 (N_1042,In_1540,In_2799);
or U1043 (N_1043,In_151,In_2584);
xor U1044 (N_1044,In_655,In_753);
nand U1045 (N_1045,In_1561,In_409);
nand U1046 (N_1046,In_671,In_1253);
or U1047 (N_1047,In_2956,In_1705);
nand U1048 (N_1048,In_560,In_2918);
nand U1049 (N_1049,In_1221,In_1051);
nand U1050 (N_1050,In_2531,In_929);
xor U1051 (N_1051,In_1958,In_2121);
or U1052 (N_1052,In_1401,In_2308);
and U1053 (N_1053,In_1048,In_67);
nand U1054 (N_1054,In_1382,In_222);
and U1055 (N_1055,In_529,In_74);
nor U1056 (N_1056,In_1275,In_622);
and U1057 (N_1057,In_233,In_1216);
nor U1058 (N_1058,In_2936,In_839);
xnor U1059 (N_1059,In_782,In_674);
or U1060 (N_1060,In_1052,In_2098);
xnor U1061 (N_1061,In_1846,In_2970);
and U1062 (N_1062,In_783,In_2447);
nand U1063 (N_1063,In_103,In_291);
nand U1064 (N_1064,In_1044,In_1084);
nand U1065 (N_1065,In_491,In_2692);
nor U1066 (N_1066,In_1210,In_2181);
and U1067 (N_1067,In_2538,In_1741);
xnor U1068 (N_1068,In_2891,In_2795);
or U1069 (N_1069,In_787,In_93);
nor U1070 (N_1070,In_2926,In_2094);
nor U1071 (N_1071,In_1965,In_98);
and U1072 (N_1072,In_1737,In_2992);
and U1073 (N_1073,In_803,In_664);
or U1074 (N_1074,In_2633,In_2585);
nand U1075 (N_1075,In_1381,In_2407);
nor U1076 (N_1076,In_2007,In_2490);
xnor U1077 (N_1077,In_2781,In_2466);
nand U1078 (N_1078,In_2522,In_281);
nor U1079 (N_1079,In_2837,In_1294);
or U1080 (N_1080,In_2903,In_1289);
and U1081 (N_1081,In_319,In_2474);
xnor U1082 (N_1082,In_2717,In_1265);
or U1083 (N_1083,In_2569,In_2276);
or U1084 (N_1084,In_285,In_2946);
or U1085 (N_1085,In_1395,In_1856);
nor U1086 (N_1086,In_1584,In_1005);
nand U1087 (N_1087,In_1920,In_1348);
nor U1088 (N_1088,In_1301,In_1978);
nor U1089 (N_1089,In_2187,In_188);
nor U1090 (N_1090,In_2178,In_2167);
nand U1091 (N_1091,In_2222,In_2610);
xor U1092 (N_1092,In_1075,In_1948);
or U1093 (N_1093,In_2081,In_2770);
and U1094 (N_1094,In_1185,In_1919);
nand U1095 (N_1095,In_398,In_2141);
and U1096 (N_1096,In_115,In_2306);
xor U1097 (N_1097,In_628,In_1400);
nand U1098 (N_1098,In_1181,In_2262);
or U1099 (N_1099,In_1595,In_2024);
xnor U1100 (N_1100,In_2258,In_129);
nor U1101 (N_1101,In_40,In_273);
and U1102 (N_1102,In_495,In_191);
or U1103 (N_1103,In_1544,In_1003);
nand U1104 (N_1104,In_2988,In_994);
xor U1105 (N_1105,In_620,In_2928);
or U1106 (N_1106,In_776,In_2227);
xor U1107 (N_1107,In_2116,In_1362);
nand U1108 (N_1108,In_2902,In_1421);
or U1109 (N_1109,In_935,In_1935);
nor U1110 (N_1110,In_820,In_1574);
or U1111 (N_1111,In_2327,In_1056);
nand U1112 (N_1112,In_2639,In_2484);
and U1113 (N_1113,In_2752,In_1704);
nor U1114 (N_1114,In_2205,In_2023);
nor U1115 (N_1115,In_1774,In_1853);
and U1116 (N_1116,In_2005,In_1399);
xnor U1117 (N_1117,In_499,In_691);
nand U1118 (N_1118,In_584,In_1378);
or U1119 (N_1119,In_1589,In_738);
or U1120 (N_1120,In_2204,In_802);
xnor U1121 (N_1121,In_31,In_1921);
xor U1122 (N_1122,In_2231,In_1925);
or U1123 (N_1123,In_195,In_644);
nor U1124 (N_1124,In_480,In_95);
nor U1125 (N_1125,In_2202,In_452);
or U1126 (N_1126,In_1286,In_2022);
nor U1127 (N_1127,In_1778,In_2924);
nor U1128 (N_1128,In_719,In_2606);
and U1129 (N_1129,In_1670,In_2515);
nand U1130 (N_1130,In_189,In_2562);
nand U1131 (N_1131,In_2274,In_926);
xnor U1132 (N_1132,In_648,In_90);
or U1133 (N_1133,In_118,In_1269);
and U1134 (N_1134,In_1970,In_2849);
and U1135 (N_1135,In_1170,In_1255);
and U1136 (N_1136,In_2780,In_577);
nor U1137 (N_1137,In_2954,In_2751);
and U1138 (N_1138,In_1207,In_1534);
or U1139 (N_1139,In_1007,In_1538);
nor U1140 (N_1140,In_2250,In_443);
xor U1141 (N_1141,In_1488,In_9);
or U1142 (N_1142,In_2080,In_19);
nor U1143 (N_1143,In_1424,In_2806);
nor U1144 (N_1144,In_2336,In_1263);
nor U1145 (N_1145,In_199,In_23);
xnor U1146 (N_1146,In_2713,In_2097);
or U1147 (N_1147,In_771,In_1247);
or U1148 (N_1148,In_52,In_2414);
and U1149 (N_1149,In_1150,In_2134);
and U1150 (N_1150,In_160,In_1085);
and U1151 (N_1151,In_2660,In_1940);
nor U1152 (N_1152,In_2416,In_936);
and U1153 (N_1153,In_540,In_899);
xnor U1154 (N_1154,In_1658,In_433);
nand U1155 (N_1155,In_301,In_2487);
and U1156 (N_1156,In_1665,In_755);
or U1157 (N_1157,In_832,In_416);
nand U1158 (N_1158,In_2419,In_290);
xor U1159 (N_1159,In_262,In_2609);
nor U1160 (N_1160,In_2870,In_2995);
xor U1161 (N_1161,In_1332,In_215);
and U1162 (N_1162,In_714,In_2852);
nor U1163 (N_1163,In_2835,In_2380);
xor U1164 (N_1164,In_1691,In_327);
or U1165 (N_1165,In_2331,In_2284);
xnor U1166 (N_1166,In_631,In_1644);
xnor U1167 (N_1167,In_377,In_1239);
or U1168 (N_1168,In_932,In_2033);
or U1169 (N_1169,In_2636,In_550);
nor U1170 (N_1170,In_939,In_2745);
or U1171 (N_1171,In_326,In_1428);
xnor U1172 (N_1172,In_228,In_721);
nor U1173 (N_1173,In_1463,In_2131);
nor U1174 (N_1174,In_965,In_589);
and U1175 (N_1175,In_2982,In_2934);
nand U1176 (N_1176,In_2854,In_1717);
xnor U1177 (N_1177,In_1427,In_2114);
nand U1178 (N_1178,In_1725,In_815);
nor U1179 (N_1179,In_662,In_1493);
nor U1180 (N_1180,In_1548,In_2229);
and U1181 (N_1181,In_737,In_1684);
xor U1182 (N_1182,In_2809,In_59);
and U1183 (N_1183,In_1232,In_2055);
and U1184 (N_1184,In_2617,In_1646);
and U1185 (N_1185,In_1770,In_2271);
nand U1186 (N_1186,In_2152,In_1897);
xnor U1187 (N_1187,In_451,In_658);
nor U1188 (N_1188,In_1660,In_2310);
xor U1189 (N_1189,In_1807,In_1888);
or U1190 (N_1190,In_2807,In_1852);
or U1191 (N_1191,In_411,In_2942);
xor U1192 (N_1192,In_2237,In_2216);
xor U1193 (N_1193,In_2857,In_2963);
nor U1194 (N_1194,In_2311,In_2503);
xor U1195 (N_1195,In_1028,In_2039);
and U1196 (N_1196,In_943,In_2137);
nand U1197 (N_1197,In_2400,In_1199);
nand U1198 (N_1198,In_1870,In_2530);
and U1199 (N_1199,In_57,In_2135);
nand U1200 (N_1200,In_1547,In_1957);
nand U1201 (N_1201,In_2550,In_1780);
xnor U1202 (N_1202,In_1936,In_2298);
nor U1203 (N_1203,In_2329,In_1523);
nand U1204 (N_1204,In_2476,In_1878);
and U1205 (N_1205,In_2402,In_1898);
or U1206 (N_1206,In_961,In_2960);
xnor U1207 (N_1207,In_2169,In_2144);
nor U1208 (N_1208,In_1058,In_1059);
and U1209 (N_1209,In_712,In_2316);
nor U1210 (N_1210,In_1785,In_623);
nor U1211 (N_1211,In_2226,In_1248);
nand U1212 (N_1212,In_2163,In_2048);
nor U1213 (N_1213,In_2154,In_937);
and U1214 (N_1214,In_56,In_300);
xor U1215 (N_1215,In_1131,In_1616);
or U1216 (N_1216,In_123,In_1649);
nand U1217 (N_1217,In_2355,In_2090);
xnor U1218 (N_1218,In_2600,In_2282);
or U1219 (N_1219,In_61,In_659);
nand U1220 (N_1220,In_579,In_1683);
nor U1221 (N_1221,In_2259,In_2917);
or U1222 (N_1222,In_2680,In_1754);
xor U1223 (N_1223,In_1394,In_759);
or U1224 (N_1224,In_767,In_2570);
nand U1225 (N_1225,In_886,In_1375);
and U1226 (N_1226,In_476,In_2518);
or U1227 (N_1227,In_184,In_1555);
xnor U1228 (N_1228,In_1188,In_1955);
nor U1229 (N_1229,In_974,In_1143);
and U1230 (N_1230,In_372,In_1097);
or U1231 (N_1231,In_2959,In_2099);
nand U1232 (N_1232,In_154,In_249);
and U1233 (N_1233,In_1585,In_441);
and U1234 (N_1234,In_2910,In_934);
and U1235 (N_1235,In_2559,In_1582);
and U1236 (N_1236,In_2927,In_2776);
or U1237 (N_1237,In_2092,In_1153);
xnor U1238 (N_1238,In_799,In_1677);
and U1239 (N_1239,In_1602,In_2718);
or U1240 (N_1240,In_2122,In_1656);
and U1241 (N_1241,In_508,In_722);
nor U1242 (N_1242,In_1671,In_349);
and U1243 (N_1243,In_1697,In_2200);
nand U1244 (N_1244,In_950,In_1065);
or U1245 (N_1245,In_2901,In_666);
nand U1246 (N_1246,In_1251,In_1322);
or U1247 (N_1247,In_2539,In_457);
xor U1248 (N_1248,In_161,In_2603);
or U1249 (N_1249,In_1361,In_102);
xor U1250 (N_1250,In_574,In_1485);
or U1251 (N_1251,In_71,In_314);
and U1252 (N_1252,In_611,In_845);
xnor U1253 (N_1253,In_1033,In_2508);
xnor U1254 (N_1254,In_255,In_28);
nor U1255 (N_1255,In_2967,In_2079);
nor U1256 (N_1256,In_1331,In_2663);
nand U1257 (N_1257,In_2196,In_1105);
and U1258 (N_1258,In_516,In_2485);
nor U1259 (N_1259,In_2555,In_1437);
and U1260 (N_1260,In_1735,In_1484);
and U1261 (N_1261,In_1129,In_698);
nor U1262 (N_1262,In_2685,In_1511);
nor U1263 (N_1263,In_1360,In_2296);
or U1264 (N_1264,In_1996,In_769);
xnor U1265 (N_1265,In_485,In_728);
or U1266 (N_1266,In_785,In_245);
xnor U1267 (N_1267,In_2052,In_2243);
nor U1268 (N_1268,In_1894,In_2965);
and U1269 (N_1269,In_1183,In_561);
nand U1270 (N_1270,In_1223,In_1798);
or U1271 (N_1271,In_1046,In_248);
or U1272 (N_1272,In_1368,In_1501);
nor U1273 (N_1273,In_2602,In_2315);
and U1274 (N_1274,In_2241,In_122);
and U1275 (N_1275,In_466,In_1298);
xor U1276 (N_1276,In_1768,In_75);
xnor U1277 (N_1277,In_897,In_1539);
nand U1278 (N_1278,In_2339,In_53);
and U1279 (N_1279,In_2844,In_660);
nand U1280 (N_1280,In_1580,In_324);
xor U1281 (N_1281,In_94,In_1278);
nand U1282 (N_1282,In_605,In_166);
and U1283 (N_1283,In_616,In_131);
nor U1284 (N_1284,In_2777,In_1693);
xnor U1285 (N_1285,In_2649,In_1629);
nand U1286 (N_1286,In_1858,In_1465);
nor U1287 (N_1287,In_1392,In_633);
or U1288 (N_1288,In_17,In_351);
xor U1289 (N_1289,In_1287,In_2232);
nor U1290 (N_1290,In_120,In_488);
nor U1291 (N_1291,In_2040,In_2669);
or U1292 (N_1292,In_2709,In_1177);
and U1293 (N_1293,In_179,In_813);
nand U1294 (N_1294,In_1201,In_700);
or U1295 (N_1295,In_369,In_1947);
nor U1296 (N_1296,In_1163,In_535);
nand U1297 (N_1297,In_2846,In_1961);
nand U1298 (N_1298,In_983,In_1518);
nand U1299 (N_1299,In_1072,In_2762);
or U1300 (N_1300,In_2697,In_696);
nand U1301 (N_1301,In_2545,In_63);
or U1302 (N_1302,In_2253,In_2066);
or U1303 (N_1303,In_76,In_866);
and U1304 (N_1304,In_1992,In_343);
xnor U1305 (N_1305,In_1886,In_373);
or U1306 (N_1306,In_1604,In_2176);
nor U1307 (N_1307,In_176,In_1608);
and U1308 (N_1308,In_772,In_1943);
xnor U1309 (N_1309,In_1110,In_2921);
and U1310 (N_1310,In_1826,In_938);
or U1311 (N_1311,In_1789,In_352);
nor U1312 (N_1312,In_1586,In_1963);
nand U1313 (N_1313,In_527,In_1099);
xnor U1314 (N_1314,In_2213,In_2156);
xor U1315 (N_1315,In_336,In_2438);
or U1316 (N_1316,In_586,In_1173);
or U1317 (N_1317,In_2356,In_912);
and U1318 (N_1318,In_2638,In_2665);
and U1319 (N_1319,In_2498,In_183);
and U1320 (N_1320,In_2164,In_2285);
xor U1321 (N_1321,In_2330,In_101);
nand U1322 (N_1322,In_602,In_367);
xor U1323 (N_1323,In_732,In_2108);
and U1324 (N_1324,In_1942,In_2017);
xor U1325 (N_1325,In_447,In_600);
xor U1326 (N_1326,In_1619,In_66);
nand U1327 (N_1327,In_822,In_2577);
xor U1328 (N_1328,In_1655,In_814);
nand U1329 (N_1329,In_399,In_669);
xnor U1330 (N_1330,In_2653,In_144);
nand U1331 (N_1331,In_2637,In_2789);
or U1332 (N_1332,In_2608,In_1652);
xnor U1333 (N_1333,In_1064,In_2627);
and U1334 (N_1334,In_155,In_1008);
and U1335 (N_1335,In_2873,In_524);
and U1336 (N_1336,In_1080,In_1135);
or U1337 (N_1337,In_1551,In_2056);
or U1338 (N_1338,In_1849,In_1531);
nor U1339 (N_1339,In_1119,In_1480);
nand U1340 (N_1340,In_2897,In_1711);
nor U1341 (N_1341,In_2769,In_853);
nor U1342 (N_1342,In_1845,In_1814);
nor U1343 (N_1343,In_1885,In_2818);
xor U1344 (N_1344,In_1837,In_2670);
xnor U1345 (N_1345,In_1166,In_2479);
xor U1346 (N_1346,In_2314,In_358);
nand U1347 (N_1347,In_895,In_2465);
nand U1348 (N_1348,In_2595,In_1631);
xnor U1349 (N_1349,In_1108,In_2184);
or U1350 (N_1350,In_1231,In_2463);
xnor U1351 (N_1351,In_2399,In_966);
and U1352 (N_1352,In_2561,In_2684);
nand U1353 (N_1353,In_1558,In_1431);
and U1354 (N_1354,In_2915,In_1407);
nand U1355 (N_1355,In_2553,In_435);
nand U1356 (N_1356,In_1019,In_587);
and U1357 (N_1357,In_2297,In_1874);
or U1358 (N_1358,In_1443,In_1726);
nor U1359 (N_1359,In_1690,In_2369);
xnor U1360 (N_1360,In_341,In_1869);
nor U1361 (N_1361,In_2110,In_212);
nand U1362 (N_1362,In_1764,In_763);
and U1363 (N_1363,In_1402,In_390);
nor U1364 (N_1364,In_2149,In_2783);
nor U1365 (N_1365,In_650,In_1680);
and U1366 (N_1366,In_668,In_442);
xnor U1367 (N_1367,In_969,In_569);
xor U1368 (N_1368,In_681,In_2840);
xnor U1369 (N_1369,In_2991,In_1969);
nor U1370 (N_1370,In_2313,In_1598);
nand U1371 (N_1371,In_756,In_2077);
nand U1372 (N_1372,In_2576,In_1111);
nor U1373 (N_1373,In_2009,In_1220);
and U1374 (N_1374,In_2725,In_1820);
or U1375 (N_1375,In_1355,In_2906);
xnor U1376 (N_1376,In_2403,In_2689);
xor U1377 (N_1377,In_613,In_487);
xor U1378 (N_1378,In_4,In_1669);
nand U1379 (N_1379,In_597,In_1102);
nor U1380 (N_1380,In_2343,In_1613);
or U1381 (N_1381,In_1079,In_2365);
nor U1382 (N_1382,In_1720,In_2454);
or U1383 (N_1383,In_478,In_2261);
or U1384 (N_1384,In_1374,In_1423);
xnor U1385 (N_1385,In_810,In_2504);
nand U1386 (N_1386,In_2175,In_1036);
nor U1387 (N_1387,In_553,In_2859);
nor U1388 (N_1388,In_197,In_1988);
or U1389 (N_1389,In_2878,In_148);
nand U1390 (N_1390,In_1479,In_2381);
xor U1391 (N_1391,In_878,In_2188);
or U1392 (N_1392,In_1288,In_137);
nor U1393 (N_1393,In_330,In_2139);
nand U1394 (N_1394,In_157,In_241);
nand U1395 (N_1395,In_1159,In_2168);
or U1396 (N_1396,In_2047,In_543);
nand U1397 (N_1397,In_1093,In_1601);
or U1398 (N_1398,In_298,In_2724);
or U1399 (N_1399,In_2502,In_909);
or U1400 (N_1400,In_370,In_6);
nor U1401 (N_1401,In_48,In_169);
nand U1402 (N_1402,In_368,In_355);
and U1403 (N_1403,In_1617,In_1304);
or U1404 (N_1404,In_2059,In_68);
xor U1405 (N_1405,In_1324,In_2876);
xor U1406 (N_1406,In_1293,In_2699);
nor U1407 (N_1407,In_1184,In_1330);
or U1408 (N_1408,In_2120,In_1449);
and U1409 (N_1409,In_130,In_1161);
or U1410 (N_1410,In_392,In_2534);
nor U1411 (N_1411,In_216,In_2749);
xor U1412 (N_1412,In_1387,In_479);
xnor U1413 (N_1413,In_831,In_2333);
nor U1414 (N_1414,In_2326,In_754);
nand U1415 (N_1415,In_2049,In_1284);
and U1416 (N_1416,In_2755,In_835);
xnor U1417 (N_1417,In_2119,In_32);
nand U1418 (N_1418,In_984,In_1687);
or U1419 (N_1419,In_2494,In_564);
and U1420 (N_1420,In_640,In_2757);
xnor U1421 (N_1421,In_2714,In_2772);
nand U1422 (N_1422,In_1516,In_1828);
xor U1423 (N_1423,In_2073,In_1759);
nand U1424 (N_1424,In_1204,In_229);
and U1425 (N_1425,In_2428,In_1313);
nor U1426 (N_1426,In_1889,In_134);
nor U1427 (N_1427,In_1219,In_2816);
xor U1428 (N_1428,In_1250,In_1712);
nand U1429 (N_1429,In_2836,In_335);
nor U1430 (N_1430,In_2368,In_1739);
nand U1431 (N_1431,In_2269,In_407);
nor U1432 (N_1432,In_2754,In_1367);
nor U1433 (N_1433,In_1235,In_1292);
or U1434 (N_1434,In_672,In_1408);
or U1435 (N_1435,In_2591,In_2408);
and U1436 (N_1436,In_2879,In_2672);
or U1437 (N_1437,In_1903,In_43);
and U1438 (N_1438,In_2011,In_2650);
and U1439 (N_1439,In_1949,In_2133);
xnor U1440 (N_1440,In_2111,In_312);
xor U1441 (N_1441,In_1746,In_1045);
nand U1442 (N_1442,In_1938,In_953);
xnor U1443 (N_1443,In_2057,In_1043);
or U1444 (N_1444,In_1557,In_100);
nand U1445 (N_1445,In_279,In_1070);
xnor U1446 (N_1446,In_2728,In_1977);
nor U1447 (N_1447,In_920,In_514);
nor U1448 (N_1448,In_1939,In_2832);
nand U1449 (N_1449,In_1388,In_1588);
nand U1450 (N_1450,In_596,In_483);
nand U1451 (N_1451,In_1196,In_2433);
xor U1452 (N_1452,In_58,In_617);
and U1453 (N_1453,In_1810,In_266);
or U1454 (N_1454,In_494,In_2393);
xor U1455 (N_1455,In_132,In_1444);
nor U1456 (N_1456,In_401,In_261);
and U1457 (N_1457,In_1901,In_812);
nor U1458 (N_1458,In_1927,In_305);
nand U1459 (N_1459,In_2904,In_1982);
and U1460 (N_1460,In_1422,In_114);
or U1461 (N_1461,In_1319,In_2351);
nand U1462 (N_1462,In_1716,In_709);
nor U1463 (N_1463,In_1187,In_1098);
nor U1464 (N_1464,In_900,In_1502);
and U1465 (N_1465,In_1447,In_2532);
nand U1466 (N_1466,In_239,In_928);
and U1467 (N_1467,In_1560,In_987);
or U1468 (N_1468,In_2342,In_15);
nand U1469 (N_1469,In_1318,In_2294);
and U1470 (N_1470,In_2911,In_792);
or U1471 (N_1471,In_1386,In_875);
nand U1472 (N_1472,In_2729,In_317);
and U1473 (N_1473,In_2029,In_1663);
and U1474 (N_1474,In_2843,In_387);
or U1475 (N_1475,In_1165,In_2850);
or U1476 (N_1476,In_1832,In_2497);
nand U1477 (N_1477,In_2086,In_2574);
xor U1478 (N_1478,In_384,In_556);
nand U1479 (N_1479,In_632,In_1017);
xnor U1480 (N_1480,In_178,In_959);
nor U1481 (N_1481,In_855,In_2735);
nor U1482 (N_1482,In_1605,In_2881);
and U1483 (N_1483,In_2082,In_283);
or U1484 (N_1484,In_2523,In_2349);
or U1485 (N_1485,In_2829,In_2838);
xnor U1486 (N_1486,In_2914,In_711);
or U1487 (N_1487,In_2654,In_981);
and U1488 (N_1488,In_1104,In_1508);
or U1489 (N_1489,In_501,In_1559);
and U1490 (N_1490,In_2155,In_278);
nor U1491 (N_1491,In_1179,In_2387);
nand U1492 (N_1492,In_1779,In_911);
or U1493 (N_1493,In_1475,In_689);
xnor U1494 (N_1494,In_2051,In_2866);
nand U1495 (N_1495,In_2431,In_1799);
nor U1496 (N_1496,In_1537,In_429);
nand U1497 (N_1497,In_2019,In_1808);
nor U1498 (N_1498,In_1642,In_2760);
nand U1499 (N_1499,In_227,In_1543);
xnor U1500 (N_1500,In_2525,In_302);
or U1501 (N_1501,In_2113,In_652);
nand U1502 (N_1502,In_2470,In_276);
and U1503 (N_1503,In_2188,In_1524);
nand U1504 (N_1504,In_580,In_225);
nand U1505 (N_1505,In_2628,In_2327);
and U1506 (N_1506,In_2316,In_215);
and U1507 (N_1507,In_1260,In_2111);
and U1508 (N_1508,In_2936,In_96);
and U1509 (N_1509,In_721,In_2612);
and U1510 (N_1510,In_149,In_2534);
nor U1511 (N_1511,In_2658,In_2154);
nor U1512 (N_1512,In_392,In_1998);
xnor U1513 (N_1513,In_904,In_1727);
or U1514 (N_1514,In_1733,In_1157);
or U1515 (N_1515,In_2208,In_2312);
xnor U1516 (N_1516,In_1697,In_1786);
nand U1517 (N_1517,In_1814,In_1184);
xnor U1518 (N_1518,In_783,In_2541);
or U1519 (N_1519,In_798,In_1428);
nor U1520 (N_1520,In_2231,In_864);
nor U1521 (N_1521,In_169,In_2602);
nand U1522 (N_1522,In_1147,In_2979);
nand U1523 (N_1523,In_2647,In_102);
xnor U1524 (N_1524,In_2588,In_957);
or U1525 (N_1525,In_2521,In_1011);
nand U1526 (N_1526,In_1547,In_2276);
xor U1527 (N_1527,In_1637,In_716);
xnor U1528 (N_1528,In_196,In_846);
xnor U1529 (N_1529,In_181,In_1251);
nor U1530 (N_1530,In_124,In_1055);
or U1531 (N_1531,In_838,In_2895);
or U1532 (N_1532,In_2903,In_379);
nor U1533 (N_1533,In_151,In_1685);
xor U1534 (N_1534,In_1476,In_1559);
and U1535 (N_1535,In_1160,In_1003);
xnor U1536 (N_1536,In_2218,In_2471);
xnor U1537 (N_1537,In_196,In_1544);
and U1538 (N_1538,In_1773,In_2791);
xor U1539 (N_1539,In_1821,In_773);
or U1540 (N_1540,In_2868,In_532);
xnor U1541 (N_1541,In_1506,In_961);
nand U1542 (N_1542,In_2808,In_296);
xor U1543 (N_1543,In_44,In_1717);
or U1544 (N_1544,In_736,In_828);
and U1545 (N_1545,In_31,In_1868);
nand U1546 (N_1546,In_1758,In_1893);
nor U1547 (N_1547,In_2187,In_2952);
nor U1548 (N_1548,In_2866,In_1257);
and U1549 (N_1549,In_948,In_2365);
xor U1550 (N_1550,In_162,In_2496);
or U1551 (N_1551,In_2806,In_2934);
xor U1552 (N_1552,In_1573,In_1000);
or U1553 (N_1553,In_4,In_2239);
xor U1554 (N_1554,In_186,In_2851);
nor U1555 (N_1555,In_1659,In_725);
or U1556 (N_1556,In_1665,In_1462);
nand U1557 (N_1557,In_2448,In_2563);
xor U1558 (N_1558,In_876,In_1350);
and U1559 (N_1559,In_2544,In_164);
nand U1560 (N_1560,In_2810,In_1066);
xnor U1561 (N_1561,In_465,In_888);
nor U1562 (N_1562,In_2820,In_1532);
xnor U1563 (N_1563,In_1243,In_8);
xor U1564 (N_1564,In_394,In_531);
or U1565 (N_1565,In_1854,In_223);
or U1566 (N_1566,In_340,In_2739);
xnor U1567 (N_1567,In_945,In_1773);
nand U1568 (N_1568,In_2592,In_1760);
xnor U1569 (N_1569,In_1171,In_37);
nand U1570 (N_1570,In_1443,In_2642);
or U1571 (N_1571,In_2561,In_663);
or U1572 (N_1572,In_502,In_828);
nand U1573 (N_1573,In_1689,In_1087);
and U1574 (N_1574,In_1363,In_1085);
nand U1575 (N_1575,In_1808,In_2471);
xor U1576 (N_1576,In_1766,In_870);
and U1577 (N_1577,In_2872,In_1531);
xor U1578 (N_1578,In_11,In_2170);
xnor U1579 (N_1579,In_757,In_652);
nand U1580 (N_1580,In_2627,In_86);
or U1581 (N_1581,In_2977,In_2681);
or U1582 (N_1582,In_1160,In_2465);
xor U1583 (N_1583,In_2652,In_1787);
xor U1584 (N_1584,In_1007,In_279);
nand U1585 (N_1585,In_427,In_2066);
and U1586 (N_1586,In_1201,In_1355);
nor U1587 (N_1587,In_1009,In_758);
nand U1588 (N_1588,In_990,In_230);
and U1589 (N_1589,In_2115,In_385);
or U1590 (N_1590,In_1135,In_2013);
nand U1591 (N_1591,In_2224,In_1949);
nand U1592 (N_1592,In_2162,In_33);
nor U1593 (N_1593,In_417,In_577);
xor U1594 (N_1594,In_576,In_2409);
nand U1595 (N_1595,In_966,In_107);
nand U1596 (N_1596,In_2262,In_225);
and U1597 (N_1597,In_1051,In_2948);
or U1598 (N_1598,In_632,In_404);
and U1599 (N_1599,In_637,In_2532);
xnor U1600 (N_1600,In_1354,In_755);
nor U1601 (N_1601,In_55,In_1726);
xnor U1602 (N_1602,In_2472,In_2548);
xor U1603 (N_1603,In_140,In_99);
xor U1604 (N_1604,In_2183,In_1135);
nor U1605 (N_1605,In_2794,In_2521);
nand U1606 (N_1606,In_1820,In_1172);
or U1607 (N_1607,In_1662,In_2941);
or U1608 (N_1608,In_2887,In_2002);
nor U1609 (N_1609,In_2800,In_2541);
or U1610 (N_1610,In_2667,In_2168);
and U1611 (N_1611,In_2580,In_1993);
xnor U1612 (N_1612,In_2341,In_659);
xor U1613 (N_1613,In_2497,In_2992);
or U1614 (N_1614,In_2202,In_142);
or U1615 (N_1615,In_1877,In_643);
or U1616 (N_1616,In_1434,In_2426);
and U1617 (N_1617,In_1240,In_908);
or U1618 (N_1618,In_892,In_2611);
and U1619 (N_1619,In_2036,In_722);
nand U1620 (N_1620,In_2112,In_2456);
xor U1621 (N_1621,In_1245,In_2093);
nand U1622 (N_1622,In_789,In_2602);
and U1623 (N_1623,In_2252,In_2577);
and U1624 (N_1624,In_1559,In_1319);
or U1625 (N_1625,In_2134,In_2495);
or U1626 (N_1626,In_2123,In_1518);
nand U1627 (N_1627,In_1058,In_454);
or U1628 (N_1628,In_2471,In_860);
xor U1629 (N_1629,In_252,In_874);
nor U1630 (N_1630,In_98,In_2805);
nor U1631 (N_1631,In_803,In_1053);
nand U1632 (N_1632,In_1662,In_1923);
or U1633 (N_1633,In_2431,In_106);
nand U1634 (N_1634,In_14,In_2571);
nand U1635 (N_1635,In_2751,In_1623);
nor U1636 (N_1636,In_660,In_2173);
or U1637 (N_1637,In_1331,In_2274);
and U1638 (N_1638,In_2223,In_157);
xor U1639 (N_1639,In_2008,In_693);
nand U1640 (N_1640,In_1082,In_2436);
nor U1641 (N_1641,In_1656,In_2262);
and U1642 (N_1642,In_1143,In_2571);
and U1643 (N_1643,In_2679,In_2321);
nor U1644 (N_1644,In_1675,In_849);
or U1645 (N_1645,In_529,In_1036);
xor U1646 (N_1646,In_2529,In_294);
and U1647 (N_1647,In_395,In_2761);
and U1648 (N_1648,In_2432,In_1368);
and U1649 (N_1649,In_1912,In_506);
xor U1650 (N_1650,In_360,In_1164);
xnor U1651 (N_1651,In_2434,In_1754);
or U1652 (N_1652,In_446,In_1169);
nor U1653 (N_1653,In_2599,In_1159);
nor U1654 (N_1654,In_2268,In_2633);
xnor U1655 (N_1655,In_1989,In_1441);
or U1656 (N_1656,In_209,In_232);
nand U1657 (N_1657,In_1783,In_2043);
nor U1658 (N_1658,In_2261,In_1050);
or U1659 (N_1659,In_1103,In_586);
xnor U1660 (N_1660,In_2894,In_1709);
nor U1661 (N_1661,In_863,In_2125);
nand U1662 (N_1662,In_1541,In_718);
or U1663 (N_1663,In_2544,In_1225);
nand U1664 (N_1664,In_2379,In_932);
nand U1665 (N_1665,In_1587,In_15);
nand U1666 (N_1666,In_1424,In_1405);
nor U1667 (N_1667,In_1225,In_793);
nor U1668 (N_1668,In_1932,In_2661);
nor U1669 (N_1669,In_848,In_1435);
xnor U1670 (N_1670,In_190,In_2358);
and U1671 (N_1671,In_1823,In_2349);
nor U1672 (N_1672,In_487,In_609);
nor U1673 (N_1673,In_1473,In_2774);
nor U1674 (N_1674,In_2161,In_2565);
nor U1675 (N_1675,In_1624,In_1233);
nand U1676 (N_1676,In_2073,In_638);
xnor U1677 (N_1677,In_1179,In_608);
or U1678 (N_1678,In_1805,In_739);
nand U1679 (N_1679,In_739,In_2124);
or U1680 (N_1680,In_2719,In_1471);
xnor U1681 (N_1681,In_696,In_683);
nor U1682 (N_1682,In_289,In_671);
or U1683 (N_1683,In_1012,In_1676);
nand U1684 (N_1684,In_994,In_1487);
xor U1685 (N_1685,In_1880,In_2363);
nand U1686 (N_1686,In_831,In_1922);
nor U1687 (N_1687,In_1791,In_2004);
or U1688 (N_1688,In_2667,In_2131);
nand U1689 (N_1689,In_2723,In_844);
xor U1690 (N_1690,In_656,In_1060);
nand U1691 (N_1691,In_733,In_1684);
or U1692 (N_1692,In_2786,In_2658);
xor U1693 (N_1693,In_1876,In_839);
or U1694 (N_1694,In_45,In_1028);
nand U1695 (N_1695,In_2347,In_1660);
nand U1696 (N_1696,In_1508,In_2379);
nor U1697 (N_1697,In_1871,In_832);
and U1698 (N_1698,In_1650,In_769);
nor U1699 (N_1699,In_1187,In_1687);
xnor U1700 (N_1700,In_490,In_1886);
and U1701 (N_1701,In_2815,In_739);
xor U1702 (N_1702,In_2958,In_2699);
or U1703 (N_1703,In_125,In_1544);
or U1704 (N_1704,In_712,In_965);
xnor U1705 (N_1705,In_1136,In_2781);
and U1706 (N_1706,In_405,In_2746);
or U1707 (N_1707,In_1476,In_37);
nor U1708 (N_1708,In_1471,In_1241);
nor U1709 (N_1709,In_2014,In_1360);
nor U1710 (N_1710,In_2970,In_1112);
and U1711 (N_1711,In_2659,In_1500);
xnor U1712 (N_1712,In_1405,In_2775);
xor U1713 (N_1713,In_2480,In_853);
and U1714 (N_1714,In_38,In_33);
nand U1715 (N_1715,In_2539,In_2009);
nor U1716 (N_1716,In_1695,In_1269);
or U1717 (N_1717,In_2853,In_1400);
nand U1718 (N_1718,In_1675,In_2236);
xor U1719 (N_1719,In_2487,In_2622);
nor U1720 (N_1720,In_770,In_1671);
and U1721 (N_1721,In_1515,In_636);
nor U1722 (N_1722,In_1534,In_1745);
and U1723 (N_1723,In_2208,In_1019);
nor U1724 (N_1724,In_1566,In_2810);
or U1725 (N_1725,In_2873,In_931);
and U1726 (N_1726,In_1782,In_469);
nor U1727 (N_1727,In_1924,In_2366);
or U1728 (N_1728,In_2000,In_2154);
and U1729 (N_1729,In_2172,In_735);
xor U1730 (N_1730,In_1859,In_428);
xnor U1731 (N_1731,In_2779,In_575);
or U1732 (N_1732,In_1184,In_36);
nor U1733 (N_1733,In_2091,In_117);
or U1734 (N_1734,In_2917,In_2626);
nand U1735 (N_1735,In_2522,In_2933);
and U1736 (N_1736,In_2079,In_2928);
nand U1737 (N_1737,In_1187,In_1398);
xnor U1738 (N_1738,In_79,In_2126);
nand U1739 (N_1739,In_798,In_1986);
nor U1740 (N_1740,In_203,In_86);
or U1741 (N_1741,In_543,In_712);
and U1742 (N_1742,In_253,In_1003);
nor U1743 (N_1743,In_1891,In_1951);
nor U1744 (N_1744,In_360,In_17);
nor U1745 (N_1745,In_148,In_202);
and U1746 (N_1746,In_1990,In_2248);
or U1747 (N_1747,In_1217,In_1753);
or U1748 (N_1748,In_1717,In_2208);
and U1749 (N_1749,In_1361,In_1653);
and U1750 (N_1750,In_1477,In_2337);
xnor U1751 (N_1751,In_2475,In_142);
nor U1752 (N_1752,In_1286,In_656);
or U1753 (N_1753,In_25,In_772);
nor U1754 (N_1754,In_1900,In_1420);
and U1755 (N_1755,In_1697,In_896);
nand U1756 (N_1756,In_2261,In_941);
and U1757 (N_1757,In_2318,In_1744);
xnor U1758 (N_1758,In_1871,In_456);
and U1759 (N_1759,In_2332,In_2281);
and U1760 (N_1760,In_2284,In_398);
and U1761 (N_1761,In_1708,In_154);
nor U1762 (N_1762,In_838,In_948);
xnor U1763 (N_1763,In_1118,In_1706);
nor U1764 (N_1764,In_1014,In_1968);
nand U1765 (N_1765,In_2126,In_255);
nor U1766 (N_1766,In_1138,In_1448);
or U1767 (N_1767,In_72,In_1513);
xor U1768 (N_1768,In_1030,In_1848);
and U1769 (N_1769,In_2997,In_1726);
or U1770 (N_1770,In_43,In_1667);
nand U1771 (N_1771,In_10,In_1196);
or U1772 (N_1772,In_2976,In_735);
xnor U1773 (N_1773,In_2811,In_2056);
nand U1774 (N_1774,In_743,In_811);
nand U1775 (N_1775,In_2388,In_849);
nand U1776 (N_1776,In_2621,In_1174);
nor U1777 (N_1777,In_1309,In_735);
or U1778 (N_1778,In_37,In_1079);
and U1779 (N_1779,In_117,In_2751);
nand U1780 (N_1780,In_895,In_1439);
nor U1781 (N_1781,In_1899,In_2946);
nand U1782 (N_1782,In_591,In_1212);
nor U1783 (N_1783,In_162,In_2046);
nand U1784 (N_1784,In_2868,In_2547);
xnor U1785 (N_1785,In_1097,In_1647);
xnor U1786 (N_1786,In_2695,In_1439);
nand U1787 (N_1787,In_1541,In_74);
xnor U1788 (N_1788,In_1088,In_1621);
nor U1789 (N_1789,In_506,In_2753);
and U1790 (N_1790,In_2863,In_2325);
xnor U1791 (N_1791,In_2825,In_2515);
and U1792 (N_1792,In_1951,In_908);
and U1793 (N_1793,In_165,In_2031);
and U1794 (N_1794,In_2760,In_1989);
xor U1795 (N_1795,In_816,In_2101);
nor U1796 (N_1796,In_1607,In_49);
nand U1797 (N_1797,In_2358,In_266);
nor U1798 (N_1798,In_921,In_2390);
or U1799 (N_1799,In_1684,In_998);
xnor U1800 (N_1800,In_405,In_1770);
or U1801 (N_1801,In_2524,In_2622);
or U1802 (N_1802,In_2235,In_2504);
nor U1803 (N_1803,In_609,In_2643);
or U1804 (N_1804,In_1009,In_348);
or U1805 (N_1805,In_1727,In_1889);
or U1806 (N_1806,In_2271,In_2044);
xor U1807 (N_1807,In_1354,In_2367);
xnor U1808 (N_1808,In_2978,In_2987);
nand U1809 (N_1809,In_2126,In_2001);
nor U1810 (N_1810,In_2489,In_215);
nor U1811 (N_1811,In_1181,In_1137);
nand U1812 (N_1812,In_1699,In_1529);
and U1813 (N_1813,In_1962,In_866);
nor U1814 (N_1814,In_1533,In_1500);
xor U1815 (N_1815,In_1833,In_219);
or U1816 (N_1816,In_604,In_1812);
nand U1817 (N_1817,In_118,In_2082);
and U1818 (N_1818,In_1093,In_454);
nor U1819 (N_1819,In_1352,In_2095);
xor U1820 (N_1820,In_1553,In_123);
or U1821 (N_1821,In_1310,In_2072);
xnor U1822 (N_1822,In_1160,In_2136);
and U1823 (N_1823,In_1844,In_2283);
nor U1824 (N_1824,In_58,In_850);
xor U1825 (N_1825,In_2389,In_2990);
nand U1826 (N_1826,In_2681,In_266);
nor U1827 (N_1827,In_2037,In_651);
or U1828 (N_1828,In_2444,In_755);
nand U1829 (N_1829,In_1115,In_2108);
xor U1830 (N_1830,In_2587,In_1032);
nor U1831 (N_1831,In_2277,In_1230);
or U1832 (N_1832,In_519,In_322);
or U1833 (N_1833,In_2433,In_593);
nand U1834 (N_1834,In_2445,In_684);
xnor U1835 (N_1835,In_1298,In_959);
nand U1836 (N_1836,In_158,In_789);
and U1837 (N_1837,In_509,In_94);
and U1838 (N_1838,In_1164,In_2689);
nor U1839 (N_1839,In_1446,In_2626);
and U1840 (N_1840,In_1780,In_2185);
and U1841 (N_1841,In_160,In_212);
nor U1842 (N_1842,In_2386,In_1022);
nor U1843 (N_1843,In_125,In_1704);
nor U1844 (N_1844,In_1119,In_2761);
nand U1845 (N_1845,In_141,In_1441);
or U1846 (N_1846,In_161,In_520);
or U1847 (N_1847,In_831,In_1324);
nor U1848 (N_1848,In_1986,In_68);
nand U1849 (N_1849,In_2574,In_351);
xnor U1850 (N_1850,In_2588,In_2112);
nand U1851 (N_1851,In_1833,In_1469);
or U1852 (N_1852,In_272,In_118);
xnor U1853 (N_1853,In_1635,In_1708);
nor U1854 (N_1854,In_177,In_2054);
or U1855 (N_1855,In_1593,In_2461);
or U1856 (N_1856,In_973,In_2300);
and U1857 (N_1857,In_1924,In_622);
nor U1858 (N_1858,In_621,In_2044);
and U1859 (N_1859,In_2451,In_468);
and U1860 (N_1860,In_2737,In_1303);
and U1861 (N_1861,In_24,In_2647);
or U1862 (N_1862,In_641,In_1435);
or U1863 (N_1863,In_337,In_443);
nand U1864 (N_1864,In_805,In_1608);
nor U1865 (N_1865,In_305,In_1834);
nand U1866 (N_1866,In_412,In_150);
or U1867 (N_1867,In_1647,In_29);
and U1868 (N_1868,In_2060,In_948);
nand U1869 (N_1869,In_2586,In_1388);
nor U1870 (N_1870,In_504,In_737);
xor U1871 (N_1871,In_1119,In_291);
xor U1872 (N_1872,In_1648,In_2634);
nor U1873 (N_1873,In_1076,In_1396);
nand U1874 (N_1874,In_2707,In_2867);
or U1875 (N_1875,In_1127,In_2127);
and U1876 (N_1876,In_2778,In_2770);
xnor U1877 (N_1877,In_2164,In_222);
and U1878 (N_1878,In_1519,In_2006);
nor U1879 (N_1879,In_1814,In_2460);
or U1880 (N_1880,In_2520,In_2176);
nor U1881 (N_1881,In_2395,In_1543);
nand U1882 (N_1882,In_2639,In_2361);
nand U1883 (N_1883,In_14,In_721);
xnor U1884 (N_1884,In_1724,In_359);
and U1885 (N_1885,In_456,In_125);
xor U1886 (N_1886,In_1172,In_1598);
xnor U1887 (N_1887,In_1111,In_187);
nor U1888 (N_1888,In_105,In_2461);
xnor U1889 (N_1889,In_1597,In_783);
and U1890 (N_1890,In_392,In_2590);
xor U1891 (N_1891,In_1690,In_2971);
and U1892 (N_1892,In_2641,In_1574);
nand U1893 (N_1893,In_2518,In_1160);
or U1894 (N_1894,In_1416,In_2074);
and U1895 (N_1895,In_2865,In_2719);
nor U1896 (N_1896,In_2876,In_1252);
and U1897 (N_1897,In_912,In_719);
xor U1898 (N_1898,In_689,In_2248);
and U1899 (N_1899,In_512,In_2212);
nor U1900 (N_1900,In_401,In_1640);
xor U1901 (N_1901,In_2243,In_2244);
or U1902 (N_1902,In_2924,In_142);
or U1903 (N_1903,In_10,In_2441);
and U1904 (N_1904,In_514,In_804);
xor U1905 (N_1905,In_1349,In_2212);
or U1906 (N_1906,In_1583,In_645);
and U1907 (N_1907,In_2936,In_462);
xor U1908 (N_1908,In_951,In_1936);
nand U1909 (N_1909,In_1022,In_1123);
nor U1910 (N_1910,In_2185,In_2496);
and U1911 (N_1911,In_2921,In_2493);
or U1912 (N_1912,In_554,In_1538);
or U1913 (N_1913,In_1234,In_2481);
nor U1914 (N_1914,In_1077,In_1635);
and U1915 (N_1915,In_23,In_1985);
nand U1916 (N_1916,In_2317,In_2889);
nand U1917 (N_1917,In_353,In_1140);
xor U1918 (N_1918,In_842,In_1911);
nand U1919 (N_1919,In_1102,In_2842);
nand U1920 (N_1920,In_2397,In_720);
xnor U1921 (N_1921,In_485,In_679);
or U1922 (N_1922,In_832,In_2651);
and U1923 (N_1923,In_755,In_2656);
xor U1924 (N_1924,In_2613,In_2515);
xnor U1925 (N_1925,In_1356,In_1973);
and U1926 (N_1926,In_718,In_457);
nor U1927 (N_1927,In_521,In_2404);
nor U1928 (N_1928,In_1358,In_25);
nor U1929 (N_1929,In_2788,In_1289);
xor U1930 (N_1930,In_2172,In_2808);
or U1931 (N_1931,In_634,In_1558);
or U1932 (N_1932,In_2861,In_25);
nand U1933 (N_1933,In_822,In_596);
nor U1934 (N_1934,In_2704,In_2297);
nand U1935 (N_1935,In_350,In_2522);
xor U1936 (N_1936,In_2578,In_212);
or U1937 (N_1937,In_932,In_2394);
and U1938 (N_1938,In_2639,In_648);
nor U1939 (N_1939,In_1731,In_560);
xnor U1940 (N_1940,In_2334,In_2754);
or U1941 (N_1941,In_1858,In_1742);
nand U1942 (N_1942,In_1675,In_1824);
and U1943 (N_1943,In_946,In_2398);
nor U1944 (N_1944,In_181,In_1172);
and U1945 (N_1945,In_654,In_869);
nand U1946 (N_1946,In_1204,In_2140);
xor U1947 (N_1947,In_2309,In_2187);
and U1948 (N_1948,In_2282,In_2772);
or U1949 (N_1949,In_827,In_2971);
or U1950 (N_1950,In_1642,In_548);
or U1951 (N_1951,In_1859,In_2450);
and U1952 (N_1952,In_769,In_2867);
and U1953 (N_1953,In_1853,In_186);
nor U1954 (N_1954,In_790,In_2642);
nor U1955 (N_1955,In_11,In_675);
nand U1956 (N_1956,In_2128,In_2315);
and U1957 (N_1957,In_1716,In_1981);
xor U1958 (N_1958,In_2951,In_629);
and U1959 (N_1959,In_1930,In_2665);
and U1960 (N_1960,In_1254,In_2262);
nor U1961 (N_1961,In_234,In_902);
nor U1962 (N_1962,In_2950,In_225);
nand U1963 (N_1963,In_2970,In_1389);
nor U1964 (N_1964,In_23,In_295);
nor U1965 (N_1965,In_1394,In_1213);
nand U1966 (N_1966,In_1638,In_343);
xnor U1967 (N_1967,In_2630,In_71);
nand U1968 (N_1968,In_2986,In_195);
and U1969 (N_1969,In_1922,In_2746);
xnor U1970 (N_1970,In_2162,In_637);
nand U1971 (N_1971,In_1531,In_1468);
xnor U1972 (N_1972,In_826,In_368);
nor U1973 (N_1973,In_1788,In_655);
nand U1974 (N_1974,In_2522,In_1824);
xnor U1975 (N_1975,In_1838,In_2150);
xnor U1976 (N_1976,In_918,In_98);
and U1977 (N_1977,In_2291,In_2536);
nor U1978 (N_1978,In_705,In_1050);
nand U1979 (N_1979,In_1215,In_2488);
xor U1980 (N_1980,In_2978,In_363);
xor U1981 (N_1981,In_1600,In_1726);
xor U1982 (N_1982,In_466,In_467);
nand U1983 (N_1983,In_2299,In_2857);
nor U1984 (N_1984,In_2544,In_1445);
and U1985 (N_1985,In_766,In_2026);
xnor U1986 (N_1986,In_2530,In_687);
nand U1987 (N_1987,In_619,In_1112);
xor U1988 (N_1988,In_1648,In_1387);
nor U1989 (N_1989,In_744,In_1248);
and U1990 (N_1990,In_247,In_1058);
nand U1991 (N_1991,In_2231,In_2921);
nand U1992 (N_1992,In_1284,In_2733);
nor U1993 (N_1993,In_2694,In_1805);
nor U1994 (N_1994,In_2821,In_1871);
xnor U1995 (N_1995,In_2595,In_1649);
and U1996 (N_1996,In_2124,In_956);
nor U1997 (N_1997,In_1686,In_2826);
nand U1998 (N_1998,In_2263,In_2064);
nor U1999 (N_1999,In_1766,In_1503);
xnor U2000 (N_2000,N_507,N_1070);
nand U2001 (N_2001,N_1027,N_1023);
nor U2002 (N_2002,N_974,N_723);
nor U2003 (N_2003,N_1943,N_428);
xor U2004 (N_2004,N_14,N_1372);
nand U2005 (N_2005,N_365,N_1002);
and U2006 (N_2006,N_31,N_1537);
nand U2007 (N_2007,N_1307,N_1813);
and U2008 (N_2008,N_991,N_1631);
nor U2009 (N_2009,N_205,N_1935);
and U2010 (N_2010,N_608,N_1486);
xnor U2011 (N_2011,N_1086,N_1033);
and U2012 (N_2012,N_874,N_1433);
xor U2013 (N_2013,N_1696,N_165);
or U2014 (N_2014,N_1069,N_1755);
nand U2015 (N_2015,N_923,N_89);
nand U2016 (N_2016,N_795,N_569);
or U2017 (N_2017,N_1513,N_20);
and U2018 (N_2018,N_1300,N_143);
xor U2019 (N_2019,N_1548,N_1677);
and U2020 (N_2020,N_1559,N_130);
xnor U2021 (N_2021,N_60,N_1480);
or U2022 (N_2022,N_34,N_1355);
and U2023 (N_2023,N_40,N_1093);
and U2024 (N_2024,N_439,N_1493);
or U2025 (N_2025,N_1672,N_707);
and U2026 (N_2026,N_1226,N_1990);
and U2027 (N_2027,N_1325,N_1890);
nor U2028 (N_2028,N_551,N_851);
or U2029 (N_2029,N_884,N_588);
nand U2030 (N_2030,N_218,N_1974);
nor U2031 (N_2031,N_761,N_1186);
xor U2032 (N_2032,N_499,N_1338);
nor U2033 (N_2033,N_1152,N_1629);
xnor U2034 (N_2034,N_125,N_1892);
xor U2035 (N_2035,N_987,N_1722);
nand U2036 (N_2036,N_191,N_1075);
or U2037 (N_2037,N_582,N_1636);
and U2038 (N_2038,N_1921,N_1041);
nand U2039 (N_2039,N_1013,N_1438);
nor U2040 (N_2040,N_198,N_533);
nor U2041 (N_2041,N_1572,N_455);
nand U2042 (N_2042,N_378,N_1727);
xor U2043 (N_2043,N_1085,N_999);
and U2044 (N_2044,N_759,N_638);
nand U2045 (N_2045,N_45,N_916);
and U2046 (N_2046,N_1485,N_1663);
xor U2047 (N_2047,N_249,N_654);
nand U2048 (N_2048,N_1803,N_1605);
nor U2049 (N_2049,N_937,N_1136);
or U2050 (N_2050,N_1847,N_285);
nand U2051 (N_2051,N_809,N_726);
nor U2052 (N_2052,N_810,N_1394);
or U2053 (N_2053,N_6,N_212);
or U2054 (N_2054,N_966,N_1877);
nor U2055 (N_2055,N_1331,N_280);
or U2056 (N_2056,N_1774,N_1397);
xnor U2057 (N_2057,N_340,N_1945);
and U2058 (N_2058,N_1930,N_1637);
xor U2059 (N_2059,N_714,N_599);
xnor U2060 (N_2060,N_1362,N_1496);
or U2061 (N_2061,N_1745,N_1734);
xor U2062 (N_2062,N_752,N_716);
xnor U2063 (N_2063,N_1241,N_734);
xnor U2064 (N_2064,N_605,N_467);
or U2065 (N_2065,N_66,N_9);
nor U2066 (N_2066,N_1467,N_1098);
xnor U2067 (N_2067,N_1639,N_393);
or U2068 (N_2068,N_1167,N_1873);
xnor U2069 (N_2069,N_49,N_1077);
nor U2070 (N_2070,N_406,N_1757);
or U2071 (N_2071,N_837,N_1809);
nor U2072 (N_2072,N_1043,N_1267);
or U2073 (N_2073,N_1244,N_1794);
xor U2074 (N_2074,N_990,N_1827);
nand U2075 (N_2075,N_1673,N_237);
and U2076 (N_2076,N_529,N_414);
and U2077 (N_2077,N_836,N_606);
or U2078 (N_2078,N_811,N_894);
or U2079 (N_2079,N_275,N_166);
nand U2080 (N_2080,N_401,N_179);
nand U2081 (N_2081,N_1179,N_1343);
or U2082 (N_2082,N_637,N_1284);
nor U2083 (N_2083,N_1643,N_1991);
nand U2084 (N_2084,N_1345,N_671);
or U2085 (N_2085,N_120,N_1595);
xnor U2086 (N_2086,N_1795,N_1099);
and U2087 (N_2087,N_519,N_308);
nand U2088 (N_2088,N_498,N_1765);
nand U2089 (N_2089,N_772,N_1110);
nand U2090 (N_2090,N_1683,N_902);
nor U2091 (N_2091,N_583,N_1649);
nor U2092 (N_2092,N_971,N_15);
and U2093 (N_2093,N_1109,N_388);
and U2094 (N_2094,N_1501,N_636);
xor U2095 (N_2095,N_1232,N_1478);
nand U2096 (N_2096,N_1315,N_1071);
and U2097 (N_2097,N_33,N_1889);
nor U2098 (N_2098,N_1546,N_1497);
nand U2099 (N_2099,N_980,N_411);
nor U2100 (N_2100,N_173,N_552);
nor U2101 (N_2101,N_348,N_889);
and U2102 (N_2102,N_1804,N_1034);
nand U2103 (N_2103,N_1653,N_438);
nor U2104 (N_2104,N_791,N_230);
and U2105 (N_2105,N_538,N_950);
nor U2106 (N_2106,N_402,N_591);
or U2107 (N_2107,N_1260,N_1404);
nor U2108 (N_2108,N_537,N_1705);
xnor U2109 (N_2109,N_883,N_970);
and U2110 (N_2110,N_1088,N_1703);
nand U2111 (N_2111,N_832,N_1272);
nand U2112 (N_2112,N_598,N_1849);
xor U2113 (N_2113,N_1008,N_1756);
and U2114 (N_2114,N_871,N_592);
nand U2115 (N_2115,N_1479,N_596);
or U2116 (N_2116,N_1987,N_663);
or U2117 (N_2117,N_483,N_964);
nand U2118 (N_2118,N_1276,N_1781);
nand U2119 (N_2119,N_1866,N_463);
nor U2120 (N_2120,N_126,N_209);
nor U2121 (N_2121,N_559,N_859);
nand U2122 (N_2122,N_724,N_254);
and U2123 (N_2123,N_1905,N_119);
or U2124 (N_2124,N_926,N_1992);
nand U2125 (N_2125,N_226,N_914);
and U2126 (N_2126,N_1932,N_1435);
nor U2127 (N_2127,N_1399,N_133);
or U2128 (N_2128,N_641,N_1668);
and U2129 (N_2129,N_407,N_459);
nor U2130 (N_2130,N_1953,N_704);
xor U2131 (N_2131,N_1254,N_1661);
nand U2132 (N_2132,N_376,N_164);
nor U2133 (N_2133,N_1379,N_1100);
xnor U2134 (N_2134,N_381,N_247);
xor U2135 (N_2135,N_202,N_1514);
xnor U2136 (N_2136,N_1360,N_593);
and U2137 (N_2137,N_140,N_1862);
xnor U2138 (N_2138,N_1221,N_302);
or U2139 (N_2139,N_992,N_1725);
nor U2140 (N_2140,N_62,N_52);
nor U2141 (N_2141,N_786,N_1861);
nor U2142 (N_2142,N_925,N_1997);
nand U2143 (N_2143,N_615,N_1224);
nor U2144 (N_2144,N_828,N_1441);
nor U2145 (N_2145,N_1555,N_1724);
nor U2146 (N_2146,N_377,N_1);
and U2147 (N_2147,N_855,N_972);
nor U2148 (N_2148,N_509,N_193);
nand U2149 (N_2149,N_135,N_1912);
or U2150 (N_2150,N_1623,N_1451);
and U2151 (N_2151,N_610,N_154);
and U2152 (N_2152,N_566,N_354);
or U2153 (N_2153,N_805,N_118);
nor U2154 (N_2154,N_703,N_1090);
and U2155 (N_2155,N_1528,N_1747);
nor U2156 (N_2156,N_760,N_693);
or U2157 (N_2157,N_635,N_1334);
xnor U2158 (N_2158,N_907,N_272);
and U2159 (N_2159,N_1908,N_1996);
and U2160 (N_2160,N_1837,N_576);
or U2161 (N_2161,N_690,N_1038);
xnor U2162 (N_2162,N_1556,N_1481);
or U2163 (N_2163,N_1453,N_211);
nor U2164 (N_2164,N_1011,N_763);
nand U2165 (N_2165,N_1473,N_260);
and U2166 (N_2166,N_1440,N_1679);
or U2167 (N_2167,N_784,N_90);
nor U2168 (N_2168,N_67,N_1158);
or U2169 (N_2169,N_1302,N_341);
nand U2170 (N_2170,N_417,N_661);
and U2171 (N_2171,N_124,N_520);
nand U2172 (N_2172,N_1618,N_542);
nand U2173 (N_2173,N_651,N_1091);
and U2174 (N_2174,N_1922,N_1194);
nand U2175 (N_2175,N_1193,N_187);
and U2176 (N_2176,N_1601,N_1906);
or U2177 (N_2177,N_122,N_1238);
or U2178 (N_2178,N_1891,N_1460);
xor U2179 (N_2179,N_1462,N_1475);
xor U2180 (N_2180,N_1979,N_1249);
nand U2181 (N_2181,N_1561,N_1352);
nand U2182 (N_2182,N_1660,N_539);
xnor U2183 (N_2183,N_514,N_1762);
nand U2184 (N_2184,N_944,N_601);
xnor U2185 (N_2185,N_1412,N_330);
and U2186 (N_2186,N_276,N_684);
or U2187 (N_2187,N_1170,N_1856);
or U2188 (N_2188,N_829,N_976);
or U2189 (N_2189,N_584,N_833);
nand U2190 (N_2190,N_785,N_1309);
xnor U2191 (N_2191,N_258,N_1209);
or U2192 (N_2192,N_76,N_936);
nand U2193 (N_2193,N_1916,N_1426);
xnor U2194 (N_2194,N_1955,N_1045);
nor U2195 (N_2195,N_1645,N_149);
xnor U2196 (N_2196,N_962,N_1787);
and U2197 (N_2197,N_602,N_336);
nand U2198 (N_2198,N_528,N_818);
nor U2199 (N_2199,N_1106,N_735);
xnor U2200 (N_2200,N_148,N_400);
and U2201 (N_2201,N_1285,N_982);
or U2202 (N_2202,N_1468,N_1036);
and U2203 (N_2203,N_623,N_1865);
nand U2204 (N_2204,N_312,N_327);
nand U2205 (N_2205,N_462,N_1223);
and U2206 (N_2206,N_452,N_1584);
nor U2207 (N_2207,N_1278,N_1189);
and U2208 (N_2208,N_1699,N_587);
xnor U2209 (N_2209,N_632,N_1753);
nor U2210 (N_2210,N_117,N_1658);
nor U2211 (N_2211,N_287,N_1929);
nor U2212 (N_2212,N_857,N_41);
and U2213 (N_2213,N_465,N_1899);
or U2214 (N_2214,N_956,N_969);
nand U2215 (N_2215,N_1886,N_109);
xnor U2216 (N_2216,N_78,N_207);
or U2217 (N_2217,N_614,N_367);
and U2218 (N_2218,N_1554,N_384);
nor U2219 (N_2219,N_274,N_1293);
nand U2220 (N_2220,N_756,N_255);
nor U2221 (N_2221,N_178,N_1967);
and U2222 (N_2222,N_310,N_780);
nor U2223 (N_2223,N_93,N_1700);
nand U2224 (N_2224,N_1926,N_328);
nand U2225 (N_2225,N_1835,N_850);
nor U2226 (N_2226,N_466,N_804);
nand U2227 (N_2227,N_282,N_1469);
or U2228 (N_2228,N_1978,N_1744);
xor U2229 (N_2229,N_170,N_1061);
or U2230 (N_2230,N_1571,N_432);
nand U2231 (N_2231,N_1078,N_29);
xor U2232 (N_2232,N_374,N_113);
or U2233 (N_2233,N_1614,N_1680);
xnor U2234 (N_2234,N_199,N_1058);
or U2235 (N_2235,N_418,N_182);
or U2236 (N_2236,N_1855,N_397);
xor U2237 (N_2237,N_1081,N_560);
and U2238 (N_2238,N_293,N_256);
xnor U2239 (N_2239,N_572,N_1321);
nand U2240 (N_2240,N_1918,N_1398);
nand U2241 (N_2241,N_1946,N_94);
nand U2242 (N_2242,N_168,N_1901);
and U2243 (N_2243,N_1697,N_186);
and U2244 (N_2244,N_891,N_1723);
nor U2245 (N_2245,N_561,N_1796);
nor U2246 (N_2246,N_317,N_1743);
nand U2247 (N_2247,N_1826,N_860);
xor U2248 (N_2248,N_856,N_1143);
nor U2249 (N_2249,N_1569,N_821);
or U2250 (N_2250,N_161,N_1124);
xnor U2251 (N_2251,N_1080,N_1247);
nand U2252 (N_2252,N_22,N_1739);
nand U2253 (N_2253,N_547,N_1760);
xnor U2254 (N_2254,N_382,N_1429);
nor U2255 (N_2255,N_17,N_1993);
nand U2256 (N_2256,N_1121,N_1025);
xor U2257 (N_2257,N_1472,N_426);
xnor U2258 (N_2258,N_1502,N_1576);
nand U2259 (N_2259,N_1879,N_872);
and U2260 (N_2260,N_18,N_975);
xor U2261 (N_2261,N_1609,N_796);
nor U2262 (N_2262,N_32,N_1356);
xor U2263 (N_2263,N_567,N_908);
nor U2264 (N_2264,N_394,N_160);
nor U2265 (N_2265,N_1103,N_1000);
nand U2266 (N_2266,N_46,N_1834);
xnor U2267 (N_2267,N_421,N_441);
or U2268 (N_2268,N_611,N_176);
and U2269 (N_2269,N_121,N_1937);
xor U2270 (N_2270,N_1188,N_1597);
and U2271 (N_2271,N_677,N_1965);
or U2272 (N_2272,N_1730,N_298);
nand U2273 (N_2273,N_1126,N_1268);
and U2274 (N_2274,N_217,N_1793);
nor U2275 (N_2275,N_666,N_398);
and U2276 (N_2276,N_1816,N_1613);
xnor U2277 (N_2277,N_1659,N_1802);
nor U2278 (N_2278,N_1195,N_1196);
and U2279 (N_2279,N_817,N_1893);
and U2280 (N_2280,N_744,N_129);
nand U2281 (N_2281,N_1424,N_842);
nand U2282 (N_2282,N_1752,N_720);
nor U2283 (N_2283,N_1652,N_1526);
nand U2284 (N_2284,N_1940,N_1369);
xnor U2285 (N_2285,N_1120,N_1366);
or U2286 (N_2286,N_1140,N_831);
xor U2287 (N_2287,N_502,N_1748);
xnor U2288 (N_2288,N_1135,N_1148);
nor U2289 (N_2289,N_1494,N_1552);
nand U2290 (N_2290,N_1329,N_1430);
or U2291 (N_2291,N_453,N_1344);
or U2292 (N_2292,N_138,N_1602);
or U2293 (N_2293,N_82,N_1067);
xor U2294 (N_2294,N_688,N_1262);
and U2295 (N_2295,N_100,N_1570);
nor U2296 (N_2296,N_1544,N_1159);
nand U2297 (N_2297,N_997,N_319);
xnor U2298 (N_2298,N_482,N_912);
or U2299 (N_2299,N_1138,N_409);
and U2300 (N_2300,N_977,N_7);
or U2301 (N_2301,N_1966,N_655);
or U2302 (N_2302,N_1387,N_574);
and U2303 (N_2303,N_1587,N_1780);
and U2304 (N_2304,N_19,N_675);
or U2305 (N_2305,N_151,N_1704);
xor U2306 (N_2306,N_996,N_1647);
and U2307 (N_2307,N_579,N_669);
xor U2308 (N_2308,N_361,N_1201);
xor U2309 (N_2309,N_1280,N_1934);
and U2310 (N_2310,N_1779,N_174);
nand U2311 (N_2311,N_1985,N_722);
nand U2312 (N_2312,N_1784,N_1145);
nor U2313 (N_2313,N_1422,N_815);
or U2314 (N_2314,N_1667,N_150);
xnor U2315 (N_2315,N_223,N_1206);
nor U2316 (N_2316,N_934,N_1589);
nor U2317 (N_2317,N_64,N_47);
or U2318 (N_2318,N_779,N_85);
and U2319 (N_2319,N_1844,N_1577);
xor U2320 (N_2320,N_1738,N_948);
nand U2321 (N_2321,N_1001,N_1821);
nand U2322 (N_2322,N_1731,N_156);
nand U2323 (N_2323,N_612,N_927);
xnor U2324 (N_2324,N_493,N_1068);
nand U2325 (N_2325,N_1251,N_471);
and U2326 (N_2326,N_77,N_988);
nor U2327 (N_2327,N_812,N_1217);
xor U2328 (N_2328,N_291,N_718);
or U2329 (N_2329,N_1212,N_711);
nor U2330 (N_2330,N_834,N_1388);
and U2331 (N_2331,N_1341,N_1060);
xor U2332 (N_2332,N_1686,N_581);
and U2333 (N_2333,N_227,N_946);
nor U2334 (N_2334,N_1644,N_861);
xor U2335 (N_2335,N_1348,N_38);
xnor U2336 (N_2336,N_290,N_503);
and U2337 (N_2337,N_864,N_682);
or U2338 (N_2338,N_43,N_1007);
or U2339 (N_2339,N_803,N_512);
or U2340 (N_2340,N_571,N_1550);
nand U2341 (N_2341,N_712,N_1600);
and U2342 (N_2342,N_292,N_1994);
xor U2343 (N_2343,N_717,N_757);
nor U2344 (N_2344,N_774,N_1326);
nand U2345 (N_2345,N_307,N_1621);
nand U2346 (N_2346,N_639,N_656);
xnor U2347 (N_2347,N_534,N_1530);
nor U2348 (N_2348,N_771,N_3);
xnor U2349 (N_2349,N_1289,N_316);
nor U2350 (N_2350,N_306,N_1487);
or U2351 (N_2351,N_412,N_108);
xor U2352 (N_2352,N_96,N_158);
or U2353 (N_2353,N_981,N_281);
or U2354 (N_2354,N_1028,N_1056);
and U2355 (N_2355,N_103,N_1638);
and U2356 (N_2356,N_123,N_1250);
or U2357 (N_2357,N_269,N_1287);
nor U2358 (N_2358,N_1153,N_1852);
nand U2359 (N_2359,N_391,N_1761);
and U2360 (N_2360,N_1928,N_349);
nand U2361 (N_2361,N_1482,N_1392);
nand U2362 (N_2362,N_955,N_1541);
nand U2363 (N_2363,N_284,N_1845);
nor U2364 (N_2364,N_1476,N_1671);
and U2365 (N_2365,N_345,N_208);
nand U2366 (N_2366,N_216,N_668);
or U2367 (N_2367,N_928,N_886);
or U2368 (N_2368,N_1830,N_777);
and U2369 (N_2369,N_1707,N_1773);
nand U2370 (N_2370,N_1735,N_1583);
nand U2371 (N_2371,N_603,N_1690);
and U2372 (N_2372,N_16,N_144);
nor U2373 (N_2373,N_568,N_892);
nor U2374 (N_2374,N_1228,N_359);
or U2375 (N_2375,N_1057,N_1311);
and U2376 (N_2376,N_1783,N_525);
or U2377 (N_2377,N_913,N_1831);
and U2378 (N_2378,N_1895,N_1346);
xor U2379 (N_2379,N_650,N_1452);
nor U2380 (N_2380,N_1829,N_1176);
nor U2381 (N_2381,N_1192,N_1792);
xor U2382 (N_2382,N_1168,N_1778);
and U2383 (N_2383,N_1558,N_800);
xnor U2384 (N_2384,N_515,N_1029);
or U2385 (N_2385,N_301,N_1535);
nand U2386 (N_2386,N_480,N_672);
and U2387 (N_2387,N_1858,N_196);
nand U2388 (N_2388,N_1962,N_1187);
xnor U2389 (N_2389,N_1048,N_1182);
and U2390 (N_2390,N_827,N_1233);
xnor U2391 (N_2391,N_1459,N_372);
nor U2392 (N_2392,N_536,N_1938);
or U2393 (N_2393,N_686,N_1466);
and U2394 (N_2394,N_1364,N_396);
xnor U2395 (N_2395,N_609,N_1712);
xnor U2396 (N_2396,N_145,N_1790);
nor U2397 (N_2397,N_1777,N_524);
nor U2398 (N_2398,N_1371,N_39);
xor U2399 (N_2399,N_1305,N_1290);
nor U2400 (N_2400,N_573,N_1620);
or U2401 (N_2401,N_825,N_732);
nand U2402 (N_2402,N_1218,N_705);
or U2403 (N_2403,N_945,N_887);
nand U2404 (N_2404,N_1910,N_1566);
and U2405 (N_2405,N_1654,N_911);
xor U2406 (N_2406,N_1913,N_127);
nor U2407 (N_2407,N_1205,N_339);
and U2408 (N_2408,N_1624,N_1439);
nor U2409 (N_2409,N_770,N_1678);
and U2410 (N_2410,N_1031,N_1857);
nor U2411 (N_2411,N_128,N_1177);
nor U2412 (N_2412,N_408,N_1490);
xor U2413 (N_2413,N_1574,N_1763);
xor U2414 (N_2414,N_575,N_344);
xor U2415 (N_2415,N_564,N_1178);
xor U2416 (N_2416,N_1607,N_768);
and U2417 (N_2417,N_983,N_1022);
xor U2418 (N_2418,N_1052,N_1204);
xnor U2419 (N_2419,N_882,N_1919);
xor U2420 (N_2420,N_1622,N_1791);
or U2421 (N_2421,N_157,N_1592);
xnor U2422 (N_2422,N_1415,N_236);
nand U2423 (N_2423,N_337,N_1959);
nor U2424 (N_2424,N_875,N_1651);
nand U2425 (N_2425,N_511,N_1180);
and U2426 (N_2426,N_315,N_1181);
or U2427 (N_2427,N_1044,N_530);
and U2428 (N_2428,N_1824,N_826);
nor U2429 (N_2429,N_358,N_1785);
nand U2430 (N_2430,N_1894,N_364);
and U2431 (N_2431,N_200,N_58);
nor U2432 (N_2432,N_862,N_1538);
or U2433 (N_2433,N_1606,N_1411);
xnor U2434 (N_2434,N_1568,N_1079);
nor U2435 (N_2435,N_1391,N_1005);
xor U2436 (N_2436,N_797,N_1635);
nand U2437 (N_2437,N_824,N_1484);
nor U2438 (N_2438,N_1681,N_895);
and U2439 (N_2439,N_1715,N_674);
nor U2440 (N_2440,N_1619,N_1114);
or U2441 (N_2441,N_457,N_740);
xor U2442 (N_2442,N_965,N_680);
and U2443 (N_2443,N_1258,N_527);
or U2444 (N_2444,N_590,N_848);
xnor U2445 (N_2445,N_1450,N_1173);
xnor U2446 (N_2446,N_286,N_116);
and U2447 (N_2447,N_1129,N_1581);
xor U2448 (N_2448,N_1308,N_1340);
xnor U2449 (N_2449,N_1656,N_295);
nor U2450 (N_2450,N_1642,N_1531);
xnor U2451 (N_2451,N_477,N_1872);
and U2452 (N_2452,N_1925,N_1259);
and U2453 (N_2453,N_44,N_1694);
xor U2454 (N_2454,N_472,N_1952);
or U2455 (N_2455,N_1693,N_648);
nor U2456 (N_2456,N_183,N_775);
nand U2457 (N_2457,N_373,N_1508);
xor U2458 (N_2458,N_1236,N_268);
and U2459 (N_2459,N_699,N_1936);
or U2460 (N_2460,N_368,N_429);
nor U2461 (N_2461,N_985,N_748);
xnor U2462 (N_2462,N_496,N_1611);
nor U2463 (N_2463,N_1104,N_1567);
nor U2464 (N_2464,N_1983,N_1527);
nor U2465 (N_2465,N_1215,N_1417);
xnor U2466 (N_2466,N_0,N_1819);
nor U2467 (N_2467,N_1039,N_1522);
xor U2468 (N_2468,N_1449,N_673);
and U2469 (N_2469,N_1507,N_1580);
and U2470 (N_2470,N_334,N_177);
or U2471 (N_2471,N_1949,N_1225);
nor U2472 (N_2472,N_1732,N_630);
and U2473 (N_2473,N_1786,N_1207);
nand U2474 (N_2474,N_1718,N_30);
nand U2475 (N_2475,N_180,N_1339);
xor U2476 (N_2476,N_1320,N_808);
or U2477 (N_2477,N_246,N_1630);
and U2478 (N_2478,N_194,N_1702);
or U2479 (N_2479,N_1533,N_1046);
nor U2480 (N_2480,N_1270,N_355);
xnor U2481 (N_2481,N_504,N_1134);
or U2482 (N_2482,N_930,N_68);
or U2483 (N_2483,N_185,N_1463);
xnor U2484 (N_2484,N_210,N_1939);
nand U2485 (N_2485,N_1483,N_963);
xor U2486 (N_2486,N_231,N_1948);
nand U2487 (N_2487,N_1020,N_1385);
xnor U2488 (N_2488,N_1701,N_1876);
or U2489 (N_2489,N_1403,N_220);
or U2490 (N_2490,N_1303,N_434);
nor U2491 (N_2491,N_941,N_1971);
xor U2492 (N_2492,N_1669,N_1018);
or U2493 (N_2493,N_1853,N_1884);
nand U2494 (N_2494,N_1503,N_369);
nor U2495 (N_2495,N_715,N_877);
nand U2496 (N_2496,N_80,N_1767);
or U2497 (N_2497,N_189,N_1163);
xor U2498 (N_2498,N_313,N_681);
xor U2499 (N_2499,N_206,N_1933);
nand U2500 (N_2500,N_846,N_197);
or U2501 (N_2501,N_1736,N_1279);
nand U2502 (N_2502,N_1634,N_1573);
or U2503 (N_2503,N_1900,N_1274);
xor U2504 (N_2504,N_1401,N_618);
xor U2505 (N_2505,N_1982,N_1828);
xor U2506 (N_2506,N_697,N_1184);
nand U2507 (N_2507,N_261,N_169);
nor U2508 (N_2508,N_456,N_1812);
xor U2509 (N_2509,N_1425,N_1814);
xnor U2510 (N_2510,N_203,N_1456);
nand U2511 (N_2511,N_1617,N_321);
xor U2512 (N_2512,N_1917,N_1771);
nand U2513 (N_2513,N_565,N_1454);
and U2514 (N_2514,N_435,N_729);
nor U2515 (N_2515,N_470,N_132);
and U2516 (N_2516,N_823,N_1800);
or U2517 (N_2517,N_224,N_21);
nor U2518 (N_2518,N_1208,N_517);
or U2519 (N_2519,N_83,N_691);
xnor U2520 (N_2520,N_1575,N_1019);
xnor U2521 (N_2521,N_181,N_1214);
nor U2522 (N_2522,N_1942,N_1427);
nor U2523 (N_2523,N_1295,N_776);
nand U2524 (N_2524,N_1864,N_1604);
xor U2525 (N_2525,N_957,N_56);
and U2526 (N_2526,N_324,N_737);
nor U2527 (N_2527,N_153,N_1868);
nand U2528 (N_2528,N_1594,N_1860);
or U2529 (N_2529,N_175,N_713);
nand U2530 (N_2530,N_1788,N_544);
and U2531 (N_2531,N_640,N_1410);
and U2532 (N_2532,N_1665,N_12);
nand U2533 (N_2533,N_1534,N_1275);
nor U2534 (N_2534,N_570,N_1640);
and U2535 (N_2535,N_1365,N_1689);
or U2536 (N_2536,N_1157,N_192);
nand U2537 (N_2537,N_1695,N_589);
or U2538 (N_2538,N_343,N_1119);
or U2539 (N_2539,N_562,N_1968);
nor U2540 (N_2540,N_1687,N_736);
or U2541 (N_2541,N_1393,N_868);
nor U2542 (N_2542,N_943,N_1520);
nor U2543 (N_2543,N_1875,N_1414);
nand U2544 (N_2544,N_1003,N_1729);
and U2545 (N_2545,N_35,N_1565);
nor U2546 (N_2546,N_695,N_1842);
nand U2547 (N_2547,N_1229,N_619);
and U2548 (N_2548,N_142,N_676);
and U2549 (N_2549,N_787,N_1495);
or U2550 (N_2550,N_1969,N_847);
or U2551 (N_2551,N_1909,N_799);
nor U2552 (N_2552,N_1342,N_1840);
and U2553 (N_2553,N_248,N_1907);
or U2554 (N_2554,N_1964,N_1582);
and U2555 (N_2555,N_664,N_1301);
nor U2556 (N_2556,N_1286,N_1769);
and U2557 (N_2557,N_305,N_112);
nand U2558 (N_2558,N_1162,N_1065);
nand U2559 (N_2559,N_1655,N_1318);
xnor U2560 (N_2560,N_251,N_1749);
nand U2561 (N_2561,N_451,N_893);
or U2562 (N_2562,N_1082,N_917);
nand U2563 (N_2563,N_1474,N_554);
xnor U2564 (N_2564,N_1625,N_867);
xor U2565 (N_2565,N_1132,N_201);
xor U2566 (N_2566,N_993,N_1458);
xor U2567 (N_2567,N_61,N_240);
xnor U2568 (N_2568,N_1728,N_1980);
xor U2569 (N_2569,N_1257,N_333);
nor U2570 (N_2570,N_652,N_1579);
nand U2571 (N_2571,N_431,N_450);
and U2572 (N_2572,N_422,N_342);
nor U2573 (N_2573,N_228,N_1130);
nor U2574 (N_2574,N_243,N_702);
and U2575 (N_2575,N_1396,N_131);
or U2576 (N_2576,N_1676,N_1944);
nand U2577 (N_2577,N_1759,N_1553);
nor U2578 (N_2578,N_214,N_755);
and U2579 (N_2579,N_1198,N_765);
nand U2580 (N_2580,N_1822,N_91);
and U2581 (N_2581,N_1095,N_1549);
and U2582 (N_2582,N_219,N_1742);
nor U2583 (N_2583,N_1758,N_403);
nand U2584 (N_2584,N_1294,N_1235);
or U2585 (N_2585,N_900,N_215);
nor U2586 (N_2586,N_338,N_844);
and U2587 (N_2587,N_580,N_549);
nor U2588 (N_2588,N_629,N_1989);
and U2589 (N_2589,N_1436,N_70);
xor U2590 (N_2590,N_1107,N_1200);
nand U2591 (N_2591,N_696,N_81);
or U2592 (N_2592,N_709,N_513);
or U2593 (N_2593,N_1096,N_1073);
and U2594 (N_2594,N_1199,N_766);
nor U2595 (N_2595,N_1141,N_819);
and U2596 (N_2596,N_1525,N_420);
and U2597 (N_2597,N_1710,N_1423);
nand U2598 (N_2598,N_852,N_806);
and U2599 (N_2599,N_624,N_1838);
xor U2600 (N_2600,N_25,N_822);
and U2601 (N_2601,N_1820,N_1882);
or U2602 (N_2602,N_213,N_404);
nor U2603 (N_2603,N_1256,N_238);
nand U2604 (N_2604,N_942,N_959);
nor U2605 (N_2605,N_1871,N_1915);
nor U2606 (N_2606,N_1789,N_622);
or U2607 (N_2607,N_814,N_95);
nor U2608 (N_2608,N_1288,N_1375);
or U2609 (N_2609,N_1947,N_389);
or U2610 (N_2610,N_516,N_1243);
nand U2611 (N_2611,N_141,N_1142);
nand U2612 (N_2612,N_1878,N_678);
xor U2613 (N_2613,N_1363,N_1444);
and U2614 (N_2614,N_162,N_933);
or U2615 (N_2615,N_1183,N_289);
and U2616 (N_2616,N_727,N_721);
or U2617 (N_2617,N_1445,N_1833);
or U2618 (N_2618,N_461,N_27);
or U2619 (N_2619,N_1632,N_473);
nand U2620 (N_2620,N_947,N_665);
or U2621 (N_2621,N_1519,N_523);
nor U2622 (N_2622,N_440,N_577);
or U2623 (N_2623,N_1951,N_74);
or U2624 (N_2624,N_1010,N_845);
and U2625 (N_2625,N_508,N_1304);
nor U2626 (N_2626,N_989,N_1708);
nor U2627 (N_2627,N_1407,N_1431);
nor U2628 (N_2628,N_898,N_1691);
or U2629 (N_2629,N_557,N_1815);
xor U2630 (N_2630,N_1313,N_1202);
and U2631 (N_2631,N_5,N_1155);
nand U2632 (N_2632,N_1354,N_53);
or U2633 (N_2633,N_8,N_423);
or U2634 (N_2634,N_1190,N_679);
or U2635 (N_2635,N_444,N_1941);
or U2636 (N_2636,N_88,N_1818);
nand U2637 (N_2637,N_634,N_1488);
xnor U2638 (N_2638,N_1863,N_555);
nor U2639 (N_2639,N_437,N_628);
xnor U2640 (N_2640,N_1832,N_1506);
nor U2641 (N_2641,N_489,N_1032);
xnor U2642 (N_2642,N_481,N_436);
or U2643 (N_2643,N_870,N_488);
or U2644 (N_2644,N_1648,N_938);
nand U2645 (N_2645,N_753,N_1977);
or U2646 (N_2646,N_951,N_1543);
nand U2647 (N_2647,N_1986,N_1477);
and U2648 (N_2648,N_79,N_521);
xor U2649 (N_2649,N_1102,N_1805);
and U2650 (N_2650,N_546,N_204);
xor U2651 (N_2651,N_1998,N_163);
and U2652 (N_2652,N_167,N_813);
and U2653 (N_2653,N_105,N_1386);
nor U2654 (N_2654,N_474,N_357);
nor U2655 (N_2655,N_1657,N_1245);
xnor U2656 (N_2656,N_257,N_1035);
nor U2657 (N_2657,N_1911,N_1087);
nand U2658 (N_2658,N_1612,N_413);
and U2659 (N_2659,N_1706,N_505);
nor U2660 (N_2660,N_931,N_1317);
or U2661 (N_2661,N_1113,N_1675);
and U2662 (N_2662,N_1185,N_1314);
or U2663 (N_2663,N_1359,N_1266);
nor U2664 (N_2664,N_229,N_1563);
xnor U2665 (N_2665,N_1012,N_1172);
nand U2666 (N_2666,N_1381,N_1242);
nand U2667 (N_2667,N_1234,N_1101);
xnor U2668 (N_2668,N_314,N_278);
and U2669 (N_2669,N_1536,N_518);
and U2670 (N_2670,N_954,N_1521);
and U2671 (N_2671,N_1817,N_1169);
or U2672 (N_2672,N_356,N_1666);
or U2673 (N_2673,N_1248,N_1511);
and U2674 (N_2674,N_1171,N_479);
and U2675 (N_2675,N_1400,N_1246);
nor U2676 (N_2676,N_1150,N_863);
and U2677 (N_2677,N_586,N_1801);
nor U2678 (N_2678,N_57,N_37);
and U2679 (N_2679,N_751,N_147);
or U2680 (N_2680,N_840,N_1263);
nor U2681 (N_2681,N_1291,N_152);
or U2682 (N_2682,N_1021,N_1292);
nand U2683 (N_2683,N_627,N_1147);
and U2684 (N_2684,N_10,N_1973);
nand U2685 (N_2685,N_932,N_110);
and U2686 (N_2686,N_758,N_347);
nand U2687 (N_2687,N_1419,N_1455);
or U2688 (N_2688,N_532,N_1903);
xnor U2689 (N_2689,N_395,N_1118);
and U2690 (N_2690,N_778,N_1733);
nand U2691 (N_2691,N_487,N_1351);
and U2692 (N_2692,N_670,N_1596);
xor U2693 (N_2693,N_1265,N_1867);
and U2694 (N_2694,N_890,N_492);
xor U2695 (N_2695,N_522,N_1564);
or U2696 (N_2696,N_233,N_738);
nor U2697 (N_2697,N_816,N_616);
or U2698 (N_2698,N_1599,N_299);
and U2699 (N_2699,N_48,N_1297);
nand U2700 (N_2700,N_1881,N_694);
nand U2701 (N_2701,N_1633,N_1316);
nor U2702 (N_2702,N_195,N_995);
nor U2703 (N_2703,N_415,N_1956);
xor U2704 (N_2704,N_794,N_643);
or U2705 (N_2705,N_1322,N_1721);
xnor U2706 (N_2706,N_1846,N_1428);
nor U2707 (N_2707,N_710,N_728);
nand U2708 (N_2708,N_485,N_392);
or U2709 (N_2709,N_1766,N_172);
or U2710 (N_2710,N_1823,N_1395);
and U2711 (N_2711,N_708,N_2);
xor U2712 (N_2712,N_458,N_190);
xnor U2713 (N_2713,N_657,N_111);
nand U2714 (N_2714,N_749,N_1711);
nand U2715 (N_2715,N_1854,N_69);
or U2716 (N_2716,N_73,N_594);
or U2717 (N_2717,N_841,N_351);
nand U2718 (N_2718,N_1808,N_320);
nor U2719 (N_2719,N_1064,N_1122);
nand U2720 (N_2720,N_1586,N_332);
xor U2721 (N_2721,N_897,N_1888);
xor U2722 (N_2722,N_1457,N_115);
xor U2723 (N_2723,N_1750,N_1353);
nand U2724 (N_2724,N_1500,N_585);
or U2725 (N_2725,N_424,N_1447);
and U2726 (N_2726,N_1017,N_1239);
xnor U2727 (N_2727,N_1255,N_1545);
or U2728 (N_2728,N_790,N_1957);
or U2729 (N_2729,N_788,N_448);
xnor U2730 (N_2730,N_1972,N_1499);
and U2731 (N_2731,N_1836,N_380);
xnor U2732 (N_2732,N_1551,N_921);
and U2733 (N_2733,N_1442,N_1434);
nand U2734 (N_2734,N_1810,N_952);
and U2735 (N_2735,N_1981,N_1330);
or U2736 (N_2736,N_1726,N_1999);
and U2737 (N_2737,N_259,N_13);
nand U2738 (N_2738,N_362,N_1146);
or U2739 (N_2739,N_769,N_1641);
nand U2740 (N_2740,N_297,N_23);
or U2741 (N_2741,N_706,N_28);
and U2742 (N_2742,N_460,N_1963);
nor U2743 (N_2743,N_888,N_288);
or U2744 (N_2744,N_1598,N_387);
or U2745 (N_2745,N_647,N_910);
or U2746 (N_2746,N_901,N_1139);
or U2747 (N_2747,N_1333,N_309);
nor U2748 (N_2748,N_1376,N_1220);
and U2749 (N_2749,N_263,N_700);
and U2750 (N_2750,N_1015,N_658);
xnor U2751 (N_2751,N_1841,N_484);
nand U2752 (N_2752,N_906,N_478);
and U2753 (N_2753,N_26,N_1839);
nor U2754 (N_2754,N_323,N_51);
nand U2755 (N_2755,N_1053,N_1950);
or U2756 (N_2756,N_86,N_294);
or U2757 (N_2757,N_97,N_1688);
nand U2758 (N_2758,N_1125,N_159);
xor U2759 (N_2759,N_1253,N_1324);
xor U2760 (N_2760,N_101,N_820);
nor U2761 (N_2761,N_692,N_1283);
xnor U2762 (N_2762,N_866,N_683);
xor U2763 (N_2763,N_265,N_476);
nor U2764 (N_2764,N_979,N_1014);
nand U2765 (N_2765,N_922,N_1874);
xnor U2766 (N_2766,N_865,N_935);
and U2767 (N_2767,N_99,N_659);
xnor U2768 (N_2768,N_1350,N_1807);
or U2769 (N_2769,N_1437,N_445);
and U2770 (N_2770,N_1885,N_1927);
xnor U2771 (N_2771,N_667,N_1509);
xor U2772 (N_2772,N_1464,N_245);
xnor U2773 (N_2773,N_1931,N_242);
nor U2774 (N_2774,N_188,N_1115);
nand U2775 (N_2775,N_1377,N_1588);
nor U2776 (N_2776,N_65,N_698);
or U2777 (N_2777,N_978,N_915);
or U2778 (N_2778,N_642,N_802);
xnor U2779 (N_2779,N_1261,N_1737);
and U2780 (N_2780,N_1421,N_495);
and U2781 (N_2781,N_1323,N_1799);
or U2782 (N_2782,N_1156,N_1518);
nor U2783 (N_2783,N_1674,N_1740);
and U2784 (N_2784,N_1896,N_416);
or U2785 (N_2785,N_442,N_1465);
and U2786 (N_2786,N_835,N_134);
nor U2787 (N_2787,N_491,N_613);
nor U2788 (N_2788,N_1319,N_318);
xor U2789 (N_2789,N_1510,N_731);
and U2790 (N_2790,N_858,N_644);
nand U2791 (N_2791,N_621,N_1374);
or U2792 (N_2792,N_1776,N_548);
or U2793 (N_2793,N_1505,N_903);
nand U2794 (N_2794,N_880,N_1231);
and U2795 (N_2795,N_1111,N_961);
or U2796 (N_2796,N_1843,N_55);
xor U2797 (N_2797,N_541,N_1337);
nor U2798 (N_2798,N_1072,N_1133);
or U2799 (N_2799,N_1175,N_1047);
or U2800 (N_2800,N_1850,N_750);
xnor U2801 (N_2801,N_1970,N_1898);
or U2802 (N_2802,N_379,N_107);
and U2803 (N_2803,N_1367,N_1117);
nand U2804 (N_2804,N_277,N_1529);
nor U2805 (N_2805,N_446,N_1650);
xor U2806 (N_2806,N_1306,N_754);
nor U2807 (N_2807,N_84,N_1416);
xnor U2808 (N_2808,N_994,N_494);
nand U2809 (N_2809,N_1976,N_1076);
xnor U2810 (N_2810,N_1382,N_1562);
nor U2811 (N_2811,N_1380,N_1213);
nor U2812 (N_2812,N_1515,N_526);
xnor U2813 (N_2813,N_350,N_1995);
or U2814 (N_2814,N_685,N_1273);
and U2815 (N_2815,N_1084,N_1361);
nor U2816 (N_2816,N_486,N_843);
or U2817 (N_2817,N_1591,N_304);
or U2818 (N_2818,N_1009,N_960);
or U2819 (N_2819,N_1349,N_653);
nor U2820 (N_2820,N_1923,N_1492);
xnor U2821 (N_2821,N_1357,N_1074);
nor U2822 (N_2822,N_1165,N_879);
or U2823 (N_2823,N_620,N_625);
xor U2824 (N_2824,N_1203,N_1191);
and U2825 (N_2825,N_1402,N_1517);
or U2826 (N_2826,N_662,N_390);
nand U2827 (N_2827,N_1768,N_1089);
or U2828 (N_2828,N_36,N_1682);
and U2829 (N_2829,N_885,N_1798);
nand U2830 (N_2830,N_1960,N_250);
and U2831 (N_2831,N_1664,N_604);
xnor U2832 (N_2832,N_375,N_1924);
xor U2833 (N_2833,N_1578,N_146);
nor U2834 (N_2834,N_1608,N_279);
or U2835 (N_2835,N_1859,N_649);
nand U2836 (N_2836,N_746,N_1560);
or U2837 (N_2837,N_1174,N_370);
or U2838 (N_2838,N_1252,N_1389);
nand U2839 (N_2839,N_1277,N_1887);
nand U2840 (N_2840,N_1904,N_449);
and U2841 (N_2841,N_1312,N_940);
nor U2842 (N_2842,N_63,N_443);
nor U2843 (N_2843,N_1037,N_1006);
and U2844 (N_2844,N_475,N_873);
nand U2845 (N_2845,N_600,N_1358);
xor U2846 (N_2846,N_743,N_1116);
and U2847 (N_2847,N_929,N_425);
or U2848 (N_2848,N_1050,N_155);
and U2849 (N_2849,N_1764,N_1281);
xor U2850 (N_2850,N_878,N_1049);
nor U2851 (N_2851,N_854,N_793);
or U2852 (N_2852,N_1975,N_1378);
or U2853 (N_2853,N_1627,N_1542);
nand U2854 (N_2854,N_1557,N_42);
xnor U2855 (N_2855,N_973,N_1083);
nor U2856 (N_2856,N_830,N_1685);
and U2857 (N_2857,N_1539,N_1016);
xnor U2858 (N_2858,N_1405,N_1628);
xnor U2859 (N_2859,N_535,N_986);
nor U2860 (N_2860,N_497,N_447);
nand U2861 (N_2861,N_578,N_1112);
and U2862 (N_2862,N_1471,N_136);
xnor U2863 (N_2863,N_558,N_701);
nor U2864 (N_2864,N_1698,N_556);
nor U2865 (N_2865,N_1988,N_839);
and U2866 (N_2866,N_239,N_725);
nor U2867 (N_2867,N_783,N_924);
and U2868 (N_2868,N_1149,N_1327);
nand U2869 (N_2869,N_631,N_1470);
nor U2870 (N_2870,N_1851,N_789);
xnor U2871 (N_2871,N_1775,N_919);
or U2872 (N_2872,N_1237,N_1219);
xor U2873 (N_2873,N_464,N_747);
nor U2874 (N_2874,N_984,N_1825);
nand U2875 (N_2875,N_1166,N_1489);
and U2876 (N_2876,N_798,N_1448);
nand U2877 (N_2877,N_733,N_501);
xor U2878 (N_2878,N_1160,N_264);
nor U2879 (N_2879,N_267,N_1540);
or U2880 (N_2880,N_1092,N_331);
xor U2881 (N_2881,N_1797,N_171);
and U2882 (N_2882,N_1051,N_1024);
or U2883 (N_2883,N_184,N_1042);
nor U2884 (N_2884,N_1512,N_597);
nor U2885 (N_2885,N_235,N_92);
nand U2886 (N_2886,N_54,N_1504);
and U2887 (N_2887,N_1984,N_545);
and U2888 (N_2888,N_1717,N_1054);
nand U2889 (N_2889,N_234,N_270);
and U2890 (N_2890,N_326,N_1593);
nor U2891 (N_2891,N_399,N_1282);
nand U2892 (N_2892,N_303,N_59);
nor U2893 (N_2893,N_454,N_1626);
nand U2894 (N_2894,N_385,N_410);
xnor U2895 (N_2895,N_1914,N_1413);
and U2896 (N_2896,N_1216,N_1713);
nand U2897 (N_2897,N_1128,N_1719);
nand U2898 (N_2898,N_1336,N_1030);
and U2899 (N_2899,N_1746,N_1197);
nor U2900 (N_2900,N_510,N_1491);
or U2901 (N_2901,N_490,N_1806);
xor U2902 (N_2902,N_1211,N_1230);
and U2903 (N_2903,N_1920,N_1298);
or U2904 (N_2904,N_1271,N_967);
nand U2905 (N_2905,N_114,N_773);
nand U2906 (N_2906,N_553,N_506);
xnor U2907 (N_2907,N_1222,N_1869);
xor U2908 (N_2908,N_1055,N_633);
nor U2909 (N_2909,N_1059,N_283);
nor U2910 (N_2910,N_1716,N_1094);
and U2911 (N_2911,N_607,N_137);
nand U2912 (N_2912,N_360,N_660);
nand U2913 (N_2913,N_232,N_1161);
nor U2914 (N_2914,N_563,N_719);
and U2915 (N_2915,N_1432,N_998);
or U2916 (N_2916,N_366,N_1240);
nor U2917 (N_2917,N_543,N_782);
or U2918 (N_2918,N_1741,N_1227);
and U2919 (N_2919,N_1516,N_1585);
xor U2920 (N_2920,N_849,N_469);
nor U2921 (N_2921,N_762,N_252);
xnor U2922 (N_2922,N_4,N_24);
and U2923 (N_2923,N_102,N_1961);
nor U2924 (N_2924,N_500,N_905);
and U2925 (N_2925,N_322,N_1123);
xor U2926 (N_2926,N_325,N_1347);
or U2927 (N_2927,N_1264,N_909);
or U2928 (N_2928,N_1383,N_1590);
and U2929 (N_2929,N_1408,N_72);
or U2930 (N_2930,N_329,N_1720);
xnor U2931 (N_2931,N_335,N_1684);
or U2932 (N_2932,N_300,N_1390);
or U2933 (N_2933,N_1210,N_1269);
or U2934 (N_2934,N_1137,N_626);
nand U2935 (N_2935,N_1902,N_241);
or U2936 (N_2936,N_953,N_75);
nand U2937 (N_2937,N_104,N_433);
and U2938 (N_2938,N_792,N_244);
xnor U2939 (N_2939,N_71,N_1004);
or U2940 (N_2940,N_311,N_262);
nand U2941 (N_2941,N_1880,N_346);
xor U2942 (N_2942,N_1409,N_1954);
and U2943 (N_2943,N_949,N_1709);
and U2944 (N_2944,N_838,N_253);
or U2945 (N_2945,N_266,N_87);
xnor U2946 (N_2946,N_98,N_271);
nand U2947 (N_2947,N_427,N_1108);
or U2948 (N_2948,N_296,N_1848);
nand U2949 (N_2949,N_1370,N_1131);
or U2950 (N_2950,N_363,N_1714);
xor U2951 (N_2951,N_1547,N_1870);
nor U2952 (N_2952,N_1420,N_1616);
or U2953 (N_2953,N_1692,N_1040);
and U2954 (N_2954,N_273,N_1335);
xor U2955 (N_2955,N_1670,N_1299);
or U2956 (N_2956,N_50,N_1662);
nor U2957 (N_2957,N_876,N_896);
xnor U2958 (N_2958,N_881,N_801);
nor U2959 (N_2959,N_1026,N_139);
nor U2960 (N_2960,N_1811,N_853);
nand U2961 (N_2961,N_1144,N_1958);
xnor U2962 (N_2962,N_1523,N_918);
nand U2963 (N_2963,N_1296,N_1418);
nand U2964 (N_2964,N_1328,N_807);
and U2965 (N_2965,N_468,N_386);
xnor U2966 (N_2966,N_1897,N_1151);
xnor U2967 (N_2967,N_595,N_353);
nor U2968 (N_2968,N_1127,N_1105);
nor U2969 (N_2969,N_222,N_1524);
or U2970 (N_2970,N_1772,N_531);
nand U2971 (N_2971,N_920,N_1782);
nand U2972 (N_2972,N_1610,N_1310);
xnor U2973 (N_2973,N_1461,N_1646);
and U2974 (N_2974,N_352,N_617);
nand U2975 (N_2975,N_904,N_745);
xnor U2976 (N_2976,N_1097,N_11);
nor U2977 (N_2977,N_869,N_645);
nor U2978 (N_2978,N_1406,N_430);
nand U2979 (N_2979,N_899,N_1164);
and U2980 (N_2980,N_958,N_383);
and U2981 (N_2981,N_767,N_687);
nor U2982 (N_2982,N_1751,N_1446);
and U2983 (N_2983,N_781,N_1883);
xor U2984 (N_2984,N_646,N_1498);
nand U2985 (N_2985,N_225,N_1770);
and U2986 (N_2986,N_106,N_1332);
and U2987 (N_2987,N_1154,N_742);
nand U2988 (N_2988,N_371,N_419);
and U2989 (N_2989,N_540,N_550);
or U2990 (N_2990,N_1066,N_1603);
nand U2991 (N_2991,N_1443,N_405);
nor U2992 (N_2992,N_764,N_730);
and U2993 (N_2993,N_1368,N_1373);
nand U2994 (N_2994,N_939,N_741);
xor U2995 (N_2995,N_739,N_1063);
xor U2996 (N_2996,N_1532,N_1062);
xor U2997 (N_2997,N_1615,N_689);
and U2998 (N_2998,N_1754,N_1384);
and U2999 (N_2999,N_968,N_221);
nor U3000 (N_3000,N_1852,N_614);
xor U3001 (N_3001,N_1334,N_1015);
xnor U3002 (N_3002,N_929,N_1302);
xnor U3003 (N_3003,N_1772,N_1766);
nand U3004 (N_3004,N_1288,N_461);
xor U3005 (N_3005,N_1974,N_725);
nand U3006 (N_3006,N_339,N_1442);
and U3007 (N_3007,N_486,N_1472);
or U3008 (N_3008,N_1477,N_327);
xnor U3009 (N_3009,N_136,N_596);
and U3010 (N_3010,N_1146,N_334);
or U3011 (N_3011,N_86,N_1521);
nand U3012 (N_3012,N_1100,N_1859);
nor U3013 (N_3013,N_1773,N_829);
or U3014 (N_3014,N_1060,N_1902);
or U3015 (N_3015,N_358,N_117);
nor U3016 (N_3016,N_1734,N_77);
or U3017 (N_3017,N_1870,N_1004);
and U3018 (N_3018,N_1552,N_1035);
nor U3019 (N_3019,N_988,N_206);
nand U3020 (N_3020,N_1725,N_147);
or U3021 (N_3021,N_356,N_1892);
nor U3022 (N_3022,N_1740,N_555);
and U3023 (N_3023,N_768,N_698);
xnor U3024 (N_3024,N_430,N_1932);
xor U3025 (N_3025,N_1282,N_1601);
and U3026 (N_3026,N_1058,N_459);
or U3027 (N_3027,N_1004,N_1985);
xor U3028 (N_3028,N_143,N_1464);
or U3029 (N_3029,N_1009,N_1683);
and U3030 (N_3030,N_1835,N_198);
and U3031 (N_3031,N_1412,N_323);
or U3032 (N_3032,N_1613,N_1771);
and U3033 (N_3033,N_955,N_1962);
and U3034 (N_3034,N_1609,N_303);
and U3035 (N_3035,N_692,N_737);
or U3036 (N_3036,N_1432,N_349);
xnor U3037 (N_3037,N_501,N_257);
and U3038 (N_3038,N_451,N_981);
nor U3039 (N_3039,N_528,N_451);
nand U3040 (N_3040,N_703,N_1697);
nor U3041 (N_3041,N_622,N_1998);
xnor U3042 (N_3042,N_91,N_1542);
xnor U3043 (N_3043,N_641,N_1277);
xor U3044 (N_3044,N_1516,N_828);
nor U3045 (N_3045,N_266,N_1046);
and U3046 (N_3046,N_1595,N_605);
or U3047 (N_3047,N_863,N_1977);
xor U3048 (N_3048,N_1282,N_885);
or U3049 (N_3049,N_256,N_939);
or U3050 (N_3050,N_1139,N_1512);
xnor U3051 (N_3051,N_1940,N_1855);
nand U3052 (N_3052,N_998,N_1253);
xor U3053 (N_3053,N_1545,N_963);
or U3054 (N_3054,N_901,N_1004);
xor U3055 (N_3055,N_1897,N_1559);
and U3056 (N_3056,N_481,N_722);
or U3057 (N_3057,N_1594,N_412);
and U3058 (N_3058,N_1926,N_1126);
and U3059 (N_3059,N_750,N_1031);
nand U3060 (N_3060,N_507,N_1220);
or U3061 (N_3061,N_280,N_1992);
and U3062 (N_3062,N_1637,N_174);
or U3063 (N_3063,N_269,N_1411);
or U3064 (N_3064,N_1128,N_1461);
nand U3065 (N_3065,N_330,N_1570);
or U3066 (N_3066,N_1229,N_1814);
or U3067 (N_3067,N_737,N_591);
or U3068 (N_3068,N_1167,N_1653);
and U3069 (N_3069,N_561,N_1921);
or U3070 (N_3070,N_1584,N_1229);
nand U3071 (N_3071,N_1005,N_1924);
nand U3072 (N_3072,N_1192,N_893);
xor U3073 (N_3073,N_162,N_838);
or U3074 (N_3074,N_144,N_746);
xnor U3075 (N_3075,N_1817,N_1313);
nand U3076 (N_3076,N_1863,N_1445);
or U3077 (N_3077,N_255,N_1483);
nand U3078 (N_3078,N_873,N_28);
nand U3079 (N_3079,N_921,N_1996);
or U3080 (N_3080,N_1743,N_1470);
or U3081 (N_3081,N_333,N_997);
nor U3082 (N_3082,N_271,N_1979);
and U3083 (N_3083,N_1313,N_656);
xor U3084 (N_3084,N_208,N_970);
and U3085 (N_3085,N_827,N_900);
or U3086 (N_3086,N_1274,N_404);
nand U3087 (N_3087,N_458,N_957);
xnor U3088 (N_3088,N_1725,N_907);
or U3089 (N_3089,N_262,N_133);
or U3090 (N_3090,N_913,N_443);
xnor U3091 (N_3091,N_1431,N_1770);
and U3092 (N_3092,N_309,N_28);
nand U3093 (N_3093,N_1851,N_1798);
nor U3094 (N_3094,N_662,N_145);
or U3095 (N_3095,N_896,N_657);
and U3096 (N_3096,N_951,N_1411);
or U3097 (N_3097,N_1849,N_1000);
nand U3098 (N_3098,N_1849,N_1171);
nor U3099 (N_3099,N_1824,N_323);
nand U3100 (N_3100,N_329,N_1794);
and U3101 (N_3101,N_781,N_518);
xor U3102 (N_3102,N_289,N_438);
xnor U3103 (N_3103,N_1207,N_17);
xor U3104 (N_3104,N_1447,N_1115);
and U3105 (N_3105,N_485,N_152);
nand U3106 (N_3106,N_1069,N_1202);
xnor U3107 (N_3107,N_605,N_851);
nor U3108 (N_3108,N_1009,N_1931);
or U3109 (N_3109,N_1884,N_1741);
xor U3110 (N_3110,N_1401,N_1822);
and U3111 (N_3111,N_1380,N_1794);
or U3112 (N_3112,N_217,N_1292);
xor U3113 (N_3113,N_1487,N_807);
nand U3114 (N_3114,N_728,N_1417);
xnor U3115 (N_3115,N_663,N_424);
nand U3116 (N_3116,N_246,N_701);
nand U3117 (N_3117,N_982,N_608);
nor U3118 (N_3118,N_1672,N_1382);
or U3119 (N_3119,N_853,N_1826);
xnor U3120 (N_3120,N_1661,N_263);
or U3121 (N_3121,N_921,N_1269);
nor U3122 (N_3122,N_508,N_215);
or U3123 (N_3123,N_186,N_1565);
or U3124 (N_3124,N_868,N_220);
or U3125 (N_3125,N_1063,N_1085);
xor U3126 (N_3126,N_1081,N_1159);
and U3127 (N_3127,N_1058,N_1985);
and U3128 (N_3128,N_1094,N_74);
nor U3129 (N_3129,N_1347,N_1817);
or U3130 (N_3130,N_1128,N_88);
and U3131 (N_3131,N_1007,N_1578);
nor U3132 (N_3132,N_1652,N_524);
or U3133 (N_3133,N_1379,N_1146);
nand U3134 (N_3134,N_1255,N_750);
nor U3135 (N_3135,N_1848,N_1071);
xnor U3136 (N_3136,N_1696,N_706);
and U3137 (N_3137,N_1693,N_449);
xnor U3138 (N_3138,N_1453,N_620);
and U3139 (N_3139,N_747,N_255);
nor U3140 (N_3140,N_854,N_45);
nor U3141 (N_3141,N_1449,N_457);
or U3142 (N_3142,N_266,N_522);
nand U3143 (N_3143,N_1412,N_80);
or U3144 (N_3144,N_1199,N_740);
nor U3145 (N_3145,N_1721,N_201);
and U3146 (N_3146,N_839,N_1447);
nand U3147 (N_3147,N_1950,N_424);
nor U3148 (N_3148,N_223,N_116);
xor U3149 (N_3149,N_1032,N_774);
and U3150 (N_3150,N_392,N_1502);
nand U3151 (N_3151,N_586,N_1497);
nand U3152 (N_3152,N_1467,N_1588);
and U3153 (N_3153,N_1768,N_725);
nand U3154 (N_3154,N_1228,N_1287);
nand U3155 (N_3155,N_1437,N_1804);
nand U3156 (N_3156,N_1731,N_950);
nor U3157 (N_3157,N_1104,N_1614);
nor U3158 (N_3158,N_1750,N_1055);
nand U3159 (N_3159,N_101,N_773);
nor U3160 (N_3160,N_676,N_442);
and U3161 (N_3161,N_372,N_860);
nor U3162 (N_3162,N_1729,N_733);
nor U3163 (N_3163,N_119,N_1612);
or U3164 (N_3164,N_101,N_1486);
nand U3165 (N_3165,N_684,N_551);
nand U3166 (N_3166,N_446,N_555);
or U3167 (N_3167,N_198,N_1895);
xor U3168 (N_3168,N_1850,N_1412);
and U3169 (N_3169,N_975,N_1717);
or U3170 (N_3170,N_241,N_1451);
xnor U3171 (N_3171,N_1897,N_1808);
or U3172 (N_3172,N_784,N_523);
nor U3173 (N_3173,N_114,N_1557);
nand U3174 (N_3174,N_663,N_988);
xor U3175 (N_3175,N_1576,N_874);
and U3176 (N_3176,N_633,N_1898);
and U3177 (N_3177,N_1814,N_483);
or U3178 (N_3178,N_111,N_1621);
nand U3179 (N_3179,N_1842,N_1503);
and U3180 (N_3180,N_984,N_1087);
nor U3181 (N_3181,N_1771,N_1348);
and U3182 (N_3182,N_786,N_146);
xor U3183 (N_3183,N_293,N_1162);
and U3184 (N_3184,N_671,N_434);
nand U3185 (N_3185,N_936,N_52);
nand U3186 (N_3186,N_1218,N_1691);
nor U3187 (N_3187,N_1503,N_1670);
nand U3188 (N_3188,N_69,N_282);
or U3189 (N_3189,N_1355,N_1764);
nor U3190 (N_3190,N_112,N_1992);
or U3191 (N_3191,N_1551,N_1891);
and U3192 (N_3192,N_1326,N_1167);
xor U3193 (N_3193,N_1337,N_1858);
and U3194 (N_3194,N_342,N_1171);
nor U3195 (N_3195,N_348,N_750);
nand U3196 (N_3196,N_1131,N_851);
and U3197 (N_3197,N_786,N_851);
and U3198 (N_3198,N_1492,N_1484);
nand U3199 (N_3199,N_1153,N_532);
xor U3200 (N_3200,N_578,N_20);
nor U3201 (N_3201,N_464,N_976);
xor U3202 (N_3202,N_737,N_1104);
xnor U3203 (N_3203,N_959,N_101);
and U3204 (N_3204,N_1324,N_1744);
nor U3205 (N_3205,N_1035,N_985);
or U3206 (N_3206,N_1947,N_1633);
or U3207 (N_3207,N_47,N_1390);
and U3208 (N_3208,N_608,N_1889);
nor U3209 (N_3209,N_682,N_975);
or U3210 (N_3210,N_1316,N_280);
xor U3211 (N_3211,N_1144,N_1908);
nand U3212 (N_3212,N_340,N_437);
nand U3213 (N_3213,N_1685,N_1275);
and U3214 (N_3214,N_269,N_1036);
nand U3215 (N_3215,N_83,N_1702);
or U3216 (N_3216,N_1824,N_1160);
and U3217 (N_3217,N_1654,N_1549);
xor U3218 (N_3218,N_160,N_979);
or U3219 (N_3219,N_1410,N_1937);
xor U3220 (N_3220,N_242,N_149);
nor U3221 (N_3221,N_629,N_1206);
nand U3222 (N_3222,N_1720,N_1902);
nand U3223 (N_3223,N_670,N_1135);
and U3224 (N_3224,N_1827,N_1006);
xor U3225 (N_3225,N_1880,N_228);
nor U3226 (N_3226,N_1661,N_716);
nand U3227 (N_3227,N_429,N_964);
nand U3228 (N_3228,N_1248,N_1520);
nor U3229 (N_3229,N_299,N_1891);
nand U3230 (N_3230,N_72,N_1090);
and U3231 (N_3231,N_1812,N_1777);
nor U3232 (N_3232,N_672,N_1337);
xor U3233 (N_3233,N_736,N_1680);
xnor U3234 (N_3234,N_30,N_1896);
xor U3235 (N_3235,N_21,N_1421);
nor U3236 (N_3236,N_1649,N_1193);
and U3237 (N_3237,N_1984,N_616);
xor U3238 (N_3238,N_1724,N_394);
xnor U3239 (N_3239,N_611,N_597);
nor U3240 (N_3240,N_1412,N_154);
xor U3241 (N_3241,N_864,N_1100);
nand U3242 (N_3242,N_632,N_42);
nand U3243 (N_3243,N_392,N_327);
nor U3244 (N_3244,N_874,N_1508);
nand U3245 (N_3245,N_1477,N_401);
nand U3246 (N_3246,N_841,N_697);
and U3247 (N_3247,N_287,N_582);
xnor U3248 (N_3248,N_215,N_1821);
or U3249 (N_3249,N_1452,N_901);
nor U3250 (N_3250,N_557,N_101);
or U3251 (N_3251,N_365,N_1383);
or U3252 (N_3252,N_1376,N_1940);
and U3253 (N_3253,N_1276,N_69);
and U3254 (N_3254,N_1270,N_944);
and U3255 (N_3255,N_616,N_783);
nand U3256 (N_3256,N_400,N_1793);
and U3257 (N_3257,N_611,N_184);
nand U3258 (N_3258,N_1852,N_1265);
nor U3259 (N_3259,N_317,N_1614);
and U3260 (N_3260,N_685,N_964);
nor U3261 (N_3261,N_1931,N_571);
or U3262 (N_3262,N_1348,N_508);
or U3263 (N_3263,N_1193,N_527);
nor U3264 (N_3264,N_863,N_1991);
nor U3265 (N_3265,N_461,N_360);
xnor U3266 (N_3266,N_401,N_1755);
or U3267 (N_3267,N_167,N_1724);
and U3268 (N_3268,N_1585,N_925);
xnor U3269 (N_3269,N_98,N_1420);
nor U3270 (N_3270,N_713,N_203);
xnor U3271 (N_3271,N_1536,N_64);
and U3272 (N_3272,N_1978,N_1655);
nand U3273 (N_3273,N_97,N_209);
or U3274 (N_3274,N_750,N_968);
and U3275 (N_3275,N_874,N_1319);
xor U3276 (N_3276,N_464,N_1056);
or U3277 (N_3277,N_1193,N_342);
nand U3278 (N_3278,N_1302,N_1779);
and U3279 (N_3279,N_1724,N_668);
xnor U3280 (N_3280,N_812,N_1440);
nand U3281 (N_3281,N_600,N_1472);
nand U3282 (N_3282,N_1367,N_350);
xnor U3283 (N_3283,N_212,N_910);
nand U3284 (N_3284,N_457,N_1866);
or U3285 (N_3285,N_677,N_1952);
nor U3286 (N_3286,N_1477,N_284);
and U3287 (N_3287,N_1713,N_861);
xnor U3288 (N_3288,N_827,N_402);
and U3289 (N_3289,N_141,N_510);
nand U3290 (N_3290,N_288,N_490);
nor U3291 (N_3291,N_478,N_414);
xor U3292 (N_3292,N_1250,N_1391);
or U3293 (N_3293,N_652,N_1392);
and U3294 (N_3294,N_423,N_47);
nor U3295 (N_3295,N_256,N_664);
nor U3296 (N_3296,N_976,N_1220);
xor U3297 (N_3297,N_1552,N_825);
nand U3298 (N_3298,N_86,N_1084);
nor U3299 (N_3299,N_875,N_900);
or U3300 (N_3300,N_565,N_1440);
xnor U3301 (N_3301,N_1383,N_1896);
xnor U3302 (N_3302,N_488,N_427);
nand U3303 (N_3303,N_1911,N_881);
nor U3304 (N_3304,N_807,N_650);
and U3305 (N_3305,N_1239,N_70);
nor U3306 (N_3306,N_1081,N_1801);
and U3307 (N_3307,N_1833,N_678);
nor U3308 (N_3308,N_1253,N_655);
or U3309 (N_3309,N_531,N_1953);
nand U3310 (N_3310,N_1124,N_1728);
nor U3311 (N_3311,N_748,N_161);
nand U3312 (N_3312,N_1925,N_1914);
xor U3313 (N_3313,N_134,N_1554);
or U3314 (N_3314,N_1524,N_32);
xor U3315 (N_3315,N_489,N_1971);
nand U3316 (N_3316,N_1885,N_291);
nor U3317 (N_3317,N_639,N_182);
and U3318 (N_3318,N_568,N_441);
xor U3319 (N_3319,N_35,N_1131);
and U3320 (N_3320,N_338,N_1750);
and U3321 (N_3321,N_639,N_288);
and U3322 (N_3322,N_72,N_1776);
xnor U3323 (N_3323,N_1743,N_1851);
or U3324 (N_3324,N_656,N_887);
nand U3325 (N_3325,N_1762,N_1460);
xnor U3326 (N_3326,N_1213,N_670);
or U3327 (N_3327,N_298,N_202);
nand U3328 (N_3328,N_1372,N_1805);
nand U3329 (N_3329,N_708,N_501);
or U3330 (N_3330,N_770,N_613);
or U3331 (N_3331,N_1982,N_292);
and U3332 (N_3332,N_843,N_108);
and U3333 (N_3333,N_370,N_1284);
xnor U3334 (N_3334,N_687,N_817);
nand U3335 (N_3335,N_123,N_206);
nand U3336 (N_3336,N_761,N_920);
xnor U3337 (N_3337,N_1696,N_769);
and U3338 (N_3338,N_435,N_1119);
nand U3339 (N_3339,N_1896,N_146);
nor U3340 (N_3340,N_902,N_1511);
nand U3341 (N_3341,N_1785,N_1924);
or U3342 (N_3342,N_549,N_1025);
nor U3343 (N_3343,N_957,N_554);
nand U3344 (N_3344,N_839,N_124);
nand U3345 (N_3345,N_1677,N_401);
and U3346 (N_3346,N_1651,N_878);
or U3347 (N_3347,N_26,N_897);
nor U3348 (N_3348,N_1578,N_1085);
and U3349 (N_3349,N_159,N_1474);
xnor U3350 (N_3350,N_746,N_855);
nand U3351 (N_3351,N_234,N_874);
or U3352 (N_3352,N_1445,N_477);
xnor U3353 (N_3353,N_1576,N_1358);
and U3354 (N_3354,N_1227,N_1180);
or U3355 (N_3355,N_879,N_614);
nand U3356 (N_3356,N_1793,N_1079);
and U3357 (N_3357,N_616,N_1873);
and U3358 (N_3358,N_133,N_362);
xor U3359 (N_3359,N_745,N_1336);
nand U3360 (N_3360,N_1290,N_1985);
and U3361 (N_3361,N_757,N_18);
xor U3362 (N_3362,N_1055,N_1006);
and U3363 (N_3363,N_737,N_1730);
and U3364 (N_3364,N_200,N_1757);
nand U3365 (N_3365,N_1869,N_655);
nor U3366 (N_3366,N_1653,N_802);
or U3367 (N_3367,N_1310,N_1820);
nand U3368 (N_3368,N_249,N_942);
nand U3369 (N_3369,N_1610,N_1734);
or U3370 (N_3370,N_226,N_769);
nand U3371 (N_3371,N_1441,N_1364);
and U3372 (N_3372,N_815,N_737);
or U3373 (N_3373,N_219,N_101);
nor U3374 (N_3374,N_1041,N_1654);
nand U3375 (N_3375,N_1963,N_151);
nand U3376 (N_3376,N_931,N_386);
nor U3377 (N_3377,N_1288,N_27);
xor U3378 (N_3378,N_1871,N_770);
or U3379 (N_3379,N_1371,N_1649);
xnor U3380 (N_3380,N_141,N_1774);
or U3381 (N_3381,N_783,N_152);
nor U3382 (N_3382,N_62,N_1526);
and U3383 (N_3383,N_12,N_924);
and U3384 (N_3384,N_1095,N_1479);
or U3385 (N_3385,N_242,N_389);
nand U3386 (N_3386,N_1720,N_1854);
nor U3387 (N_3387,N_1187,N_1872);
xnor U3388 (N_3388,N_372,N_906);
nor U3389 (N_3389,N_1584,N_322);
or U3390 (N_3390,N_1301,N_1379);
and U3391 (N_3391,N_1352,N_1699);
xnor U3392 (N_3392,N_1255,N_1266);
or U3393 (N_3393,N_37,N_644);
nand U3394 (N_3394,N_1038,N_1877);
and U3395 (N_3395,N_193,N_342);
nor U3396 (N_3396,N_577,N_762);
nor U3397 (N_3397,N_290,N_1011);
or U3398 (N_3398,N_153,N_805);
xnor U3399 (N_3399,N_418,N_1351);
nor U3400 (N_3400,N_36,N_1310);
nand U3401 (N_3401,N_509,N_216);
nor U3402 (N_3402,N_128,N_1042);
nor U3403 (N_3403,N_1074,N_1569);
or U3404 (N_3404,N_299,N_702);
nor U3405 (N_3405,N_1715,N_1153);
or U3406 (N_3406,N_892,N_187);
nor U3407 (N_3407,N_749,N_437);
nand U3408 (N_3408,N_791,N_948);
nor U3409 (N_3409,N_1805,N_1099);
and U3410 (N_3410,N_909,N_604);
xnor U3411 (N_3411,N_969,N_473);
xor U3412 (N_3412,N_1773,N_52);
nor U3413 (N_3413,N_527,N_434);
xor U3414 (N_3414,N_21,N_1678);
xor U3415 (N_3415,N_924,N_1734);
and U3416 (N_3416,N_371,N_1118);
nor U3417 (N_3417,N_698,N_1552);
nor U3418 (N_3418,N_1221,N_733);
or U3419 (N_3419,N_1702,N_426);
and U3420 (N_3420,N_1031,N_834);
and U3421 (N_3421,N_1244,N_909);
xor U3422 (N_3422,N_570,N_575);
nor U3423 (N_3423,N_741,N_971);
xnor U3424 (N_3424,N_920,N_1756);
nor U3425 (N_3425,N_938,N_745);
nor U3426 (N_3426,N_1612,N_716);
nor U3427 (N_3427,N_1600,N_1266);
xnor U3428 (N_3428,N_1478,N_1200);
nor U3429 (N_3429,N_1828,N_1351);
and U3430 (N_3430,N_113,N_403);
and U3431 (N_3431,N_1447,N_733);
or U3432 (N_3432,N_740,N_455);
xnor U3433 (N_3433,N_106,N_1158);
xor U3434 (N_3434,N_1297,N_336);
xor U3435 (N_3435,N_1314,N_1858);
xor U3436 (N_3436,N_1442,N_504);
or U3437 (N_3437,N_97,N_277);
nand U3438 (N_3438,N_534,N_622);
nand U3439 (N_3439,N_1628,N_351);
and U3440 (N_3440,N_1720,N_554);
xnor U3441 (N_3441,N_669,N_156);
or U3442 (N_3442,N_359,N_1197);
nand U3443 (N_3443,N_558,N_1607);
nand U3444 (N_3444,N_237,N_329);
xnor U3445 (N_3445,N_1783,N_1126);
xor U3446 (N_3446,N_637,N_1316);
nor U3447 (N_3447,N_99,N_1411);
or U3448 (N_3448,N_165,N_1933);
or U3449 (N_3449,N_394,N_1191);
or U3450 (N_3450,N_1913,N_1411);
or U3451 (N_3451,N_833,N_677);
nand U3452 (N_3452,N_1676,N_1325);
nor U3453 (N_3453,N_242,N_787);
nor U3454 (N_3454,N_1128,N_1746);
nor U3455 (N_3455,N_475,N_1277);
nand U3456 (N_3456,N_507,N_1168);
nand U3457 (N_3457,N_947,N_1393);
xor U3458 (N_3458,N_213,N_1188);
nand U3459 (N_3459,N_1577,N_869);
xor U3460 (N_3460,N_346,N_1105);
xor U3461 (N_3461,N_1301,N_154);
nor U3462 (N_3462,N_593,N_1203);
xor U3463 (N_3463,N_153,N_1986);
or U3464 (N_3464,N_1738,N_1228);
xor U3465 (N_3465,N_769,N_1695);
xor U3466 (N_3466,N_1015,N_1696);
or U3467 (N_3467,N_1900,N_1754);
nor U3468 (N_3468,N_1516,N_689);
xor U3469 (N_3469,N_1325,N_1307);
xnor U3470 (N_3470,N_1958,N_1946);
nand U3471 (N_3471,N_508,N_97);
xor U3472 (N_3472,N_1972,N_247);
xor U3473 (N_3473,N_1357,N_508);
nand U3474 (N_3474,N_1858,N_1370);
and U3475 (N_3475,N_412,N_1953);
nor U3476 (N_3476,N_1829,N_1923);
nand U3477 (N_3477,N_1777,N_1624);
and U3478 (N_3478,N_1502,N_572);
or U3479 (N_3479,N_1037,N_302);
nand U3480 (N_3480,N_1585,N_1452);
nor U3481 (N_3481,N_432,N_1426);
xnor U3482 (N_3482,N_405,N_1477);
nand U3483 (N_3483,N_715,N_967);
xor U3484 (N_3484,N_1759,N_1748);
nand U3485 (N_3485,N_1905,N_1060);
and U3486 (N_3486,N_12,N_382);
or U3487 (N_3487,N_1494,N_688);
nor U3488 (N_3488,N_51,N_32);
and U3489 (N_3489,N_598,N_728);
xnor U3490 (N_3490,N_1698,N_203);
nand U3491 (N_3491,N_1812,N_1559);
nor U3492 (N_3492,N_156,N_1487);
nand U3493 (N_3493,N_198,N_1588);
nor U3494 (N_3494,N_960,N_1110);
or U3495 (N_3495,N_122,N_842);
and U3496 (N_3496,N_75,N_1243);
and U3497 (N_3497,N_1903,N_895);
nand U3498 (N_3498,N_1588,N_1820);
xor U3499 (N_3499,N_785,N_1512);
and U3500 (N_3500,N_949,N_1239);
or U3501 (N_3501,N_1182,N_213);
xor U3502 (N_3502,N_1639,N_1476);
or U3503 (N_3503,N_1852,N_1860);
nor U3504 (N_3504,N_1821,N_1359);
xor U3505 (N_3505,N_300,N_646);
and U3506 (N_3506,N_220,N_349);
nor U3507 (N_3507,N_1831,N_1531);
nand U3508 (N_3508,N_1188,N_882);
nand U3509 (N_3509,N_776,N_981);
nand U3510 (N_3510,N_1637,N_1229);
and U3511 (N_3511,N_269,N_1703);
nor U3512 (N_3512,N_738,N_1513);
nor U3513 (N_3513,N_890,N_1536);
or U3514 (N_3514,N_890,N_1307);
or U3515 (N_3515,N_505,N_1619);
or U3516 (N_3516,N_1547,N_1658);
nor U3517 (N_3517,N_445,N_1998);
nand U3518 (N_3518,N_1084,N_45);
nand U3519 (N_3519,N_696,N_981);
nand U3520 (N_3520,N_1332,N_1802);
or U3521 (N_3521,N_42,N_1680);
nor U3522 (N_3522,N_1166,N_1009);
nand U3523 (N_3523,N_949,N_191);
and U3524 (N_3524,N_842,N_1120);
nand U3525 (N_3525,N_605,N_612);
and U3526 (N_3526,N_1706,N_302);
nand U3527 (N_3527,N_1182,N_435);
nor U3528 (N_3528,N_1062,N_840);
nor U3529 (N_3529,N_1125,N_1233);
or U3530 (N_3530,N_1340,N_1857);
and U3531 (N_3531,N_1603,N_1288);
or U3532 (N_3532,N_685,N_325);
nor U3533 (N_3533,N_1070,N_414);
nand U3534 (N_3534,N_1915,N_1648);
and U3535 (N_3535,N_1004,N_323);
nor U3536 (N_3536,N_1861,N_331);
xor U3537 (N_3537,N_430,N_1049);
and U3538 (N_3538,N_1361,N_63);
nor U3539 (N_3539,N_982,N_1529);
or U3540 (N_3540,N_991,N_372);
or U3541 (N_3541,N_895,N_1587);
and U3542 (N_3542,N_1384,N_15);
xnor U3543 (N_3543,N_719,N_1602);
and U3544 (N_3544,N_681,N_774);
or U3545 (N_3545,N_984,N_1782);
or U3546 (N_3546,N_822,N_937);
nor U3547 (N_3547,N_574,N_488);
nand U3548 (N_3548,N_1555,N_605);
nand U3549 (N_3549,N_1319,N_1158);
or U3550 (N_3550,N_102,N_1329);
nand U3551 (N_3551,N_1194,N_934);
nor U3552 (N_3552,N_1471,N_1468);
or U3553 (N_3553,N_781,N_81);
nor U3554 (N_3554,N_1642,N_932);
nor U3555 (N_3555,N_1124,N_613);
xor U3556 (N_3556,N_977,N_1862);
nor U3557 (N_3557,N_1735,N_843);
or U3558 (N_3558,N_1066,N_1280);
nand U3559 (N_3559,N_407,N_1331);
or U3560 (N_3560,N_1803,N_1697);
nor U3561 (N_3561,N_444,N_926);
and U3562 (N_3562,N_703,N_150);
or U3563 (N_3563,N_1244,N_1054);
xor U3564 (N_3564,N_1293,N_1377);
nor U3565 (N_3565,N_315,N_1984);
or U3566 (N_3566,N_816,N_798);
nand U3567 (N_3567,N_254,N_1427);
or U3568 (N_3568,N_980,N_1941);
and U3569 (N_3569,N_1219,N_1838);
nand U3570 (N_3570,N_1131,N_1069);
and U3571 (N_3571,N_762,N_553);
or U3572 (N_3572,N_9,N_492);
and U3573 (N_3573,N_1522,N_1471);
and U3574 (N_3574,N_899,N_1228);
or U3575 (N_3575,N_1454,N_630);
and U3576 (N_3576,N_1427,N_1961);
or U3577 (N_3577,N_961,N_1891);
and U3578 (N_3578,N_1954,N_1010);
xor U3579 (N_3579,N_1529,N_1316);
or U3580 (N_3580,N_369,N_1714);
nor U3581 (N_3581,N_1074,N_1124);
nand U3582 (N_3582,N_1505,N_1608);
nor U3583 (N_3583,N_43,N_1723);
and U3584 (N_3584,N_559,N_520);
xnor U3585 (N_3585,N_960,N_594);
xor U3586 (N_3586,N_1374,N_1378);
nand U3587 (N_3587,N_866,N_1946);
nor U3588 (N_3588,N_1958,N_823);
xor U3589 (N_3589,N_1236,N_386);
and U3590 (N_3590,N_195,N_1151);
xor U3591 (N_3591,N_671,N_1260);
xnor U3592 (N_3592,N_1148,N_865);
nor U3593 (N_3593,N_622,N_605);
nand U3594 (N_3594,N_597,N_1348);
and U3595 (N_3595,N_1418,N_84);
or U3596 (N_3596,N_1911,N_83);
xor U3597 (N_3597,N_1300,N_1413);
nand U3598 (N_3598,N_931,N_1564);
and U3599 (N_3599,N_363,N_274);
and U3600 (N_3600,N_752,N_544);
or U3601 (N_3601,N_1979,N_81);
nand U3602 (N_3602,N_489,N_1320);
nand U3603 (N_3603,N_986,N_748);
nor U3604 (N_3604,N_1487,N_1642);
nor U3605 (N_3605,N_1060,N_49);
nor U3606 (N_3606,N_921,N_1163);
nor U3607 (N_3607,N_1307,N_685);
nor U3608 (N_3608,N_1686,N_1704);
xor U3609 (N_3609,N_724,N_1170);
and U3610 (N_3610,N_563,N_763);
nor U3611 (N_3611,N_156,N_434);
or U3612 (N_3612,N_1196,N_1787);
xor U3613 (N_3613,N_1322,N_1371);
or U3614 (N_3614,N_216,N_1277);
nor U3615 (N_3615,N_1068,N_205);
nor U3616 (N_3616,N_80,N_229);
nor U3617 (N_3617,N_1577,N_243);
nand U3618 (N_3618,N_1880,N_1192);
or U3619 (N_3619,N_347,N_677);
nand U3620 (N_3620,N_949,N_311);
nor U3621 (N_3621,N_170,N_335);
and U3622 (N_3622,N_1737,N_1146);
or U3623 (N_3623,N_346,N_523);
and U3624 (N_3624,N_259,N_492);
nor U3625 (N_3625,N_402,N_1598);
nand U3626 (N_3626,N_1906,N_1837);
or U3627 (N_3627,N_821,N_1713);
and U3628 (N_3628,N_422,N_1181);
nand U3629 (N_3629,N_1465,N_1038);
nor U3630 (N_3630,N_0,N_1547);
xnor U3631 (N_3631,N_1891,N_479);
nand U3632 (N_3632,N_547,N_498);
xor U3633 (N_3633,N_1569,N_1052);
or U3634 (N_3634,N_1828,N_1461);
xnor U3635 (N_3635,N_645,N_630);
and U3636 (N_3636,N_334,N_537);
and U3637 (N_3637,N_1769,N_233);
nand U3638 (N_3638,N_381,N_765);
and U3639 (N_3639,N_1463,N_1715);
or U3640 (N_3640,N_1447,N_823);
nor U3641 (N_3641,N_1075,N_1925);
nand U3642 (N_3642,N_262,N_397);
nor U3643 (N_3643,N_494,N_1017);
or U3644 (N_3644,N_1664,N_798);
xor U3645 (N_3645,N_1827,N_490);
and U3646 (N_3646,N_1504,N_729);
and U3647 (N_3647,N_69,N_126);
nor U3648 (N_3648,N_832,N_753);
and U3649 (N_3649,N_1398,N_1790);
or U3650 (N_3650,N_649,N_379);
or U3651 (N_3651,N_7,N_780);
and U3652 (N_3652,N_1947,N_1139);
or U3653 (N_3653,N_658,N_374);
and U3654 (N_3654,N_131,N_1674);
xnor U3655 (N_3655,N_871,N_1924);
or U3656 (N_3656,N_796,N_280);
xnor U3657 (N_3657,N_1775,N_2);
and U3658 (N_3658,N_824,N_671);
or U3659 (N_3659,N_1188,N_1208);
or U3660 (N_3660,N_1686,N_1619);
nor U3661 (N_3661,N_325,N_96);
nand U3662 (N_3662,N_531,N_181);
and U3663 (N_3663,N_126,N_1152);
and U3664 (N_3664,N_720,N_690);
or U3665 (N_3665,N_1681,N_944);
xor U3666 (N_3666,N_174,N_1849);
xor U3667 (N_3667,N_255,N_593);
nor U3668 (N_3668,N_1579,N_269);
or U3669 (N_3669,N_837,N_1852);
or U3670 (N_3670,N_1940,N_1021);
and U3671 (N_3671,N_473,N_573);
xor U3672 (N_3672,N_1612,N_330);
nor U3673 (N_3673,N_1874,N_923);
nor U3674 (N_3674,N_1227,N_1104);
nor U3675 (N_3675,N_1919,N_614);
nand U3676 (N_3676,N_2,N_1553);
and U3677 (N_3677,N_1504,N_1506);
nor U3678 (N_3678,N_1502,N_912);
nand U3679 (N_3679,N_1618,N_808);
xor U3680 (N_3680,N_62,N_1112);
or U3681 (N_3681,N_84,N_996);
and U3682 (N_3682,N_256,N_1951);
nand U3683 (N_3683,N_91,N_1116);
and U3684 (N_3684,N_58,N_1844);
nor U3685 (N_3685,N_114,N_546);
xnor U3686 (N_3686,N_1948,N_792);
nand U3687 (N_3687,N_50,N_696);
nor U3688 (N_3688,N_110,N_759);
and U3689 (N_3689,N_1019,N_1568);
xor U3690 (N_3690,N_591,N_729);
nor U3691 (N_3691,N_942,N_1925);
xor U3692 (N_3692,N_513,N_814);
nand U3693 (N_3693,N_1178,N_522);
nand U3694 (N_3694,N_171,N_1354);
and U3695 (N_3695,N_1906,N_1643);
xor U3696 (N_3696,N_961,N_1272);
and U3697 (N_3697,N_1193,N_44);
nor U3698 (N_3698,N_1145,N_627);
and U3699 (N_3699,N_1241,N_1841);
or U3700 (N_3700,N_731,N_363);
nand U3701 (N_3701,N_1504,N_489);
nand U3702 (N_3702,N_429,N_1670);
nor U3703 (N_3703,N_1007,N_347);
nand U3704 (N_3704,N_1110,N_878);
xnor U3705 (N_3705,N_463,N_1300);
nand U3706 (N_3706,N_1128,N_1883);
or U3707 (N_3707,N_108,N_1944);
or U3708 (N_3708,N_207,N_177);
xnor U3709 (N_3709,N_451,N_544);
xnor U3710 (N_3710,N_733,N_482);
nor U3711 (N_3711,N_1882,N_1206);
nor U3712 (N_3712,N_1032,N_1445);
and U3713 (N_3713,N_368,N_1021);
and U3714 (N_3714,N_730,N_439);
or U3715 (N_3715,N_1720,N_238);
or U3716 (N_3716,N_1448,N_1883);
and U3717 (N_3717,N_1134,N_1421);
and U3718 (N_3718,N_617,N_1763);
nand U3719 (N_3719,N_461,N_948);
or U3720 (N_3720,N_1890,N_1439);
nor U3721 (N_3721,N_269,N_1269);
or U3722 (N_3722,N_1868,N_847);
nand U3723 (N_3723,N_1769,N_930);
or U3724 (N_3724,N_683,N_1921);
nand U3725 (N_3725,N_1915,N_1273);
nand U3726 (N_3726,N_1022,N_411);
nand U3727 (N_3727,N_102,N_1669);
nand U3728 (N_3728,N_1300,N_1097);
xnor U3729 (N_3729,N_602,N_1040);
or U3730 (N_3730,N_1647,N_529);
and U3731 (N_3731,N_757,N_524);
or U3732 (N_3732,N_631,N_1608);
xnor U3733 (N_3733,N_372,N_1297);
xnor U3734 (N_3734,N_1686,N_1965);
xor U3735 (N_3735,N_1082,N_1383);
and U3736 (N_3736,N_1552,N_1995);
and U3737 (N_3737,N_1506,N_1027);
nand U3738 (N_3738,N_1821,N_1952);
and U3739 (N_3739,N_1697,N_679);
nor U3740 (N_3740,N_1733,N_115);
xor U3741 (N_3741,N_601,N_1960);
and U3742 (N_3742,N_889,N_984);
nor U3743 (N_3743,N_1630,N_1403);
nand U3744 (N_3744,N_1881,N_1711);
or U3745 (N_3745,N_463,N_932);
nand U3746 (N_3746,N_1303,N_56);
nand U3747 (N_3747,N_211,N_894);
nor U3748 (N_3748,N_615,N_221);
nor U3749 (N_3749,N_405,N_1939);
nor U3750 (N_3750,N_344,N_1699);
nor U3751 (N_3751,N_18,N_161);
and U3752 (N_3752,N_403,N_1178);
nor U3753 (N_3753,N_829,N_260);
and U3754 (N_3754,N_755,N_1397);
xnor U3755 (N_3755,N_771,N_1086);
nand U3756 (N_3756,N_1737,N_1148);
nor U3757 (N_3757,N_1084,N_1055);
xnor U3758 (N_3758,N_326,N_1378);
nand U3759 (N_3759,N_1354,N_1673);
and U3760 (N_3760,N_1395,N_267);
nor U3761 (N_3761,N_1993,N_175);
and U3762 (N_3762,N_757,N_1306);
nand U3763 (N_3763,N_339,N_182);
xor U3764 (N_3764,N_867,N_1673);
or U3765 (N_3765,N_446,N_1913);
or U3766 (N_3766,N_1207,N_1717);
nand U3767 (N_3767,N_739,N_537);
or U3768 (N_3768,N_1727,N_183);
nor U3769 (N_3769,N_8,N_828);
xnor U3770 (N_3770,N_948,N_156);
and U3771 (N_3771,N_616,N_762);
xnor U3772 (N_3772,N_1956,N_845);
nand U3773 (N_3773,N_563,N_470);
nand U3774 (N_3774,N_700,N_547);
nor U3775 (N_3775,N_686,N_302);
xor U3776 (N_3776,N_1372,N_369);
nor U3777 (N_3777,N_1938,N_1900);
nand U3778 (N_3778,N_1347,N_95);
nor U3779 (N_3779,N_27,N_325);
nor U3780 (N_3780,N_332,N_608);
or U3781 (N_3781,N_1588,N_1500);
and U3782 (N_3782,N_637,N_1501);
xor U3783 (N_3783,N_1411,N_873);
nor U3784 (N_3784,N_783,N_53);
nor U3785 (N_3785,N_1715,N_1467);
nand U3786 (N_3786,N_1876,N_564);
and U3787 (N_3787,N_1899,N_1492);
xor U3788 (N_3788,N_1917,N_1836);
or U3789 (N_3789,N_359,N_783);
nand U3790 (N_3790,N_1844,N_1377);
and U3791 (N_3791,N_1267,N_1809);
xor U3792 (N_3792,N_845,N_503);
nand U3793 (N_3793,N_1903,N_1078);
nand U3794 (N_3794,N_1509,N_1106);
and U3795 (N_3795,N_483,N_766);
or U3796 (N_3796,N_1421,N_769);
and U3797 (N_3797,N_1494,N_946);
nand U3798 (N_3798,N_793,N_1275);
xor U3799 (N_3799,N_138,N_1111);
xnor U3800 (N_3800,N_1727,N_430);
or U3801 (N_3801,N_1474,N_582);
xnor U3802 (N_3802,N_738,N_198);
nor U3803 (N_3803,N_1722,N_1868);
nand U3804 (N_3804,N_1796,N_1261);
or U3805 (N_3805,N_760,N_1517);
xnor U3806 (N_3806,N_727,N_781);
or U3807 (N_3807,N_774,N_852);
xor U3808 (N_3808,N_854,N_1704);
or U3809 (N_3809,N_116,N_815);
and U3810 (N_3810,N_546,N_423);
and U3811 (N_3811,N_1826,N_1799);
and U3812 (N_3812,N_1972,N_61);
or U3813 (N_3813,N_220,N_889);
or U3814 (N_3814,N_1640,N_1220);
or U3815 (N_3815,N_187,N_353);
nor U3816 (N_3816,N_1134,N_583);
nand U3817 (N_3817,N_235,N_1048);
nand U3818 (N_3818,N_1880,N_1077);
or U3819 (N_3819,N_1482,N_1654);
xnor U3820 (N_3820,N_98,N_970);
xnor U3821 (N_3821,N_1655,N_1692);
nor U3822 (N_3822,N_68,N_1595);
xnor U3823 (N_3823,N_1485,N_887);
or U3824 (N_3824,N_340,N_1185);
or U3825 (N_3825,N_147,N_616);
nor U3826 (N_3826,N_1513,N_832);
or U3827 (N_3827,N_148,N_1073);
nor U3828 (N_3828,N_1655,N_563);
nor U3829 (N_3829,N_1252,N_1044);
and U3830 (N_3830,N_836,N_1283);
or U3831 (N_3831,N_195,N_736);
or U3832 (N_3832,N_674,N_1736);
or U3833 (N_3833,N_784,N_1113);
xor U3834 (N_3834,N_1988,N_1831);
xnor U3835 (N_3835,N_503,N_943);
nand U3836 (N_3836,N_1244,N_656);
or U3837 (N_3837,N_1983,N_1997);
nor U3838 (N_3838,N_1817,N_120);
nor U3839 (N_3839,N_726,N_866);
nand U3840 (N_3840,N_869,N_844);
or U3841 (N_3841,N_1366,N_1604);
nand U3842 (N_3842,N_610,N_1908);
or U3843 (N_3843,N_1859,N_646);
xor U3844 (N_3844,N_1140,N_1731);
and U3845 (N_3845,N_1458,N_327);
nand U3846 (N_3846,N_687,N_1216);
and U3847 (N_3847,N_106,N_1452);
nor U3848 (N_3848,N_1572,N_630);
and U3849 (N_3849,N_1579,N_760);
nand U3850 (N_3850,N_77,N_1204);
and U3851 (N_3851,N_1696,N_1312);
nor U3852 (N_3852,N_1021,N_1581);
nor U3853 (N_3853,N_1038,N_826);
and U3854 (N_3854,N_391,N_1650);
nor U3855 (N_3855,N_314,N_1663);
nand U3856 (N_3856,N_1724,N_1747);
or U3857 (N_3857,N_331,N_261);
nor U3858 (N_3858,N_1943,N_1245);
xor U3859 (N_3859,N_1541,N_938);
nor U3860 (N_3860,N_783,N_231);
xor U3861 (N_3861,N_1432,N_661);
xnor U3862 (N_3862,N_177,N_1603);
or U3863 (N_3863,N_1926,N_534);
nor U3864 (N_3864,N_1170,N_1719);
or U3865 (N_3865,N_214,N_1054);
xnor U3866 (N_3866,N_389,N_625);
and U3867 (N_3867,N_272,N_11);
or U3868 (N_3868,N_387,N_1665);
nor U3869 (N_3869,N_1275,N_1709);
or U3870 (N_3870,N_1247,N_943);
nor U3871 (N_3871,N_1201,N_1896);
and U3872 (N_3872,N_219,N_1409);
xnor U3873 (N_3873,N_752,N_494);
nand U3874 (N_3874,N_1831,N_1845);
and U3875 (N_3875,N_376,N_1884);
nor U3876 (N_3876,N_1691,N_1328);
nand U3877 (N_3877,N_734,N_1177);
and U3878 (N_3878,N_1705,N_627);
nor U3879 (N_3879,N_681,N_1562);
and U3880 (N_3880,N_1249,N_893);
and U3881 (N_3881,N_601,N_269);
xor U3882 (N_3882,N_1614,N_1991);
and U3883 (N_3883,N_267,N_303);
or U3884 (N_3884,N_1078,N_1891);
nor U3885 (N_3885,N_830,N_1665);
xnor U3886 (N_3886,N_1470,N_1977);
or U3887 (N_3887,N_500,N_48);
and U3888 (N_3888,N_1297,N_1550);
and U3889 (N_3889,N_1706,N_1817);
nand U3890 (N_3890,N_1428,N_289);
or U3891 (N_3891,N_1158,N_669);
and U3892 (N_3892,N_166,N_1037);
xor U3893 (N_3893,N_521,N_44);
or U3894 (N_3894,N_383,N_557);
nand U3895 (N_3895,N_188,N_1882);
nor U3896 (N_3896,N_318,N_510);
and U3897 (N_3897,N_1540,N_1341);
xor U3898 (N_3898,N_40,N_1715);
nor U3899 (N_3899,N_831,N_1011);
or U3900 (N_3900,N_788,N_1204);
xor U3901 (N_3901,N_650,N_216);
xor U3902 (N_3902,N_833,N_251);
or U3903 (N_3903,N_345,N_623);
or U3904 (N_3904,N_1758,N_862);
nor U3905 (N_3905,N_1810,N_155);
nand U3906 (N_3906,N_1642,N_1004);
and U3907 (N_3907,N_1946,N_12);
nand U3908 (N_3908,N_819,N_1992);
nor U3909 (N_3909,N_1625,N_642);
xnor U3910 (N_3910,N_424,N_912);
nand U3911 (N_3911,N_1540,N_507);
or U3912 (N_3912,N_1138,N_118);
and U3913 (N_3913,N_435,N_1527);
xnor U3914 (N_3914,N_48,N_1268);
or U3915 (N_3915,N_1863,N_1488);
nor U3916 (N_3916,N_39,N_1370);
nor U3917 (N_3917,N_452,N_847);
nand U3918 (N_3918,N_69,N_1160);
nor U3919 (N_3919,N_1020,N_1241);
nand U3920 (N_3920,N_1091,N_1090);
and U3921 (N_3921,N_591,N_1797);
nor U3922 (N_3922,N_492,N_416);
nor U3923 (N_3923,N_1806,N_1154);
or U3924 (N_3924,N_408,N_1347);
xnor U3925 (N_3925,N_393,N_797);
nor U3926 (N_3926,N_899,N_911);
xnor U3927 (N_3927,N_717,N_97);
or U3928 (N_3928,N_1002,N_1679);
or U3929 (N_3929,N_1021,N_801);
nor U3930 (N_3930,N_447,N_1368);
xor U3931 (N_3931,N_1353,N_1865);
xnor U3932 (N_3932,N_1566,N_648);
nor U3933 (N_3933,N_749,N_1167);
xor U3934 (N_3934,N_1690,N_1822);
xnor U3935 (N_3935,N_679,N_424);
or U3936 (N_3936,N_1384,N_772);
nor U3937 (N_3937,N_553,N_324);
or U3938 (N_3938,N_1837,N_91);
and U3939 (N_3939,N_218,N_1847);
nand U3940 (N_3940,N_1997,N_578);
nand U3941 (N_3941,N_119,N_526);
and U3942 (N_3942,N_933,N_1978);
nand U3943 (N_3943,N_1644,N_1485);
xor U3944 (N_3944,N_150,N_439);
or U3945 (N_3945,N_440,N_67);
and U3946 (N_3946,N_1997,N_522);
xnor U3947 (N_3947,N_1585,N_1926);
or U3948 (N_3948,N_688,N_1399);
and U3949 (N_3949,N_134,N_1271);
nand U3950 (N_3950,N_445,N_203);
and U3951 (N_3951,N_1204,N_546);
xnor U3952 (N_3952,N_1620,N_502);
or U3953 (N_3953,N_66,N_778);
xor U3954 (N_3954,N_385,N_1670);
xor U3955 (N_3955,N_1127,N_1915);
xnor U3956 (N_3956,N_107,N_1300);
nor U3957 (N_3957,N_468,N_1482);
and U3958 (N_3958,N_968,N_367);
or U3959 (N_3959,N_1230,N_1206);
xnor U3960 (N_3960,N_946,N_674);
nand U3961 (N_3961,N_228,N_617);
xor U3962 (N_3962,N_1767,N_862);
and U3963 (N_3963,N_1420,N_1545);
and U3964 (N_3964,N_1291,N_1395);
or U3965 (N_3965,N_341,N_1501);
and U3966 (N_3966,N_1399,N_1972);
xor U3967 (N_3967,N_55,N_605);
nand U3968 (N_3968,N_1363,N_765);
and U3969 (N_3969,N_421,N_1840);
or U3970 (N_3970,N_1064,N_946);
nand U3971 (N_3971,N_142,N_162);
nor U3972 (N_3972,N_1224,N_325);
xor U3973 (N_3973,N_171,N_1593);
or U3974 (N_3974,N_1522,N_170);
xnor U3975 (N_3975,N_1531,N_1771);
nor U3976 (N_3976,N_580,N_681);
and U3977 (N_3977,N_1470,N_1709);
nand U3978 (N_3978,N_1124,N_749);
nand U3979 (N_3979,N_1711,N_1417);
nand U3980 (N_3980,N_1145,N_1571);
nand U3981 (N_3981,N_266,N_1278);
nand U3982 (N_3982,N_693,N_717);
nand U3983 (N_3983,N_1843,N_281);
or U3984 (N_3984,N_139,N_714);
nand U3985 (N_3985,N_813,N_859);
nor U3986 (N_3986,N_160,N_889);
xor U3987 (N_3987,N_506,N_1097);
and U3988 (N_3988,N_457,N_145);
nor U3989 (N_3989,N_1675,N_1704);
xnor U3990 (N_3990,N_1480,N_1702);
nor U3991 (N_3991,N_277,N_954);
nor U3992 (N_3992,N_534,N_1499);
xor U3993 (N_3993,N_654,N_1624);
nor U3994 (N_3994,N_1020,N_0);
or U3995 (N_3995,N_585,N_314);
and U3996 (N_3996,N_1817,N_1640);
xor U3997 (N_3997,N_1963,N_190);
xor U3998 (N_3998,N_1902,N_1540);
and U3999 (N_3999,N_1373,N_1254);
and U4000 (N_4000,N_3949,N_2568);
and U4001 (N_4001,N_3198,N_2224);
nand U4002 (N_4002,N_3181,N_2400);
nand U4003 (N_4003,N_3764,N_3218);
nor U4004 (N_4004,N_2064,N_2134);
or U4005 (N_4005,N_3752,N_2550);
or U4006 (N_4006,N_2390,N_3479);
xor U4007 (N_4007,N_2884,N_2947);
or U4008 (N_4008,N_2930,N_2563);
xnor U4009 (N_4009,N_3262,N_2066);
xnor U4010 (N_4010,N_2758,N_2438);
and U4011 (N_4011,N_3936,N_2079);
or U4012 (N_4012,N_3056,N_2045);
nand U4013 (N_4013,N_2242,N_3843);
and U4014 (N_4014,N_3363,N_2889);
xor U4015 (N_4015,N_2048,N_3509);
nor U4016 (N_4016,N_3478,N_3623);
xor U4017 (N_4017,N_2398,N_3840);
or U4018 (N_4018,N_2312,N_2248);
nand U4019 (N_4019,N_3951,N_3639);
xor U4020 (N_4020,N_3435,N_2547);
xnor U4021 (N_4021,N_2310,N_2073);
or U4022 (N_4022,N_3127,N_3605);
nand U4023 (N_4023,N_3595,N_3396);
xnor U4024 (N_4024,N_3297,N_2342);
or U4025 (N_4025,N_2567,N_3737);
xor U4026 (N_4026,N_2611,N_2839);
or U4027 (N_4027,N_2043,N_3770);
nor U4028 (N_4028,N_3966,N_3771);
xnor U4029 (N_4029,N_3142,N_3367);
and U4030 (N_4030,N_3909,N_2120);
and U4031 (N_4031,N_2991,N_3229);
xnor U4032 (N_4032,N_3295,N_3985);
or U4033 (N_4033,N_3634,N_3612);
nor U4034 (N_4034,N_2363,N_3233);
xor U4035 (N_4035,N_3819,N_3400);
nor U4036 (N_4036,N_3282,N_3473);
nor U4037 (N_4037,N_2492,N_3934);
and U4038 (N_4038,N_2650,N_2440);
and U4039 (N_4039,N_3266,N_3824);
xor U4040 (N_4040,N_3372,N_2419);
or U4041 (N_4041,N_2628,N_3258);
or U4042 (N_4042,N_3947,N_2745);
or U4043 (N_4043,N_2574,N_3038);
xnor U4044 (N_4044,N_3861,N_2952);
nor U4045 (N_4045,N_2171,N_2725);
or U4046 (N_4046,N_3059,N_3796);
nor U4047 (N_4047,N_3418,N_3125);
nor U4048 (N_4048,N_2843,N_2649);
xnor U4049 (N_4049,N_2881,N_2226);
and U4050 (N_4050,N_3350,N_3781);
and U4051 (N_4051,N_2380,N_3802);
nand U4052 (N_4052,N_3371,N_2987);
or U4053 (N_4053,N_2526,N_2504);
and U4054 (N_4054,N_2521,N_2957);
nand U4055 (N_4055,N_2657,N_3621);
nor U4056 (N_4056,N_2127,N_2821);
or U4057 (N_4057,N_3070,N_2227);
xnor U4058 (N_4058,N_3289,N_3535);
nor U4059 (N_4059,N_3719,N_2466);
nand U4060 (N_4060,N_3483,N_3585);
or U4061 (N_4061,N_2265,N_3669);
or U4062 (N_4062,N_2922,N_2002);
nand U4063 (N_4063,N_3943,N_2395);
xnor U4064 (N_4064,N_3183,N_2690);
nor U4065 (N_4065,N_3196,N_2644);
and U4066 (N_4066,N_2793,N_3434);
nand U4067 (N_4067,N_3139,N_3041);
nand U4068 (N_4068,N_2050,N_2605);
and U4069 (N_4069,N_3128,N_3228);
nand U4070 (N_4070,N_2182,N_3477);
nor U4071 (N_4071,N_3880,N_3083);
xnor U4072 (N_4072,N_3078,N_3531);
nand U4073 (N_4073,N_3954,N_2092);
nor U4074 (N_4074,N_2473,N_3376);
xnor U4075 (N_4075,N_2875,N_3748);
xnor U4076 (N_4076,N_3699,N_3809);
or U4077 (N_4077,N_2237,N_3785);
nor U4078 (N_4078,N_2966,N_3582);
nand U4079 (N_4079,N_3867,N_2715);
nand U4080 (N_4080,N_2365,N_2424);
nor U4081 (N_4081,N_3285,N_2943);
nor U4082 (N_4082,N_3518,N_3447);
and U4083 (N_4083,N_3377,N_3865);
xnor U4084 (N_4084,N_2378,N_2070);
nor U4085 (N_4085,N_2019,N_2137);
or U4086 (N_4086,N_2594,N_2458);
nor U4087 (N_4087,N_2729,N_3104);
and U4088 (N_4088,N_2586,N_3787);
xor U4089 (N_4089,N_2445,N_3030);
xnor U4090 (N_4090,N_3932,N_2435);
and U4091 (N_4091,N_3797,N_2882);
nand U4092 (N_4092,N_3099,N_2340);
xnor U4093 (N_4093,N_2232,N_3587);
and U4094 (N_4094,N_2996,N_3711);
and U4095 (N_4095,N_2308,N_3720);
and U4096 (N_4096,N_3302,N_3792);
nand U4097 (N_4097,N_2921,N_3501);
nor U4098 (N_4098,N_3899,N_3525);
or U4099 (N_4099,N_2710,N_2155);
nand U4100 (N_4100,N_3293,N_3604);
nor U4101 (N_4101,N_3015,N_3722);
xor U4102 (N_4102,N_3217,N_2476);
and U4103 (N_4103,N_2447,N_3742);
and U4104 (N_4104,N_2785,N_3517);
and U4105 (N_4105,N_2795,N_2280);
and U4106 (N_4106,N_3321,N_3608);
and U4107 (N_4107,N_2302,N_2416);
nor U4108 (N_4108,N_3897,N_3859);
xor U4109 (N_4109,N_3607,N_3050);
nand U4110 (N_4110,N_2756,N_3622);
nor U4111 (N_4111,N_3158,N_3715);
or U4112 (N_4112,N_2728,N_2203);
nor U4113 (N_4113,N_3378,N_3788);
nor U4114 (N_4114,N_3355,N_3731);
xnor U4115 (N_4115,N_2080,N_2722);
xnor U4116 (N_4116,N_2152,N_3270);
nor U4117 (N_4117,N_3693,N_3666);
nor U4118 (N_4118,N_2746,N_2848);
or U4119 (N_4119,N_2626,N_2772);
nand U4120 (N_4120,N_3594,N_3994);
or U4121 (N_4121,N_3221,N_2115);
nand U4122 (N_4122,N_2510,N_3998);
or U4123 (N_4123,N_2888,N_3893);
and U4124 (N_4124,N_3095,N_2298);
and U4125 (N_4125,N_3468,N_2714);
nor U4126 (N_4126,N_3387,N_3098);
xnor U4127 (N_4127,N_3432,N_3779);
xor U4128 (N_4128,N_3138,N_2251);
xor U4129 (N_4129,N_3598,N_2621);
or U4130 (N_4130,N_2235,N_2779);
nand U4131 (N_4131,N_2275,N_2643);
xor U4132 (N_4132,N_2544,N_3904);
nor U4133 (N_4133,N_3987,N_2844);
xnor U4134 (N_4134,N_2300,N_3090);
xor U4135 (N_4135,N_3444,N_2011);
or U4136 (N_4136,N_3741,N_2314);
nand U4137 (N_4137,N_2800,N_2318);
and U4138 (N_4138,N_3045,N_3386);
xor U4139 (N_4139,N_2030,N_3273);
or U4140 (N_4140,N_3858,N_2478);
nand U4141 (N_4141,N_3398,N_2929);
nand U4142 (N_4142,N_2332,N_2420);
or U4143 (N_4143,N_2076,N_3401);
and U4144 (N_4144,N_3870,N_3251);
nand U4145 (N_4145,N_3414,N_2838);
nor U4146 (N_4146,N_2106,N_2260);
nand U4147 (N_4147,N_3991,N_2322);
nand U4148 (N_4148,N_3499,N_3529);
or U4149 (N_4149,N_3431,N_2055);
xor U4150 (N_4150,N_2439,N_3766);
xnor U4151 (N_4151,N_2486,N_2387);
nor U4152 (N_4152,N_3135,N_2956);
or U4153 (N_4153,N_3010,N_3492);
nand U4154 (N_4154,N_2743,N_3680);
xnor U4155 (N_4155,N_3922,N_3278);
and U4156 (N_4156,N_3397,N_2924);
nor U4157 (N_4157,N_2598,N_2412);
and U4158 (N_4158,N_2170,N_3872);
or U4159 (N_4159,N_2289,N_2602);
or U4160 (N_4160,N_2427,N_3163);
nor U4161 (N_4161,N_2978,N_3537);
and U4162 (N_4162,N_3487,N_3189);
nand U4163 (N_4163,N_3765,N_2484);
and U4164 (N_4164,N_2601,N_3505);
xnor U4165 (N_4165,N_2078,N_2908);
or U4166 (N_4166,N_3154,N_3878);
nand U4167 (N_4167,N_2951,N_2151);
nand U4168 (N_4168,N_2680,N_3426);
and U4169 (N_4169,N_3596,N_2121);
or U4170 (N_4170,N_2075,N_2249);
or U4171 (N_4171,N_2971,N_2358);
or U4172 (N_4172,N_3354,N_2907);
or U4173 (N_4173,N_2430,N_3245);
nor U4174 (N_4174,N_2708,N_3438);
nand U4175 (N_4175,N_2692,N_2652);
nor U4176 (N_4176,N_3724,N_3006);
nor U4177 (N_4177,N_2571,N_2784);
nor U4178 (N_4178,N_3694,N_3250);
nand U4179 (N_4179,N_3451,N_2349);
and U4180 (N_4180,N_3649,N_3532);
or U4181 (N_4181,N_2899,N_3567);
nor U4182 (N_4182,N_3283,N_3881);
and U4183 (N_4183,N_2126,N_3199);
and U4184 (N_4184,N_3343,N_3891);
xor U4185 (N_4185,N_3094,N_3412);
and U4186 (N_4186,N_2897,N_3352);
nand U4187 (N_4187,N_2753,N_3082);
nor U4188 (N_4188,N_3981,N_3330);
and U4189 (N_4189,N_3032,N_2836);
nand U4190 (N_4190,N_3915,N_3068);
or U4191 (N_4191,N_2191,N_3905);
nor U4192 (N_4192,N_2056,N_2503);
and U4193 (N_4193,N_2431,N_3241);
nor U4194 (N_4194,N_2781,N_3149);
and U4195 (N_4195,N_2536,N_2317);
xor U4196 (N_4196,N_2590,N_3803);
or U4197 (N_4197,N_2997,N_2004);
xor U4198 (N_4198,N_2861,N_3761);
or U4199 (N_4199,N_3342,N_3838);
xnor U4200 (N_4200,N_3676,N_2767);
and U4201 (N_4201,N_3296,N_2067);
nand U4202 (N_4202,N_2456,N_3854);
nor U4203 (N_4203,N_2969,N_3417);
nand U4204 (N_4204,N_3557,N_3713);
nor U4205 (N_4205,N_2580,N_2009);
or U4206 (N_4206,N_2000,N_2118);
xor U4207 (N_4207,N_3945,N_3613);
or U4208 (N_4208,N_2663,N_3144);
and U4209 (N_4209,N_2864,N_3804);
nor U4210 (N_4210,N_3333,N_3236);
xnor U4211 (N_4211,N_2297,N_2948);
nor U4212 (N_4212,N_2341,N_3207);
xor U4213 (N_4213,N_3661,N_2255);
and U4214 (N_4214,N_2560,N_2119);
or U4215 (N_4215,N_2388,N_2968);
nand U4216 (N_4216,N_2196,N_3561);
or U4217 (N_4217,N_2188,N_3392);
and U4218 (N_4218,N_3203,N_2411);
nor U4219 (N_4219,N_2519,N_2407);
xnor U4220 (N_4220,N_2805,N_2937);
xor U4221 (N_4221,N_2647,N_2160);
nand U4222 (N_4222,N_2344,N_3406);
nor U4223 (N_4223,N_3055,N_3572);
nor U4224 (N_4224,N_3000,N_3800);
and U4225 (N_4225,N_3408,N_3222);
or U4226 (N_4226,N_3807,N_2423);
nand U4227 (N_4227,N_3977,N_2443);
xnor U4228 (N_4228,N_3433,N_3209);
nor U4229 (N_4229,N_2624,N_2288);
and U4230 (N_4230,N_2741,N_3982);
or U4231 (N_4231,N_2665,N_3996);
nand U4232 (N_4232,N_3832,N_2819);
or U4233 (N_4233,N_3374,N_3690);
nor U4234 (N_4234,N_3860,N_3303);
nor U4235 (N_4235,N_2213,N_3717);
or U4236 (N_4236,N_2989,N_2931);
or U4237 (N_4237,N_3555,N_2459);
xor U4238 (N_4238,N_2404,N_3573);
and U4239 (N_4239,N_2866,N_2285);
xnor U4240 (N_4240,N_3329,N_2012);
nand U4241 (N_4241,N_2813,N_3110);
or U4242 (N_4242,N_3405,N_2862);
nor U4243 (N_4243,N_2027,N_3002);
and U4244 (N_4244,N_2629,N_3362);
or U4245 (N_4245,N_3153,N_2942);
or U4246 (N_4246,N_2667,N_2166);
and U4247 (N_4247,N_2790,N_2986);
xnor U4248 (N_4248,N_3235,N_3076);
nand U4249 (N_4249,N_2099,N_2198);
nor U4250 (N_4250,N_3618,N_2422);
xor U4251 (N_4251,N_3472,N_3575);
or U4252 (N_4252,N_2316,N_3581);
or U4253 (N_4253,N_3710,N_2920);
or U4254 (N_4254,N_2052,N_2592);
xnor U4255 (N_4255,N_2186,N_3663);
or U4256 (N_4256,N_2108,N_3026);
or U4257 (N_4257,N_2900,N_2306);
and U4258 (N_4258,N_2675,N_2259);
and U4259 (N_4259,N_2522,N_3786);
nand U4260 (N_4260,N_3545,N_2671);
nor U4261 (N_4261,N_2225,N_2085);
nor U4262 (N_4262,N_3332,N_2071);
xnor U4263 (N_4263,N_2549,N_3044);
nand U4264 (N_4264,N_3877,N_2190);
and U4265 (N_4265,N_2311,N_2591);
xor U4266 (N_4266,N_2293,N_3320);
xor U4267 (N_4267,N_3570,N_3062);
and U4268 (N_4268,N_2373,N_2946);
nor U4269 (N_4269,N_2001,N_3016);
xnor U4270 (N_4270,N_3475,N_2918);
nand U4271 (N_4271,N_2670,N_3052);
xnor U4272 (N_4272,N_3071,N_2169);
or U4273 (N_4273,N_3830,N_3265);
nor U4274 (N_4274,N_3656,N_2891);
and U4275 (N_4275,N_3856,N_2672);
and U4276 (N_4276,N_3459,N_2719);
or U4277 (N_4277,N_3349,N_3725);
nor U4278 (N_4278,N_3769,N_2286);
nor U4279 (N_4279,N_2938,N_3419);
or U4280 (N_4280,N_3974,N_3166);
nor U4281 (N_4281,N_3577,N_2381);
nand U4282 (N_4282,N_3997,N_2425);
xor U4283 (N_4283,N_2187,N_2666);
or U4284 (N_4284,N_3541,N_3004);
or U4285 (N_4285,N_2578,N_3772);
and U4286 (N_4286,N_3616,N_2513);
nor U4287 (N_4287,N_3970,N_2802);
nand U4288 (N_4288,N_3674,N_2554);
xnor U4289 (N_4289,N_3540,N_3727);
nor U4290 (N_4290,N_3176,N_3976);
and U4291 (N_4291,N_2887,N_2041);
nor U4292 (N_4292,N_2777,N_2944);
and U4293 (N_4293,N_2535,N_3448);
nand U4294 (N_4294,N_2877,N_3122);
and U4295 (N_4295,N_2765,N_2069);
nor U4296 (N_4296,N_3884,N_2327);
nand U4297 (N_4297,N_3200,N_2616);
or U4298 (N_4298,N_2494,N_3558);
nand U4299 (N_4299,N_3850,N_2036);
or U4300 (N_4300,N_3630,N_3365);
nor U4301 (N_4301,N_2180,N_2637);
nor U4302 (N_4302,N_2252,N_2434);
nor U4303 (N_4303,N_2183,N_3047);
nor U4304 (N_4304,N_3500,N_2214);
and U4305 (N_4305,N_3167,N_3436);
xnor U4306 (N_4306,N_3822,N_3703);
or U4307 (N_4307,N_2525,N_2818);
xnor U4308 (N_4308,N_3257,N_2524);
nand U4309 (N_4309,N_2654,N_3020);
or U4310 (N_4310,N_3827,N_3467);
and U4311 (N_4311,N_3667,N_2832);
or U4312 (N_4312,N_3999,N_2148);
and U4313 (N_4313,N_3526,N_2613);
and U4314 (N_4314,N_2321,N_2769);
nand U4315 (N_4315,N_2366,N_2829);
nor U4316 (N_4316,N_3873,N_3952);
nand U4317 (N_4317,N_2982,N_2147);
nand U4318 (N_4318,N_2748,N_2913);
nor U4319 (N_4319,N_3043,N_3294);
nand U4320 (N_4320,N_3248,N_3197);
nor U4321 (N_4321,N_3276,N_2046);
xnor U4322 (N_4322,N_3601,N_2354);
nand U4323 (N_4323,N_2051,N_2515);
xnor U4324 (N_4324,N_3346,N_2974);
xnor U4325 (N_4325,N_3390,N_3931);
xnor U4326 (N_4326,N_2122,N_2172);
and U4327 (N_4327,N_3721,N_2263);
and U4328 (N_4328,N_3394,N_2017);
nor U4329 (N_4329,N_2348,N_3161);
xor U4330 (N_4330,N_3373,N_3140);
nor U4331 (N_4331,N_3341,N_2361);
nand U4332 (N_4332,N_2809,N_3627);
or U4333 (N_4333,N_3688,N_2408);
nor U4334 (N_4334,N_2206,N_2631);
and U4335 (N_4335,N_3496,N_2759);
xor U4336 (N_4336,N_2697,N_3316);
xor U4337 (N_4337,N_3995,N_3061);
xnor U4338 (N_4338,N_2735,N_3280);
xor U4339 (N_4339,N_3718,N_3370);
nor U4340 (N_4340,N_2678,N_3464);
nor U4341 (N_4341,N_2406,N_3421);
or U4342 (N_4342,N_2061,N_2682);
or U4343 (N_4343,N_3253,N_3215);
or U4344 (N_4344,N_3136,N_2863);
nand U4345 (N_4345,N_3389,N_3143);
nor U4346 (N_4346,N_2016,N_2333);
and U4347 (N_4347,N_2330,N_3599);
and U4348 (N_4348,N_3449,N_2295);
nor U4349 (N_4349,N_2860,N_2737);
nor U4350 (N_4350,N_3677,N_2038);
and U4351 (N_4351,N_2977,N_2757);
or U4352 (N_4352,N_2744,N_2830);
and U4353 (N_4353,N_2250,N_3420);
nand U4354 (N_4354,N_2964,N_3036);
or U4355 (N_4355,N_2551,N_3527);
xnor U4356 (N_4356,N_2548,N_3851);
and U4357 (N_4357,N_3456,N_2385);
and U4358 (N_4358,N_3279,N_2796);
nand U4359 (N_4359,N_2794,N_3455);
xnor U4360 (N_4360,N_3442,N_2615);
nand U4361 (N_4361,N_2975,N_3675);
xnor U4362 (N_4362,N_2619,N_2498);
nand U4363 (N_4363,N_2337,N_2869);
xor U4364 (N_4364,N_2681,N_3410);
nor U4365 (N_4365,N_3120,N_3428);
nand U4366 (N_4366,N_3441,N_3654);
xor U4367 (N_4367,N_3211,N_2386);
or U4368 (N_4368,N_2552,N_3182);
and U4369 (N_4369,N_2717,N_2060);
xnor U4370 (N_4370,N_2357,N_2904);
nand U4371 (N_4371,N_3275,N_2676);
or U4372 (N_4372,N_3988,N_2851);
nor U4373 (N_4373,N_2970,N_2609);
nor U4374 (N_4374,N_2556,N_2668);
xor U4375 (N_4375,N_3466,N_2846);
and U4376 (N_4376,N_3723,N_2688);
xor U4377 (N_4377,N_3544,N_2402);
and U4378 (N_4378,N_2584,N_2895);
xor U4379 (N_4379,N_2527,N_2367);
nor U4380 (N_4380,N_3190,N_2197);
nand U4381 (N_4381,N_3668,N_2362);
nor U4382 (N_4382,N_3866,N_3583);
nor U4383 (N_4383,N_2648,N_3755);
nand U4384 (N_4384,N_3898,N_2468);
nand U4385 (N_4385,N_3053,N_2502);
nand U4386 (N_4386,N_2645,N_3430);
and U4387 (N_4387,N_3172,N_3829);
nor U4388 (N_4388,N_3782,N_3214);
nand U4389 (N_4389,N_2501,N_2480);
nor U4390 (N_4390,N_2094,N_3510);
xor U4391 (N_4391,N_3543,N_3778);
nand U4392 (N_4392,N_3784,N_2896);
nand U4393 (N_4393,N_3488,N_3437);
xor U4394 (N_4394,N_2117,N_2764);
and U4395 (N_4395,N_3029,N_2471);
or U4396 (N_4396,N_2077,N_2216);
and U4397 (N_4397,N_2927,N_2919);
nand U4398 (N_4398,N_3151,N_3252);
and U4399 (N_4399,N_2426,N_3048);
nor U4400 (N_4400,N_2816,N_2014);
nor U4401 (N_4401,N_2910,N_2393);
nor U4402 (N_4402,N_2441,N_2095);
and U4403 (N_4403,N_3660,N_3628);
and U4404 (N_4404,N_2256,N_2024);
xnor U4405 (N_4405,N_3284,N_2988);
nand U4406 (N_4406,N_2985,N_2158);
xnor U4407 (N_4407,N_2335,N_2161);
or U4408 (N_4408,N_3027,N_3923);
and U4409 (N_4409,N_2999,N_3476);
xnor U4410 (N_4410,N_2025,N_2489);
nor U4411 (N_4411,N_3744,N_2980);
and U4412 (N_4412,N_3009,N_3042);
nand U4413 (N_4413,N_3092,N_3566);
or U4414 (N_4414,N_3695,N_2033);
and U4415 (N_4415,N_3465,N_2762);
nor U4416 (N_4416,N_3754,N_3471);
nor U4417 (N_4417,N_3051,N_3632);
or U4418 (N_4418,N_3534,N_2105);
and U4419 (N_4419,N_3638,N_2053);
and U4420 (N_4420,N_2143,N_2482);
and U4421 (N_4421,N_2808,N_2042);
xnor U4422 (N_4422,N_3298,N_2916);
or U4423 (N_4423,N_2520,N_3067);
nor U4424 (N_4424,N_3460,N_3486);
nor U4425 (N_4425,N_2261,N_3249);
nor U4426 (N_4426,N_3767,N_3935);
and U4427 (N_4427,N_2129,N_3559);
and U4428 (N_4428,N_3131,N_2834);
nand U4429 (N_4429,N_2890,N_2448);
xnor U4430 (N_4430,N_2313,N_3168);
nand U4431 (N_4431,N_2465,N_3446);
nand U4432 (N_4432,N_3485,N_3673);
nor U4433 (N_4433,N_2343,N_2063);
and U4434 (N_4434,N_3763,N_3357);
and U4435 (N_4435,N_3963,N_3910);
nor U4436 (N_4436,N_2325,N_2353);
nand U4437 (N_4437,N_3696,N_3890);
nand U4438 (N_4438,N_3833,N_2683);
nand U4439 (N_4439,N_2189,N_3857);
xor U4440 (N_4440,N_3202,N_3777);
or U4441 (N_4441,N_3037,N_2955);
xor U4442 (N_4442,N_3708,N_3889);
and U4443 (N_4443,N_2491,N_3416);
nor U4444 (N_4444,N_2278,N_2040);
nand U4445 (N_4445,N_2181,N_2806);
nor U4446 (N_4446,N_2479,N_3242);
and U4447 (N_4447,N_2693,N_2368);
nor U4448 (N_4448,N_3692,N_3759);
and U4449 (N_4449,N_2810,N_3733);
nor U4450 (N_4450,N_3232,N_2352);
nor U4451 (N_4451,N_3173,N_3220);
nand U4452 (N_4452,N_2842,N_2537);
nand U4453 (N_4453,N_3237,N_2451);
and U4454 (N_4454,N_3790,N_2273);
nor U4455 (N_4455,N_2347,N_3109);
nand U4456 (N_4456,N_2081,N_3576);
or U4457 (N_4457,N_3641,N_2589);
or U4458 (N_4458,N_2309,N_3930);
and U4459 (N_4459,N_3938,N_2096);
xor U4460 (N_4460,N_2469,N_3498);
nand U4461 (N_4461,N_3698,N_3735);
xor U4462 (N_4462,N_3075,N_3972);
and U4463 (N_4463,N_3883,N_2461);
nand U4464 (N_4464,N_2374,N_3597);
and U4465 (N_4465,N_2359,N_3848);
or U4466 (N_4466,N_2664,N_3239);
nand U4467 (N_4467,N_3569,N_2215);
nand U4468 (N_4468,N_3334,N_3863);
nand U4469 (N_4469,N_2691,N_3074);
nand U4470 (N_4470,N_3916,N_3491);
nand U4471 (N_4471,N_2820,N_2562);
or U4472 (N_4472,N_2801,N_2209);
nand U4473 (N_4473,N_3150,N_2057);
or U4474 (N_4474,N_2138,N_3753);
nand U4475 (N_4475,N_2903,N_2059);
xor U4476 (N_4476,N_3129,N_2642);
or U4477 (N_4477,N_3012,N_3568);
xor U4478 (N_4478,N_2013,N_2211);
xor U4479 (N_4479,N_2369,N_3908);
xor U4480 (N_4480,N_3423,N_2817);
and U4481 (N_4481,N_3216,N_2886);
nor U4482 (N_4482,N_3462,N_2267);
nor U4483 (N_4483,N_2290,N_2506);
nand U4484 (N_4484,N_3705,N_2018);
nand U4485 (N_4485,N_3609,N_2831);
nor U4486 (N_4486,N_3516,N_3747);
and U4487 (N_4487,N_3826,N_3980);
nor U4488 (N_4488,N_2130,N_3642);
nor U4489 (N_4489,N_3671,N_2032);
nand U4490 (N_4490,N_3750,N_2727);
xor U4491 (N_4491,N_2540,N_3014);
xnor U4492 (N_4492,N_2339,N_3204);
and U4493 (N_4493,N_2375,N_3152);
or U4494 (N_4494,N_3846,N_3162);
or U4495 (N_4495,N_2814,N_3480);
or U4496 (N_4496,N_2703,N_3939);
nand U4497 (N_4497,N_2852,N_3385);
and U4498 (N_4498,N_2518,N_3077);
and U4499 (N_4499,N_3689,N_2301);
xnor U4500 (N_4500,N_2659,N_2008);
nand U4501 (N_4501,N_2163,N_3658);
nor U4502 (N_4502,N_3664,N_2803);
and U4503 (N_4503,N_3105,N_2338);
xnor U4504 (N_4504,N_2505,N_2539);
or U4505 (N_4505,N_3402,N_3709);
xnor U4506 (N_4506,N_3672,N_3137);
nand U4507 (N_4507,N_2700,N_2088);
xor U4508 (N_4508,N_2559,N_2721);
or U4509 (N_4509,N_3812,N_2754);
nand U4510 (N_4510,N_3941,N_2516);
or U4511 (N_4511,N_2835,N_3841);
and U4512 (N_4512,N_2604,N_2442);
nor U4513 (N_4513,N_3968,N_3917);
or U4514 (N_4514,N_2558,N_2168);
nand U4515 (N_4515,N_3992,N_2822);
or U4516 (N_4516,N_2065,N_3834);
or U4517 (N_4517,N_2090,N_3679);
xnor U4518 (N_4518,N_2892,N_3358);
xor U4519 (N_4519,N_2379,N_3046);
or U4520 (N_4520,N_2773,N_3697);
xor U4521 (N_4521,N_2054,N_2768);
and U4522 (N_4522,N_3331,N_3361);
nor U4523 (N_4523,N_2315,N_2857);
and U4524 (N_4524,N_2086,N_3729);
or U4525 (N_4525,N_2883,N_2973);
nor U4526 (N_4526,N_3828,N_3403);
nor U4527 (N_4527,N_3290,N_3281);
and U4528 (N_4528,N_3413,N_3901);
or U4529 (N_4529,N_3180,N_2015);
and U4530 (N_4530,N_3712,N_3637);
and U4531 (N_4531,N_3590,N_2771);
nor U4532 (N_4532,N_3762,N_3603);
and U4533 (N_4533,N_2911,N_3887);
or U4534 (N_4534,N_3508,N_2238);
and U4535 (N_4535,N_2142,N_2859);
nand U4536 (N_4536,N_3339,N_2320);
or U4537 (N_4537,N_2413,N_3903);
xor U4538 (N_4538,N_2872,N_3886);
and U4539 (N_4539,N_3682,N_2173);
nand U4540 (N_4540,N_3017,N_2894);
nor U4541 (N_4541,N_3079,N_3523);
and U4542 (N_4542,N_3538,N_2135);
or U4543 (N_4543,N_3123,N_2110);
nand U4544 (N_4544,N_2268,N_2928);
or U4545 (N_4545,N_3549,N_2454);
nor U4546 (N_4546,N_2625,N_3457);
nor U4547 (N_4547,N_3645,N_2608);
and U4548 (N_4548,N_2274,N_2185);
xnor U4549 (N_4549,N_3574,N_2087);
nand U4550 (N_4550,N_3539,N_3502);
xnor U4551 (N_4551,N_3876,N_2326);
or U4552 (N_4552,N_3458,N_2926);
or U4553 (N_4553,N_2370,N_3793);
or U4554 (N_4554,N_3962,N_3328);
nand U4555 (N_4555,N_2915,N_3101);
or U4556 (N_4556,N_3187,N_2689);
and U4557 (N_4557,N_2739,N_2940);
xor U4558 (N_4558,N_3452,N_2695);
nand U4559 (N_4559,N_3900,N_3964);
or U4560 (N_4560,N_2245,N_3814);
and U4561 (N_4561,N_2202,N_3184);
and U4562 (N_4562,N_3315,N_3023);
and U4563 (N_4563,N_3324,N_2778);
nor U4564 (N_4564,N_3269,N_3978);
nand U4565 (N_4565,N_3989,N_2564);
or U4566 (N_4566,N_2512,N_3686);
nand U4567 (N_4567,N_3164,N_2749);
nand U4568 (N_4568,N_2194,N_3337);
xor U4569 (N_4569,N_2270,N_2391);
or U4570 (N_4570,N_2673,N_2847);
and U4571 (N_4571,N_3835,N_3178);
and U4572 (N_4572,N_3513,N_2112);
or U4573 (N_4573,N_3836,N_3121);
xor U4574 (N_4574,N_3979,N_3234);
and U4575 (N_4575,N_2463,N_2623);
nand U4576 (N_4576,N_2264,N_3111);
or U4577 (N_4577,N_3443,N_2994);
nand U4578 (N_4578,N_2706,N_3906);
and U4579 (N_4579,N_3065,N_2418);
or U4580 (N_4580,N_3847,N_2219);
xnor U4581 (N_4581,N_2350,N_2236);
and U4582 (N_4582,N_2319,N_3493);
nand U4583 (N_4583,N_3054,N_2953);
nor U4584 (N_4584,N_2156,N_2107);
or U4585 (N_4585,N_2874,N_3615);
nor U4586 (N_4586,N_2935,N_3732);
xnor U4587 (N_4587,N_3309,N_2677);
nand U4588 (N_4588,N_2934,N_3929);
or U4589 (N_4589,N_2638,N_3469);
and U4590 (N_4590,N_3805,N_3107);
xnor U4591 (N_4591,N_3288,N_3586);
or U4592 (N_4592,N_3126,N_3560);
and U4593 (N_4593,N_2035,N_3356);
and U4594 (N_4594,N_2356,N_2597);
or U4595 (N_4595,N_2139,N_2660);
xnor U4596 (N_4596,N_2641,N_3519);
nand U4597 (N_4597,N_2020,N_2993);
or U4598 (N_4598,N_2210,N_2507);
nand U4599 (N_4599,N_2072,N_2849);
nor U4600 (N_4600,N_3625,N_3990);
and U4601 (N_4601,N_3381,N_3894);
xnor U4602 (N_4602,N_2091,N_3192);
and U4603 (N_4603,N_2579,N_3201);
nand U4604 (N_4604,N_3461,N_2833);
and U4605 (N_4605,N_2639,N_2058);
and U4606 (N_4606,N_3040,N_2201);
xor U4607 (N_4607,N_3146,N_2279);
nor U4608 (N_4608,N_2429,N_2855);
xor U4609 (N_4609,N_3058,N_3636);
nor U4610 (N_4610,N_3340,N_3427);
or U4611 (N_4611,N_2799,N_2724);
or U4612 (N_4612,N_2195,N_2470);
nor U4613 (N_4613,N_3463,N_3657);
xnor U4614 (N_4614,N_2167,N_3961);
nand U4615 (N_4615,N_2392,N_3003);
and U4616 (N_4616,N_2364,N_2736);
nor U4617 (N_4617,N_3593,N_3205);
or U4618 (N_4618,N_3028,N_3415);
nand U4619 (N_4619,N_2824,N_3844);
nor U4620 (N_4620,N_3681,N_3305);
and U4621 (N_4621,N_3259,N_2208);
nor U4622 (N_4622,N_2698,N_2726);
or U4623 (N_4623,N_3975,N_2243);
xor U4624 (N_4624,N_3959,N_2958);
nor U4625 (N_4625,N_3195,N_3034);
and U4626 (N_4626,N_3351,N_2788);
xor U4627 (N_4627,N_3301,N_2912);
or U4628 (N_4628,N_2932,N_3097);
nor U4629 (N_4629,N_2811,N_2389);
xor U4630 (N_4630,N_3287,N_3825);
or U4631 (N_4631,N_3399,N_3611);
and U4632 (N_4632,N_3422,N_3955);
xor U4633 (N_4633,N_2854,N_2346);
nand U4634 (N_4634,N_3626,N_2109);
and U4635 (N_4635,N_2179,N_2959);
and U4636 (N_4636,N_2104,N_3823);
xor U4637 (N_4637,N_2394,N_3528);
nor U4638 (N_4638,N_2377,N_3018);
xor U4639 (N_4639,N_2184,N_3918);
and U4640 (N_4640,N_3852,N_2098);
xor U4641 (N_4641,N_2674,N_2410);
or U4642 (N_4642,N_3277,N_2783);
nor U4643 (N_4643,N_2546,N_3610);
and U4644 (N_4644,N_3141,N_2662);
nand U4645 (N_4645,N_2444,N_2967);
nand U4646 (N_4646,N_2789,N_3384);
or U4647 (N_4647,N_2807,N_3326);
xnor U4648 (N_4648,N_2157,N_2026);
nor U4649 (N_4649,N_2747,N_2610);
and U4650 (N_4650,N_3393,N_3547);
or U4651 (N_4651,N_2841,N_2917);
and U4652 (N_4652,N_2514,N_3546);
nor U4653 (N_4653,N_2401,N_3862);
nand U4654 (N_4654,N_3885,N_3080);
nand U4655 (N_4655,N_2532,N_2871);
or U4656 (N_4656,N_3633,N_2508);
nand U4657 (N_4657,N_2292,N_2296);
nand U4658 (N_4658,N_3914,N_2557);
xor U4659 (N_4659,N_2257,N_2382);
and U4660 (N_4660,N_2711,N_3148);
nand U4661 (N_4661,N_3177,N_2089);
or U4662 (N_4662,N_2751,N_3319);
and U4663 (N_4663,N_3210,N_3085);
xor U4664 (N_4664,N_3564,N_2720);
and U4665 (N_4665,N_2763,N_2240);
or U4666 (N_4666,N_3274,N_3662);
and U4667 (N_4667,N_3704,N_2617);
or U4668 (N_4668,N_3219,N_3347);
nor U4669 (N_4669,N_3993,N_3839);
nand U4670 (N_4670,N_2331,N_2607);
and U4671 (N_4671,N_3619,N_2797);
nand U4672 (N_4672,N_2705,N_3132);
or U4673 (N_4673,N_2812,N_3179);
or U4674 (N_4674,N_2475,N_3606);
nand U4675 (N_4675,N_3286,N_3069);
nor U4676 (N_4676,N_2084,N_2282);
nand U4677 (N_4677,N_3327,N_2113);
xnor U4678 (N_4678,N_2217,N_3650);
xor U4679 (N_4679,N_3481,N_2658);
nor U4680 (N_4680,N_3255,N_3145);
or U4681 (N_4681,N_2124,N_2481);
xnor U4682 (N_4682,N_2254,N_3511);
or U4683 (N_4683,N_3013,N_3185);
nand U4684 (N_4684,N_3300,N_3306);
and U4685 (N_4685,N_3260,N_2154);
or U4686 (N_4686,N_2867,N_2174);
nand U4687 (N_4687,N_3169,N_2511);
nor U4688 (N_4688,N_2984,N_2409);
and U4689 (N_4689,N_3631,N_3556);
xnor U4690 (N_4690,N_3317,N_2945);
nor U4691 (N_4691,N_2023,N_3159);
or U4692 (N_4692,N_2840,N_2983);
or U4693 (N_4693,N_3652,N_3308);
and U4694 (N_4694,N_2488,N_2414);
or U4695 (N_4695,N_2123,N_2543);
xor U4696 (N_4696,N_2272,N_2165);
nor U4697 (N_4697,N_3757,N_3942);
or U4698 (N_4698,N_3614,N_3060);
xnor U4699 (N_4699,N_3780,N_3548);
nand U4700 (N_4700,N_3325,N_3494);
or U4701 (N_4701,N_3360,N_2307);
xor U4702 (N_4702,N_2878,N_2399);
nor U4703 (N_4703,N_2823,N_3445);
and U4704 (N_4704,N_3551,N_3226);
nor U4705 (N_4705,N_3871,N_2581);
xnor U4706 (N_4706,N_2730,N_3089);
nand U4707 (N_4707,N_3902,N_3271);
nand U4708 (N_4708,N_2774,N_3504);
or U4709 (N_4709,N_2701,N_3243);
xor U4710 (N_4710,N_3019,N_3382);
xor U4711 (N_4711,N_3629,N_3700);
nand U4712 (N_4712,N_3102,N_2656);
nand U4713 (N_4713,N_3007,N_3520);
nor U4714 (N_4714,N_2230,N_3773);
nor U4715 (N_4715,N_2704,N_2450);
xor U4716 (N_4716,N_2258,N_3714);
nand U4717 (N_4717,N_3440,N_3268);
xor U4718 (N_4718,N_2655,N_2786);
nor U4719 (N_4719,N_2962,N_3230);
nor U4720 (N_4720,N_2775,N_2329);
xnor U4721 (N_4721,N_3624,N_2200);
and U4722 (N_4722,N_3892,N_3971);
xnor U4723 (N_4723,N_3768,N_3924);
or U4724 (N_4724,N_2576,N_3049);
or U4725 (N_4725,N_2879,N_2291);
xor U4726 (N_4726,N_2039,N_3379);
or U4727 (N_4727,N_2716,N_2477);
xor U4728 (N_4728,N_3292,N_3359);
and U4729 (N_4729,N_2755,N_3170);
xor U4730 (N_4730,N_3117,N_3025);
xnor U4731 (N_4731,N_2003,N_2865);
xor U4732 (N_4732,N_2132,N_3743);
nand U4733 (N_4733,N_3100,N_2457);
nor U4734 (N_4734,N_2893,N_2464);
xnor U4735 (N_4735,N_2583,N_3113);
nor U4736 (N_4736,N_2281,N_3081);
or U4737 (N_4737,N_3592,N_3648);
xor U4738 (N_4738,N_2880,N_2593);
and U4739 (N_4739,N_2588,N_3864);
nor U4740 (N_4740,N_3946,N_2684);
nor U4741 (N_4741,N_3291,N_2405);
nor U4742 (N_4742,N_2467,N_3208);
nand U4743 (N_4743,N_3375,N_3484);
nand U4744 (N_4744,N_2141,N_2493);
or U4745 (N_4745,N_2752,N_3967);
or U4746 (N_4746,N_3849,N_2100);
and U4747 (N_4747,N_2262,N_3212);
or U4748 (N_4748,N_3522,N_3175);
nand U4749 (N_4749,N_2495,N_2712);
or U4750 (N_4750,N_3311,N_3454);
or U4751 (N_4751,N_3707,N_2114);
or U4752 (N_4752,N_2460,N_2868);
and U4753 (N_4753,N_3869,N_2738);
nand U4754 (N_4754,N_3240,N_3001);
and U4755 (N_4755,N_2474,N_3096);
and U4756 (N_4756,N_2572,N_2787);
nor U4757 (N_4757,N_2804,N_3746);
nand U4758 (N_4758,N_3868,N_3550);
nor U4759 (N_4759,N_2634,N_2247);
nand U4760 (N_4760,N_2707,N_3106);
xor U4761 (N_4761,N_2825,N_2614);
xnor U4762 (N_4762,N_3791,N_2324);
xnor U4763 (N_4763,N_2760,N_3031);
xnor U4764 (N_4764,N_3655,N_3497);
and U4765 (N_4765,N_2199,N_2630);
xnor U4766 (N_4766,N_3617,N_3227);
and U4767 (N_4767,N_2517,N_2925);
and U4768 (N_4768,N_3116,N_3921);
xnor U4769 (N_4769,N_2177,N_3815);
nand U4770 (N_4770,N_2573,N_2047);
xnor U4771 (N_4771,N_2500,N_2283);
or U4772 (N_4772,N_3530,N_2204);
xnor U4773 (N_4773,N_3318,N_3119);
nand U4774 (N_4774,N_2149,N_2334);
xnor U4775 (N_4775,N_3653,N_3256);
or U4776 (N_4776,N_2218,N_2632);
or U4777 (N_4777,N_2082,N_2276);
xor U4778 (N_4778,N_2487,N_3853);
or U4779 (N_4779,N_2145,N_2679);
and U4780 (N_4780,N_3659,N_2661);
and U4781 (N_4781,N_2193,N_2485);
nor U4782 (N_4782,N_2622,N_3687);
xnor U4783 (N_4783,N_2269,N_3338);
and U4784 (N_4784,N_2653,N_2131);
and U4785 (N_4785,N_3620,N_3818);
or U4786 (N_4786,N_3740,N_3383);
nand U4787 (N_4787,N_2093,N_2566);
or U4788 (N_4788,N_3751,N_3191);
and U4789 (N_4789,N_3810,N_3588);
nor U4790 (N_4790,N_3064,N_3811);
nor U4791 (N_4791,N_3643,N_3758);
and U4792 (N_4792,N_2923,N_2998);
nor U4793 (N_4793,N_2403,N_3299);
xor U4794 (N_4794,N_2497,N_3973);
and U4795 (N_4795,N_2914,N_2599);
xnor U4796 (N_4796,N_3874,N_2146);
or U4797 (N_4797,N_3745,N_3395);
or U4798 (N_4798,N_3039,N_2028);
nor U4799 (N_4799,N_2555,N_2029);
nand U4800 (N_4800,N_2990,N_2336);
or U4801 (N_4801,N_2351,N_2898);
nor U4802 (N_4802,N_3369,N_2207);
and U4803 (N_4803,N_3115,N_2133);
or U4804 (N_4804,N_3310,N_2241);
nand U4805 (N_4805,N_3756,N_2529);
or U4806 (N_4806,N_2153,N_2372);
and U4807 (N_4807,N_3108,N_3247);
or U4808 (N_4808,N_2223,N_2627);
xor U4809 (N_4809,N_3304,N_3155);
nor U4810 (N_4810,N_2873,N_2446);
or U4811 (N_4811,N_2533,N_2415);
or U4812 (N_4812,N_2101,N_2853);
or U4813 (N_4813,N_3407,N_2792);
and U4814 (N_4814,N_2421,N_3091);
or U4815 (N_4815,N_3490,N_3685);
and U4816 (N_4816,N_3644,N_2253);
or U4817 (N_4817,N_2782,N_2221);
and U4818 (N_4818,N_2294,N_2150);
or U4819 (N_4819,N_3103,N_2178);
and U4820 (N_4820,N_2694,N_2575);
nand U4821 (N_4821,N_2620,N_2483);
nand U4822 (N_4822,N_2733,N_3507);
nor U4823 (N_4823,N_2561,N_3171);
nand U4824 (N_4824,N_2709,N_2284);
xor U4825 (N_4825,N_3087,N_3584);
or U4826 (N_4826,N_2428,N_2600);
nand U4827 (N_4827,N_2192,N_2531);
and U4828 (N_4828,N_3005,N_3646);
nor U4829 (N_4829,N_3368,N_3533);
and U4830 (N_4830,N_2901,N_3760);
nand U4831 (N_4831,N_2885,N_3950);
nor U4832 (N_4832,N_3691,N_2205);
xnor U4833 (N_4833,N_3429,N_2305);
nand U4834 (N_4834,N_3882,N_3837);
nor U4835 (N_4835,N_2452,N_2909);
nand U4836 (N_4836,N_2074,N_2740);
nor U4837 (N_4837,N_2538,N_2936);
nand U4838 (N_4838,N_2595,N_3345);
nand U4839 (N_4839,N_3156,N_2376);
nor U4840 (N_4840,N_3600,N_3035);
nand U4841 (N_4841,N_2596,N_3193);
xnor U4842 (N_4842,N_2176,N_2976);
xor U4843 (N_4843,N_3896,N_3157);
or U4844 (N_4844,N_3937,N_3969);
xnor U4845 (N_4845,N_3736,N_3578);
nor U4846 (N_4846,N_2827,N_2702);
nand U4847 (N_4847,N_2229,N_3927);
and U4848 (N_4848,N_2570,N_2826);
nand U4849 (N_4849,N_3795,N_3821);
nor U4850 (N_4850,N_2222,N_3801);
nand U4851 (N_4851,N_2103,N_2770);
or U4852 (N_4852,N_3022,N_2646);
nor U4853 (N_4853,N_2696,N_3133);
nor U4854 (N_4854,N_3928,N_2530);
nor U4855 (N_4855,N_2954,N_3174);
or U4856 (N_4856,N_3057,N_2164);
or U4857 (N_4857,N_3684,N_3323);
xnor U4858 (N_4858,N_2034,N_2355);
nand U4859 (N_4859,N_3879,N_3965);
nand U4860 (N_4860,N_2828,N_2972);
or U4861 (N_4861,N_2635,N_3855);
nor U4862 (N_4862,N_2144,N_3960);
and U4863 (N_4863,N_3702,N_3008);
nor U4864 (N_4864,N_2116,N_3738);
nor U4865 (N_4865,N_3453,N_3913);
or U4866 (N_4866,N_3514,N_3380);
nand U4867 (N_4867,N_2949,N_2271);
nor U4868 (N_4868,N_2162,N_3799);
xor U4869 (N_4869,N_2761,N_2287);
nor U4870 (N_4870,N_3875,N_3118);
xnor U4871 (N_4871,N_2102,N_2858);
and U4872 (N_4872,N_2603,N_2582);
nor U4873 (N_4873,N_2455,N_3424);
and U4874 (N_4874,N_2545,N_3470);
xnor U4875 (N_4875,N_3983,N_2397);
xor U4876 (N_4876,N_3775,N_3086);
or U4877 (N_4877,N_2780,N_3322);
nor U4878 (N_4878,N_3958,N_3602);
or U4879 (N_4879,N_3474,N_2791);
nor U4880 (N_4880,N_2699,N_2384);
or U4881 (N_4881,N_3783,N_2128);
xor U4882 (N_4882,N_2618,N_2523);
or U4883 (N_4883,N_3895,N_3957);
xor U4884 (N_4884,N_3084,N_2233);
nor U4885 (N_4885,N_2731,N_3580);
and U4886 (N_4886,N_3231,N_3940);
nor U4887 (N_4887,N_2577,N_3033);
or U4888 (N_4888,N_2433,N_2750);
or U4889 (N_4889,N_2010,N_2062);
and U4890 (N_4890,N_3263,N_3344);
and U4891 (N_4891,N_2111,N_2449);
or U4892 (N_4892,N_3391,N_2553);
and U4893 (N_4893,N_3589,N_3147);
nor U4894 (N_4894,N_3774,N_3789);
nand U4895 (N_4895,N_2640,N_3353);
xor U4896 (N_4896,N_3842,N_3186);
or U4897 (N_4897,N_3261,N_2856);
nand U4898 (N_4898,N_3845,N_2140);
nor U4899 (N_4899,N_2766,N_2231);
nand U4900 (N_4900,N_3820,N_3536);
xor U4901 (N_4901,N_3907,N_2950);
xnor U4902 (N_4902,N_2246,N_3093);
and U4903 (N_4903,N_2837,N_2304);
xnor U4904 (N_4904,N_2021,N_3706);
and U4905 (N_4905,N_3831,N_2905);
nor U4906 (N_4906,N_3194,N_3554);
nand U4907 (N_4907,N_3563,N_2175);
xnor U4908 (N_4908,N_2961,N_2906);
and U4909 (N_4909,N_2541,N_3238);
or U4910 (N_4910,N_2815,N_3562);
or U4911 (N_4911,N_3307,N_2396);
xnor U4912 (N_4912,N_3506,N_3919);
nor U4913 (N_4913,N_3640,N_3024);
and U4914 (N_4914,N_3364,N_2587);
xor U4915 (N_4915,N_3651,N_3272);
or U4916 (N_4916,N_3225,N_2732);
or U4917 (N_4917,N_2436,N_3670);
or U4918 (N_4918,N_3524,N_2432);
nor U4919 (N_4919,N_3542,N_3552);
xnor U4920 (N_4920,N_3716,N_3246);
nor U4921 (N_4921,N_2277,N_2159);
xor U4922 (N_4922,N_2850,N_3411);
and U4923 (N_4923,N_2303,N_3011);
xor U4924 (N_4924,N_2496,N_3073);
nor U4925 (N_4925,N_3647,N_3726);
and U4926 (N_4926,N_2585,N_3911);
or U4927 (N_4927,N_3130,N_3066);
nor U4928 (N_4928,N_3948,N_3482);
xnor U4929 (N_4929,N_2125,N_2685);
and U4930 (N_4930,N_3335,N_2417);
nand U4931 (N_4931,N_2499,N_3683);
and U4932 (N_4932,N_2902,N_2845);
and U4933 (N_4933,N_2490,N_2963);
nand U4934 (N_4934,N_2636,N_2723);
and U4935 (N_4935,N_2323,N_2965);
xor U4936 (N_4936,N_2606,N_2068);
or U4937 (N_4937,N_3388,N_3313);
or U4938 (N_4938,N_3348,N_3264);
and U4939 (N_4939,N_2266,N_2713);
or U4940 (N_4940,N_3515,N_3739);
nor U4941 (N_4941,N_2136,N_3813);
xnor U4942 (N_4942,N_3450,N_3021);
nand U4943 (N_4943,N_2462,N_3489);
nand U4944 (N_4944,N_3749,N_3072);
or U4945 (N_4945,N_2669,N_3114);
and U4946 (N_4946,N_2734,N_3244);
nand U4947 (N_4947,N_3404,N_2437);
nand U4948 (N_4948,N_3366,N_2565);
nand U4949 (N_4949,N_3565,N_2742);
nor U4950 (N_4950,N_2212,N_3806);
nor U4951 (N_4951,N_2979,N_3165);
or U4952 (N_4952,N_2569,N_3798);
nand U4953 (N_4953,N_2528,N_3254);
nand U4954 (N_4954,N_2939,N_3920);
xor U4955 (N_4955,N_2234,N_2044);
and U4956 (N_4956,N_3591,N_3088);
or U4957 (N_4957,N_3336,N_2981);
nand U4958 (N_4958,N_3267,N_3223);
xnor U4959 (N_4959,N_2049,N_3160);
xnor U4960 (N_4960,N_3734,N_3888);
and U4961 (N_4961,N_2031,N_2633);
nor U4962 (N_4962,N_2239,N_3314);
nor U4963 (N_4963,N_3635,N_2083);
nor U4964 (N_4964,N_2612,N_2534);
xor U4965 (N_4965,N_3503,N_3925);
nand U4966 (N_4966,N_2360,N_2345);
nand U4967 (N_4967,N_2007,N_3933);
nor U4968 (N_4968,N_2651,N_3728);
nand U4969 (N_4969,N_3926,N_2022);
nor U4970 (N_4970,N_3124,N_2941);
xor U4971 (N_4971,N_3808,N_3816);
xnor U4972 (N_4972,N_3678,N_2006);
or U4973 (N_4973,N_3409,N_2371);
xor U4974 (N_4974,N_2472,N_3224);
nand U4975 (N_4975,N_2299,N_3730);
nand U4976 (N_4976,N_3984,N_3439);
and U4977 (N_4977,N_2798,N_3206);
or U4978 (N_4978,N_3956,N_2870);
xnor U4979 (N_4979,N_3063,N_3188);
and U4980 (N_4980,N_3112,N_2244);
nor U4981 (N_4981,N_3701,N_3776);
nand U4982 (N_4982,N_2037,N_2995);
or U4983 (N_4983,N_3817,N_3521);
nand U4984 (N_4984,N_2097,N_2005);
xnor U4985 (N_4985,N_2960,N_2686);
nand U4986 (N_4986,N_3571,N_2776);
xnor U4987 (N_4987,N_3944,N_3213);
xnor U4988 (N_4988,N_3912,N_2876);
nor U4989 (N_4989,N_3553,N_2687);
xnor U4990 (N_4990,N_3665,N_2453);
and U4991 (N_4991,N_2542,N_2933);
and U4992 (N_4992,N_3312,N_3134);
xnor U4993 (N_4993,N_3579,N_2220);
xnor U4994 (N_4994,N_3495,N_2992);
nor U4995 (N_4995,N_3794,N_2383);
nor U4996 (N_4996,N_3986,N_2509);
nand U4997 (N_4997,N_3512,N_3953);
nor U4998 (N_4998,N_2228,N_2718);
and U4999 (N_4999,N_2328,N_3425);
or U5000 (N_5000,N_3814,N_3333);
nor U5001 (N_5001,N_2115,N_2808);
and U5002 (N_5002,N_2556,N_2046);
xor U5003 (N_5003,N_2956,N_3356);
or U5004 (N_5004,N_2375,N_3608);
and U5005 (N_5005,N_3011,N_2261);
xor U5006 (N_5006,N_2004,N_2859);
xnor U5007 (N_5007,N_3618,N_2709);
nor U5008 (N_5008,N_2719,N_3697);
nor U5009 (N_5009,N_2185,N_2149);
or U5010 (N_5010,N_2649,N_2422);
and U5011 (N_5011,N_2769,N_2632);
or U5012 (N_5012,N_2089,N_2124);
or U5013 (N_5013,N_3858,N_2476);
nor U5014 (N_5014,N_2991,N_3090);
xnor U5015 (N_5015,N_3486,N_3744);
xnor U5016 (N_5016,N_2100,N_2758);
xnor U5017 (N_5017,N_2231,N_2152);
xor U5018 (N_5018,N_2229,N_3337);
or U5019 (N_5019,N_3489,N_3699);
or U5020 (N_5020,N_3559,N_3428);
xor U5021 (N_5021,N_2912,N_2029);
or U5022 (N_5022,N_2809,N_2955);
nor U5023 (N_5023,N_2102,N_2764);
or U5024 (N_5024,N_3164,N_3416);
xor U5025 (N_5025,N_3899,N_2172);
or U5026 (N_5026,N_2257,N_2183);
xnor U5027 (N_5027,N_3488,N_2131);
and U5028 (N_5028,N_2396,N_2897);
and U5029 (N_5029,N_2367,N_2396);
nand U5030 (N_5030,N_2170,N_2831);
nand U5031 (N_5031,N_3062,N_3884);
nor U5032 (N_5032,N_3851,N_2742);
or U5033 (N_5033,N_2331,N_2964);
nor U5034 (N_5034,N_3158,N_2623);
and U5035 (N_5035,N_3574,N_3290);
and U5036 (N_5036,N_2130,N_3795);
xor U5037 (N_5037,N_3390,N_2367);
xor U5038 (N_5038,N_3273,N_2767);
or U5039 (N_5039,N_3706,N_2579);
xnor U5040 (N_5040,N_3338,N_3892);
nor U5041 (N_5041,N_2861,N_3553);
nor U5042 (N_5042,N_3499,N_3403);
xnor U5043 (N_5043,N_2594,N_3693);
nor U5044 (N_5044,N_2167,N_2806);
xnor U5045 (N_5045,N_2125,N_3888);
or U5046 (N_5046,N_3468,N_3867);
and U5047 (N_5047,N_3061,N_3724);
xor U5048 (N_5048,N_3330,N_2241);
xor U5049 (N_5049,N_3773,N_2683);
nor U5050 (N_5050,N_2053,N_2729);
or U5051 (N_5051,N_2594,N_2425);
xnor U5052 (N_5052,N_2926,N_3672);
nor U5053 (N_5053,N_2948,N_3263);
nand U5054 (N_5054,N_2592,N_2254);
xnor U5055 (N_5055,N_3501,N_3634);
nor U5056 (N_5056,N_2479,N_3810);
xnor U5057 (N_5057,N_2028,N_3116);
xnor U5058 (N_5058,N_3798,N_2775);
nor U5059 (N_5059,N_2755,N_3129);
and U5060 (N_5060,N_3898,N_3057);
and U5061 (N_5061,N_2178,N_3106);
or U5062 (N_5062,N_2193,N_3017);
nand U5063 (N_5063,N_2893,N_2896);
nand U5064 (N_5064,N_3908,N_2705);
or U5065 (N_5065,N_2044,N_3923);
or U5066 (N_5066,N_2089,N_3038);
and U5067 (N_5067,N_3874,N_3970);
nand U5068 (N_5068,N_3214,N_2221);
and U5069 (N_5069,N_2149,N_3455);
xor U5070 (N_5070,N_2304,N_3282);
nor U5071 (N_5071,N_3307,N_3686);
or U5072 (N_5072,N_3455,N_3203);
or U5073 (N_5073,N_2817,N_2792);
xor U5074 (N_5074,N_3063,N_2532);
xnor U5075 (N_5075,N_3419,N_3444);
or U5076 (N_5076,N_3419,N_3344);
or U5077 (N_5077,N_2591,N_2431);
xor U5078 (N_5078,N_3097,N_2515);
nor U5079 (N_5079,N_2981,N_2882);
nand U5080 (N_5080,N_3512,N_2492);
nand U5081 (N_5081,N_2359,N_2744);
nor U5082 (N_5082,N_2231,N_2851);
nor U5083 (N_5083,N_2941,N_3351);
nand U5084 (N_5084,N_2641,N_3474);
nor U5085 (N_5085,N_3805,N_3810);
nand U5086 (N_5086,N_2826,N_2600);
or U5087 (N_5087,N_2610,N_2589);
nor U5088 (N_5088,N_3741,N_2077);
and U5089 (N_5089,N_3043,N_2279);
xnor U5090 (N_5090,N_2878,N_2949);
nor U5091 (N_5091,N_2728,N_2055);
xnor U5092 (N_5092,N_3017,N_2482);
xor U5093 (N_5093,N_2342,N_2925);
nor U5094 (N_5094,N_2028,N_3593);
or U5095 (N_5095,N_3029,N_3333);
xnor U5096 (N_5096,N_2343,N_3255);
nand U5097 (N_5097,N_2670,N_2783);
and U5098 (N_5098,N_2073,N_2543);
or U5099 (N_5099,N_2805,N_3949);
and U5100 (N_5100,N_3219,N_2574);
nor U5101 (N_5101,N_3701,N_3617);
nor U5102 (N_5102,N_2695,N_3860);
or U5103 (N_5103,N_3224,N_3291);
and U5104 (N_5104,N_2077,N_2247);
xor U5105 (N_5105,N_3271,N_3807);
nand U5106 (N_5106,N_3954,N_2948);
nor U5107 (N_5107,N_3095,N_3832);
and U5108 (N_5108,N_2599,N_2035);
nor U5109 (N_5109,N_2563,N_2669);
and U5110 (N_5110,N_2538,N_3494);
and U5111 (N_5111,N_2695,N_3098);
nand U5112 (N_5112,N_2637,N_2444);
nand U5113 (N_5113,N_3568,N_2669);
nand U5114 (N_5114,N_2267,N_3943);
nor U5115 (N_5115,N_2133,N_3427);
nand U5116 (N_5116,N_3313,N_2931);
or U5117 (N_5117,N_2845,N_2840);
nor U5118 (N_5118,N_3912,N_3904);
or U5119 (N_5119,N_3555,N_3865);
xnor U5120 (N_5120,N_2852,N_3405);
or U5121 (N_5121,N_3711,N_3515);
nor U5122 (N_5122,N_3203,N_3584);
nor U5123 (N_5123,N_3067,N_3645);
nor U5124 (N_5124,N_3134,N_2895);
nand U5125 (N_5125,N_2772,N_3312);
xnor U5126 (N_5126,N_2981,N_2194);
and U5127 (N_5127,N_2085,N_3018);
nand U5128 (N_5128,N_3252,N_2840);
or U5129 (N_5129,N_3393,N_3252);
xnor U5130 (N_5130,N_3282,N_2578);
nor U5131 (N_5131,N_2679,N_3362);
and U5132 (N_5132,N_2197,N_2465);
nor U5133 (N_5133,N_2761,N_3589);
or U5134 (N_5134,N_2119,N_2713);
xnor U5135 (N_5135,N_3920,N_3294);
and U5136 (N_5136,N_2511,N_3976);
nand U5137 (N_5137,N_3606,N_2105);
and U5138 (N_5138,N_2402,N_2828);
or U5139 (N_5139,N_3108,N_3003);
nand U5140 (N_5140,N_3912,N_3670);
xor U5141 (N_5141,N_3594,N_3946);
nand U5142 (N_5142,N_3783,N_2840);
xnor U5143 (N_5143,N_3074,N_2686);
or U5144 (N_5144,N_3872,N_2408);
or U5145 (N_5145,N_2994,N_2035);
and U5146 (N_5146,N_3096,N_2904);
nand U5147 (N_5147,N_2000,N_2426);
and U5148 (N_5148,N_3299,N_3221);
and U5149 (N_5149,N_3653,N_2278);
or U5150 (N_5150,N_3123,N_2280);
and U5151 (N_5151,N_3423,N_2985);
or U5152 (N_5152,N_2112,N_3336);
nand U5153 (N_5153,N_2850,N_2183);
or U5154 (N_5154,N_2514,N_3508);
xnor U5155 (N_5155,N_2824,N_3705);
xor U5156 (N_5156,N_2553,N_2437);
nor U5157 (N_5157,N_3993,N_3384);
nand U5158 (N_5158,N_2448,N_3900);
nor U5159 (N_5159,N_2022,N_2819);
nand U5160 (N_5160,N_3722,N_2779);
nand U5161 (N_5161,N_2104,N_3197);
xor U5162 (N_5162,N_2308,N_3153);
nand U5163 (N_5163,N_2153,N_3571);
xor U5164 (N_5164,N_2080,N_2617);
nor U5165 (N_5165,N_2807,N_3466);
xnor U5166 (N_5166,N_2460,N_3909);
or U5167 (N_5167,N_3719,N_3192);
xor U5168 (N_5168,N_2702,N_2639);
and U5169 (N_5169,N_2432,N_2752);
nor U5170 (N_5170,N_3772,N_2911);
xor U5171 (N_5171,N_3075,N_3403);
xor U5172 (N_5172,N_3336,N_2452);
xor U5173 (N_5173,N_3792,N_2362);
or U5174 (N_5174,N_3406,N_2385);
and U5175 (N_5175,N_3275,N_2957);
and U5176 (N_5176,N_3057,N_3551);
nand U5177 (N_5177,N_3168,N_3326);
nand U5178 (N_5178,N_2980,N_3761);
or U5179 (N_5179,N_3787,N_3154);
and U5180 (N_5180,N_2461,N_2281);
nand U5181 (N_5181,N_2406,N_2419);
and U5182 (N_5182,N_3388,N_2352);
nor U5183 (N_5183,N_3098,N_2369);
nor U5184 (N_5184,N_2768,N_3724);
and U5185 (N_5185,N_3598,N_2753);
and U5186 (N_5186,N_2893,N_3787);
and U5187 (N_5187,N_2157,N_3330);
or U5188 (N_5188,N_3010,N_3636);
nand U5189 (N_5189,N_3192,N_3236);
xor U5190 (N_5190,N_2933,N_3422);
and U5191 (N_5191,N_3641,N_3588);
and U5192 (N_5192,N_3847,N_2250);
xnor U5193 (N_5193,N_2865,N_3762);
and U5194 (N_5194,N_3052,N_2721);
xor U5195 (N_5195,N_3477,N_3307);
xor U5196 (N_5196,N_3521,N_3364);
or U5197 (N_5197,N_2185,N_3878);
and U5198 (N_5198,N_2519,N_3701);
xor U5199 (N_5199,N_2886,N_2252);
nor U5200 (N_5200,N_3100,N_2942);
and U5201 (N_5201,N_2547,N_2224);
and U5202 (N_5202,N_3020,N_3532);
or U5203 (N_5203,N_2116,N_2095);
nor U5204 (N_5204,N_3006,N_2716);
nor U5205 (N_5205,N_3522,N_3788);
or U5206 (N_5206,N_2403,N_3105);
and U5207 (N_5207,N_3237,N_3147);
or U5208 (N_5208,N_2228,N_2999);
nor U5209 (N_5209,N_3561,N_2952);
and U5210 (N_5210,N_2863,N_2149);
nor U5211 (N_5211,N_2257,N_3082);
xnor U5212 (N_5212,N_2133,N_2604);
and U5213 (N_5213,N_3362,N_3956);
nand U5214 (N_5214,N_2340,N_2589);
or U5215 (N_5215,N_3075,N_2246);
nand U5216 (N_5216,N_2359,N_2763);
nor U5217 (N_5217,N_2472,N_2438);
nand U5218 (N_5218,N_3531,N_2095);
nand U5219 (N_5219,N_3406,N_2639);
nor U5220 (N_5220,N_3923,N_3498);
and U5221 (N_5221,N_3055,N_2437);
xor U5222 (N_5222,N_3810,N_3042);
and U5223 (N_5223,N_3495,N_3386);
nand U5224 (N_5224,N_2231,N_3290);
and U5225 (N_5225,N_3779,N_2104);
nand U5226 (N_5226,N_3132,N_3670);
xor U5227 (N_5227,N_3468,N_3193);
xnor U5228 (N_5228,N_2209,N_3547);
and U5229 (N_5229,N_2458,N_3139);
nand U5230 (N_5230,N_3826,N_3046);
xnor U5231 (N_5231,N_2210,N_3319);
nand U5232 (N_5232,N_2321,N_2151);
xnor U5233 (N_5233,N_2170,N_3595);
nor U5234 (N_5234,N_3053,N_3079);
xor U5235 (N_5235,N_2509,N_2695);
nand U5236 (N_5236,N_2689,N_2729);
nor U5237 (N_5237,N_3677,N_3095);
and U5238 (N_5238,N_2318,N_3780);
nor U5239 (N_5239,N_2099,N_3839);
xor U5240 (N_5240,N_2462,N_2670);
nand U5241 (N_5241,N_2013,N_2924);
xnor U5242 (N_5242,N_3372,N_2251);
xnor U5243 (N_5243,N_2411,N_2936);
nand U5244 (N_5244,N_3421,N_2838);
nand U5245 (N_5245,N_2245,N_3527);
nor U5246 (N_5246,N_3584,N_2556);
nand U5247 (N_5247,N_2684,N_2490);
xnor U5248 (N_5248,N_3305,N_3118);
or U5249 (N_5249,N_3057,N_2660);
or U5250 (N_5250,N_3407,N_2952);
nand U5251 (N_5251,N_3339,N_3220);
and U5252 (N_5252,N_3985,N_3840);
xor U5253 (N_5253,N_3425,N_2469);
and U5254 (N_5254,N_2706,N_2905);
and U5255 (N_5255,N_2794,N_3471);
nand U5256 (N_5256,N_3115,N_3285);
xor U5257 (N_5257,N_3574,N_3045);
nor U5258 (N_5258,N_2730,N_2057);
nand U5259 (N_5259,N_3276,N_3174);
nand U5260 (N_5260,N_2500,N_3320);
or U5261 (N_5261,N_3465,N_2409);
xor U5262 (N_5262,N_3322,N_2821);
or U5263 (N_5263,N_3782,N_2964);
xor U5264 (N_5264,N_2272,N_2671);
or U5265 (N_5265,N_2956,N_3396);
nor U5266 (N_5266,N_3771,N_3366);
nand U5267 (N_5267,N_3754,N_3978);
xnor U5268 (N_5268,N_2021,N_2290);
nand U5269 (N_5269,N_2780,N_3506);
nand U5270 (N_5270,N_2397,N_2140);
and U5271 (N_5271,N_3962,N_3446);
or U5272 (N_5272,N_3265,N_2197);
and U5273 (N_5273,N_3944,N_3011);
nand U5274 (N_5274,N_3172,N_2964);
and U5275 (N_5275,N_3531,N_2791);
or U5276 (N_5276,N_3739,N_2980);
nand U5277 (N_5277,N_2707,N_2875);
or U5278 (N_5278,N_3755,N_2664);
and U5279 (N_5279,N_3491,N_3075);
or U5280 (N_5280,N_3310,N_2786);
or U5281 (N_5281,N_3840,N_3704);
and U5282 (N_5282,N_3285,N_3766);
nor U5283 (N_5283,N_3787,N_2334);
nand U5284 (N_5284,N_2649,N_2258);
xor U5285 (N_5285,N_2969,N_3772);
xnor U5286 (N_5286,N_3738,N_2403);
or U5287 (N_5287,N_2010,N_2596);
and U5288 (N_5288,N_3335,N_3547);
nor U5289 (N_5289,N_2696,N_3523);
nor U5290 (N_5290,N_2865,N_3436);
and U5291 (N_5291,N_3554,N_3074);
xor U5292 (N_5292,N_3634,N_3060);
nand U5293 (N_5293,N_2148,N_3685);
nand U5294 (N_5294,N_3754,N_2343);
and U5295 (N_5295,N_2834,N_2729);
xor U5296 (N_5296,N_3469,N_3291);
xnor U5297 (N_5297,N_3882,N_2133);
nor U5298 (N_5298,N_3149,N_2256);
nor U5299 (N_5299,N_2313,N_2388);
xnor U5300 (N_5300,N_3741,N_2694);
nand U5301 (N_5301,N_3921,N_2211);
nand U5302 (N_5302,N_3588,N_3530);
nor U5303 (N_5303,N_2626,N_3764);
nor U5304 (N_5304,N_3699,N_3653);
nor U5305 (N_5305,N_3866,N_3930);
nor U5306 (N_5306,N_2243,N_3883);
nand U5307 (N_5307,N_3835,N_3476);
xnor U5308 (N_5308,N_3644,N_3091);
nand U5309 (N_5309,N_3927,N_3839);
or U5310 (N_5310,N_3881,N_2019);
nand U5311 (N_5311,N_3805,N_2953);
or U5312 (N_5312,N_2799,N_2631);
or U5313 (N_5313,N_3349,N_3435);
or U5314 (N_5314,N_3776,N_2187);
or U5315 (N_5315,N_3602,N_3033);
nand U5316 (N_5316,N_2807,N_3600);
or U5317 (N_5317,N_3949,N_3564);
nand U5318 (N_5318,N_2646,N_2961);
or U5319 (N_5319,N_2314,N_2244);
xor U5320 (N_5320,N_3474,N_2044);
nand U5321 (N_5321,N_3550,N_2778);
and U5322 (N_5322,N_3287,N_3313);
and U5323 (N_5323,N_2561,N_3603);
or U5324 (N_5324,N_2571,N_3221);
nand U5325 (N_5325,N_2771,N_3862);
nand U5326 (N_5326,N_2967,N_3726);
or U5327 (N_5327,N_3276,N_2081);
xnor U5328 (N_5328,N_3022,N_2550);
nor U5329 (N_5329,N_2761,N_2572);
or U5330 (N_5330,N_2854,N_3287);
and U5331 (N_5331,N_2268,N_2100);
nand U5332 (N_5332,N_3884,N_3633);
or U5333 (N_5333,N_2504,N_2656);
nand U5334 (N_5334,N_3932,N_3666);
nor U5335 (N_5335,N_2274,N_3107);
and U5336 (N_5336,N_3032,N_3280);
nand U5337 (N_5337,N_2877,N_2002);
nand U5338 (N_5338,N_2864,N_3371);
xor U5339 (N_5339,N_2567,N_2310);
nor U5340 (N_5340,N_3030,N_2786);
xor U5341 (N_5341,N_3363,N_2677);
nor U5342 (N_5342,N_3279,N_2272);
nor U5343 (N_5343,N_2455,N_3332);
nor U5344 (N_5344,N_3155,N_2858);
nand U5345 (N_5345,N_3231,N_2502);
xnor U5346 (N_5346,N_2939,N_3934);
nor U5347 (N_5347,N_2358,N_2102);
or U5348 (N_5348,N_2005,N_2911);
nor U5349 (N_5349,N_3509,N_3639);
nor U5350 (N_5350,N_3027,N_3821);
and U5351 (N_5351,N_3991,N_2221);
and U5352 (N_5352,N_3131,N_2078);
or U5353 (N_5353,N_2766,N_2233);
nor U5354 (N_5354,N_2768,N_2157);
and U5355 (N_5355,N_2390,N_2822);
nand U5356 (N_5356,N_3909,N_2316);
nand U5357 (N_5357,N_2381,N_2907);
or U5358 (N_5358,N_2986,N_2057);
nand U5359 (N_5359,N_2674,N_2128);
nand U5360 (N_5360,N_2512,N_2454);
nand U5361 (N_5361,N_2312,N_2747);
nand U5362 (N_5362,N_3947,N_2901);
xor U5363 (N_5363,N_3099,N_2266);
nand U5364 (N_5364,N_3743,N_3025);
and U5365 (N_5365,N_3966,N_2620);
nand U5366 (N_5366,N_2260,N_2313);
nand U5367 (N_5367,N_3256,N_2553);
and U5368 (N_5368,N_2330,N_2574);
and U5369 (N_5369,N_2857,N_2248);
and U5370 (N_5370,N_2103,N_3372);
and U5371 (N_5371,N_2140,N_2841);
nand U5372 (N_5372,N_2485,N_2159);
nand U5373 (N_5373,N_2495,N_2397);
and U5374 (N_5374,N_3914,N_2465);
xor U5375 (N_5375,N_2706,N_3656);
nand U5376 (N_5376,N_3294,N_3181);
or U5377 (N_5377,N_3500,N_2854);
and U5378 (N_5378,N_3959,N_2699);
and U5379 (N_5379,N_2811,N_3368);
nand U5380 (N_5380,N_2537,N_2112);
nand U5381 (N_5381,N_2211,N_2451);
nor U5382 (N_5382,N_2634,N_2608);
or U5383 (N_5383,N_3540,N_3725);
or U5384 (N_5384,N_2385,N_3756);
nor U5385 (N_5385,N_2925,N_2500);
or U5386 (N_5386,N_2192,N_3217);
nor U5387 (N_5387,N_2136,N_2528);
xor U5388 (N_5388,N_3349,N_2018);
and U5389 (N_5389,N_2921,N_3682);
xnor U5390 (N_5390,N_2913,N_2015);
nor U5391 (N_5391,N_3627,N_2839);
nor U5392 (N_5392,N_3514,N_3609);
nand U5393 (N_5393,N_2211,N_3020);
nand U5394 (N_5394,N_2507,N_2464);
nor U5395 (N_5395,N_3862,N_2175);
xor U5396 (N_5396,N_3410,N_3249);
and U5397 (N_5397,N_2204,N_2081);
xnor U5398 (N_5398,N_2942,N_3370);
xor U5399 (N_5399,N_2545,N_3512);
or U5400 (N_5400,N_2805,N_3968);
nor U5401 (N_5401,N_3794,N_2508);
nand U5402 (N_5402,N_3213,N_3767);
nand U5403 (N_5403,N_3244,N_2660);
and U5404 (N_5404,N_3510,N_3227);
nor U5405 (N_5405,N_3918,N_3766);
and U5406 (N_5406,N_2092,N_2314);
and U5407 (N_5407,N_3471,N_2927);
and U5408 (N_5408,N_3215,N_3322);
and U5409 (N_5409,N_2571,N_2529);
or U5410 (N_5410,N_3782,N_3525);
xnor U5411 (N_5411,N_2010,N_3949);
nand U5412 (N_5412,N_2913,N_2476);
nand U5413 (N_5413,N_2586,N_2042);
and U5414 (N_5414,N_3826,N_3080);
nor U5415 (N_5415,N_3272,N_2158);
or U5416 (N_5416,N_3525,N_2175);
or U5417 (N_5417,N_3155,N_2983);
nand U5418 (N_5418,N_2244,N_2921);
nand U5419 (N_5419,N_3223,N_3085);
xor U5420 (N_5420,N_2843,N_2370);
and U5421 (N_5421,N_3215,N_2085);
or U5422 (N_5422,N_2760,N_3384);
nor U5423 (N_5423,N_3155,N_2397);
or U5424 (N_5424,N_3728,N_2207);
nand U5425 (N_5425,N_3407,N_2098);
or U5426 (N_5426,N_3973,N_3178);
and U5427 (N_5427,N_2634,N_3438);
nand U5428 (N_5428,N_2360,N_3239);
xnor U5429 (N_5429,N_3323,N_3480);
and U5430 (N_5430,N_2261,N_3392);
or U5431 (N_5431,N_2576,N_2297);
nor U5432 (N_5432,N_2693,N_2644);
nand U5433 (N_5433,N_2767,N_2341);
nor U5434 (N_5434,N_2377,N_3208);
or U5435 (N_5435,N_2799,N_3149);
xor U5436 (N_5436,N_2192,N_2294);
xor U5437 (N_5437,N_2104,N_3492);
xor U5438 (N_5438,N_3264,N_2328);
and U5439 (N_5439,N_3341,N_2646);
and U5440 (N_5440,N_3261,N_2921);
xnor U5441 (N_5441,N_3659,N_2429);
or U5442 (N_5442,N_3577,N_3594);
nor U5443 (N_5443,N_2010,N_2919);
xnor U5444 (N_5444,N_3861,N_2526);
xor U5445 (N_5445,N_2762,N_2020);
xor U5446 (N_5446,N_3049,N_2071);
nor U5447 (N_5447,N_2035,N_2749);
nor U5448 (N_5448,N_3316,N_2856);
or U5449 (N_5449,N_3335,N_3984);
or U5450 (N_5450,N_2062,N_2636);
nor U5451 (N_5451,N_2328,N_2521);
nor U5452 (N_5452,N_2170,N_2147);
or U5453 (N_5453,N_2036,N_3488);
xor U5454 (N_5454,N_2154,N_3859);
nor U5455 (N_5455,N_3519,N_3255);
and U5456 (N_5456,N_2860,N_2155);
or U5457 (N_5457,N_2196,N_2031);
nand U5458 (N_5458,N_3376,N_3587);
xor U5459 (N_5459,N_3674,N_2043);
nor U5460 (N_5460,N_3342,N_2731);
or U5461 (N_5461,N_2501,N_3780);
or U5462 (N_5462,N_2799,N_3318);
or U5463 (N_5463,N_3620,N_3753);
nand U5464 (N_5464,N_3539,N_3479);
and U5465 (N_5465,N_3013,N_2351);
nor U5466 (N_5466,N_2232,N_3008);
xnor U5467 (N_5467,N_3200,N_3930);
or U5468 (N_5468,N_2781,N_3146);
and U5469 (N_5469,N_2520,N_2295);
xnor U5470 (N_5470,N_3274,N_2353);
xor U5471 (N_5471,N_3038,N_2168);
nand U5472 (N_5472,N_2217,N_3741);
nor U5473 (N_5473,N_2330,N_3114);
nor U5474 (N_5474,N_2075,N_3597);
nand U5475 (N_5475,N_3931,N_3604);
and U5476 (N_5476,N_2782,N_3772);
nand U5477 (N_5477,N_3740,N_2838);
nand U5478 (N_5478,N_3606,N_3707);
nand U5479 (N_5479,N_2333,N_2233);
nand U5480 (N_5480,N_3107,N_2172);
or U5481 (N_5481,N_3970,N_2999);
nand U5482 (N_5482,N_3557,N_3701);
and U5483 (N_5483,N_2895,N_3102);
nand U5484 (N_5484,N_3046,N_3191);
and U5485 (N_5485,N_3596,N_3913);
xor U5486 (N_5486,N_2621,N_3197);
nor U5487 (N_5487,N_3317,N_2505);
or U5488 (N_5488,N_2919,N_2130);
xnor U5489 (N_5489,N_3372,N_3139);
nor U5490 (N_5490,N_3967,N_2685);
nand U5491 (N_5491,N_2761,N_2664);
nor U5492 (N_5492,N_2641,N_3267);
and U5493 (N_5493,N_2994,N_3103);
xor U5494 (N_5494,N_3143,N_3782);
xor U5495 (N_5495,N_2301,N_3191);
nand U5496 (N_5496,N_3812,N_2915);
and U5497 (N_5497,N_2697,N_2972);
xor U5498 (N_5498,N_3634,N_2798);
xnor U5499 (N_5499,N_3279,N_3881);
or U5500 (N_5500,N_3096,N_2658);
xnor U5501 (N_5501,N_3915,N_2740);
and U5502 (N_5502,N_3009,N_2790);
nor U5503 (N_5503,N_3408,N_3319);
xnor U5504 (N_5504,N_3019,N_3102);
xor U5505 (N_5505,N_3289,N_2232);
xnor U5506 (N_5506,N_2440,N_2134);
nand U5507 (N_5507,N_2902,N_3877);
xor U5508 (N_5508,N_3788,N_2343);
nor U5509 (N_5509,N_3714,N_3282);
or U5510 (N_5510,N_3619,N_3612);
nor U5511 (N_5511,N_3962,N_3501);
xnor U5512 (N_5512,N_3827,N_2277);
xnor U5513 (N_5513,N_3784,N_3930);
nand U5514 (N_5514,N_2935,N_2246);
nand U5515 (N_5515,N_3216,N_2985);
nor U5516 (N_5516,N_2136,N_2686);
xor U5517 (N_5517,N_3051,N_3263);
nand U5518 (N_5518,N_2855,N_3260);
nand U5519 (N_5519,N_2693,N_3119);
xnor U5520 (N_5520,N_3994,N_3213);
nand U5521 (N_5521,N_3619,N_3168);
nor U5522 (N_5522,N_2383,N_2765);
and U5523 (N_5523,N_2755,N_2423);
or U5524 (N_5524,N_2133,N_3420);
nor U5525 (N_5525,N_2183,N_3361);
nor U5526 (N_5526,N_3662,N_2826);
nand U5527 (N_5527,N_3914,N_3464);
and U5528 (N_5528,N_2496,N_2678);
xnor U5529 (N_5529,N_2687,N_2429);
xnor U5530 (N_5530,N_2611,N_2580);
nand U5531 (N_5531,N_3282,N_2828);
and U5532 (N_5532,N_3121,N_3872);
and U5533 (N_5533,N_3381,N_2422);
or U5534 (N_5534,N_3183,N_2516);
or U5535 (N_5535,N_2572,N_2427);
and U5536 (N_5536,N_2627,N_3301);
and U5537 (N_5537,N_3270,N_3835);
xor U5538 (N_5538,N_3409,N_2389);
nand U5539 (N_5539,N_2986,N_3506);
nand U5540 (N_5540,N_2475,N_3539);
or U5541 (N_5541,N_2915,N_2893);
and U5542 (N_5542,N_2935,N_2946);
or U5543 (N_5543,N_3245,N_3557);
and U5544 (N_5544,N_3163,N_2780);
nand U5545 (N_5545,N_3699,N_2351);
xor U5546 (N_5546,N_2435,N_3422);
nor U5547 (N_5547,N_2911,N_2872);
and U5548 (N_5548,N_3394,N_2936);
xor U5549 (N_5549,N_2337,N_3895);
nor U5550 (N_5550,N_3687,N_3305);
or U5551 (N_5551,N_3875,N_3033);
and U5552 (N_5552,N_2213,N_2588);
and U5553 (N_5553,N_2686,N_2443);
and U5554 (N_5554,N_3263,N_2466);
and U5555 (N_5555,N_2919,N_3654);
or U5556 (N_5556,N_3631,N_3475);
nand U5557 (N_5557,N_3973,N_2135);
xor U5558 (N_5558,N_3948,N_2512);
nor U5559 (N_5559,N_2075,N_3544);
or U5560 (N_5560,N_3227,N_2379);
nor U5561 (N_5561,N_2698,N_3672);
nor U5562 (N_5562,N_2356,N_2446);
or U5563 (N_5563,N_2806,N_2098);
nand U5564 (N_5564,N_2321,N_3779);
xnor U5565 (N_5565,N_2314,N_2236);
or U5566 (N_5566,N_3626,N_2041);
xnor U5567 (N_5567,N_2335,N_3417);
nand U5568 (N_5568,N_2367,N_3322);
xnor U5569 (N_5569,N_2205,N_2960);
xnor U5570 (N_5570,N_3504,N_2343);
xor U5571 (N_5571,N_3391,N_3269);
xor U5572 (N_5572,N_3982,N_2941);
xor U5573 (N_5573,N_3417,N_3511);
and U5574 (N_5574,N_2928,N_2117);
nor U5575 (N_5575,N_2644,N_3397);
nor U5576 (N_5576,N_2390,N_2664);
nand U5577 (N_5577,N_2793,N_3348);
or U5578 (N_5578,N_2703,N_2022);
nand U5579 (N_5579,N_2535,N_2720);
xnor U5580 (N_5580,N_3382,N_2853);
or U5581 (N_5581,N_2459,N_2798);
or U5582 (N_5582,N_2794,N_2090);
nor U5583 (N_5583,N_3728,N_2543);
or U5584 (N_5584,N_2997,N_2657);
nand U5585 (N_5585,N_2052,N_2510);
nand U5586 (N_5586,N_3323,N_2530);
and U5587 (N_5587,N_2182,N_3785);
nand U5588 (N_5588,N_2289,N_3239);
xnor U5589 (N_5589,N_3596,N_3389);
xor U5590 (N_5590,N_3387,N_2134);
nand U5591 (N_5591,N_2769,N_3759);
nand U5592 (N_5592,N_3801,N_3196);
nor U5593 (N_5593,N_3110,N_2953);
nor U5594 (N_5594,N_2725,N_3529);
and U5595 (N_5595,N_3782,N_2626);
xor U5596 (N_5596,N_2920,N_3703);
and U5597 (N_5597,N_2054,N_3871);
or U5598 (N_5598,N_2147,N_3699);
or U5599 (N_5599,N_2800,N_2547);
nor U5600 (N_5600,N_2253,N_3151);
and U5601 (N_5601,N_2279,N_3886);
xor U5602 (N_5602,N_2821,N_3265);
xor U5603 (N_5603,N_2382,N_3272);
nor U5604 (N_5604,N_3981,N_2462);
or U5605 (N_5605,N_3132,N_3852);
nor U5606 (N_5606,N_3290,N_2972);
and U5607 (N_5607,N_3176,N_2909);
nor U5608 (N_5608,N_3586,N_2735);
nor U5609 (N_5609,N_2675,N_3852);
and U5610 (N_5610,N_3117,N_3532);
nor U5611 (N_5611,N_3666,N_2958);
nor U5612 (N_5612,N_3444,N_2198);
or U5613 (N_5613,N_3943,N_3984);
nor U5614 (N_5614,N_3971,N_3645);
and U5615 (N_5615,N_3494,N_3406);
nor U5616 (N_5616,N_3735,N_2771);
and U5617 (N_5617,N_3479,N_2724);
and U5618 (N_5618,N_3527,N_3081);
and U5619 (N_5619,N_2104,N_3399);
and U5620 (N_5620,N_2561,N_3738);
xor U5621 (N_5621,N_3568,N_3705);
and U5622 (N_5622,N_2396,N_2682);
xnor U5623 (N_5623,N_3525,N_3597);
and U5624 (N_5624,N_2684,N_3688);
nand U5625 (N_5625,N_3539,N_3554);
or U5626 (N_5626,N_2183,N_2992);
and U5627 (N_5627,N_2165,N_2840);
nand U5628 (N_5628,N_3600,N_2936);
and U5629 (N_5629,N_2237,N_3746);
and U5630 (N_5630,N_3098,N_2452);
and U5631 (N_5631,N_3635,N_3763);
and U5632 (N_5632,N_3862,N_2544);
nor U5633 (N_5633,N_3069,N_3172);
nor U5634 (N_5634,N_2223,N_2966);
or U5635 (N_5635,N_3492,N_2941);
and U5636 (N_5636,N_2889,N_2505);
nor U5637 (N_5637,N_3499,N_2733);
and U5638 (N_5638,N_3400,N_2110);
or U5639 (N_5639,N_3375,N_3411);
nand U5640 (N_5640,N_3324,N_2831);
nand U5641 (N_5641,N_3643,N_3376);
and U5642 (N_5642,N_3534,N_2826);
nand U5643 (N_5643,N_3890,N_2273);
nor U5644 (N_5644,N_3323,N_2910);
xor U5645 (N_5645,N_2535,N_2763);
nor U5646 (N_5646,N_3095,N_3325);
xor U5647 (N_5647,N_2717,N_3961);
nor U5648 (N_5648,N_3704,N_2673);
xor U5649 (N_5649,N_3819,N_3732);
nand U5650 (N_5650,N_2949,N_3615);
and U5651 (N_5651,N_3514,N_2871);
nand U5652 (N_5652,N_3405,N_2608);
nand U5653 (N_5653,N_3243,N_2622);
nor U5654 (N_5654,N_3753,N_2985);
or U5655 (N_5655,N_2300,N_3798);
or U5656 (N_5656,N_3205,N_2634);
xnor U5657 (N_5657,N_3762,N_2786);
xor U5658 (N_5658,N_2076,N_3540);
and U5659 (N_5659,N_2589,N_2313);
and U5660 (N_5660,N_2737,N_2741);
nand U5661 (N_5661,N_3237,N_3141);
and U5662 (N_5662,N_3081,N_3348);
nor U5663 (N_5663,N_3870,N_3119);
nor U5664 (N_5664,N_3952,N_2947);
nor U5665 (N_5665,N_3234,N_3378);
and U5666 (N_5666,N_2222,N_2465);
xnor U5667 (N_5667,N_3669,N_3595);
xnor U5668 (N_5668,N_2352,N_3793);
nand U5669 (N_5669,N_3302,N_2667);
and U5670 (N_5670,N_3953,N_2012);
or U5671 (N_5671,N_2364,N_3497);
and U5672 (N_5672,N_3684,N_2209);
nor U5673 (N_5673,N_3776,N_2773);
nand U5674 (N_5674,N_2720,N_2597);
and U5675 (N_5675,N_3679,N_2828);
xnor U5676 (N_5676,N_2056,N_3443);
nor U5677 (N_5677,N_2311,N_3222);
or U5678 (N_5678,N_3780,N_3767);
xnor U5679 (N_5679,N_2979,N_3519);
or U5680 (N_5680,N_3115,N_2398);
and U5681 (N_5681,N_3162,N_3265);
nor U5682 (N_5682,N_3962,N_2290);
nor U5683 (N_5683,N_2094,N_2194);
or U5684 (N_5684,N_2437,N_2490);
nand U5685 (N_5685,N_2715,N_2664);
or U5686 (N_5686,N_2193,N_2022);
and U5687 (N_5687,N_3173,N_2659);
nand U5688 (N_5688,N_2938,N_3019);
and U5689 (N_5689,N_2744,N_3464);
nor U5690 (N_5690,N_3355,N_2295);
or U5691 (N_5691,N_2916,N_3528);
and U5692 (N_5692,N_3664,N_3279);
xor U5693 (N_5693,N_3801,N_3754);
xnor U5694 (N_5694,N_2276,N_2940);
xor U5695 (N_5695,N_3796,N_3971);
nand U5696 (N_5696,N_3308,N_3067);
or U5697 (N_5697,N_3938,N_3810);
nand U5698 (N_5698,N_3126,N_3032);
nor U5699 (N_5699,N_2248,N_2357);
nand U5700 (N_5700,N_2590,N_3135);
and U5701 (N_5701,N_2868,N_3651);
xnor U5702 (N_5702,N_2215,N_3568);
or U5703 (N_5703,N_2400,N_2132);
nor U5704 (N_5704,N_2624,N_2349);
and U5705 (N_5705,N_3511,N_3752);
and U5706 (N_5706,N_3078,N_3583);
nand U5707 (N_5707,N_2631,N_2553);
nor U5708 (N_5708,N_3691,N_3469);
nand U5709 (N_5709,N_2182,N_2392);
and U5710 (N_5710,N_3514,N_2311);
xnor U5711 (N_5711,N_3703,N_2280);
nand U5712 (N_5712,N_3769,N_3243);
and U5713 (N_5713,N_3169,N_3951);
xor U5714 (N_5714,N_2114,N_2913);
xor U5715 (N_5715,N_2275,N_2711);
or U5716 (N_5716,N_2929,N_3405);
or U5717 (N_5717,N_3050,N_2653);
and U5718 (N_5718,N_3203,N_3106);
or U5719 (N_5719,N_3834,N_2145);
nor U5720 (N_5720,N_2379,N_2062);
or U5721 (N_5721,N_3678,N_3683);
nand U5722 (N_5722,N_3124,N_2366);
or U5723 (N_5723,N_3381,N_3493);
nor U5724 (N_5724,N_2160,N_3692);
and U5725 (N_5725,N_3557,N_2113);
xnor U5726 (N_5726,N_3223,N_2428);
and U5727 (N_5727,N_3329,N_3179);
or U5728 (N_5728,N_2244,N_2743);
or U5729 (N_5729,N_3218,N_3405);
nor U5730 (N_5730,N_2886,N_3972);
and U5731 (N_5731,N_3628,N_3164);
xnor U5732 (N_5732,N_3007,N_2006);
nand U5733 (N_5733,N_3091,N_3673);
nand U5734 (N_5734,N_2016,N_3140);
xnor U5735 (N_5735,N_2935,N_3897);
or U5736 (N_5736,N_3919,N_3206);
xor U5737 (N_5737,N_3787,N_2674);
xnor U5738 (N_5738,N_2146,N_2909);
nand U5739 (N_5739,N_3395,N_2567);
or U5740 (N_5740,N_2468,N_2498);
or U5741 (N_5741,N_3200,N_2352);
nor U5742 (N_5742,N_2525,N_2988);
or U5743 (N_5743,N_3768,N_3417);
nor U5744 (N_5744,N_2168,N_2260);
nand U5745 (N_5745,N_2397,N_3370);
or U5746 (N_5746,N_2556,N_3012);
nand U5747 (N_5747,N_3184,N_3360);
and U5748 (N_5748,N_3841,N_2152);
nor U5749 (N_5749,N_3020,N_2551);
xnor U5750 (N_5750,N_2888,N_2414);
or U5751 (N_5751,N_3998,N_2534);
nand U5752 (N_5752,N_3783,N_3337);
nor U5753 (N_5753,N_2627,N_2839);
or U5754 (N_5754,N_3821,N_3167);
nor U5755 (N_5755,N_2820,N_3457);
nand U5756 (N_5756,N_2089,N_3568);
xnor U5757 (N_5757,N_3265,N_2616);
or U5758 (N_5758,N_3752,N_2515);
nand U5759 (N_5759,N_2797,N_2650);
and U5760 (N_5760,N_2034,N_2922);
xnor U5761 (N_5761,N_2992,N_2810);
nor U5762 (N_5762,N_2790,N_3982);
nor U5763 (N_5763,N_3428,N_2760);
or U5764 (N_5764,N_3266,N_2105);
xnor U5765 (N_5765,N_3127,N_3788);
xnor U5766 (N_5766,N_2713,N_3247);
and U5767 (N_5767,N_2598,N_2194);
nor U5768 (N_5768,N_2767,N_2650);
nand U5769 (N_5769,N_2161,N_3636);
nor U5770 (N_5770,N_3975,N_3488);
or U5771 (N_5771,N_2844,N_2688);
and U5772 (N_5772,N_2292,N_3430);
and U5773 (N_5773,N_3856,N_3194);
or U5774 (N_5774,N_3909,N_2707);
nor U5775 (N_5775,N_3927,N_2919);
nor U5776 (N_5776,N_2344,N_2015);
nor U5777 (N_5777,N_2540,N_3979);
xor U5778 (N_5778,N_3920,N_2848);
or U5779 (N_5779,N_2184,N_2016);
nand U5780 (N_5780,N_3292,N_3964);
and U5781 (N_5781,N_3057,N_3770);
nand U5782 (N_5782,N_3211,N_3943);
and U5783 (N_5783,N_3011,N_2128);
or U5784 (N_5784,N_2614,N_2822);
or U5785 (N_5785,N_2932,N_2442);
and U5786 (N_5786,N_2851,N_3717);
xnor U5787 (N_5787,N_2385,N_3327);
and U5788 (N_5788,N_2501,N_3873);
nor U5789 (N_5789,N_2965,N_3052);
xnor U5790 (N_5790,N_2385,N_3269);
and U5791 (N_5791,N_2873,N_2155);
nor U5792 (N_5792,N_2718,N_2419);
nor U5793 (N_5793,N_3426,N_2422);
and U5794 (N_5794,N_2479,N_3456);
nand U5795 (N_5795,N_2291,N_2607);
nor U5796 (N_5796,N_2591,N_2068);
nand U5797 (N_5797,N_3436,N_2760);
and U5798 (N_5798,N_3680,N_2707);
or U5799 (N_5799,N_3157,N_3322);
and U5800 (N_5800,N_3426,N_3735);
and U5801 (N_5801,N_2685,N_3592);
and U5802 (N_5802,N_2960,N_2558);
nor U5803 (N_5803,N_2852,N_3679);
nand U5804 (N_5804,N_3506,N_2578);
and U5805 (N_5805,N_3222,N_2108);
nand U5806 (N_5806,N_3587,N_2771);
or U5807 (N_5807,N_2522,N_2392);
and U5808 (N_5808,N_3390,N_2968);
or U5809 (N_5809,N_2775,N_3163);
and U5810 (N_5810,N_2717,N_3489);
nor U5811 (N_5811,N_3904,N_2472);
or U5812 (N_5812,N_3564,N_2793);
nor U5813 (N_5813,N_3231,N_3520);
nand U5814 (N_5814,N_2611,N_3150);
nand U5815 (N_5815,N_3000,N_3992);
nor U5816 (N_5816,N_2746,N_3645);
or U5817 (N_5817,N_2967,N_3885);
or U5818 (N_5818,N_2071,N_3387);
or U5819 (N_5819,N_2404,N_2490);
nor U5820 (N_5820,N_2221,N_2965);
nand U5821 (N_5821,N_3914,N_3230);
nor U5822 (N_5822,N_2095,N_3146);
nor U5823 (N_5823,N_3587,N_3488);
or U5824 (N_5824,N_3053,N_2652);
and U5825 (N_5825,N_2036,N_3699);
xor U5826 (N_5826,N_3763,N_2949);
nand U5827 (N_5827,N_3011,N_3128);
nand U5828 (N_5828,N_3253,N_2661);
or U5829 (N_5829,N_3372,N_3579);
and U5830 (N_5830,N_2485,N_3362);
nor U5831 (N_5831,N_2058,N_3820);
or U5832 (N_5832,N_2019,N_2058);
xnor U5833 (N_5833,N_2142,N_3596);
and U5834 (N_5834,N_2239,N_2077);
nor U5835 (N_5835,N_3192,N_3264);
xor U5836 (N_5836,N_3499,N_3102);
and U5837 (N_5837,N_3452,N_3964);
or U5838 (N_5838,N_2497,N_2542);
xor U5839 (N_5839,N_3673,N_2891);
nand U5840 (N_5840,N_2874,N_2193);
xor U5841 (N_5841,N_3892,N_3993);
nor U5842 (N_5842,N_3504,N_2675);
nor U5843 (N_5843,N_3360,N_3629);
xor U5844 (N_5844,N_2358,N_2221);
xnor U5845 (N_5845,N_2893,N_3479);
and U5846 (N_5846,N_3118,N_3691);
and U5847 (N_5847,N_3145,N_3227);
and U5848 (N_5848,N_2038,N_2299);
nand U5849 (N_5849,N_2883,N_2033);
xnor U5850 (N_5850,N_3343,N_3577);
and U5851 (N_5851,N_2436,N_3740);
nand U5852 (N_5852,N_2366,N_3485);
or U5853 (N_5853,N_3026,N_3291);
or U5854 (N_5854,N_2238,N_3228);
nor U5855 (N_5855,N_3076,N_3389);
nand U5856 (N_5856,N_2297,N_3340);
xnor U5857 (N_5857,N_3522,N_3758);
nor U5858 (N_5858,N_3658,N_2692);
and U5859 (N_5859,N_2428,N_3081);
nor U5860 (N_5860,N_2698,N_2834);
nor U5861 (N_5861,N_3560,N_2900);
nor U5862 (N_5862,N_2612,N_3572);
nand U5863 (N_5863,N_2973,N_3965);
xor U5864 (N_5864,N_2752,N_2800);
nand U5865 (N_5865,N_2461,N_2579);
nand U5866 (N_5866,N_2979,N_3603);
nand U5867 (N_5867,N_2201,N_2220);
xor U5868 (N_5868,N_3527,N_2773);
and U5869 (N_5869,N_2082,N_2657);
nor U5870 (N_5870,N_2588,N_2643);
or U5871 (N_5871,N_3205,N_3603);
xnor U5872 (N_5872,N_2258,N_2396);
nand U5873 (N_5873,N_3749,N_2333);
nand U5874 (N_5874,N_3601,N_2087);
nand U5875 (N_5875,N_3590,N_3922);
or U5876 (N_5876,N_3739,N_2243);
or U5877 (N_5877,N_2114,N_2933);
and U5878 (N_5878,N_3750,N_2616);
xnor U5879 (N_5879,N_2685,N_3435);
xor U5880 (N_5880,N_2805,N_2132);
xor U5881 (N_5881,N_2520,N_2450);
and U5882 (N_5882,N_3052,N_2870);
nor U5883 (N_5883,N_3439,N_2062);
xor U5884 (N_5884,N_3184,N_2017);
and U5885 (N_5885,N_2130,N_2010);
or U5886 (N_5886,N_2332,N_3241);
or U5887 (N_5887,N_3862,N_3729);
xor U5888 (N_5888,N_2992,N_2979);
nor U5889 (N_5889,N_3063,N_2189);
nand U5890 (N_5890,N_2702,N_3133);
and U5891 (N_5891,N_3019,N_2519);
and U5892 (N_5892,N_3535,N_2460);
xor U5893 (N_5893,N_3812,N_2827);
and U5894 (N_5894,N_3742,N_3162);
and U5895 (N_5895,N_2669,N_2492);
xnor U5896 (N_5896,N_2150,N_2968);
nor U5897 (N_5897,N_2272,N_2286);
or U5898 (N_5898,N_3794,N_2407);
xnor U5899 (N_5899,N_2346,N_3022);
and U5900 (N_5900,N_3152,N_2688);
xnor U5901 (N_5901,N_3224,N_2363);
nor U5902 (N_5902,N_3310,N_2900);
and U5903 (N_5903,N_3024,N_3552);
nand U5904 (N_5904,N_3207,N_2085);
or U5905 (N_5905,N_3809,N_2531);
nor U5906 (N_5906,N_3140,N_3138);
or U5907 (N_5907,N_3670,N_3525);
xnor U5908 (N_5908,N_2395,N_2310);
and U5909 (N_5909,N_2888,N_3914);
xnor U5910 (N_5910,N_3757,N_3277);
xnor U5911 (N_5911,N_2840,N_3264);
xor U5912 (N_5912,N_3150,N_3828);
and U5913 (N_5913,N_2026,N_3642);
and U5914 (N_5914,N_3957,N_3282);
nor U5915 (N_5915,N_3518,N_3962);
and U5916 (N_5916,N_3375,N_3796);
xnor U5917 (N_5917,N_3888,N_3833);
xnor U5918 (N_5918,N_3995,N_3093);
xnor U5919 (N_5919,N_3416,N_3145);
nand U5920 (N_5920,N_3760,N_3091);
and U5921 (N_5921,N_2022,N_2199);
and U5922 (N_5922,N_2054,N_3057);
or U5923 (N_5923,N_3228,N_3364);
or U5924 (N_5924,N_2851,N_2019);
and U5925 (N_5925,N_2567,N_3270);
nand U5926 (N_5926,N_3916,N_3804);
xor U5927 (N_5927,N_3452,N_3107);
nor U5928 (N_5928,N_3302,N_2026);
or U5929 (N_5929,N_3596,N_3851);
or U5930 (N_5930,N_3708,N_3136);
and U5931 (N_5931,N_3098,N_3588);
xnor U5932 (N_5932,N_3151,N_2217);
or U5933 (N_5933,N_3505,N_2305);
xor U5934 (N_5934,N_2197,N_3830);
xnor U5935 (N_5935,N_2183,N_3118);
nor U5936 (N_5936,N_3028,N_2461);
and U5937 (N_5937,N_3021,N_3671);
xor U5938 (N_5938,N_3483,N_3825);
nor U5939 (N_5939,N_2141,N_3230);
nor U5940 (N_5940,N_3560,N_3624);
xor U5941 (N_5941,N_3561,N_3212);
or U5942 (N_5942,N_3080,N_2002);
and U5943 (N_5943,N_2780,N_3681);
nor U5944 (N_5944,N_3566,N_3986);
and U5945 (N_5945,N_2542,N_3189);
nor U5946 (N_5946,N_2168,N_3873);
nand U5947 (N_5947,N_2437,N_3119);
and U5948 (N_5948,N_3375,N_2721);
or U5949 (N_5949,N_2241,N_2702);
xnor U5950 (N_5950,N_3629,N_2996);
nand U5951 (N_5951,N_3093,N_3814);
or U5952 (N_5952,N_2868,N_2697);
nor U5953 (N_5953,N_3923,N_3580);
or U5954 (N_5954,N_2865,N_2877);
nand U5955 (N_5955,N_3324,N_2370);
nor U5956 (N_5956,N_3104,N_3013);
nor U5957 (N_5957,N_2432,N_2634);
xnor U5958 (N_5958,N_2294,N_2938);
nor U5959 (N_5959,N_2027,N_2801);
nor U5960 (N_5960,N_3575,N_3366);
nand U5961 (N_5961,N_3854,N_2192);
nor U5962 (N_5962,N_3135,N_2660);
or U5963 (N_5963,N_3722,N_3878);
and U5964 (N_5964,N_2353,N_3800);
xnor U5965 (N_5965,N_3342,N_3285);
nand U5966 (N_5966,N_2064,N_2401);
nor U5967 (N_5967,N_3834,N_3770);
nor U5968 (N_5968,N_2144,N_3097);
nand U5969 (N_5969,N_3289,N_2309);
nand U5970 (N_5970,N_2336,N_3729);
xor U5971 (N_5971,N_3112,N_2210);
nor U5972 (N_5972,N_3251,N_3804);
or U5973 (N_5973,N_2094,N_3247);
nand U5974 (N_5974,N_2556,N_3822);
or U5975 (N_5975,N_2517,N_3258);
nand U5976 (N_5976,N_2035,N_3034);
xor U5977 (N_5977,N_3427,N_3621);
or U5978 (N_5978,N_2803,N_2757);
nand U5979 (N_5979,N_2721,N_3793);
nor U5980 (N_5980,N_2216,N_2082);
and U5981 (N_5981,N_2925,N_2131);
and U5982 (N_5982,N_3666,N_3486);
nand U5983 (N_5983,N_2704,N_2779);
xnor U5984 (N_5984,N_2695,N_2656);
xnor U5985 (N_5985,N_2344,N_2932);
nor U5986 (N_5986,N_3464,N_2735);
and U5987 (N_5987,N_3597,N_2679);
and U5988 (N_5988,N_2905,N_3515);
and U5989 (N_5989,N_2039,N_3729);
or U5990 (N_5990,N_3139,N_2272);
nand U5991 (N_5991,N_3468,N_2319);
and U5992 (N_5992,N_3097,N_2305);
nor U5993 (N_5993,N_2152,N_3911);
nand U5994 (N_5994,N_3459,N_3323);
nor U5995 (N_5995,N_2938,N_2796);
nand U5996 (N_5996,N_3154,N_3766);
xnor U5997 (N_5997,N_2176,N_3799);
nand U5998 (N_5998,N_2302,N_2772);
nor U5999 (N_5999,N_2550,N_3920);
nand U6000 (N_6000,N_5539,N_4777);
nor U6001 (N_6001,N_5808,N_4087);
xor U6002 (N_6002,N_4694,N_5378);
nand U6003 (N_6003,N_4944,N_5165);
nor U6004 (N_6004,N_5101,N_5752);
or U6005 (N_6005,N_4269,N_4957);
nor U6006 (N_6006,N_4824,N_5576);
xor U6007 (N_6007,N_4823,N_5900);
or U6008 (N_6008,N_4207,N_5942);
nor U6009 (N_6009,N_5409,N_4245);
nand U6010 (N_6010,N_4666,N_4853);
nand U6011 (N_6011,N_5063,N_5919);
xor U6012 (N_6012,N_5184,N_5369);
xor U6013 (N_6013,N_4599,N_5018);
nand U6014 (N_6014,N_5178,N_5312);
and U6015 (N_6015,N_4125,N_5334);
nor U6016 (N_6016,N_5427,N_5742);
xor U6017 (N_6017,N_5273,N_5897);
and U6018 (N_6018,N_4936,N_5297);
and U6019 (N_6019,N_4438,N_4050);
or U6020 (N_6020,N_5182,N_4955);
or U6021 (N_6021,N_5666,N_5110);
xnor U6022 (N_6022,N_4831,N_4295);
and U6023 (N_6023,N_4258,N_4371);
nand U6024 (N_6024,N_5092,N_4165);
xor U6025 (N_6025,N_4890,N_4031);
nor U6026 (N_6026,N_4619,N_4387);
xnor U6027 (N_6027,N_5392,N_5499);
nor U6028 (N_6028,N_4586,N_5336);
nand U6029 (N_6029,N_5558,N_5848);
and U6030 (N_6030,N_4945,N_4391);
xor U6031 (N_6031,N_4151,N_4718);
xnor U6032 (N_6032,N_4605,N_4393);
nor U6033 (N_6033,N_5533,N_5448);
and U6034 (N_6034,N_4849,N_4174);
nor U6035 (N_6035,N_5434,N_5335);
and U6036 (N_6036,N_5798,N_4389);
or U6037 (N_6037,N_4642,N_4836);
and U6038 (N_6038,N_5710,N_5955);
or U6039 (N_6039,N_5037,N_5021);
and U6040 (N_6040,N_4896,N_4287);
or U6041 (N_6041,N_5795,N_5344);
nor U6042 (N_6042,N_5598,N_5714);
or U6043 (N_6043,N_5245,N_4638);
and U6044 (N_6044,N_4872,N_4439);
or U6045 (N_6045,N_5729,N_4120);
nor U6046 (N_6046,N_5768,N_5121);
and U6047 (N_6047,N_5503,N_5132);
nand U6048 (N_6048,N_4555,N_4613);
nand U6049 (N_6049,N_5609,N_5460);
or U6050 (N_6050,N_4964,N_5876);
nand U6051 (N_6051,N_5888,N_5472);
xor U6052 (N_6052,N_4437,N_4693);
and U6053 (N_6053,N_5176,N_4710);
nor U6054 (N_6054,N_4539,N_4339);
or U6055 (N_6055,N_5356,N_5571);
nor U6056 (N_6056,N_4152,N_5200);
xnor U6057 (N_6057,N_4624,N_5089);
or U6058 (N_6058,N_4700,N_5163);
or U6059 (N_6059,N_5424,N_4812);
and U6060 (N_6060,N_4435,N_5801);
nand U6061 (N_6061,N_4311,N_4792);
or U6062 (N_6062,N_4829,N_5115);
nor U6063 (N_6063,N_5407,N_5148);
xor U6064 (N_6064,N_5947,N_5974);
xnor U6065 (N_6065,N_5720,N_4526);
or U6066 (N_6066,N_5331,N_5152);
nand U6067 (N_6067,N_4141,N_4067);
and U6068 (N_6068,N_4013,N_5168);
nand U6069 (N_6069,N_5998,N_5903);
nand U6070 (N_6070,N_4430,N_4161);
and U6071 (N_6071,N_4279,N_5096);
xnor U6072 (N_6072,N_4464,N_4550);
or U6073 (N_6073,N_5253,N_5939);
and U6074 (N_6074,N_4720,N_4815);
xnor U6075 (N_6075,N_4881,N_4545);
nand U6076 (N_6076,N_5582,N_5570);
or U6077 (N_6077,N_5451,N_4509);
nor U6078 (N_6078,N_4768,N_5177);
and U6079 (N_6079,N_5195,N_5034);
or U6080 (N_6080,N_4932,N_4787);
xnor U6081 (N_6081,N_4755,N_5299);
and U6082 (N_6082,N_4959,N_5347);
and U6083 (N_6083,N_5726,N_5305);
and U6084 (N_6084,N_4711,N_4782);
nor U6085 (N_6085,N_5102,N_4901);
nand U6086 (N_6086,N_4482,N_4257);
xor U6087 (N_6087,N_4969,N_4521);
or U6088 (N_6088,N_4578,N_4754);
and U6089 (N_6089,N_5327,N_4562);
nand U6090 (N_6090,N_4956,N_4119);
and U6091 (N_6091,N_5716,N_5862);
nand U6092 (N_6092,N_5358,N_4556);
xnor U6093 (N_6093,N_4088,N_4805);
nand U6094 (N_6094,N_5512,N_4401);
and U6095 (N_6095,N_4200,N_5519);
or U6096 (N_6096,N_4885,N_4770);
or U6097 (N_6097,N_4380,N_4227);
or U6098 (N_6098,N_5401,N_5890);
or U6099 (N_6099,N_5703,N_5529);
nand U6100 (N_6100,N_4024,N_5678);
and U6101 (N_6101,N_5161,N_4834);
xnor U6102 (N_6102,N_5119,N_4445);
and U6103 (N_6103,N_4403,N_5643);
and U6104 (N_6104,N_5107,N_4073);
xnor U6105 (N_6105,N_4297,N_5559);
xor U6106 (N_6106,N_5639,N_4789);
nor U6107 (N_6107,N_4867,N_4377);
nor U6108 (N_6108,N_4116,N_4835);
xor U6109 (N_6109,N_5692,N_4669);
nor U6110 (N_6110,N_5926,N_4347);
nand U6111 (N_6111,N_4988,N_5035);
nand U6112 (N_6112,N_5129,N_5659);
nand U6113 (N_6113,N_5541,N_5540);
xnor U6114 (N_6114,N_5206,N_4358);
and U6115 (N_6115,N_5717,N_4048);
and U6116 (N_6116,N_5288,N_4123);
and U6117 (N_6117,N_5563,N_4267);
nor U6118 (N_6118,N_5008,N_4385);
xnor U6119 (N_6119,N_4290,N_4360);
nand U6120 (N_6120,N_5332,N_5295);
or U6121 (N_6121,N_5945,N_4589);
nand U6122 (N_6122,N_4863,N_5581);
xor U6123 (N_6123,N_5186,N_4035);
and U6124 (N_6124,N_4884,N_5954);
nor U6125 (N_6125,N_4156,N_4410);
nand U6126 (N_6126,N_4384,N_4177);
nor U6127 (N_6127,N_4967,N_4612);
and U6128 (N_6128,N_5470,N_5383);
or U6129 (N_6129,N_4514,N_5938);
xor U6130 (N_6130,N_4176,N_4242);
nand U6131 (N_6131,N_5621,N_5611);
xor U6132 (N_6132,N_5773,N_5341);
or U6133 (N_6133,N_4256,N_5817);
nor U6134 (N_6134,N_5836,N_4193);
or U6135 (N_6135,N_5811,N_4054);
and U6136 (N_6136,N_4595,N_4785);
and U6137 (N_6137,N_5619,N_4293);
xnor U6138 (N_6138,N_4981,N_5647);
and U6139 (N_6139,N_5125,N_5651);
and U6140 (N_6140,N_4454,N_4844);
or U6141 (N_6141,N_5397,N_4052);
and U6142 (N_6142,N_4366,N_4852);
and U6143 (N_6143,N_4738,N_5158);
nand U6144 (N_6144,N_5661,N_5964);
nand U6145 (N_6145,N_4921,N_5108);
and U6146 (N_6146,N_4549,N_4222);
nor U6147 (N_6147,N_4497,N_4034);
nand U6148 (N_6148,N_5595,N_4906);
and U6149 (N_6149,N_5761,N_5737);
nor U6150 (N_6150,N_5544,N_5914);
nand U6151 (N_6151,N_5930,N_4596);
xor U6152 (N_6152,N_4064,N_4517);
nand U6153 (N_6153,N_5793,N_4576);
or U6154 (N_6154,N_5188,N_5046);
and U6155 (N_6155,N_4786,N_4171);
and U6156 (N_6156,N_4271,N_5654);
xnor U6157 (N_6157,N_5216,N_5875);
xnor U6158 (N_6158,N_4124,N_5260);
and U6159 (N_6159,N_5244,N_5412);
or U6160 (N_6160,N_5650,N_5302);
nor U6161 (N_6161,N_5083,N_4224);
nand U6162 (N_6162,N_4900,N_5461);
or U6163 (N_6163,N_4658,N_4769);
or U6164 (N_6164,N_5003,N_5185);
xor U6165 (N_6165,N_4218,N_5638);
nand U6166 (N_6166,N_4799,N_4922);
nor U6167 (N_6167,N_5859,N_5174);
and U6168 (N_6168,N_5498,N_5975);
nand U6169 (N_6169,N_5916,N_4062);
or U6170 (N_6170,N_4065,N_5738);
or U6171 (N_6171,N_5749,N_5991);
xnor U6172 (N_6172,N_4089,N_5880);
xnor U6173 (N_6173,N_4428,N_4028);
xnor U6174 (N_6174,N_4995,N_4551);
and U6175 (N_6175,N_4818,N_4895);
xnor U6176 (N_6176,N_4351,N_4663);
nor U6177 (N_6177,N_5951,N_4682);
nand U6178 (N_6178,N_5311,N_4928);
nand U6179 (N_6179,N_4966,N_4811);
or U6180 (N_6180,N_4870,N_4312);
and U6181 (N_6181,N_5522,N_5950);
xor U6182 (N_6182,N_4727,N_4847);
and U6183 (N_6183,N_4983,N_5677);
xor U6184 (N_6184,N_5193,N_5632);
or U6185 (N_6185,N_4903,N_5791);
xnor U6186 (N_6186,N_5814,N_4471);
nand U6187 (N_6187,N_5599,N_4668);
nor U6188 (N_6188,N_5387,N_5100);
or U6189 (N_6189,N_4997,N_5746);
nor U6190 (N_6190,N_5391,N_4732);
and U6191 (N_6191,N_4661,N_4505);
or U6192 (N_6192,N_4146,N_5725);
xor U6193 (N_6193,N_4577,N_4973);
nor U6194 (N_6194,N_4272,N_5170);
or U6195 (N_6195,N_4275,N_5553);
or U6196 (N_6196,N_4701,N_5143);
or U6197 (N_6197,N_5385,N_5411);
nor U6198 (N_6198,N_4976,N_4513);
or U6199 (N_6199,N_4080,N_5285);
nand U6200 (N_6200,N_5354,N_4652);
nand U6201 (N_6201,N_5094,N_5220);
or U6202 (N_6202,N_5247,N_5361);
or U6203 (N_6203,N_5010,N_5007);
and U6204 (N_6204,N_4862,N_4296);
nor U6205 (N_6205,N_4571,N_4677);
or U6206 (N_6206,N_4457,N_5999);
nand U6207 (N_6207,N_5464,N_5410);
nor U6208 (N_6208,N_4373,N_5296);
nand U6209 (N_6209,N_5779,N_4761);
nor U6210 (N_6210,N_5405,N_4283);
or U6211 (N_6211,N_5022,N_5204);
and U6212 (N_6212,N_5906,N_4570);
or U6213 (N_6213,N_5868,N_4098);
nor U6214 (N_6214,N_4343,N_5976);
and U6215 (N_6215,N_4179,N_5166);
or U6216 (N_6216,N_4208,N_4408);
nor U6217 (N_6217,N_5180,N_4203);
nand U6218 (N_6218,N_4778,N_5386);
nand U6219 (N_6219,N_5538,N_5851);
xnor U6220 (N_6220,N_4491,N_4075);
or U6221 (N_6221,N_5524,N_5287);
nand U6222 (N_6222,N_4802,N_4210);
and U6223 (N_6223,N_4164,N_5755);
nor U6224 (N_6224,N_5794,N_5648);
nor U6225 (N_6225,N_5600,N_5040);
nand U6226 (N_6226,N_5835,N_4680);
nor U6227 (N_6227,N_5702,N_5751);
nand U6228 (N_6228,N_4078,N_5493);
nand U6229 (N_6229,N_5685,N_5882);
or U6230 (N_6230,N_5421,N_5282);
or U6231 (N_6231,N_4306,N_4608);
and U6232 (N_6232,N_5612,N_5658);
nand U6233 (N_6233,N_4560,N_5854);
or U6234 (N_6234,N_4051,N_5915);
or U6235 (N_6235,N_5970,N_5471);
or U6236 (N_6236,N_5437,N_4460);
and U6237 (N_6237,N_4473,N_4458);
and U6238 (N_6238,N_5363,N_4247);
and U6239 (N_6239,N_4322,N_5633);
or U6240 (N_6240,N_5248,N_5899);
nand U6241 (N_6241,N_4592,N_5987);
nor U6242 (N_6242,N_4425,N_5274);
or U6243 (N_6243,N_4929,N_5966);
or U6244 (N_6244,N_4868,N_5775);
xnor U6245 (N_6245,N_4121,N_5218);
nand U6246 (N_6246,N_5227,N_5453);
and U6247 (N_6247,N_4991,N_5649);
nand U6248 (N_6248,N_4828,N_4593);
nand U6249 (N_6249,N_5045,N_5479);
xor U6250 (N_6250,N_4664,N_4135);
xnor U6251 (N_6251,N_4305,N_5554);
and U6252 (N_6252,N_5229,N_4108);
and U6253 (N_6253,N_5514,N_5318);
nor U6254 (N_6254,N_5754,N_4859);
nand U6255 (N_6255,N_4766,N_4633);
or U6256 (N_6256,N_4243,N_5160);
xnor U6257 (N_6257,N_4039,N_5236);
nor U6258 (N_6258,N_4490,N_4582);
xnor U6259 (N_6259,N_5001,N_5797);
nand U6260 (N_6260,N_5694,N_5940);
and U6261 (N_6261,N_5199,N_5281);
or U6262 (N_6262,N_5672,N_4202);
nor U6263 (N_6263,N_4648,N_4688);
xnor U6264 (N_6264,N_4538,N_5815);
nand U6265 (N_6265,N_4790,N_5074);
nand U6266 (N_6266,N_4702,N_5187);
xor U6267 (N_6267,N_5044,N_5958);
nand U6268 (N_6268,N_4486,N_4166);
xnor U6269 (N_6269,N_4014,N_4563);
nand U6270 (N_6270,N_5719,N_5556);
xor U6271 (N_6271,N_5225,N_5442);
nand U6272 (N_6272,N_5727,N_5925);
or U6273 (N_6273,N_5164,N_5144);
xor U6274 (N_6274,N_5137,N_4318);
nand U6275 (N_6275,N_4059,N_5333);
xnor U6276 (N_6276,N_5821,N_5809);
xor U6277 (N_6277,N_5126,N_4912);
nor U6278 (N_6278,N_5262,N_5413);
and U6279 (N_6279,N_4255,N_5239);
or U6280 (N_6280,N_5252,N_4703);
nand U6281 (N_6281,N_4470,N_5111);
nor U6282 (N_6282,N_5896,N_5603);
or U6283 (N_6283,N_5766,N_4573);
or U6284 (N_6284,N_5587,N_4617);
nor U6285 (N_6285,N_5436,N_4234);
nor U6286 (N_6286,N_4451,N_5861);
and U6287 (N_6287,N_4249,N_4449);
nand U6288 (N_6288,N_5476,N_5231);
xor U6289 (N_6289,N_5760,N_4984);
and U6290 (N_6290,N_4813,N_5824);
or U6291 (N_6291,N_5475,N_4525);
nand U6292 (N_6292,N_4914,N_5934);
xnor U6293 (N_6293,N_5446,N_5605);
nand U6294 (N_6294,N_5626,N_5078);
xnor U6295 (N_6295,N_5447,N_4420);
nand U6296 (N_6296,N_5028,N_4583);
nand U6297 (N_6297,N_5723,N_5969);
or U6298 (N_6298,N_4467,N_4848);
and U6299 (N_6299,N_4076,N_4554);
nand U6300 (N_6300,N_4447,N_4341);
or U6301 (N_6301,N_4620,N_4531);
nor U6302 (N_6302,N_5860,N_5822);
nand U6303 (N_6303,N_4797,N_4114);
nor U6304 (N_6304,N_5933,N_4641);
nor U6305 (N_6305,N_4559,N_5850);
xor U6306 (N_6306,N_4697,N_4337);
nor U6307 (N_6307,N_5292,N_5316);
nor U6308 (N_6308,N_4947,N_4806);
and U6309 (N_6309,N_4016,N_5776);
xnor U6310 (N_6310,N_5031,N_4219);
nor U6311 (N_6311,N_5732,N_4396);
nand U6312 (N_6312,N_5763,N_4000);
or U6313 (N_6313,N_5557,N_4071);
nand U6314 (N_6314,N_4026,N_5445);
nor U6315 (N_6315,N_4047,N_5384);
xor U6316 (N_6316,N_4845,N_5173);
or U6317 (N_6317,N_5994,N_5560);
or U6318 (N_6318,N_5482,N_4647);
xor U6319 (N_6319,N_4581,N_4044);
or U6320 (N_6320,N_5415,N_5601);
xnor U6321 (N_6321,N_5128,N_4502);
and U6322 (N_6322,N_4692,N_4736);
xor U6323 (N_6323,N_5712,N_5147);
xor U6324 (N_6324,N_5833,N_5474);
xor U6325 (N_6325,N_4137,N_5511);
nand U6326 (N_6326,N_5543,N_5771);
or U6327 (N_6327,N_5085,N_5660);
xnor U6328 (N_6328,N_5490,N_5076);
or U6329 (N_6329,N_5614,N_4771);
and U6330 (N_6330,N_5064,N_5124);
nand U6331 (N_6331,N_4147,N_4791);
xnor U6332 (N_6332,N_4740,N_4518);
xnor U6333 (N_6333,N_5623,N_5346);
nand U6334 (N_6334,N_4394,N_5531);
nand U6335 (N_6335,N_5033,N_5462);
and U6336 (N_6336,N_5172,N_4418);
nand U6337 (N_6337,N_4023,N_4625);
nor U6338 (N_6338,N_5566,N_5644);
or U6339 (N_6339,N_5910,N_4270);
and U6340 (N_6340,N_5904,N_4367);
or U6341 (N_6341,N_5912,N_4540);
or U6342 (N_6342,N_5443,N_5151);
and U6343 (N_6343,N_4169,N_4734);
and U6344 (N_6344,N_5131,N_5374);
nor U6345 (N_6345,N_4160,N_4898);
nor U6346 (N_6346,N_5155,N_4499);
nand U6347 (N_6347,N_5050,N_4977);
and U6348 (N_6348,N_5799,N_4996);
and U6349 (N_6349,N_5535,N_4332);
and U6350 (N_6350,N_5527,N_5264);
nand U6351 (N_6351,N_5205,N_4604);
nor U6352 (N_6352,N_5487,N_4474);
xor U6353 (N_6353,N_5834,N_4130);
nand U6354 (N_6354,N_4992,N_4522);
nor U6355 (N_6355,N_5960,N_5812);
xor U6356 (N_6356,N_5329,N_4468);
xor U6357 (N_6357,N_5425,N_4724);
xor U6358 (N_6358,N_5463,N_5241);
and U6359 (N_6359,N_4235,N_5234);
nand U6360 (N_6360,N_5982,N_4299);
or U6361 (N_6361,N_4580,N_4049);
nor U6362 (N_6362,N_4622,N_4086);
or U6363 (N_6363,N_4291,N_4484);
nand U6364 (N_6364,N_4767,N_5408);
or U6365 (N_6365,N_5961,N_5189);
xor U6366 (N_6366,N_4905,N_5709);
or U6367 (N_6367,N_4175,N_5081);
or U6368 (N_6368,N_5291,N_4342);
or U6369 (N_6369,N_4060,N_4877);
and U6370 (N_6370,N_5841,N_4747);
and U6371 (N_6371,N_4731,N_5140);
or U6372 (N_6372,N_5098,N_4310);
or U6373 (N_6373,N_4561,N_4386);
and U6374 (N_6374,N_5782,N_5303);
or U6375 (N_6375,N_5466,N_4572);
and U6376 (N_6376,N_4241,N_5853);
nand U6377 (N_6377,N_5546,N_5803);
and U6378 (N_6378,N_5497,N_4574);
nor U6379 (N_6379,N_4676,N_5084);
or U6380 (N_6380,N_4359,N_5774);
or U6381 (N_6381,N_4276,N_4558);
xor U6382 (N_6382,N_4354,N_4597);
and U6383 (N_6383,N_5058,N_5240);
nand U6384 (N_6384,N_5207,N_4833);
nor U6385 (N_6385,N_4433,N_4012);
nor U6386 (N_6386,N_5665,N_4307);
nand U6387 (N_6387,N_5502,N_5596);
and U6388 (N_6388,N_5597,N_5887);
nor U6389 (N_6389,N_4917,N_5713);
or U6390 (N_6390,N_4808,N_4240);
nand U6391 (N_6391,N_5990,N_4409);
nand U6392 (N_6392,N_4092,N_5894);
or U6393 (N_6393,N_5985,N_4372);
xnor U6394 (N_6394,N_4838,N_4935);
nand U6395 (N_6395,N_4729,N_4244);
or U6396 (N_6396,N_5388,N_5201);
nor U6397 (N_6397,N_4285,N_5069);
nand U6398 (N_6398,N_5259,N_4102);
or U6399 (N_6399,N_4238,N_5704);
and U6400 (N_6400,N_5406,N_4205);
and U6401 (N_6401,N_4330,N_5375);
and U6402 (N_6402,N_4980,N_5872);
nand U6403 (N_6403,N_5550,N_5562);
nand U6404 (N_6404,N_4500,N_5509);
and U6405 (N_6405,N_4636,N_4780);
and U6406 (N_6406,N_4609,N_5454);
nor U6407 (N_6407,N_5818,N_4519);
nand U6408 (N_6408,N_4998,N_5222);
xnor U6409 (N_6409,N_4392,N_4897);
xnor U6410 (N_6410,N_5534,N_4252);
and U6411 (N_6411,N_4429,N_4335);
or U6412 (N_6412,N_5065,N_4716);
xor U6413 (N_6413,N_4534,N_4541);
xnor U6414 (N_6414,N_5283,N_5099);
nand U6415 (N_6415,N_5864,N_5831);
nor U6416 (N_6416,N_5747,N_5845);
nor U6417 (N_6417,N_5636,N_5551);
xor U6418 (N_6418,N_5625,N_5324);
xnor U6419 (N_6419,N_4376,N_4284);
nand U6420 (N_6420,N_5526,N_5922);
nand U6421 (N_6421,N_5153,N_4374);
and U6422 (N_6422,N_5898,N_5515);
or U6423 (N_6423,N_5181,N_5414);
nand U6424 (N_6424,N_4423,N_4159);
nor U6425 (N_6425,N_5000,N_4348);
nor U6426 (N_6426,N_4397,N_4002);
nor U6427 (N_6427,N_4704,N_4653);
nand U6428 (N_6428,N_4631,N_4678);
nand U6429 (N_6429,N_4629,N_5030);
nand U6430 (N_6430,N_4431,N_5149);
xnor U6431 (N_6431,N_4046,N_5592);
nand U6432 (N_6432,N_4079,N_5986);
or U6433 (N_6433,N_4960,N_5983);
or U6434 (N_6434,N_5968,N_5457);
xnor U6435 (N_6435,N_4209,N_5146);
or U6436 (N_6436,N_4855,N_4657);
nand U6437 (N_6437,N_4153,N_4814);
and U6438 (N_6438,N_5017,N_4887);
and U6439 (N_6439,N_4524,N_4093);
and U6440 (N_6440,N_4744,N_4839);
and U6441 (N_6441,N_4452,N_5150);
nor U6442 (N_6442,N_4266,N_4850);
xor U6443 (N_6443,N_4939,N_5846);
nand U6444 (N_6444,N_4830,N_4781);
and U6445 (N_6445,N_4616,N_5591);
nand U6446 (N_6446,N_4118,N_4331);
xor U6447 (N_6447,N_5212,N_5908);
nand U6448 (N_6448,N_5362,N_4606);
xnor U6449 (N_6449,N_4810,N_4999);
nor U6450 (N_6450,N_4197,N_5674);
or U6451 (N_6451,N_4715,N_4533);
nor U6452 (N_6452,N_4494,N_5029);
nand U6453 (N_6453,N_4399,N_5469);
and U6454 (N_6454,N_5988,N_4691);
and U6455 (N_6455,N_4378,N_5893);
nand U6456 (N_6456,N_5006,N_5567);
nor U6457 (N_6457,N_4507,N_4301);
xnor U6458 (N_6458,N_5748,N_4195);
and U6459 (N_6459,N_4492,N_4298);
or U6460 (N_6460,N_5060,N_5767);
and U6461 (N_6461,N_4091,N_4404);
and U6462 (N_6462,N_5807,N_5655);
nor U6463 (N_6463,N_4909,N_4741);
and U6464 (N_6464,N_4199,N_4520);
xnor U6465 (N_6465,N_5077,N_4753);
xnor U6466 (N_6466,N_5870,N_4925);
or U6467 (N_6467,N_4112,N_5931);
xnor U6468 (N_6468,N_4547,N_5744);
nor U6469 (N_6469,N_4598,N_4294);
or U6470 (N_6470,N_5032,N_5989);
xnor U6471 (N_6471,N_4730,N_4673);
nor U6472 (N_6472,N_5048,N_4557);
nor U6473 (N_6473,N_4488,N_5491);
xnor U6474 (N_6474,N_5604,N_5428);
and U6475 (N_6475,N_5321,N_5480);
nor U6476 (N_6476,N_4379,N_5456);
and U6477 (N_6477,N_5284,N_5404);
and U6478 (N_6478,N_5417,N_5352);
nand U6479 (N_6479,N_5242,N_4751);
or U6480 (N_6480,N_4798,N_5431);
nor U6481 (N_6481,N_5120,N_4292);
and U6482 (N_6482,N_5444,N_5772);
or U6483 (N_6483,N_5663,N_4178);
or U6484 (N_6484,N_4854,N_4874);
nor U6485 (N_6485,N_4304,N_4614);
and U6486 (N_6486,N_5485,N_4889);
and U6487 (N_6487,N_4695,N_5440);
nor U6488 (N_6488,N_5235,N_5909);
or U6489 (N_6489,N_4004,N_5832);
xor U6490 (N_6490,N_4809,N_5459);
xnor U6491 (N_6491,N_5267,N_4325);
and U6492 (N_6492,N_4183,N_5123);
xor U6493 (N_6493,N_5090,N_4816);
or U6494 (N_6494,N_5328,N_4032);
xor U6495 (N_6495,N_5043,N_4878);
nand U6496 (N_6496,N_5097,N_4113);
or U6497 (N_6497,N_5923,N_4154);
nor U6498 (N_6498,N_5802,N_4434);
or U6499 (N_6499,N_5932,N_5630);
and U6500 (N_6500,N_4419,N_5373);
nor U6501 (N_6501,N_5902,N_4068);
xnor U6502 (N_6502,N_4214,N_4543);
xor U6503 (N_6503,N_4587,N_5095);
nor U6504 (N_6504,N_5657,N_5686);
and U6505 (N_6505,N_5676,N_5357);
xnor U6506 (N_6506,N_5399,N_4248);
and U6507 (N_6507,N_4565,N_4876);
nand U6508 (N_6508,N_5504,N_5217);
or U6509 (N_6509,N_5827,N_4223);
xnor U6510 (N_6510,N_5135,N_4020);
and U6511 (N_6511,N_4277,N_5279);
and U6512 (N_6512,N_4970,N_4066);
nand U6513 (N_6513,N_5465,N_4355);
or U6514 (N_6514,N_5696,N_5602);
xnor U6515 (N_6515,N_4455,N_4516);
nand U6516 (N_6516,N_5731,N_4313);
nor U6517 (N_6517,N_4097,N_5300);
nor U6518 (N_6518,N_5588,N_4552);
nor U6519 (N_6519,N_5027,N_4145);
nand U6520 (N_6520,N_5277,N_4607);
or U6521 (N_6521,N_4400,N_4229);
and U6522 (N_6522,N_5145,N_5169);
nor U6523 (N_6523,N_5885,N_5025);
or U6524 (N_6524,N_4254,N_4228);
and U6525 (N_6525,N_4634,N_5268);
or U6526 (N_6526,N_5769,N_5730);
or U6527 (N_6527,N_5805,N_4784);
nor U6528 (N_6528,N_4601,N_5707);
xnor U6529 (N_6529,N_5082,N_4941);
and U6530 (N_6530,N_4940,N_5418);
nand U6531 (N_6531,N_4149,N_4542);
and U6532 (N_6532,N_4264,N_5056);
xor U6533 (N_6533,N_5739,N_4143);
xnor U6534 (N_6534,N_4323,N_5977);
nor U6535 (N_6535,N_5722,N_5946);
nor U6536 (N_6536,N_5856,N_5957);
and U6537 (N_6537,N_4649,N_4709);
nor U6538 (N_6538,N_5495,N_4671);
xor U6539 (N_6539,N_4170,N_4546);
nand U6540 (N_6540,N_4989,N_5314);
nand U6541 (N_6541,N_5345,N_4111);
or U6542 (N_6542,N_5080,N_4259);
nor U6543 (N_6543,N_4459,N_4172);
xnor U6544 (N_6544,N_5432,N_5866);
nor U6545 (N_6545,N_5340,N_5765);
and U6546 (N_6546,N_4487,N_4674);
nand U6547 (N_6547,N_5039,N_5757);
xor U6548 (N_6548,N_5372,N_4101);
xor U6549 (N_6549,N_4320,N_5104);
nand U6550 (N_6550,N_5380,N_4196);
or U6551 (N_6551,N_4057,N_4742);
xnor U6552 (N_6552,N_4480,N_4303);
nor U6553 (N_6553,N_5389,N_5517);
or U6554 (N_6554,N_5395,N_4588);
xnor U6555 (N_6555,N_5616,N_5343);
and U6556 (N_6556,N_4356,N_5396);
xor U6557 (N_6557,N_5359,N_5036);
nand U6558 (N_6558,N_5756,N_4192);
and U6559 (N_6559,N_4278,N_5670);
or U6560 (N_6560,N_4405,N_5594);
and U6561 (N_6561,N_5093,N_4979);
xor U6562 (N_6562,N_4107,N_4886);
xor U6563 (N_6563,N_4142,N_4381);
xor U6564 (N_6564,N_5023,N_5701);
and U6565 (N_6565,N_4036,N_5133);
nand U6566 (N_6566,N_4752,N_5233);
nand U6567 (N_6567,N_4022,N_4640);
nand U6568 (N_6568,N_5325,N_4157);
and U6569 (N_6569,N_4483,N_5467);
or U6570 (N_6570,N_4643,N_5113);
xnor U6571 (N_6571,N_5269,N_4626);
and U6572 (N_6572,N_4496,N_4489);
and U6573 (N_6573,N_4918,N_4690);
or U6574 (N_6574,N_4892,N_4030);
and U6575 (N_6575,N_4338,N_4472);
or U6576 (N_6576,N_4345,N_5935);
or U6577 (N_6577,N_5024,N_4462);
nand U6578 (N_6578,N_4033,N_4382);
or U6579 (N_6579,N_4158,N_5130);
xnor U6580 (N_6580,N_4180,N_5640);
and U6581 (N_6581,N_5452,N_4875);
or U6582 (N_6582,N_4369,N_4726);
nor U6583 (N_6583,N_5826,N_5667);
xnor U6584 (N_6584,N_5047,N_5828);
nor U6585 (N_6585,N_5258,N_5971);
and U6586 (N_6586,N_5441,N_5891);
and U6587 (N_6587,N_4985,N_5243);
or U6588 (N_6588,N_5561,N_4722);
nor U6589 (N_6589,N_4216,N_4590);
and U6590 (N_6590,N_4600,N_5690);
nor U6591 (N_6591,N_5753,N_5154);
nor U6592 (N_6592,N_4646,N_4436);
xnor U6593 (N_6593,N_4943,N_4840);
or U6594 (N_6594,N_5873,N_4685);
xnor U6595 (N_6595,N_5266,N_4915);
xnor U6596 (N_6596,N_4651,N_4846);
or U6597 (N_6597,N_4994,N_5585);
or U6598 (N_6598,N_5507,N_5628);
nand U6599 (N_6599,N_5705,N_4645);
or U6600 (N_6600,N_4413,N_5552);
xor U6601 (N_6601,N_5484,N_5537);
nor U6602 (N_6602,N_5278,N_4719);
nor U6603 (N_6603,N_5059,N_5593);
nor U6604 (N_6604,N_5532,N_4485);
nor U6605 (N_6605,N_4532,N_4029);
and U6606 (N_6606,N_4281,N_4982);
and U6607 (N_6607,N_4221,N_5068);
or U6608 (N_6608,N_5687,N_4975);
nor U6609 (N_6609,N_5041,N_5481);
nand U6610 (N_6610,N_5353,N_4190);
and U6611 (N_6611,N_4758,N_5255);
nand U6612 (N_6612,N_5778,N_5995);
or U6613 (N_6613,N_4253,N_5157);
xnor U6614 (N_6614,N_4104,N_5310);
nor U6615 (N_6615,N_4204,N_5483);
nor U6616 (N_6616,N_4450,N_4503);
xnor U6617 (N_6617,N_4913,N_5992);
xnor U6618 (N_6618,N_4795,N_4096);
or U6619 (N_6619,N_4796,N_4743);
or U6620 (N_6620,N_4591,N_5675);
nand U6621 (N_6621,N_5367,N_4843);
xnor U6622 (N_6622,N_4045,N_5579);
nor U6623 (N_6623,N_4891,N_4053);
xor U6624 (N_6624,N_5478,N_4289);
xnor U6625 (N_6625,N_4904,N_4061);
nand U6626 (N_6626,N_4122,N_4510);
and U6627 (N_6627,N_5290,N_5280);
nand U6628 (N_6628,N_4136,N_4411);
nor U6629 (N_6629,N_4368,N_5963);
nor U6630 (N_6630,N_5492,N_5838);
nand U6631 (N_6631,N_5905,N_5214);
nor U6632 (N_6632,N_5542,N_5190);
nor U6633 (N_6633,N_4564,N_4803);
xor U6634 (N_6634,N_5669,N_5276);
nand U6635 (N_6635,N_5997,N_4858);
nand U6636 (N_6636,N_4537,N_4656);
nand U6637 (N_6637,N_5622,N_5646);
nor U6638 (N_6638,N_5978,N_4788);
or U6639 (N_6639,N_5656,N_4110);
xor U6640 (N_6640,N_4686,N_5052);
or U6641 (N_6641,N_4128,N_5011);
or U6642 (N_6642,N_4553,N_4860);
xnor U6643 (N_6643,N_4748,N_4733);
nor U6644 (N_6644,N_4861,N_5867);
or U6645 (N_6645,N_5348,N_4910);
xnor U6646 (N_6646,N_4453,N_4251);
and U6647 (N_6647,N_4946,N_4018);
or U6648 (N_6648,N_5298,N_5613);
or U6649 (N_6649,N_5924,N_5637);
and U6650 (N_6650,N_4696,N_4336);
or U6651 (N_6651,N_5879,N_4764);
and U6652 (N_6652,N_5790,N_4931);
xor U6653 (N_6653,N_4759,N_5878);
and U6654 (N_6654,N_5250,N_4611);
xor U6655 (N_6655,N_4962,N_4422);
and U6656 (N_6656,N_5364,N_4933);
xnor U6657 (N_6657,N_5122,N_4350);
nand U6658 (N_6658,N_4584,N_5263);
or U6659 (N_6659,N_4273,N_4465);
or U6660 (N_6660,N_5688,N_4851);
nor U6661 (N_6661,N_4402,N_5038);
nand U6662 (N_6662,N_5641,N_5918);
and U6663 (N_6663,N_4760,N_5020);
or U6664 (N_6664,N_5584,N_4015);
nand U6665 (N_6665,N_5668,N_5350);
nor U6666 (N_6666,N_4011,N_4282);
or U6667 (N_6667,N_4038,N_4566);
xnor U6668 (N_6668,N_5307,N_4406);
or U6669 (N_6669,N_4201,N_4585);
xor U6670 (N_6670,N_4705,N_4515);
or U6671 (N_6671,N_4493,N_4757);
nand U6672 (N_6672,N_5759,N_5486);
nand U6673 (N_6673,N_4188,N_5547);
nand U6674 (N_6674,N_5496,N_5683);
nand U6675 (N_6675,N_5293,N_4129);
nor U6676 (N_6676,N_5740,N_4953);
nand U6677 (N_6677,N_4019,N_4801);
xor U6678 (N_6678,N_4099,N_4009);
xnor U6679 (N_6679,N_4005,N_5877);
and U6680 (N_6680,N_4508,N_5804);
xnor U6681 (N_6681,N_5500,N_5844);
nor U6682 (N_6682,N_4055,N_5330);
nor U6683 (N_6683,N_4894,N_5192);
and U6684 (N_6684,N_5927,N_4821);
xor U6685 (N_6685,N_4424,N_4040);
nor U6686 (N_6686,N_5067,N_5393);
and U6687 (N_6687,N_4466,N_4390);
nor U6688 (N_6688,N_4706,N_4630);
and U6689 (N_6689,N_5741,N_5439);
or U6690 (N_6690,N_4427,N_4817);
xor U6691 (N_6691,N_5884,N_4527);
nor U6692 (N_6692,N_4961,N_5523);
nor U6693 (N_6693,N_4043,N_4100);
and U6694 (N_6694,N_5366,N_4186);
xor U6695 (N_6695,N_5319,N_4138);
nand U6696 (N_6696,N_5365,N_5351);
nor U6697 (N_6697,N_5627,N_5272);
and U6698 (N_6698,N_4444,N_5071);
xnor U6699 (N_6699,N_4414,N_4978);
and U6700 (N_6700,N_4728,N_4417);
xor U6701 (N_6701,N_4478,N_5787);
xnor U6702 (N_6702,N_4226,N_5265);
nor U6703 (N_6703,N_4621,N_4662);
nor U6704 (N_6704,N_5770,N_4003);
xor U6705 (N_6705,N_4106,N_4268);
or U6706 (N_6706,N_5777,N_4213);
or U6707 (N_6707,N_5568,N_4911);
nor U6708 (N_6708,N_4783,N_5715);
or U6709 (N_6709,N_4286,N_5711);
nand U6710 (N_6710,N_5134,N_5863);
and U6711 (N_6711,N_4191,N_4511);
xor U6712 (N_6712,N_5196,N_5171);
or U6713 (N_6713,N_4974,N_4569);
or U6714 (N_6714,N_5208,N_5271);
and U6715 (N_6715,N_4528,N_5762);
or U6716 (N_6716,N_5226,N_5013);
and U6717 (N_6717,N_4168,N_5062);
xor U6718 (N_6718,N_5698,N_5416);
or U6719 (N_6719,N_5820,N_5323);
nor U6720 (N_6720,N_5339,N_5306);
or U6721 (N_6721,N_5583,N_5572);
or U6722 (N_6722,N_5943,N_5070);
nand U6723 (N_6723,N_4103,N_4856);
nor U6724 (N_6724,N_5049,N_5806);
and U6725 (N_6725,N_4344,N_4986);
xor U6726 (N_6726,N_4529,N_5138);
and U6727 (N_6727,N_4628,N_5518);
and U6728 (N_6728,N_5257,N_4324);
nor U6729 (N_6729,N_5355,N_5607);
xor U6730 (N_6730,N_5662,N_5780);
nand U6731 (N_6731,N_4893,N_4866);
nand U6732 (N_6732,N_4665,N_4681);
xnor U6733 (N_6733,N_5944,N_4644);
nand U6734 (N_6734,N_4603,N_5959);
nand U6735 (N_6735,N_5842,N_5142);
nor U6736 (N_6736,N_5796,N_4037);
xor U6737 (N_6737,N_4660,N_4328);
nand U6738 (N_6738,N_4481,N_5743);
xor U6739 (N_6739,N_4069,N_4105);
nand U6740 (N_6740,N_4948,N_5016);
nor U6741 (N_6741,N_5578,N_4883);
xor U6742 (N_6742,N_4225,N_4415);
nand U6743 (N_6743,N_4949,N_5326);
nand U6744 (N_6744,N_4794,N_4842);
and U6745 (N_6745,N_5590,N_4077);
nor U6746 (N_6746,N_4650,N_4233);
nor U6747 (N_6747,N_5631,N_5764);
nand U6748 (N_6748,N_4010,N_5400);
nor U6749 (N_6749,N_4938,N_4395);
nand U6750 (N_6750,N_4362,N_5889);
xnor U6751 (N_6751,N_5981,N_4250);
and U6752 (N_6752,N_4865,N_4919);
or U6753 (N_6753,N_4775,N_4699);
and U6754 (N_6754,N_4908,N_5342);
nor U6755 (N_6755,N_5869,N_4081);
nor U6756 (N_6756,N_5936,N_4416);
or U6757 (N_6757,N_4315,N_4185);
nand U6758 (N_6758,N_4370,N_5075);
and U6759 (N_6759,N_4627,N_5610);
nand U6760 (N_6760,N_4346,N_5073);
and U6761 (N_6761,N_5901,N_4426);
nand U6762 (N_6762,N_5061,N_4461);
nand U6763 (N_6763,N_4687,N_4001);
nor U6764 (N_6764,N_4126,N_4602);
or U6765 (N_6765,N_5430,N_5026);
nor U6766 (N_6766,N_4765,N_5874);
or U6767 (N_6767,N_5917,N_5617);
nor U6768 (N_6768,N_5606,N_5458);
and U6769 (N_6769,N_5304,N_4357);
and U6770 (N_6770,N_5105,N_4027);
or U6771 (N_6771,N_5055,N_5429);
or U6772 (N_6772,N_5865,N_5642);
xor U6773 (N_6773,N_4737,N_4951);
or U6774 (N_6774,N_5139,N_4042);
nand U6775 (N_6775,N_4746,N_5892);
or U6776 (N_6776,N_5895,N_5308);
nand U6777 (N_6777,N_4217,N_5564);
or U6778 (N_6778,N_4888,N_4713);
or U6779 (N_6779,N_5019,N_5695);
xor U6780 (N_6780,N_4144,N_5219);
xnor U6781 (N_6781,N_5839,N_5213);
nand U6782 (N_6782,N_5468,N_5015);
nor U6783 (N_6783,N_5009,N_4321);
nor U6784 (N_6784,N_4215,N_5002);
and U6785 (N_6785,N_5881,N_4383);
and U6786 (N_6786,N_4683,N_4512);
and U6787 (N_6787,N_5937,N_5103);
nand U6788 (N_6788,N_4567,N_4288);
and U6789 (N_6789,N_4707,N_5750);
xnor U6790 (N_6790,N_4442,N_4448);
or U6791 (N_6791,N_4363,N_4329);
nor U6792 (N_6792,N_4826,N_5575);
xor U6793 (N_6793,N_4316,N_4610);
xor U6794 (N_6794,N_4127,N_4326);
xnor U6795 (N_6795,N_5338,N_5634);
nor U6796 (N_6796,N_4058,N_4309);
xor U6797 (N_6797,N_5371,N_5574);
nand U6798 (N_6798,N_4873,N_4773);
xnor U6799 (N_6799,N_5315,N_4041);
xnor U6800 (N_6800,N_5091,N_5758);
and U6801 (N_6801,N_4440,N_5980);
nand U6802 (N_6802,N_5736,N_5455);
or U6803 (N_6803,N_4594,N_4920);
nand U6804 (N_6804,N_4927,N_4820);
xnor U6805 (N_6805,N_4793,N_4237);
and U6806 (N_6806,N_5508,N_5057);
nor U6807 (N_6807,N_4672,N_4774);
or U6808 (N_6808,N_4025,N_5224);
nand U6809 (N_6809,N_4637,N_5054);
and U6810 (N_6810,N_4659,N_5645);
nor U6811 (N_6811,N_4968,N_5112);
nand U6812 (N_6812,N_4443,N_4469);
nor U6813 (N_6813,N_5569,N_4954);
nand U6814 (N_6814,N_5246,N_4148);
nor U6815 (N_6815,N_5781,N_4349);
nand U6816 (N_6816,N_5520,N_4475);
or U6817 (N_6817,N_4779,N_4302);
nor U6818 (N_6818,N_5198,N_5624);
and U6819 (N_6819,N_5141,N_5435);
nand U6820 (N_6820,N_4056,N_5555);
nand U6821 (N_6821,N_4163,N_4084);
and U6822 (N_6822,N_4618,N_5156);
nor U6823 (N_6823,N_5337,N_5116);
nand U6824 (N_6824,N_5684,N_4523);
and U6825 (N_6825,N_4864,N_4530);
nor U6826 (N_6826,N_4934,N_4708);
or U6827 (N_6827,N_5855,N_5608);
nand U6828 (N_6828,N_4083,N_4155);
xor U6829 (N_6829,N_5573,N_5792);
and U6830 (N_6830,N_4667,N_5849);
nand U6831 (N_6831,N_5816,N_5438);
nand U6832 (N_6832,N_5829,N_4398);
nand U6833 (N_6833,N_4070,N_4095);
or U6834 (N_6834,N_5072,N_5728);
xor U6835 (N_6835,N_5317,N_4880);
nand U6836 (N_6836,N_4990,N_4832);
nand U6837 (N_6837,N_4182,N_4937);
xnor U6838 (N_6838,N_4698,N_4712);
and U6839 (N_6839,N_4131,N_5313);
and U6840 (N_6840,N_5261,N_4745);
and U6841 (N_6841,N_4902,N_5379);
xnor U6842 (N_6842,N_4090,N_5005);
nand U6843 (N_6843,N_5516,N_4446);
nand U6844 (N_6844,N_5251,N_5489);
nor U6845 (N_6845,N_4007,N_5194);
nor U6846 (N_6846,N_4749,N_5286);
xor U6847 (N_6847,N_4807,N_4739);
nor U6848 (N_6848,N_5920,N_4334);
nor U6849 (N_6849,N_4008,N_4575);
nor U6850 (N_6850,N_4952,N_5949);
nor U6851 (N_6851,N_4140,N_4432);
or U6852 (N_6852,N_4265,N_5420);
xnor U6853 (N_6853,N_4689,N_4924);
nor U6854 (N_6854,N_5403,N_4548);
xnor U6855 (N_6855,N_4333,N_5202);
nor U6856 (N_6856,N_5785,N_4670);
nand U6857 (N_6857,N_5681,N_4074);
xnor U6858 (N_6858,N_4308,N_4762);
and U6859 (N_6859,N_4879,N_4463);
nor U6860 (N_6860,N_4804,N_5086);
xnor U6861 (N_6861,N_5615,N_4639);
xor U6862 (N_6862,N_5377,N_4340);
or U6863 (N_6863,N_4987,N_4184);
nor U6864 (N_6864,N_5004,N_4837);
or U6865 (N_6865,N_5228,N_4211);
or U6866 (N_6866,N_4239,N_5586);
nand U6867 (N_6867,N_5117,N_4717);
xnor U6868 (N_6868,N_5270,N_5394);
xor U6869 (N_6869,N_5721,N_5679);
xor U6870 (N_6870,N_4871,N_4963);
or U6871 (N_6871,N_4412,N_4364);
nor U6872 (N_6872,N_5368,N_5635);
xor U6873 (N_6873,N_5813,N_5505);
or U6874 (N_6874,N_5360,N_5620);
xor U6875 (N_6875,N_5238,N_5810);
and U6876 (N_6876,N_5823,N_4675);
nor U6877 (N_6877,N_4198,N_4115);
and U6878 (N_6878,N_4133,N_5577);
nand U6879 (N_6879,N_5473,N_5993);
xnor U6880 (N_6880,N_5525,N_5800);
or U6881 (N_6881,N_5254,N_4916);
xnor U6882 (N_6882,N_5653,N_5680);
xor U6883 (N_6883,N_4260,N_5819);
nand U6884 (N_6884,N_5249,N_5913);
and U6885 (N_6885,N_5528,N_5221);
nor U6886 (N_6886,N_4232,N_5952);
nor U6887 (N_6887,N_4477,N_4479);
or U6888 (N_6888,N_4721,N_4535);
and U6889 (N_6889,N_4972,N_4085);
nand U6890 (N_6890,N_5501,N_4763);
xnor U6891 (N_6891,N_4750,N_4261);
or U6892 (N_6892,N_5956,N_5053);
xor U6893 (N_6893,N_4725,N_4262);
nor U6894 (N_6894,N_5109,N_5294);
or U6895 (N_6895,N_4958,N_5494);
nor U6896 (N_6896,N_4679,N_4134);
and U6897 (N_6897,N_5786,N_4498);
nor U6898 (N_6898,N_4365,N_5256);
nor U6899 (N_6899,N_5419,N_4869);
or U6900 (N_6900,N_4800,N_5376);
nor U6901 (N_6901,N_5197,N_4714);
nand U6902 (N_6902,N_5223,N_4006);
or U6903 (N_6903,N_4825,N_5422);
and U6904 (N_6904,N_5106,N_4971);
or U6905 (N_6905,N_5301,N_5965);
nand U6906 (N_6906,N_5847,N_5530);
and U6907 (N_6907,N_5232,N_5536);
or U6908 (N_6908,N_4506,N_5673);
nor U6909 (N_6909,N_4827,N_4684);
and U6910 (N_6910,N_4212,N_5699);
nand U6911 (N_6911,N_5079,N_4181);
or U6912 (N_6912,N_4361,N_5734);
nand U6913 (N_6913,N_5488,N_4300);
nand U6914 (N_6914,N_4654,N_5230);
and U6915 (N_6915,N_4236,N_4822);
or U6916 (N_6916,N_5671,N_4926);
or U6917 (N_6917,N_5708,N_5209);
nor U6918 (N_6918,N_5953,N_4017);
nor U6919 (N_6919,N_5979,N_5215);
xor U6920 (N_6920,N_4504,N_5549);
or U6921 (N_6921,N_4220,N_5788);
nand U6922 (N_6922,N_5962,N_4841);
nand U6923 (N_6923,N_5911,N_4194);
nor U6924 (N_6924,N_4723,N_5589);
nand U6925 (N_6925,N_4407,N_5477);
nand U6926 (N_6926,N_4615,N_5700);
xor U6927 (N_6927,N_4117,N_4632);
nand U6928 (N_6928,N_5565,N_4993);
nand U6929 (N_6929,N_4495,N_5423);
nor U6930 (N_6930,N_4501,N_4139);
nor U6931 (N_6931,N_4536,N_5928);
and U6932 (N_6932,N_4735,N_5381);
and U6933 (N_6933,N_4544,N_4930);
and U6934 (N_6934,N_5289,N_4072);
xor U6935 (N_6935,N_5691,N_5167);
and U6936 (N_6936,N_5159,N_4109);
nand U6937 (N_6937,N_5693,N_5506);
and U6938 (N_6938,N_5510,N_5183);
and U6939 (N_6939,N_5275,N_5718);
or U6940 (N_6940,N_4206,N_5682);
xor U6941 (N_6941,N_4776,N_4353);
nor U6942 (N_6942,N_5697,N_5733);
nor U6943 (N_6943,N_4317,N_5629);
nand U6944 (N_6944,N_5191,N_5941);
nor U6945 (N_6945,N_4274,N_5179);
or U6946 (N_6946,N_4965,N_5907);
nor U6947 (N_6947,N_5871,N_4375);
xnor U6948 (N_6948,N_5175,N_5996);
and U6949 (N_6949,N_4063,N_5840);
xor U6950 (N_6950,N_4623,N_5652);
nand U6951 (N_6951,N_5789,N_4942);
xor U6952 (N_6952,N_4263,N_4857);
nand U6953 (N_6953,N_4476,N_4456);
or U6954 (N_6954,N_5066,N_5320);
nor U6955 (N_6955,N_5857,N_5114);
nand U6956 (N_6956,N_4162,N_5837);
and U6957 (N_6957,N_5136,N_5398);
and U6958 (N_6958,N_5210,N_5118);
nor U6959 (N_6959,N_5051,N_4352);
or U6960 (N_6960,N_4907,N_4021);
nand U6961 (N_6961,N_5972,N_5309);
and U6962 (N_6962,N_4899,N_4280);
and U6963 (N_6963,N_4923,N_5042);
nand U6964 (N_6964,N_5967,N_5783);
and U6965 (N_6965,N_5433,N_5449);
xor U6966 (N_6966,N_4950,N_4167);
nand U6967 (N_6967,N_5370,N_5127);
or U6968 (N_6968,N_4327,N_4189);
nand U6969 (N_6969,N_4421,N_5858);
or U6970 (N_6970,N_5580,N_4635);
xnor U6971 (N_6971,N_5706,N_5886);
xor U6972 (N_6972,N_4230,N_5203);
nand U6973 (N_6973,N_4756,N_5162);
nand U6974 (N_6974,N_5426,N_4579);
nand U6975 (N_6975,N_4772,N_5012);
and U6976 (N_6976,N_5237,N_5548);
nor U6977 (N_6977,N_5784,N_4231);
and U6978 (N_6978,N_5382,N_5211);
or U6979 (N_6979,N_4882,N_5852);
nand U6980 (N_6980,N_5618,N_4082);
xor U6981 (N_6981,N_5929,N_5322);
xor U6982 (N_6982,N_5689,N_5349);
nand U6983 (N_6983,N_5724,N_5513);
or U6984 (N_6984,N_5521,N_5825);
or U6985 (N_6985,N_4819,N_5921);
xnor U6986 (N_6986,N_5735,N_4319);
or U6987 (N_6987,N_5545,N_4246);
xnor U6988 (N_6988,N_5984,N_4094);
and U6989 (N_6989,N_5402,N_4132);
or U6990 (N_6990,N_5088,N_5014);
and U6991 (N_6991,N_4187,N_5973);
xor U6992 (N_6992,N_5745,N_5664);
xnor U6993 (N_6993,N_5883,N_4150);
and U6994 (N_6994,N_4655,N_5843);
xor U6995 (N_6995,N_5450,N_5087);
or U6996 (N_6996,N_4388,N_5390);
xnor U6997 (N_6997,N_4173,N_4314);
nor U6998 (N_6998,N_4568,N_5948);
nor U6999 (N_6999,N_4441,N_5830);
nand U7000 (N_7000,N_4938,N_4268);
nand U7001 (N_7001,N_5529,N_4344);
nor U7002 (N_7002,N_5905,N_5109);
and U7003 (N_7003,N_4030,N_5038);
or U7004 (N_7004,N_5677,N_4763);
and U7005 (N_7005,N_5172,N_5019);
nor U7006 (N_7006,N_4951,N_4512);
and U7007 (N_7007,N_4935,N_4198);
nand U7008 (N_7008,N_4458,N_5340);
xor U7009 (N_7009,N_4343,N_5107);
or U7010 (N_7010,N_5660,N_4037);
or U7011 (N_7011,N_5975,N_4501);
or U7012 (N_7012,N_4134,N_5566);
and U7013 (N_7013,N_4605,N_5037);
xnor U7014 (N_7014,N_5281,N_5265);
nand U7015 (N_7015,N_4208,N_4808);
or U7016 (N_7016,N_5430,N_4820);
and U7017 (N_7017,N_5543,N_4486);
xnor U7018 (N_7018,N_4823,N_5467);
and U7019 (N_7019,N_4596,N_4343);
and U7020 (N_7020,N_5320,N_4415);
and U7021 (N_7021,N_4434,N_5860);
or U7022 (N_7022,N_4665,N_5198);
nor U7023 (N_7023,N_4267,N_5557);
or U7024 (N_7024,N_5545,N_5468);
and U7025 (N_7025,N_4660,N_5617);
and U7026 (N_7026,N_5078,N_5699);
xnor U7027 (N_7027,N_4377,N_5776);
nand U7028 (N_7028,N_5183,N_4348);
nor U7029 (N_7029,N_4618,N_5981);
xnor U7030 (N_7030,N_4952,N_5034);
nor U7031 (N_7031,N_5636,N_5325);
and U7032 (N_7032,N_4396,N_5032);
and U7033 (N_7033,N_5455,N_5142);
xnor U7034 (N_7034,N_4563,N_4778);
and U7035 (N_7035,N_5709,N_5896);
nand U7036 (N_7036,N_5325,N_4393);
nand U7037 (N_7037,N_4096,N_5372);
nand U7038 (N_7038,N_4468,N_4700);
xnor U7039 (N_7039,N_5010,N_4297);
and U7040 (N_7040,N_4224,N_4707);
xor U7041 (N_7041,N_4584,N_4967);
and U7042 (N_7042,N_4310,N_5768);
nor U7043 (N_7043,N_5788,N_5504);
or U7044 (N_7044,N_5313,N_4958);
or U7045 (N_7045,N_5551,N_4107);
and U7046 (N_7046,N_4431,N_4059);
and U7047 (N_7047,N_4470,N_5832);
xor U7048 (N_7048,N_4242,N_5319);
or U7049 (N_7049,N_5425,N_4536);
nand U7050 (N_7050,N_5835,N_4522);
nand U7051 (N_7051,N_4019,N_5772);
and U7052 (N_7052,N_5127,N_4372);
or U7053 (N_7053,N_4001,N_5335);
nand U7054 (N_7054,N_4311,N_4844);
and U7055 (N_7055,N_5884,N_4738);
nand U7056 (N_7056,N_5949,N_4972);
nor U7057 (N_7057,N_4120,N_5289);
and U7058 (N_7058,N_4684,N_5879);
nor U7059 (N_7059,N_4129,N_4002);
nor U7060 (N_7060,N_5815,N_5661);
and U7061 (N_7061,N_4052,N_5385);
and U7062 (N_7062,N_4646,N_5973);
and U7063 (N_7063,N_5880,N_4268);
nor U7064 (N_7064,N_4748,N_4843);
xor U7065 (N_7065,N_5824,N_5992);
or U7066 (N_7066,N_5166,N_5143);
and U7067 (N_7067,N_5460,N_5876);
nand U7068 (N_7068,N_4014,N_5619);
nand U7069 (N_7069,N_4951,N_5955);
or U7070 (N_7070,N_5865,N_5186);
nor U7071 (N_7071,N_5183,N_5515);
nand U7072 (N_7072,N_5616,N_5130);
nand U7073 (N_7073,N_4791,N_4370);
and U7074 (N_7074,N_5450,N_5250);
xnor U7075 (N_7075,N_4457,N_5588);
nand U7076 (N_7076,N_5584,N_5474);
nand U7077 (N_7077,N_4796,N_5110);
nor U7078 (N_7078,N_4730,N_5713);
nand U7079 (N_7079,N_5462,N_4334);
xnor U7080 (N_7080,N_4637,N_5007);
nor U7081 (N_7081,N_4340,N_5056);
nor U7082 (N_7082,N_5616,N_5003);
nor U7083 (N_7083,N_5468,N_4838);
xnor U7084 (N_7084,N_4373,N_4116);
or U7085 (N_7085,N_5405,N_5348);
or U7086 (N_7086,N_4841,N_4977);
nand U7087 (N_7087,N_5650,N_5716);
nand U7088 (N_7088,N_4279,N_4566);
nand U7089 (N_7089,N_5054,N_4519);
or U7090 (N_7090,N_4962,N_4760);
or U7091 (N_7091,N_4430,N_4227);
xnor U7092 (N_7092,N_5496,N_5018);
xor U7093 (N_7093,N_5348,N_5741);
or U7094 (N_7094,N_5903,N_5848);
nor U7095 (N_7095,N_4567,N_5618);
nand U7096 (N_7096,N_4576,N_4903);
xor U7097 (N_7097,N_5140,N_5182);
nand U7098 (N_7098,N_5444,N_5417);
or U7099 (N_7099,N_4717,N_5004);
and U7100 (N_7100,N_4832,N_4345);
nor U7101 (N_7101,N_5185,N_4011);
xor U7102 (N_7102,N_4093,N_4203);
nand U7103 (N_7103,N_5936,N_4875);
xnor U7104 (N_7104,N_4388,N_5299);
xor U7105 (N_7105,N_4816,N_4054);
xnor U7106 (N_7106,N_4535,N_4245);
or U7107 (N_7107,N_4568,N_5670);
and U7108 (N_7108,N_5965,N_4689);
xor U7109 (N_7109,N_4778,N_5891);
or U7110 (N_7110,N_4265,N_4781);
xnor U7111 (N_7111,N_4537,N_4472);
or U7112 (N_7112,N_4104,N_5193);
and U7113 (N_7113,N_4490,N_4226);
nor U7114 (N_7114,N_4860,N_5000);
xor U7115 (N_7115,N_4116,N_5890);
nor U7116 (N_7116,N_5955,N_4174);
nor U7117 (N_7117,N_5726,N_4061);
nor U7118 (N_7118,N_4660,N_5839);
nor U7119 (N_7119,N_4437,N_4462);
xnor U7120 (N_7120,N_4035,N_4968);
nand U7121 (N_7121,N_4111,N_5645);
or U7122 (N_7122,N_4807,N_5159);
nor U7123 (N_7123,N_5938,N_5710);
and U7124 (N_7124,N_5544,N_5205);
nand U7125 (N_7125,N_4713,N_4848);
and U7126 (N_7126,N_5451,N_4610);
nor U7127 (N_7127,N_4673,N_5414);
or U7128 (N_7128,N_4721,N_4119);
and U7129 (N_7129,N_4699,N_4070);
and U7130 (N_7130,N_5201,N_4664);
or U7131 (N_7131,N_4816,N_4846);
xnor U7132 (N_7132,N_5231,N_5827);
and U7133 (N_7133,N_4598,N_4059);
nand U7134 (N_7134,N_5321,N_5454);
or U7135 (N_7135,N_4567,N_5827);
and U7136 (N_7136,N_5812,N_4838);
xor U7137 (N_7137,N_4244,N_5958);
xnor U7138 (N_7138,N_5408,N_5557);
and U7139 (N_7139,N_5409,N_4053);
and U7140 (N_7140,N_4375,N_5882);
and U7141 (N_7141,N_5175,N_4303);
or U7142 (N_7142,N_4780,N_4814);
nand U7143 (N_7143,N_5192,N_4845);
nor U7144 (N_7144,N_5575,N_5837);
and U7145 (N_7145,N_5387,N_4321);
nand U7146 (N_7146,N_5967,N_5341);
xor U7147 (N_7147,N_4102,N_4804);
nand U7148 (N_7148,N_4487,N_4802);
nand U7149 (N_7149,N_4255,N_4881);
or U7150 (N_7150,N_5042,N_5079);
xnor U7151 (N_7151,N_4405,N_4685);
xor U7152 (N_7152,N_5970,N_5352);
xnor U7153 (N_7153,N_4060,N_5585);
and U7154 (N_7154,N_5717,N_5590);
and U7155 (N_7155,N_5424,N_4499);
xnor U7156 (N_7156,N_4254,N_4463);
xnor U7157 (N_7157,N_5991,N_4882);
nand U7158 (N_7158,N_5302,N_4007);
and U7159 (N_7159,N_5855,N_4511);
or U7160 (N_7160,N_5406,N_4949);
nor U7161 (N_7161,N_5952,N_4846);
nand U7162 (N_7162,N_4980,N_5433);
nor U7163 (N_7163,N_4382,N_5172);
nand U7164 (N_7164,N_5713,N_5465);
or U7165 (N_7165,N_5779,N_4749);
xor U7166 (N_7166,N_5850,N_4111);
nand U7167 (N_7167,N_4036,N_5471);
nand U7168 (N_7168,N_5117,N_5139);
nor U7169 (N_7169,N_4858,N_4495);
nor U7170 (N_7170,N_4381,N_5767);
and U7171 (N_7171,N_5321,N_5292);
xor U7172 (N_7172,N_4709,N_5717);
nor U7173 (N_7173,N_4120,N_5017);
or U7174 (N_7174,N_4689,N_5391);
nor U7175 (N_7175,N_4903,N_5888);
or U7176 (N_7176,N_5966,N_5020);
nand U7177 (N_7177,N_5643,N_4775);
nor U7178 (N_7178,N_4458,N_4655);
or U7179 (N_7179,N_4237,N_5031);
and U7180 (N_7180,N_5080,N_4109);
xnor U7181 (N_7181,N_4146,N_5706);
xor U7182 (N_7182,N_5299,N_5568);
xnor U7183 (N_7183,N_4110,N_5337);
nor U7184 (N_7184,N_4064,N_5075);
or U7185 (N_7185,N_5381,N_5939);
xnor U7186 (N_7186,N_5874,N_5417);
nor U7187 (N_7187,N_4718,N_4801);
nand U7188 (N_7188,N_4363,N_4995);
nand U7189 (N_7189,N_4404,N_5845);
or U7190 (N_7190,N_4600,N_4798);
and U7191 (N_7191,N_5702,N_4290);
nand U7192 (N_7192,N_4042,N_5254);
xor U7193 (N_7193,N_5807,N_4068);
and U7194 (N_7194,N_4632,N_4938);
nand U7195 (N_7195,N_4775,N_5560);
or U7196 (N_7196,N_5102,N_4239);
xor U7197 (N_7197,N_4420,N_4726);
and U7198 (N_7198,N_5094,N_5036);
nor U7199 (N_7199,N_5393,N_5198);
nor U7200 (N_7200,N_4200,N_4014);
and U7201 (N_7201,N_5968,N_4459);
and U7202 (N_7202,N_4778,N_4186);
nor U7203 (N_7203,N_5146,N_5257);
nor U7204 (N_7204,N_5075,N_4854);
xnor U7205 (N_7205,N_4026,N_4627);
or U7206 (N_7206,N_4087,N_4106);
nand U7207 (N_7207,N_5507,N_5956);
nor U7208 (N_7208,N_5489,N_4923);
and U7209 (N_7209,N_5027,N_4957);
and U7210 (N_7210,N_4865,N_4599);
nand U7211 (N_7211,N_4492,N_5694);
nand U7212 (N_7212,N_4107,N_5323);
and U7213 (N_7213,N_4374,N_5084);
nand U7214 (N_7214,N_5070,N_4660);
xor U7215 (N_7215,N_5167,N_5072);
nand U7216 (N_7216,N_4251,N_4892);
and U7217 (N_7217,N_5386,N_5278);
xor U7218 (N_7218,N_5978,N_5324);
or U7219 (N_7219,N_5360,N_4876);
and U7220 (N_7220,N_4248,N_5818);
nand U7221 (N_7221,N_5056,N_4841);
xnor U7222 (N_7222,N_4865,N_4713);
nor U7223 (N_7223,N_5248,N_4593);
and U7224 (N_7224,N_4554,N_4002);
nand U7225 (N_7225,N_4271,N_4409);
nand U7226 (N_7226,N_4892,N_5803);
or U7227 (N_7227,N_5092,N_5597);
and U7228 (N_7228,N_5357,N_4640);
or U7229 (N_7229,N_4439,N_5267);
or U7230 (N_7230,N_5496,N_4686);
nand U7231 (N_7231,N_5497,N_4026);
and U7232 (N_7232,N_5524,N_4738);
xnor U7233 (N_7233,N_5468,N_5995);
and U7234 (N_7234,N_5061,N_5388);
nor U7235 (N_7235,N_5081,N_4555);
and U7236 (N_7236,N_5175,N_4863);
nand U7237 (N_7237,N_4003,N_5721);
and U7238 (N_7238,N_4760,N_5878);
nand U7239 (N_7239,N_5262,N_4090);
or U7240 (N_7240,N_5592,N_4755);
and U7241 (N_7241,N_5795,N_5782);
or U7242 (N_7242,N_5131,N_4543);
and U7243 (N_7243,N_4323,N_4801);
nand U7244 (N_7244,N_4549,N_4317);
and U7245 (N_7245,N_4738,N_5491);
nand U7246 (N_7246,N_4202,N_5358);
xnor U7247 (N_7247,N_4819,N_5509);
nor U7248 (N_7248,N_5164,N_4557);
and U7249 (N_7249,N_4228,N_5660);
nor U7250 (N_7250,N_5000,N_4176);
and U7251 (N_7251,N_5533,N_5902);
and U7252 (N_7252,N_4654,N_4689);
and U7253 (N_7253,N_5204,N_4194);
nand U7254 (N_7254,N_4223,N_4702);
xnor U7255 (N_7255,N_5814,N_4101);
and U7256 (N_7256,N_4545,N_4566);
nand U7257 (N_7257,N_5776,N_4091);
nor U7258 (N_7258,N_5969,N_5539);
and U7259 (N_7259,N_4645,N_5981);
xnor U7260 (N_7260,N_5176,N_4878);
and U7261 (N_7261,N_4217,N_5954);
xor U7262 (N_7262,N_5455,N_5502);
or U7263 (N_7263,N_5468,N_4402);
nor U7264 (N_7264,N_5201,N_4107);
nor U7265 (N_7265,N_4374,N_4454);
nand U7266 (N_7266,N_5611,N_4303);
xor U7267 (N_7267,N_4177,N_5870);
and U7268 (N_7268,N_4072,N_5699);
nor U7269 (N_7269,N_5858,N_5350);
nor U7270 (N_7270,N_4270,N_4953);
and U7271 (N_7271,N_5163,N_5867);
and U7272 (N_7272,N_4083,N_5871);
or U7273 (N_7273,N_5951,N_4987);
or U7274 (N_7274,N_4136,N_4820);
or U7275 (N_7275,N_4105,N_4656);
xor U7276 (N_7276,N_4783,N_4429);
nand U7277 (N_7277,N_5305,N_5386);
nand U7278 (N_7278,N_4934,N_4552);
nand U7279 (N_7279,N_4630,N_5320);
and U7280 (N_7280,N_4113,N_5280);
xnor U7281 (N_7281,N_4206,N_4676);
and U7282 (N_7282,N_4027,N_5753);
or U7283 (N_7283,N_5344,N_5416);
nor U7284 (N_7284,N_4936,N_5386);
nor U7285 (N_7285,N_4470,N_4047);
nor U7286 (N_7286,N_4581,N_5587);
or U7287 (N_7287,N_4958,N_5296);
nor U7288 (N_7288,N_5141,N_5160);
nand U7289 (N_7289,N_4160,N_4045);
and U7290 (N_7290,N_4887,N_5720);
nand U7291 (N_7291,N_4692,N_4905);
or U7292 (N_7292,N_4346,N_5819);
nand U7293 (N_7293,N_5267,N_4285);
nor U7294 (N_7294,N_4141,N_5405);
xnor U7295 (N_7295,N_4291,N_4842);
xor U7296 (N_7296,N_4291,N_5337);
xor U7297 (N_7297,N_4391,N_5082);
or U7298 (N_7298,N_5751,N_4050);
xnor U7299 (N_7299,N_4062,N_4380);
and U7300 (N_7300,N_5364,N_5360);
and U7301 (N_7301,N_5997,N_4257);
or U7302 (N_7302,N_4995,N_4026);
nor U7303 (N_7303,N_5225,N_4527);
xor U7304 (N_7304,N_5982,N_4285);
nor U7305 (N_7305,N_4892,N_4432);
and U7306 (N_7306,N_5659,N_5206);
xor U7307 (N_7307,N_4070,N_4931);
nor U7308 (N_7308,N_5871,N_5883);
and U7309 (N_7309,N_5834,N_5809);
and U7310 (N_7310,N_5720,N_4435);
and U7311 (N_7311,N_5461,N_4721);
nand U7312 (N_7312,N_5862,N_4778);
nand U7313 (N_7313,N_4550,N_4450);
or U7314 (N_7314,N_5802,N_5250);
nor U7315 (N_7315,N_4642,N_5689);
and U7316 (N_7316,N_5582,N_4672);
xnor U7317 (N_7317,N_5843,N_4555);
nor U7318 (N_7318,N_5211,N_4353);
and U7319 (N_7319,N_5692,N_5413);
xnor U7320 (N_7320,N_4889,N_5559);
and U7321 (N_7321,N_5316,N_4483);
xor U7322 (N_7322,N_4818,N_4213);
or U7323 (N_7323,N_5022,N_5218);
or U7324 (N_7324,N_4134,N_5060);
nand U7325 (N_7325,N_4511,N_4591);
and U7326 (N_7326,N_5405,N_4448);
nor U7327 (N_7327,N_5884,N_4725);
and U7328 (N_7328,N_4184,N_5878);
and U7329 (N_7329,N_5525,N_5544);
nor U7330 (N_7330,N_5765,N_4201);
and U7331 (N_7331,N_4748,N_5891);
nor U7332 (N_7332,N_5563,N_5074);
xnor U7333 (N_7333,N_5689,N_5014);
and U7334 (N_7334,N_4219,N_4018);
and U7335 (N_7335,N_4844,N_4538);
and U7336 (N_7336,N_5552,N_4836);
or U7337 (N_7337,N_4551,N_4038);
xor U7338 (N_7338,N_5456,N_4150);
nor U7339 (N_7339,N_4300,N_5426);
or U7340 (N_7340,N_5594,N_5345);
xor U7341 (N_7341,N_5155,N_4475);
nand U7342 (N_7342,N_4938,N_5343);
nand U7343 (N_7343,N_4503,N_4133);
xor U7344 (N_7344,N_5226,N_5488);
or U7345 (N_7345,N_4361,N_5789);
xnor U7346 (N_7346,N_5109,N_5219);
and U7347 (N_7347,N_4224,N_5772);
xor U7348 (N_7348,N_5983,N_4703);
or U7349 (N_7349,N_4676,N_4294);
nor U7350 (N_7350,N_5553,N_4721);
xor U7351 (N_7351,N_5077,N_5939);
and U7352 (N_7352,N_5395,N_4884);
xnor U7353 (N_7353,N_4300,N_5576);
nor U7354 (N_7354,N_4873,N_5671);
and U7355 (N_7355,N_5236,N_5491);
nand U7356 (N_7356,N_5723,N_5063);
nor U7357 (N_7357,N_4091,N_5997);
or U7358 (N_7358,N_5387,N_5988);
or U7359 (N_7359,N_4785,N_5583);
or U7360 (N_7360,N_5128,N_4026);
nand U7361 (N_7361,N_4783,N_5114);
or U7362 (N_7362,N_4921,N_4087);
or U7363 (N_7363,N_5002,N_5824);
xor U7364 (N_7364,N_5349,N_4590);
or U7365 (N_7365,N_5815,N_4016);
or U7366 (N_7366,N_5876,N_4944);
or U7367 (N_7367,N_5371,N_4054);
xor U7368 (N_7368,N_4295,N_4210);
or U7369 (N_7369,N_4597,N_4619);
or U7370 (N_7370,N_5017,N_5787);
xnor U7371 (N_7371,N_5822,N_4362);
nor U7372 (N_7372,N_4145,N_5293);
or U7373 (N_7373,N_4657,N_5241);
nor U7374 (N_7374,N_5003,N_4660);
and U7375 (N_7375,N_4924,N_5346);
or U7376 (N_7376,N_5058,N_4523);
xor U7377 (N_7377,N_5139,N_5065);
nand U7378 (N_7378,N_5875,N_4430);
xnor U7379 (N_7379,N_5966,N_4522);
nand U7380 (N_7380,N_5991,N_5407);
nor U7381 (N_7381,N_5758,N_4705);
xor U7382 (N_7382,N_4300,N_4052);
xor U7383 (N_7383,N_4302,N_5833);
xor U7384 (N_7384,N_5571,N_5156);
xnor U7385 (N_7385,N_5448,N_5497);
nand U7386 (N_7386,N_5908,N_4616);
xnor U7387 (N_7387,N_5890,N_4087);
xor U7388 (N_7388,N_5925,N_5691);
or U7389 (N_7389,N_4792,N_5062);
xnor U7390 (N_7390,N_4113,N_4120);
and U7391 (N_7391,N_4771,N_4202);
xor U7392 (N_7392,N_5209,N_4971);
nand U7393 (N_7393,N_5217,N_5255);
or U7394 (N_7394,N_4559,N_4369);
nor U7395 (N_7395,N_4689,N_4024);
nor U7396 (N_7396,N_5657,N_5677);
nor U7397 (N_7397,N_5622,N_4305);
nand U7398 (N_7398,N_5225,N_5129);
and U7399 (N_7399,N_5949,N_5842);
nor U7400 (N_7400,N_5001,N_4423);
or U7401 (N_7401,N_4410,N_5584);
nor U7402 (N_7402,N_4902,N_4450);
nand U7403 (N_7403,N_5623,N_5020);
or U7404 (N_7404,N_5450,N_5771);
nor U7405 (N_7405,N_4109,N_5637);
nand U7406 (N_7406,N_5199,N_5295);
nor U7407 (N_7407,N_4479,N_5946);
or U7408 (N_7408,N_4062,N_4667);
and U7409 (N_7409,N_5056,N_5335);
and U7410 (N_7410,N_5348,N_5634);
nand U7411 (N_7411,N_4403,N_5418);
nand U7412 (N_7412,N_4947,N_5234);
nor U7413 (N_7413,N_5214,N_5704);
xnor U7414 (N_7414,N_4916,N_4222);
and U7415 (N_7415,N_5136,N_5549);
nor U7416 (N_7416,N_5400,N_5410);
nor U7417 (N_7417,N_5463,N_4198);
nor U7418 (N_7418,N_5944,N_4519);
nor U7419 (N_7419,N_5664,N_5369);
nand U7420 (N_7420,N_5265,N_5881);
nand U7421 (N_7421,N_4764,N_5307);
and U7422 (N_7422,N_5163,N_4234);
nor U7423 (N_7423,N_5463,N_5291);
nand U7424 (N_7424,N_4837,N_4416);
nand U7425 (N_7425,N_4845,N_5822);
xor U7426 (N_7426,N_5861,N_4377);
nand U7427 (N_7427,N_4222,N_5811);
and U7428 (N_7428,N_4012,N_4561);
and U7429 (N_7429,N_4221,N_5122);
or U7430 (N_7430,N_4261,N_5866);
xnor U7431 (N_7431,N_4212,N_4484);
xor U7432 (N_7432,N_5353,N_5510);
xnor U7433 (N_7433,N_5862,N_4027);
and U7434 (N_7434,N_5140,N_4380);
nor U7435 (N_7435,N_4958,N_4316);
nand U7436 (N_7436,N_4147,N_4641);
xnor U7437 (N_7437,N_5167,N_5223);
xor U7438 (N_7438,N_4610,N_5407);
and U7439 (N_7439,N_5956,N_5633);
nor U7440 (N_7440,N_4122,N_4249);
nand U7441 (N_7441,N_5198,N_4101);
and U7442 (N_7442,N_4880,N_4774);
and U7443 (N_7443,N_4333,N_4744);
xnor U7444 (N_7444,N_5447,N_5611);
nand U7445 (N_7445,N_4982,N_5671);
or U7446 (N_7446,N_5996,N_4549);
or U7447 (N_7447,N_5579,N_4341);
xor U7448 (N_7448,N_4173,N_4601);
nand U7449 (N_7449,N_5443,N_4877);
or U7450 (N_7450,N_5074,N_4029);
and U7451 (N_7451,N_4221,N_5727);
and U7452 (N_7452,N_4603,N_5563);
xnor U7453 (N_7453,N_5343,N_5035);
or U7454 (N_7454,N_5247,N_4969);
nor U7455 (N_7455,N_4515,N_5803);
or U7456 (N_7456,N_5840,N_4658);
nor U7457 (N_7457,N_4141,N_4661);
or U7458 (N_7458,N_5058,N_4710);
xnor U7459 (N_7459,N_5758,N_4472);
xor U7460 (N_7460,N_5666,N_4807);
xor U7461 (N_7461,N_4671,N_5054);
xnor U7462 (N_7462,N_4943,N_4402);
nand U7463 (N_7463,N_4016,N_5885);
nand U7464 (N_7464,N_4550,N_4917);
nand U7465 (N_7465,N_4938,N_4277);
nor U7466 (N_7466,N_4606,N_4029);
nand U7467 (N_7467,N_5772,N_4294);
nand U7468 (N_7468,N_4422,N_5008);
nand U7469 (N_7469,N_5702,N_5115);
and U7470 (N_7470,N_4753,N_5114);
nand U7471 (N_7471,N_4039,N_5489);
nand U7472 (N_7472,N_4082,N_5036);
and U7473 (N_7473,N_5403,N_5367);
nor U7474 (N_7474,N_5861,N_5188);
xor U7475 (N_7475,N_5130,N_4050);
or U7476 (N_7476,N_4908,N_4901);
or U7477 (N_7477,N_4771,N_4323);
nor U7478 (N_7478,N_5846,N_4298);
nand U7479 (N_7479,N_4965,N_5522);
nor U7480 (N_7480,N_4910,N_4594);
and U7481 (N_7481,N_4582,N_4194);
and U7482 (N_7482,N_5963,N_4824);
nand U7483 (N_7483,N_4219,N_5300);
and U7484 (N_7484,N_4779,N_4372);
nand U7485 (N_7485,N_4361,N_5485);
or U7486 (N_7486,N_5070,N_5630);
or U7487 (N_7487,N_5127,N_5431);
and U7488 (N_7488,N_4078,N_5304);
xor U7489 (N_7489,N_4550,N_5644);
nand U7490 (N_7490,N_4146,N_4058);
or U7491 (N_7491,N_4885,N_5647);
and U7492 (N_7492,N_5325,N_5347);
and U7493 (N_7493,N_5914,N_4859);
nor U7494 (N_7494,N_4861,N_5619);
xor U7495 (N_7495,N_4830,N_4420);
and U7496 (N_7496,N_4746,N_4442);
xnor U7497 (N_7497,N_4629,N_5885);
and U7498 (N_7498,N_5803,N_5817);
nor U7499 (N_7499,N_4377,N_4509);
nor U7500 (N_7500,N_4858,N_5599);
or U7501 (N_7501,N_5086,N_5189);
nor U7502 (N_7502,N_4218,N_4191);
and U7503 (N_7503,N_4880,N_4229);
nand U7504 (N_7504,N_5778,N_5044);
nor U7505 (N_7505,N_5977,N_5419);
nand U7506 (N_7506,N_4948,N_5416);
and U7507 (N_7507,N_4513,N_5180);
nand U7508 (N_7508,N_4443,N_5545);
nor U7509 (N_7509,N_4319,N_5324);
nor U7510 (N_7510,N_4010,N_4044);
or U7511 (N_7511,N_4265,N_5363);
xor U7512 (N_7512,N_4046,N_5936);
nor U7513 (N_7513,N_5683,N_5913);
nor U7514 (N_7514,N_4083,N_5425);
or U7515 (N_7515,N_5453,N_5817);
and U7516 (N_7516,N_4337,N_5171);
nor U7517 (N_7517,N_5846,N_5336);
and U7518 (N_7518,N_5434,N_5706);
xor U7519 (N_7519,N_5339,N_4155);
or U7520 (N_7520,N_5105,N_5262);
nor U7521 (N_7521,N_5119,N_4494);
xnor U7522 (N_7522,N_5412,N_5377);
nand U7523 (N_7523,N_5763,N_5827);
nand U7524 (N_7524,N_5658,N_4832);
or U7525 (N_7525,N_5826,N_5014);
xnor U7526 (N_7526,N_5736,N_4722);
xor U7527 (N_7527,N_4814,N_5114);
and U7528 (N_7528,N_4780,N_5460);
nor U7529 (N_7529,N_4420,N_4292);
or U7530 (N_7530,N_5024,N_4194);
and U7531 (N_7531,N_5888,N_5913);
nand U7532 (N_7532,N_4870,N_4920);
nor U7533 (N_7533,N_5732,N_5222);
and U7534 (N_7534,N_4059,N_4269);
nor U7535 (N_7535,N_4363,N_5123);
or U7536 (N_7536,N_4471,N_5939);
xnor U7537 (N_7537,N_4037,N_5122);
or U7538 (N_7538,N_5485,N_4053);
or U7539 (N_7539,N_5817,N_5295);
nand U7540 (N_7540,N_4622,N_5654);
nand U7541 (N_7541,N_4590,N_4558);
nand U7542 (N_7542,N_5228,N_4274);
nor U7543 (N_7543,N_4593,N_4400);
nor U7544 (N_7544,N_4572,N_4559);
nand U7545 (N_7545,N_4189,N_4138);
nand U7546 (N_7546,N_4642,N_4602);
and U7547 (N_7547,N_5078,N_4620);
or U7548 (N_7548,N_5972,N_5548);
nor U7549 (N_7549,N_4747,N_5427);
and U7550 (N_7550,N_4940,N_4872);
nand U7551 (N_7551,N_5477,N_5738);
and U7552 (N_7552,N_5056,N_4964);
nor U7553 (N_7553,N_5041,N_4334);
nor U7554 (N_7554,N_4287,N_5997);
nand U7555 (N_7555,N_4947,N_4282);
xor U7556 (N_7556,N_4411,N_5946);
nor U7557 (N_7557,N_5122,N_4316);
or U7558 (N_7558,N_4648,N_5740);
and U7559 (N_7559,N_5123,N_4972);
xnor U7560 (N_7560,N_4677,N_4108);
or U7561 (N_7561,N_5222,N_4630);
or U7562 (N_7562,N_4986,N_5374);
and U7563 (N_7563,N_5784,N_4682);
nand U7564 (N_7564,N_4599,N_5525);
or U7565 (N_7565,N_5785,N_4930);
and U7566 (N_7566,N_4970,N_5695);
xor U7567 (N_7567,N_5523,N_5702);
nand U7568 (N_7568,N_4018,N_5475);
nand U7569 (N_7569,N_4213,N_5523);
or U7570 (N_7570,N_5635,N_5295);
and U7571 (N_7571,N_4003,N_4508);
nand U7572 (N_7572,N_5229,N_4033);
nand U7573 (N_7573,N_4490,N_4447);
and U7574 (N_7574,N_5419,N_4213);
nand U7575 (N_7575,N_4007,N_5106);
xnor U7576 (N_7576,N_5598,N_4615);
nand U7577 (N_7577,N_5833,N_5022);
and U7578 (N_7578,N_5834,N_4217);
or U7579 (N_7579,N_4066,N_4213);
or U7580 (N_7580,N_4334,N_5587);
xnor U7581 (N_7581,N_4805,N_4123);
or U7582 (N_7582,N_5468,N_4667);
nor U7583 (N_7583,N_4851,N_5551);
nor U7584 (N_7584,N_4961,N_4655);
and U7585 (N_7585,N_5230,N_5986);
nand U7586 (N_7586,N_4441,N_5536);
nor U7587 (N_7587,N_4979,N_5569);
and U7588 (N_7588,N_5829,N_5885);
nand U7589 (N_7589,N_5778,N_4655);
and U7590 (N_7590,N_4068,N_4095);
or U7591 (N_7591,N_4620,N_4320);
xor U7592 (N_7592,N_4660,N_4933);
xor U7593 (N_7593,N_5219,N_5428);
and U7594 (N_7594,N_5652,N_4347);
or U7595 (N_7595,N_4474,N_5731);
nor U7596 (N_7596,N_4011,N_5926);
xor U7597 (N_7597,N_4743,N_4994);
or U7598 (N_7598,N_5924,N_4031);
nand U7599 (N_7599,N_5636,N_4086);
xnor U7600 (N_7600,N_4621,N_4155);
and U7601 (N_7601,N_4914,N_5196);
nor U7602 (N_7602,N_5598,N_5493);
nand U7603 (N_7603,N_5433,N_4813);
and U7604 (N_7604,N_5260,N_4342);
and U7605 (N_7605,N_5618,N_5444);
and U7606 (N_7606,N_5145,N_5315);
nor U7607 (N_7607,N_4920,N_4945);
nor U7608 (N_7608,N_5902,N_5308);
nand U7609 (N_7609,N_4476,N_5446);
and U7610 (N_7610,N_4020,N_5414);
nor U7611 (N_7611,N_4379,N_4514);
nor U7612 (N_7612,N_5830,N_5836);
or U7613 (N_7613,N_5320,N_5874);
nand U7614 (N_7614,N_4069,N_4243);
and U7615 (N_7615,N_5843,N_4760);
xnor U7616 (N_7616,N_4189,N_5817);
nor U7617 (N_7617,N_5918,N_5492);
nor U7618 (N_7618,N_4700,N_5712);
nor U7619 (N_7619,N_5886,N_4715);
and U7620 (N_7620,N_4520,N_5573);
nand U7621 (N_7621,N_4162,N_4475);
nor U7622 (N_7622,N_4241,N_4501);
and U7623 (N_7623,N_5613,N_4003);
and U7624 (N_7624,N_4872,N_4924);
nand U7625 (N_7625,N_5744,N_4676);
nand U7626 (N_7626,N_4481,N_4215);
and U7627 (N_7627,N_5557,N_4922);
xnor U7628 (N_7628,N_5659,N_4620);
and U7629 (N_7629,N_4236,N_4324);
nand U7630 (N_7630,N_5291,N_4960);
and U7631 (N_7631,N_4236,N_4794);
nand U7632 (N_7632,N_4837,N_4881);
nand U7633 (N_7633,N_4814,N_5225);
nand U7634 (N_7634,N_4422,N_4423);
and U7635 (N_7635,N_5514,N_5320);
and U7636 (N_7636,N_5152,N_5197);
nor U7637 (N_7637,N_4625,N_5782);
xnor U7638 (N_7638,N_5641,N_4162);
and U7639 (N_7639,N_5827,N_4483);
and U7640 (N_7640,N_5660,N_4363);
xor U7641 (N_7641,N_5984,N_4250);
or U7642 (N_7642,N_4469,N_4333);
or U7643 (N_7643,N_4803,N_5062);
and U7644 (N_7644,N_5863,N_4807);
nor U7645 (N_7645,N_4838,N_4102);
nor U7646 (N_7646,N_4065,N_5461);
nor U7647 (N_7647,N_5378,N_4015);
and U7648 (N_7648,N_5993,N_5476);
nand U7649 (N_7649,N_5465,N_4800);
or U7650 (N_7650,N_4720,N_4990);
xnor U7651 (N_7651,N_5264,N_5554);
or U7652 (N_7652,N_5587,N_5904);
and U7653 (N_7653,N_4865,N_5977);
nand U7654 (N_7654,N_4451,N_5370);
nand U7655 (N_7655,N_4675,N_5931);
xnor U7656 (N_7656,N_5622,N_4609);
nand U7657 (N_7657,N_4871,N_5443);
nand U7658 (N_7658,N_5206,N_5497);
nand U7659 (N_7659,N_5468,N_4762);
nor U7660 (N_7660,N_5141,N_4182);
and U7661 (N_7661,N_5222,N_5595);
nor U7662 (N_7662,N_4356,N_5037);
nor U7663 (N_7663,N_5526,N_5679);
and U7664 (N_7664,N_4778,N_5139);
and U7665 (N_7665,N_5584,N_4391);
nand U7666 (N_7666,N_5757,N_4183);
or U7667 (N_7667,N_5227,N_4895);
xnor U7668 (N_7668,N_4214,N_5728);
xnor U7669 (N_7669,N_5617,N_4826);
and U7670 (N_7670,N_4840,N_4001);
nand U7671 (N_7671,N_4951,N_5610);
nor U7672 (N_7672,N_5214,N_5398);
xnor U7673 (N_7673,N_5390,N_5186);
nand U7674 (N_7674,N_4345,N_4602);
nand U7675 (N_7675,N_5211,N_4787);
xnor U7676 (N_7676,N_4733,N_4466);
or U7677 (N_7677,N_4315,N_5617);
and U7678 (N_7678,N_5550,N_5806);
or U7679 (N_7679,N_5057,N_4585);
xor U7680 (N_7680,N_4929,N_4990);
or U7681 (N_7681,N_4096,N_5919);
or U7682 (N_7682,N_5669,N_5445);
xnor U7683 (N_7683,N_5180,N_5761);
nand U7684 (N_7684,N_4464,N_4981);
nand U7685 (N_7685,N_4881,N_4906);
nor U7686 (N_7686,N_5877,N_4788);
or U7687 (N_7687,N_5506,N_5472);
or U7688 (N_7688,N_5807,N_4149);
nand U7689 (N_7689,N_5364,N_5420);
xnor U7690 (N_7690,N_5134,N_5627);
xnor U7691 (N_7691,N_5630,N_5219);
or U7692 (N_7692,N_4585,N_5951);
nand U7693 (N_7693,N_4234,N_5586);
xor U7694 (N_7694,N_5656,N_4556);
nand U7695 (N_7695,N_5245,N_4104);
xor U7696 (N_7696,N_4481,N_5904);
nand U7697 (N_7697,N_5813,N_5542);
nand U7698 (N_7698,N_5195,N_5920);
and U7699 (N_7699,N_5897,N_4034);
or U7700 (N_7700,N_5563,N_5831);
xnor U7701 (N_7701,N_4485,N_5202);
or U7702 (N_7702,N_5756,N_5427);
and U7703 (N_7703,N_5305,N_4620);
xnor U7704 (N_7704,N_4910,N_4038);
nor U7705 (N_7705,N_4676,N_5974);
nor U7706 (N_7706,N_5379,N_4355);
or U7707 (N_7707,N_4339,N_5558);
nor U7708 (N_7708,N_4931,N_4764);
and U7709 (N_7709,N_4039,N_5963);
nand U7710 (N_7710,N_5063,N_4290);
nor U7711 (N_7711,N_4559,N_4554);
xor U7712 (N_7712,N_5928,N_5075);
nor U7713 (N_7713,N_4211,N_5140);
xor U7714 (N_7714,N_5626,N_5733);
or U7715 (N_7715,N_4437,N_5527);
nand U7716 (N_7716,N_5109,N_4577);
nand U7717 (N_7717,N_5722,N_4634);
nand U7718 (N_7718,N_4476,N_4006);
and U7719 (N_7719,N_5727,N_4593);
xor U7720 (N_7720,N_4194,N_4462);
and U7721 (N_7721,N_5056,N_5064);
nor U7722 (N_7722,N_4288,N_5556);
nand U7723 (N_7723,N_4410,N_5927);
nor U7724 (N_7724,N_4610,N_5438);
or U7725 (N_7725,N_5772,N_4536);
or U7726 (N_7726,N_5682,N_4643);
and U7727 (N_7727,N_5500,N_4210);
xor U7728 (N_7728,N_4101,N_5625);
nor U7729 (N_7729,N_5892,N_4797);
and U7730 (N_7730,N_5570,N_5321);
and U7731 (N_7731,N_4809,N_4901);
and U7732 (N_7732,N_4164,N_4287);
or U7733 (N_7733,N_5878,N_5304);
and U7734 (N_7734,N_4212,N_5902);
nor U7735 (N_7735,N_4027,N_4788);
or U7736 (N_7736,N_5793,N_5148);
and U7737 (N_7737,N_4804,N_5736);
nand U7738 (N_7738,N_4209,N_4072);
nor U7739 (N_7739,N_4152,N_4194);
and U7740 (N_7740,N_4921,N_4609);
nand U7741 (N_7741,N_4723,N_4053);
nor U7742 (N_7742,N_5126,N_4338);
nor U7743 (N_7743,N_4255,N_5754);
nand U7744 (N_7744,N_5482,N_5340);
nand U7745 (N_7745,N_4198,N_4083);
or U7746 (N_7746,N_5940,N_5821);
and U7747 (N_7747,N_5770,N_4358);
and U7748 (N_7748,N_5765,N_5158);
nand U7749 (N_7749,N_5913,N_5464);
or U7750 (N_7750,N_5255,N_5916);
and U7751 (N_7751,N_5081,N_5097);
or U7752 (N_7752,N_5877,N_5452);
xnor U7753 (N_7753,N_5965,N_4789);
or U7754 (N_7754,N_5212,N_5952);
xnor U7755 (N_7755,N_4759,N_5206);
or U7756 (N_7756,N_5229,N_5644);
or U7757 (N_7757,N_5749,N_5935);
nor U7758 (N_7758,N_4833,N_4966);
xnor U7759 (N_7759,N_5348,N_5029);
nand U7760 (N_7760,N_4873,N_4348);
xor U7761 (N_7761,N_5840,N_4374);
and U7762 (N_7762,N_5597,N_4900);
and U7763 (N_7763,N_5867,N_5842);
nand U7764 (N_7764,N_4301,N_5929);
nand U7765 (N_7765,N_4984,N_5786);
nand U7766 (N_7766,N_5381,N_4866);
and U7767 (N_7767,N_5633,N_4467);
xor U7768 (N_7768,N_5209,N_4281);
and U7769 (N_7769,N_4429,N_5273);
xor U7770 (N_7770,N_5436,N_5398);
nor U7771 (N_7771,N_4924,N_4844);
or U7772 (N_7772,N_5368,N_5173);
or U7773 (N_7773,N_4170,N_5055);
and U7774 (N_7774,N_4846,N_5926);
nand U7775 (N_7775,N_4629,N_4360);
xor U7776 (N_7776,N_5304,N_5482);
and U7777 (N_7777,N_4569,N_5524);
nor U7778 (N_7778,N_5203,N_4606);
and U7779 (N_7779,N_5331,N_5070);
and U7780 (N_7780,N_5152,N_4347);
and U7781 (N_7781,N_5434,N_4299);
nor U7782 (N_7782,N_5138,N_5767);
nor U7783 (N_7783,N_4348,N_5726);
nand U7784 (N_7784,N_5546,N_5086);
or U7785 (N_7785,N_4588,N_4319);
xnor U7786 (N_7786,N_4373,N_4345);
and U7787 (N_7787,N_4924,N_4690);
xnor U7788 (N_7788,N_4364,N_5832);
nor U7789 (N_7789,N_4471,N_4374);
nand U7790 (N_7790,N_5840,N_5768);
nor U7791 (N_7791,N_5341,N_5265);
nand U7792 (N_7792,N_5903,N_4524);
and U7793 (N_7793,N_5324,N_5179);
nand U7794 (N_7794,N_4250,N_4191);
and U7795 (N_7795,N_4264,N_4627);
nand U7796 (N_7796,N_5489,N_4689);
nor U7797 (N_7797,N_4533,N_4686);
and U7798 (N_7798,N_4409,N_4004);
nand U7799 (N_7799,N_5059,N_4040);
and U7800 (N_7800,N_5433,N_5916);
or U7801 (N_7801,N_4257,N_5036);
and U7802 (N_7802,N_4869,N_5214);
nand U7803 (N_7803,N_4746,N_5915);
nor U7804 (N_7804,N_5993,N_4738);
nor U7805 (N_7805,N_4228,N_4992);
or U7806 (N_7806,N_5960,N_5277);
and U7807 (N_7807,N_5490,N_5745);
nand U7808 (N_7808,N_5493,N_5921);
or U7809 (N_7809,N_4562,N_4367);
nor U7810 (N_7810,N_5517,N_5170);
and U7811 (N_7811,N_5816,N_5745);
xnor U7812 (N_7812,N_5448,N_5051);
nor U7813 (N_7813,N_5643,N_4157);
or U7814 (N_7814,N_4429,N_5805);
xnor U7815 (N_7815,N_5901,N_5418);
xnor U7816 (N_7816,N_5591,N_5101);
nor U7817 (N_7817,N_4662,N_5462);
and U7818 (N_7818,N_4316,N_5938);
or U7819 (N_7819,N_5509,N_4679);
or U7820 (N_7820,N_5799,N_4014);
nand U7821 (N_7821,N_5063,N_5061);
or U7822 (N_7822,N_4801,N_4597);
xnor U7823 (N_7823,N_4136,N_4527);
and U7824 (N_7824,N_5757,N_4329);
and U7825 (N_7825,N_4385,N_4423);
nand U7826 (N_7826,N_5462,N_4635);
nor U7827 (N_7827,N_4839,N_4356);
nor U7828 (N_7828,N_4725,N_5526);
and U7829 (N_7829,N_5219,N_4444);
xor U7830 (N_7830,N_4484,N_5990);
and U7831 (N_7831,N_4463,N_5558);
and U7832 (N_7832,N_5556,N_5271);
nand U7833 (N_7833,N_4725,N_5795);
xnor U7834 (N_7834,N_5745,N_4340);
and U7835 (N_7835,N_4242,N_5444);
or U7836 (N_7836,N_4712,N_5266);
xnor U7837 (N_7837,N_4250,N_5119);
or U7838 (N_7838,N_5764,N_5197);
nor U7839 (N_7839,N_5034,N_4161);
xor U7840 (N_7840,N_5467,N_5021);
xnor U7841 (N_7841,N_4771,N_5153);
and U7842 (N_7842,N_4145,N_4846);
nor U7843 (N_7843,N_5293,N_5632);
or U7844 (N_7844,N_4932,N_5750);
nand U7845 (N_7845,N_5263,N_5047);
and U7846 (N_7846,N_4464,N_5239);
nor U7847 (N_7847,N_4127,N_5641);
and U7848 (N_7848,N_4525,N_4538);
and U7849 (N_7849,N_5190,N_4637);
xnor U7850 (N_7850,N_4874,N_5250);
nor U7851 (N_7851,N_5136,N_4791);
and U7852 (N_7852,N_4478,N_5291);
and U7853 (N_7853,N_5712,N_4286);
nand U7854 (N_7854,N_5258,N_5444);
nor U7855 (N_7855,N_5449,N_5405);
and U7856 (N_7856,N_5903,N_4487);
xor U7857 (N_7857,N_4931,N_4195);
xnor U7858 (N_7858,N_4478,N_4201);
nor U7859 (N_7859,N_4128,N_5826);
nand U7860 (N_7860,N_4950,N_5711);
nand U7861 (N_7861,N_4178,N_5353);
and U7862 (N_7862,N_5340,N_5269);
or U7863 (N_7863,N_5298,N_4273);
and U7864 (N_7864,N_4424,N_5310);
xor U7865 (N_7865,N_5380,N_5069);
xnor U7866 (N_7866,N_4173,N_4492);
xor U7867 (N_7867,N_5229,N_5196);
nand U7868 (N_7868,N_5687,N_5189);
or U7869 (N_7869,N_5816,N_4121);
and U7870 (N_7870,N_4804,N_4233);
nand U7871 (N_7871,N_4429,N_5539);
nand U7872 (N_7872,N_4477,N_5019);
nor U7873 (N_7873,N_4585,N_5343);
nor U7874 (N_7874,N_4051,N_5058);
xnor U7875 (N_7875,N_5056,N_4452);
xor U7876 (N_7876,N_4669,N_4433);
nand U7877 (N_7877,N_4511,N_5861);
and U7878 (N_7878,N_5802,N_5729);
nor U7879 (N_7879,N_4760,N_5148);
xor U7880 (N_7880,N_4042,N_4270);
xor U7881 (N_7881,N_4583,N_4883);
and U7882 (N_7882,N_4631,N_4449);
nor U7883 (N_7883,N_5950,N_4936);
xor U7884 (N_7884,N_4428,N_5555);
nand U7885 (N_7885,N_4653,N_5908);
and U7886 (N_7886,N_5658,N_5684);
or U7887 (N_7887,N_4917,N_5739);
nand U7888 (N_7888,N_4282,N_5100);
or U7889 (N_7889,N_5350,N_4329);
or U7890 (N_7890,N_4605,N_4523);
xor U7891 (N_7891,N_5971,N_5253);
or U7892 (N_7892,N_5103,N_4738);
nand U7893 (N_7893,N_4702,N_5973);
and U7894 (N_7894,N_4890,N_5669);
nor U7895 (N_7895,N_4880,N_5810);
nand U7896 (N_7896,N_5183,N_5987);
and U7897 (N_7897,N_5133,N_5937);
nand U7898 (N_7898,N_5902,N_4529);
nor U7899 (N_7899,N_4355,N_4446);
and U7900 (N_7900,N_5246,N_5334);
nand U7901 (N_7901,N_4317,N_5934);
and U7902 (N_7902,N_4170,N_5487);
xor U7903 (N_7903,N_4390,N_5713);
nand U7904 (N_7904,N_5157,N_4780);
nand U7905 (N_7905,N_4216,N_4258);
and U7906 (N_7906,N_4789,N_4134);
nor U7907 (N_7907,N_5424,N_5582);
and U7908 (N_7908,N_5747,N_4857);
nand U7909 (N_7909,N_5490,N_4084);
and U7910 (N_7910,N_4090,N_5762);
and U7911 (N_7911,N_5061,N_4234);
xnor U7912 (N_7912,N_5396,N_4375);
and U7913 (N_7913,N_5627,N_5070);
and U7914 (N_7914,N_5964,N_5962);
nor U7915 (N_7915,N_4078,N_5752);
or U7916 (N_7916,N_4504,N_4287);
and U7917 (N_7917,N_5767,N_5036);
or U7918 (N_7918,N_4006,N_5706);
xnor U7919 (N_7919,N_5705,N_5932);
xnor U7920 (N_7920,N_4686,N_5186);
or U7921 (N_7921,N_5104,N_5284);
and U7922 (N_7922,N_5312,N_5367);
or U7923 (N_7923,N_5414,N_5935);
xnor U7924 (N_7924,N_5693,N_5218);
and U7925 (N_7925,N_5937,N_4295);
nor U7926 (N_7926,N_4073,N_5253);
nand U7927 (N_7927,N_5523,N_4128);
or U7928 (N_7928,N_5610,N_4407);
xnor U7929 (N_7929,N_4236,N_5031);
and U7930 (N_7930,N_5521,N_5068);
xnor U7931 (N_7931,N_4779,N_4190);
nor U7932 (N_7932,N_4868,N_4032);
xnor U7933 (N_7933,N_4625,N_4823);
nand U7934 (N_7934,N_5696,N_5913);
and U7935 (N_7935,N_5546,N_5149);
and U7936 (N_7936,N_5378,N_5929);
and U7937 (N_7937,N_4955,N_5133);
or U7938 (N_7938,N_5034,N_4731);
nor U7939 (N_7939,N_5792,N_5012);
nor U7940 (N_7940,N_5456,N_5655);
or U7941 (N_7941,N_5427,N_4376);
and U7942 (N_7942,N_5492,N_4484);
or U7943 (N_7943,N_5014,N_5992);
xor U7944 (N_7944,N_4627,N_4157);
and U7945 (N_7945,N_5456,N_4805);
and U7946 (N_7946,N_5743,N_5201);
and U7947 (N_7947,N_4814,N_4968);
nand U7948 (N_7948,N_4824,N_4526);
nor U7949 (N_7949,N_4627,N_5880);
and U7950 (N_7950,N_4451,N_4022);
nand U7951 (N_7951,N_5038,N_5848);
and U7952 (N_7952,N_4674,N_4339);
or U7953 (N_7953,N_5908,N_5536);
xor U7954 (N_7954,N_5619,N_5677);
nand U7955 (N_7955,N_4436,N_4103);
and U7956 (N_7956,N_4824,N_5440);
xor U7957 (N_7957,N_4878,N_5968);
xor U7958 (N_7958,N_5753,N_5536);
nor U7959 (N_7959,N_4813,N_5116);
nand U7960 (N_7960,N_5161,N_4626);
or U7961 (N_7961,N_4290,N_4446);
nor U7962 (N_7962,N_4007,N_4652);
and U7963 (N_7963,N_4604,N_5013);
and U7964 (N_7964,N_5529,N_4315);
and U7965 (N_7965,N_4433,N_4118);
and U7966 (N_7966,N_5309,N_5481);
nor U7967 (N_7967,N_4439,N_4021);
nor U7968 (N_7968,N_5407,N_5051);
and U7969 (N_7969,N_5830,N_4984);
nor U7970 (N_7970,N_5146,N_5161);
xor U7971 (N_7971,N_4950,N_4937);
nand U7972 (N_7972,N_4599,N_4172);
and U7973 (N_7973,N_4077,N_4154);
nand U7974 (N_7974,N_5897,N_4350);
or U7975 (N_7975,N_5455,N_5253);
nand U7976 (N_7976,N_5571,N_4684);
xor U7977 (N_7977,N_5280,N_5149);
and U7978 (N_7978,N_5054,N_5503);
or U7979 (N_7979,N_4791,N_5877);
and U7980 (N_7980,N_5716,N_4884);
nand U7981 (N_7981,N_4332,N_4711);
and U7982 (N_7982,N_4740,N_5878);
nand U7983 (N_7983,N_5968,N_4847);
nor U7984 (N_7984,N_5192,N_4030);
and U7985 (N_7985,N_5029,N_5551);
nor U7986 (N_7986,N_4883,N_5502);
nor U7987 (N_7987,N_4886,N_5926);
nand U7988 (N_7988,N_4605,N_5855);
xnor U7989 (N_7989,N_5417,N_4444);
and U7990 (N_7990,N_5727,N_5978);
nor U7991 (N_7991,N_5345,N_4314);
nand U7992 (N_7992,N_4425,N_5051);
nor U7993 (N_7993,N_5514,N_5745);
xnor U7994 (N_7994,N_4596,N_5029);
and U7995 (N_7995,N_4185,N_4241);
and U7996 (N_7996,N_4338,N_4706);
nor U7997 (N_7997,N_4439,N_5360);
or U7998 (N_7998,N_5228,N_5106);
nor U7999 (N_7999,N_4968,N_5239);
and U8000 (N_8000,N_6913,N_7268);
nor U8001 (N_8001,N_6749,N_7193);
nor U8002 (N_8002,N_6510,N_7617);
nand U8003 (N_8003,N_6147,N_7367);
nand U8004 (N_8004,N_6944,N_7350);
nor U8005 (N_8005,N_6728,N_6567);
xnor U8006 (N_8006,N_7642,N_7124);
nand U8007 (N_8007,N_6844,N_7245);
and U8008 (N_8008,N_7991,N_6186);
nor U8009 (N_8009,N_6921,N_6910);
or U8010 (N_8010,N_7799,N_7498);
or U8011 (N_8011,N_6899,N_6055);
xnor U8012 (N_8012,N_7577,N_7125);
and U8013 (N_8013,N_7242,N_7394);
nand U8014 (N_8014,N_7345,N_6314);
xnor U8015 (N_8015,N_7397,N_6941);
nor U8016 (N_8016,N_6650,N_6018);
and U8017 (N_8017,N_6908,N_7916);
xnor U8018 (N_8018,N_7385,N_7552);
or U8019 (N_8019,N_6383,N_6570);
xnor U8020 (N_8020,N_6402,N_7536);
and U8021 (N_8021,N_6995,N_7770);
nand U8022 (N_8022,N_7418,N_6025);
nor U8023 (N_8023,N_6451,N_6571);
nor U8024 (N_8024,N_6107,N_6263);
and U8025 (N_8025,N_6460,N_6133);
nand U8026 (N_8026,N_6699,N_7514);
or U8027 (N_8027,N_7836,N_6445);
nor U8028 (N_8028,N_7297,N_6869);
or U8029 (N_8029,N_6351,N_6824);
nor U8030 (N_8030,N_6439,N_6686);
or U8031 (N_8031,N_6931,N_7704);
xnor U8032 (N_8032,N_6333,N_6523);
nor U8033 (N_8033,N_7290,N_7884);
and U8034 (N_8034,N_6750,N_6718);
and U8035 (N_8035,N_7275,N_7671);
nor U8036 (N_8036,N_6323,N_6034);
or U8037 (N_8037,N_6374,N_7669);
and U8038 (N_8038,N_7547,N_6932);
nand U8039 (N_8039,N_6377,N_6244);
xnor U8040 (N_8040,N_7389,N_7187);
xor U8041 (N_8041,N_6796,N_7220);
or U8042 (N_8042,N_6030,N_6215);
xor U8043 (N_8043,N_7155,N_7545);
nor U8044 (N_8044,N_7171,N_7630);
xor U8045 (N_8045,N_7833,N_6836);
xnor U8046 (N_8046,N_6717,N_6363);
and U8047 (N_8047,N_7056,N_6493);
nor U8048 (N_8048,N_6057,N_7148);
or U8049 (N_8049,N_6959,N_7018);
nand U8050 (N_8050,N_7743,N_6403);
and U8051 (N_8051,N_6662,N_6741);
xor U8052 (N_8052,N_6894,N_6066);
nand U8053 (N_8053,N_7004,N_7601);
nor U8054 (N_8054,N_6070,N_6754);
or U8055 (N_8055,N_6652,N_6211);
and U8056 (N_8056,N_7249,N_7925);
nor U8057 (N_8057,N_6457,N_6840);
and U8058 (N_8058,N_7771,N_7428);
or U8059 (N_8059,N_7106,N_7184);
nand U8060 (N_8060,N_6655,N_6121);
or U8061 (N_8061,N_7113,N_7908);
nand U8062 (N_8062,N_7659,N_6256);
nor U8063 (N_8063,N_6350,N_7570);
nand U8064 (N_8064,N_7595,N_7938);
and U8065 (N_8065,N_6349,N_7217);
and U8066 (N_8066,N_6587,N_7892);
and U8067 (N_8067,N_6243,N_6809);
or U8068 (N_8068,N_6605,N_7431);
nand U8069 (N_8069,N_7519,N_7083);
or U8070 (N_8070,N_6636,N_6156);
or U8071 (N_8071,N_7639,N_7383);
and U8072 (N_8072,N_7696,N_6812);
or U8073 (N_8073,N_7543,N_6731);
nor U8074 (N_8074,N_7751,N_7172);
or U8075 (N_8075,N_7827,N_7014);
and U8076 (N_8076,N_6723,N_6250);
xor U8077 (N_8077,N_7561,N_6238);
nor U8078 (N_8078,N_7854,N_7824);
nor U8079 (N_8079,N_7086,N_6416);
or U8080 (N_8080,N_6278,N_6001);
nand U8081 (N_8081,N_7537,N_7831);
nand U8082 (N_8082,N_7323,N_7948);
and U8083 (N_8083,N_6930,N_6659);
and U8084 (N_8084,N_7594,N_6409);
xnor U8085 (N_8085,N_7711,N_6434);
and U8086 (N_8086,N_6837,N_6372);
xnor U8087 (N_8087,N_6893,N_7352);
and U8088 (N_8088,N_7997,N_7044);
xnor U8089 (N_8089,N_6863,N_6775);
xor U8090 (N_8090,N_6562,N_7301);
or U8091 (N_8091,N_6142,N_6850);
nor U8092 (N_8092,N_7463,N_7645);
nor U8093 (N_8093,N_7666,N_6617);
xor U8094 (N_8094,N_7979,N_6239);
nand U8095 (N_8095,N_7413,N_6230);
and U8096 (N_8096,N_6739,N_6534);
or U8097 (N_8097,N_6481,N_6786);
nor U8098 (N_8098,N_7282,N_7493);
nor U8099 (N_8099,N_7952,N_6037);
nand U8100 (N_8100,N_7214,N_7749);
or U8101 (N_8101,N_7656,N_7073);
nand U8102 (N_8102,N_7729,N_6900);
and U8103 (N_8103,N_6705,N_7528);
nor U8104 (N_8104,N_6233,N_6252);
and U8105 (N_8105,N_6407,N_7538);
and U8106 (N_8106,N_6572,N_6242);
or U8107 (N_8107,N_7093,N_7091);
nor U8108 (N_8108,N_6014,N_7660);
xnor U8109 (N_8109,N_7199,N_7551);
xnor U8110 (N_8110,N_6656,N_6385);
or U8111 (N_8111,N_6581,N_6588);
or U8112 (N_8112,N_6952,N_6148);
or U8113 (N_8113,N_6956,N_6648);
nand U8114 (N_8114,N_7655,N_6890);
nand U8115 (N_8115,N_7638,N_7706);
and U8116 (N_8116,N_7949,N_7364);
nor U8117 (N_8117,N_7472,N_6074);
xnor U8118 (N_8118,N_6499,N_7135);
nand U8119 (N_8119,N_6294,N_6821);
nor U8120 (N_8120,N_6543,N_7393);
xor U8121 (N_8121,N_6738,N_6110);
xor U8122 (N_8122,N_6486,N_7310);
xnor U8123 (N_8123,N_7374,N_6473);
nand U8124 (N_8124,N_6024,N_7255);
nand U8125 (N_8125,N_6906,N_7196);
nand U8126 (N_8126,N_7508,N_7340);
nand U8127 (N_8127,N_6094,N_7085);
and U8128 (N_8128,N_6404,N_6764);
nor U8129 (N_8129,N_7975,N_7777);
or U8130 (N_8130,N_7879,N_6820);
nand U8131 (N_8131,N_6266,N_7795);
nand U8132 (N_8132,N_6180,N_7988);
xor U8133 (N_8133,N_6261,N_7930);
nor U8134 (N_8134,N_6756,N_6971);
nor U8135 (N_8135,N_6545,N_6803);
nor U8136 (N_8136,N_6847,N_6702);
nand U8137 (N_8137,N_6725,N_7679);
and U8138 (N_8138,N_7286,N_6965);
nand U8139 (N_8139,N_6732,N_7410);
xnor U8140 (N_8140,N_6124,N_7969);
xor U8141 (N_8141,N_7684,N_6068);
and U8142 (N_8142,N_7865,N_6284);
xnor U8143 (N_8143,N_7610,N_7919);
nor U8144 (N_8144,N_6139,N_6685);
or U8145 (N_8145,N_7848,N_7238);
nand U8146 (N_8146,N_7998,N_6022);
and U8147 (N_8147,N_7661,N_7077);
or U8148 (N_8148,N_7134,N_6815);
and U8149 (N_8149,N_6283,N_7246);
nand U8150 (N_8150,N_6287,N_6841);
xnor U8151 (N_8151,N_6277,N_7976);
or U8152 (N_8152,N_6199,N_6524);
nor U8153 (N_8153,N_7548,N_6084);
nor U8154 (N_8154,N_6217,N_7276);
xor U8155 (N_8155,N_7072,N_7980);
and U8156 (N_8156,N_7596,N_7046);
nor U8157 (N_8157,N_7181,N_6787);
or U8158 (N_8158,N_7120,N_7070);
and U8159 (N_8159,N_7223,N_7691);
xnor U8160 (N_8160,N_7424,N_6131);
and U8161 (N_8161,N_6067,N_6989);
nor U8162 (N_8162,N_6637,N_6979);
xnor U8163 (N_8163,N_6802,N_7445);
and U8164 (N_8164,N_6673,N_6414);
nor U8165 (N_8165,N_7226,N_7562);
nand U8166 (N_8166,N_7259,N_7612);
and U8167 (N_8167,N_7504,N_6173);
nor U8168 (N_8168,N_7296,N_6376);
or U8169 (N_8169,N_6682,N_6538);
nand U8170 (N_8170,N_7168,N_6661);
nand U8171 (N_8171,N_7872,N_6390);
nand U8172 (N_8172,N_7312,N_6794);
nand U8173 (N_8173,N_6257,N_7423);
and U8174 (N_8174,N_6663,N_7623);
or U8175 (N_8175,N_6059,N_7037);
or U8176 (N_8176,N_6969,N_7745);
xor U8177 (N_8177,N_6942,N_6479);
nor U8178 (N_8178,N_7675,N_7322);
nor U8179 (N_8179,N_7657,N_7859);
xor U8180 (N_8180,N_6429,N_6565);
xnor U8181 (N_8181,N_6957,N_6514);
xor U8182 (N_8182,N_7897,N_6053);
or U8183 (N_8183,N_6209,N_7447);
or U8184 (N_8184,N_6255,N_6964);
or U8185 (N_8185,N_6099,N_7420);
xnor U8186 (N_8186,N_6861,N_6146);
or U8187 (N_8187,N_7329,N_6365);
or U8188 (N_8188,N_7235,N_7721);
and U8189 (N_8189,N_6619,N_6370);
xnor U8190 (N_8190,N_6128,N_6483);
xor U8191 (N_8191,N_7328,N_6010);
nand U8192 (N_8192,N_6399,N_7588);
xor U8193 (N_8193,N_7990,N_7355);
nand U8194 (N_8194,N_7597,N_6842);
nand U8195 (N_8195,N_7989,N_7754);
nand U8196 (N_8196,N_6496,N_7392);
nor U8197 (N_8197,N_6838,N_6219);
xnor U8198 (N_8198,N_7287,N_7057);
nand U8199 (N_8199,N_7593,N_7400);
or U8200 (N_8200,N_6886,N_7280);
or U8201 (N_8201,N_6624,N_7169);
or U8202 (N_8202,N_6462,N_6651);
nand U8203 (N_8203,N_6017,N_6553);
nand U8204 (N_8204,N_7146,N_6202);
and U8205 (N_8205,N_6270,N_7521);
nand U8206 (N_8206,N_7198,N_7643);
or U8207 (N_8207,N_6746,N_6996);
and U8208 (N_8208,N_6081,N_6688);
or U8209 (N_8209,N_7294,N_6785);
xor U8210 (N_8210,N_7417,N_7186);
xor U8211 (N_8211,N_6225,N_7794);
nor U8212 (N_8212,N_6406,N_7421);
or U8213 (N_8213,N_6293,N_7395);
or U8214 (N_8214,N_7730,N_6159);
nand U8215 (N_8215,N_7658,N_6212);
nor U8216 (N_8216,N_7587,N_6143);
xor U8217 (N_8217,N_7358,N_7183);
and U8218 (N_8218,N_6367,N_6945);
and U8219 (N_8219,N_6733,N_6231);
xnor U8220 (N_8220,N_6320,N_6246);
or U8221 (N_8221,N_6911,N_7152);
or U8222 (N_8222,N_6990,N_7786);
nor U8223 (N_8223,N_7133,N_6623);
xor U8224 (N_8224,N_6751,N_7663);
xor U8225 (N_8225,N_7864,N_6031);
xnor U8226 (N_8226,N_7550,N_6338);
nor U8227 (N_8227,N_6129,N_6249);
nand U8228 (N_8228,N_7111,N_7667);
nor U8229 (N_8229,N_6340,N_6526);
xor U8230 (N_8230,N_7986,N_6214);
nor U8231 (N_8231,N_6719,N_7909);
xnor U8232 (N_8232,N_7614,N_7869);
nand U8233 (N_8233,N_6606,N_7703);
nand U8234 (N_8234,N_7019,N_7629);
and U8235 (N_8235,N_7026,N_7775);
or U8236 (N_8236,N_7160,N_7518);
nand U8237 (N_8237,N_6771,N_7132);
xnor U8238 (N_8238,N_7260,N_6817);
or U8239 (N_8239,N_7441,N_6985);
nor U8240 (N_8240,N_6026,N_7122);
and U8241 (N_8241,N_6634,N_7257);
or U8242 (N_8242,N_7142,N_6192);
and U8243 (N_8243,N_7103,N_6105);
or U8244 (N_8244,N_7460,N_6912);
nand U8245 (N_8245,N_7946,N_6917);
and U8246 (N_8246,N_6715,N_7603);
nor U8247 (N_8247,N_7676,N_7708);
nand U8248 (N_8248,N_6568,N_6830);
nor U8249 (N_8249,N_6851,N_6477);
nand U8250 (N_8250,N_7945,N_6926);
xnor U8251 (N_8251,N_6345,N_7839);
nand U8252 (N_8252,N_7935,N_6378);
nor U8253 (N_8253,N_7698,N_6454);
nand U8254 (N_8254,N_7736,N_6806);
nand U8255 (N_8255,N_6324,N_7632);
and U8256 (N_8256,N_6355,N_6521);
and U8257 (N_8257,N_7499,N_7448);
nand U8258 (N_8258,N_6576,N_6282);
or U8259 (N_8259,N_6210,N_7572);
xnor U8260 (N_8260,N_7201,N_6308);
nand U8261 (N_8261,N_6229,N_7524);
nand U8262 (N_8262,N_7497,N_6127);
nand U8263 (N_8263,N_6152,N_7295);
xor U8264 (N_8264,N_7654,N_6469);
or U8265 (N_8265,N_6613,N_7112);
and U8266 (N_8266,N_7608,N_7313);
nand U8267 (N_8267,N_6674,N_6115);
and U8268 (N_8268,N_6177,N_6714);
or U8269 (N_8269,N_7722,N_6729);
nand U8270 (N_8270,N_7525,N_6466);
xor U8271 (N_8271,N_7531,N_6927);
and U8272 (N_8272,N_7856,N_6111);
nand U8273 (N_8273,N_6801,N_7564);
and U8274 (N_8274,N_6835,N_7893);
nor U8275 (N_8275,N_6860,N_7241);
and U8276 (N_8276,N_7810,N_6958);
and U8277 (N_8277,N_7584,N_7375);
xnor U8278 (N_8278,N_6042,N_7779);
nand U8279 (N_8279,N_7953,N_7918);
nand U8280 (N_8280,N_6972,N_7163);
nand U8281 (N_8281,N_6792,N_7024);
and U8282 (N_8282,N_7816,N_7955);
or U8283 (N_8283,N_7549,N_6864);
nand U8284 (N_8284,N_6175,N_6168);
nand U8285 (N_8285,N_6819,N_7150);
xor U8286 (N_8286,N_7911,N_6566);
nor U8287 (N_8287,N_6816,N_7141);
nor U8288 (N_8288,N_6833,N_7422);
nand U8289 (N_8289,N_7047,N_6788);
or U8290 (N_8290,N_6694,N_7049);
or U8291 (N_8291,N_6316,N_6050);
nor U8292 (N_8292,N_7407,N_6432);
nor U8293 (N_8293,N_6218,N_6716);
nand U8294 (N_8294,N_7672,N_6144);
or U8295 (N_8295,N_6155,N_7359);
or U8296 (N_8296,N_7715,N_6870);
and U8297 (N_8297,N_7624,N_6698);
nand U8298 (N_8298,N_6991,N_7067);
nand U8299 (N_8299,N_7641,N_7759);
xor U8300 (N_8300,N_6875,N_7211);
and U8301 (N_8301,N_6839,N_7347);
or U8302 (N_8302,N_7139,N_7003);
xnor U8303 (N_8303,N_6504,N_6446);
nor U8304 (N_8304,N_6450,N_7600);
xnor U8305 (N_8305,N_7533,N_6398);
and U8306 (N_8306,N_6896,N_7559);
or U8307 (N_8307,N_7923,N_7899);
and U8308 (N_8308,N_6807,N_6391);
xor U8309 (N_8309,N_6118,N_6003);
and U8310 (N_8310,N_6711,N_6923);
xor U8311 (N_8311,N_7127,N_7941);
xnor U8312 (N_8312,N_6734,N_6895);
or U8313 (N_8313,N_7118,N_6411);
nand U8314 (N_8314,N_7495,N_6354);
nand U8315 (N_8315,N_6339,N_6343);
nand U8316 (N_8316,N_7331,N_7351);
or U8317 (N_8317,N_6914,N_7109);
nand U8318 (N_8318,N_6268,N_6500);
nor U8319 (N_8319,N_6922,N_6664);
nor U8320 (N_8320,N_7651,N_7688);
nand U8321 (N_8321,N_6721,N_7627);
xor U8322 (N_8322,N_6043,N_7228);
xor U8323 (N_8323,N_6119,N_7012);
nor U8324 (N_8324,N_7857,N_6428);
nor U8325 (N_8325,N_7811,N_7076);
nor U8326 (N_8326,N_7905,N_6799);
nand U8327 (N_8327,N_7471,N_7457);
xnor U8328 (N_8328,N_7291,N_6488);
nor U8329 (N_8329,N_7088,N_7677);
and U8330 (N_8330,N_7804,N_7089);
nor U8331 (N_8331,N_7232,N_7720);
xor U8332 (N_8332,N_6130,N_6038);
or U8333 (N_8333,N_6328,N_7693);
or U8334 (N_8334,N_6396,N_6936);
nor U8335 (N_8335,N_6831,N_6963);
and U8336 (N_8336,N_6978,N_6464);
nor U8337 (N_8337,N_6061,N_6184);
and U8338 (N_8338,N_6907,N_7732);
nor U8339 (N_8339,N_7269,N_7903);
nand U8340 (N_8340,N_6549,N_6480);
and U8341 (N_8341,N_7311,N_7866);
nor U8342 (N_8342,N_6049,N_6056);
and U8343 (N_8343,N_6271,N_7568);
xnor U8344 (N_8344,N_6440,N_7818);
and U8345 (N_8345,N_6435,N_6665);
xnor U8346 (N_8346,N_7336,N_6166);
or U8347 (N_8347,N_7425,N_6677);
nand U8348 (N_8348,N_7216,N_7567);
and U8349 (N_8349,N_7041,N_7022);
and U8350 (N_8350,N_7443,N_6949);
or U8351 (N_8351,N_7886,N_7335);
and U8352 (N_8352,N_7064,N_6631);
nor U8353 (N_8353,N_7176,N_6925);
nor U8354 (N_8354,N_7405,N_7136);
and U8355 (N_8355,N_7687,N_6116);
nand U8356 (N_8356,N_6086,N_7815);
xor U8357 (N_8357,N_6994,N_6253);
nor U8358 (N_8358,N_6132,N_7262);
xor U8359 (N_8359,N_6341,N_7440);
nor U8360 (N_8360,N_6418,N_7558);
nand U8361 (N_8361,N_7481,N_7931);
nand U8362 (N_8362,N_7496,N_7517);
and U8363 (N_8363,N_7921,N_7030);
and U8364 (N_8364,N_7878,N_7308);
and U8365 (N_8365,N_7622,N_7914);
and U8366 (N_8366,N_7192,N_7734);
nor U8367 (N_8367,N_7784,N_6096);
or U8368 (N_8368,N_6981,N_6200);
xnor U8369 (N_8369,N_6234,N_7270);
nand U8370 (N_8370,N_6670,N_6019);
or U8371 (N_8371,N_7470,N_6950);
nand U8372 (N_8372,N_7605,N_6501);
nand U8373 (N_8373,N_6555,N_6903);
nand U8374 (N_8374,N_6482,N_7348);
or U8375 (N_8375,N_7149,N_6898);
or U8376 (N_8376,N_7293,N_7305);
nand U8377 (N_8377,N_6470,N_7750);
or U8378 (N_8378,N_6574,N_6427);
or U8379 (N_8379,N_7444,N_6109);
nor U8380 (N_8380,N_6575,N_7673);
nor U8381 (N_8381,N_6783,N_6251);
nand U8382 (N_8382,N_6160,N_7361);
and U8383 (N_8383,N_7680,N_6304);
xor U8384 (N_8384,N_7084,N_7212);
nand U8385 (N_8385,N_7048,N_6381);
nand U8386 (N_8386,N_7994,N_7402);
nor U8387 (N_8387,N_7438,N_7271);
and U8388 (N_8388,N_6938,N_7243);
and U8389 (N_8389,N_6491,N_7333);
nand U8390 (N_8390,N_6629,N_7636);
or U8391 (N_8391,N_6782,N_7382);
nand U8392 (N_8392,N_7712,N_7723);
or U8393 (N_8393,N_6973,N_6584);
and U8394 (N_8394,N_6077,N_7221);
xor U8395 (N_8395,N_6497,N_6827);
or U8396 (N_8396,N_6704,N_7179);
and U8397 (N_8397,N_6630,N_6879);
nor U8398 (N_8398,N_6425,N_6984);
and U8399 (N_8399,N_6171,N_6091);
nor U8400 (N_8400,N_6098,N_7360);
or U8401 (N_8401,N_6442,N_6093);
or U8402 (N_8402,N_6600,N_7074);
nand U8403 (N_8403,N_6335,N_6178);
and U8404 (N_8404,N_6612,N_7415);
nand U8405 (N_8405,N_6458,N_7609);
nand U8406 (N_8406,N_6054,N_7871);
and U8407 (N_8407,N_6307,N_6855);
or U8408 (N_8408,N_6977,N_6492);
xor U8409 (N_8409,N_7901,N_7963);
nor U8410 (N_8410,N_6583,N_6627);
xnor U8411 (N_8411,N_6048,N_6185);
xnor U8412 (N_8412,N_6935,N_7265);
nand U8413 (N_8413,N_6036,N_7231);
nand U8414 (N_8414,N_6009,N_6639);
nor U8415 (N_8415,N_6970,N_7469);
xor U8416 (N_8416,N_6279,N_7716);
or U8417 (N_8417,N_7835,N_6306);
nand U8418 (N_8418,N_7430,N_6360);
nand U8419 (N_8419,N_7384,N_7554);
nand U8420 (N_8420,N_6577,N_7522);
nor U8421 (N_8421,N_7808,N_7512);
nor U8422 (N_8422,N_7121,N_6172);
or U8423 (N_8423,N_7523,N_7061);
and U8424 (N_8424,N_7222,N_7842);
and U8425 (N_8425,N_7834,N_7138);
or U8426 (N_8426,N_7461,N_6193);
or U8427 (N_8427,N_7204,N_6700);
and U8428 (N_8428,N_7819,N_7509);
nand U8429 (N_8429,N_7036,N_7913);
and U8430 (N_8430,N_6352,N_6982);
nor U8431 (N_8431,N_7797,N_6097);
nor U8432 (N_8432,N_7747,N_7690);
and U8433 (N_8433,N_7962,N_7167);
nor U8434 (N_8434,N_7256,N_6849);
xor U8435 (N_8435,N_7320,N_7855);
nor U8436 (N_8436,N_7248,N_7081);
nor U8437 (N_8437,N_7500,N_7803);
nand U8438 (N_8438,N_6573,N_6537);
and U8439 (N_8439,N_7563,N_6597);
nand U8440 (N_8440,N_7583,N_7526);
and U8441 (N_8441,N_6060,N_7058);
nand U8442 (N_8442,N_7363,N_7852);
or U8443 (N_8443,N_7613,N_6342);
xor U8444 (N_8444,N_6305,N_7040);
nor U8445 (N_8445,N_7929,N_7427);
nor U8446 (N_8446,N_6196,N_7957);
or U8447 (N_8447,N_7028,N_7841);
or U8448 (N_8448,N_7515,N_7094);
nand U8449 (N_8449,N_7546,N_7474);
and U8450 (N_8450,N_7621,N_6322);
nand U8451 (N_8451,N_6312,N_7733);
nor U8452 (N_8452,N_6805,N_6736);
and U8453 (N_8453,N_6134,N_6602);
or U8454 (N_8454,N_6955,N_6884);
xor U8455 (N_8455,N_7801,N_7874);
nor U8456 (N_8456,N_7466,N_6962);
xnor U8457 (N_8457,N_7477,N_6095);
nor U8458 (N_8458,N_6591,N_7116);
and U8459 (N_8459,N_6405,N_6763);
or U8460 (N_8460,N_7792,N_6919);
nor U8461 (N_8461,N_7476,N_6883);
nand U8462 (N_8462,N_7218,N_6596);
nor U8463 (N_8463,N_6852,N_7023);
and U8464 (N_8464,N_6592,N_6853);
or U8465 (N_8465,N_6525,N_6027);
and U8466 (N_8466,N_6675,N_6236);
and U8467 (N_8467,N_6106,N_6811);
and U8468 (N_8468,N_7261,N_7426);
nor U8469 (N_8469,N_6548,N_7452);
and U8470 (N_8470,N_7544,N_7740);
and U8471 (N_8471,N_7011,N_6635);
or U8472 (N_8472,N_7379,N_7707);
nor U8473 (N_8473,N_6413,N_7556);
nand U8474 (N_8474,N_7783,N_7387);
or U8475 (N_8475,N_7202,N_6203);
nand U8476 (N_8476,N_7450,N_7302);
or U8477 (N_8477,N_6103,N_7664);
and U8478 (N_8478,N_6162,N_7306);
and U8479 (N_8479,N_6286,N_6968);
nand U8480 (N_8480,N_6915,N_7459);
or U8481 (N_8481,N_7928,N_6625);
or U8482 (N_8482,N_7119,N_7412);
xor U8483 (N_8483,N_7891,N_6452);
or U8484 (N_8484,N_6437,N_7153);
nor U8485 (N_8485,N_6045,N_6706);
nor U8486 (N_8486,N_6720,N_7876);
xnor U8487 (N_8487,N_7009,N_7902);
or U8488 (N_8488,N_7180,N_6433);
and U8489 (N_8489,N_7480,N_6529);
nand U8490 (N_8490,N_7279,N_6871);
or U8491 (N_8491,N_7814,N_7668);
and U8492 (N_8492,N_7285,N_7739);
nor U8493 (N_8493,N_6297,N_7565);
nor U8494 (N_8494,N_6221,N_6033);
nor U8495 (N_8495,N_6288,N_6974);
nor U8496 (N_8496,N_7369,N_7177);
and U8497 (N_8497,N_6387,N_7475);
or U8498 (N_8498,N_7873,N_6485);
and U8499 (N_8499,N_6456,N_6509);
or U8500 (N_8500,N_6204,N_6325);
xnor U8501 (N_8501,N_6189,N_6846);
or U8502 (N_8502,N_7850,N_7840);
nand U8503 (N_8503,N_7887,N_6946);
nand U8504 (N_8504,N_7025,N_6518);
nor U8505 (N_8505,N_6028,N_7705);
nand U8506 (N_8506,N_6490,N_7051);
nor U8507 (N_8507,N_7458,N_6532);
nor U8508 (N_8508,N_7154,N_6594);
or U8509 (N_8509,N_6393,N_7889);
or U8510 (N_8510,N_6317,N_7123);
or U8511 (N_8511,N_6709,N_7370);
nand U8512 (N_8512,N_6085,N_7213);
nand U8513 (N_8513,N_7315,N_7974);
nor U8514 (N_8514,N_7230,N_7832);
nand U8515 (N_8515,N_6310,N_6161);
nor U8516 (N_8516,N_6015,N_7010);
nor U8517 (N_8517,N_6220,N_6000);
and U8518 (N_8518,N_7798,N_7386);
xor U8519 (N_8519,N_6887,N_6951);
xor U8520 (N_8520,N_6117,N_6515);
nor U8521 (N_8521,N_6885,N_7812);
xnor U8522 (N_8522,N_6857,N_7403);
or U8523 (N_8523,N_7557,N_7773);
xor U8524 (N_8524,N_7828,N_7510);
or U8525 (N_8525,N_7236,N_6643);
xnor U8526 (N_8526,N_7727,N_6854);
or U8527 (N_8527,N_7451,N_7158);
nand U8528 (N_8528,N_6375,N_7502);
nor U8529 (N_8529,N_7591,N_6589);
xnor U8530 (N_8530,N_6276,N_7607);
and U8531 (N_8531,N_6453,N_6102);
nand U8532 (N_8532,N_6511,N_7449);
xor U8533 (N_8533,N_6267,N_6713);
and U8534 (N_8534,N_6474,N_7772);
xor U8535 (N_8535,N_7728,N_7503);
and U8536 (N_8536,N_7175,N_6318);
and U8537 (N_8537,N_7757,N_7904);
or U8538 (N_8538,N_6426,N_6072);
nand U8539 (N_8539,N_7972,N_7035);
nor U8540 (N_8540,N_7882,N_7062);
nand U8541 (N_8541,N_6929,N_7059);
nand U8542 (N_8542,N_7206,N_7095);
nand U8543 (N_8543,N_6285,N_7738);
nor U8544 (N_8544,N_7362,N_6327);
nor U8545 (N_8545,N_7436,N_6601);
nand U8546 (N_8546,N_6735,N_6793);
nand U8547 (N_8547,N_6810,N_7845);
xor U8548 (N_8548,N_6859,N_6216);
nand U8549 (N_8549,N_7987,N_6336);
and U8550 (N_8550,N_7985,N_7263);
nor U8551 (N_8551,N_6680,N_7437);
nor U8552 (N_8552,N_6421,N_7042);
nor U8553 (N_8553,N_6513,N_7965);
or U8554 (N_8554,N_6112,N_7371);
nand U8555 (N_8555,N_6804,N_7589);
and U8556 (N_8556,N_7837,N_7999);
nor U8557 (N_8557,N_7092,N_6023);
nand U8558 (N_8558,N_7357,N_7604);
and U8559 (N_8559,N_6489,N_7488);
nand U8560 (N_8560,N_6726,N_7060);
and U8561 (N_8561,N_6108,N_6640);
and U8562 (N_8562,N_6522,N_7034);
nor U8563 (N_8563,N_7165,N_7339);
xor U8564 (N_8564,N_7719,N_6303);
nand U8565 (N_8565,N_7292,N_7781);
or U8566 (N_8566,N_7789,N_6882);
xnor U8567 (N_8567,N_6135,N_6315);
nor U8568 (N_8568,N_6667,N_6826);
and U8569 (N_8569,N_6141,N_7429);
xor U8570 (N_8570,N_6016,N_7731);
nand U8571 (N_8571,N_6765,N_7029);
and U8572 (N_8572,N_7096,N_7065);
nor U8573 (N_8573,N_6789,N_7020);
nor U8574 (N_8574,N_7467,N_7881);
nor U8575 (N_8575,N_6188,N_6966);
nor U8576 (N_8576,N_6207,N_6878);
nand U8577 (N_8577,N_6051,N_6431);
or U8578 (N_8578,N_7755,N_6065);
xnor U8579 (N_8579,N_7529,N_7960);
xnor U8580 (N_8580,N_7434,N_6382);
or U8581 (N_8581,N_6505,N_6448);
or U8582 (N_8582,N_7846,N_6359);
or U8583 (N_8583,N_7967,N_6006);
nor U8584 (N_8584,N_6737,N_6264);
nor U8585 (N_8585,N_6904,N_7907);
or U8586 (N_8586,N_6275,N_6073);
or U8587 (N_8587,N_7000,N_7378);
or U8588 (N_8588,N_7031,N_7768);
or U8589 (N_8589,N_7491,N_7910);
xnor U8590 (N_8590,N_7254,N_6590);
or U8591 (N_8591,N_6223,N_7513);
nor U8592 (N_8592,N_6461,N_7895);
and U8593 (N_8593,N_7943,N_6029);
xnor U8594 (N_8594,N_6550,N_6645);
nand U8595 (N_8595,N_7126,N_7700);
and U8596 (N_8596,N_7581,N_6638);
nor U8597 (N_8597,N_6013,N_6780);
xnor U8598 (N_8598,N_6240,N_6348);
and U8599 (N_8599,N_6653,N_6487);
xnor U8600 (N_8600,N_6295,N_7709);
or U8601 (N_8601,N_6632,N_7582);
and U8602 (N_8602,N_6260,N_6319);
nand U8603 (N_8603,N_6708,N_6683);
and U8604 (N_8604,N_7283,N_6388);
nor U8605 (N_8605,N_7954,N_6986);
nand U8606 (N_8606,N_6554,N_6005);
nand U8607 (N_8607,N_7494,N_7266);
or U8608 (N_8608,N_7670,N_7569);
nand U8609 (N_8609,N_6865,N_7066);
or U8610 (N_8610,N_7104,N_7115);
or U8611 (N_8611,N_7958,N_7805);
nor U8612 (N_8612,N_7486,N_6781);
and U8613 (N_8613,N_7372,N_6198);
or U8614 (N_8614,N_6397,N_6512);
xnor U8615 (N_8615,N_7346,N_7090);
and U8616 (N_8616,N_6834,N_6422);
or U8617 (N_8617,N_6364,N_7763);
nand U8618 (N_8618,N_6170,N_6976);
and U8619 (N_8619,N_7778,N_6436);
nor U8620 (N_8620,N_6140,N_7646);
nand U8621 (N_8621,N_7052,N_7356);
nor U8622 (N_8622,N_6987,N_7368);
xnor U8623 (N_8623,N_6556,N_7319);
nor U8624 (N_8624,N_6353,N_7542);
nor U8625 (N_8625,N_6621,N_6546);
or U8626 (N_8626,N_7304,N_7130);
and U8627 (N_8627,N_7373,N_6389);
nand U8628 (N_8628,N_7950,N_7327);
nor U8629 (N_8629,N_7017,N_7702);
nor U8630 (N_8630,N_7737,N_6872);
nand U8631 (N_8631,N_6347,N_7272);
nor U8632 (N_8632,N_7233,N_7682);
or U8633 (N_8633,N_6183,N_7229);
nand U8634 (N_8634,N_7129,N_7252);
and U8635 (N_8635,N_6916,N_7391);
nand U8636 (N_8636,N_7683,N_7807);
nand U8637 (N_8637,N_6710,N_6227);
xor U8638 (N_8638,N_6008,N_6478);
or U8639 (N_8639,N_7225,N_6877);
or U8640 (N_8640,N_6666,N_6862);
nor U8641 (N_8641,N_7847,N_6531);
nor U8642 (N_8642,N_7490,N_7699);
nand U8643 (N_8643,N_7966,N_6400);
or U8644 (N_8644,N_7005,N_7098);
nand U8645 (N_8645,N_7648,N_7829);
or U8646 (N_8646,N_6745,N_6933);
or U8647 (N_8647,N_7435,N_7631);
nand U8648 (N_8648,N_6776,N_7267);
and U8649 (N_8649,N_7027,N_6114);
nor U8650 (N_8650,N_6595,N_6302);
xor U8651 (N_8651,N_6100,N_7164);
xor U8652 (N_8652,N_7849,N_7932);
xor U8653 (N_8653,N_6101,N_7446);
nand U8654 (N_8654,N_7823,N_6298);
nor U8655 (N_8655,N_6104,N_7050);
and U8656 (N_8656,N_6150,N_6222);
nand U8657 (N_8657,N_6586,N_7939);
or U8658 (N_8658,N_7343,N_6158);
and U8659 (N_8659,N_6164,N_7961);
or U8660 (N_8660,N_6309,N_6742);
xor U8661 (N_8661,N_6773,N_6693);
xnor U8662 (N_8662,N_6539,N_6321);
and U8663 (N_8663,N_6087,N_7776);
or U8664 (N_8664,N_6947,N_7586);
nand U8665 (N_8665,N_7237,N_7144);
nor U8666 (N_8666,N_7432,N_6502);
and U8667 (N_8667,N_7032,N_6187);
nand U8668 (N_8668,N_7419,N_6373);
xnor U8669 (N_8669,N_6772,N_7376);
or U8670 (N_8670,N_7131,N_6058);
or U8671 (N_8671,N_6660,N_7983);
or U8672 (N_8672,N_6078,N_6004);
nand U8673 (N_8673,N_6692,N_7785);
or U8674 (N_8674,N_7002,N_6386);
xor U8675 (N_8675,N_6507,N_7830);
or U8676 (N_8676,N_6744,N_6228);
and U8677 (N_8677,N_6415,N_7615);
xor U8678 (N_8678,N_6544,N_6273);
xor U8679 (N_8679,N_6724,N_7075);
and U8680 (N_8680,N_6040,N_7043);
nor U8681 (N_8681,N_7166,N_6126);
nor U8682 (N_8682,N_7013,N_6089);
xnor U8683 (N_8683,N_7984,N_6069);
nand U8684 (N_8684,N_6424,N_7300);
xnor U8685 (N_8685,N_6615,N_7959);
nor U8686 (N_8686,N_7239,N_7482);
nand U8687 (N_8687,N_6891,N_7853);
nand U8688 (N_8688,N_7307,N_7780);
nor U8689 (N_8689,N_7107,N_7637);
and U8690 (N_8690,N_6822,N_6254);
nand U8691 (N_8691,N_6668,N_7316);
or U8692 (N_8692,N_7309,N_7264);
nand U8693 (N_8693,N_7826,N_6616);
and U8694 (N_8694,N_6443,N_7349);
xor U8695 (N_8695,N_7277,N_7501);
nand U8696 (N_8696,N_7506,N_7473);
or U8697 (N_8697,N_7861,N_6463);
and U8698 (N_8698,N_6760,N_7575);
and U8699 (N_8699,N_7108,N_6046);
nand U8700 (N_8700,N_6181,N_6384);
nor U8701 (N_8701,N_6628,N_6289);
nor U8702 (N_8702,N_7752,N_6330);
nor U8703 (N_8703,N_6075,N_7578);
nor U8704 (N_8704,N_6828,N_6292);
nand U8705 (N_8705,N_7455,N_6873);
or U8706 (N_8706,N_6618,N_7822);
and U8707 (N_8707,N_7626,N_6557);
or U8708 (N_8708,N_7598,N_7100);
nand U8709 (N_8709,N_6603,N_6248);
xor U8710 (N_8710,N_7240,N_7174);
nor U8711 (N_8711,N_6767,N_7793);
xor U8712 (N_8712,N_7971,N_6961);
xor U8713 (N_8713,N_6007,N_7162);
nor U8714 (N_8714,N_6167,N_6149);
nand U8715 (N_8715,N_7602,N_6296);
and U8716 (N_8716,N_7620,N_6552);
nand U8717 (N_8717,N_6206,N_6527);
nand U8718 (N_8718,N_7885,N_6136);
or U8719 (N_8719,N_6520,N_6998);
and U8720 (N_8720,N_7207,N_7366);
or U8721 (N_8721,N_6062,N_6191);
and U8722 (N_8722,N_7571,N_7788);
xor U8723 (N_8723,N_7681,N_6848);
nor U8724 (N_8724,N_7381,N_6671);
nor U8725 (N_8725,N_6657,N_6174);
or U8726 (N_8726,N_7298,N_6125);
and U8727 (N_8727,N_6748,N_6052);
xor U8728 (N_8728,N_6498,N_7442);
or U8729 (N_8729,N_6897,N_7762);
and U8730 (N_8730,N_6868,N_7585);
nand U8731 (N_8731,N_6120,N_7203);
nor U8732 (N_8732,N_7843,N_6547);
nand U8733 (N_8733,N_7342,N_6208);
nand U8734 (N_8734,N_6237,N_7611);
or U8735 (N_8735,N_6542,N_7970);
nor U8736 (N_8736,N_6626,N_7888);
nor U8737 (N_8737,N_6311,N_7008);
nand U8738 (N_8738,N_7860,N_6747);
nand U8739 (N_8739,N_6423,N_6696);
or U8740 (N_8740,N_6909,N_7590);
nor U8741 (N_8741,N_7208,N_7978);
nand U8742 (N_8742,N_6281,N_7520);
or U8743 (N_8743,N_7713,N_6331);
or U8744 (N_8744,N_6258,N_7053);
or U8745 (N_8745,N_6980,N_6825);
xor U8746 (N_8746,N_7398,N_6012);
nand U8747 (N_8747,N_7599,N_6730);
or U8748 (N_8748,N_6889,N_6528);
nand U8749 (N_8749,N_7995,N_6622);
or U8750 (N_8750,N_7735,N_7071);
or U8751 (N_8751,N_6122,N_7087);
and U8752 (N_8752,N_7890,N_7189);
xnor U8753 (N_8753,N_6993,N_7205);
or U8754 (N_8754,N_6468,N_6123);
nand U8755 (N_8755,N_7992,N_6948);
nor U8756 (N_8756,N_7867,N_7820);
nand U8757 (N_8757,N_6090,N_7054);
nand U8758 (N_8758,N_6361,N_6684);
nor U8759 (N_8759,N_6992,N_7191);
nand U8760 (N_8760,N_7318,N_7782);
nand U8761 (N_8761,N_6508,N_6368);
nand U8762 (N_8762,N_6369,N_6540);
and U8763 (N_8763,N_7650,N_7485);
nand U8764 (N_8764,N_7870,N_7649);
nor U8765 (N_8765,N_6169,N_7534);
xnor U8766 (N_8766,N_6444,N_6939);
xor U8767 (N_8767,N_7137,N_7388);
xor U8768 (N_8768,N_6988,N_7765);
nand U8769 (N_8769,N_6633,N_7695);
xnor U8770 (N_8770,N_6088,N_7408);
or U8771 (N_8771,N_6519,N_6274);
nand U8772 (N_8772,N_6954,N_6769);
or U8773 (N_8773,N_7741,N_7326);
or U8774 (N_8774,N_6609,N_7080);
or U8775 (N_8775,N_7251,N_6646);
and U8776 (N_8776,N_6179,N_7906);
xor U8777 (N_8777,N_7185,N_6044);
nor U8778 (N_8778,N_6564,N_6447);
nor U8779 (N_8779,N_7616,N_6494);
nand U8780 (N_8780,N_6201,N_6459);
or U8781 (N_8781,N_6960,N_7479);
and U8782 (N_8782,N_6346,N_6503);
nand U8783 (N_8783,N_7717,N_7592);
nand U8784 (N_8784,N_6163,N_7883);
or U8785 (N_8785,N_6063,N_7764);
or U8786 (N_8786,N_7063,N_7478);
nand U8787 (N_8787,N_6071,N_6357);
or U8788 (N_8788,N_7647,N_6280);
nor U8789 (N_8789,N_7644,N_7802);
xnor U8790 (N_8790,N_7933,N_6790);
and U8791 (N_8791,N_6035,N_6758);
nor U8792 (N_8792,N_7937,N_7973);
and U8793 (N_8793,N_7993,N_6642);
or U8794 (N_8794,N_7940,N_7468);
nor U8795 (N_8795,N_6813,N_7210);
or U8796 (N_8796,N_6380,N_7817);
and U8797 (N_8797,N_7685,N_7530);
xor U8798 (N_8798,N_7170,N_6241);
xnor U8799 (N_8799,N_7825,N_7151);
xnor U8800 (N_8800,N_6768,N_7303);
and U8801 (N_8801,N_7539,N_7224);
xnor U8802 (N_8802,N_6299,N_7439);
xor U8803 (N_8803,N_6814,N_6975);
xnor U8804 (N_8804,N_6614,N_7760);
or U8805 (N_8805,N_7535,N_6691);
and U8806 (N_8806,N_6658,N_7483);
xnor U8807 (N_8807,N_7744,N_7746);
and U8808 (N_8808,N_7078,N_7896);
xor U8809 (N_8809,N_7399,N_6472);
nor U8810 (N_8810,N_7021,N_7250);
or U8811 (N_8811,N_6092,N_7511);
xor U8812 (N_8812,N_6190,N_7039);
nor U8813 (N_8813,N_6843,N_7353);
nor U8814 (N_8814,N_7652,N_7492);
and U8815 (N_8815,N_7332,N_7197);
nand U8816 (N_8816,N_6727,N_6579);
or U8817 (N_8817,N_6476,N_6766);
nor U8818 (N_8818,N_6020,N_6032);
xor U8819 (N_8819,N_7686,N_6740);
nor U8820 (N_8820,N_7555,N_6265);
and U8821 (N_8821,N_7724,N_6778);
or U8822 (N_8822,N_6920,N_7748);
xnor U8823 (N_8823,N_6701,N_7464);
nor U8824 (N_8824,N_7273,N_7674);
xnor U8825 (N_8825,N_7194,N_7324);
nand U8826 (N_8826,N_6417,N_6585);
or U8827 (N_8827,N_6676,N_7209);
and U8828 (N_8828,N_7354,N_7396);
nand U8829 (N_8829,N_7574,N_7619);
or U8830 (N_8830,N_7281,N_7289);
nor U8831 (N_8831,N_7227,N_6924);
and U8832 (N_8832,N_7934,N_6937);
nand U8833 (N_8833,N_7079,N_7678);
and U8834 (N_8834,N_6301,N_6647);
nand U8835 (N_8835,N_6669,N_7097);
nor U8836 (N_8836,N_7038,N_7877);
nand U8837 (N_8837,N_6560,N_7157);
or U8838 (N_8838,N_6138,N_6197);
xor U8839 (N_8839,N_7635,N_7920);
nor U8840 (N_8840,N_7456,N_7234);
and U8841 (N_8841,N_6392,N_7337);
and U8842 (N_8842,N_7951,N_6866);
nor U8843 (N_8843,N_7219,N_7527);
nor U8844 (N_8844,N_7791,N_6678);
or U8845 (N_8845,N_7215,N_7200);
nand U8846 (N_8846,N_6759,N_7665);
nand U8847 (N_8847,N_6928,N_7787);
or U8848 (N_8848,N_7809,N_6703);
xnor U8849 (N_8849,N_7161,N_6332);
nor U8850 (N_8850,N_7532,N_7796);
xor U8851 (N_8851,N_7082,N_6762);
nand U8852 (N_8852,N_7068,N_7409);
and U8853 (N_8853,N_6041,N_6687);
and U8854 (N_8854,N_7964,N_6722);
nor U8855 (N_8855,N_6876,N_7758);
nor U8856 (N_8856,N_6002,N_7790);
nand U8857 (N_8857,N_7813,N_6449);
nor U8858 (N_8858,N_7634,N_7956);
xnor U8859 (N_8859,N_7195,N_7540);
xor U8860 (N_8860,N_6366,N_6438);
or U8861 (N_8861,N_7625,N_6083);
and U8862 (N_8862,N_6344,N_7821);
and U8863 (N_8863,N_7697,N_7182);
xor U8864 (N_8864,N_7981,N_6832);
xnor U8865 (N_8865,N_7244,N_7406);
nand U8866 (N_8866,N_6362,N_7922);
and U8867 (N_8867,N_6940,N_6580);
and U8868 (N_8868,N_7253,N_6761);
or U8869 (N_8869,N_7487,N_7718);
nand U8870 (N_8870,N_7377,N_6516);
nor U8871 (N_8871,N_6465,N_7851);
xnor U8872 (N_8872,N_6559,N_6379);
xor U8873 (N_8873,N_6784,N_6607);
and U8874 (N_8874,N_6495,N_6536);
xor U8875 (N_8875,N_7767,N_7325);
xnor U8876 (N_8876,N_6823,N_7863);
nand U8877 (N_8877,N_6829,N_7573);
nor U8878 (N_8878,N_7766,N_7936);
and U8879 (N_8879,N_7411,N_7838);
or U8880 (N_8880,N_7714,N_6791);
xnor U8881 (N_8881,N_6430,N_7926);
nor U8882 (N_8882,N_6578,N_6561);
and U8883 (N_8883,N_7507,N_7334);
nand U8884 (N_8884,N_7380,N_7338);
and U8885 (N_8885,N_6558,N_6953);
or U8886 (N_8886,N_6395,N_7114);
nand U8887 (N_8887,N_7416,N_6681);
or U8888 (N_8888,N_7453,N_6226);
or U8889 (N_8889,N_6563,N_7147);
xor U8890 (N_8890,N_6641,N_7190);
nor U8891 (N_8891,N_6697,N_7653);
or U8892 (N_8892,N_6153,N_6918);
xor U8893 (N_8893,N_6182,N_7317);
nand U8894 (N_8894,N_6441,N_7742);
nand U8895 (N_8895,N_6774,N_6154);
and U8896 (N_8896,N_7560,N_7278);
and U8897 (N_8897,N_6888,N_6329);
nor U8898 (N_8898,N_6892,N_6881);
nand U8899 (N_8899,N_6313,N_7580);
nand U8900 (N_8900,N_7178,N_7761);
nor U8901 (N_8901,N_6858,N_6967);
or U8902 (N_8902,N_6943,N_6408);
and U8903 (N_8903,N_6867,N_7055);
nand U8904 (N_8904,N_6176,N_7774);
or U8905 (N_8905,N_6983,N_6743);
nand U8906 (N_8906,N_6800,N_7101);
and U8907 (N_8907,N_6856,N_7173);
nor U8908 (N_8908,N_6420,N_6157);
and U8909 (N_8909,N_7844,N_6247);
nor U8910 (N_8910,N_6874,N_6712);
nand U8911 (N_8911,N_6475,N_6195);
or U8912 (N_8912,N_7274,N_6541);
or U8913 (N_8913,N_7404,N_7489);
and U8914 (N_8914,N_6517,N_7006);
and U8915 (N_8915,N_6999,N_6151);
xor U8916 (N_8916,N_7284,N_6326);
nor U8917 (N_8917,N_6818,N_7433);
xor U8918 (N_8918,N_7710,N_6934);
and U8919 (N_8919,N_7900,N_6551);
nor U8920 (N_8920,N_7541,N_7694);
and U8921 (N_8921,N_7145,N_6798);
or U8922 (N_8922,N_6145,N_6598);
nand U8923 (N_8923,N_7045,N_6611);
xnor U8924 (N_8924,N_7924,N_7618);
nand U8925 (N_8925,N_7247,N_7942);
nor U8926 (N_8926,N_6410,N_7894);
or U8927 (N_8927,N_6047,N_7692);
nand U8928 (N_8928,N_6707,N_7105);
or U8929 (N_8929,N_7484,N_7321);
and U8930 (N_8930,N_7505,N_6506);
xor U8931 (N_8931,N_6880,N_6113);
nor U8932 (N_8932,N_7726,N_6620);
xor U8933 (N_8933,N_7858,N_7401);
and U8934 (N_8934,N_7099,N_7128);
and U8935 (N_8935,N_6997,N_6269);
nor U8936 (N_8936,N_6695,N_7288);
nand U8937 (N_8937,N_7140,N_7102);
and U8938 (N_8938,N_6808,N_6272);
or U8939 (N_8939,N_7868,N_6412);
nand U8940 (N_8940,N_7898,N_6076);
nand U8941 (N_8941,N_6011,N_7862);
or U8942 (N_8942,N_6419,N_6679);
and U8943 (N_8943,N_7579,N_6530);
nand U8944 (N_8944,N_7968,N_7390);
and U8945 (N_8945,N_7982,N_6039);
nand U8946 (N_8946,N_6608,N_6599);
or U8947 (N_8947,N_6757,N_7662);
nor U8948 (N_8948,N_6213,N_6467);
nand U8949 (N_8949,N_7640,N_7725);
and U8950 (N_8950,N_7462,N_6471);
or U8951 (N_8951,N_7753,N_7344);
and U8952 (N_8952,N_6770,N_7917);
xor U8953 (N_8953,N_6644,N_6752);
and U8954 (N_8954,N_6082,N_6394);
xnor U8955 (N_8955,N_6755,N_7069);
nor U8956 (N_8956,N_7016,N_7143);
nor U8957 (N_8957,N_6777,N_6610);
xor U8958 (N_8958,N_7553,N_6356);
nor U8959 (N_8959,N_6064,N_6455);
nand U8960 (N_8960,N_6290,N_7566);
or U8961 (N_8961,N_6291,N_7927);
or U8962 (N_8962,N_6334,N_6194);
nor U8963 (N_8963,N_7516,N_6232);
xor U8964 (N_8964,N_7947,N_6205);
nand U8965 (N_8965,N_7365,N_7944);
nand U8966 (N_8966,N_6165,N_7001);
xor U8967 (N_8967,N_6902,N_6654);
and U8968 (N_8968,N_7628,N_6079);
and U8969 (N_8969,N_6795,N_7977);
nor U8970 (N_8970,N_6845,N_7330);
nand U8971 (N_8971,N_7800,N_6901);
nor U8972 (N_8972,N_7156,N_6779);
or U8973 (N_8973,N_7806,N_6401);
or U8974 (N_8974,N_6358,N_6371);
or U8975 (N_8975,N_7875,N_7576);
nor U8976 (N_8976,N_7701,N_6690);
nand U8977 (N_8977,N_7915,N_7159);
and U8978 (N_8978,N_7117,N_6337);
nand U8979 (N_8979,N_7314,N_6137);
or U8980 (N_8980,N_7689,N_6649);
nand U8981 (N_8981,N_7341,N_6245);
nor U8982 (N_8982,N_7110,N_7912);
and U8983 (N_8983,N_7299,N_6235);
nor U8984 (N_8984,N_6689,N_7633);
or U8985 (N_8985,N_7015,N_7258);
or U8986 (N_8986,N_6262,N_6905);
and U8987 (N_8987,N_7033,N_6224);
and U8988 (N_8988,N_7996,N_7756);
nor U8989 (N_8989,N_7188,N_6080);
and U8990 (N_8990,N_7606,N_7880);
or U8991 (N_8991,N_6484,N_6582);
nor U8992 (N_8992,N_6021,N_7465);
xor U8993 (N_8993,N_6533,N_6569);
nor U8994 (N_8994,N_7769,N_6535);
nor U8995 (N_8995,N_6259,N_7007);
xor U8996 (N_8996,N_6300,N_6593);
nor U8997 (N_8997,N_6672,N_7414);
nand U8998 (N_8998,N_6797,N_6753);
xor U8999 (N_8999,N_7454,N_6604);
nand U9000 (N_9000,N_6831,N_7773);
or U9001 (N_9001,N_6406,N_7818);
or U9002 (N_9002,N_6168,N_7983);
nor U9003 (N_9003,N_6163,N_6544);
nand U9004 (N_9004,N_7134,N_7891);
or U9005 (N_9005,N_7304,N_6735);
xor U9006 (N_9006,N_7752,N_6693);
and U9007 (N_9007,N_6535,N_6683);
or U9008 (N_9008,N_7657,N_7424);
nor U9009 (N_9009,N_6780,N_7581);
xnor U9010 (N_9010,N_7063,N_6767);
and U9011 (N_9011,N_6461,N_7744);
nand U9012 (N_9012,N_6550,N_6068);
nand U9013 (N_9013,N_7853,N_6878);
xor U9014 (N_9014,N_6048,N_7210);
nor U9015 (N_9015,N_6777,N_6505);
and U9016 (N_9016,N_7208,N_7901);
xnor U9017 (N_9017,N_7565,N_7991);
nor U9018 (N_9018,N_7775,N_7830);
and U9019 (N_9019,N_7928,N_7274);
xnor U9020 (N_9020,N_7510,N_7839);
or U9021 (N_9021,N_7081,N_6529);
or U9022 (N_9022,N_6262,N_6692);
xnor U9023 (N_9023,N_6784,N_7927);
nor U9024 (N_9024,N_6795,N_6192);
xor U9025 (N_9025,N_6858,N_7386);
or U9026 (N_9026,N_7366,N_7372);
xor U9027 (N_9027,N_6037,N_7141);
xnor U9028 (N_9028,N_7967,N_7609);
xor U9029 (N_9029,N_6069,N_7298);
xnor U9030 (N_9030,N_6491,N_6233);
nand U9031 (N_9031,N_6879,N_6727);
and U9032 (N_9032,N_6297,N_6412);
and U9033 (N_9033,N_7701,N_7853);
xor U9034 (N_9034,N_6644,N_7544);
xnor U9035 (N_9035,N_6053,N_7887);
xor U9036 (N_9036,N_7692,N_7777);
nand U9037 (N_9037,N_6839,N_6501);
nor U9038 (N_9038,N_6047,N_6737);
and U9039 (N_9039,N_7519,N_6751);
and U9040 (N_9040,N_7724,N_6999);
nand U9041 (N_9041,N_7992,N_6724);
and U9042 (N_9042,N_6190,N_6949);
nand U9043 (N_9043,N_6802,N_6747);
nand U9044 (N_9044,N_6466,N_6724);
nor U9045 (N_9045,N_6182,N_7681);
xnor U9046 (N_9046,N_7923,N_6054);
nand U9047 (N_9047,N_6038,N_7166);
and U9048 (N_9048,N_7843,N_6733);
nand U9049 (N_9049,N_6479,N_7227);
nor U9050 (N_9050,N_7594,N_7969);
nand U9051 (N_9051,N_6113,N_6226);
and U9052 (N_9052,N_6219,N_7900);
nand U9053 (N_9053,N_6785,N_7117);
nor U9054 (N_9054,N_7697,N_6375);
or U9055 (N_9055,N_6175,N_7516);
or U9056 (N_9056,N_6151,N_6225);
nor U9057 (N_9057,N_6143,N_6982);
or U9058 (N_9058,N_6566,N_6111);
xnor U9059 (N_9059,N_6288,N_6302);
xor U9060 (N_9060,N_6676,N_7220);
xor U9061 (N_9061,N_7239,N_7714);
nand U9062 (N_9062,N_7577,N_6840);
and U9063 (N_9063,N_7061,N_6342);
or U9064 (N_9064,N_6305,N_6150);
and U9065 (N_9065,N_6158,N_6788);
and U9066 (N_9066,N_7799,N_6086);
nand U9067 (N_9067,N_6670,N_6949);
nor U9068 (N_9068,N_6486,N_6423);
or U9069 (N_9069,N_7017,N_7569);
and U9070 (N_9070,N_7484,N_6542);
nor U9071 (N_9071,N_6647,N_7231);
xnor U9072 (N_9072,N_7571,N_6915);
nand U9073 (N_9073,N_7808,N_6682);
nor U9074 (N_9074,N_7593,N_6003);
and U9075 (N_9075,N_6374,N_7481);
and U9076 (N_9076,N_6402,N_6337);
or U9077 (N_9077,N_7498,N_6280);
nand U9078 (N_9078,N_7196,N_7124);
and U9079 (N_9079,N_7473,N_6511);
or U9080 (N_9080,N_6596,N_7292);
and U9081 (N_9081,N_6327,N_6317);
nand U9082 (N_9082,N_6751,N_6408);
nor U9083 (N_9083,N_7396,N_7550);
xnor U9084 (N_9084,N_7495,N_6885);
and U9085 (N_9085,N_7565,N_7833);
nor U9086 (N_9086,N_7068,N_6161);
nand U9087 (N_9087,N_6949,N_7123);
nor U9088 (N_9088,N_7952,N_6429);
and U9089 (N_9089,N_6237,N_6016);
nor U9090 (N_9090,N_6800,N_6460);
and U9091 (N_9091,N_7338,N_7033);
or U9092 (N_9092,N_6739,N_7070);
nand U9093 (N_9093,N_7097,N_6690);
nand U9094 (N_9094,N_6928,N_7565);
nand U9095 (N_9095,N_6264,N_7398);
nand U9096 (N_9096,N_6920,N_7412);
or U9097 (N_9097,N_7086,N_7134);
and U9098 (N_9098,N_7483,N_6416);
nor U9099 (N_9099,N_7757,N_6699);
xor U9100 (N_9100,N_7839,N_6766);
or U9101 (N_9101,N_6465,N_7554);
xor U9102 (N_9102,N_7590,N_7965);
or U9103 (N_9103,N_7771,N_7635);
nand U9104 (N_9104,N_6373,N_7210);
and U9105 (N_9105,N_7253,N_7689);
nand U9106 (N_9106,N_7846,N_7608);
or U9107 (N_9107,N_6597,N_6162);
or U9108 (N_9108,N_7277,N_7366);
and U9109 (N_9109,N_7485,N_6432);
and U9110 (N_9110,N_7453,N_6820);
or U9111 (N_9111,N_6388,N_6400);
or U9112 (N_9112,N_7334,N_7998);
or U9113 (N_9113,N_6142,N_6112);
or U9114 (N_9114,N_7062,N_7106);
xor U9115 (N_9115,N_7117,N_6651);
and U9116 (N_9116,N_6224,N_6186);
nand U9117 (N_9117,N_7274,N_7368);
and U9118 (N_9118,N_7710,N_6342);
or U9119 (N_9119,N_7845,N_7096);
or U9120 (N_9120,N_7220,N_7345);
nand U9121 (N_9121,N_6586,N_7254);
and U9122 (N_9122,N_6053,N_6854);
nor U9123 (N_9123,N_6375,N_7317);
nand U9124 (N_9124,N_7116,N_7105);
and U9125 (N_9125,N_6436,N_7740);
nor U9126 (N_9126,N_6531,N_6082);
or U9127 (N_9127,N_6485,N_6418);
or U9128 (N_9128,N_6728,N_7045);
or U9129 (N_9129,N_6355,N_7385);
and U9130 (N_9130,N_7424,N_7000);
or U9131 (N_9131,N_7826,N_6218);
or U9132 (N_9132,N_7096,N_6320);
and U9133 (N_9133,N_7450,N_7618);
or U9134 (N_9134,N_7398,N_6342);
or U9135 (N_9135,N_7801,N_7838);
or U9136 (N_9136,N_6239,N_6218);
and U9137 (N_9137,N_7883,N_7712);
nand U9138 (N_9138,N_6146,N_7564);
nor U9139 (N_9139,N_7167,N_7601);
and U9140 (N_9140,N_6420,N_7393);
xnor U9141 (N_9141,N_7318,N_7401);
or U9142 (N_9142,N_7224,N_7748);
nand U9143 (N_9143,N_7541,N_7307);
and U9144 (N_9144,N_7891,N_6968);
nand U9145 (N_9145,N_6663,N_6902);
nand U9146 (N_9146,N_6630,N_7906);
xnor U9147 (N_9147,N_7912,N_6672);
nor U9148 (N_9148,N_7920,N_6833);
and U9149 (N_9149,N_6551,N_7920);
nor U9150 (N_9150,N_6175,N_6298);
nand U9151 (N_9151,N_7672,N_7244);
nand U9152 (N_9152,N_6496,N_6111);
or U9153 (N_9153,N_6328,N_7082);
nand U9154 (N_9154,N_7041,N_6319);
nand U9155 (N_9155,N_6180,N_7694);
nand U9156 (N_9156,N_6778,N_6034);
and U9157 (N_9157,N_6205,N_6252);
xor U9158 (N_9158,N_7235,N_7779);
xnor U9159 (N_9159,N_6632,N_7938);
xnor U9160 (N_9160,N_7975,N_6583);
and U9161 (N_9161,N_6495,N_7676);
and U9162 (N_9162,N_6255,N_7822);
and U9163 (N_9163,N_7688,N_7821);
xor U9164 (N_9164,N_6141,N_7547);
xor U9165 (N_9165,N_7548,N_6146);
and U9166 (N_9166,N_7403,N_6841);
or U9167 (N_9167,N_6395,N_6471);
nand U9168 (N_9168,N_7877,N_6537);
nand U9169 (N_9169,N_6870,N_6611);
nor U9170 (N_9170,N_6741,N_6112);
and U9171 (N_9171,N_6848,N_6099);
and U9172 (N_9172,N_7653,N_7727);
or U9173 (N_9173,N_6606,N_7145);
nand U9174 (N_9174,N_7149,N_6382);
xnor U9175 (N_9175,N_7474,N_6813);
xor U9176 (N_9176,N_7094,N_7540);
or U9177 (N_9177,N_7445,N_6280);
xnor U9178 (N_9178,N_6364,N_6053);
nor U9179 (N_9179,N_7239,N_7522);
nand U9180 (N_9180,N_6590,N_7192);
nor U9181 (N_9181,N_7323,N_6479);
nor U9182 (N_9182,N_6998,N_6786);
xor U9183 (N_9183,N_6709,N_6017);
xnor U9184 (N_9184,N_6024,N_6337);
nand U9185 (N_9185,N_6766,N_7708);
nor U9186 (N_9186,N_6440,N_6058);
nor U9187 (N_9187,N_6555,N_7373);
nand U9188 (N_9188,N_6857,N_6864);
and U9189 (N_9189,N_7378,N_6972);
and U9190 (N_9190,N_6854,N_6513);
and U9191 (N_9191,N_7502,N_6487);
nor U9192 (N_9192,N_7384,N_7545);
nand U9193 (N_9193,N_6888,N_6462);
nand U9194 (N_9194,N_6998,N_6546);
xnor U9195 (N_9195,N_7691,N_6652);
or U9196 (N_9196,N_7512,N_6443);
or U9197 (N_9197,N_6309,N_7312);
or U9198 (N_9198,N_6774,N_6779);
nand U9199 (N_9199,N_6117,N_6607);
or U9200 (N_9200,N_7779,N_6863);
nand U9201 (N_9201,N_6916,N_6506);
xnor U9202 (N_9202,N_6464,N_6732);
and U9203 (N_9203,N_7241,N_7605);
xnor U9204 (N_9204,N_7302,N_6693);
xor U9205 (N_9205,N_7887,N_6276);
nand U9206 (N_9206,N_7060,N_7899);
or U9207 (N_9207,N_7294,N_7035);
and U9208 (N_9208,N_7870,N_7767);
xor U9209 (N_9209,N_7192,N_6703);
or U9210 (N_9210,N_7500,N_7633);
or U9211 (N_9211,N_7189,N_6252);
xnor U9212 (N_9212,N_7194,N_7407);
nor U9213 (N_9213,N_6179,N_7855);
and U9214 (N_9214,N_6743,N_6924);
and U9215 (N_9215,N_6108,N_6212);
nand U9216 (N_9216,N_6816,N_7996);
nand U9217 (N_9217,N_7613,N_6071);
nor U9218 (N_9218,N_6207,N_6048);
and U9219 (N_9219,N_6018,N_7901);
or U9220 (N_9220,N_7107,N_7523);
and U9221 (N_9221,N_6892,N_7773);
or U9222 (N_9222,N_7119,N_6916);
and U9223 (N_9223,N_6785,N_7646);
xnor U9224 (N_9224,N_6002,N_7710);
and U9225 (N_9225,N_7491,N_7954);
nor U9226 (N_9226,N_6117,N_7384);
nor U9227 (N_9227,N_6738,N_7868);
nor U9228 (N_9228,N_7449,N_7854);
xnor U9229 (N_9229,N_7693,N_7989);
xnor U9230 (N_9230,N_6116,N_7997);
nor U9231 (N_9231,N_7508,N_6399);
or U9232 (N_9232,N_6255,N_6729);
and U9233 (N_9233,N_7286,N_6459);
or U9234 (N_9234,N_7506,N_7874);
or U9235 (N_9235,N_7297,N_7446);
xor U9236 (N_9236,N_6441,N_6000);
xor U9237 (N_9237,N_6101,N_6357);
or U9238 (N_9238,N_6630,N_6949);
and U9239 (N_9239,N_6660,N_7446);
nor U9240 (N_9240,N_7642,N_6726);
or U9241 (N_9241,N_6022,N_7210);
and U9242 (N_9242,N_6594,N_7997);
nor U9243 (N_9243,N_7668,N_7633);
and U9244 (N_9244,N_6409,N_7741);
xor U9245 (N_9245,N_7508,N_7743);
nor U9246 (N_9246,N_7672,N_7980);
nor U9247 (N_9247,N_6915,N_6280);
nand U9248 (N_9248,N_7293,N_6627);
or U9249 (N_9249,N_6463,N_7215);
or U9250 (N_9250,N_7242,N_7214);
nor U9251 (N_9251,N_6923,N_7959);
nor U9252 (N_9252,N_7790,N_6350);
and U9253 (N_9253,N_7844,N_6410);
xor U9254 (N_9254,N_7596,N_6567);
nor U9255 (N_9255,N_7356,N_7120);
and U9256 (N_9256,N_6883,N_6184);
nor U9257 (N_9257,N_6079,N_6918);
xnor U9258 (N_9258,N_7057,N_6167);
nand U9259 (N_9259,N_6933,N_7037);
nor U9260 (N_9260,N_6140,N_7054);
or U9261 (N_9261,N_7250,N_7094);
and U9262 (N_9262,N_6651,N_7279);
xnor U9263 (N_9263,N_7400,N_7824);
xnor U9264 (N_9264,N_7199,N_7309);
xnor U9265 (N_9265,N_7626,N_6445);
nand U9266 (N_9266,N_7913,N_7193);
xor U9267 (N_9267,N_7081,N_7595);
nand U9268 (N_9268,N_7982,N_6507);
xnor U9269 (N_9269,N_7817,N_6594);
or U9270 (N_9270,N_6495,N_6981);
nand U9271 (N_9271,N_7579,N_6989);
nor U9272 (N_9272,N_7593,N_6250);
or U9273 (N_9273,N_6406,N_7726);
nor U9274 (N_9274,N_6181,N_7241);
xnor U9275 (N_9275,N_7979,N_6469);
nand U9276 (N_9276,N_6340,N_7703);
xor U9277 (N_9277,N_7186,N_6432);
or U9278 (N_9278,N_7473,N_6525);
nand U9279 (N_9279,N_6944,N_6804);
nand U9280 (N_9280,N_7487,N_7126);
nand U9281 (N_9281,N_7524,N_7487);
nor U9282 (N_9282,N_7767,N_6280);
nand U9283 (N_9283,N_6367,N_7278);
xor U9284 (N_9284,N_7305,N_6879);
nor U9285 (N_9285,N_7394,N_6638);
xor U9286 (N_9286,N_7304,N_6506);
nand U9287 (N_9287,N_7948,N_7465);
nor U9288 (N_9288,N_6069,N_6690);
nor U9289 (N_9289,N_7345,N_7957);
and U9290 (N_9290,N_6100,N_7491);
or U9291 (N_9291,N_7869,N_6270);
or U9292 (N_9292,N_6452,N_7203);
xnor U9293 (N_9293,N_7602,N_7908);
xor U9294 (N_9294,N_7032,N_6078);
xnor U9295 (N_9295,N_6942,N_7778);
nand U9296 (N_9296,N_6271,N_7667);
nand U9297 (N_9297,N_7613,N_6648);
or U9298 (N_9298,N_7424,N_7114);
or U9299 (N_9299,N_6574,N_6382);
nand U9300 (N_9300,N_6135,N_7478);
and U9301 (N_9301,N_7834,N_7265);
nor U9302 (N_9302,N_6709,N_6629);
nor U9303 (N_9303,N_7208,N_7522);
nand U9304 (N_9304,N_7007,N_6736);
or U9305 (N_9305,N_6002,N_7682);
nand U9306 (N_9306,N_6835,N_6748);
nor U9307 (N_9307,N_7686,N_7509);
nor U9308 (N_9308,N_6394,N_6465);
nor U9309 (N_9309,N_6219,N_7301);
xor U9310 (N_9310,N_7491,N_6235);
and U9311 (N_9311,N_6137,N_6473);
nor U9312 (N_9312,N_6257,N_7141);
nand U9313 (N_9313,N_6767,N_6805);
nand U9314 (N_9314,N_7033,N_7852);
nor U9315 (N_9315,N_6891,N_6292);
nor U9316 (N_9316,N_6445,N_7268);
xnor U9317 (N_9317,N_6909,N_7192);
nand U9318 (N_9318,N_6566,N_7294);
and U9319 (N_9319,N_6888,N_7160);
xnor U9320 (N_9320,N_6385,N_6451);
xnor U9321 (N_9321,N_7485,N_6893);
nand U9322 (N_9322,N_6395,N_6469);
nand U9323 (N_9323,N_7692,N_7917);
or U9324 (N_9324,N_7049,N_6308);
and U9325 (N_9325,N_7835,N_7453);
nand U9326 (N_9326,N_6068,N_7756);
or U9327 (N_9327,N_7734,N_6572);
and U9328 (N_9328,N_7755,N_6501);
and U9329 (N_9329,N_7705,N_7191);
nand U9330 (N_9330,N_7961,N_6700);
xor U9331 (N_9331,N_7511,N_6082);
nand U9332 (N_9332,N_6923,N_6284);
nor U9333 (N_9333,N_7061,N_7283);
nand U9334 (N_9334,N_7042,N_6976);
and U9335 (N_9335,N_6348,N_6409);
or U9336 (N_9336,N_7918,N_6693);
nor U9337 (N_9337,N_6939,N_6329);
or U9338 (N_9338,N_6072,N_7513);
xnor U9339 (N_9339,N_7616,N_6531);
nor U9340 (N_9340,N_7303,N_6733);
nor U9341 (N_9341,N_7003,N_6210);
nor U9342 (N_9342,N_7851,N_7107);
xnor U9343 (N_9343,N_6395,N_7946);
nor U9344 (N_9344,N_6262,N_7552);
nand U9345 (N_9345,N_6013,N_6955);
nand U9346 (N_9346,N_7848,N_7267);
and U9347 (N_9347,N_7388,N_6359);
and U9348 (N_9348,N_7351,N_7406);
and U9349 (N_9349,N_7257,N_6359);
nor U9350 (N_9350,N_7971,N_6904);
xor U9351 (N_9351,N_7573,N_6985);
or U9352 (N_9352,N_7523,N_6136);
xnor U9353 (N_9353,N_7905,N_6507);
or U9354 (N_9354,N_6812,N_6302);
or U9355 (N_9355,N_7200,N_7523);
or U9356 (N_9356,N_6390,N_7068);
xor U9357 (N_9357,N_7355,N_6499);
and U9358 (N_9358,N_7037,N_6761);
xnor U9359 (N_9359,N_6105,N_6042);
or U9360 (N_9360,N_7651,N_7864);
or U9361 (N_9361,N_7768,N_7780);
nand U9362 (N_9362,N_6434,N_7430);
xnor U9363 (N_9363,N_6953,N_6808);
or U9364 (N_9364,N_7486,N_6027);
xnor U9365 (N_9365,N_7771,N_6778);
xnor U9366 (N_9366,N_7945,N_7380);
nand U9367 (N_9367,N_6939,N_6573);
nor U9368 (N_9368,N_6754,N_7360);
or U9369 (N_9369,N_6216,N_7213);
nand U9370 (N_9370,N_6313,N_7091);
nor U9371 (N_9371,N_7238,N_7839);
nand U9372 (N_9372,N_7600,N_6815);
nor U9373 (N_9373,N_6332,N_6861);
nor U9374 (N_9374,N_7350,N_6062);
nand U9375 (N_9375,N_6572,N_6471);
or U9376 (N_9376,N_6649,N_6578);
and U9377 (N_9377,N_6599,N_6323);
xnor U9378 (N_9378,N_6386,N_6644);
and U9379 (N_9379,N_6096,N_7592);
or U9380 (N_9380,N_6600,N_6645);
and U9381 (N_9381,N_6216,N_6149);
and U9382 (N_9382,N_7286,N_7754);
nand U9383 (N_9383,N_7378,N_6515);
xnor U9384 (N_9384,N_6702,N_6692);
nor U9385 (N_9385,N_7719,N_6828);
and U9386 (N_9386,N_6994,N_7703);
or U9387 (N_9387,N_6680,N_7513);
nor U9388 (N_9388,N_7086,N_6571);
and U9389 (N_9389,N_7020,N_6239);
and U9390 (N_9390,N_7436,N_7816);
xnor U9391 (N_9391,N_6131,N_7624);
nor U9392 (N_9392,N_6304,N_6244);
nor U9393 (N_9393,N_7006,N_7577);
xnor U9394 (N_9394,N_6384,N_6387);
nand U9395 (N_9395,N_7661,N_6201);
nor U9396 (N_9396,N_6538,N_6576);
nor U9397 (N_9397,N_6377,N_7440);
nand U9398 (N_9398,N_6589,N_6670);
nor U9399 (N_9399,N_7471,N_6640);
xor U9400 (N_9400,N_7922,N_6600);
nand U9401 (N_9401,N_7421,N_6916);
nor U9402 (N_9402,N_6547,N_6423);
nand U9403 (N_9403,N_7702,N_7897);
xnor U9404 (N_9404,N_7013,N_6396);
or U9405 (N_9405,N_6396,N_6599);
xnor U9406 (N_9406,N_7526,N_6060);
or U9407 (N_9407,N_7451,N_6156);
and U9408 (N_9408,N_6706,N_7412);
xnor U9409 (N_9409,N_6022,N_7140);
or U9410 (N_9410,N_7473,N_6499);
and U9411 (N_9411,N_7280,N_7173);
and U9412 (N_9412,N_6801,N_7173);
xnor U9413 (N_9413,N_7348,N_7508);
nor U9414 (N_9414,N_6558,N_6258);
xor U9415 (N_9415,N_6931,N_7890);
xnor U9416 (N_9416,N_7291,N_7874);
or U9417 (N_9417,N_7092,N_7548);
or U9418 (N_9418,N_6571,N_7409);
or U9419 (N_9419,N_7256,N_6285);
nand U9420 (N_9420,N_7207,N_7460);
and U9421 (N_9421,N_6105,N_6242);
nor U9422 (N_9422,N_7208,N_6059);
and U9423 (N_9423,N_6078,N_7107);
and U9424 (N_9424,N_7913,N_7900);
nand U9425 (N_9425,N_7284,N_7231);
or U9426 (N_9426,N_6400,N_7317);
and U9427 (N_9427,N_7836,N_6184);
xnor U9428 (N_9428,N_6500,N_6843);
xor U9429 (N_9429,N_6914,N_6908);
and U9430 (N_9430,N_7392,N_6765);
and U9431 (N_9431,N_6292,N_7602);
or U9432 (N_9432,N_7862,N_6013);
nor U9433 (N_9433,N_7293,N_6781);
and U9434 (N_9434,N_6516,N_6117);
xor U9435 (N_9435,N_7030,N_6399);
nor U9436 (N_9436,N_6632,N_7031);
nand U9437 (N_9437,N_6706,N_6908);
or U9438 (N_9438,N_7179,N_7209);
nand U9439 (N_9439,N_7440,N_7653);
and U9440 (N_9440,N_7460,N_7086);
and U9441 (N_9441,N_7523,N_6999);
xnor U9442 (N_9442,N_6157,N_7611);
nor U9443 (N_9443,N_6017,N_6616);
xor U9444 (N_9444,N_7857,N_7661);
or U9445 (N_9445,N_7760,N_7386);
nor U9446 (N_9446,N_7420,N_6491);
and U9447 (N_9447,N_7165,N_7352);
or U9448 (N_9448,N_7418,N_6193);
nand U9449 (N_9449,N_7438,N_6595);
nor U9450 (N_9450,N_7536,N_7151);
and U9451 (N_9451,N_6340,N_6724);
nor U9452 (N_9452,N_7283,N_6557);
nand U9453 (N_9453,N_6330,N_6130);
xnor U9454 (N_9454,N_6579,N_7617);
or U9455 (N_9455,N_7602,N_7243);
or U9456 (N_9456,N_6572,N_7243);
or U9457 (N_9457,N_6863,N_6599);
and U9458 (N_9458,N_7633,N_7337);
nor U9459 (N_9459,N_7930,N_6180);
and U9460 (N_9460,N_6689,N_7312);
or U9461 (N_9461,N_7258,N_7812);
and U9462 (N_9462,N_6954,N_7396);
nor U9463 (N_9463,N_7560,N_7037);
or U9464 (N_9464,N_6209,N_6123);
nor U9465 (N_9465,N_6888,N_6288);
nand U9466 (N_9466,N_6004,N_6012);
nand U9467 (N_9467,N_7756,N_6137);
and U9468 (N_9468,N_7243,N_6936);
and U9469 (N_9469,N_7715,N_6375);
nand U9470 (N_9470,N_6826,N_6824);
and U9471 (N_9471,N_7494,N_7472);
xor U9472 (N_9472,N_7136,N_6839);
nand U9473 (N_9473,N_6802,N_6583);
or U9474 (N_9474,N_7644,N_7376);
nor U9475 (N_9475,N_7220,N_6414);
or U9476 (N_9476,N_7194,N_6409);
nor U9477 (N_9477,N_7288,N_6511);
nor U9478 (N_9478,N_6051,N_7486);
nor U9479 (N_9479,N_6212,N_6307);
nand U9480 (N_9480,N_6015,N_7138);
nor U9481 (N_9481,N_7746,N_6982);
or U9482 (N_9482,N_7207,N_6661);
and U9483 (N_9483,N_7997,N_6667);
and U9484 (N_9484,N_7751,N_6125);
and U9485 (N_9485,N_6023,N_6484);
xor U9486 (N_9486,N_6659,N_7717);
nand U9487 (N_9487,N_7730,N_6926);
and U9488 (N_9488,N_6055,N_7775);
nand U9489 (N_9489,N_6448,N_6989);
and U9490 (N_9490,N_7978,N_6907);
and U9491 (N_9491,N_7423,N_6252);
nor U9492 (N_9492,N_7492,N_6513);
nor U9493 (N_9493,N_6569,N_7929);
and U9494 (N_9494,N_7850,N_7008);
and U9495 (N_9495,N_6407,N_6873);
and U9496 (N_9496,N_6613,N_7113);
nor U9497 (N_9497,N_6190,N_7243);
xnor U9498 (N_9498,N_7213,N_7265);
and U9499 (N_9499,N_7039,N_7653);
or U9500 (N_9500,N_7705,N_7036);
nor U9501 (N_9501,N_6248,N_6336);
or U9502 (N_9502,N_6627,N_7462);
and U9503 (N_9503,N_7582,N_7454);
and U9504 (N_9504,N_7758,N_6947);
nor U9505 (N_9505,N_7462,N_6362);
xor U9506 (N_9506,N_6434,N_6773);
or U9507 (N_9507,N_7154,N_6434);
and U9508 (N_9508,N_7117,N_6061);
xnor U9509 (N_9509,N_7654,N_6138);
nand U9510 (N_9510,N_6797,N_7190);
and U9511 (N_9511,N_6890,N_7600);
nand U9512 (N_9512,N_6517,N_6528);
xnor U9513 (N_9513,N_6876,N_6268);
nand U9514 (N_9514,N_7108,N_6027);
or U9515 (N_9515,N_7738,N_6200);
or U9516 (N_9516,N_7563,N_6698);
or U9517 (N_9517,N_6719,N_7779);
and U9518 (N_9518,N_6135,N_6832);
nand U9519 (N_9519,N_7603,N_6045);
or U9520 (N_9520,N_6539,N_6066);
xnor U9521 (N_9521,N_7902,N_7448);
or U9522 (N_9522,N_7111,N_7659);
and U9523 (N_9523,N_6880,N_6001);
nor U9524 (N_9524,N_7710,N_6844);
nor U9525 (N_9525,N_7126,N_6932);
nor U9526 (N_9526,N_7601,N_7977);
nand U9527 (N_9527,N_7995,N_6387);
xor U9528 (N_9528,N_6773,N_7304);
and U9529 (N_9529,N_7085,N_6604);
xor U9530 (N_9530,N_7831,N_7435);
xnor U9531 (N_9531,N_6691,N_7475);
and U9532 (N_9532,N_6173,N_6384);
or U9533 (N_9533,N_6840,N_6377);
nor U9534 (N_9534,N_7141,N_6398);
nand U9535 (N_9535,N_6818,N_6891);
nor U9536 (N_9536,N_6694,N_6528);
xnor U9537 (N_9537,N_6826,N_7578);
xnor U9538 (N_9538,N_7388,N_6585);
nor U9539 (N_9539,N_7229,N_7961);
nor U9540 (N_9540,N_7731,N_7420);
xor U9541 (N_9541,N_7643,N_7160);
nand U9542 (N_9542,N_6529,N_6353);
xor U9543 (N_9543,N_6341,N_6002);
or U9544 (N_9544,N_6114,N_7316);
or U9545 (N_9545,N_7126,N_7071);
nor U9546 (N_9546,N_7472,N_6193);
xor U9547 (N_9547,N_6570,N_6298);
and U9548 (N_9548,N_7640,N_6909);
nand U9549 (N_9549,N_6866,N_7381);
nor U9550 (N_9550,N_7354,N_7417);
nand U9551 (N_9551,N_7203,N_6628);
and U9552 (N_9552,N_6184,N_6506);
nand U9553 (N_9553,N_6087,N_6050);
xnor U9554 (N_9554,N_6999,N_7623);
or U9555 (N_9555,N_7528,N_7631);
nor U9556 (N_9556,N_6575,N_6423);
nor U9557 (N_9557,N_7042,N_7678);
nand U9558 (N_9558,N_7495,N_6077);
nor U9559 (N_9559,N_6607,N_6138);
nor U9560 (N_9560,N_6012,N_6954);
or U9561 (N_9561,N_7383,N_6076);
nor U9562 (N_9562,N_6495,N_6878);
nand U9563 (N_9563,N_7193,N_6287);
and U9564 (N_9564,N_7251,N_7238);
xnor U9565 (N_9565,N_6343,N_6142);
or U9566 (N_9566,N_7417,N_6599);
xnor U9567 (N_9567,N_6145,N_6759);
and U9568 (N_9568,N_7327,N_7463);
nor U9569 (N_9569,N_7911,N_6775);
nor U9570 (N_9570,N_6364,N_7099);
xor U9571 (N_9571,N_6782,N_6588);
nor U9572 (N_9572,N_7120,N_6681);
xnor U9573 (N_9573,N_7706,N_6608);
xor U9574 (N_9574,N_7159,N_6843);
nor U9575 (N_9575,N_7121,N_7933);
and U9576 (N_9576,N_6212,N_7197);
nand U9577 (N_9577,N_7358,N_6061);
nor U9578 (N_9578,N_6972,N_7577);
xnor U9579 (N_9579,N_7191,N_7631);
xnor U9580 (N_9580,N_6211,N_7849);
or U9581 (N_9581,N_6862,N_6784);
nor U9582 (N_9582,N_6324,N_6991);
xor U9583 (N_9583,N_6769,N_6165);
and U9584 (N_9584,N_6530,N_6112);
and U9585 (N_9585,N_6654,N_7576);
nand U9586 (N_9586,N_7205,N_6875);
nand U9587 (N_9587,N_6954,N_7143);
xnor U9588 (N_9588,N_6960,N_6967);
nand U9589 (N_9589,N_6601,N_7712);
and U9590 (N_9590,N_7606,N_7630);
or U9591 (N_9591,N_7060,N_7531);
nor U9592 (N_9592,N_6554,N_7745);
xnor U9593 (N_9593,N_7441,N_7253);
nor U9594 (N_9594,N_7149,N_7585);
nand U9595 (N_9595,N_6302,N_6310);
or U9596 (N_9596,N_7270,N_6397);
and U9597 (N_9597,N_7679,N_6568);
nand U9598 (N_9598,N_7529,N_6054);
nor U9599 (N_9599,N_7937,N_6464);
nand U9600 (N_9600,N_7355,N_7339);
and U9601 (N_9601,N_7354,N_6283);
nor U9602 (N_9602,N_6904,N_6913);
nor U9603 (N_9603,N_7907,N_7065);
xnor U9604 (N_9604,N_6326,N_7779);
and U9605 (N_9605,N_6501,N_7791);
or U9606 (N_9606,N_7436,N_6376);
xor U9607 (N_9607,N_6200,N_7369);
nor U9608 (N_9608,N_6086,N_7430);
xnor U9609 (N_9609,N_7063,N_7884);
nor U9610 (N_9610,N_6580,N_6311);
nand U9611 (N_9611,N_6627,N_6784);
and U9612 (N_9612,N_6505,N_7644);
nand U9613 (N_9613,N_7004,N_6899);
or U9614 (N_9614,N_7513,N_7913);
and U9615 (N_9615,N_6870,N_6593);
or U9616 (N_9616,N_7527,N_6273);
xor U9617 (N_9617,N_6934,N_6819);
or U9618 (N_9618,N_7976,N_6356);
nand U9619 (N_9619,N_6021,N_6422);
or U9620 (N_9620,N_6065,N_6395);
and U9621 (N_9621,N_7077,N_7706);
xor U9622 (N_9622,N_7844,N_7460);
and U9623 (N_9623,N_6399,N_7671);
or U9624 (N_9624,N_6835,N_6888);
or U9625 (N_9625,N_7325,N_6819);
nor U9626 (N_9626,N_7011,N_7813);
and U9627 (N_9627,N_6211,N_6203);
and U9628 (N_9628,N_7794,N_7199);
xnor U9629 (N_9629,N_7976,N_7885);
nor U9630 (N_9630,N_6299,N_7659);
xor U9631 (N_9631,N_6624,N_6804);
nand U9632 (N_9632,N_6770,N_6787);
xor U9633 (N_9633,N_7875,N_7261);
nor U9634 (N_9634,N_6572,N_6662);
or U9635 (N_9635,N_6931,N_7647);
nor U9636 (N_9636,N_6725,N_7914);
nor U9637 (N_9637,N_6782,N_7259);
or U9638 (N_9638,N_6796,N_6551);
nand U9639 (N_9639,N_6322,N_7225);
nand U9640 (N_9640,N_6831,N_6772);
nor U9641 (N_9641,N_6098,N_7152);
nand U9642 (N_9642,N_7510,N_6701);
and U9643 (N_9643,N_7468,N_7210);
or U9644 (N_9644,N_6648,N_7733);
or U9645 (N_9645,N_7535,N_7059);
and U9646 (N_9646,N_7171,N_6865);
xnor U9647 (N_9647,N_6485,N_6781);
nand U9648 (N_9648,N_6024,N_6933);
and U9649 (N_9649,N_6485,N_6712);
xnor U9650 (N_9650,N_7816,N_7482);
xor U9651 (N_9651,N_6688,N_7532);
xnor U9652 (N_9652,N_6341,N_7578);
nand U9653 (N_9653,N_7270,N_6469);
or U9654 (N_9654,N_7459,N_6328);
xor U9655 (N_9655,N_7142,N_6553);
or U9656 (N_9656,N_6174,N_6239);
and U9657 (N_9657,N_7507,N_7952);
xnor U9658 (N_9658,N_7309,N_7841);
or U9659 (N_9659,N_7163,N_7870);
or U9660 (N_9660,N_7069,N_6080);
nor U9661 (N_9661,N_6241,N_7791);
xnor U9662 (N_9662,N_6664,N_6413);
nand U9663 (N_9663,N_6413,N_7469);
nand U9664 (N_9664,N_6094,N_7253);
nand U9665 (N_9665,N_6744,N_7251);
xor U9666 (N_9666,N_6739,N_7821);
xor U9667 (N_9667,N_6251,N_6005);
nand U9668 (N_9668,N_7211,N_7731);
and U9669 (N_9669,N_6118,N_7090);
or U9670 (N_9670,N_7395,N_6147);
nor U9671 (N_9671,N_7304,N_7356);
or U9672 (N_9672,N_6852,N_6909);
nor U9673 (N_9673,N_6944,N_6809);
nand U9674 (N_9674,N_6748,N_6381);
xnor U9675 (N_9675,N_6763,N_6059);
nor U9676 (N_9676,N_7527,N_7391);
and U9677 (N_9677,N_7330,N_6582);
nor U9678 (N_9678,N_6589,N_7332);
and U9679 (N_9679,N_7327,N_6302);
nand U9680 (N_9680,N_7460,N_7343);
xor U9681 (N_9681,N_7388,N_6793);
xnor U9682 (N_9682,N_6033,N_6044);
xnor U9683 (N_9683,N_7348,N_7120);
and U9684 (N_9684,N_7228,N_6336);
xnor U9685 (N_9685,N_6308,N_6397);
and U9686 (N_9686,N_7050,N_6943);
or U9687 (N_9687,N_7148,N_7090);
or U9688 (N_9688,N_6297,N_7878);
xor U9689 (N_9689,N_6319,N_7217);
or U9690 (N_9690,N_7713,N_7533);
and U9691 (N_9691,N_7749,N_6803);
or U9692 (N_9692,N_6958,N_6621);
or U9693 (N_9693,N_7109,N_7725);
xnor U9694 (N_9694,N_7202,N_7852);
nand U9695 (N_9695,N_6773,N_6941);
xor U9696 (N_9696,N_7529,N_7025);
xor U9697 (N_9697,N_6418,N_7768);
or U9698 (N_9698,N_7064,N_7509);
nor U9699 (N_9699,N_7488,N_7305);
nand U9700 (N_9700,N_6874,N_6733);
or U9701 (N_9701,N_6941,N_7204);
nor U9702 (N_9702,N_6226,N_7568);
and U9703 (N_9703,N_6715,N_6415);
xor U9704 (N_9704,N_6424,N_6698);
nand U9705 (N_9705,N_7352,N_7559);
nand U9706 (N_9706,N_6213,N_6628);
or U9707 (N_9707,N_6408,N_6527);
nor U9708 (N_9708,N_6878,N_7253);
or U9709 (N_9709,N_6835,N_7582);
nand U9710 (N_9710,N_6748,N_7277);
xor U9711 (N_9711,N_7400,N_7493);
and U9712 (N_9712,N_7875,N_6829);
and U9713 (N_9713,N_7831,N_7358);
or U9714 (N_9714,N_7838,N_6096);
nand U9715 (N_9715,N_6451,N_6993);
or U9716 (N_9716,N_7762,N_7694);
nor U9717 (N_9717,N_7232,N_6033);
nor U9718 (N_9718,N_7161,N_7436);
and U9719 (N_9719,N_7904,N_6863);
and U9720 (N_9720,N_7189,N_7741);
nor U9721 (N_9721,N_6710,N_6244);
and U9722 (N_9722,N_6127,N_7423);
or U9723 (N_9723,N_6104,N_7596);
or U9724 (N_9724,N_7874,N_7740);
nand U9725 (N_9725,N_7361,N_6582);
or U9726 (N_9726,N_7069,N_6757);
nand U9727 (N_9727,N_7129,N_7248);
and U9728 (N_9728,N_7360,N_7934);
or U9729 (N_9729,N_6358,N_6431);
and U9730 (N_9730,N_7458,N_6732);
nand U9731 (N_9731,N_7067,N_6989);
nand U9732 (N_9732,N_6129,N_7403);
or U9733 (N_9733,N_7921,N_6226);
or U9734 (N_9734,N_6268,N_7536);
xor U9735 (N_9735,N_7160,N_7830);
and U9736 (N_9736,N_6955,N_7992);
nor U9737 (N_9737,N_6844,N_6860);
or U9738 (N_9738,N_7351,N_6937);
and U9739 (N_9739,N_6910,N_6896);
or U9740 (N_9740,N_7202,N_7090);
xnor U9741 (N_9741,N_7293,N_6319);
nor U9742 (N_9742,N_6758,N_6821);
nand U9743 (N_9743,N_6338,N_7228);
nand U9744 (N_9744,N_7827,N_6326);
nand U9745 (N_9745,N_6390,N_6365);
nor U9746 (N_9746,N_7274,N_6881);
nor U9747 (N_9747,N_7415,N_6832);
nand U9748 (N_9748,N_7840,N_7679);
nand U9749 (N_9749,N_6493,N_7333);
or U9750 (N_9750,N_6740,N_6056);
and U9751 (N_9751,N_7650,N_6029);
nor U9752 (N_9752,N_6323,N_6339);
nand U9753 (N_9753,N_7808,N_6110);
nor U9754 (N_9754,N_7528,N_6264);
and U9755 (N_9755,N_7257,N_7950);
or U9756 (N_9756,N_7637,N_6058);
nand U9757 (N_9757,N_6579,N_6667);
or U9758 (N_9758,N_6287,N_6307);
nand U9759 (N_9759,N_6738,N_6815);
and U9760 (N_9760,N_6212,N_7912);
and U9761 (N_9761,N_7639,N_6602);
xnor U9762 (N_9762,N_7887,N_7958);
nor U9763 (N_9763,N_7957,N_6540);
and U9764 (N_9764,N_6866,N_7982);
nand U9765 (N_9765,N_7939,N_7417);
and U9766 (N_9766,N_7300,N_6751);
or U9767 (N_9767,N_6457,N_6282);
nand U9768 (N_9768,N_7253,N_7068);
nor U9769 (N_9769,N_7567,N_6078);
nand U9770 (N_9770,N_6066,N_6702);
or U9771 (N_9771,N_7128,N_6253);
nand U9772 (N_9772,N_6969,N_6134);
xnor U9773 (N_9773,N_6793,N_6756);
and U9774 (N_9774,N_6533,N_7801);
nand U9775 (N_9775,N_6089,N_6248);
nand U9776 (N_9776,N_6288,N_7084);
nand U9777 (N_9777,N_6473,N_6401);
or U9778 (N_9778,N_7180,N_6171);
and U9779 (N_9779,N_7176,N_7781);
nand U9780 (N_9780,N_7154,N_7233);
nand U9781 (N_9781,N_7690,N_7709);
or U9782 (N_9782,N_7568,N_7934);
and U9783 (N_9783,N_7518,N_6426);
and U9784 (N_9784,N_6412,N_7970);
nand U9785 (N_9785,N_7225,N_7356);
or U9786 (N_9786,N_7647,N_6469);
nor U9787 (N_9787,N_6663,N_7721);
or U9788 (N_9788,N_6885,N_6301);
and U9789 (N_9789,N_7676,N_7296);
xor U9790 (N_9790,N_6519,N_6240);
nand U9791 (N_9791,N_7890,N_7070);
or U9792 (N_9792,N_7990,N_7224);
or U9793 (N_9793,N_6594,N_6281);
nand U9794 (N_9794,N_6732,N_6040);
nand U9795 (N_9795,N_7879,N_6455);
or U9796 (N_9796,N_6147,N_6334);
xor U9797 (N_9797,N_6112,N_7721);
xor U9798 (N_9798,N_6499,N_6568);
nand U9799 (N_9799,N_6051,N_6586);
nor U9800 (N_9800,N_6819,N_7589);
and U9801 (N_9801,N_6143,N_7308);
and U9802 (N_9802,N_7933,N_6353);
nor U9803 (N_9803,N_6257,N_7606);
nand U9804 (N_9804,N_6504,N_6659);
xor U9805 (N_9805,N_7917,N_6515);
and U9806 (N_9806,N_6905,N_7529);
xor U9807 (N_9807,N_6263,N_7996);
or U9808 (N_9808,N_6836,N_6896);
nand U9809 (N_9809,N_6102,N_6336);
or U9810 (N_9810,N_7478,N_6642);
or U9811 (N_9811,N_7212,N_7566);
nor U9812 (N_9812,N_6393,N_7439);
nand U9813 (N_9813,N_7355,N_6849);
nor U9814 (N_9814,N_6181,N_6844);
nor U9815 (N_9815,N_6145,N_6979);
or U9816 (N_9816,N_7195,N_7930);
or U9817 (N_9817,N_7193,N_7005);
and U9818 (N_9818,N_7101,N_6035);
or U9819 (N_9819,N_7918,N_7413);
nor U9820 (N_9820,N_7237,N_7921);
and U9821 (N_9821,N_6807,N_6008);
and U9822 (N_9822,N_7903,N_7592);
xor U9823 (N_9823,N_6048,N_7473);
and U9824 (N_9824,N_7869,N_7346);
or U9825 (N_9825,N_7566,N_7021);
nor U9826 (N_9826,N_7691,N_7807);
nand U9827 (N_9827,N_6216,N_6253);
or U9828 (N_9828,N_7186,N_6706);
xor U9829 (N_9829,N_6904,N_6971);
and U9830 (N_9830,N_7280,N_7006);
nor U9831 (N_9831,N_6296,N_7933);
xor U9832 (N_9832,N_6847,N_7766);
or U9833 (N_9833,N_7239,N_6435);
nor U9834 (N_9834,N_6472,N_6586);
nor U9835 (N_9835,N_7435,N_7013);
nor U9836 (N_9836,N_7683,N_7767);
and U9837 (N_9837,N_6753,N_6244);
or U9838 (N_9838,N_7585,N_6497);
and U9839 (N_9839,N_7534,N_6862);
and U9840 (N_9840,N_7775,N_6527);
nor U9841 (N_9841,N_6301,N_6356);
or U9842 (N_9842,N_6589,N_6793);
nor U9843 (N_9843,N_7762,N_6977);
and U9844 (N_9844,N_6299,N_6369);
or U9845 (N_9845,N_7610,N_7078);
or U9846 (N_9846,N_6922,N_6777);
xor U9847 (N_9847,N_7431,N_7918);
nor U9848 (N_9848,N_6140,N_7522);
nor U9849 (N_9849,N_6944,N_6069);
and U9850 (N_9850,N_6479,N_6478);
and U9851 (N_9851,N_7456,N_6321);
nand U9852 (N_9852,N_7425,N_6540);
nand U9853 (N_9853,N_6665,N_7783);
nor U9854 (N_9854,N_6587,N_7346);
and U9855 (N_9855,N_6108,N_6575);
nor U9856 (N_9856,N_7725,N_6575);
nand U9857 (N_9857,N_6783,N_6147);
nand U9858 (N_9858,N_6677,N_6365);
nor U9859 (N_9859,N_7246,N_7536);
xor U9860 (N_9860,N_7780,N_6388);
nand U9861 (N_9861,N_7297,N_7733);
or U9862 (N_9862,N_7947,N_7636);
and U9863 (N_9863,N_6485,N_6005);
nor U9864 (N_9864,N_6441,N_6403);
or U9865 (N_9865,N_7950,N_7831);
nand U9866 (N_9866,N_7856,N_6738);
nor U9867 (N_9867,N_6113,N_7714);
nand U9868 (N_9868,N_7098,N_6279);
xor U9869 (N_9869,N_7589,N_6687);
nor U9870 (N_9870,N_6883,N_6543);
nand U9871 (N_9871,N_7286,N_7170);
nand U9872 (N_9872,N_7117,N_6332);
and U9873 (N_9873,N_6015,N_7362);
or U9874 (N_9874,N_6771,N_7953);
nor U9875 (N_9875,N_7432,N_7780);
and U9876 (N_9876,N_6282,N_6161);
and U9877 (N_9877,N_6776,N_6565);
xor U9878 (N_9878,N_7525,N_7656);
nor U9879 (N_9879,N_7948,N_7475);
and U9880 (N_9880,N_7890,N_6766);
nand U9881 (N_9881,N_6918,N_7286);
and U9882 (N_9882,N_6292,N_7488);
nor U9883 (N_9883,N_7817,N_7211);
or U9884 (N_9884,N_6997,N_6587);
nand U9885 (N_9885,N_6227,N_7787);
xor U9886 (N_9886,N_7627,N_6359);
and U9887 (N_9887,N_6772,N_6647);
and U9888 (N_9888,N_6487,N_7481);
xor U9889 (N_9889,N_7330,N_7148);
and U9890 (N_9890,N_6642,N_6870);
nand U9891 (N_9891,N_6725,N_7018);
and U9892 (N_9892,N_6521,N_7698);
or U9893 (N_9893,N_7722,N_7827);
nor U9894 (N_9894,N_7801,N_6639);
nor U9895 (N_9895,N_7891,N_7488);
and U9896 (N_9896,N_7408,N_6915);
xor U9897 (N_9897,N_7439,N_6789);
and U9898 (N_9898,N_6966,N_7778);
and U9899 (N_9899,N_6339,N_7125);
xor U9900 (N_9900,N_7031,N_7379);
nor U9901 (N_9901,N_6348,N_7203);
or U9902 (N_9902,N_6760,N_6631);
nand U9903 (N_9903,N_6589,N_7686);
nor U9904 (N_9904,N_6462,N_7755);
nor U9905 (N_9905,N_6207,N_6362);
xor U9906 (N_9906,N_7609,N_6551);
or U9907 (N_9907,N_7515,N_7007);
nand U9908 (N_9908,N_7636,N_7261);
nand U9909 (N_9909,N_7462,N_6424);
nor U9910 (N_9910,N_6687,N_6115);
nand U9911 (N_9911,N_6835,N_7113);
xor U9912 (N_9912,N_6212,N_7114);
or U9913 (N_9913,N_6016,N_7725);
or U9914 (N_9914,N_6123,N_6496);
nand U9915 (N_9915,N_7841,N_6285);
or U9916 (N_9916,N_7360,N_6084);
or U9917 (N_9917,N_7535,N_7455);
and U9918 (N_9918,N_7384,N_7923);
nor U9919 (N_9919,N_7235,N_6313);
nand U9920 (N_9920,N_6521,N_7139);
nand U9921 (N_9921,N_6116,N_6518);
nor U9922 (N_9922,N_6524,N_7595);
xor U9923 (N_9923,N_7401,N_6892);
or U9924 (N_9924,N_6387,N_6851);
nor U9925 (N_9925,N_7605,N_7887);
nor U9926 (N_9926,N_6614,N_7291);
or U9927 (N_9927,N_6570,N_6807);
and U9928 (N_9928,N_6021,N_7316);
xnor U9929 (N_9929,N_6148,N_7864);
and U9930 (N_9930,N_7501,N_7318);
nand U9931 (N_9931,N_7790,N_7035);
or U9932 (N_9932,N_6167,N_7932);
and U9933 (N_9933,N_7863,N_6934);
nand U9934 (N_9934,N_6543,N_6793);
and U9935 (N_9935,N_6746,N_6446);
nand U9936 (N_9936,N_6081,N_6146);
nor U9937 (N_9937,N_6444,N_7170);
nor U9938 (N_9938,N_6215,N_6158);
nor U9939 (N_9939,N_6819,N_6464);
xor U9940 (N_9940,N_7768,N_6390);
nand U9941 (N_9941,N_7645,N_7178);
xor U9942 (N_9942,N_6398,N_7591);
and U9943 (N_9943,N_7622,N_6508);
nand U9944 (N_9944,N_7512,N_6900);
and U9945 (N_9945,N_6787,N_6093);
nand U9946 (N_9946,N_7149,N_6939);
nand U9947 (N_9947,N_6284,N_6942);
xor U9948 (N_9948,N_6828,N_6806);
nand U9949 (N_9949,N_7284,N_6242);
or U9950 (N_9950,N_6092,N_7964);
nor U9951 (N_9951,N_6257,N_7337);
nor U9952 (N_9952,N_6862,N_7724);
or U9953 (N_9953,N_6946,N_7231);
nor U9954 (N_9954,N_7619,N_6678);
xnor U9955 (N_9955,N_6758,N_6043);
xnor U9956 (N_9956,N_7148,N_6706);
and U9957 (N_9957,N_7514,N_7896);
nor U9958 (N_9958,N_6333,N_6520);
or U9959 (N_9959,N_7123,N_7844);
nand U9960 (N_9960,N_7419,N_7071);
and U9961 (N_9961,N_6056,N_7042);
nand U9962 (N_9962,N_6411,N_7681);
and U9963 (N_9963,N_6037,N_7951);
nor U9964 (N_9964,N_6874,N_6820);
nand U9965 (N_9965,N_6690,N_7590);
xnor U9966 (N_9966,N_7838,N_7994);
and U9967 (N_9967,N_6701,N_6086);
and U9968 (N_9968,N_6612,N_7931);
xor U9969 (N_9969,N_7781,N_7730);
nand U9970 (N_9970,N_7786,N_6116);
xor U9971 (N_9971,N_6459,N_7174);
nor U9972 (N_9972,N_7111,N_6543);
xor U9973 (N_9973,N_7537,N_7744);
xor U9974 (N_9974,N_6345,N_6084);
or U9975 (N_9975,N_7409,N_7685);
xor U9976 (N_9976,N_7743,N_6869);
or U9977 (N_9977,N_6829,N_6860);
xnor U9978 (N_9978,N_6266,N_7682);
xnor U9979 (N_9979,N_6294,N_6063);
xnor U9980 (N_9980,N_7055,N_7414);
nand U9981 (N_9981,N_6011,N_6734);
nor U9982 (N_9982,N_7212,N_7753);
and U9983 (N_9983,N_6031,N_6575);
xor U9984 (N_9984,N_6164,N_6560);
and U9985 (N_9985,N_7697,N_7221);
and U9986 (N_9986,N_6670,N_7224);
or U9987 (N_9987,N_7135,N_6021);
nand U9988 (N_9988,N_6457,N_6320);
nand U9989 (N_9989,N_7692,N_7134);
nor U9990 (N_9990,N_6706,N_6956);
and U9991 (N_9991,N_6377,N_6108);
and U9992 (N_9992,N_7061,N_6632);
nand U9993 (N_9993,N_7052,N_7059);
and U9994 (N_9994,N_7428,N_7937);
nor U9995 (N_9995,N_6906,N_6573);
nor U9996 (N_9996,N_6260,N_6407);
nand U9997 (N_9997,N_7340,N_6337);
nor U9998 (N_9998,N_6257,N_7087);
and U9999 (N_9999,N_6545,N_7871);
nand U10000 (N_10000,N_9260,N_8020);
nor U10001 (N_10001,N_9841,N_9502);
nor U10002 (N_10002,N_9479,N_9089);
xor U10003 (N_10003,N_8737,N_9995);
nand U10004 (N_10004,N_9946,N_9092);
nor U10005 (N_10005,N_8132,N_9126);
and U10006 (N_10006,N_9111,N_8895);
nor U10007 (N_10007,N_9748,N_9333);
xor U10008 (N_10008,N_9085,N_9736);
nand U10009 (N_10009,N_9977,N_8182);
xnor U10010 (N_10010,N_8559,N_8011);
or U10011 (N_10011,N_9945,N_8119);
nand U10012 (N_10012,N_9372,N_8812);
xnor U10013 (N_10013,N_9005,N_8898);
and U10014 (N_10014,N_9919,N_9883);
and U10015 (N_10015,N_8708,N_8497);
or U10016 (N_10016,N_8344,N_9076);
nor U10017 (N_10017,N_9271,N_8078);
nor U10018 (N_10018,N_9644,N_8406);
and U10019 (N_10019,N_9710,N_8069);
or U10020 (N_10020,N_9322,N_9061);
xor U10021 (N_10021,N_8310,N_8545);
or U10022 (N_10022,N_8756,N_8338);
nand U10023 (N_10023,N_8611,N_9589);
and U10024 (N_10024,N_9412,N_9454);
xnor U10025 (N_10025,N_9519,N_8588);
and U10026 (N_10026,N_9593,N_8177);
xor U10027 (N_10027,N_9052,N_8876);
nor U10028 (N_10028,N_8472,N_8946);
and U10029 (N_10029,N_8195,N_8867);
and U10030 (N_10030,N_8672,N_8924);
or U10031 (N_10031,N_9912,N_8302);
nor U10032 (N_10032,N_9166,N_8139);
and U10033 (N_10033,N_8724,N_8998);
and U10034 (N_10034,N_8114,N_8115);
nand U10035 (N_10035,N_8465,N_8087);
nand U10036 (N_10036,N_8145,N_8595);
xor U10037 (N_10037,N_8467,N_9828);
or U10038 (N_10038,N_9933,N_8795);
xnor U10039 (N_10039,N_9444,N_8318);
nor U10040 (N_10040,N_9928,N_9048);
nand U10041 (N_10041,N_9926,N_8009);
and U10042 (N_10042,N_9304,N_9764);
xor U10043 (N_10043,N_9953,N_9623);
nor U10044 (N_10044,N_8024,N_9442);
and U10045 (N_10045,N_8074,N_9493);
nand U10046 (N_10046,N_9836,N_9905);
and U10047 (N_10047,N_8646,N_9208);
or U10048 (N_10048,N_9701,N_8824);
nor U10049 (N_10049,N_8975,N_8710);
xor U10050 (N_10050,N_8235,N_9998);
nor U10051 (N_10051,N_9996,N_9607);
or U10052 (N_10052,N_9433,N_8413);
or U10053 (N_10053,N_9878,N_9962);
nor U10054 (N_10054,N_8520,N_8977);
nand U10055 (N_10055,N_9820,N_9272);
xor U10056 (N_10056,N_8927,N_9706);
or U10057 (N_10057,N_9730,N_9573);
nand U10058 (N_10058,N_9380,N_8333);
xnor U10059 (N_10059,N_8689,N_9936);
or U10060 (N_10060,N_9687,N_8326);
or U10061 (N_10061,N_9394,N_8916);
xnor U10062 (N_10062,N_9608,N_8965);
xor U10063 (N_10063,N_9338,N_9232);
and U10064 (N_10064,N_8905,N_8103);
xor U10065 (N_10065,N_9053,N_9938);
and U10066 (N_10066,N_8436,N_9478);
and U10067 (N_10067,N_8202,N_8381);
xor U10068 (N_10068,N_8889,N_8675);
nand U10069 (N_10069,N_9080,N_8397);
nand U10070 (N_10070,N_8451,N_9787);
or U10071 (N_10071,N_8800,N_8627);
or U10072 (N_10072,N_9167,N_8586);
xor U10073 (N_10073,N_9075,N_8297);
xnor U10074 (N_10074,N_8967,N_8726);
and U10075 (N_10075,N_9255,N_9657);
xor U10076 (N_10076,N_8232,N_9050);
nand U10077 (N_10077,N_8718,N_8517);
and U10078 (N_10078,N_8912,N_8222);
nor U10079 (N_10079,N_9279,N_8692);
nor U10080 (N_10080,N_8906,N_9062);
and U10081 (N_10081,N_8879,N_8862);
xnor U10082 (N_10082,N_9723,N_9885);
xnor U10083 (N_10083,N_8529,N_8493);
or U10084 (N_10084,N_9678,N_9504);
and U10085 (N_10085,N_8201,N_8623);
nor U10086 (N_10086,N_8254,N_9428);
nor U10087 (N_10087,N_9758,N_8051);
nor U10088 (N_10088,N_8583,N_8854);
nand U10089 (N_10089,N_9720,N_8825);
or U10090 (N_10090,N_9219,N_8942);
xor U10091 (N_10091,N_8709,N_8711);
or U10092 (N_10092,N_8606,N_8416);
nor U10093 (N_10093,N_8341,N_9567);
nor U10094 (N_10094,N_8037,N_8964);
nand U10095 (N_10095,N_8666,N_8094);
or U10096 (N_10096,N_8288,N_9940);
xor U10097 (N_10097,N_9273,N_9671);
and U10098 (N_10098,N_8358,N_8766);
and U10099 (N_10099,N_9106,N_9339);
nor U10100 (N_10100,N_9491,N_8925);
or U10101 (N_10101,N_8379,N_9588);
nand U10102 (N_10102,N_9229,N_9328);
nand U10103 (N_10103,N_8619,N_9527);
xor U10104 (N_10104,N_8022,N_9420);
xor U10105 (N_10105,N_9004,N_8872);
xor U10106 (N_10106,N_8340,N_9287);
and U10107 (N_10107,N_9530,N_8356);
nand U10108 (N_10108,N_8374,N_8429);
xor U10109 (N_10109,N_8440,N_9030);
xnor U10110 (N_10110,N_9526,N_9713);
nor U10111 (N_10111,N_8732,N_9976);
nand U10112 (N_10112,N_8866,N_9244);
or U10113 (N_10113,N_8231,N_9595);
or U10114 (N_10114,N_8079,N_9199);
xnor U10115 (N_10115,N_9741,N_9384);
or U10116 (N_10116,N_8439,N_8161);
nand U10117 (N_10117,N_9195,N_8597);
nand U10118 (N_10118,N_8428,N_9019);
xor U10119 (N_10119,N_8016,N_8739);
nor U10120 (N_10120,N_9297,N_8803);
or U10121 (N_10121,N_8410,N_8747);
xor U10122 (N_10122,N_9856,N_8057);
nand U10123 (N_10123,N_9397,N_8607);
xor U10124 (N_10124,N_8881,N_8170);
nand U10125 (N_10125,N_8295,N_8658);
nor U10126 (N_10126,N_8647,N_9869);
and U10127 (N_10127,N_8938,N_9499);
nand U10128 (N_10128,N_9174,N_8313);
nor U10129 (N_10129,N_8858,N_8105);
xnor U10130 (N_10130,N_9042,N_9973);
and U10131 (N_10131,N_9664,N_9991);
nor U10132 (N_10132,N_9718,N_9555);
or U10133 (N_10133,N_9746,N_8503);
nor U10134 (N_10134,N_9637,N_8043);
xnor U10135 (N_10135,N_8352,N_8407);
nand U10136 (N_10136,N_8420,N_9214);
and U10137 (N_10137,N_9296,N_8637);
nor U10138 (N_10138,N_8990,N_8499);
nand U10139 (N_10139,N_8549,N_8697);
nor U10140 (N_10140,N_9190,N_9942);
and U10141 (N_10141,N_9847,N_9717);
and U10142 (N_10142,N_9781,N_9377);
nor U10143 (N_10143,N_9268,N_8631);
or U10144 (N_10144,N_9543,N_8952);
nand U10145 (N_10145,N_9362,N_9775);
nor U10146 (N_10146,N_8515,N_9778);
or U10147 (N_10147,N_8426,N_8822);
or U10148 (N_10148,N_8994,N_9979);
nor U10149 (N_10149,N_9823,N_9385);
xnor U10150 (N_10150,N_9686,N_9675);
nor U10151 (N_10151,N_8810,N_9763);
nand U10152 (N_10152,N_8980,N_8495);
xor U10153 (N_10153,N_8017,N_9586);
nor U10154 (N_10154,N_9674,N_8956);
xnor U10155 (N_10155,N_9321,N_8028);
and U10156 (N_10156,N_8554,N_8186);
nor U10157 (N_10157,N_8284,N_9127);
or U10158 (N_10158,N_8518,N_9281);
nor U10159 (N_10159,N_8476,N_9342);
or U10160 (N_10160,N_9165,N_8477);
nor U10161 (N_10161,N_9063,N_9306);
nor U10162 (N_10162,N_9120,N_8189);
xor U10163 (N_10163,N_8620,N_9189);
nor U10164 (N_10164,N_8757,N_9057);
or U10165 (N_10165,N_9269,N_9348);
xor U10166 (N_10166,N_8243,N_9753);
nor U10167 (N_10167,N_9603,N_9851);
or U10168 (N_10168,N_9920,N_9997);
or U10169 (N_10169,N_9114,N_8802);
nor U10170 (N_10170,N_8579,N_9197);
and U10171 (N_10171,N_8147,N_9719);
nor U10172 (N_10172,N_9970,N_8897);
and U10173 (N_10173,N_9295,N_8015);
or U10174 (N_10174,N_8578,N_9669);
or U10175 (N_10175,N_9735,N_9954);
xor U10176 (N_10176,N_8963,N_8856);
nand U10177 (N_10177,N_8274,N_9855);
xor U10178 (N_10178,N_9797,N_8699);
nand U10179 (N_10179,N_9066,N_8608);
xor U10180 (N_10180,N_8509,N_9662);
or U10181 (N_10181,N_8304,N_9916);
xnor U10182 (N_10182,N_8062,N_9568);
nand U10183 (N_10183,N_9756,N_9474);
xnor U10184 (N_10184,N_9274,N_9750);
xor U10185 (N_10185,N_8883,N_9948);
xor U10186 (N_10186,N_8654,N_8151);
or U10187 (N_10187,N_9960,N_8328);
xnor U10188 (N_10188,N_8514,N_9186);
and U10189 (N_10189,N_8593,N_8817);
or U10190 (N_10190,N_9356,N_8797);
and U10191 (N_10191,N_8601,N_8749);
and U10192 (N_10192,N_9776,N_9814);
and U10193 (N_10193,N_9248,N_9233);
and U10194 (N_10194,N_9346,N_9284);
and U10195 (N_10195,N_8865,N_9930);
nor U10196 (N_10196,N_8241,N_8835);
or U10197 (N_10197,N_9622,N_9947);
nand U10198 (N_10198,N_9032,N_8798);
nor U10199 (N_10199,N_8969,N_9350);
and U10200 (N_10200,N_9316,N_9635);
xor U10201 (N_10201,N_9015,N_8142);
nand U10202 (N_10202,N_9286,N_9925);
and U10203 (N_10203,N_9477,N_9007);
nand U10204 (N_10204,N_9819,N_8134);
xnor U10205 (N_10205,N_8863,N_8226);
and U10206 (N_10206,N_8774,N_9860);
nand U10207 (N_10207,N_8199,N_8108);
nand U10208 (N_10208,N_8633,N_8783);
or U10209 (N_10209,N_8536,N_9138);
and U10210 (N_10210,N_9506,N_9508);
and U10211 (N_10211,N_8796,N_8026);
and U10212 (N_10212,N_8471,N_8175);
nor U10213 (N_10213,N_9927,N_8792);
xnor U10214 (N_10214,N_9411,N_9204);
nor U10215 (N_10215,N_8673,N_9722);
or U10216 (N_10216,N_8148,N_8890);
nor U10217 (N_10217,N_9359,N_8433);
nand U10218 (N_10218,N_8459,N_8861);
nor U10219 (N_10219,N_9067,N_8042);
nor U10220 (N_10220,N_8126,N_8808);
xnor U10221 (N_10221,N_8978,N_9108);
xor U10222 (N_10222,N_9026,N_8716);
or U10223 (N_10223,N_9312,N_9002);
xor U10224 (N_10224,N_9207,N_8355);
nor U10225 (N_10225,N_8248,N_8762);
xor U10226 (N_10226,N_9645,N_9517);
nor U10227 (N_10227,N_9949,N_8256);
or U10228 (N_10228,N_8287,N_8268);
and U10229 (N_10229,N_9223,N_8784);
and U10230 (N_10230,N_8286,N_9198);
xor U10231 (N_10231,N_8930,N_9305);
nor U10232 (N_10232,N_8887,N_8704);
and U10233 (N_10233,N_8408,N_9613);
xnor U10234 (N_10234,N_8933,N_8342);
nor U10235 (N_10235,N_9658,N_8884);
nand U10236 (N_10236,N_8204,N_8192);
xor U10237 (N_10237,N_9886,N_9768);
nand U10238 (N_10238,N_8343,N_9472);
nor U10239 (N_10239,N_9914,N_9971);
nor U10240 (N_10240,N_9587,N_8306);
or U10241 (N_10241,N_9760,N_8748);
nand U10242 (N_10242,N_9931,N_8188);
xnor U10243 (N_10243,N_9033,N_8706);
and U10244 (N_10244,N_9740,N_9465);
nor U10245 (N_10245,N_8090,N_9476);
nor U10246 (N_10246,N_9447,N_9558);
nand U10247 (N_10247,N_8077,N_9632);
nor U10248 (N_10248,N_8533,N_8713);
xor U10249 (N_10249,N_9395,N_9239);
xnor U10250 (N_10250,N_8655,N_8375);
and U10251 (N_10251,N_9553,N_9352);
or U10252 (N_10252,N_8357,N_8568);
xnor U10253 (N_10253,N_8215,N_9090);
nand U10254 (N_10254,N_9105,N_8164);
nand U10255 (N_10255,N_8460,N_9020);
and U10256 (N_10256,N_8855,N_8537);
and U10257 (N_10257,N_8411,N_9659);
and U10258 (N_10258,N_9791,N_9135);
or U10259 (N_10259,N_8903,N_8380);
nand U10260 (N_10260,N_8733,N_9488);
xor U10261 (N_10261,N_9959,N_9404);
or U10262 (N_10262,N_8991,N_9749);
nand U10263 (N_10263,N_9974,N_9552);
and U10264 (N_10264,N_8255,N_9993);
nand U10265 (N_10265,N_9846,N_9620);
and U10266 (N_10266,N_8725,N_9141);
nand U10267 (N_10267,N_8829,N_9745);
and U10268 (N_10268,N_8849,N_8636);
nand U10269 (N_10269,N_8085,N_9184);
xnor U10270 (N_10270,N_9387,N_8919);
and U10271 (N_10271,N_9879,N_9254);
and U10272 (N_10272,N_9142,N_9857);
or U10273 (N_10273,N_8104,N_8316);
xor U10274 (N_10274,N_9439,N_8169);
nand U10275 (N_10275,N_9897,N_8320);
or U10276 (N_10276,N_9899,N_8298);
nor U10277 (N_10277,N_8183,N_9624);
or U10278 (N_10278,N_8639,N_9731);
nor U10279 (N_10279,N_8129,N_8837);
nor U10280 (N_10280,N_9770,N_8038);
and U10281 (N_10281,N_9179,N_9688);
and U10282 (N_10282,N_9450,N_8696);
and U10283 (N_10283,N_9824,N_8047);
or U10284 (N_10284,N_8594,N_8642);
xnor U10285 (N_10285,N_8546,N_8613);
and U10286 (N_10286,N_9086,N_8029);
xnor U10287 (N_10287,N_8216,N_9018);
nor U10288 (N_10288,N_9596,N_8084);
or U10289 (N_10289,N_8973,N_9460);
or U10290 (N_10290,N_8446,N_8957);
xor U10291 (N_10291,N_8360,N_8441);
nand U10292 (N_10292,N_8698,N_8067);
nor U10293 (N_10293,N_9400,N_8768);
or U10294 (N_10294,N_8213,N_8736);
or U10295 (N_10295,N_9652,N_8896);
nand U10296 (N_10296,N_9732,N_8144);
xnor U10297 (N_10297,N_8913,N_8682);
nand U10298 (N_10298,N_9503,N_8609);
nand U10299 (N_10299,N_9351,N_9044);
nand U10300 (N_10300,N_8684,N_9743);
or U10301 (N_10301,N_8772,N_8412);
nor U10302 (N_10302,N_9366,N_9434);
or U10303 (N_10303,N_8048,N_9803);
nand U10304 (N_10304,N_9577,N_9104);
or U10305 (N_10305,N_8120,N_9369);
xor U10306 (N_10306,N_9882,N_8309);
or U10307 (N_10307,N_9839,N_8442);
and U10308 (N_10308,N_8150,N_8353);
nor U10309 (N_10309,N_8373,N_8218);
xor U10310 (N_10310,N_8519,N_8418);
or U10311 (N_10311,N_9655,N_9525);
and U10312 (N_10312,N_8308,N_9415);
and U10313 (N_10313,N_9110,N_9694);
nand U10314 (N_10314,N_9677,N_8700);
xor U10315 (N_10315,N_8670,N_9148);
and U10316 (N_10316,N_9969,N_9193);
xnor U10317 (N_10317,N_9082,N_9074);
nor U10318 (N_10318,N_8417,N_9944);
xnor U10319 (N_10319,N_9070,N_9457);
nand U10320 (N_10320,N_9073,N_8163);
xnor U10321 (N_10321,N_8900,N_9950);
nor U10322 (N_10322,N_9807,N_9131);
nor U10323 (N_10323,N_9462,N_8832);
or U10324 (N_10324,N_9319,N_8247);
nand U10325 (N_10325,N_8367,N_9896);
and U10326 (N_10326,N_8096,N_8667);
xor U10327 (N_10327,N_9203,N_9418);
nand U10328 (N_10328,N_9924,N_9837);
xnor U10329 (N_10329,N_9246,N_9784);
or U10330 (N_10330,N_8886,N_8563);
or U10331 (N_10331,N_9226,N_9425);
or U10332 (N_10332,N_9314,N_9582);
nor U10333 (N_10333,N_8458,N_9072);
nand U10334 (N_10334,N_8888,N_9303);
or U10335 (N_10335,N_9782,N_8760);
nand U10336 (N_10336,N_9794,N_8560);
nand U10337 (N_10337,N_8530,N_8409);
and U10338 (N_10338,N_9103,N_9689);
and U10339 (N_10339,N_9697,N_8901);
and U10340 (N_10340,N_9739,N_9529);
xnor U10341 (N_10341,N_9864,N_9382);
and U10342 (N_10342,N_9792,N_9448);
or U10343 (N_10343,N_8066,N_9225);
or U10344 (N_10344,N_8382,N_8006);
nor U10345 (N_10345,N_8492,N_9468);
and U10346 (N_10346,N_8926,N_9334);
or U10347 (N_10347,N_8225,N_8434);
or U10348 (N_10348,N_8645,N_8127);
or U10349 (N_10349,N_9160,N_9642);
nand U10350 (N_10350,N_8448,N_9266);
and U10351 (N_10351,N_8996,N_8311);
nor U10352 (N_10352,N_8983,N_8676);
or U10353 (N_10353,N_9887,N_8180);
or U10354 (N_10354,N_9585,N_9222);
and U10355 (N_10355,N_8109,N_9000);
or U10356 (N_10356,N_9917,N_8270);
or U10357 (N_10357,N_9065,N_8664);
xnor U10358 (N_10358,N_8880,N_9559);
nand U10359 (N_10359,N_8101,N_9829);
nor U10360 (N_10360,N_9040,N_8331);
and U10361 (N_10361,N_9317,N_9150);
xnor U10362 (N_10362,N_9188,N_8075);
nor U10363 (N_10363,N_9871,N_8622);
and U10364 (N_10364,N_8053,N_9614);
nor U10365 (N_10365,N_8694,N_9805);
and U10366 (N_10366,N_8683,N_9877);
nor U10367 (N_10367,N_8209,N_9592);
xor U10368 (N_10368,N_9569,N_8117);
xnor U10369 (N_10369,N_8040,N_8007);
and U10370 (N_10370,N_8997,N_8551);
xor U10371 (N_10371,N_9475,N_9337);
or U10372 (N_10372,N_9137,N_8369);
nor U10373 (N_10373,N_8394,N_8512);
xor U10374 (N_10374,N_8294,N_8227);
or U10375 (N_10375,N_9999,N_8258);
nand U10376 (N_10376,N_8740,N_9035);
or U10377 (N_10377,N_9838,N_8317);
nand U10378 (N_10378,N_8157,N_8059);
nor U10379 (N_10379,N_9421,N_8377);
and U10380 (N_10380,N_9438,N_9544);
and U10381 (N_10381,N_9789,N_9496);
xnor U10382 (N_10382,N_9531,N_9084);
nor U10383 (N_10383,N_8485,N_8031);
and U10384 (N_10384,N_9754,N_9320);
and U10385 (N_10385,N_8771,N_9663);
or U10386 (N_10386,N_8091,N_9604);
xor U10387 (N_10387,N_8572,N_9602);
and U10388 (N_10388,N_9844,N_8220);
xor U10389 (N_10389,N_8845,N_8196);
nand U10390 (N_10390,N_9874,N_8234);
or U10391 (N_10391,N_8457,N_8014);
nor U10392 (N_10392,N_8521,N_9935);
or U10393 (N_10393,N_9473,N_8712);
and U10394 (N_10394,N_9984,N_8640);
or U10395 (N_10395,N_9849,N_8018);
nor U10396 (N_10396,N_8794,N_8769);
or U10397 (N_10397,N_8136,N_9145);
nand U10398 (N_10398,N_8454,N_8873);
nor U10399 (N_10399,N_8634,N_9615);
and U10400 (N_10400,N_9815,N_9034);
nand U10401 (N_10401,N_8187,N_9703);
nand U10402 (N_10402,N_9629,N_8072);
nand U10403 (N_10403,N_8404,N_9576);
nand U10404 (N_10404,N_8972,N_9393);
nor U10405 (N_10405,N_8197,N_8244);
nor U10406 (N_10406,N_8878,N_9392);
nand U10407 (N_10407,N_9283,N_8035);
nor U10408 (N_10408,N_8624,N_8722);
and U10409 (N_10409,N_8252,N_8758);
nand U10410 (N_10410,N_8325,N_9060);
nor U10411 (N_10411,N_8652,N_9361);
nand U10412 (N_10412,N_9547,N_8221);
xor U10413 (N_10413,N_8219,N_9099);
nor U10414 (N_10414,N_9676,N_8488);
nand U10415 (N_10415,N_8135,N_9264);
or U10416 (N_10416,N_9095,N_9485);
nand U10417 (N_10417,N_9812,N_9458);
nand U10418 (N_10418,N_9452,N_8882);
or U10419 (N_10419,N_9389,N_8577);
and U10420 (N_10420,N_9584,N_8668);
or U10421 (N_10421,N_8966,N_9275);
nand U10422 (N_10422,N_8319,N_9031);
nor U10423 (N_10423,N_8553,N_8951);
or U10424 (N_10424,N_8931,N_9096);
and U10425 (N_10425,N_8552,N_8937);
xor U10426 (N_10426,N_8461,N_8399);
nand U10427 (N_10427,N_8954,N_9516);
nor U10428 (N_10428,N_8131,N_8787);
and U10429 (N_10429,N_8437,N_8266);
xnor U10430 (N_10430,N_8172,N_9408);
or U10431 (N_10431,N_9766,N_8463);
nor U10432 (N_10432,N_8686,N_8171);
or U10433 (N_10433,N_9240,N_8238);
nand U10434 (N_10434,N_8780,N_8267);
xor U10435 (N_10435,N_9518,N_8501);
xor U10436 (N_10436,N_9660,N_8125);
and U10437 (N_10437,N_8746,N_8596);
and U10438 (N_10438,N_8050,N_8778);
nand U10439 (N_10439,N_8717,N_8765);
xor U10440 (N_10440,N_9591,N_8555);
nor U10441 (N_10441,N_9939,N_8527);
xor U10442 (N_10442,N_8984,N_9980);
xor U10443 (N_10443,N_8469,N_9436);
and U10444 (N_10444,N_8036,N_9046);
xor U10445 (N_10445,N_8838,N_8566);
or U10446 (N_10446,N_9524,N_8615);
or U10447 (N_10447,N_9381,N_9008);
and U10448 (N_10448,N_8004,N_9181);
and U10449 (N_10449,N_8790,N_9978);
and U10450 (N_10450,N_8818,N_9884);
and U10451 (N_10451,N_8681,N_8576);
nor U10452 (N_10452,N_9045,N_8893);
xnor U10453 (N_10453,N_9130,N_9619);
nor U10454 (N_10454,N_8402,N_9115);
nand U10455 (N_10455,N_8763,N_9565);
nor U10456 (N_10456,N_8981,N_8959);
nor U10457 (N_10457,N_9483,N_9560);
xor U10458 (N_10458,N_8617,N_9118);
or U10459 (N_10459,N_8293,N_9453);
or U10460 (N_10460,N_9843,N_9597);
nand U10461 (N_10461,N_9876,N_8727);
xnor U10462 (N_10462,N_9907,N_8001);
nor U10463 (N_10463,N_9765,N_9056);
and U10464 (N_10464,N_8573,N_9551);
xnor U10465 (N_10465,N_8030,N_8229);
xnor U10466 (N_10466,N_8693,N_8474);
and U10467 (N_10467,N_9025,N_9449);
xnor U10468 (N_10468,N_8741,N_8523);
xnor U10469 (N_10469,N_9112,N_8809);
nand U10470 (N_10470,N_9888,N_9481);
or U10471 (N_10471,N_8806,N_9910);
and U10472 (N_10472,N_9290,N_9616);
or U10473 (N_10473,N_9277,N_8657);
nor U10474 (N_10474,N_8614,N_9129);
nand U10475 (N_10475,N_9416,N_8111);
xor U10476 (N_10476,N_8005,N_9424);
or U10477 (N_10477,N_8974,N_8095);
nor U10478 (N_10478,N_9249,N_9238);
nand U10479 (N_10479,N_8445,N_9043);
xor U10480 (N_10480,N_8941,N_8289);
nor U10481 (N_10481,N_9302,N_9094);
nor U10482 (N_10482,N_9548,N_9932);
nand U10483 (N_10483,N_9028,N_9113);
xnor U10484 (N_10484,N_9326,N_8932);
or U10485 (N_10485,N_9673,N_9097);
xor U10486 (N_10486,N_9398,N_8307);
and U10487 (N_10487,N_9014,N_8390);
nand U10488 (N_10488,N_9300,N_8242);
nand U10489 (N_10489,N_8376,N_8339);
or U10490 (N_10490,N_9528,N_8021);
or U10491 (N_10491,N_9695,N_8616);
or U10492 (N_10492,N_9378,N_9200);
and U10493 (N_10493,N_9175,N_8857);
or U10494 (N_10494,N_8690,N_8971);
and U10495 (N_10495,N_8531,N_8324);
nor U10496 (N_10496,N_8943,N_9402);
nor U10497 (N_10497,N_8859,N_9536);
nor U10498 (N_10498,N_9638,N_8470);
nand U10499 (N_10499,N_9810,N_9786);
or U10500 (N_10500,N_8190,N_9647);
xnor U10501 (N_10501,N_9867,N_9501);
and U10502 (N_10502,N_9367,N_8604);
nand U10503 (N_10503,N_9217,N_9383);
nand U10504 (N_10504,N_9407,N_9598);
nand U10505 (N_10505,N_8923,N_8278);
and U10506 (N_10506,N_8415,N_8032);
and U10507 (N_10507,N_9601,N_9231);
or U10508 (N_10508,N_8265,N_9988);
xnor U10509 (N_10509,N_9059,N_8960);
and U10510 (N_10510,N_9430,N_9800);
nor U10511 (N_10511,N_9806,N_9510);
nor U10512 (N_10512,N_8123,N_9021);
xnor U10513 (N_10513,N_8714,N_8124);
and U10514 (N_10514,N_9540,N_9866);
xor U10515 (N_10515,N_8776,N_9728);
and U10516 (N_10516,N_9711,N_9003);
nand U10517 (N_10517,N_9036,N_8449);
nor U10518 (N_10518,N_8562,N_9301);
nand U10519 (N_10519,N_8071,N_8253);
and U10520 (N_10520,N_8999,N_8950);
xnor U10521 (N_10521,N_9835,N_9679);
nor U10522 (N_10522,N_9737,N_9667);
and U10523 (N_10523,N_8403,N_8116);
nand U10524 (N_10524,N_8508,N_8143);
and U10525 (N_10525,N_8070,N_9833);
or U10526 (N_10526,N_8705,N_9774);
and U10527 (N_10527,N_9215,N_9017);
and U10528 (N_10528,N_9311,N_8141);
nand U10529 (N_10529,N_8010,N_9136);
xor U10530 (N_10530,N_9618,N_8055);
and U10531 (N_10531,N_8612,N_8400);
nor U10532 (N_10532,N_8506,N_9064);
nor U10533 (N_10533,N_8083,N_9466);
nand U10534 (N_10534,N_9834,N_8589);
and U10535 (N_10535,N_9282,N_8605);
xnor U10536 (N_10536,N_8386,N_8743);
nor U10537 (N_10537,N_9440,N_8100);
or U10538 (N_10538,N_8921,N_9773);
nand U10539 (N_10539,N_8643,N_8102);
or U10540 (N_10540,N_9724,N_8277);
nand U10541 (N_10541,N_9895,N_9868);
and U10542 (N_10542,N_8025,N_9955);
nor U10543 (N_10543,N_8368,N_8582);
nand U10544 (N_10544,N_8788,N_8922);
nand U10545 (N_10545,N_8166,N_9865);
and U10546 (N_10546,N_9357,N_8635);
or U10547 (N_10547,N_9854,N_8431);
xnor U10548 (N_10548,N_9813,N_8332);
and U10549 (N_10549,N_8154,N_9221);
or U10550 (N_10550,N_9759,N_9353);
nor U10551 (N_10551,N_8371,N_8453);
xnor U10552 (N_10552,N_8539,N_8013);
xor U10553 (N_10553,N_9818,N_8337);
or U10554 (N_10554,N_8773,N_8505);
or U10555 (N_10555,N_9102,N_9480);
xor U10556 (N_10556,N_9822,N_9934);
nor U10557 (N_10557,N_8419,N_8260);
xor U10558 (N_10558,N_8968,N_9890);
or U10559 (N_10559,N_8731,N_9164);
or U10560 (N_10560,N_9058,N_9826);
or U10561 (N_10561,N_8688,N_8299);
or U10562 (N_10562,N_9327,N_9410);
nand U10563 (N_10563,N_9318,N_9470);
and U10564 (N_10564,N_9832,N_8936);
nand U10565 (N_10565,N_8068,N_8603);
and U10566 (N_10566,N_8233,N_9267);
and U10567 (N_10567,N_8826,N_8421);
nand U10568 (N_10568,N_8940,N_9777);
xnor U10569 (N_10569,N_8535,N_8848);
nor U10570 (N_10570,N_8259,N_9168);
nor U10571 (N_10571,N_9227,N_9599);
nand U10572 (N_10572,N_9666,N_8868);
xor U10573 (N_10573,N_9594,N_9291);
nand U10574 (N_10574,N_8513,N_8816);
and U10575 (N_10575,N_9534,N_9921);
and U10576 (N_10576,N_8628,N_9013);
nand U10577 (N_10577,N_9989,N_9492);
nor U10578 (N_10578,N_8167,N_8847);
nand U10579 (N_10579,N_9790,N_9811);
nand U10580 (N_10580,N_9633,N_9427);
nor U10581 (N_10581,N_9733,N_9561);
xnor U10582 (N_10582,N_9107,N_9690);
nor U10583 (N_10583,N_9253,N_8528);
and U10584 (N_10584,N_9606,N_8482);
nor U10585 (N_10585,N_9881,N_9464);
xnor U10586 (N_10586,N_8480,N_8836);
and U10587 (N_10587,N_8869,N_8587);
nand U10588 (N_10588,N_8581,N_9636);
xnor U10589 (N_10589,N_9681,N_8301);
nor U10590 (N_10590,N_8444,N_8540);
or U10591 (N_10591,N_8750,N_8290);
nand U10592 (N_10592,N_9725,N_8982);
nor U10593 (N_10593,N_8264,N_8819);
and U10594 (N_10594,N_8153,N_8228);
nand U10595 (N_10595,N_9396,N_9049);
nor U10596 (N_10596,N_9985,N_8852);
nand U10597 (N_10597,N_9132,N_9702);
nor U10598 (N_10598,N_9964,N_9729);
xnor U10599 (N_10599,N_9423,N_9259);
nor U10600 (N_10600,N_8500,N_9943);
or U10601 (N_10601,N_9220,N_9682);
xor U10602 (N_10602,N_8846,N_8345);
nor U10603 (N_10603,N_8130,N_8249);
xnor U10604 (N_10604,N_8073,N_8392);
nand U10605 (N_10605,N_8263,N_8944);
xor U10606 (N_10606,N_8775,N_9600);
or U10607 (N_10607,N_8860,N_9469);
or U10608 (N_10608,N_8811,N_9109);
or U10609 (N_10609,N_9742,N_8466);
and U10610 (N_10610,N_9101,N_9523);
nor U10611 (N_10611,N_9643,N_8224);
nor U10612 (N_10612,N_8393,N_8565);
or U10613 (N_10613,N_8907,N_8584);
nor U10614 (N_10614,N_9872,N_8695);
xnor U10615 (N_10615,N_9609,N_9243);
and U10616 (N_10616,N_8894,N_9692);
and U10617 (N_10617,N_9213,N_9344);
or U10618 (N_10618,N_9590,N_8911);
or U10619 (N_10619,N_8162,N_8305);
xor U10620 (N_10620,N_8456,N_9391);
or U10621 (N_10621,N_8351,N_8468);
nor U10622 (N_10622,N_8430,N_9566);
xor U10623 (N_10623,N_8099,N_8522);
or U10624 (N_10624,N_8200,N_8250);
xnor U10625 (N_10625,N_8455,N_9006);
xnor U10626 (N_10626,N_8785,N_8823);
xnor U10627 (N_10627,N_9263,N_8279);
nor U10628 (N_10628,N_8909,N_8580);
and U10629 (N_10629,N_9990,N_8744);
or U10630 (N_10630,N_9875,N_8012);
nor U10631 (N_10631,N_9451,N_9176);
and U10632 (N_10632,N_8719,N_8874);
or U10633 (N_10633,N_9994,N_8207);
xor U10634 (N_10634,N_8844,N_9780);
or U10635 (N_10635,N_9545,N_8828);
nand U10636 (N_10636,N_9761,N_9691);
or U10637 (N_10637,N_8159,N_9646);
xnor U10638 (N_10638,N_8827,N_9125);
and U10639 (N_10639,N_9705,N_8359);
or U10640 (N_10640,N_9187,N_9987);
nand U10641 (N_10641,N_8063,N_9831);
nand U10642 (N_10642,N_9708,N_8550);
nand U10643 (N_10643,N_9349,N_8184);
and U10644 (N_10644,N_8834,N_9192);
or U10645 (N_10645,N_8486,N_8185);
or U10646 (N_10646,N_8044,N_8269);
or U10647 (N_10647,N_8592,N_8805);
nand U10648 (N_10648,N_8076,N_9653);
nand U10649 (N_10649,N_8106,N_8113);
nand U10650 (N_10650,N_9751,N_8665);
and U10651 (N_10651,N_8291,N_9325);
xor U10652 (N_10652,N_9767,N_8496);
and U10653 (N_10653,N_8585,N_9963);
or U10654 (N_10654,N_8915,N_9489);
nor U10655 (N_10655,N_9230,N_8058);
xor U10656 (N_10656,N_9941,N_8821);
nor U10657 (N_10657,N_8752,N_8098);
nand U10658 (N_10658,N_8165,N_9413);
and U10659 (N_10659,N_9641,N_8052);
and U10660 (N_10660,N_8650,N_9915);
and U10661 (N_10661,N_9639,N_9680);
xor U10662 (N_10662,N_9908,N_9900);
nor U10663 (N_10663,N_9185,N_8314);
nand U10664 (N_10664,N_8391,N_8958);
nor U10665 (N_10665,N_8534,N_9194);
nor U10666 (N_10666,N_8452,N_9549);
nand U10667 (N_10667,N_9027,N_9299);
or U10668 (N_10668,N_9795,N_8251);
nor U10669 (N_10669,N_9016,N_9251);
and U10670 (N_10670,N_9323,N_8137);
or U10671 (N_10671,N_8272,N_9648);
xor U10672 (N_10672,N_9435,N_9902);
or U10673 (N_10673,N_9649,N_8193);
nor U10674 (N_10674,N_9892,N_8086);
xor U10675 (N_10675,N_8979,N_8178);
nand U10676 (N_10676,N_8962,N_9541);
nand U10677 (N_10677,N_8786,N_9047);
nor U10678 (N_10678,N_8877,N_8110);
or U10679 (N_10679,N_9414,N_8378);
nor U10680 (N_10680,N_8149,N_9419);
nor U10681 (N_10681,N_8600,N_8364);
nor U10682 (N_10682,N_9484,N_9612);
nand U10683 (N_10683,N_9307,N_9171);
or U10684 (N_10684,N_9262,N_8217);
nand U10685 (N_10685,N_9037,N_9521);
nand U10686 (N_10686,N_8490,N_8908);
and U10687 (N_10687,N_9571,N_9625);
nor U10688 (N_10688,N_9081,N_9234);
nor U10689 (N_10689,N_8427,N_8648);
xnor U10690 (N_10690,N_8961,N_8659);
or U10691 (N_10691,N_9308,N_9514);
or U10692 (N_10692,N_9557,N_8677);
and U10693 (N_10693,N_8179,N_9495);
nand U10694 (N_10694,N_9656,N_9533);
or U10695 (N_10695,N_8644,N_8435);
and U10696 (N_10696,N_9801,N_9289);
xnor U10697 (N_10697,N_8507,N_9443);
or U10698 (N_10698,N_8663,N_9191);
xnor U10699 (N_10699,N_9023,N_9172);
and U10700 (N_10700,N_9029,N_8312);
xnor U10701 (N_10701,N_8257,N_9276);
nor U10702 (N_10702,N_8638,N_9873);
xnor U10703 (N_10703,N_8236,N_9889);
nor U10704 (N_10704,N_9288,N_8093);
nor U10705 (N_10705,N_8282,N_8065);
and U10706 (N_10706,N_8475,N_9961);
nand U10707 (N_10707,N_9515,N_9009);
and U10708 (N_10708,N_8801,N_9821);
nor U10709 (N_10709,N_9952,N_9683);
or U10710 (N_10710,N_8155,N_8557);
or U10711 (N_10711,N_8107,N_8425);
xnor U10712 (N_10712,N_9406,N_9578);
nor U10713 (N_10713,N_9752,N_9360);
or U10714 (N_10714,N_9852,N_9909);
nor U10715 (N_10715,N_9661,N_8625);
xnor U10716 (N_10716,N_8955,N_9574);
xor U10717 (N_10717,N_8547,N_8498);
and U10718 (N_10718,N_8146,N_8904);
nor U10719 (N_10719,N_8989,N_8097);
and U10720 (N_10720,N_8208,N_8405);
and U10721 (N_10721,N_8049,N_9498);
or U10722 (N_10722,N_8088,N_8807);
xor U10723 (N_10723,N_9241,N_8396);
xor U10724 (N_10724,N_9012,N_9563);
nand U10725 (N_10725,N_9509,N_9727);
nand U10726 (N_10726,N_9842,N_8121);
nor U10727 (N_10727,N_9211,N_9429);
nand U10728 (N_10728,N_8918,N_8363);
nand U10729 (N_10729,N_8567,N_8479);
and U10730 (N_10730,N_9788,N_9324);
or U10731 (N_10731,N_9699,N_9918);
xor U10732 (N_10732,N_9796,N_9071);
and U10733 (N_10733,N_9685,N_9224);
nand U10734 (N_10734,N_9651,N_9461);
and U10735 (N_10735,N_8296,N_9078);
xnor U10736 (N_10736,N_8610,N_8602);
and U10737 (N_10737,N_9169,N_9022);
nand U10738 (N_10738,N_8347,N_9605);
nand U10739 (N_10739,N_9783,N_8728);
nor U10740 (N_10740,N_8128,N_9294);
nand U10741 (N_10741,N_8483,N_8240);
or U10742 (N_10742,N_9762,N_8543);
or U10743 (N_10743,N_8885,N_8680);
and U10744 (N_10744,N_8422,N_8494);
xor U10745 (N_10745,N_8591,N_8753);
xnor U10746 (N_10746,N_8703,N_9355);
or U10747 (N_10747,N_8395,N_9486);
and U10748 (N_10748,N_9441,N_9247);
nor U10749 (N_10749,N_9310,N_8152);
and U10750 (N_10750,N_8275,N_9100);
nor U10751 (N_10751,N_8212,N_9177);
nand U10752 (N_10752,N_8280,N_8532);
nand U10753 (N_10753,N_9155,N_9937);
xnor U10754 (N_10754,N_9827,N_9968);
nor U10755 (N_10755,N_9734,N_9986);
and U10756 (N_10756,N_9511,N_8970);
xor U10757 (N_10757,N_9817,N_9845);
nand U10758 (N_10758,N_9922,N_8510);
and U10759 (N_10759,N_9329,N_8366);
nor U10760 (N_10760,N_9863,N_8935);
xor U10761 (N_10761,N_9982,N_8158);
nor U10762 (N_10762,N_9714,N_9830);
nand U10763 (N_10763,N_8081,N_9401);
or U10764 (N_10764,N_8564,N_8365);
or U10765 (N_10765,N_8992,N_9278);
or U10766 (N_10766,N_9668,N_8156);
nor U10767 (N_10767,N_8526,N_8194);
xor U10768 (N_10768,N_8671,N_9672);
xor U10769 (N_10769,N_9202,N_8820);
nand U10770 (N_10770,N_9456,N_8687);
nand U10771 (N_10771,N_8558,N_8372);
nor U10772 (N_10772,N_9001,N_8561);
or U10773 (N_10773,N_9270,N_8542);
nand U10774 (N_10774,N_9292,N_9494);
xor U10775 (N_10775,N_8745,N_9610);
xnor U10776 (N_10776,N_9245,N_8782);
xnor U10777 (N_10777,N_9956,N_9738);
xor U10778 (N_10778,N_8571,N_9375);
and U10779 (N_10779,N_8761,N_8777);
nand U10780 (N_10780,N_9772,N_9696);
and U10781 (N_10781,N_8245,N_9542);
nor U10782 (N_10782,N_8599,N_8779);
nor U10783 (N_10783,N_9972,N_9151);
nand U10784 (N_10784,N_8423,N_8928);
or U10785 (N_10785,N_8570,N_9816);
xor U10786 (N_10786,N_9923,N_9124);
or U10787 (N_10787,N_9859,N_8398);
nor U10788 (N_10788,N_8019,N_8755);
nor U10789 (N_10789,N_9716,N_9757);
xor U10790 (N_10790,N_8953,N_9123);
nand U10791 (N_10791,N_9965,N_9898);
and U10792 (N_10792,N_9799,N_8789);
or U10793 (N_10793,N_9583,N_9347);
and U10794 (N_10794,N_9182,N_9146);
xnor U10795 (N_10795,N_8598,N_9654);
or U10796 (N_10796,N_9228,N_8721);
xor U10797 (N_10797,N_8685,N_9861);
nor U10798 (N_10798,N_8138,N_8754);
nor U10799 (N_10799,N_8323,N_9376);
xor U10800 (N_10800,N_9280,N_9358);
xnor U10801 (N_10801,N_9236,N_9975);
nand U10802 (N_10802,N_9546,N_8618);
xor U10803 (N_10803,N_8892,N_9252);
xnor U10804 (N_10804,N_8329,N_8330);
xor U10805 (N_10805,N_9537,N_9721);
or U10806 (N_10806,N_8734,N_9405);
nand U10807 (N_10807,N_9373,N_9399);
and U10808 (N_10808,N_9522,N_8516);
or U10809 (N_10809,N_8875,N_9929);
nand U10810 (N_10810,N_8830,N_8262);
xor U10811 (N_10811,N_9951,N_9913);
nor U10812 (N_10812,N_8387,N_9698);
xor U10813 (N_10813,N_9482,N_8061);
or U10814 (N_10814,N_8089,N_8853);
nor U10815 (N_10815,N_9880,N_8118);
nor U10816 (N_10816,N_9665,N_9209);
and U10817 (N_10817,N_9122,N_9068);
nor U10818 (N_10818,N_8002,N_8140);
xnor U10819 (N_10819,N_8626,N_8491);
nand U10820 (N_10820,N_9850,N_9715);
and U10821 (N_10821,N_8210,N_9802);
nor U10822 (N_10822,N_8759,N_8205);
or U10823 (N_10823,N_9265,N_8349);
and U10824 (N_10824,N_9785,N_8590);
nor U10825 (N_10825,N_9178,N_8976);
nor U10826 (N_10826,N_8261,N_8730);
nand U10827 (N_10827,N_9157,N_8034);
nand U10828 (N_10828,N_9992,N_9098);
and U10829 (N_10829,N_8871,N_8917);
xor U10830 (N_10830,N_9051,N_8237);
or U10831 (N_10831,N_8176,N_9870);
nand U10832 (N_10832,N_9116,N_9156);
xor U10833 (N_10833,N_9437,N_8674);
xor U10834 (N_10834,N_8230,N_8046);
or U10835 (N_10835,N_9631,N_8841);
nand U10836 (N_10836,N_9513,N_8947);
xnor U10837 (N_10837,N_9556,N_9550);
xnor U10838 (N_10838,N_9139,N_8715);
nand U10839 (N_10839,N_8315,N_9809);
nand U10840 (N_10840,N_9432,N_9370);
and U10841 (N_10841,N_9862,N_9256);
or U10842 (N_10842,N_8321,N_9779);
and U10843 (N_10843,N_9298,N_9332);
nand U10844 (N_10844,N_9170,N_8556);
nor U10845 (N_10845,N_9196,N_8008);
xor U10846 (N_10846,N_9539,N_9083);
and U10847 (N_10847,N_9487,N_8929);
nor U10848 (N_10848,N_9374,N_9149);
xnor U10849 (N_10849,N_8487,N_8767);
or U10850 (N_10850,N_9134,N_9077);
and U10851 (N_10851,N_9261,N_9611);
or U10852 (N_10852,N_9431,N_8920);
nor U10853 (N_10853,N_9147,N_8276);
or U10854 (N_10854,N_8840,N_8948);
nand U10855 (N_10855,N_9966,N_9379);
or U10856 (N_10856,N_8939,N_8701);
and U10857 (N_10857,N_9459,N_9575);
and U10858 (N_10858,N_9581,N_9793);
or U10859 (N_10859,N_9363,N_9445);
xor U10860 (N_10860,N_9634,N_9554);
or U10861 (N_10861,N_8041,N_8060);
nand U10862 (N_10862,N_8334,N_8383);
nor U10863 (N_10863,N_8168,N_8544);
and U10864 (N_10864,N_9315,N_8133);
nand U10865 (N_10865,N_9455,N_9390);
nand U10866 (N_10866,N_9365,N_9981);
nor U10867 (N_10867,N_8362,N_8902);
nor U10868 (N_10868,N_9755,N_9039);
nand U10869 (N_10869,N_8285,N_9630);
xnor U10870 (N_10870,N_9210,N_9386);
nor U10871 (N_10871,N_9538,N_8348);
or U10872 (N_10872,N_8033,N_8484);
nand U10873 (N_10873,N_8039,N_9309);
or U10874 (N_10874,N_8793,N_8524);
nor U10875 (N_10875,N_9313,N_9257);
or U10876 (N_10876,N_8723,N_8864);
or U10877 (N_10877,N_9626,N_8831);
and U10878 (N_10878,N_8720,N_9206);
nand U10879 (N_10879,N_8092,N_8742);
and U10880 (N_10880,N_9335,N_9520);
or U10881 (N_10881,N_9798,N_9368);
and U10882 (N_10882,N_9904,N_9467);
or U10883 (N_10883,N_9579,N_8945);
and U10884 (N_10884,N_9684,N_9038);
and U10885 (N_10885,N_8450,N_8995);
nor U10886 (N_10886,N_9617,N_9161);
nand U10887 (N_10887,N_8191,N_9144);
nor U10888 (N_10888,N_8679,N_8401);
or U10889 (N_10889,N_9218,N_9340);
nor U10890 (N_10890,N_8181,N_8064);
nand U10891 (N_10891,N_8833,N_9640);
nor U10892 (N_10892,N_8080,N_9825);
xnor U10893 (N_10893,N_9422,N_9957);
nor U10894 (N_10894,N_8246,N_8056);
nor U10895 (N_10895,N_9403,N_9152);
nand U10896 (N_10896,N_8283,N_9507);
and U10897 (N_10897,N_8641,N_8899);
nor U10898 (N_10898,N_9967,N_9808);
or U10899 (N_10899,N_9388,N_8629);
or U10900 (N_10900,N_9163,N_9128);
nand U10901 (N_10901,N_8738,N_8669);
xor U10902 (N_10902,N_9345,N_9497);
or U10903 (N_10903,N_9650,N_9848);
xnor U10904 (N_10904,N_9535,N_8489);
xor U10905 (N_10905,N_9958,N_9010);
or U10906 (N_10906,N_8271,N_9894);
or U10907 (N_10907,N_8003,N_9055);
xnor U10908 (N_10908,N_8630,N_8443);
or U10909 (N_10909,N_8575,N_8292);
or U10910 (N_10910,N_9903,N_9893);
nor U10911 (N_10911,N_8203,N_8335);
nand U10912 (N_10912,N_8350,N_9853);
or U10913 (N_10913,N_8112,N_8336);
and U10914 (N_10914,N_8045,N_9891);
nor U10915 (N_10915,N_8206,N_9471);
nand U10916 (N_10916,N_8839,N_9709);
xor U10917 (N_10917,N_8986,N_8910);
nor U10918 (N_10918,N_8388,N_9117);
or U10919 (N_10919,N_9804,N_8198);
nand U10920 (N_10920,N_8851,N_9771);
nand U10921 (N_10921,N_9173,N_9911);
xor U10922 (N_10922,N_8843,N_9079);
and U10923 (N_10923,N_9490,N_9133);
and U10924 (N_10924,N_8511,N_8322);
xor U10925 (N_10925,N_9354,N_8764);
nor U10926 (N_10926,N_8993,N_8462);
nor U10927 (N_10927,N_9628,N_8914);
nand U10928 (N_10928,N_9087,N_8370);
or U10929 (N_10929,N_9143,N_8850);
xor U10930 (N_10930,N_9242,N_8384);
or U10931 (N_10931,N_8751,N_8389);
xor U10932 (N_10932,N_8354,N_8653);
nand U10933 (N_10933,N_9180,N_8985);
or U10934 (N_10934,N_9564,N_8438);
nor U10935 (N_10935,N_8842,N_8160);
xor U10936 (N_10936,N_8174,N_8729);
nor U10937 (N_10937,N_8000,N_9371);
xor U10938 (N_10938,N_8424,N_9670);
nor U10939 (N_10939,N_9201,N_9707);
xor U10940 (N_10940,N_8870,N_9285);
and U10941 (N_10941,N_8464,N_8781);
nand U10942 (N_10942,N_8891,N_9091);
nor U10943 (N_10943,N_8223,N_8478);
and U10944 (N_10944,N_9341,N_8481);
or U10945 (N_10945,N_9159,N_8814);
and U10946 (N_10946,N_9235,N_9906);
xor U10947 (N_10947,N_8303,N_8621);
nand U10948 (N_10948,N_8273,N_9154);
and U10949 (N_10949,N_8541,N_8023);
nand U10950 (N_10950,N_9446,N_8678);
nor U10951 (N_10951,N_8361,N_8661);
or U10952 (N_10952,N_8656,N_9205);
nor U10953 (N_10953,N_9840,N_9426);
nor U10954 (N_10954,N_9417,N_8385);
nand U10955 (N_10955,N_8770,N_8211);
or U10956 (N_10956,N_9505,N_9983);
or U10957 (N_10957,N_9093,N_9500);
xor U10958 (N_10958,N_9726,N_9088);
or U10959 (N_10959,N_8281,N_9158);
nand U10960 (N_10960,N_8122,N_8707);
nand U10961 (N_10961,N_8702,N_8735);
and U10962 (N_10962,N_8504,N_9700);
xnor U10963 (N_10963,N_8987,N_9069);
nand U10964 (N_10964,N_8173,N_9212);
and U10965 (N_10965,N_9901,N_8538);
nor U10966 (N_10966,N_9183,N_9162);
xnor U10967 (N_10967,N_8054,N_8791);
or U10968 (N_10968,N_8813,N_8569);
nand U10969 (N_10969,N_8214,N_9769);
and U10970 (N_10970,N_9747,N_8804);
xor U10971 (N_10971,N_8632,N_8432);
and U10972 (N_10972,N_8660,N_8949);
nand U10973 (N_10973,N_8473,N_8082);
xor U10974 (N_10974,N_9121,N_8815);
or U10975 (N_10975,N_9580,N_8300);
nand U10976 (N_10976,N_8447,N_8691);
nand U10977 (N_10977,N_9570,N_8651);
or U10978 (N_10978,N_9693,N_9250);
and U10979 (N_10979,N_9336,N_9463);
and U10980 (N_10980,N_8574,N_9330);
nand U10981 (N_10981,N_9293,N_9627);
nand U10982 (N_10982,N_9532,N_9621);
and U10983 (N_10983,N_9258,N_8502);
nor U10984 (N_10984,N_8027,N_9712);
xor U10985 (N_10985,N_8548,N_9054);
nand U10986 (N_10986,N_8327,N_8934);
and U10987 (N_10987,N_8525,N_9024);
xor U10988 (N_10988,N_8414,N_9153);
and U10989 (N_10989,N_9364,N_8649);
or U10990 (N_10990,N_9409,N_9858);
or U10991 (N_10991,N_9041,N_9119);
nand U10992 (N_10992,N_9512,N_8346);
xnor U10993 (N_10993,N_9562,N_8239);
xor U10994 (N_10994,N_9237,N_8662);
nor U10995 (N_10995,N_9572,N_9704);
or U10996 (N_10996,N_9011,N_9343);
xor U10997 (N_10997,N_9744,N_9331);
nor U10998 (N_10998,N_8799,N_9140);
and U10999 (N_10999,N_8988,N_9216);
or U11000 (N_11000,N_9366,N_8856);
nor U11001 (N_11001,N_8856,N_8757);
or U11002 (N_11002,N_9055,N_9747);
xnor U11003 (N_11003,N_8156,N_9784);
and U11004 (N_11004,N_8640,N_9212);
nand U11005 (N_11005,N_8399,N_9490);
or U11006 (N_11006,N_9589,N_8131);
nand U11007 (N_11007,N_9084,N_9383);
xnor U11008 (N_11008,N_9249,N_8588);
nand U11009 (N_11009,N_8569,N_8673);
and U11010 (N_11010,N_8465,N_9306);
xnor U11011 (N_11011,N_9023,N_9197);
and U11012 (N_11012,N_8618,N_9793);
nor U11013 (N_11013,N_9851,N_8460);
and U11014 (N_11014,N_9460,N_8539);
xnor U11015 (N_11015,N_8859,N_8084);
and U11016 (N_11016,N_8379,N_8874);
or U11017 (N_11017,N_8571,N_8217);
xor U11018 (N_11018,N_9631,N_8802);
nor U11019 (N_11019,N_9638,N_8243);
xor U11020 (N_11020,N_8278,N_9510);
and U11021 (N_11021,N_9939,N_9533);
or U11022 (N_11022,N_9469,N_9194);
nor U11023 (N_11023,N_8337,N_8574);
or U11024 (N_11024,N_8732,N_9948);
and U11025 (N_11025,N_8316,N_9002);
and U11026 (N_11026,N_9016,N_9538);
or U11027 (N_11027,N_9997,N_8825);
nand U11028 (N_11028,N_9220,N_8428);
xnor U11029 (N_11029,N_9088,N_9552);
nand U11030 (N_11030,N_9368,N_9727);
xor U11031 (N_11031,N_8991,N_9393);
nand U11032 (N_11032,N_8300,N_8849);
and U11033 (N_11033,N_8717,N_9840);
xor U11034 (N_11034,N_9465,N_8462);
nand U11035 (N_11035,N_8316,N_8684);
and U11036 (N_11036,N_8306,N_9648);
nor U11037 (N_11037,N_8353,N_8989);
nor U11038 (N_11038,N_8743,N_9079);
or U11039 (N_11039,N_8787,N_8611);
xnor U11040 (N_11040,N_9084,N_8872);
nand U11041 (N_11041,N_9389,N_8742);
xnor U11042 (N_11042,N_9084,N_9967);
xor U11043 (N_11043,N_9645,N_9298);
or U11044 (N_11044,N_8106,N_9557);
and U11045 (N_11045,N_8967,N_8939);
or U11046 (N_11046,N_9748,N_9171);
or U11047 (N_11047,N_9711,N_8850);
nor U11048 (N_11048,N_9170,N_9202);
nand U11049 (N_11049,N_9559,N_8987);
nand U11050 (N_11050,N_9674,N_8399);
or U11051 (N_11051,N_9881,N_8953);
xnor U11052 (N_11052,N_8793,N_8238);
xnor U11053 (N_11053,N_9110,N_8133);
xor U11054 (N_11054,N_9090,N_8706);
xor U11055 (N_11055,N_8484,N_9360);
xnor U11056 (N_11056,N_8984,N_9789);
nor U11057 (N_11057,N_9150,N_8840);
and U11058 (N_11058,N_9479,N_8232);
nor U11059 (N_11059,N_9740,N_9276);
xnor U11060 (N_11060,N_8987,N_9263);
nor U11061 (N_11061,N_8388,N_8435);
xor U11062 (N_11062,N_9726,N_8640);
or U11063 (N_11063,N_8224,N_8030);
nor U11064 (N_11064,N_9182,N_9206);
nor U11065 (N_11065,N_8903,N_8362);
or U11066 (N_11066,N_8103,N_9744);
nand U11067 (N_11067,N_8651,N_8206);
xnor U11068 (N_11068,N_8865,N_8213);
xnor U11069 (N_11069,N_8415,N_8849);
nor U11070 (N_11070,N_8100,N_8400);
xor U11071 (N_11071,N_9817,N_8439);
nand U11072 (N_11072,N_9588,N_9759);
or U11073 (N_11073,N_8944,N_9746);
and U11074 (N_11074,N_9523,N_8097);
xor U11075 (N_11075,N_8274,N_8471);
nand U11076 (N_11076,N_8292,N_9322);
nor U11077 (N_11077,N_9499,N_8005);
xnor U11078 (N_11078,N_9993,N_9140);
and U11079 (N_11079,N_9506,N_9708);
nand U11080 (N_11080,N_8856,N_9433);
or U11081 (N_11081,N_8709,N_8054);
and U11082 (N_11082,N_9321,N_9288);
or U11083 (N_11083,N_9272,N_9139);
or U11084 (N_11084,N_9099,N_8147);
and U11085 (N_11085,N_8553,N_8390);
nor U11086 (N_11086,N_8760,N_8003);
or U11087 (N_11087,N_8904,N_8337);
nor U11088 (N_11088,N_8397,N_8529);
xor U11089 (N_11089,N_8588,N_8528);
or U11090 (N_11090,N_8874,N_8356);
xnor U11091 (N_11091,N_8869,N_9596);
and U11092 (N_11092,N_8342,N_9140);
nor U11093 (N_11093,N_9389,N_9626);
xnor U11094 (N_11094,N_8690,N_8844);
xor U11095 (N_11095,N_8683,N_8704);
or U11096 (N_11096,N_9953,N_9359);
nand U11097 (N_11097,N_8343,N_9488);
nand U11098 (N_11098,N_8001,N_9882);
nand U11099 (N_11099,N_9235,N_9405);
or U11100 (N_11100,N_9704,N_8522);
nand U11101 (N_11101,N_9769,N_8314);
nand U11102 (N_11102,N_9417,N_8952);
nor U11103 (N_11103,N_8841,N_9376);
nor U11104 (N_11104,N_9923,N_9772);
nand U11105 (N_11105,N_8246,N_9989);
nand U11106 (N_11106,N_9991,N_8712);
nor U11107 (N_11107,N_9697,N_8965);
nand U11108 (N_11108,N_8839,N_8128);
xnor U11109 (N_11109,N_8032,N_8236);
nor U11110 (N_11110,N_8730,N_8481);
xor U11111 (N_11111,N_9369,N_8842);
and U11112 (N_11112,N_9371,N_8721);
and U11113 (N_11113,N_8377,N_8466);
or U11114 (N_11114,N_9469,N_8756);
nand U11115 (N_11115,N_8647,N_8103);
nor U11116 (N_11116,N_8930,N_8989);
xor U11117 (N_11117,N_8984,N_8166);
or U11118 (N_11118,N_9889,N_8649);
nand U11119 (N_11119,N_9551,N_8206);
xnor U11120 (N_11120,N_9096,N_8887);
or U11121 (N_11121,N_8391,N_8393);
xnor U11122 (N_11122,N_8752,N_9427);
and U11123 (N_11123,N_8160,N_9659);
or U11124 (N_11124,N_8315,N_8466);
nor U11125 (N_11125,N_8928,N_8675);
xor U11126 (N_11126,N_8969,N_9140);
nor U11127 (N_11127,N_9940,N_8282);
nor U11128 (N_11128,N_8173,N_9841);
xnor U11129 (N_11129,N_9781,N_8327);
or U11130 (N_11130,N_8851,N_8815);
xor U11131 (N_11131,N_9574,N_9287);
nand U11132 (N_11132,N_8895,N_9754);
and U11133 (N_11133,N_9424,N_9264);
and U11134 (N_11134,N_9834,N_8270);
xor U11135 (N_11135,N_9669,N_8842);
nand U11136 (N_11136,N_8468,N_8710);
nand U11137 (N_11137,N_9993,N_8234);
nor U11138 (N_11138,N_8937,N_9948);
nand U11139 (N_11139,N_9026,N_8237);
nor U11140 (N_11140,N_8371,N_8737);
nand U11141 (N_11141,N_9824,N_9915);
xnor U11142 (N_11142,N_8289,N_9531);
and U11143 (N_11143,N_8000,N_8214);
nand U11144 (N_11144,N_8341,N_9724);
and U11145 (N_11145,N_9436,N_8005);
or U11146 (N_11146,N_8515,N_9379);
and U11147 (N_11147,N_8074,N_9344);
or U11148 (N_11148,N_9547,N_8451);
or U11149 (N_11149,N_9619,N_9364);
nor U11150 (N_11150,N_8576,N_9674);
nor U11151 (N_11151,N_8391,N_8969);
xor U11152 (N_11152,N_9436,N_9271);
nand U11153 (N_11153,N_9249,N_9074);
or U11154 (N_11154,N_9315,N_8095);
nand U11155 (N_11155,N_9312,N_8482);
xor U11156 (N_11156,N_8137,N_9337);
and U11157 (N_11157,N_8828,N_9996);
and U11158 (N_11158,N_9994,N_8187);
nor U11159 (N_11159,N_9078,N_8411);
xnor U11160 (N_11160,N_9590,N_9024);
nand U11161 (N_11161,N_9721,N_8536);
xor U11162 (N_11162,N_8646,N_9784);
nand U11163 (N_11163,N_9988,N_8854);
or U11164 (N_11164,N_8398,N_8619);
nor U11165 (N_11165,N_8123,N_8594);
and U11166 (N_11166,N_8992,N_9435);
or U11167 (N_11167,N_9891,N_9247);
nand U11168 (N_11168,N_9979,N_9147);
nand U11169 (N_11169,N_8732,N_9023);
nor U11170 (N_11170,N_9685,N_9687);
and U11171 (N_11171,N_9565,N_9612);
or U11172 (N_11172,N_9994,N_8573);
and U11173 (N_11173,N_8898,N_8883);
or U11174 (N_11174,N_8942,N_8593);
xnor U11175 (N_11175,N_8542,N_9842);
and U11176 (N_11176,N_9282,N_8786);
or U11177 (N_11177,N_9138,N_9808);
nand U11178 (N_11178,N_8702,N_8990);
xor U11179 (N_11179,N_9155,N_8957);
nand U11180 (N_11180,N_9503,N_8209);
nor U11181 (N_11181,N_9430,N_9813);
nor U11182 (N_11182,N_8793,N_8967);
xnor U11183 (N_11183,N_9372,N_8038);
and U11184 (N_11184,N_8667,N_8748);
nor U11185 (N_11185,N_8815,N_8985);
xnor U11186 (N_11186,N_9117,N_9154);
nor U11187 (N_11187,N_9805,N_8373);
and U11188 (N_11188,N_9798,N_8217);
xor U11189 (N_11189,N_9459,N_9738);
nand U11190 (N_11190,N_9512,N_8659);
xnor U11191 (N_11191,N_9367,N_9308);
or U11192 (N_11192,N_9130,N_8907);
nand U11193 (N_11193,N_9920,N_8583);
and U11194 (N_11194,N_8600,N_9237);
nand U11195 (N_11195,N_8543,N_8482);
nand U11196 (N_11196,N_9454,N_8743);
or U11197 (N_11197,N_9706,N_9316);
or U11198 (N_11198,N_8246,N_8973);
nand U11199 (N_11199,N_8395,N_8675);
nor U11200 (N_11200,N_8813,N_8704);
and U11201 (N_11201,N_9238,N_9710);
nor U11202 (N_11202,N_9867,N_9391);
xor U11203 (N_11203,N_9373,N_9784);
and U11204 (N_11204,N_9395,N_9271);
xor U11205 (N_11205,N_9758,N_9086);
nand U11206 (N_11206,N_9920,N_9638);
and U11207 (N_11207,N_8139,N_8217);
or U11208 (N_11208,N_9198,N_8693);
nand U11209 (N_11209,N_8711,N_8212);
nor U11210 (N_11210,N_8473,N_8003);
xor U11211 (N_11211,N_9353,N_9913);
xnor U11212 (N_11212,N_9551,N_9868);
or U11213 (N_11213,N_8418,N_8047);
and U11214 (N_11214,N_9343,N_9468);
or U11215 (N_11215,N_8866,N_9926);
and U11216 (N_11216,N_8204,N_9111);
xnor U11217 (N_11217,N_9822,N_9379);
nand U11218 (N_11218,N_9891,N_8157);
nand U11219 (N_11219,N_9559,N_9050);
nor U11220 (N_11220,N_8497,N_8792);
nand U11221 (N_11221,N_8693,N_8692);
or U11222 (N_11222,N_9104,N_8724);
xor U11223 (N_11223,N_9198,N_9106);
nand U11224 (N_11224,N_9668,N_8726);
nor U11225 (N_11225,N_8212,N_9178);
xnor U11226 (N_11226,N_8652,N_9616);
nand U11227 (N_11227,N_8559,N_8572);
nor U11228 (N_11228,N_9193,N_8742);
or U11229 (N_11229,N_8867,N_8500);
or U11230 (N_11230,N_9168,N_8206);
nand U11231 (N_11231,N_8468,N_8486);
xnor U11232 (N_11232,N_9393,N_9907);
xor U11233 (N_11233,N_8499,N_9398);
nand U11234 (N_11234,N_8325,N_8006);
and U11235 (N_11235,N_8556,N_8925);
and U11236 (N_11236,N_8981,N_8028);
and U11237 (N_11237,N_9701,N_9854);
nor U11238 (N_11238,N_9839,N_8962);
xnor U11239 (N_11239,N_8430,N_9202);
xnor U11240 (N_11240,N_8492,N_9692);
nor U11241 (N_11241,N_8854,N_8545);
nor U11242 (N_11242,N_8788,N_9574);
nor U11243 (N_11243,N_9353,N_8419);
nand U11244 (N_11244,N_9594,N_9399);
and U11245 (N_11245,N_9806,N_9615);
and U11246 (N_11246,N_9846,N_9800);
xor U11247 (N_11247,N_8266,N_9946);
nor U11248 (N_11248,N_9101,N_8570);
or U11249 (N_11249,N_8145,N_8851);
xor U11250 (N_11250,N_8093,N_8163);
xor U11251 (N_11251,N_9839,N_9725);
and U11252 (N_11252,N_9556,N_8029);
or U11253 (N_11253,N_9646,N_9039);
nand U11254 (N_11254,N_8117,N_8518);
xor U11255 (N_11255,N_9560,N_8116);
and U11256 (N_11256,N_9975,N_9274);
nand U11257 (N_11257,N_9869,N_9968);
or U11258 (N_11258,N_8151,N_9572);
nand U11259 (N_11259,N_9100,N_9452);
nor U11260 (N_11260,N_9573,N_8943);
and U11261 (N_11261,N_9382,N_8954);
nor U11262 (N_11262,N_8302,N_8027);
nand U11263 (N_11263,N_9077,N_8027);
nor U11264 (N_11264,N_9658,N_9282);
nor U11265 (N_11265,N_9391,N_8534);
or U11266 (N_11266,N_8730,N_9104);
xnor U11267 (N_11267,N_9423,N_9080);
xor U11268 (N_11268,N_9716,N_8104);
or U11269 (N_11269,N_9565,N_8021);
xor U11270 (N_11270,N_8830,N_9057);
xnor U11271 (N_11271,N_8047,N_8011);
nand U11272 (N_11272,N_8584,N_9620);
nor U11273 (N_11273,N_9602,N_8200);
nor U11274 (N_11274,N_8444,N_8621);
or U11275 (N_11275,N_8177,N_8536);
nand U11276 (N_11276,N_9860,N_9363);
and U11277 (N_11277,N_9321,N_9614);
and U11278 (N_11278,N_8206,N_8213);
or U11279 (N_11279,N_8151,N_8572);
or U11280 (N_11280,N_9489,N_8268);
xnor U11281 (N_11281,N_9775,N_9512);
xor U11282 (N_11282,N_9472,N_9158);
or U11283 (N_11283,N_8813,N_9293);
or U11284 (N_11284,N_9994,N_9689);
xnor U11285 (N_11285,N_8257,N_8394);
nor U11286 (N_11286,N_8136,N_8119);
xnor U11287 (N_11287,N_8221,N_9027);
nand U11288 (N_11288,N_9810,N_9323);
and U11289 (N_11289,N_9191,N_9981);
nor U11290 (N_11290,N_9134,N_9571);
or U11291 (N_11291,N_9307,N_8748);
or U11292 (N_11292,N_8822,N_8361);
nand U11293 (N_11293,N_9844,N_9885);
xor U11294 (N_11294,N_8496,N_8351);
and U11295 (N_11295,N_9863,N_8779);
or U11296 (N_11296,N_9268,N_9284);
xnor U11297 (N_11297,N_8232,N_8252);
nor U11298 (N_11298,N_9207,N_9014);
xnor U11299 (N_11299,N_8855,N_8232);
nor U11300 (N_11300,N_9588,N_8818);
nand U11301 (N_11301,N_8486,N_9725);
nor U11302 (N_11302,N_8736,N_9224);
or U11303 (N_11303,N_9482,N_9801);
xor U11304 (N_11304,N_8203,N_8640);
or U11305 (N_11305,N_9149,N_9938);
nor U11306 (N_11306,N_9434,N_9609);
nor U11307 (N_11307,N_9668,N_8097);
and U11308 (N_11308,N_8548,N_9044);
nand U11309 (N_11309,N_9807,N_8482);
or U11310 (N_11310,N_8331,N_9739);
nor U11311 (N_11311,N_9123,N_9665);
and U11312 (N_11312,N_8337,N_9774);
and U11313 (N_11313,N_8098,N_8785);
and U11314 (N_11314,N_9456,N_8082);
and U11315 (N_11315,N_8977,N_9370);
nand U11316 (N_11316,N_8409,N_8844);
nand U11317 (N_11317,N_9176,N_9141);
nor U11318 (N_11318,N_9184,N_9830);
and U11319 (N_11319,N_8724,N_8328);
or U11320 (N_11320,N_9921,N_9813);
and U11321 (N_11321,N_8925,N_8630);
nand U11322 (N_11322,N_9963,N_9711);
or U11323 (N_11323,N_9198,N_9367);
nor U11324 (N_11324,N_8568,N_8220);
xor U11325 (N_11325,N_9933,N_9679);
or U11326 (N_11326,N_9205,N_8699);
nor U11327 (N_11327,N_9228,N_9337);
nand U11328 (N_11328,N_8353,N_9356);
and U11329 (N_11329,N_8812,N_9073);
and U11330 (N_11330,N_9390,N_8963);
and U11331 (N_11331,N_9657,N_8298);
nand U11332 (N_11332,N_8575,N_9560);
or U11333 (N_11333,N_9086,N_8598);
xor U11334 (N_11334,N_9625,N_8602);
and U11335 (N_11335,N_8647,N_8859);
and U11336 (N_11336,N_9581,N_9321);
and U11337 (N_11337,N_9923,N_9838);
and U11338 (N_11338,N_8906,N_8640);
xnor U11339 (N_11339,N_9411,N_8020);
nand U11340 (N_11340,N_9624,N_8086);
nand U11341 (N_11341,N_9146,N_8163);
or U11342 (N_11342,N_8907,N_8990);
xor U11343 (N_11343,N_8847,N_8748);
nor U11344 (N_11344,N_8885,N_8109);
xor U11345 (N_11345,N_8558,N_8447);
xnor U11346 (N_11346,N_9733,N_8060);
nor U11347 (N_11347,N_8050,N_9448);
nor U11348 (N_11348,N_8416,N_9663);
and U11349 (N_11349,N_8827,N_9472);
nand U11350 (N_11350,N_9595,N_8295);
xor U11351 (N_11351,N_9763,N_8451);
nor U11352 (N_11352,N_8648,N_9116);
xnor U11353 (N_11353,N_9941,N_9554);
nor U11354 (N_11354,N_9080,N_8344);
or U11355 (N_11355,N_9167,N_9040);
xnor U11356 (N_11356,N_9105,N_9381);
xor U11357 (N_11357,N_8930,N_9040);
or U11358 (N_11358,N_8683,N_8655);
nor U11359 (N_11359,N_9106,N_9506);
xnor U11360 (N_11360,N_8062,N_8140);
or U11361 (N_11361,N_9095,N_8357);
xnor U11362 (N_11362,N_9690,N_8406);
nand U11363 (N_11363,N_8692,N_9777);
nor U11364 (N_11364,N_9492,N_9069);
nor U11365 (N_11365,N_8540,N_9799);
nor U11366 (N_11366,N_8401,N_9831);
and U11367 (N_11367,N_8408,N_9290);
nor U11368 (N_11368,N_9800,N_9175);
xor U11369 (N_11369,N_9328,N_8611);
nand U11370 (N_11370,N_9807,N_9495);
xor U11371 (N_11371,N_9531,N_8023);
xnor U11372 (N_11372,N_9057,N_8271);
nor U11373 (N_11373,N_8815,N_9137);
xnor U11374 (N_11374,N_8311,N_8988);
xnor U11375 (N_11375,N_8125,N_8110);
nand U11376 (N_11376,N_9959,N_9769);
nand U11377 (N_11377,N_8315,N_8207);
xor U11378 (N_11378,N_8108,N_8369);
or U11379 (N_11379,N_9794,N_9203);
nand U11380 (N_11380,N_8860,N_9761);
xnor U11381 (N_11381,N_9494,N_8580);
and U11382 (N_11382,N_9103,N_8920);
nor U11383 (N_11383,N_9198,N_9168);
and U11384 (N_11384,N_8413,N_9884);
nor U11385 (N_11385,N_8679,N_9816);
xor U11386 (N_11386,N_9873,N_9377);
nand U11387 (N_11387,N_8352,N_9481);
or U11388 (N_11388,N_8551,N_8399);
nand U11389 (N_11389,N_8077,N_9831);
or U11390 (N_11390,N_8577,N_9753);
nor U11391 (N_11391,N_9262,N_9941);
nand U11392 (N_11392,N_9652,N_8151);
nor U11393 (N_11393,N_8736,N_8065);
nand U11394 (N_11394,N_9695,N_9930);
xor U11395 (N_11395,N_9902,N_9039);
nor U11396 (N_11396,N_9066,N_8643);
nor U11397 (N_11397,N_8032,N_9999);
or U11398 (N_11398,N_9066,N_8908);
xor U11399 (N_11399,N_8954,N_8676);
or U11400 (N_11400,N_9772,N_8199);
nand U11401 (N_11401,N_9126,N_9634);
and U11402 (N_11402,N_9631,N_8980);
xor U11403 (N_11403,N_8945,N_9833);
and U11404 (N_11404,N_8238,N_9847);
nor U11405 (N_11405,N_9593,N_8316);
nand U11406 (N_11406,N_9176,N_9605);
xor U11407 (N_11407,N_9939,N_8277);
and U11408 (N_11408,N_8048,N_8180);
or U11409 (N_11409,N_8227,N_9277);
nor U11410 (N_11410,N_8936,N_9847);
xnor U11411 (N_11411,N_9291,N_8766);
xnor U11412 (N_11412,N_8084,N_8364);
nand U11413 (N_11413,N_8336,N_8699);
or U11414 (N_11414,N_8475,N_9897);
nor U11415 (N_11415,N_8962,N_9984);
nand U11416 (N_11416,N_9041,N_9255);
and U11417 (N_11417,N_9244,N_8443);
xor U11418 (N_11418,N_9685,N_9731);
xor U11419 (N_11419,N_9253,N_8086);
or U11420 (N_11420,N_9514,N_9021);
xnor U11421 (N_11421,N_8177,N_8370);
nand U11422 (N_11422,N_8079,N_9938);
nand U11423 (N_11423,N_9055,N_9482);
nand U11424 (N_11424,N_9509,N_9107);
or U11425 (N_11425,N_8584,N_9667);
xor U11426 (N_11426,N_8145,N_8702);
nor U11427 (N_11427,N_9812,N_8259);
nor U11428 (N_11428,N_8731,N_8361);
nand U11429 (N_11429,N_9304,N_8910);
and U11430 (N_11430,N_9494,N_9118);
xor U11431 (N_11431,N_9944,N_8130);
and U11432 (N_11432,N_8416,N_8539);
and U11433 (N_11433,N_8766,N_8112);
or U11434 (N_11434,N_9624,N_9678);
nor U11435 (N_11435,N_9314,N_9658);
xor U11436 (N_11436,N_9034,N_8219);
and U11437 (N_11437,N_8570,N_8016);
xor U11438 (N_11438,N_9736,N_8064);
nor U11439 (N_11439,N_9256,N_8115);
nor U11440 (N_11440,N_8561,N_8254);
xnor U11441 (N_11441,N_8207,N_8340);
xor U11442 (N_11442,N_9180,N_8249);
and U11443 (N_11443,N_9891,N_9325);
and U11444 (N_11444,N_9034,N_9751);
or U11445 (N_11445,N_9257,N_9638);
nand U11446 (N_11446,N_8483,N_9441);
nor U11447 (N_11447,N_9248,N_8607);
nor U11448 (N_11448,N_9983,N_9161);
xor U11449 (N_11449,N_9830,N_8542);
or U11450 (N_11450,N_9223,N_9685);
nand U11451 (N_11451,N_8340,N_8284);
xor U11452 (N_11452,N_9570,N_8476);
nor U11453 (N_11453,N_8799,N_8142);
and U11454 (N_11454,N_9286,N_9331);
or U11455 (N_11455,N_9021,N_9373);
nand U11456 (N_11456,N_9000,N_8017);
nor U11457 (N_11457,N_8045,N_9518);
or U11458 (N_11458,N_9004,N_8438);
and U11459 (N_11459,N_8672,N_9083);
and U11460 (N_11460,N_9802,N_8915);
nor U11461 (N_11461,N_8053,N_9739);
nor U11462 (N_11462,N_8285,N_8792);
nand U11463 (N_11463,N_8643,N_8086);
and U11464 (N_11464,N_9543,N_9534);
xnor U11465 (N_11465,N_8509,N_9349);
and U11466 (N_11466,N_9482,N_8214);
or U11467 (N_11467,N_8089,N_9355);
xor U11468 (N_11468,N_8952,N_8820);
nand U11469 (N_11469,N_9288,N_9076);
nand U11470 (N_11470,N_9236,N_9838);
nand U11471 (N_11471,N_9899,N_9349);
and U11472 (N_11472,N_8858,N_9165);
nor U11473 (N_11473,N_9792,N_8331);
or U11474 (N_11474,N_9193,N_9923);
and U11475 (N_11475,N_8224,N_9642);
xnor U11476 (N_11476,N_9393,N_8181);
xor U11477 (N_11477,N_9524,N_8790);
and U11478 (N_11478,N_9289,N_8883);
nand U11479 (N_11479,N_9072,N_8035);
nor U11480 (N_11480,N_9497,N_8052);
or U11481 (N_11481,N_9425,N_9925);
xnor U11482 (N_11482,N_8836,N_9329);
or U11483 (N_11483,N_9756,N_8228);
xnor U11484 (N_11484,N_9544,N_8176);
nand U11485 (N_11485,N_8211,N_8895);
xor U11486 (N_11486,N_9951,N_9034);
nor U11487 (N_11487,N_8588,N_9781);
or U11488 (N_11488,N_9926,N_9872);
xnor U11489 (N_11489,N_9355,N_9646);
or U11490 (N_11490,N_9335,N_8845);
nand U11491 (N_11491,N_9992,N_9523);
xor U11492 (N_11492,N_8067,N_8047);
nor U11493 (N_11493,N_9525,N_8532);
nor U11494 (N_11494,N_8308,N_9019);
nor U11495 (N_11495,N_9598,N_8091);
nand U11496 (N_11496,N_8051,N_8521);
xnor U11497 (N_11497,N_9176,N_9887);
and U11498 (N_11498,N_9495,N_9508);
nand U11499 (N_11499,N_8469,N_8759);
or U11500 (N_11500,N_9398,N_8108);
nand U11501 (N_11501,N_8819,N_8547);
nand U11502 (N_11502,N_8295,N_9452);
or U11503 (N_11503,N_8880,N_8644);
xnor U11504 (N_11504,N_9738,N_8678);
and U11505 (N_11505,N_8455,N_8691);
nor U11506 (N_11506,N_8447,N_8896);
and U11507 (N_11507,N_9351,N_8068);
and U11508 (N_11508,N_8707,N_8053);
and U11509 (N_11509,N_9386,N_9828);
nand U11510 (N_11510,N_8828,N_8091);
xnor U11511 (N_11511,N_9085,N_9557);
and U11512 (N_11512,N_8383,N_8666);
and U11513 (N_11513,N_8862,N_8512);
or U11514 (N_11514,N_9447,N_8885);
xor U11515 (N_11515,N_8907,N_9690);
or U11516 (N_11516,N_8184,N_8430);
and U11517 (N_11517,N_8515,N_8152);
xor U11518 (N_11518,N_8675,N_8519);
nand U11519 (N_11519,N_8560,N_9980);
nor U11520 (N_11520,N_9337,N_8536);
nand U11521 (N_11521,N_9727,N_9818);
nand U11522 (N_11522,N_9764,N_8167);
or U11523 (N_11523,N_9893,N_9577);
nand U11524 (N_11524,N_9675,N_9392);
nand U11525 (N_11525,N_8142,N_9934);
nor U11526 (N_11526,N_8237,N_9560);
xor U11527 (N_11527,N_9536,N_9548);
or U11528 (N_11528,N_9195,N_9545);
and U11529 (N_11529,N_8639,N_9514);
or U11530 (N_11530,N_8250,N_8376);
nand U11531 (N_11531,N_9898,N_9463);
or U11532 (N_11532,N_8810,N_9192);
and U11533 (N_11533,N_8525,N_9737);
or U11534 (N_11534,N_9568,N_8700);
xor U11535 (N_11535,N_8281,N_8029);
xor U11536 (N_11536,N_9363,N_8403);
nor U11537 (N_11537,N_9514,N_9285);
and U11538 (N_11538,N_8678,N_9062);
nor U11539 (N_11539,N_8358,N_9662);
xor U11540 (N_11540,N_8644,N_8997);
or U11541 (N_11541,N_8025,N_9616);
and U11542 (N_11542,N_8724,N_9498);
xor U11543 (N_11543,N_9542,N_9125);
nand U11544 (N_11544,N_9751,N_8165);
xnor U11545 (N_11545,N_8984,N_9461);
or U11546 (N_11546,N_8328,N_9148);
or U11547 (N_11547,N_8777,N_8752);
nor U11548 (N_11548,N_8520,N_9247);
nor U11549 (N_11549,N_8196,N_9286);
nand U11550 (N_11550,N_8978,N_9814);
or U11551 (N_11551,N_8120,N_9589);
and U11552 (N_11552,N_9164,N_9582);
and U11553 (N_11553,N_8098,N_9551);
xnor U11554 (N_11554,N_9740,N_9062);
or U11555 (N_11555,N_9500,N_8816);
nand U11556 (N_11556,N_8738,N_9594);
nor U11557 (N_11557,N_8598,N_8433);
xnor U11558 (N_11558,N_8972,N_9441);
or U11559 (N_11559,N_9451,N_9973);
nand U11560 (N_11560,N_9039,N_9268);
nand U11561 (N_11561,N_8217,N_9584);
and U11562 (N_11562,N_9703,N_9177);
nor U11563 (N_11563,N_8102,N_9849);
or U11564 (N_11564,N_8282,N_8344);
and U11565 (N_11565,N_9463,N_9511);
or U11566 (N_11566,N_8087,N_8842);
and U11567 (N_11567,N_9188,N_8705);
or U11568 (N_11568,N_8208,N_8225);
xnor U11569 (N_11569,N_9651,N_9245);
nor U11570 (N_11570,N_9221,N_9495);
or U11571 (N_11571,N_9115,N_8011);
or U11572 (N_11572,N_9404,N_8407);
nand U11573 (N_11573,N_9708,N_9532);
nor U11574 (N_11574,N_8813,N_9067);
nor U11575 (N_11575,N_8356,N_9762);
or U11576 (N_11576,N_9450,N_9567);
or U11577 (N_11577,N_8201,N_8456);
or U11578 (N_11578,N_9277,N_8375);
nor U11579 (N_11579,N_8361,N_8335);
xor U11580 (N_11580,N_8642,N_8114);
nand U11581 (N_11581,N_8312,N_8999);
xor U11582 (N_11582,N_8771,N_9533);
nand U11583 (N_11583,N_9629,N_9620);
nor U11584 (N_11584,N_8254,N_8977);
and U11585 (N_11585,N_8543,N_9505);
nor U11586 (N_11586,N_9622,N_8108);
xor U11587 (N_11587,N_8602,N_9707);
or U11588 (N_11588,N_9262,N_8261);
nand U11589 (N_11589,N_8801,N_9865);
xor U11590 (N_11590,N_9566,N_8360);
or U11591 (N_11591,N_8769,N_9139);
nor U11592 (N_11592,N_9598,N_8277);
xor U11593 (N_11593,N_9096,N_8923);
or U11594 (N_11594,N_8070,N_8735);
nand U11595 (N_11595,N_8843,N_9382);
nor U11596 (N_11596,N_9086,N_9406);
nand U11597 (N_11597,N_9561,N_8850);
xnor U11598 (N_11598,N_8065,N_8617);
nand U11599 (N_11599,N_9878,N_9857);
xnor U11600 (N_11600,N_9616,N_9825);
or U11601 (N_11601,N_9238,N_8946);
xor U11602 (N_11602,N_8025,N_9330);
xnor U11603 (N_11603,N_8503,N_8310);
or U11604 (N_11604,N_9363,N_9765);
xnor U11605 (N_11605,N_8083,N_8171);
nand U11606 (N_11606,N_8891,N_9482);
nor U11607 (N_11607,N_9424,N_8422);
or U11608 (N_11608,N_8872,N_8698);
nand U11609 (N_11609,N_9511,N_8143);
or U11610 (N_11610,N_9056,N_9676);
and U11611 (N_11611,N_9764,N_8117);
or U11612 (N_11612,N_8693,N_9957);
xnor U11613 (N_11613,N_8472,N_9273);
nand U11614 (N_11614,N_9429,N_8149);
nand U11615 (N_11615,N_8580,N_8040);
nor U11616 (N_11616,N_9236,N_8462);
nand U11617 (N_11617,N_9588,N_9010);
nand U11618 (N_11618,N_9368,N_9814);
or U11619 (N_11619,N_8377,N_9223);
nor U11620 (N_11620,N_8710,N_8772);
or U11621 (N_11621,N_8745,N_8853);
nand U11622 (N_11622,N_9023,N_9162);
and U11623 (N_11623,N_9780,N_8263);
or U11624 (N_11624,N_8034,N_9449);
or U11625 (N_11625,N_9740,N_8098);
or U11626 (N_11626,N_8255,N_8825);
nor U11627 (N_11627,N_8539,N_9199);
nand U11628 (N_11628,N_8611,N_9938);
nor U11629 (N_11629,N_8659,N_8446);
nand U11630 (N_11630,N_9280,N_9355);
nand U11631 (N_11631,N_8564,N_8147);
and U11632 (N_11632,N_9326,N_8219);
xor U11633 (N_11633,N_8338,N_8915);
nand U11634 (N_11634,N_8879,N_8625);
nand U11635 (N_11635,N_8158,N_9929);
and U11636 (N_11636,N_9416,N_8861);
or U11637 (N_11637,N_8989,N_9489);
nand U11638 (N_11638,N_8655,N_8064);
nand U11639 (N_11639,N_8880,N_8239);
nand U11640 (N_11640,N_8250,N_9148);
and U11641 (N_11641,N_8985,N_8638);
and U11642 (N_11642,N_8950,N_8378);
nor U11643 (N_11643,N_9218,N_9358);
xnor U11644 (N_11644,N_9887,N_9781);
nor U11645 (N_11645,N_9499,N_8876);
xor U11646 (N_11646,N_8358,N_9569);
xnor U11647 (N_11647,N_8102,N_9656);
nor U11648 (N_11648,N_9691,N_9439);
nand U11649 (N_11649,N_9916,N_8258);
xor U11650 (N_11650,N_9450,N_9687);
nand U11651 (N_11651,N_8870,N_8625);
xnor U11652 (N_11652,N_9460,N_8576);
nor U11653 (N_11653,N_9209,N_9457);
or U11654 (N_11654,N_8253,N_8574);
and U11655 (N_11655,N_9903,N_8052);
nor U11656 (N_11656,N_9273,N_8674);
xor U11657 (N_11657,N_9556,N_9429);
and U11658 (N_11658,N_8865,N_9278);
nor U11659 (N_11659,N_9856,N_8507);
xor U11660 (N_11660,N_8820,N_8801);
xnor U11661 (N_11661,N_9174,N_9614);
xor U11662 (N_11662,N_9514,N_8787);
or U11663 (N_11663,N_8503,N_9618);
or U11664 (N_11664,N_8408,N_9968);
or U11665 (N_11665,N_8723,N_8467);
nand U11666 (N_11666,N_9097,N_9844);
and U11667 (N_11667,N_9247,N_8613);
nor U11668 (N_11668,N_9294,N_8959);
or U11669 (N_11669,N_8396,N_8222);
xor U11670 (N_11670,N_9781,N_8010);
or U11671 (N_11671,N_8817,N_9333);
and U11672 (N_11672,N_8623,N_9426);
and U11673 (N_11673,N_8153,N_8972);
nand U11674 (N_11674,N_8404,N_9644);
nand U11675 (N_11675,N_8016,N_8058);
nor U11676 (N_11676,N_9752,N_8923);
xor U11677 (N_11677,N_9794,N_9137);
and U11678 (N_11678,N_8004,N_8788);
or U11679 (N_11679,N_9546,N_9525);
nor U11680 (N_11680,N_9499,N_9636);
and U11681 (N_11681,N_8764,N_8433);
or U11682 (N_11682,N_8791,N_8081);
nand U11683 (N_11683,N_9865,N_9168);
nand U11684 (N_11684,N_8978,N_9281);
or U11685 (N_11685,N_9565,N_9759);
and U11686 (N_11686,N_8689,N_8597);
or U11687 (N_11687,N_9197,N_8576);
and U11688 (N_11688,N_9739,N_8464);
and U11689 (N_11689,N_8844,N_9219);
xor U11690 (N_11690,N_9078,N_8162);
and U11691 (N_11691,N_9545,N_9280);
and U11692 (N_11692,N_8105,N_9675);
nor U11693 (N_11693,N_8942,N_9218);
and U11694 (N_11694,N_9486,N_8589);
nand U11695 (N_11695,N_8065,N_8645);
or U11696 (N_11696,N_9411,N_8560);
and U11697 (N_11697,N_9031,N_9456);
nor U11698 (N_11698,N_8797,N_8107);
nand U11699 (N_11699,N_8405,N_8863);
and U11700 (N_11700,N_9668,N_8322);
nor U11701 (N_11701,N_9363,N_8831);
xor U11702 (N_11702,N_8613,N_8073);
nand U11703 (N_11703,N_8747,N_9269);
or U11704 (N_11704,N_8074,N_9137);
or U11705 (N_11705,N_9049,N_9512);
nand U11706 (N_11706,N_9502,N_8245);
nor U11707 (N_11707,N_8531,N_9428);
nand U11708 (N_11708,N_9460,N_9387);
and U11709 (N_11709,N_8440,N_8007);
and U11710 (N_11710,N_9073,N_8951);
nand U11711 (N_11711,N_8206,N_9752);
nand U11712 (N_11712,N_8294,N_8477);
xnor U11713 (N_11713,N_8893,N_9701);
nand U11714 (N_11714,N_8955,N_8565);
or U11715 (N_11715,N_8520,N_8267);
or U11716 (N_11716,N_8776,N_8539);
nand U11717 (N_11717,N_9789,N_8820);
xnor U11718 (N_11718,N_8322,N_9001);
or U11719 (N_11719,N_8583,N_8971);
nand U11720 (N_11720,N_9019,N_9538);
xor U11721 (N_11721,N_8985,N_9493);
nand U11722 (N_11722,N_8083,N_9960);
xnor U11723 (N_11723,N_8179,N_8023);
and U11724 (N_11724,N_8281,N_8730);
and U11725 (N_11725,N_9801,N_9281);
nor U11726 (N_11726,N_9430,N_9626);
nor U11727 (N_11727,N_9153,N_8611);
nand U11728 (N_11728,N_9501,N_8543);
nand U11729 (N_11729,N_8474,N_9574);
and U11730 (N_11730,N_8585,N_9991);
nor U11731 (N_11731,N_8734,N_8865);
nor U11732 (N_11732,N_9265,N_9014);
nor U11733 (N_11733,N_8604,N_8943);
or U11734 (N_11734,N_8496,N_8220);
or U11735 (N_11735,N_8660,N_8709);
or U11736 (N_11736,N_9456,N_8820);
nor U11737 (N_11737,N_8080,N_9307);
xor U11738 (N_11738,N_8707,N_9368);
nor U11739 (N_11739,N_8284,N_8568);
and U11740 (N_11740,N_9610,N_8596);
nand U11741 (N_11741,N_9905,N_8402);
nor U11742 (N_11742,N_9577,N_8581);
nand U11743 (N_11743,N_8579,N_8207);
nor U11744 (N_11744,N_9070,N_9076);
or U11745 (N_11745,N_9528,N_9600);
nand U11746 (N_11746,N_9492,N_8805);
nand U11747 (N_11747,N_8258,N_8334);
or U11748 (N_11748,N_9949,N_9867);
xor U11749 (N_11749,N_9724,N_8540);
or U11750 (N_11750,N_9151,N_8668);
nor U11751 (N_11751,N_9421,N_9319);
or U11752 (N_11752,N_8776,N_9493);
and U11753 (N_11753,N_8394,N_9273);
or U11754 (N_11754,N_8786,N_8557);
or U11755 (N_11755,N_8512,N_8470);
nand U11756 (N_11756,N_8009,N_9233);
xnor U11757 (N_11757,N_9627,N_9479);
or U11758 (N_11758,N_8909,N_9251);
or U11759 (N_11759,N_9551,N_9997);
xnor U11760 (N_11760,N_8860,N_9645);
xnor U11761 (N_11761,N_9530,N_9103);
and U11762 (N_11762,N_9641,N_8159);
xnor U11763 (N_11763,N_8300,N_9949);
or U11764 (N_11764,N_8498,N_8457);
or U11765 (N_11765,N_8613,N_8616);
and U11766 (N_11766,N_9587,N_9766);
nor U11767 (N_11767,N_9316,N_9231);
xnor U11768 (N_11768,N_8858,N_8584);
nand U11769 (N_11769,N_9808,N_8847);
nor U11770 (N_11770,N_9532,N_9191);
and U11771 (N_11771,N_9619,N_8196);
xnor U11772 (N_11772,N_9420,N_8899);
nor U11773 (N_11773,N_9785,N_8694);
nand U11774 (N_11774,N_9229,N_8101);
or U11775 (N_11775,N_8455,N_8935);
nand U11776 (N_11776,N_8204,N_9588);
nand U11777 (N_11777,N_8526,N_8282);
xnor U11778 (N_11778,N_8926,N_9187);
and U11779 (N_11779,N_9689,N_9698);
and U11780 (N_11780,N_8079,N_9367);
and U11781 (N_11781,N_9602,N_9932);
xnor U11782 (N_11782,N_9005,N_8831);
or U11783 (N_11783,N_8174,N_8635);
xnor U11784 (N_11784,N_9977,N_8794);
or U11785 (N_11785,N_8879,N_8526);
and U11786 (N_11786,N_8715,N_9431);
or U11787 (N_11787,N_8936,N_9523);
or U11788 (N_11788,N_9927,N_8971);
nand U11789 (N_11789,N_9105,N_8932);
xnor U11790 (N_11790,N_9337,N_9736);
nor U11791 (N_11791,N_9072,N_8006);
xor U11792 (N_11792,N_8604,N_8122);
nand U11793 (N_11793,N_9063,N_9152);
and U11794 (N_11794,N_8421,N_9741);
or U11795 (N_11795,N_8861,N_9065);
xor U11796 (N_11796,N_9115,N_9601);
xor U11797 (N_11797,N_9027,N_9021);
nand U11798 (N_11798,N_9647,N_8819);
xor U11799 (N_11799,N_9783,N_8032);
and U11800 (N_11800,N_9135,N_8211);
nor U11801 (N_11801,N_9640,N_9781);
or U11802 (N_11802,N_8976,N_8678);
or U11803 (N_11803,N_9191,N_9167);
and U11804 (N_11804,N_8706,N_8748);
and U11805 (N_11805,N_8596,N_9131);
or U11806 (N_11806,N_8965,N_8503);
and U11807 (N_11807,N_9491,N_8335);
nor U11808 (N_11808,N_9562,N_9633);
and U11809 (N_11809,N_9166,N_8843);
nor U11810 (N_11810,N_9821,N_8997);
or U11811 (N_11811,N_9598,N_9659);
or U11812 (N_11812,N_8825,N_8319);
nor U11813 (N_11813,N_8762,N_9332);
and U11814 (N_11814,N_8120,N_9274);
nand U11815 (N_11815,N_9229,N_9176);
nand U11816 (N_11816,N_9951,N_8226);
or U11817 (N_11817,N_8632,N_9330);
xor U11818 (N_11818,N_8439,N_9201);
xor U11819 (N_11819,N_9608,N_8029);
or U11820 (N_11820,N_9516,N_8037);
xor U11821 (N_11821,N_8627,N_9116);
xor U11822 (N_11822,N_8476,N_9021);
or U11823 (N_11823,N_9097,N_9715);
nor U11824 (N_11824,N_9128,N_8047);
nor U11825 (N_11825,N_8437,N_8441);
xor U11826 (N_11826,N_8360,N_8659);
or U11827 (N_11827,N_8885,N_9152);
or U11828 (N_11828,N_8789,N_8462);
nor U11829 (N_11829,N_8856,N_8145);
and U11830 (N_11830,N_9604,N_9639);
nand U11831 (N_11831,N_8284,N_9432);
nor U11832 (N_11832,N_9659,N_8223);
or U11833 (N_11833,N_9024,N_9930);
nor U11834 (N_11834,N_9281,N_9699);
xnor U11835 (N_11835,N_9917,N_8119);
nand U11836 (N_11836,N_9900,N_8366);
nor U11837 (N_11837,N_9860,N_9508);
and U11838 (N_11838,N_8020,N_8130);
nand U11839 (N_11839,N_8144,N_9169);
nand U11840 (N_11840,N_9720,N_8081);
nor U11841 (N_11841,N_9839,N_9763);
nor U11842 (N_11842,N_9430,N_8755);
nor U11843 (N_11843,N_8840,N_9040);
nor U11844 (N_11844,N_8044,N_9494);
nor U11845 (N_11845,N_8824,N_8395);
xor U11846 (N_11846,N_9277,N_9679);
or U11847 (N_11847,N_9995,N_8002);
or U11848 (N_11848,N_8020,N_8910);
and U11849 (N_11849,N_9639,N_9523);
nor U11850 (N_11850,N_8486,N_9136);
xor U11851 (N_11851,N_8957,N_8419);
nor U11852 (N_11852,N_8358,N_8596);
nand U11853 (N_11853,N_9478,N_9856);
nor U11854 (N_11854,N_9019,N_9194);
or U11855 (N_11855,N_9593,N_8849);
xor U11856 (N_11856,N_8307,N_9543);
or U11857 (N_11857,N_8857,N_8597);
and U11858 (N_11858,N_9807,N_8327);
and U11859 (N_11859,N_9265,N_9158);
and U11860 (N_11860,N_8560,N_9284);
and U11861 (N_11861,N_9121,N_9289);
or U11862 (N_11862,N_8645,N_9697);
nor U11863 (N_11863,N_8407,N_9253);
and U11864 (N_11864,N_9377,N_9954);
and U11865 (N_11865,N_9145,N_8777);
nand U11866 (N_11866,N_8928,N_9881);
xnor U11867 (N_11867,N_8264,N_8197);
nand U11868 (N_11868,N_9627,N_8585);
nand U11869 (N_11869,N_9408,N_9333);
and U11870 (N_11870,N_8849,N_9654);
or U11871 (N_11871,N_8166,N_8746);
and U11872 (N_11872,N_8033,N_8717);
and U11873 (N_11873,N_8203,N_8329);
or U11874 (N_11874,N_8344,N_8953);
nand U11875 (N_11875,N_8848,N_9152);
nand U11876 (N_11876,N_8345,N_8385);
xnor U11877 (N_11877,N_9076,N_9207);
nor U11878 (N_11878,N_8919,N_9532);
nand U11879 (N_11879,N_8300,N_8631);
or U11880 (N_11880,N_9034,N_9817);
nor U11881 (N_11881,N_9813,N_9298);
nor U11882 (N_11882,N_9215,N_8727);
nor U11883 (N_11883,N_9820,N_9243);
nor U11884 (N_11884,N_8135,N_9662);
xor U11885 (N_11885,N_8745,N_8649);
nor U11886 (N_11886,N_8349,N_8662);
nand U11887 (N_11887,N_9866,N_8330);
and U11888 (N_11888,N_8875,N_8988);
nor U11889 (N_11889,N_9902,N_8276);
nand U11890 (N_11890,N_8605,N_8848);
nand U11891 (N_11891,N_9830,N_9521);
xor U11892 (N_11892,N_9454,N_9468);
nand U11893 (N_11893,N_8867,N_9259);
nand U11894 (N_11894,N_8886,N_8826);
nor U11895 (N_11895,N_8267,N_8251);
xor U11896 (N_11896,N_8685,N_8153);
xnor U11897 (N_11897,N_8415,N_8474);
nand U11898 (N_11898,N_9161,N_9073);
nand U11899 (N_11899,N_9732,N_8674);
nand U11900 (N_11900,N_9667,N_9615);
and U11901 (N_11901,N_8780,N_9194);
xnor U11902 (N_11902,N_8778,N_8875);
xnor U11903 (N_11903,N_8935,N_8478);
or U11904 (N_11904,N_8841,N_9851);
nor U11905 (N_11905,N_9196,N_9418);
or U11906 (N_11906,N_8139,N_9139);
or U11907 (N_11907,N_9175,N_9465);
or U11908 (N_11908,N_8670,N_8026);
or U11909 (N_11909,N_8871,N_8033);
nand U11910 (N_11910,N_8210,N_9059);
nor U11911 (N_11911,N_8042,N_8203);
nor U11912 (N_11912,N_8068,N_9759);
or U11913 (N_11913,N_8189,N_8335);
nand U11914 (N_11914,N_8702,N_9058);
nand U11915 (N_11915,N_8550,N_9188);
nand U11916 (N_11916,N_8669,N_8999);
nand U11917 (N_11917,N_9560,N_8240);
nand U11918 (N_11918,N_8086,N_9674);
or U11919 (N_11919,N_8087,N_9823);
or U11920 (N_11920,N_8662,N_8386);
and U11921 (N_11921,N_9398,N_8233);
xnor U11922 (N_11922,N_9696,N_8487);
nor U11923 (N_11923,N_9871,N_8331);
nand U11924 (N_11924,N_9286,N_9885);
or U11925 (N_11925,N_9473,N_8433);
or U11926 (N_11926,N_9061,N_8135);
or U11927 (N_11927,N_9929,N_9260);
nand U11928 (N_11928,N_8190,N_8518);
or U11929 (N_11929,N_9246,N_9215);
nor U11930 (N_11930,N_8033,N_8339);
xor U11931 (N_11931,N_9340,N_9138);
xnor U11932 (N_11932,N_9106,N_8668);
xnor U11933 (N_11933,N_9718,N_8900);
and U11934 (N_11934,N_8544,N_8500);
nand U11935 (N_11935,N_9708,N_9318);
nor U11936 (N_11936,N_8429,N_9189);
nand U11937 (N_11937,N_9764,N_8148);
xnor U11938 (N_11938,N_8562,N_9181);
or U11939 (N_11939,N_9192,N_9676);
xor U11940 (N_11940,N_8426,N_8268);
nor U11941 (N_11941,N_9503,N_9087);
or U11942 (N_11942,N_8508,N_9461);
xor U11943 (N_11943,N_8513,N_9620);
nand U11944 (N_11944,N_8178,N_8834);
or U11945 (N_11945,N_9399,N_9557);
nand U11946 (N_11946,N_9109,N_9216);
or U11947 (N_11947,N_9709,N_9238);
and U11948 (N_11948,N_8888,N_9357);
nand U11949 (N_11949,N_8407,N_9256);
and U11950 (N_11950,N_8929,N_9240);
or U11951 (N_11951,N_9865,N_9614);
nor U11952 (N_11952,N_9258,N_9082);
and U11953 (N_11953,N_9232,N_8658);
nor U11954 (N_11954,N_9804,N_8999);
xor U11955 (N_11955,N_8952,N_9895);
xnor U11956 (N_11956,N_9617,N_9753);
nand U11957 (N_11957,N_9856,N_8428);
or U11958 (N_11958,N_9442,N_9274);
nand U11959 (N_11959,N_9115,N_9634);
xnor U11960 (N_11960,N_9384,N_9936);
or U11961 (N_11961,N_9460,N_8133);
or U11962 (N_11962,N_9113,N_8649);
nor U11963 (N_11963,N_9350,N_8310);
or U11964 (N_11964,N_8329,N_9917);
nand U11965 (N_11965,N_8194,N_8282);
and U11966 (N_11966,N_8821,N_9491);
nand U11967 (N_11967,N_9645,N_8522);
xnor U11968 (N_11968,N_9209,N_9808);
or U11969 (N_11969,N_8495,N_8341);
and U11970 (N_11970,N_9555,N_8778);
or U11971 (N_11971,N_9109,N_8768);
nand U11972 (N_11972,N_8116,N_8570);
nand U11973 (N_11973,N_8483,N_9748);
xor U11974 (N_11974,N_8393,N_8550);
nor U11975 (N_11975,N_9135,N_8987);
nand U11976 (N_11976,N_8255,N_8799);
and U11977 (N_11977,N_8049,N_8348);
nor U11978 (N_11978,N_9200,N_9564);
xnor U11979 (N_11979,N_8078,N_8124);
xor U11980 (N_11980,N_9415,N_8364);
nor U11981 (N_11981,N_9231,N_9879);
xnor U11982 (N_11982,N_8543,N_9473);
xor U11983 (N_11983,N_8774,N_9072);
xor U11984 (N_11984,N_9850,N_9282);
or U11985 (N_11985,N_8359,N_9467);
or U11986 (N_11986,N_8676,N_8995);
nor U11987 (N_11987,N_9317,N_8399);
and U11988 (N_11988,N_9666,N_8090);
xnor U11989 (N_11989,N_8644,N_8661);
and U11990 (N_11990,N_8323,N_8723);
xnor U11991 (N_11991,N_8619,N_8986);
or U11992 (N_11992,N_8417,N_9239);
and U11993 (N_11993,N_9737,N_9754);
nand U11994 (N_11994,N_8847,N_8683);
xor U11995 (N_11995,N_8183,N_8773);
or U11996 (N_11996,N_9472,N_8322);
nor U11997 (N_11997,N_9210,N_9023);
or U11998 (N_11998,N_8464,N_8466);
xnor U11999 (N_11999,N_8699,N_9631);
nand U12000 (N_12000,N_10365,N_10646);
and U12001 (N_12001,N_11181,N_11782);
and U12002 (N_12002,N_11477,N_11584);
nand U12003 (N_12003,N_11301,N_11257);
and U12004 (N_12004,N_10504,N_11825);
or U12005 (N_12005,N_11734,N_11211);
nor U12006 (N_12006,N_11580,N_11576);
nand U12007 (N_12007,N_10501,N_10438);
nand U12008 (N_12008,N_10554,N_10741);
or U12009 (N_12009,N_11235,N_10856);
xor U12010 (N_12010,N_10650,N_10642);
nor U12011 (N_12011,N_11546,N_11493);
xnor U12012 (N_12012,N_10989,N_11896);
or U12013 (N_12013,N_10923,N_10335);
nand U12014 (N_12014,N_10291,N_11041);
and U12015 (N_12015,N_11661,N_10000);
xor U12016 (N_12016,N_11070,N_10657);
xor U12017 (N_12017,N_11474,N_11590);
xnor U12018 (N_12018,N_10510,N_10987);
and U12019 (N_12019,N_10878,N_11586);
and U12020 (N_12020,N_10742,N_11357);
or U12021 (N_12021,N_11884,N_10697);
nand U12022 (N_12022,N_11690,N_11682);
and U12023 (N_12023,N_11623,N_11753);
nand U12024 (N_12024,N_11908,N_10991);
or U12025 (N_12025,N_10986,N_11891);
nor U12026 (N_12026,N_11605,N_11127);
and U12027 (N_12027,N_10421,N_10071);
nand U12028 (N_12028,N_11379,N_10324);
or U12029 (N_12029,N_10933,N_10505);
or U12030 (N_12030,N_10569,N_11579);
and U12031 (N_12031,N_11885,N_11361);
or U12032 (N_12032,N_11777,N_10435);
xor U12033 (N_12033,N_10561,N_11221);
xor U12034 (N_12034,N_11043,N_10731);
xor U12035 (N_12035,N_11273,N_10252);
xor U12036 (N_12036,N_10573,N_11748);
nand U12037 (N_12037,N_10468,N_10683);
xnor U12038 (N_12038,N_11616,N_10436);
or U12039 (N_12039,N_11323,N_11241);
nand U12040 (N_12040,N_10549,N_10350);
xnor U12041 (N_12041,N_11478,N_10068);
and U12042 (N_12042,N_11010,N_10928);
or U12043 (N_12043,N_10719,N_11383);
and U12044 (N_12044,N_11700,N_10883);
xnor U12045 (N_12045,N_11621,N_10442);
nor U12046 (N_12046,N_10298,N_11141);
nor U12047 (N_12047,N_10248,N_11712);
nor U12048 (N_12048,N_10607,N_10728);
and U12049 (N_12049,N_10242,N_10775);
nor U12050 (N_12050,N_11069,N_10149);
nand U12051 (N_12051,N_11762,N_10545);
nand U12052 (N_12052,N_10823,N_10179);
and U12053 (N_12053,N_10694,N_11089);
or U12054 (N_12054,N_11341,N_11485);
xnor U12055 (N_12055,N_11557,N_10849);
or U12056 (N_12056,N_11467,N_10391);
xnor U12057 (N_12057,N_11456,N_10144);
xnor U12058 (N_12058,N_10115,N_11611);
or U12059 (N_12059,N_11677,N_11191);
or U12060 (N_12060,N_10089,N_10379);
or U12061 (N_12061,N_11658,N_11511);
nor U12062 (N_12062,N_10571,N_10723);
nor U12063 (N_12063,N_11374,N_11567);
xor U12064 (N_12064,N_11130,N_11465);
nor U12065 (N_12065,N_11669,N_10401);
and U12066 (N_12066,N_10613,N_11154);
or U12067 (N_12067,N_10825,N_10114);
xnor U12068 (N_12068,N_10695,N_10205);
xnor U12069 (N_12069,N_11117,N_11376);
and U12070 (N_12070,N_10811,N_11801);
and U12071 (N_12071,N_11670,N_11166);
or U12072 (N_12072,N_11932,N_11672);
xnor U12073 (N_12073,N_10389,N_10272);
and U12074 (N_12074,N_11197,N_10603);
and U12075 (N_12075,N_11327,N_10032);
or U12076 (N_12076,N_11086,N_10629);
nor U12077 (N_12077,N_10537,N_10064);
nor U12078 (N_12078,N_11495,N_10790);
xor U12079 (N_12079,N_11346,N_11104);
nand U12080 (N_12080,N_10460,N_11156);
or U12081 (N_12081,N_10711,N_11920);
nand U12082 (N_12082,N_11432,N_11992);
or U12083 (N_12083,N_11308,N_11209);
xnor U12084 (N_12084,N_11299,N_11916);
nor U12085 (N_12085,N_11863,N_10950);
and U12086 (N_12086,N_10146,N_11125);
and U12087 (N_12087,N_10922,N_11022);
and U12088 (N_12088,N_10511,N_11890);
and U12089 (N_12089,N_11736,N_11851);
xor U12090 (N_12090,N_10925,N_10340);
xor U12091 (N_12091,N_10069,N_10768);
xor U12092 (N_12092,N_11516,N_11168);
nor U12093 (N_12093,N_11123,N_10698);
nand U12094 (N_12094,N_11552,N_10231);
or U12095 (N_12095,N_10875,N_11872);
nand U12096 (N_12096,N_10927,N_10541);
nand U12097 (N_12097,N_10832,N_10263);
xnor U12098 (N_12098,N_11926,N_11237);
or U12099 (N_12099,N_11936,N_11554);
nand U12100 (N_12100,N_11260,N_10100);
nor U12101 (N_12101,N_11899,N_11424);
nand U12102 (N_12102,N_10227,N_11082);
nand U12103 (N_12103,N_10975,N_10137);
or U12104 (N_12104,N_10173,N_11155);
and U12105 (N_12105,N_10011,N_11088);
nor U12106 (N_12106,N_10470,N_10949);
nor U12107 (N_12107,N_11225,N_11226);
nand U12108 (N_12108,N_10465,N_10192);
xnor U12109 (N_12109,N_10117,N_11881);
nor U12110 (N_12110,N_11266,N_11913);
or U12111 (N_12111,N_10632,N_10955);
or U12112 (N_12112,N_11060,N_10439);
xnor U12113 (N_12113,N_11846,N_11101);
and U12114 (N_12114,N_10361,N_11282);
or U12115 (N_12115,N_10551,N_10310);
nand U12116 (N_12116,N_11230,N_11947);
or U12117 (N_12117,N_11791,N_11000);
nand U12118 (N_12118,N_10871,N_11223);
xnor U12119 (N_12119,N_11038,N_10373);
and U12120 (N_12120,N_11519,N_11131);
nand U12121 (N_12121,N_11622,N_11759);
and U12122 (N_12122,N_11343,N_10303);
and U12123 (N_12123,N_10641,N_10544);
nand U12124 (N_12124,N_10672,N_10602);
nor U12125 (N_12125,N_11012,N_11927);
nand U12126 (N_12126,N_11385,N_10752);
xor U12127 (N_12127,N_11574,N_10585);
xor U12128 (N_12128,N_11149,N_11693);
or U12129 (N_12129,N_11109,N_10065);
nor U12130 (N_12130,N_11460,N_10469);
nor U12131 (N_12131,N_11382,N_11262);
nand U12132 (N_12132,N_11135,N_11642);
xnor U12133 (N_12133,N_11165,N_10516);
nor U12134 (N_12134,N_11268,N_10055);
nand U12135 (N_12135,N_11161,N_10054);
and U12136 (N_12136,N_11776,N_11861);
nand U12137 (N_12137,N_11429,N_11402);
or U12138 (N_12138,N_10186,N_11820);
or U12139 (N_12139,N_11443,N_10720);
and U12140 (N_12140,N_10351,N_10402);
or U12141 (N_12141,N_11528,N_10488);
or U12142 (N_12142,N_11923,N_11520);
nor U12143 (N_12143,N_10206,N_11042);
nor U12144 (N_12144,N_11632,N_11003);
nand U12145 (N_12145,N_11666,N_10512);
or U12146 (N_12146,N_11969,N_10036);
nor U12147 (N_12147,N_11758,N_10946);
nor U12148 (N_12148,N_10266,N_11120);
nor U12149 (N_12149,N_10398,N_11111);
and U12150 (N_12150,N_10221,N_10563);
xnor U12151 (N_12151,N_10387,N_11604);
xnor U12152 (N_12152,N_10847,N_11019);
and U12153 (N_12153,N_10228,N_11401);
nor U12154 (N_12154,N_10577,N_10647);
or U12155 (N_12155,N_10852,N_11811);
nand U12156 (N_12156,N_11978,N_11079);
or U12157 (N_12157,N_11321,N_10334);
nor U12158 (N_12158,N_11367,N_10778);
and U12159 (N_12159,N_10450,N_11059);
nand U12160 (N_12160,N_10658,N_10084);
nand U12161 (N_12161,N_11352,N_10893);
nor U12162 (N_12162,N_11534,N_10860);
nand U12163 (N_12163,N_10882,N_11106);
nor U12164 (N_12164,N_10558,N_10256);
nor U12165 (N_12165,N_11084,N_11681);
nand U12166 (N_12166,N_10321,N_11178);
or U12167 (N_12167,N_10670,N_10574);
nand U12168 (N_12168,N_11723,N_10410);
or U12169 (N_12169,N_11606,N_11340);
nand U12170 (N_12170,N_10330,N_11549);
or U12171 (N_12171,N_11659,N_11955);
and U12172 (N_12172,N_11097,N_11011);
nor U12173 (N_12173,N_11431,N_11005);
xor U12174 (N_12174,N_11423,N_11963);
nand U12175 (N_12175,N_11842,N_11451);
or U12176 (N_12176,N_11684,N_10111);
nor U12177 (N_12177,N_11232,N_10748);
nor U12178 (N_12178,N_11806,N_10406);
xor U12179 (N_12179,N_10456,N_11826);
and U12180 (N_12180,N_11134,N_11175);
nand U12181 (N_12181,N_11648,N_11906);
xnor U12182 (N_12182,N_10087,N_10165);
or U12183 (N_12183,N_11598,N_10663);
or U12184 (N_12184,N_10736,N_10411);
xor U12185 (N_12185,N_10845,N_11537);
or U12186 (N_12186,N_11635,N_10140);
nor U12187 (N_12187,N_10336,N_10645);
or U12188 (N_12188,N_11405,N_10322);
or U12189 (N_12189,N_10496,N_10276);
nor U12190 (N_12190,N_11983,N_10476);
and U12191 (N_12191,N_11269,N_10042);
nand U12192 (N_12192,N_10175,N_10153);
nor U12193 (N_12193,N_11347,N_11889);
or U12194 (N_12194,N_10214,N_11362);
nor U12195 (N_12195,N_11540,N_10333);
or U12196 (N_12196,N_11768,N_10265);
or U12197 (N_12197,N_11153,N_11668);
or U12198 (N_12198,N_10887,N_11695);
nand U12199 (N_12199,N_10145,N_11862);
or U12200 (N_12200,N_10854,N_11822);
or U12201 (N_12201,N_11238,N_11835);
nor U12202 (N_12202,N_11317,N_10522);
and U12203 (N_12203,N_10648,N_10855);
xnor U12204 (N_12204,N_10606,N_10564);
nand U12205 (N_12205,N_11351,N_11683);
xor U12206 (N_12206,N_10770,N_10708);
or U12207 (N_12207,N_11244,N_10444);
or U12208 (N_12208,N_11675,N_10457);
and U12209 (N_12209,N_11210,N_10918);
or U12210 (N_12210,N_10753,N_10277);
xor U12211 (N_12211,N_10188,N_11619);
and U12212 (N_12212,N_10896,N_11745);
and U12213 (N_12213,N_10834,N_10200);
nor U12214 (N_12214,N_10837,N_10939);
nor U12215 (N_12215,N_10581,N_10938);
or U12216 (N_12216,N_11102,N_10077);
nor U12217 (N_12217,N_10785,N_11322);
nand U12218 (N_12218,N_11763,N_11802);
and U12219 (N_12219,N_11037,N_10264);
and U12220 (N_12220,N_10609,N_11600);
or U12221 (N_12221,N_10814,N_10267);
or U12222 (N_12222,N_10026,N_11702);
nand U12223 (N_12223,N_11800,N_11170);
and U12224 (N_12224,N_10312,N_10682);
xnor U12225 (N_12225,N_10980,N_11620);
nand U12226 (N_12226,N_10020,N_10189);
nand U12227 (N_12227,N_10374,N_10518);
nand U12228 (N_12228,N_10381,N_10836);
and U12229 (N_12229,N_11137,N_10792);
nor U12230 (N_12230,N_11373,N_11286);
xnor U12231 (N_12231,N_10128,N_10744);
and U12232 (N_12232,N_11334,N_10363);
and U12233 (N_12233,N_10500,N_10472);
or U12234 (N_12234,N_11051,N_11199);
nor U12235 (N_12235,N_10174,N_10169);
nor U12236 (N_12236,N_10956,N_11486);
nand U12237 (N_12237,N_10123,N_11370);
nor U12238 (N_12238,N_10945,N_11187);
or U12239 (N_12239,N_10777,N_10142);
nand U12240 (N_12240,N_11293,N_10907);
nor U12241 (N_12241,N_10217,N_10515);
xnor U12242 (N_12242,N_11426,N_11463);
or U12243 (N_12243,N_11617,N_11544);
and U12244 (N_12244,N_10782,N_11787);
xnor U12245 (N_12245,N_10876,N_10879);
and U12246 (N_12246,N_11428,N_11653);
nand U12247 (N_12247,N_11345,N_11821);
xor U12248 (N_12248,N_11095,N_11510);
and U12249 (N_12249,N_10497,N_11028);
nor U12250 (N_12250,N_10828,N_10440);
and U12251 (N_12251,N_10023,N_10431);
and U12252 (N_12252,N_10684,N_11212);
nor U12253 (N_12253,N_11942,N_11314);
and U12254 (N_12254,N_11065,N_10678);
xnor U12255 (N_12255,N_10130,N_10167);
nor U12256 (N_12256,N_10304,N_10195);
nand U12257 (N_12257,N_10345,N_11836);
nor U12258 (N_12258,N_10013,N_10019);
xor U12259 (N_12259,N_10637,N_10325);
nor U12260 (N_12260,N_10316,N_10972);
nand U12261 (N_12261,N_10044,N_11246);
and U12262 (N_12262,N_11338,N_11815);
nor U12263 (N_12263,N_11179,N_11311);
nor U12264 (N_12264,N_10086,N_10232);
xor U12265 (N_12265,N_10354,N_10685);
or U12266 (N_12266,N_11609,N_10323);
nand U12267 (N_12267,N_10234,N_11289);
nor U12268 (N_12268,N_10717,N_11922);
and U12269 (N_12269,N_10491,N_11180);
and U12270 (N_12270,N_10700,N_11816);
xnor U12271 (N_12271,N_10244,N_11208);
nand U12272 (N_12272,N_10788,N_10817);
and U12273 (N_12273,N_11336,N_11096);
nand U12274 (N_12274,N_11928,N_10041);
xnor U12275 (N_12275,N_11613,N_11172);
nor U12276 (N_12276,N_10908,N_11018);
nand U12277 (N_12277,N_10001,N_11738);
nand U12278 (N_12278,N_10954,N_10403);
and U12279 (N_12279,N_10301,N_10668);
or U12280 (N_12280,N_10568,N_10487);
or U12281 (N_12281,N_11368,N_10358);
nand U12282 (N_12282,N_10029,N_10953);
or U12283 (N_12283,N_10249,N_11403);
xor U12284 (N_12284,N_11784,N_10969);
or U12285 (N_12285,N_11739,N_11183);
nand U12286 (N_12286,N_10957,N_11631);
or U12287 (N_12287,N_11522,N_10935);
nor U12288 (N_12288,N_11421,N_10447);
and U12289 (N_12289,N_10521,N_10058);
nor U12290 (N_12290,N_10126,N_10937);
nand U12291 (N_12291,N_11680,N_10095);
nor U12292 (N_12292,N_10735,N_10166);
nand U12293 (N_12293,N_11457,N_10343);
and U12294 (N_12294,N_10547,N_10014);
nor U12295 (N_12295,N_11017,N_11960);
or U12296 (N_12296,N_10375,N_11177);
nand U12297 (N_12297,N_11895,N_11091);
xor U12298 (N_12298,N_10176,N_10160);
and U12299 (N_12299,N_11227,N_11742);
and U12300 (N_12300,N_11450,N_10884);
or U12301 (N_12301,N_10125,N_11182);
nor U12302 (N_12302,N_11535,N_10508);
and U12303 (N_12303,N_10962,N_11977);
xor U12304 (N_12304,N_11350,N_10833);
nor U12305 (N_12305,N_10034,N_10618);
nor U12306 (N_12306,N_11744,N_11917);
nand U12307 (N_12307,N_11792,N_10634);
or U12308 (N_12308,N_11594,N_10288);
nand U12309 (N_12309,N_11686,N_10493);
xnor U12310 (N_12310,N_11302,N_10548);
or U12311 (N_12311,N_11303,N_10921);
and U12312 (N_12312,N_10215,N_11229);
xnor U12313 (N_12313,N_11276,N_11687);
xnor U12314 (N_12314,N_11435,N_10791);
xnor U12315 (N_12315,N_10572,N_11407);
nand U12316 (N_12316,N_11892,N_10138);
nor U12317 (N_12317,N_11638,N_11053);
nor U12318 (N_12318,N_10870,N_11393);
and U12319 (N_12319,N_11650,N_10886);
xnor U12320 (N_12320,N_11730,N_10317);
nand U12321 (N_12321,N_11797,N_11640);
xor U12322 (N_12322,N_11961,N_10046);
or U12323 (N_12323,N_11389,N_10262);
nand U12324 (N_12324,N_11869,N_10897);
xnor U12325 (N_12325,N_10012,N_11985);
nand U12326 (N_12326,N_11214,N_11691);
and U12327 (N_12327,N_10342,N_11581);
or U12328 (N_12328,N_11310,N_10112);
nand U12329 (N_12329,N_11838,N_11419);
xnor U12330 (N_12330,N_10484,N_10434);
or U12331 (N_12331,N_11092,N_10693);
nor U12332 (N_12332,N_10480,N_10449);
nand U12333 (N_12333,N_10164,N_10948);
nand U12334 (N_12334,N_10666,N_10830);
nor U12335 (N_12335,N_10070,N_11562);
and U12336 (N_12336,N_10218,N_11422);
nor U12337 (N_12337,N_10526,N_11551);
and U12338 (N_12338,N_10766,N_11318);
nand U12339 (N_12339,N_10525,N_10096);
nand U12340 (N_12340,N_10566,N_10024);
nor U12341 (N_12341,N_11470,N_10677);
and U12342 (N_12342,N_11476,N_11664);
xnor U12343 (N_12343,N_11848,N_10229);
xor U12344 (N_12344,N_10073,N_10857);
or U12345 (N_12345,N_11396,N_11773);
nand U12346 (N_12346,N_10669,N_10543);
or U12347 (N_12347,N_11628,N_10813);
nand U12348 (N_12348,N_11381,N_10755);
xnor U12349 (N_12349,N_10540,N_10005);
xor U12350 (N_12350,N_10616,N_10710);
or U12351 (N_12351,N_10513,N_10798);
nand U12352 (N_12352,N_11957,N_11271);
nor U12353 (N_12353,N_11025,N_10831);
nand U12354 (N_12354,N_11387,N_10580);
or U12355 (N_12355,N_11943,N_11697);
and U12356 (N_12356,N_11900,N_10261);
xnor U12357 (N_12357,N_10062,N_11312);
xnor U12358 (N_12358,N_11860,N_10437);
or U12359 (N_12359,N_11538,N_11727);
nand U12360 (N_12360,N_11678,N_11258);
nand U12361 (N_12361,N_10492,N_11786);
xnor U12362 (N_12362,N_11867,N_10453);
nand U12363 (N_12363,N_11305,N_10461);
nor U12364 (N_12364,N_11277,N_11555);
xor U12365 (N_12365,N_10253,N_10210);
and U12366 (N_12366,N_11205,N_10995);
xnor U12367 (N_12367,N_11883,N_11337);
and U12368 (N_12368,N_10797,N_10846);
or U12369 (N_12369,N_10066,N_11532);
nand U12370 (N_12370,N_10978,N_10279);
or U12371 (N_12371,N_11840,N_10356);
nand U12372 (N_12372,N_11414,N_10425);
or U12373 (N_12373,N_11970,N_10102);
or U12374 (N_12374,N_10360,N_11708);
nand U12375 (N_12375,N_10162,N_11918);
nand U12376 (N_12376,N_11254,N_11563);
or U12377 (N_12377,N_11855,N_10756);
or U12378 (N_12378,N_10101,N_11694);
and U12379 (N_12379,N_11805,N_11548);
nand U12380 (N_12380,N_11626,N_11796);
nor U12381 (N_12381,N_11601,N_10659);
nand U12382 (N_12382,N_11794,N_10287);
xnor U12383 (N_12383,N_11831,N_11643);
nor U12384 (N_12384,N_11854,N_10584);
nand U12385 (N_12385,N_10459,N_11795);
nand U12386 (N_12386,N_10517,N_11560);
or U12387 (N_12387,N_10092,N_10865);
and U12388 (N_12388,N_10789,N_11026);
or U12389 (N_12389,N_10399,N_11339);
nand U12390 (N_12390,N_10239,N_11886);
and U12391 (N_12391,N_10691,N_10074);
nor U12392 (N_12392,N_10419,N_11220);
nor U12393 (N_12393,N_11406,N_10180);
nor U12394 (N_12394,N_10794,N_10751);
and U12395 (N_12395,N_10369,N_11112);
and U12396 (N_12396,N_11843,N_11163);
nand U12397 (N_12397,N_10331,N_11912);
and U12398 (N_12398,N_11394,N_10219);
nor U12399 (N_12399,N_11441,N_11188);
nand U12400 (N_12400,N_11754,N_10254);
xnor U12401 (N_12401,N_11094,N_11243);
xor U12402 (N_12402,N_11756,N_10660);
and U12403 (N_12403,N_10926,N_11715);
and U12404 (N_12404,N_11479,N_10097);
or U12405 (N_12405,N_10635,N_10308);
nand U12406 (N_12406,N_10467,N_10626);
or U12407 (N_12407,N_11201,N_11901);
nand U12408 (N_12408,N_11909,N_10981);
or U12409 (N_12409,N_10850,N_10815);
and U12410 (N_12410,N_10844,N_10204);
or U12411 (N_12411,N_10652,N_11817);
or U12412 (N_12412,N_10082,N_11481);
nor U12413 (N_12413,N_10201,N_10233);
xor U12414 (N_12414,N_11875,N_10392);
or U12415 (N_12415,N_11915,N_10536);
nor U12416 (N_12416,N_11893,N_10786);
or U12417 (N_12417,N_10801,N_11571);
and U12418 (N_12418,N_11436,N_10429);
nor U12419 (N_12419,N_11329,N_11705);
nand U12420 (N_12420,N_10455,N_10018);
xor U12421 (N_12421,N_11769,N_11075);
xor U12422 (N_12422,N_11124,N_11716);
xnor U12423 (N_12423,N_11072,N_11722);
or U12424 (N_12424,N_11965,N_11703);
or U12425 (N_12425,N_11050,N_10839);
nand U12426 (N_12426,N_11068,N_10826);
or U12427 (N_12427,N_10732,N_10527);
nor U12428 (N_12428,N_11767,N_10104);
nand U12429 (N_12429,N_11195,N_11793);
and U12430 (N_12430,N_10305,N_11315);
xnor U12431 (N_12431,N_11743,N_10902);
xnor U12432 (N_12432,N_11981,N_10339);
or U12433 (N_12433,N_11570,N_10905);
xor U12434 (N_12434,N_11935,N_11319);
nor U12435 (N_12435,N_10901,N_11625);
xnor U12436 (N_12436,N_11133,N_11234);
and U12437 (N_12437,N_10157,N_10724);
nor U12438 (N_12438,N_11627,N_11719);
nor U12439 (N_12439,N_10567,N_10498);
or U12440 (N_12440,N_10979,N_10413);
xnor U12441 (N_12441,N_10929,N_11029);
or U12442 (N_12442,N_11231,N_11189);
xnor U12443 (N_12443,N_11192,N_11378);
or U12444 (N_12444,N_10235,N_11894);
xnor U12445 (N_12445,N_11056,N_11568);
xor U12446 (N_12446,N_10390,N_10795);
nor U12447 (N_12447,N_10835,N_11449);
nand U12448 (N_12448,N_11607,N_11500);
or U12449 (N_12449,N_10594,N_11996);
and U12450 (N_12450,N_11509,N_11046);
and U12451 (N_12451,N_11902,N_10947);
nand U12452 (N_12452,N_11866,N_11228);
or U12453 (N_12453,N_11434,N_11365);
or U12454 (N_12454,N_11704,N_10627);
nand U12455 (N_12455,N_11062,N_10393);
nor U12456 (N_12456,N_11993,N_11966);
and U12457 (N_12457,N_10885,N_11278);
nor U12458 (N_12458,N_11785,N_10273);
nor U12459 (N_12459,N_11602,N_11033);
nor U12460 (N_12460,N_10190,N_10783);
xnor U12461 (N_12461,N_11328,N_10478);
or U12462 (N_12462,N_11749,N_11342);
or U12463 (N_12463,N_10395,N_11647);
xor U12464 (N_12464,N_10750,N_10213);
xnor U12465 (N_12465,N_10426,N_11774);
nand U12466 (N_12466,N_10990,N_11433);
nand U12467 (N_12467,N_11215,N_11873);
or U12468 (N_12468,N_11386,N_11651);
nand U12469 (N_12469,N_10282,N_10076);
nand U12470 (N_12470,N_10533,N_11780);
nand U12471 (N_12471,N_10621,N_10984);
or U12472 (N_12472,N_11397,N_10386);
or U12473 (N_12473,N_10730,N_11444);
nor U12474 (N_12474,N_11255,N_10328);
and U12475 (N_12475,N_11275,N_11972);
nor U12476 (N_12476,N_11185,N_11986);
and U12477 (N_12477,N_10983,N_10132);
nor U12478 (N_12478,N_11071,N_10445);
and U12479 (N_12479,N_10964,N_11020);
or U12480 (N_12480,N_11770,N_11331);
xor U12481 (N_12481,N_11100,N_11973);
and U12482 (N_12482,N_11371,N_10881);
nor U12483 (N_12483,N_11982,N_10623);
nand U12484 (N_12484,N_11559,N_11790);
and U12485 (N_12485,N_11504,N_10630);
or U12486 (N_12486,N_11764,N_11203);
xor U12487 (N_12487,N_10519,N_10904);
or U12488 (N_12488,N_11462,N_11924);
nand U12489 (N_12489,N_10129,N_11948);
and U12490 (N_12490,N_11655,N_11914);
or U12491 (N_12491,N_10355,N_11021);
xnor U12492 (N_12492,N_11250,N_11484);
or U12493 (N_12493,N_10209,N_11176);
nand U12494 (N_12494,N_11066,N_10963);
nand U12495 (N_12495,N_11143,N_10614);
nor U12496 (N_12496,N_11533,N_11596);
nor U12497 (N_12497,N_11610,N_10805);
xor U12498 (N_12498,N_11253,N_11248);
nor U12499 (N_12499,N_10890,N_10827);
or U12500 (N_12500,N_10349,N_10368);
or U12501 (N_12501,N_11523,N_11849);
or U12502 (N_12502,N_11939,N_11698);
nand U12503 (N_12503,N_11313,N_11633);
nor U12504 (N_12504,N_10787,N_10799);
xor U12505 (N_12505,N_11556,N_11921);
xnor U12506 (N_12506,N_10237,N_10269);
xor U12507 (N_12507,N_11747,N_10848);
nor U12508 (N_12508,N_10052,N_10631);
nor U12509 (N_12509,N_11296,N_10576);
and U12510 (N_12510,N_11292,N_10382);
and U12511 (N_12511,N_10593,N_10713);
nor U12512 (N_12512,N_10141,N_11440);
nor U12513 (N_12513,N_11761,N_11827);
xor U12514 (N_12514,N_10091,N_10286);
nand U12515 (N_12515,N_10552,N_10207);
nor U12516 (N_12516,N_10808,N_11724);
and U12517 (N_12517,N_11788,N_11304);
nor U12518 (N_12518,N_11578,N_10458);
nor U12519 (N_12519,N_11122,N_10407);
nand U12520 (N_12520,N_11597,N_11058);
and U12521 (N_12521,N_10679,N_10477);
nor U12522 (N_12522,N_10376,N_11202);
nand U12523 (N_12523,N_10337,N_10171);
nor U12524 (N_12524,N_11591,N_11823);
nand U12525 (N_12525,N_10706,N_11455);
or U12526 (N_12526,N_11765,N_10415);
and U12527 (N_12527,N_10412,N_11380);
nor U12528 (N_12528,N_11987,N_11689);
nand U12529 (N_12529,N_11471,N_10598);
nor U12530 (N_12530,N_10313,N_10454);
xor U12531 (N_12531,N_10113,N_11007);
nand U12532 (N_12532,N_10639,N_10628);
and U12533 (N_12533,N_11819,N_10346);
or U12534 (N_12534,N_11850,N_11839);
or U12535 (N_12535,N_10531,N_11667);
or U12536 (N_12536,N_10873,N_11151);
and U12537 (N_12537,N_11905,N_10638);
nand U12538 (N_12538,N_10428,N_10452);
xor U12539 (N_12539,N_10622,N_10589);
xnor U12540 (N_12540,N_10037,N_10941);
or U12541 (N_12541,N_11472,N_10017);
and U12542 (N_12542,N_10661,N_10243);
nor U12543 (N_12543,N_11356,N_10681);
nor U12544 (N_12544,N_11585,N_10320);
nor U12545 (N_12545,N_10043,N_11469);
nor U12546 (N_12546,N_10260,N_10985);
nand U12547 (N_12547,N_10721,N_10781);
or U12548 (N_12548,N_10191,N_10915);
xor U12549 (N_12549,N_11494,N_11014);
nor U12550 (N_12550,N_10867,N_10704);
or U12551 (N_12551,N_10357,N_10633);
xor U12552 (N_12552,N_10600,N_11288);
nor U12553 (N_12553,N_10542,N_11636);
nand U12554 (N_12554,N_11644,N_10579);
or U12555 (N_12555,N_11045,N_10804);
or U12556 (N_12556,N_11270,N_11879);
nand U12557 (N_12557,N_10423,N_11498);
nor U12558 (N_12558,N_10223,N_10583);
nand U12559 (N_12559,N_10274,N_11711);
nand U12560 (N_12560,N_10422,N_10520);
or U12561 (N_12561,N_10003,N_10874);
nand U12562 (N_12562,N_11575,N_11663);
and U12563 (N_12563,N_11959,N_10654);
and U12564 (N_12564,N_11573,N_11040);
and U12565 (N_12565,N_10977,N_11291);
or U12566 (N_12566,N_11259,N_11565);
or U12567 (N_12567,N_10643,N_10996);
nor U12568 (N_12568,N_11662,N_10341);
xor U12569 (N_12569,N_10872,N_10420);
nor U12570 (N_12570,N_10967,N_10919);
xnor U12571 (N_12571,N_10462,N_11503);
nor U12572 (N_12572,N_10106,N_10562);
and U12573 (N_12573,N_11852,N_10676);
nand U12574 (N_12574,N_10578,N_11824);
nand U12575 (N_12575,N_10035,N_11750);
nor U12576 (N_12576,N_11355,N_10898);
or U12577 (N_12577,N_10992,N_10546);
xor U12578 (N_12578,N_10644,N_10912);
nor U12579 (N_12579,N_11105,N_11771);
or U12580 (N_12580,N_11507,N_10432);
or U12581 (N_12581,N_10383,N_10098);
nand U12582 (N_12582,N_10107,N_11333);
or U12583 (N_12583,N_11039,N_10203);
or U12584 (N_12584,N_11649,N_10959);
nand U12585 (N_12585,N_11944,N_11713);
and U12586 (N_12586,N_11139,N_10212);
nand U12587 (N_12587,N_11710,N_10482);
nor U12588 (N_12588,N_11654,N_11236);
xnor U12589 (N_12589,N_10197,N_10247);
nor U12590 (N_12590,N_10771,N_11502);
nand U12591 (N_12591,N_10725,N_11297);
nand U12592 (N_12592,N_11218,N_11264);
xnor U12593 (N_12593,N_11542,N_10976);
xor U12594 (N_12594,N_11512,N_11006);
nor U12595 (N_12595,N_10575,N_11144);
xor U12596 (N_12596,N_10025,N_11833);
and U12597 (N_12597,N_11729,N_11778);
or U12598 (N_12598,N_11964,N_10481);
and U12599 (N_12599,N_10168,N_10779);
or U12600 (N_12600,N_11968,N_10534);
xnor U12601 (N_12601,N_10754,N_11152);
xnor U12602 (N_12602,N_11870,N_10920);
or U12603 (N_12603,N_11354,N_10769);
and U12604 (N_12604,N_11882,N_10430);
and U12605 (N_12605,N_10424,N_11061);
xnor U12606 (N_12606,N_11971,N_10810);
or U12607 (N_12607,N_11353,N_11466);
nand U12608 (N_12608,N_10767,N_11593);
xor U12609 (N_12609,N_11897,N_11717);
and U12610 (N_12610,N_11344,N_10255);
nor U12611 (N_12611,N_11330,N_10952);
xor U12612 (N_12612,N_10712,N_11430);
and U12613 (N_12613,N_10490,N_11164);
xor U12614 (N_12614,N_10673,N_10692);
nor U12615 (N_12615,N_11398,N_10246);
xnor U12616 (N_12616,N_11416,N_11015);
nand U12617 (N_12617,N_10078,N_10559);
xnor U12618 (N_12618,N_11999,N_10371);
and U12619 (N_12619,N_11527,N_10033);
nor U12620 (N_12620,N_10707,N_11147);
nor U12621 (N_12621,N_10757,N_11804);
and U12622 (N_12622,N_11196,N_10093);
nand U12623 (N_12623,N_11290,N_10841);
or U12624 (N_12624,N_11903,N_11464);
or U12625 (N_12625,N_11217,N_11263);
nand U12626 (N_12626,N_10888,N_10414);
and U12627 (N_12627,N_10726,N_10495);
nor U12628 (N_12628,N_10284,N_10268);
xor U12629 (N_12629,N_11775,N_10009);
or U12630 (N_12630,N_11145,N_11646);
nand U12631 (N_12631,N_11492,N_11247);
and U12632 (N_12632,N_11207,N_10943);
and U12633 (N_12633,N_10194,N_11358);
nor U12634 (N_12634,N_10994,N_10951);
xor U12635 (N_12635,N_10858,N_10690);
nor U12636 (N_12636,N_11725,N_10451);
nor U12637 (N_12637,N_11272,N_10982);
xnor U12638 (N_12638,N_11044,N_11907);
and U12639 (N_12639,N_10746,N_10615);
xor U12640 (N_12640,N_10966,N_10793);
and U12641 (N_12641,N_11408,N_11910);
nand U12642 (N_12642,N_10418,N_10958);
xnor U12643 (N_12643,N_11989,N_10022);
and U12644 (N_12644,N_10198,N_10582);
and U12645 (N_12645,N_10002,N_10134);
or U12646 (N_12646,N_10021,N_10385);
xnor U12647 (N_12647,N_11265,N_11904);
xor U12648 (N_12648,N_10611,N_10259);
nor U12649 (N_12649,N_11415,N_11024);
nand U12650 (N_12650,N_10557,N_11233);
xor U12651 (N_12651,N_10238,N_10936);
xnor U12652 (N_12652,N_10586,N_11335);
nand U12653 (N_12653,N_10999,N_10932);
or U12654 (N_12654,N_10299,N_11036);
or U12655 (N_12655,N_11475,N_10965);
and U12656 (N_12656,N_10765,N_11174);
and U12657 (N_12657,N_10103,N_11665);
nand U12658 (N_12658,N_10039,N_10258);
xor U12659 (N_12659,N_10702,N_10853);
nor U12660 (N_12660,N_11023,N_10090);
nor U12661 (N_12661,N_11118,N_10840);
nand U12662 (N_12662,N_11834,N_10155);
xnor U12663 (N_12663,N_11103,N_11940);
and U12664 (N_12664,N_10530,N_10776);
nor U12665 (N_12665,N_11009,N_10281);
nand U12666 (N_12666,N_10961,N_11173);
xor U12667 (N_12667,N_11731,N_10057);
nand U12668 (N_12668,N_10539,N_10532);
and U12669 (N_12669,N_10662,N_11865);
nand U12670 (N_12670,N_10524,N_11728);
nand U12671 (N_12671,N_11699,N_11198);
nand U12672 (N_12672,N_10147,N_11813);
nand U12673 (N_12673,N_10088,N_11976);
xor U12674 (N_12674,N_10913,N_10332);
or U12675 (N_12675,N_11709,N_10619);
or U12676 (N_12676,N_11309,N_10245);
nand U12677 (N_12677,N_10348,N_10716);
and U12678 (N_12678,N_10220,N_11589);
or U12679 (N_12679,N_11047,N_10914);
nor U12680 (N_12680,N_10818,N_11332);
and U12681 (N_12681,N_10202,N_11952);
xnor U12682 (N_12682,N_11857,N_11369);
xnor U12683 (N_12683,N_10745,N_10705);
or U12684 (N_12684,N_10974,N_10471);
and U12685 (N_12685,N_11934,N_11349);
and U12686 (N_12686,N_11461,N_10473);
nor U12687 (N_12687,N_10441,N_11974);
nor U12688 (N_12688,N_11515,N_10079);
xor U12689 (N_12689,N_10257,N_10050);
and U12690 (N_12690,N_11366,N_10061);
or U12691 (N_12691,N_10122,N_10636);
xor U12692 (N_12692,N_11789,N_11108);
and U12693 (N_12693,N_10226,N_11298);
and U12694 (N_12694,N_10466,N_10931);
xor U12695 (N_12695,N_11696,N_11438);
xor U12696 (N_12696,N_11048,N_10565);
nor U12697 (N_12697,N_11454,N_10295);
nor U12698 (N_12698,N_11064,N_11035);
and U12699 (N_12699,N_10314,N_11735);
xor U12700 (N_12700,N_11830,N_11488);
xnor U12701 (N_12701,N_10780,N_11437);
or U12702 (N_12702,N_11692,N_11081);
nand U12703 (N_12703,N_10010,N_10380);
xor U12704 (N_12704,N_10802,N_10733);
and U12705 (N_12705,N_10183,N_10655);
xor U12706 (N_12706,N_10293,N_10820);
or U12707 (N_12707,N_10667,N_11513);
xnor U12708 (N_12708,N_11425,N_10821);
nand U12709 (N_12709,N_10760,N_10278);
xnor U12710 (N_12710,N_10127,N_11858);
and U12711 (N_12711,N_11400,N_11013);
or U12712 (N_12712,N_10135,N_10417);
or U12713 (N_12713,N_10800,N_10347);
nand U12714 (N_12714,N_10822,N_11614);
nand U12715 (N_12715,N_11306,N_11295);
nor U12716 (N_12716,N_10699,N_11074);
or U12717 (N_12717,N_10463,N_11107);
nand U12718 (N_12718,N_11733,N_10665);
and U12719 (N_12719,N_10997,N_11737);
and U12720 (N_12720,N_10152,N_10599);
and U12721 (N_12721,N_10120,N_11930);
nand U12722 (N_12722,N_11239,N_11245);
and U12723 (N_12723,N_11720,N_10729);
nor U12724 (N_12724,N_11931,N_11204);
and U12725 (N_12725,N_11452,N_11224);
nand U12726 (N_12726,N_11518,N_11395);
and U12727 (N_12727,N_11937,N_10696);
nand U12728 (N_12728,N_10409,N_11547);
nand U12729 (N_12729,N_10910,N_10774);
nor U12730 (N_12730,N_11445,N_11740);
or U12731 (N_12731,N_10105,N_10971);
or U12732 (N_12732,N_10251,N_11132);
nand U12733 (N_12733,N_11721,N_11637);
nor U12734 (N_12734,N_11701,N_10004);
or U12735 (N_12735,N_11639,N_11929);
or U12736 (N_12736,N_11877,N_10494);
xor U12737 (N_12737,N_11281,N_10714);
and U12738 (N_12738,N_10911,N_11030);
or U12739 (N_12739,N_11671,N_10028);
or U12740 (N_12740,N_10523,N_11279);
nor U12741 (N_12741,N_10384,N_10764);
nand U12742 (N_12742,N_10686,N_10185);
or U12743 (N_12743,N_10182,N_10761);
and U12744 (N_12744,N_10159,N_10051);
nand U12745 (N_12745,N_10674,N_11676);
nand U12746 (N_12746,N_10224,N_11031);
xnor U12747 (N_12747,N_11925,N_11219);
nand U12748 (N_12748,N_10124,N_10624);
xor U12749 (N_12749,N_11517,N_10027);
and U12750 (N_12750,N_11055,N_10556);
and U12751 (N_12751,N_10877,N_11240);
nor U12752 (N_12752,N_11569,N_11384);
and U12753 (N_12753,N_11577,N_10030);
nor U12754 (N_12754,N_11967,N_11949);
nand U12755 (N_12755,N_11388,N_11377);
or U12756 (N_12756,N_10806,N_11190);
or U12757 (N_12757,N_10404,N_10156);
nand U12758 (N_12758,N_10352,N_10784);
nor U12759 (N_12759,N_11508,N_11411);
or U12760 (N_12760,N_10502,N_10285);
xnor U12761 (N_12761,N_10485,N_10006);
xor U12762 (N_12762,N_10475,N_10049);
or U12763 (N_12763,N_10075,N_10099);
and U12764 (N_12764,N_11798,N_11200);
nor U12765 (N_12765,N_10590,N_10608);
nand U12766 (N_12766,N_10319,N_11448);
and U12767 (N_12767,N_11656,N_11781);
or U12768 (N_12768,N_11249,N_10080);
xnor U12769 (N_12769,N_11446,N_11158);
xnor U12770 (N_12770,N_11624,N_11988);
nand U12771 (N_12771,N_10338,N_10772);
xnor U12772 (N_12772,N_10158,N_10446);
and U12773 (N_12773,N_10408,N_11529);
nand U12774 (N_12774,N_11032,N_10843);
xnor U12775 (N_12775,N_11480,N_11612);
nor U12776 (N_12776,N_10143,N_10015);
and U12777 (N_12777,N_10464,N_10688);
or U12778 (N_12778,N_11660,N_11553);
xnor U12779 (N_12779,N_11285,N_10236);
nand U12780 (N_12780,N_11073,N_10895);
nor U12781 (N_12781,N_11148,N_10740);
and U12782 (N_12782,N_10150,N_11859);
nand U12783 (N_12783,N_11483,N_11564);
and U12784 (N_12784,N_11946,N_11167);
nand U12785 (N_12785,N_10550,N_10909);
nand U12786 (N_12786,N_10300,N_10110);
or U12787 (N_12787,N_11726,N_10722);
and U12788 (N_12788,N_10738,N_10193);
and U12789 (N_12789,N_11887,N_11634);
and U12790 (N_12790,N_11812,N_11184);
nand U12791 (N_12791,N_11294,N_10184);
or U12792 (N_12792,N_11076,N_10829);
and U12793 (N_12793,N_11115,N_10222);
nand U12794 (N_12794,N_10172,N_10116);
xor U12795 (N_12795,N_10998,N_11324);
and U12796 (N_12796,N_10715,N_10045);
nand U12797 (N_12797,N_10448,N_10400);
or U12798 (N_12798,N_11359,N_10085);
nor U12799 (N_12799,N_11162,N_11583);
and U12800 (N_12800,N_10056,N_11803);
nor U12801 (N_12801,N_10514,N_11809);
and U12802 (N_12802,N_11718,N_10397);
nand U12803 (N_12803,N_11307,N_10486);
or U12804 (N_12804,N_10394,N_11630);
nand U12805 (N_12805,N_10047,N_11751);
or U12806 (N_12806,N_10290,N_11618);
nand U12807 (N_12807,N_11984,N_11439);
nand U12808 (N_12808,N_10108,N_10747);
xor U12809 (N_12809,N_11090,N_10063);
and U12810 (N_12810,N_11536,N_10934);
nand U12811 (N_12811,N_10081,N_11364);
and U12812 (N_12812,N_11499,N_11572);
nand U12813 (N_12813,N_10059,N_11008);
nand U12814 (N_12814,N_11049,N_11757);
xor U12815 (N_12815,N_11489,N_11994);
and U12816 (N_12816,N_11052,N_10803);
xor U12817 (N_12817,N_10587,N_10894);
and U12818 (N_12818,N_10591,N_10177);
and U12819 (N_12819,N_11417,N_11213);
and U12820 (N_12820,N_11325,N_11592);
nor U12821 (N_12821,N_11543,N_11746);
or U12822 (N_12822,N_10535,N_10366);
or U12823 (N_12823,N_11962,N_10187);
nor U12824 (N_12824,N_11099,N_10170);
or U12825 (N_12825,N_10506,N_11599);
and U12826 (N_12826,N_11458,N_10329);
nor U12827 (N_12827,N_10489,N_10538);
nor U12828 (N_12828,N_11372,N_11808);
and U12829 (N_12829,N_11531,N_11501);
nand U12830 (N_12830,N_11951,N_11027);
nand U12831 (N_12831,N_11975,N_11468);
or U12832 (N_12832,N_10359,N_10743);
xnor U12833 (N_12833,N_10866,N_10294);
and U12834 (N_12834,N_10280,N_10924);
and U12835 (N_12835,N_11004,N_11077);
or U12836 (N_12836,N_11078,N_10796);
xnor U12837 (N_12837,N_11399,N_10862);
xnor U12838 (N_12838,N_11876,N_10230);
and U12839 (N_12839,N_10275,N_10891);
or U12840 (N_12840,N_10199,N_10759);
and U12841 (N_12841,N_11818,N_10283);
xor U12842 (N_12842,N_11979,N_10211);
nand U12843 (N_12843,N_11841,N_11685);
or U12844 (N_12844,N_10528,N_10163);
and U12845 (N_12845,N_10315,N_11958);
nor U12846 (N_12846,N_10916,N_10388);
nand U12847 (N_12847,N_10701,N_11087);
nand U12848 (N_12848,N_10758,N_11413);
and U12849 (N_12849,N_11524,N_11657);
and U12850 (N_12850,N_10592,N_11222);
and U12851 (N_12851,N_10121,N_10326);
and U12852 (N_12852,N_11652,N_11525);
nand U12853 (N_12853,N_11561,N_11083);
nor U12854 (N_12854,N_11128,N_11880);
and U12855 (N_12855,N_10809,N_10307);
nor U12856 (N_12856,N_11280,N_11615);
nand U12857 (N_12857,N_11016,N_11998);
nor U12858 (N_12858,N_10889,N_11063);
and U12859 (N_12859,N_10309,N_10292);
xor U12860 (N_12860,N_10154,N_10181);
and U12861 (N_12861,N_11375,N_10892);
nor U12862 (N_12862,N_11054,N_11760);
and U12863 (N_12863,N_11491,N_11645);
nor U12864 (N_12864,N_11194,N_11779);
or U12865 (N_12865,N_10344,N_11093);
xor U12866 (N_12866,N_11283,N_11002);
nor U12867 (N_12867,N_11814,N_11363);
or U12868 (N_12868,N_11261,N_11473);
or U12869 (N_12869,N_10553,N_11390);
nand U12870 (N_12870,N_10031,N_11997);
xor U12871 (N_12871,N_11828,N_10503);
nor U12872 (N_12872,N_11274,N_10362);
xor U12873 (N_12873,N_11113,N_11898);
xnor U12874 (N_12874,N_11409,N_11216);
nand U12875 (N_12875,N_11911,N_11169);
xnor U12876 (N_12876,N_11146,N_10296);
and U12877 (N_12877,N_10604,N_10016);
and U12878 (N_12878,N_10318,N_10709);
or U12879 (N_12879,N_10649,N_10588);
nor U12880 (N_12880,N_11844,N_11956);
or U12881 (N_12881,N_11539,N_11832);
or U12882 (N_12882,N_11530,N_11541);
nor U12883 (N_12883,N_10327,N_11545);
nand U12884 (N_12884,N_10595,N_10008);
nand U12885 (N_12885,N_10824,N_11954);
nor U12886 (N_12886,N_10094,N_11566);
xor U12887 (N_12887,N_11829,N_11783);
nor U12888 (N_12888,N_10842,N_10689);
or U12889 (N_12889,N_10651,N_11418);
nor U12890 (N_12890,N_11980,N_11121);
and U12891 (N_12891,N_11496,N_11582);
and U12892 (N_12892,N_11588,N_10656);
nor U12893 (N_12893,N_10763,N_10664);
nand U12894 (N_12894,N_10109,N_11871);
and U12895 (N_12895,N_10083,N_11442);
xor U12896 (N_12896,N_10240,N_11766);
xnor U12897 (N_12897,N_11034,N_11707);
xnor U12898 (N_12898,N_11252,N_11300);
nand U12899 (N_12899,N_11256,N_11420);
and U12900 (N_12900,N_10968,N_11490);
xnor U12901 (N_12901,N_10859,N_10612);
and U12902 (N_12902,N_11608,N_10930);
nor U12903 (N_12903,N_11487,N_10917);
nor U12904 (N_12904,N_11799,N_11868);
and U12905 (N_12905,N_11080,N_10762);
nand U12906 (N_12906,N_10396,N_11067);
and U12907 (N_12907,N_11242,N_11447);
nand U12908 (N_12908,N_11140,N_10529);
or U12909 (N_12909,N_10509,N_10861);
or U12910 (N_12910,N_11919,N_11284);
xnor U12911 (N_12911,N_10718,N_10139);
xnor U12912 (N_12912,N_10970,N_10289);
or U12913 (N_12913,N_11316,N_10940);
nor U12914 (N_12914,N_10067,N_11990);
nor U12915 (N_12915,N_10241,N_11206);
or U12916 (N_12916,N_11085,N_10370);
and U12917 (N_12917,N_10499,N_11837);
xor U12918 (N_12918,N_10973,N_10734);
or U12919 (N_12919,N_10703,N_11142);
and U12920 (N_12920,N_11404,N_10773);
xor U12921 (N_12921,N_10899,N_10605);
xnor U12922 (N_12922,N_10868,N_10560);
or U12923 (N_12923,N_10372,N_10942);
or U12924 (N_12924,N_10483,N_11098);
or U12925 (N_12925,N_11810,N_10416);
or U12926 (N_12926,N_10863,N_11412);
or U12927 (N_12927,N_11732,N_10405);
and U12928 (N_12928,N_10807,N_11392);
and U12929 (N_12929,N_11950,N_11845);
xor U12930 (N_12930,N_11410,N_10864);
nor U12931 (N_12931,N_10988,N_10687);
nand U12932 (N_12932,N_11847,N_11320);
nor U12933 (N_12933,N_11497,N_10960);
and U12934 (N_12934,N_10151,N_11752);
nor U12935 (N_12935,N_11267,N_11888);
and U12936 (N_12936,N_11482,N_11057);
nand U12937 (N_12937,N_11391,N_10306);
nand U12938 (N_12938,N_10270,N_11953);
nand U12939 (N_12939,N_11171,N_11506);
nor U12940 (N_12940,N_10880,N_10353);
xor U12941 (N_12941,N_10072,N_11119);
and U12942 (N_12942,N_10555,N_10680);
nor U12943 (N_12943,N_11348,N_10378);
and U12944 (N_12944,N_11595,N_10297);
nor U12945 (N_12945,N_10196,N_10311);
nor U12946 (N_12946,N_10443,N_10597);
or U12947 (N_12947,N_11287,N_10601);
and U12948 (N_12948,N_11853,N_10816);
nand U12949 (N_12949,N_10474,N_10161);
or U12950 (N_12950,N_10640,N_11587);
xor U12951 (N_12951,N_10610,N_10838);
nor U12952 (N_12952,N_11326,N_11933);
nand U12953 (N_12953,N_11945,N_10250);
nand U12954 (N_12954,N_10208,N_10225);
nand U12955 (N_12955,N_11550,N_11514);
xnor U12956 (N_12956,N_10133,N_11360);
and U12957 (N_12957,N_11941,N_11864);
or U12958 (N_12958,N_10507,N_10007);
nand U12959 (N_12959,N_11938,N_11874);
nand U12960 (N_12960,N_11114,N_10053);
nand U12961 (N_12961,N_11251,N_10119);
nand U12962 (N_12962,N_10038,N_10302);
nor U12963 (N_12963,N_10851,N_10653);
and U12964 (N_12964,N_11741,N_10131);
or U12965 (N_12965,N_11772,N_10048);
nor U12966 (N_12966,N_11136,N_10819);
nor U12967 (N_12967,N_10148,N_10620);
nor U12968 (N_12968,N_11526,N_11714);
xor U12969 (N_12969,N_11186,N_11558);
nand U12970 (N_12970,N_10671,N_10040);
and U12971 (N_12971,N_10903,N_10367);
xnor U12972 (N_12972,N_10427,N_10271);
nand U12973 (N_12973,N_10906,N_10812);
and U12974 (N_12974,N_11427,N_10617);
nor U12975 (N_12975,N_11755,N_11603);
and U12976 (N_12976,N_11459,N_11129);
and U12977 (N_12977,N_10479,N_11160);
nand U12978 (N_12978,N_11629,N_11673);
and U12979 (N_12979,N_10944,N_11110);
nor U12980 (N_12980,N_11001,N_11116);
and U12981 (N_12981,N_11157,N_10570);
or U12982 (N_12982,N_11641,N_10993);
and U12983 (N_12983,N_11521,N_11159);
nand U12984 (N_12984,N_11807,N_11674);
nor U12985 (N_12985,N_10596,N_11193);
or U12986 (N_12986,N_10060,N_10178);
nand U12987 (N_12987,N_11679,N_11995);
xnor U12988 (N_12988,N_11856,N_11706);
nand U12989 (N_12989,N_10900,N_11150);
or U12990 (N_12990,N_11453,N_10118);
nand U12991 (N_12991,N_10216,N_10433);
xor U12992 (N_12992,N_11878,N_10136);
or U12993 (N_12993,N_10675,N_11138);
nand U12994 (N_12994,N_11688,N_10625);
and U12995 (N_12995,N_10364,N_11991);
nand U12996 (N_12996,N_11505,N_10727);
and U12997 (N_12997,N_11126,N_10869);
nor U12998 (N_12998,N_10377,N_10749);
nor U12999 (N_12999,N_10737,N_10739);
nor U13000 (N_13000,N_10370,N_11161);
and U13001 (N_13001,N_11950,N_11788);
and U13002 (N_13002,N_11410,N_10113);
nand U13003 (N_13003,N_11886,N_11389);
nor U13004 (N_13004,N_10699,N_11717);
or U13005 (N_13005,N_11103,N_11511);
and U13006 (N_13006,N_11412,N_11737);
nor U13007 (N_13007,N_11848,N_11923);
nand U13008 (N_13008,N_10658,N_11192);
xnor U13009 (N_13009,N_10660,N_11098);
xor U13010 (N_13010,N_10600,N_11640);
nor U13011 (N_13011,N_11452,N_11000);
or U13012 (N_13012,N_10371,N_10249);
and U13013 (N_13013,N_10223,N_11684);
or U13014 (N_13014,N_11767,N_10042);
and U13015 (N_13015,N_11103,N_10264);
nor U13016 (N_13016,N_10126,N_11655);
and U13017 (N_13017,N_11114,N_11625);
nor U13018 (N_13018,N_10380,N_11333);
or U13019 (N_13019,N_10291,N_10484);
xnor U13020 (N_13020,N_11179,N_11536);
and U13021 (N_13021,N_11069,N_11534);
nand U13022 (N_13022,N_10381,N_11185);
nor U13023 (N_13023,N_11685,N_10818);
nor U13024 (N_13024,N_11769,N_11248);
nor U13025 (N_13025,N_11828,N_10881);
nor U13026 (N_13026,N_11168,N_10909);
and U13027 (N_13027,N_11867,N_11619);
nor U13028 (N_13028,N_10653,N_10373);
nor U13029 (N_13029,N_11650,N_10190);
and U13030 (N_13030,N_10642,N_10567);
xor U13031 (N_13031,N_11197,N_10724);
or U13032 (N_13032,N_11173,N_11400);
nor U13033 (N_13033,N_10656,N_11371);
xor U13034 (N_13034,N_10203,N_10503);
or U13035 (N_13035,N_10982,N_10627);
xor U13036 (N_13036,N_10524,N_11976);
nand U13037 (N_13037,N_11493,N_11139);
nand U13038 (N_13038,N_10874,N_10737);
xor U13039 (N_13039,N_11919,N_11841);
xnor U13040 (N_13040,N_10256,N_11677);
nand U13041 (N_13041,N_10238,N_10133);
nor U13042 (N_13042,N_11673,N_11499);
or U13043 (N_13043,N_11379,N_10670);
xor U13044 (N_13044,N_11858,N_10933);
nor U13045 (N_13045,N_11215,N_11263);
nand U13046 (N_13046,N_11130,N_11017);
xnor U13047 (N_13047,N_11246,N_11512);
nor U13048 (N_13048,N_11458,N_10340);
and U13049 (N_13049,N_11629,N_10885);
and U13050 (N_13050,N_11329,N_10455);
xor U13051 (N_13051,N_10468,N_11290);
nand U13052 (N_13052,N_11649,N_10173);
or U13053 (N_13053,N_11128,N_10225);
nor U13054 (N_13054,N_10175,N_10254);
and U13055 (N_13055,N_10183,N_10419);
or U13056 (N_13056,N_11992,N_11920);
and U13057 (N_13057,N_11276,N_10673);
xnor U13058 (N_13058,N_11954,N_10582);
or U13059 (N_13059,N_10826,N_10269);
xnor U13060 (N_13060,N_10032,N_10993);
xnor U13061 (N_13061,N_11409,N_11168);
nor U13062 (N_13062,N_11933,N_10467);
nor U13063 (N_13063,N_11564,N_11926);
and U13064 (N_13064,N_10813,N_11770);
xor U13065 (N_13065,N_11384,N_10960);
xnor U13066 (N_13066,N_10755,N_10002);
and U13067 (N_13067,N_10687,N_10705);
xnor U13068 (N_13068,N_10014,N_11980);
and U13069 (N_13069,N_10687,N_11720);
or U13070 (N_13070,N_10831,N_11283);
or U13071 (N_13071,N_10049,N_11660);
xor U13072 (N_13072,N_11611,N_11693);
and U13073 (N_13073,N_11268,N_10204);
or U13074 (N_13074,N_10467,N_10288);
nand U13075 (N_13075,N_10260,N_10691);
and U13076 (N_13076,N_11564,N_11736);
xnor U13077 (N_13077,N_10573,N_11894);
or U13078 (N_13078,N_10624,N_10768);
or U13079 (N_13079,N_11365,N_11052);
and U13080 (N_13080,N_10532,N_10473);
xnor U13081 (N_13081,N_11680,N_11176);
or U13082 (N_13082,N_10102,N_10400);
xnor U13083 (N_13083,N_10221,N_11750);
xnor U13084 (N_13084,N_11730,N_11038);
nor U13085 (N_13085,N_11568,N_10237);
nor U13086 (N_13086,N_10709,N_10742);
and U13087 (N_13087,N_10582,N_10225);
nand U13088 (N_13088,N_11470,N_11873);
nor U13089 (N_13089,N_10005,N_10296);
and U13090 (N_13090,N_11676,N_11217);
or U13091 (N_13091,N_10691,N_10940);
nand U13092 (N_13092,N_10362,N_10093);
xnor U13093 (N_13093,N_11151,N_11158);
xor U13094 (N_13094,N_10038,N_10913);
nand U13095 (N_13095,N_11627,N_11364);
and U13096 (N_13096,N_11846,N_10368);
and U13097 (N_13097,N_11358,N_11107);
xnor U13098 (N_13098,N_11410,N_10381);
and U13099 (N_13099,N_11175,N_11719);
xnor U13100 (N_13100,N_11491,N_10091);
or U13101 (N_13101,N_10538,N_10647);
or U13102 (N_13102,N_10566,N_11078);
nand U13103 (N_13103,N_10771,N_10424);
nor U13104 (N_13104,N_11570,N_11470);
nand U13105 (N_13105,N_10382,N_11906);
and U13106 (N_13106,N_10817,N_11447);
nand U13107 (N_13107,N_10326,N_11928);
nand U13108 (N_13108,N_10561,N_10633);
xnor U13109 (N_13109,N_10418,N_10582);
or U13110 (N_13110,N_11182,N_11644);
or U13111 (N_13111,N_10119,N_10137);
nand U13112 (N_13112,N_10209,N_10103);
nand U13113 (N_13113,N_11768,N_11913);
and U13114 (N_13114,N_10378,N_10233);
xor U13115 (N_13115,N_11470,N_10437);
nor U13116 (N_13116,N_11232,N_10442);
nor U13117 (N_13117,N_10377,N_10832);
and U13118 (N_13118,N_11995,N_10441);
nand U13119 (N_13119,N_11333,N_11851);
nand U13120 (N_13120,N_10921,N_10255);
nor U13121 (N_13121,N_11973,N_10004);
nor U13122 (N_13122,N_11946,N_11686);
xor U13123 (N_13123,N_10114,N_10695);
and U13124 (N_13124,N_10020,N_11948);
or U13125 (N_13125,N_11828,N_10171);
xor U13126 (N_13126,N_11688,N_10245);
and U13127 (N_13127,N_10577,N_10447);
nand U13128 (N_13128,N_11691,N_10270);
xor U13129 (N_13129,N_11593,N_11486);
xnor U13130 (N_13130,N_10249,N_11282);
nand U13131 (N_13131,N_11207,N_11103);
nand U13132 (N_13132,N_11903,N_11732);
nor U13133 (N_13133,N_10478,N_10378);
nand U13134 (N_13134,N_10116,N_10934);
nand U13135 (N_13135,N_10710,N_11328);
and U13136 (N_13136,N_11132,N_10837);
xnor U13137 (N_13137,N_10807,N_10234);
and U13138 (N_13138,N_10575,N_11087);
or U13139 (N_13139,N_10051,N_10890);
nor U13140 (N_13140,N_11156,N_11793);
and U13141 (N_13141,N_11552,N_11907);
or U13142 (N_13142,N_11101,N_10906);
or U13143 (N_13143,N_11054,N_10900);
xnor U13144 (N_13144,N_10767,N_10280);
or U13145 (N_13145,N_10983,N_11048);
and U13146 (N_13146,N_10041,N_11687);
nor U13147 (N_13147,N_10927,N_10305);
nand U13148 (N_13148,N_10339,N_10175);
nor U13149 (N_13149,N_10818,N_11506);
nor U13150 (N_13150,N_11030,N_10044);
nand U13151 (N_13151,N_10514,N_11481);
and U13152 (N_13152,N_11822,N_11774);
and U13153 (N_13153,N_11963,N_11018);
xnor U13154 (N_13154,N_10302,N_11114);
nor U13155 (N_13155,N_10797,N_11764);
xor U13156 (N_13156,N_11884,N_11001);
and U13157 (N_13157,N_11947,N_10078);
nand U13158 (N_13158,N_11273,N_11493);
xnor U13159 (N_13159,N_10036,N_10047);
or U13160 (N_13160,N_10780,N_11386);
nor U13161 (N_13161,N_11723,N_10066);
nor U13162 (N_13162,N_10438,N_11991);
nor U13163 (N_13163,N_11248,N_11464);
xnor U13164 (N_13164,N_11815,N_11772);
or U13165 (N_13165,N_11093,N_11307);
nor U13166 (N_13166,N_11062,N_11321);
or U13167 (N_13167,N_10547,N_10310);
nor U13168 (N_13168,N_10700,N_11608);
xor U13169 (N_13169,N_10994,N_10753);
nor U13170 (N_13170,N_11726,N_11120);
nor U13171 (N_13171,N_10496,N_11358);
and U13172 (N_13172,N_11304,N_11193);
or U13173 (N_13173,N_10361,N_11890);
and U13174 (N_13174,N_11015,N_11661);
or U13175 (N_13175,N_10389,N_11892);
or U13176 (N_13176,N_11020,N_10233);
xnor U13177 (N_13177,N_11370,N_11988);
xor U13178 (N_13178,N_11949,N_11711);
xnor U13179 (N_13179,N_10562,N_10144);
and U13180 (N_13180,N_11502,N_10954);
nand U13181 (N_13181,N_10749,N_10750);
or U13182 (N_13182,N_11960,N_11672);
xnor U13183 (N_13183,N_11713,N_11205);
and U13184 (N_13184,N_11827,N_10053);
and U13185 (N_13185,N_10434,N_10673);
nand U13186 (N_13186,N_11128,N_10951);
or U13187 (N_13187,N_10211,N_11092);
nor U13188 (N_13188,N_11607,N_10782);
nor U13189 (N_13189,N_10812,N_11221);
xor U13190 (N_13190,N_11223,N_11335);
nand U13191 (N_13191,N_10764,N_11290);
or U13192 (N_13192,N_10759,N_10222);
xnor U13193 (N_13193,N_10437,N_10617);
or U13194 (N_13194,N_11251,N_10630);
nand U13195 (N_13195,N_10399,N_10099);
nand U13196 (N_13196,N_10680,N_11680);
xor U13197 (N_13197,N_11051,N_10865);
nand U13198 (N_13198,N_10981,N_10129);
nor U13199 (N_13199,N_11167,N_11385);
and U13200 (N_13200,N_10981,N_10160);
or U13201 (N_13201,N_10840,N_11754);
xnor U13202 (N_13202,N_10830,N_10852);
and U13203 (N_13203,N_10120,N_10577);
nor U13204 (N_13204,N_10792,N_10564);
and U13205 (N_13205,N_10567,N_11399);
or U13206 (N_13206,N_10448,N_11825);
nor U13207 (N_13207,N_10962,N_11639);
xor U13208 (N_13208,N_10292,N_10709);
nor U13209 (N_13209,N_11944,N_10454);
or U13210 (N_13210,N_10524,N_11907);
and U13211 (N_13211,N_10964,N_10521);
nand U13212 (N_13212,N_10123,N_10019);
xnor U13213 (N_13213,N_11624,N_10155);
or U13214 (N_13214,N_10509,N_10986);
and U13215 (N_13215,N_11329,N_10629);
xor U13216 (N_13216,N_11505,N_11608);
nor U13217 (N_13217,N_11943,N_10098);
and U13218 (N_13218,N_11496,N_11889);
nor U13219 (N_13219,N_11711,N_11029);
or U13220 (N_13220,N_10550,N_11917);
and U13221 (N_13221,N_10587,N_11926);
and U13222 (N_13222,N_11373,N_10323);
and U13223 (N_13223,N_11361,N_10688);
nand U13224 (N_13224,N_11195,N_11657);
nand U13225 (N_13225,N_10942,N_10241);
nor U13226 (N_13226,N_11873,N_10613);
nor U13227 (N_13227,N_10328,N_11351);
xnor U13228 (N_13228,N_10909,N_11336);
xnor U13229 (N_13229,N_11554,N_11426);
or U13230 (N_13230,N_11842,N_11674);
nor U13231 (N_13231,N_10322,N_11493);
or U13232 (N_13232,N_10022,N_11767);
nand U13233 (N_13233,N_10552,N_10507);
nand U13234 (N_13234,N_11343,N_10934);
xnor U13235 (N_13235,N_10177,N_11145);
xor U13236 (N_13236,N_11713,N_10733);
nand U13237 (N_13237,N_10978,N_11943);
xnor U13238 (N_13238,N_10658,N_11332);
and U13239 (N_13239,N_10021,N_10061);
or U13240 (N_13240,N_10637,N_10763);
xnor U13241 (N_13241,N_10074,N_11074);
xnor U13242 (N_13242,N_11191,N_10671);
and U13243 (N_13243,N_10437,N_11179);
nor U13244 (N_13244,N_10488,N_10335);
nor U13245 (N_13245,N_10312,N_10032);
nand U13246 (N_13246,N_10360,N_10316);
nand U13247 (N_13247,N_11104,N_11440);
and U13248 (N_13248,N_11150,N_11134);
nand U13249 (N_13249,N_11772,N_11226);
nor U13250 (N_13250,N_11036,N_11397);
xor U13251 (N_13251,N_11430,N_10236);
xor U13252 (N_13252,N_11510,N_10507);
nand U13253 (N_13253,N_11795,N_11202);
nor U13254 (N_13254,N_10642,N_10664);
or U13255 (N_13255,N_11185,N_11240);
xnor U13256 (N_13256,N_11303,N_10363);
nand U13257 (N_13257,N_10291,N_11622);
or U13258 (N_13258,N_11437,N_10715);
and U13259 (N_13259,N_11646,N_10473);
xnor U13260 (N_13260,N_11984,N_10154);
xor U13261 (N_13261,N_11630,N_10487);
and U13262 (N_13262,N_11946,N_11731);
nor U13263 (N_13263,N_11539,N_10717);
or U13264 (N_13264,N_11415,N_10030);
xnor U13265 (N_13265,N_10504,N_11049);
and U13266 (N_13266,N_10131,N_11399);
nand U13267 (N_13267,N_11586,N_11754);
or U13268 (N_13268,N_10241,N_10455);
or U13269 (N_13269,N_11687,N_10619);
nand U13270 (N_13270,N_11694,N_11160);
xnor U13271 (N_13271,N_11209,N_11857);
xor U13272 (N_13272,N_10040,N_11791);
nor U13273 (N_13273,N_10122,N_11688);
nor U13274 (N_13274,N_11940,N_10805);
nand U13275 (N_13275,N_10667,N_11659);
xor U13276 (N_13276,N_11435,N_11935);
or U13277 (N_13277,N_11847,N_11729);
xnor U13278 (N_13278,N_11424,N_11335);
or U13279 (N_13279,N_10956,N_11422);
nor U13280 (N_13280,N_11030,N_10699);
xor U13281 (N_13281,N_10855,N_10475);
nand U13282 (N_13282,N_10061,N_10494);
nand U13283 (N_13283,N_10818,N_11643);
and U13284 (N_13284,N_11948,N_10634);
xor U13285 (N_13285,N_11114,N_11311);
and U13286 (N_13286,N_11427,N_11146);
nor U13287 (N_13287,N_10584,N_11376);
nand U13288 (N_13288,N_11278,N_10676);
nor U13289 (N_13289,N_11982,N_10342);
or U13290 (N_13290,N_10266,N_11399);
nand U13291 (N_13291,N_11658,N_10741);
and U13292 (N_13292,N_10071,N_10403);
nand U13293 (N_13293,N_10384,N_11595);
xnor U13294 (N_13294,N_10831,N_10127);
nor U13295 (N_13295,N_11702,N_11965);
xnor U13296 (N_13296,N_11380,N_11860);
and U13297 (N_13297,N_10653,N_10751);
or U13298 (N_13298,N_11517,N_10887);
and U13299 (N_13299,N_11068,N_10644);
or U13300 (N_13300,N_11609,N_11750);
and U13301 (N_13301,N_10273,N_11982);
xor U13302 (N_13302,N_10647,N_10743);
xor U13303 (N_13303,N_11539,N_11723);
and U13304 (N_13304,N_11230,N_11436);
or U13305 (N_13305,N_11297,N_10187);
nor U13306 (N_13306,N_11947,N_11945);
nand U13307 (N_13307,N_11867,N_10403);
xnor U13308 (N_13308,N_11154,N_10026);
or U13309 (N_13309,N_11249,N_10567);
or U13310 (N_13310,N_10360,N_11416);
and U13311 (N_13311,N_10379,N_10636);
nand U13312 (N_13312,N_10588,N_10847);
nor U13313 (N_13313,N_11577,N_11442);
xnor U13314 (N_13314,N_10453,N_11685);
xor U13315 (N_13315,N_11644,N_10839);
nor U13316 (N_13316,N_11173,N_10284);
and U13317 (N_13317,N_10147,N_10440);
xnor U13318 (N_13318,N_11500,N_11068);
nand U13319 (N_13319,N_11325,N_11396);
nor U13320 (N_13320,N_11245,N_11438);
and U13321 (N_13321,N_10234,N_11901);
and U13322 (N_13322,N_10818,N_11803);
nand U13323 (N_13323,N_11285,N_11814);
and U13324 (N_13324,N_11895,N_11946);
or U13325 (N_13325,N_10061,N_11517);
or U13326 (N_13326,N_10880,N_10325);
or U13327 (N_13327,N_11893,N_11517);
xnor U13328 (N_13328,N_10192,N_10749);
nor U13329 (N_13329,N_11694,N_11676);
xnor U13330 (N_13330,N_11138,N_11353);
nand U13331 (N_13331,N_11940,N_11898);
nor U13332 (N_13332,N_11118,N_10871);
nor U13333 (N_13333,N_11798,N_10759);
xnor U13334 (N_13334,N_10696,N_10745);
or U13335 (N_13335,N_11166,N_11433);
nand U13336 (N_13336,N_11378,N_11579);
and U13337 (N_13337,N_10150,N_10957);
or U13338 (N_13338,N_11999,N_11018);
xnor U13339 (N_13339,N_11379,N_11148);
xor U13340 (N_13340,N_10344,N_10143);
or U13341 (N_13341,N_10317,N_11402);
xnor U13342 (N_13342,N_10791,N_10734);
nand U13343 (N_13343,N_10171,N_10800);
xnor U13344 (N_13344,N_11222,N_11409);
or U13345 (N_13345,N_11805,N_10577);
xor U13346 (N_13346,N_11308,N_11859);
nor U13347 (N_13347,N_11046,N_11918);
xnor U13348 (N_13348,N_10389,N_11269);
or U13349 (N_13349,N_10452,N_10890);
or U13350 (N_13350,N_10358,N_10233);
and U13351 (N_13351,N_10238,N_10264);
nor U13352 (N_13352,N_11214,N_10934);
nand U13353 (N_13353,N_11099,N_11611);
and U13354 (N_13354,N_11751,N_10331);
nor U13355 (N_13355,N_11492,N_11761);
nor U13356 (N_13356,N_10395,N_10890);
nor U13357 (N_13357,N_11597,N_11063);
or U13358 (N_13358,N_11008,N_11421);
nor U13359 (N_13359,N_10664,N_11005);
nor U13360 (N_13360,N_11892,N_11380);
or U13361 (N_13361,N_10668,N_11830);
nor U13362 (N_13362,N_10142,N_11809);
nor U13363 (N_13363,N_11293,N_10831);
nor U13364 (N_13364,N_10065,N_10018);
xor U13365 (N_13365,N_10161,N_11422);
or U13366 (N_13366,N_11124,N_11698);
xor U13367 (N_13367,N_10681,N_10858);
and U13368 (N_13368,N_10181,N_11297);
and U13369 (N_13369,N_10104,N_10629);
or U13370 (N_13370,N_11851,N_10410);
and U13371 (N_13371,N_11379,N_11244);
and U13372 (N_13372,N_11143,N_10903);
or U13373 (N_13373,N_11485,N_11578);
nor U13374 (N_13374,N_10174,N_10829);
and U13375 (N_13375,N_11416,N_11305);
or U13376 (N_13376,N_11919,N_11389);
nor U13377 (N_13377,N_10167,N_10063);
nand U13378 (N_13378,N_10731,N_11261);
nand U13379 (N_13379,N_10797,N_10295);
nor U13380 (N_13380,N_10038,N_10733);
xnor U13381 (N_13381,N_10428,N_11664);
and U13382 (N_13382,N_11705,N_11854);
nand U13383 (N_13383,N_10975,N_11408);
nor U13384 (N_13384,N_11687,N_10998);
and U13385 (N_13385,N_10372,N_10428);
nor U13386 (N_13386,N_11048,N_11056);
and U13387 (N_13387,N_11186,N_11720);
and U13388 (N_13388,N_10011,N_11005);
or U13389 (N_13389,N_11750,N_10600);
xnor U13390 (N_13390,N_11260,N_11829);
nand U13391 (N_13391,N_10300,N_10065);
xnor U13392 (N_13392,N_10497,N_11399);
xor U13393 (N_13393,N_10749,N_10586);
and U13394 (N_13394,N_11745,N_10189);
and U13395 (N_13395,N_10193,N_11719);
nor U13396 (N_13396,N_10994,N_10750);
nand U13397 (N_13397,N_10736,N_10365);
and U13398 (N_13398,N_10434,N_10649);
and U13399 (N_13399,N_11019,N_11766);
and U13400 (N_13400,N_10704,N_11773);
nand U13401 (N_13401,N_11114,N_11249);
and U13402 (N_13402,N_10968,N_11657);
nor U13403 (N_13403,N_10382,N_11620);
or U13404 (N_13404,N_10008,N_10370);
and U13405 (N_13405,N_10135,N_11372);
xor U13406 (N_13406,N_11699,N_10171);
and U13407 (N_13407,N_11588,N_10643);
and U13408 (N_13408,N_10637,N_10733);
nand U13409 (N_13409,N_10340,N_10974);
xnor U13410 (N_13410,N_11449,N_11415);
and U13411 (N_13411,N_10339,N_11072);
nand U13412 (N_13412,N_11857,N_10289);
nand U13413 (N_13413,N_10859,N_10428);
nand U13414 (N_13414,N_11612,N_11691);
xor U13415 (N_13415,N_10924,N_10777);
or U13416 (N_13416,N_10415,N_11624);
xnor U13417 (N_13417,N_10499,N_10217);
or U13418 (N_13418,N_11596,N_11507);
or U13419 (N_13419,N_10595,N_11942);
nor U13420 (N_13420,N_11990,N_11196);
and U13421 (N_13421,N_11922,N_11397);
nor U13422 (N_13422,N_10663,N_11893);
or U13423 (N_13423,N_10769,N_11204);
and U13424 (N_13424,N_11135,N_10956);
nor U13425 (N_13425,N_10782,N_10212);
and U13426 (N_13426,N_11969,N_10251);
xor U13427 (N_13427,N_10703,N_11023);
or U13428 (N_13428,N_10664,N_10735);
nor U13429 (N_13429,N_10429,N_10751);
or U13430 (N_13430,N_10862,N_11124);
or U13431 (N_13431,N_11379,N_10167);
nor U13432 (N_13432,N_11384,N_10422);
and U13433 (N_13433,N_11699,N_10142);
nor U13434 (N_13434,N_11003,N_11609);
and U13435 (N_13435,N_11927,N_11376);
xor U13436 (N_13436,N_11532,N_11690);
or U13437 (N_13437,N_10903,N_10812);
xor U13438 (N_13438,N_10121,N_10213);
or U13439 (N_13439,N_10536,N_11526);
nand U13440 (N_13440,N_11866,N_10025);
nor U13441 (N_13441,N_11516,N_10246);
and U13442 (N_13442,N_11683,N_10601);
nand U13443 (N_13443,N_11225,N_10109);
nand U13444 (N_13444,N_11237,N_10141);
nand U13445 (N_13445,N_10192,N_10829);
xnor U13446 (N_13446,N_10912,N_11743);
or U13447 (N_13447,N_11793,N_11868);
xor U13448 (N_13448,N_10000,N_11166);
and U13449 (N_13449,N_10551,N_11082);
nor U13450 (N_13450,N_11822,N_10214);
nor U13451 (N_13451,N_10779,N_11232);
or U13452 (N_13452,N_10911,N_10509);
nor U13453 (N_13453,N_10804,N_11889);
nand U13454 (N_13454,N_10971,N_11240);
and U13455 (N_13455,N_11697,N_10906);
nor U13456 (N_13456,N_10194,N_10261);
and U13457 (N_13457,N_11555,N_10044);
nand U13458 (N_13458,N_10445,N_11333);
xnor U13459 (N_13459,N_10526,N_10274);
xor U13460 (N_13460,N_10909,N_11236);
or U13461 (N_13461,N_10999,N_11535);
nand U13462 (N_13462,N_10244,N_10672);
nor U13463 (N_13463,N_11042,N_11177);
nor U13464 (N_13464,N_11543,N_10107);
and U13465 (N_13465,N_10518,N_10183);
xnor U13466 (N_13466,N_11723,N_11242);
nor U13467 (N_13467,N_10959,N_10708);
or U13468 (N_13468,N_11145,N_11030);
nand U13469 (N_13469,N_10639,N_10104);
and U13470 (N_13470,N_10734,N_10277);
nand U13471 (N_13471,N_11777,N_11754);
or U13472 (N_13472,N_10450,N_11587);
and U13473 (N_13473,N_11047,N_11563);
or U13474 (N_13474,N_10416,N_11543);
nand U13475 (N_13475,N_11826,N_11539);
and U13476 (N_13476,N_10804,N_11521);
nor U13477 (N_13477,N_10645,N_10844);
nand U13478 (N_13478,N_11409,N_11463);
or U13479 (N_13479,N_11395,N_10563);
and U13480 (N_13480,N_11679,N_11788);
or U13481 (N_13481,N_10044,N_11807);
nor U13482 (N_13482,N_11600,N_10780);
xor U13483 (N_13483,N_11288,N_11287);
and U13484 (N_13484,N_10720,N_10237);
nor U13485 (N_13485,N_10687,N_11770);
or U13486 (N_13486,N_10912,N_11932);
nor U13487 (N_13487,N_10360,N_10627);
nand U13488 (N_13488,N_10580,N_10222);
and U13489 (N_13489,N_10827,N_11143);
and U13490 (N_13490,N_11959,N_10231);
xnor U13491 (N_13491,N_11429,N_10409);
xnor U13492 (N_13492,N_11145,N_11350);
nor U13493 (N_13493,N_11976,N_10916);
or U13494 (N_13494,N_11562,N_10676);
or U13495 (N_13495,N_11010,N_11120);
xor U13496 (N_13496,N_10016,N_11905);
xnor U13497 (N_13497,N_10851,N_11336);
nor U13498 (N_13498,N_11609,N_10241);
or U13499 (N_13499,N_11485,N_11370);
nor U13500 (N_13500,N_11026,N_11648);
nor U13501 (N_13501,N_10660,N_10946);
or U13502 (N_13502,N_10677,N_10312);
or U13503 (N_13503,N_11968,N_11048);
and U13504 (N_13504,N_10596,N_11436);
xor U13505 (N_13505,N_10420,N_11312);
nor U13506 (N_13506,N_10265,N_11870);
nand U13507 (N_13507,N_10394,N_10684);
or U13508 (N_13508,N_11278,N_10373);
nand U13509 (N_13509,N_11532,N_10837);
nand U13510 (N_13510,N_10792,N_10278);
nand U13511 (N_13511,N_10390,N_10982);
xnor U13512 (N_13512,N_10261,N_10883);
nor U13513 (N_13513,N_10789,N_11155);
xor U13514 (N_13514,N_11945,N_11774);
and U13515 (N_13515,N_11152,N_10105);
nor U13516 (N_13516,N_10391,N_11469);
xor U13517 (N_13517,N_10652,N_11026);
nor U13518 (N_13518,N_11723,N_11031);
and U13519 (N_13519,N_10749,N_11298);
nand U13520 (N_13520,N_10600,N_10966);
nor U13521 (N_13521,N_10788,N_10534);
and U13522 (N_13522,N_11372,N_10696);
nor U13523 (N_13523,N_11433,N_10887);
nor U13524 (N_13524,N_10478,N_10967);
xor U13525 (N_13525,N_10565,N_11149);
and U13526 (N_13526,N_11927,N_10424);
and U13527 (N_13527,N_10282,N_10442);
nand U13528 (N_13528,N_11224,N_11711);
nand U13529 (N_13529,N_10331,N_10721);
and U13530 (N_13530,N_11087,N_10239);
nor U13531 (N_13531,N_11214,N_10726);
and U13532 (N_13532,N_11249,N_10357);
nand U13533 (N_13533,N_10125,N_11574);
and U13534 (N_13534,N_10729,N_11553);
or U13535 (N_13535,N_10179,N_11357);
and U13536 (N_13536,N_10567,N_11542);
nand U13537 (N_13537,N_11688,N_10066);
and U13538 (N_13538,N_11003,N_10739);
xor U13539 (N_13539,N_10873,N_10255);
nor U13540 (N_13540,N_11825,N_11505);
nand U13541 (N_13541,N_10777,N_11767);
nand U13542 (N_13542,N_10377,N_11979);
or U13543 (N_13543,N_11805,N_10717);
and U13544 (N_13544,N_11165,N_10056);
nor U13545 (N_13545,N_11148,N_11596);
and U13546 (N_13546,N_10046,N_10303);
nor U13547 (N_13547,N_11615,N_10071);
and U13548 (N_13548,N_11206,N_10348);
and U13549 (N_13549,N_11543,N_11579);
nand U13550 (N_13550,N_10612,N_11289);
or U13551 (N_13551,N_10457,N_10320);
xor U13552 (N_13552,N_10719,N_11463);
nor U13553 (N_13553,N_10195,N_10319);
nor U13554 (N_13554,N_10023,N_10388);
or U13555 (N_13555,N_11101,N_11690);
and U13556 (N_13556,N_10297,N_11152);
and U13557 (N_13557,N_10689,N_10047);
and U13558 (N_13558,N_10363,N_10202);
and U13559 (N_13559,N_10270,N_10075);
nor U13560 (N_13560,N_10020,N_10811);
xor U13561 (N_13561,N_11268,N_10019);
or U13562 (N_13562,N_10721,N_11689);
nor U13563 (N_13563,N_11112,N_10804);
nor U13564 (N_13564,N_10774,N_11025);
xor U13565 (N_13565,N_11644,N_10843);
xor U13566 (N_13566,N_11200,N_10424);
xnor U13567 (N_13567,N_11596,N_10124);
and U13568 (N_13568,N_11285,N_10830);
or U13569 (N_13569,N_10407,N_10750);
or U13570 (N_13570,N_10171,N_10267);
nor U13571 (N_13571,N_11099,N_11124);
and U13572 (N_13572,N_11730,N_11716);
xor U13573 (N_13573,N_10931,N_11994);
nand U13574 (N_13574,N_10062,N_11071);
xor U13575 (N_13575,N_11069,N_11572);
nand U13576 (N_13576,N_11395,N_10070);
or U13577 (N_13577,N_10399,N_10735);
or U13578 (N_13578,N_11788,N_10835);
nor U13579 (N_13579,N_11729,N_10518);
nand U13580 (N_13580,N_10239,N_10400);
and U13581 (N_13581,N_10979,N_10220);
nand U13582 (N_13582,N_10255,N_10983);
and U13583 (N_13583,N_11081,N_11885);
nor U13584 (N_13584,N_11475,N_11073);
or U13585 (N_13585,N_10044,N_10844);
or U13586 (N_13586,N_10294,N_11418);
and U13587 (N_13587,N_11350,N_10827);
xor U13588 (N_13588,N_10260,N_10098);
nor U13589 (N_13589,N_11879,N_11338);
nor U13590 (N_13590,N_10002,N_11721);
and U13591 (N_13591,N_11188,N_10664);
nor U13592 (N_13592,N_10516,N_11416);
nand U13593 (N_13593,N_10038,N_10537);
nor U13594 (N_13594,N_11278,N_10912);
and U13595 (N_13595,N_10767,N_11414);
or U13596 (N_13596,N_11582,N_10895);
and U13597 (N_13597,N_11169,N_11743);
and U13598 (N_13598,N_11067,N_10589);
xnor U13599 (N_13599,N_11739,N_11969);
or U13600 (N_13600,N_11840,N_10329);
xnor U13601 (N_13601,N_11489,N_11023);
xnor U13602 (N_13602,N_11268,N_11502);
and U13603 (N_13603,N_11023,N_11794);
nor U13604 (N_13604,N_10270,N_10432);
or U13605 (N_13605,N_10848,N_11131);
and U13606 (N_13606,N_10708,N_10714);
xor U13607 (N_13607,N_11602,N_11918);
nand U13608 (N_13608,N_11188,N_10870);
and U13609 (N_13609,N_10827,N_10440);
and U13610 (N_13610,N_10969,N_10670);
or U13611 (N_13611,N_11853,N_10998);
nor U13612 (N_13612,N_10762,N_10673);
or U13613 (N_13613,N_10286,N_10674);
and U13614 (N_13614,N_11792,N_10375);
xnor U13615 (N_13615,N_11286,N_10446);
and U13616 (N_13616,N_10355,N_10367);
and U13617 (N_13617,N_10016,N_11880);
and U13618 (N_13618,N_11919,N_10002);
or U13619 (N_13619,N_10251,N_11476);
or U13620 (N_13620,N_11463,N_10456);
nand U13621 (N_13621,N_11278,N_10502);
and U13622 (N_13622,N_11813,N_10447);
xor U13623 (N_13623,N_10449,N_10033);
xnor U13624 (N_13624,N_10509,N_11521);
and U13625 (N_13625,N_10263,N_10331);
nand U13626 (N_13626,N_11357,N_11565);
xor U13627 (N_13627,N_10124,N_11143);
and U13628 (N_13628,N_10187,N_10249);
or U13629 (N_13629,N_10233,N_11616);
nor U13630 (N_13630,N_10401,N_10851);
nand U13631 (N_13631,N_11492,N_10808);
xnor U13632 (N_13632,N_10363,N_11028);
nor U13633 (N_13633,N_11933,N_10199);
nor U13634 (N_13634,N_11523,N_11132);
and U13635 (N_13635,N_11389,N_10158);
nand U13636 (N_13636,N_10366,N_10886);
nor U13637 (N_13637,N_10501,N_11234);
and U13638 (N_13638,N_10927,N_11617);
nand U13639 (N_13639,N_10545,N_11664);
nand U13640 (N_13640,N_10281,N_11652);
or U13641 (N_13641,N_10260,N_11354);
nor U13642 (N_13642,N_10569,N_10754);
nand U13643 (N_13643,N_10046,N_11827);
nor U13644 (N_13644,N_11503,N_11835);
nor U13645 (N_13645,N_11029,N_10862);
nor U13646 (N_13646,N_10470,N_11029);
or U13647 (N_13647,N_10244,N_11918);
or U13648 (N_13648,N_10583,N_11727);
or U13649 (N_13649,N_10011,N_11278);
and U13650 (N_13650,N_11286,N_10453);
nor U13651 (N_13651,N_11689,N_10971);
and U13652 (N_13652,N_11719,N_10126);
and U13653 (N_13653,N_11490,N_10130);
and U13654 (N_13654,N_11322,N_11723);
or U13655 (N_13655,N_10757,N_11464);
nor U13656 (N_13656,N_10312,N_11409);
and U13657 (N_13657,N_11903,N_11831);
or U13658 (N_13658,N_10151,N_11591);
or U13659 (N_13659,N_10931,N_11763);
or U13660 (N_13660,N_11018,N_11400);
nand U13661 (N_13661,N_11210,N_10979);
and U13662 (N_13662,N_10720,N_10989);
or U13663 (N_13663,N_11444,N_11590);
or U13664 (N_13664,N_11519,N_11541);
or U13665 (N_13665,N_10028,N_11868);
nand U13666 (N_13666,N_11119,N_11430);
and U13667 (N_13667,N_10805,N_10263);
or U13668 (N_13668,N_11688,N_11518);
or U13669 (N_13669,N_10881,N_10682);
or U13670 (N_13670,N_10670,N_11921);
nand U13671 (N_13671,N_11008,N_10798);
and U13672 (N_13672,N_10125,N_11906);
or U13673 (N_13673,N_11126,N_11893);
and U13674 (N_13674,N_11444,N_11755);
and U13675 (N_13675,N_10585,N_11002);
xnor U13676 (N_13676,N_11488,N_10511);
and U13677 (N_13677,N_11628,N_10353);
and U13678 (N_13678,N_11861,N_11987);
nand U13679 (N_13679,N_10626,N_10657);
nand U13680 (N_13680,N_10050,N_11380);
xnor U13681 (N_13681,N_10406,N_10217);
nor U13682 (N_13682,N_11683,N_11329);
nand U13683 (N_13683,N_10113,N_11677);
nand U13684 (N_13684,N_10088,N_10107);
or U13685 (N_13685,N_10939,N_10189);
xnor U13686 (N_13686,N_11774,N_11471);
or U13687 (N_13687,N_10446,N_11004);
or U13688 (N_13688,N_10893,N_11840);
and U13689 (N_13689,N_10007,N_10394);
xor U13690 (N_13690,N_11451,N_11997);
xor U13691 (N_13691,N_11082,N_10388);
or U13692 (N_13692,N_10691,N_10763);
nand U13693 (N_13693,N_11347,N_11128);
xnor U13694 (N_13694,N_11559,N_10074);
nand U13695 (N_13695,N_10005,N_10607);
xor U13696 (N_13696,N_11011,N_10874);
nor U13697 (N_13697,N_10936,N_10043);
nand U13698 (N_13698,N_10724,N_10897);
or U13699 (N_13699,N_11933,N_10232);
nand U13700 (N_13700,N_11518,N_11232);
xor U13701 (N_13701,N_11027,N_11581);
and U13702 (N_13702,N_11584,N_10305);
or U13703 (N_13703,N_10875,N_11159);
or U13704 (N_13704,N_11224,N_11977);
and U13705 (N_13705,N_11888,N_11467);
or U13706 (N_13706,N_10572,N_10053);
and U13707 (N_13707,N_10216,N_10875);
or U13708 (N_13708,N_10742,N_11922);
nor U13709 (N_13709,N_10066,N_11806);
or U13710 (N_13710,N_11130,N_11831);
nand U13711 (N_13711,N_10347,N_10115);
and U13712 (N_13712,N_11866,N_10693);
or U13713 (N_13713,N_10065,N_10276);
nor U13714 (N_13714,N_10545,N_11771);
nand U13715 (N_13715,N_11994,N_10880);
or U13716 (N_13716,N_11016,N_10290);
nor U13717 (N_13717,N_11730,N_10318);
nand U13718 (N_13718,N_11033,N_10166);
or U13719 (N_13719,N_10798,N_11163);
and U13720 (N_13720,N_11429,N_10367);
nand U13721 (N_13721,N_11066,N_11352);
nor U13722 (N_13722,N_10295,N_11944);
xor U13723 (N_13723,N_11745,N_11146);
or U13724 (N_13724,N_11949,N_10029);
or U13725 (N_13725,N_10908,N_10559);
and U13726 (N_13726,N_11839,N_10147);
xnor U13727 (N_13727,N_10960,N_11357);
or U13728 (N_13728,N_10850,N_10974);
or U13729 (N_13729,N_11500,N_11759);
and U13730 (N_13730,N_11973,N_11197);
nand U13731 (N_13731,N_10575,N_10126);
xnor U13732 (N_13732,N_11813,N_11189);
or U13733 (N_13733,N_11408,N_11368);
xor U13734 (N_13734,N_11954,N_11878);
nor U13735 (N_13735,N_10342,N_10011);
xnor U13736 (N_13736,N_11221,N_11308);
nor U13737 (N_13737,N_11025,N_10718);
nor U13738 (N_13738,N_11020,N_11424);
and U13739 (N_13739,N_10850,N_10858);
or U13740 (N_13740,N_10965,N_10350);
nand U13741 (N_13741,N_10076,N_10557);
or U13742 (N_13742,N_10113,N_10252);
xnor U13743 (N_13743,N_10857,N_10660);
or U13744 (N_13744,N_11400,N_10418);
and U13745 (N_13745,N_10912,N_10138);
xor U13746 (N_13746,N_11825,N_10844);
or U13747 (N_13747,N_11091,N_10810);
and U13748 (N_13748,N_10439,N_11155);
nor U13749 (N_13749,N_11019,N_11267);
xnor U13750 (N_13750,N_11017,N_10879);
or U13751 (N_13751,N_11426,N_10145);
xor U13752 (N_13752,N_11086,N_10491);
or U13753 (N_13753,N_11905,N_10227);
or U13754 (N_13754,N_10670,N_10479);
or U13755 (N_13755,N_11591,N_11124);
nor U13756 (N_13756,N_11383,N_11493);
nand U13757 (N_13757,N_11844,N_10522);
and U13758 (N_13758,N_11042,N_10718);
or U13759 (N_13759,N_11055,N_11530);
xnor U13760 (N_13760,N_10137,N_11923);
and U13761 (N_13761,N_10935,N_11553);
nand U13762 (N_13762,N_10524,N_10439);
xor U13763 (N_13763,N_11368,N_11809);
xor U13764 (N_13764,N_11984,N_10264);
and U13765 (N_13765,N_11239,N_11857);
nand U13766 (N_13766,N_10053,N_10657);
and U13767 (N_13767,N_11667,N_11506);
nor U13768 (N_13768,N_11000,N_11724);
and U13769 (N_13769,N_11731,N_10537);
nand U13770 (N_13770,N_11935,N_10416);
nand U13771 (N_13771,N_11825,N_10508);
or U13772 (N_13772,N_10648,N_10114);
and U13773 (N_13773,N_10725,N_11212);
xnor U13774 (N_13774,N_11012,N_11033);
or U13775 (N_13775,N_10056,N_10790);
nor U13776 (N_13776,N_11444,N_11102);
or U13777 (N_13777,N_11522,N_10536);
and U13778 (N_13778,N_11279,N_10223);
nor U13779 (N_13779,N_10152,N_11814);
xnor U13780 (N_13780,N_11610,N_11840);
nor U13781 (N_13781,N_11316,N_11717);
xor U13782 (N_13782,N_11046,N_10037);
xor U13783 (N_13783,N_11612,N_11737);
and U13784 (N_13784,N_11021,N_11624);
nor U13785 (N_13785,N_10743,N_10355);
nand U13786 (N_13786,N_11763,N_10203);
xor U13787 (N_13787,N_10408,N_11904);
or U13788 (N_13788,N_10387,N_11682);
and U13789 (N_13789,N_11678,N_11140);
or U13790 (N_13790,N_11426,N_10733);
or U13791 (N_13791,N_11216,N_10632);
or U13792 (N_13792,N_10685,N_10280);
and U13793 (N_13793,N_11980,N_10184);
nand U13794 (N_13794,N_10091,N_10482);
nand U13795 (N_13795,N_10807,N_11736);
nor U13796 (N_13796,N_10958,N_10246);
nand U13797 (N_13797,N_11816,N_10789);
nor U13798 (N_13798,N_10445,N_10903);
or U13799 (N_13799,N_10536,N_11386);
nand U13800 (N_13800,N_10272,N_10499);
xor U13801 (N_13801,N_10948,N_10199);
nand U13802 (N_13802,N_10805,N_10506);
nand U13803 (N_13803,N_11161,N_11005);
and U13804 (N_13804,N_11848,N_11209);
nand U13805 (N_13805,N_10576,N_10727);
nor U13806 (N_13806,N_11174,N_11300);
nor U13807 (N_13807,N_11506,N_10738);
xor U13808 (N_13808,N_10799,N_10173);
xnor U13809 (N_13809,N_10198,N_10154);
xnor U13810 (N_13810,N_10973,N_10747);
xnor U13811 (N_13811,N_10883,N_11049);
nor U13812 (N_13812,N_11817,N_11841);
xor U13813 (N_13813,N_10157,N_10596);
or U13814 (N_13814,N_10922,N_10046);
nor U13815 (N_13815,N_11776,N_10044);
nand U13816 (N_13816,N_10075,N_10387);
and U13817 (N_13817,N_11825,N_10132);
xor U13818 (N_13818,N_10941,N_10761);
nor U13819 (N_13819,N_10151,N_10903);
and U13820 (N_13820,N_11135,N_10584);
or U13821 (N_13821,N_10204,N_11957);
and U13822 (N_13822,N_10710,N_11200);
nand U13823 (N_13823,N_10353,N_10823);
nand U13824 (N_13824,N_10592,N_10037);
nor U13825 (N_13825,N_11645,N_10676);
nand U13826 (N_13826,N_10000,N_11855);
and U13827 (N_13827,N_10086,N_10660);
or U13828 (N_13828,N_11339,N_11546);
xnor U13829 (N_13829,N_11202,N_10686);
xor U13830 (N_13830,N_10068,N_11977);
nor U13831 (N_13831,N_10507,N_11617);
xnor U13832 (N_13832,N_10357,N_10764);
nand U13833 (N_13833,N_10682,N_10861);
nor U13834 (N_13834,N_11099,N_11826);
and U13835 (N_13835,N_11169,N_11241);
nand U13836 (N_13836,N_10253,N_10848);
or U13837 (N_13837,N_10428,N_10090);
and U13838 (N_13838,N_11345,N_11421);
and U13839 (N_13839,N_11534,N_10145);
and U13840 (N_13840,N_11530,N_11619);
nand U13841 (N_13841,N_10362,N_10330);
or U13842 (N_13842,N_11452,N_10967);
nand U13843 (N_13843,N_11919,N_10106);
nand U13844 (N_13844,N_11808,N_11598);
nand U13845 (N_13845,N_10814,N_11863);
or U13846 (N_13846,N_11236,N_11607);
and U13847 (N_13847,N_11238,N_10630);
nor U13848 (N_13848,N_10349,N_11463);
nand U13849 (N_13849,N_11662,N_11747);
nand U13850 (N_13850,N_10221,N_11954);
nand U13851 (N_13851,N_11978,N_10209);
nor U13852 (N_13852,N_10289,N_10086);
nand U13853 (N_13853,N_11264,N_10580);
and U13854 (N_13854,N_10870,N_11660);
or U13855 (N_13855,N_11903,N_11731);
nor U13856 (N_13856,N_10245,N_11217);
nor U13857 (N_13857,N_10468,N_10690);
xnor U13858 (N_13858,N_10312,N_10825);
and U13859 (N_13859,N_10324,N_10557);
xnor U13860 (N_13860,N_10450,N_10580);
nand U13861 (N_13861,N_10467,N_11541);
and U13862 (N_13862,N_11015,N_11021);
and U13863 (N_13863,N_11073,N_10917);
nor U13864 (N_13864,N_11885,N_11354);
nand U13865 (N_13865,N_11032,N_11284);
and U13866 (N_13866,N_11939,N_10918);
nand U13867 (N_13867,N_10366,N_10120);
xor U13868 (N_13868,N_11578,N_11059);
xor U13869 (N_13869,N_10336,N_11591);
and U13870 (N_13870,N_10100,N_10857);
nand U13871 (N_13871,N_10978,N_10781);
nand U13872 (N_13872,N_10073,N_10357);
nor U13873 (N_13873,N_10079,N_10919);
xnor U13874 (N_13874,N_11457,N_11600);
or U13875 (N_13875,N_11227,N_10644);
nor U13876 (N_13876,N_11684,N_10498);
nor U13877 (N_13877,N_10935,N_10998);
or U13878 (N_13878,N_11448,N_10208);
and U13879 (N_13879,N_10960,N_11656);
xnor U13880 (N_13880,N_10519,N_10848);
nor U13881 (N_13881,N_10570,N_10615);
nand U13882 (N_13882,N_11033,N_11408);
xor U13883 (N_13883,N_11354,N_10823);
and U13884 (N_13884,N_11269,N_11321);
and U13885 (N_13885,N_10569,N_10122);
xor U13886 (N_13886,N_11398,N_11295);
nor U13887 (N_13887,N_11038,N_10012);
nor U13888 (N_13888,N_10021,N_11490);
xor U13889 (N_13889,N_11221,N_11142);
xor U13890 (N_13890,N_11471,N_11166);
nand U13891 (N_13891,N_11409,N_11407);
xor U13892 (N_13892,N_11717,N_11196);
or U13893 (N_13893,N_10731,N_11748);
nor U13894 (N_13894,N_11675,N_11465);
or U13895 (N_13895,N_11188,N_10042);
or U13896 (N_13896,N_11695,N_10200);
nor U13897 (N_13897,N_10243,N_11524);
nor U13898 (N_13898,N_11889,N_10884);
nand U13899 (N_13899,N_11925,N_10731);
or U13900 (N_13900,N_10782,N_11620);
and U13901 (N_13901,N_10990,N_11362);
xor U13902 (N_13902,N_11214,N_11367);
or U13903 (N_13903,N_11663,N_10310);
nor U13904 (N_13904,N_11590,N_11475);
nand U13905 (N_13905,N_10095,N_11040);
nand U13906 (N_13906,N_10601,N_11505);
nor U13907 (N_13907,N_11122,N_10545);
or U13908 (N_13908,N_10269,N_11207);
and U13909 (N_13909,N_10320,N_11986);
nor U13910 (N_13910,N_11884,N_11397);
xnor U13911 (N_13911,N_10107,N_10562);
nand U13912 (N_13912,N_10108,N_11402);
nor U13913 (N_13913,N_10098,N_11207);
nor U13914 (N_13914,N_10353,N_11800);
or U13915 (N_13915,N_10775,N_10517);
xor U13916 (N_13916,N_10471,N_10348);
nand U13917 (N_13917,N_11185,N_10656);
and U13918 (N_13918,N_11177,N_10761);
xor U13919 (N_13919,N_10091,N_10525);
nand U13920 (N_13920,N_11891,N_10708);
xor U13921 (N_13921,N_11062,N_11008);
nor U13922 (N_13922,N_11192,N_11277);
nor U13923 (N_13923,N_11376,N_10151);
nor U13924 (N_13924,N_10273,N_11956);
or U13925 (N_13925,N_11565,N_10348);
nand U13926 (N_13926,N_10489,N_11883);
nand U13927 (N_13927,N_11927,N_10044);
and U13928 (N_13928,N_10059,N_10785);
xor U13929 (N_13929,N_10791,N_11750);
nor U13930 (N_13930,N_10473,N_11015);
and U13931 (N_13931,N_11622,N_10584);
or U13932 (N_13932,N_10225,N_11403);
and U13933 (N_13933,N_11419,N_10564);
and U13934 (N_13934,N_10684,N_10250);
xor U13935 (N_13935,N_10706,N_10040);
nor U13936 (N_13936,N_10556,N_11388);
nor U13937 (N_13937,N_10664,N_10968);
or U13938 (N_13938,N_10295,N_10161);
xnor U13939 (N_13939,N_10309,N_11435);
xnor U13940 (N_13940,N_11162,N_11023);
nand U13941 (N_13941,N_11924,N_10142);
nand U13942 (N_13942,N_10527,N_11596);
or U13943 (N_13943,N_10037,N_11553);
nor U13944 (N_13944,N_11568,N_10929);
nand U13945 (N_13945,N_11538,N_10888);
nor U13946 (N_13946,N_11465,N_10242);
and U13947 (N_13947,N_10871,N_11662);
or U13948 (N_13948,N_11421,N_10200);
and U13949 (N_13949,N_11557,N_10238);
nor U13950 (N_13950,N_10634,N_10457);
or U13951 (N_13951,N_11018,N_11744);
xnor U13952 (N_13952,N_11745,N_10444);
or U13953 (N_13953,N_11526,N_11389);
nor U13954 (N_13954,N_10210,N_11040);
xor U13955 (N_13955,N_10390,N_10236);
or U13956 (N_13956,N_11073,N_11951);
nand U13957 (N_13957,N_11020,N_11607);
or U13958 (N_13958,N_10867,N_11101);
nor U13959 (N_13959,N_11549,N_10442);
nand U13960 (N_13960,N_11737,N_10299);
nand U13961 (N_13961,N_10106,N_10327);
or U13962 (N_13962,N_10457,N_10955);
and U13963 (N_13963,N_10455,N_10203);
xnor U13964 (N_13964,N_10727,N_10055);
and U13965 (N_13965,N_10625,N_11125);
nor U13966 (N_13966,N_11024,N_11801);
xnor U13967 (N_13967,N_11010,N_11261);
nor U13968 (N_13968,N_11239,N_11737);
or U13969 (N_13969,N_11859,N_11625);
or U13970 (N_13970,N_10327,N_11395);
nor U13971 (N_13971,N_11192,N_11388);
and U13972 (N_13972,N_10663,N_11314);
xnor U13973 (N_13973,N_10660,N_11863);
nor U13974 (N_13974,N_10431,N_10598);
nand U13975 (N_13975,N_11233,N_11074);
nor U13976 (N_13976,N_11489,N_11746);
xnor U13977 (N_13977,N_10131,N_11499);
and U13978 (N_13978,N_10098,N_11228);
nor U13979 (N_13979,N_10371,N_10263);
nor U13980 (N_13980,N_10508,N_10832);
and U13981 (N_13981,N_11187,N_10104);
nand U13982 (N_13982,N_11989,N_10139);
nand U13983 (N_13983,N_10887,N_10085);
xor U13984 (N_13984,N_11629,N_11879);
and U13985 (N_13985,N_10701,N_11580);
nor U13986 (N_13986,N_10912,N_11752);
xor U13987 (N_13987,N_10741,N_11826);
nand U13988 (N_13988,N_10555,N_10909);
nor U13989 (N_13989,N_11930,N_11278);
nand U13990 (N_13990,N_10835,N_11245);
nand U13991 (N_13991,N_10276,N_10494);
nand U13992 (N_13992,N_11930,N_10134);
nor U13993 (N_13993,N_11966,N_11734);
nor U13994 (N_13994,N_11322,N_11962);
and U13995 (N_13995,N_10424,N_11883);
and U13996 (N_13996,N_10418,N_11755);
xnor U13997 (N_13997,N_11875,N_11346);
and U13998 (N_13998,N_11758,N_11930);
or U13999 (N_13999,N_11907,N_10599);
nand U14000 (N_14000,N_12469,N_13166);
or U14001 (N_14001,N_12937,N_13076);
nand U14002 (N_14002,N_12644,N_12302);
and U14003 (N_14003,N_13434,N_12732);
xnor U14004 (N_14004,N_12497,N_12114);
nand U14005 (N_14005,N_13092,N_12250);
or U14006 (N_14006,N_13230,N_13521);
and U14007 (N_14007,N_13457,N_12776);
and U14008 (N_14008,N_12981,N_12213);
and U14009 (N_14009,N_12459,N_12040);
nor U14010 (N_14010,N_13644,N_12178);
nor U14011 (N_14011,N_12032,N_12803);
and U14012 (N_14012,N_13273,N_13961);
or U14013 (N_14013,N_12074,N_13259);
and U14014 (N_14014,N_13715,N_12791);
nand U14015 (N_14015,N_13677,N_13548);
or U14016 (N_14016,N_13950,N_13240);
or U14017 (N_14017,N_13889,N_13121);
nor U14018 (N_14018,N_13135,N_13160);
and U14019 (N_14019,N_12815,N_12544);
xor U14020 (N_14020,N_13806,N_12617);
xnor U14021 (N_14021,N_13069,N_13948);
or U14022 (N_14022,N_12322,N_12682);
nor U14023 (N_14023,N_12821,N_13564);
nand U14024 (N_14024,N_12916,N_12901);
or U14025 (N_14025,N_12249,N_13312);
nor U14026 (N_14026,N_12278,N_13262);
nand U14027 (N_14027,N_12387,N_13243);
and U14028 (N_14028,N_13481,N_12830);
nand U14029 (N_14029,N_12300,N_12643);
nor U14030 (N_14030,N_13223,N_13460);
nor U14031 (N_14031,N_12840,N_13971);
xor U14032 (N_14032,N_12903,N_12319);
xor U14033 (N_14033,N_12312,N_12079);
nand U14034 (N_14034,N_13790,N_12926);
nor U14035 (N_14035,N_13404,N_13744);
or U14036 (N_14036,N_12404,N_12875);
or U14037 (N_14037,N_13400,N_13826);
nor U14038 (N_14038,N_13559,N_12675);
nand U14039 (N_14039,N_12608,N_12228);
or U14040 (N_14040,N_12772,N_12487);
and U14041 (N_14041,N_12863,N_13053);
and U14042 (N_14042,N_13929,N_12296);
nor U14043 (N_14043,N_12514,N_13307);
nor U14044 (N_14044,N_12509,N_12236);
or U14045 (N_14045,N_12798,N_12021);
xnor U14046 (N_14046,N_12076,N_12508);
xnor U14047 (N_14047,N_13317,N_13784);
nand U14048 (N_14048,N_12000,N_13084);
xnor U14049 (N_14049,N_12031,N_12323);
nand U14050 (N_14050,N_12861,N_13853);
and U14051 (N_14051,N_13396,N_12072);
nor U14052 (N_14052,N_13804,N_12271);
nor U14053 (N_14053,N_13114,N_13492);
or U14054 (N_14054,N_13747,N_13174);
xnor U14055 (N_14055,N_13546,N_12671);
and U14056 (N_14056,N_12519,N_13222);
or U14057 (N_14057,N_13995,N_13242);
or U14058 (N_14058,N_12832,N_13377);
xor U14059 (N_14059,N_12719,N_12504);
nor U14060 (N_14060,N_12460,N_12596);
xnor U14061 (N_14061,N_13118,N_12698);
or U14062 (N_14062,N_13721,N_13567);
xnor U14063 (N_14063,N_12649,N_13392);
nand U14064 (N_14064,N_13869,N_13505);
or U14065 (N_14065,N_12217,N_12131);
xnor U14066 (N_14066,N_13329,N_13414);
nand U14067 (N_14067,N_12011,N_13541);
xor U14068 (N_14068,N_13027,N_12016);
nand U14069 (N_14069,N_13447,N_12789);
and U14070 (N_14070,N_13682,N_12913);
or U14071 (N_14071,N_12150,N_12727);
and U14072 (N_14072,N_13822,N_13295);
nand U14073 (N_14073,N_12570,N_13599);
or U14074 (N_14074,N_12135,N_12914);
and U14075 (N_14075,N_12951,N_13198);
and U14076 (N_14076,N_12679,N_13023);
xnor U14077 (N_14077,N_13107,N_13164);
nand U14078 (N_14078,N_12680,N_12492);
or U14079 (N_14079,N_13290,N_12355);
xor U14080 (N_14080,N_13570,N_13299);
nor U14081 (N_14081,N_13407,N_12775);
or U14082 (N_14082,N_13871,N_13241);
or U14083 (N_14083,N_13751,N_13438);
and U14084 (N_14084,N_13415,N_12491);
nand U14085 (N_14085,N_13814,N_13729);
xnor U14086 (N_14086,N_13960,N_12411);
xor U14087 (N_14087,N_12804,N_12802);
or U14088 (N_14088,N_12080,N_13476);
nor U14089 (N_14089,N_13921,N_13040);
and U14090 (N_14090,N_13805,N_13630);
nor U14091 (N_14091,N_12028,N_12851);
or U14092 (N_14092,N_12368,N_13458);
nor U14093 (N_14093,N_12026,N_12988);
nand U14094 (N_14094,N_12974,N_12320);
nor U14095 (N_14095,N_12728,N_12159);
nand U14096 (N_14096,N_13202,N_13470);
xnor U14097 (N_14097,N_13618,N_12256);
nor U14098 (N_14098,N_12234,N_13193);
and U14099 (N_14099,N_13293,N_12690);
nand U14100 (N_14100,N_12485,N_12505);
nand U14101 (N_14101,N_12102,N_12545);
and U14102 (N_14102,N_12556,N_13823);
xnor U14103 (N_14103,N_12393,N_13436);
xnor U14104 (N_14104,N_13879,N_12670);
or U14105 (N_14105,N_13776,N_12450);
xnor U14106 (N_14106,N_13713,N_12513);
nand U14107 (N_14107,N_12412,N_13339);
nand U14108 (N_14108,N_13761,N_13072);
and U14109 (N_14109,N_13621,N_12950);
nand U14110 (N_14110,N_13342,N_13659);
nand U14111 (N_14111,N_13900,N_12037);
and U14112 (N_14112,N_12154,N_12087);
nor U14113 (N_14113,N_12241,N_12876);
nor U14114 (N_14114,N_13922,N_13172);
xor U14115 (N_14115,N_13522,N_12639);
nor U14116 (N_14116,N_12085,N_13746);
xnor U14117 (N_14117,N_12609,N_13707);
or U14118 (N_14118,N_13571,N_13149);
or U14119 (N_14119,N_12543,N_12632);
or U14120 (N_14120,N_12731,N_12942);
nor U14121 (N_14121,N_12326,N_13895);
nand U14122 (N_14122,N_13066,N_13783);
and U14123 (N_14123,N_12162,N_13412);
and U14124 (N_14124,N_12814,N_12986);
xor U14125 (N_14125,N_13516,N_12663);
nand U14126 (N_14126,N_12051,N_12449);
and U14127 (N_14127,N_12052,N_13877);
xnor U14128 (N_14128,N_12893,N_12344);
or U14129 (N_14129,N_13782,N_12822);
nor U14130 (N_14130,N_12111,N_12963);
and U14131 (N_14131,N_13433,N_13647);
and U14132 (N_14132,N_13285,N_13300);
and U14133 (N_14133,N_12416,N_12027);
nor U14134 (N_14134,N_13723,N_12940);
and U14135 (N_14135,N_13777,N_13082);
and U14136 (N_14136,N_12155,N_13815);
and U14137 (N_14137,N_13423,N_12381);
xnor U14138 (N_14138,N_13833,N_12751);
nor U14139 (N_14139,N_13544,N_12467);
nand U14140 (N_14140,N_12613,N_13637);
xor U14141 (N_14141,N_12226,N_13055);
nor U14142 (N_14142,N_13552,N_13327);
nor U14143 (N_14143,N_12837,N_13781);
nor U14144 (N_14144,N_12805,N_12747);
or U14145 (N_14145,N_12142,N_13156);
and U14146 (N_14146,N_13035,N_13153);
nor U14147 (N_14147,N_12126,N_13456);
or U14148 (N_14148,N_13416,N_12269);
or U14149 (N_14149,N_13020,N_12753);
nand U14150 (N_14150,N_12436,N_13606);
xor U14151 (N_14151,N_13937,N_13945);
or U14152 (N_14152,N_12023,N_13737);
xor U14153 (N_14153,N_12253,N_13575);
and U14154 (N_14154,N_12567,N_13191);
xnor U14155 (N_14155,N_13788,N_13633);
nor U14156 (N_14156,N_13534,N_13225);
nand U14157 (N_14157,N_12985,N_12407);
nand U14158 (N_14158,N_12835,N_13827);
or U14159 (N_14159,N_12646,N_12169);
xnor U14160 (N_14160,N_13667,N_13828);
nand U14161 (N_14161,N_12859,N_13399);
or U14162 (N_14162,N_13562,N_13572);
and U14163 (N_14163,N_12633,N_12536);
nand U14164 (N_14164,N_13021,N_12919);
nor U14165 (N_14165,N_12252,N_13275);
or U14166 (N_14166,N_13305,N_12959);
xor U14167 (N_14167,N_12763,N_12336);
or U14168 (N_14168,N_12257,N_12309);
xnor U14169 (N_14169,N_13213,N_12086);
xor U14170 (N_14170,N_12419,N_12599);
xnor U14171 (N_14171,N_12677,N_12918);
nor U14172 (N_14172,N_12097,N_12168);
xor U14173 (N_14173,N_12899,N_13856);
or U14174 (N_14174,N_13897,N_13532);
nor U14175 (N_14175,N_13904,N_13626);
nor U14176 (N_14176,N_12904,N_13812);
and U14177 (N_14177,N_12780,N_12328);
xor U14178 (N_14178,N_12306,N_12025);
nand U14179 (N_14179,N_12141,N_13654);
nand U14180 (N_14180,N_12165,N_12113);
nand U14181 (N_14181,N_13585,N_13173);
nand U14182 (N_14182,N_13763,N_13170);
xnor U14183 (N_14183,N_12934,N_13311);
xor U14184 (N_14184,N_13683,N_13286);
or U14185 (N_14185,N_13801,N_13657);
nor U14186 (N_14186,N_12330,N_13254);
nand U14187 (N_14187,N_13607,N_13093);
or U14188 (N_14188,N_12321,N_13731);
xnor U14189 (N_14189,N_12554,N_13590);
nor U14190 (N_14190,N_13942,N_13378);
nand U14191 (N_14191,N_12083,N_12706);
and U14192 (N_14192,N_12542,N_13050);
xor U14193 (N_14193,N_12243,N_13270);
nand U14194 (N_14194,N_12860,N_13775);
nand U14195 (N_14195,N_12882,N_12013);
nor U14196 (N_14196,N_12635,N_13386);
nand U14197 (N_14197,N_12852,N_13966);
or U14198 (N_14198,N_12537,N_12696);
xor U14199 (N_14199,N_12069,N_12827);
and U14200 (N_14200,N_13760,N_13561);
nor U14201 (N_14201,N_12692,N_12370);
nor U14202 (N_14202,N_12809,N_13229);
nand U14203 (N_14203,N_13725,N_13450);
and U14204 (N_14204,N_12406,N_13183);
nand U14205 (N_14205,N_12889,N_12057);
or U14206 (N_14206,N_12399,N_13056);
nor U14207 (N_14207,N_13033,N_13435);
xnor U14208 (N_14208,N_12784,N_13375);
xor U14209 (N_14209,N_13287,N_13753);
or U14210 (N_14210,N_13640,N_13694);
nor U14211 (N_14211,N_13100,N_13067);
nand U14212 (N_14212,N_12693,N_13324);
nand U14213 (N_14213,N_12510,N_13990);
and U14214 (N_14214,N_12180,N_13926);
xor U14215 (N_14215,N_13261,N_12983);
or U14216 (N_14216,N_13049,N_12838);
xor U14217 (N_14217,N_12365,N_12088);
and U14218 (N_14218,N_12925,N_13113);
nand U14219 (N_14219,N_13832,N_13045);
and U14220 (N_14220,N_12287,N_12530);
or U14221 (N_14221,N_13065,N_13646);
or U14222 (N_14222,N_13750,N_13260);
or U14223 (N_14223,N_13078,N_13103);
or U14224 (N_14224,N_12230,N_12118);
xnor U14225 (N_14225,N_13870,N_12558);
nor U14226 (N_14226,N_12210,N_12045);
or U14227 (N_14227,N_12127,N_12931);
or U14228 (N_14228,N_13829,N_12396);
nor U14229 (N_14229,N_13362,N_13908);
xnor U14230 (N_14230,N_13976,N_13837);
or U14231 (N_14231,N_13130,N_12790);
nand U14232 (N_14232,N_13789,N_12261);
nand U14233 (N_14233,N_13802,N_13787);
nand U14234 (N_14234,N_13000,N_12285);
xnor U14235 (N_14235,N_12588,N_13062);
and U14236 (N_14236,N_13461,N_12035);
and U14237 (N_14237,N_12546,N_13793);
or U14238 (N_14238,N_12655,N_12310);
nand U14239 (N_14239,N_13119,N_12359);
and U14240 (N_14240,N_13664,N_12434);
xor U14241 (N_14241,N_12585,N_12055);
nor U14242 (N_14242,N_13180,N_13741);
or U14243 (N_14243,N_12066,N_13308);
nand U14244 (N_14244,N_13127,N_12157);
nor U14245 (N_14245,N_13155,N_13724);
xnor U14246 (N_14246,N_12197,N_13818);
and U14247 (N_14247,N_13611,N_13026);
or U14248 (N_14248,N_12064,N_12147);
and U14249 (N_14249,N_12200,N_12220);
nor U14250 (N_14250,N_13733,N_13722);
and U14251 (N_14251,N_13351,N_12960);
or U14252 (N_14252,N_12970,N_13419);
and U14253 (N_14253,N_13593,N_12511);
xor U14254 (N_14254,N_13304,N_13653);
and U14255 (N_14255,N_13680,N_13124);
xor U14256 (N_14256,N_13199,N_12823);
or U14257 (N_14257,N_12140,N_13573);
nand U14258 (N_14258,N_13880,N_13380);
or U14259 (N_14259,N_12561,N_13218);
nand U14260 (N_14260,N_12992,N_12977);
or U14261 (N_14261,N_13578,N_12318);
nor U14262 (N_14262,N_12722,N_12465);
and U14263 (N_14263,N_12939,N_12283);
xor U14264 (N_14264,N_13325,N_12954);
nand U14265 (N_14265,N_12070,N_13002);
nor U14266 (N_14266,N_13323,N_12255);
or U14267 (N_14267,N_12203,N_12428);
nor U14268 (N_14268,N_12922,N_13088);
nand U14269 (N_14269,N_13666,N_13201);
nand U14270 (N_14270,N_12651,N_13779);
nand U14271 (N_14271,N_12705,N_12816);
or U14272 (N_14272,N_12908,N_12844);
or U14273 (N_14273,N_13385,N_12059);
xor U14274 (N_14274,N_12186,N_12833);
xor U14275 (N_14275,N_13907,N_13686);
or U14276 (N_14276,N_12669,N_13893);
or U14277 (N_14277,N_12557,N_12195);
nor U14278 (N_14278,N_12700,N_13511);
or U14279 (N_14279,N_12817,N_12749);
nor U14280 (N_14280,N_13129,N_12628);
xnor U14281 (N_14281,N_13147,N_13167);
and U14282 (N_14282,N_12311,N_13389);
nand U14283 (N_14283,N_12892,N_12347);
nor U14284 (N_14284,N_13996,N_13690);
and U14285 (N_14285,N_12437,N_12762);
nand U14286 (N_14286,N_12806,N_12621);
or U14287 (N_14287,N_12389,N_12515);
or U14288 (N_14288,N_13219,N_13648);
and U14289 (N_14289,N_12795,N_13175);
nor U14290 (N_14290,N_12340,N_13350);
and U14291 (N_14291,N_13533,N_12291);
nor U14292 (N_14292,N_12461,N_12601);
xor U14293 (N_14293,N_12642,N_13662);
nand U14294 (N_14294,N_12998,N_12181);
nand U14295 (N_14295,N_12115,N_13528);
or U14296 (N_14296,N_13315,N_12092);
and U14297 (N_14297,N_13036,N_13489);
nor U14298 (N_14298,N_13704,N_13310);
or U14299 (N_14299,N_12448,N_12167);
and U14300 (N_14300,N_13140,N_12936);
or U14301 (N_14301,N_13268,N_12501);
and U14302 (N_14302,N_13972,N_13239);
and U14303 (N_14303,N_12648,N_12660);
or U14304 (N_14304,N_12418,N_13263);
and U14305 (N_14305,N_12123,N_13057);
and U14306 (N_14306,N_12584,N_12778);
or U14307 (N_14307,N_12474,N_12071);
and U14308 (N_14308,N_12575,N_13309);
nand U14309 (N_14309,N_12267,N_13196);
nand U14310 (N_14310,N_12125,N_13152);
and U14311 (N_14311,N_13282,N_12440);
nand U14312 (N_14312,N_13513,N_12729);
nor U14313 (N_14313,N_12033,N_13719);
nor U14314 (N_14314,N_12622,N_13594);
and U14315 (N_14315,N_13509,N_12238);
xor U14316 (N_14316,N_13137,N_12292);
nand U14317 (N_14317,N_12341,N_12752);
and U14318 (N_14318,N_13011,N_12290);
xnor U14319 (N_14319,N_12388,N_13393);
and U14320 (N_14320,N_12979,N_12522);
nor U14321 (N_14321,N_12014,N_13859);
or U14322 (N_14322,N_13558,N_12078);
and U14323 (N_14323,N_12563,N_12315);
or U14324 (N_14324,N_13452,N_12850);
xor U14325 (N_14325,N_12104,N_13817);
and U14326 (N_14326,N_12382,N_12402);
nand U14327 (N_14327,N_13501,N_12061);
or U14328 (N_14328,N_12246,N_13421);
or U14329 (N_14329,N_12653,N_12041);
xnor U14330 (N_14330,N_13864,N_12855);
or U14331 (N_14331,N_12376,N_13099);
nand U14332 (N_14332,N_13910,N_13272);
nand U14333 (N_14333,N_13264,N_12877);
nor U14334 (N_14334,N_12219,N_12552);
nor U14335 (N_14335,N_13221,N_13369);
and U14336 (N_14336,N_12880,N_13493);
nand U14337 (N_14337,N_12338,N_13244);
or U14338 (N_14338,N_12777,N_13549);
or U14339 (N_14339,N_13215,N_12204);
and U14340 (N_14340,N_13269,N_13700);
xnor U14341 (N_14341,N_13687,N_13769);
xnor U14342 (N_14342,N_13034,N_12191);
or U14343 (N_14343,N_13208,N_12075);
xor U14344 (N_14344,N_12119,N_13234);
xnor U14345 (N_14345,N_13361,N_12174);
nor U14346 (N_14346,N_12573,N_13896);
nand U14347 (N_14347,N_13437,N_12024);
and U14348 (N_14348,N_12160,N_12688);
or U14349 (N_14349,N_13906,N_13184);
nor U14350 (N_14350,N_12587,N_13515);
nand U14351 (N_14351,N_13394,N_13890);
or U14352 (N_14352,N_12152,N_13925);
nor U14353 (N_14353,N_12371,N_13774);
nand U14354 (N_14354,N_13740,N_13278);
nand U14355 (N_14355,N_13197,N_12392);
nand U14356 (N_14356,N_12483,N_12435);
nand U14357 (N_14357,N_12709,N_13614);
xor U14358 (N_14358,N_13070,N_13338);
nand U14359 (N_14359,N_13060,N_13255);
nand U14360 (N_14360,N_12484,N_13398);
nand U14361 (N_14361,N_12620,N_13531);
xnor U14362 (N_14362,N_13673,N_12030);
nor U14363 (N_14363,N_12581,N_12148);
nand U14364 (N_14364,N_12268,N_12957);
nor U14365 (N_14365,N_13624,N_13472);
nor U14366 (N_14366,N_12973,N_13671);
nand U14367 (N_14367,N_12808,N_13387);
or U14368 (N_14368,N_13809,N_13811);
nand U14369 (N_14369,N_12854,N_13109);
xnor U14370 (N_14370,N_12143,N_13794);
or U14371 (N_14371,N_13852,N_12225);
xor U14372 (N_14372,N_13795,N_12431);
xnor U14373 (N_14373,N_13987,N_12812);
nand U14374 (N_14374,N_13792,N_13917);
xor U14375 (N_14375,N_13200,N_13238);
xor U14376 (N_14376,N_12572,N_13813);
nand U14377 (N_14377,N_12503,N_12673);
or U14378 (N_14378,N_12629,N_12991);
xor U14379 (N_14379,N_12149,N_13302);
nand U14380 (N_14380,N_13185,N_12667);
xnor U14381 (N_14381,N_13181,N_13756);
nor U14382 (N_14382,N_13727,N_12579);
nor U14383 (N_14383,N_13508,N_12003);
and U14384 (N_14384,N_13402,N_13762);
nor U14385 (N_14385,N_12616,N_12886);
nor U14386 (N_14386,N_12890,N_12779);
xnor U14387 (N_14387,N_12891,N_12647);
xnor U14388 (N_14388,N_13095,N_13336);
and U14389 (N_14389,N_13898,N_12944);
nor U14390 (N_14390,N_13157,N_13353);
and U14391 (N_14391,N_12865,N_13847);
nor U14392 (N_14392,N_13554,N_13619);
nand U14393 (N_14393,N_12774,N_13656);
nand U14394 (N_14394,N_12451,N_13148);
xnor U14395 (N_14395,N_12410,N_12265);
or U14396 (N_14396,N_12116,N_13177);
nor U14397 (N_14397,N_12385,N_12718);
nand U14398 (N_14398,N_12745,N_12369);
nand U14399 (N_14399,N_12993,N_12361);
xor U14400 (N_14400,N_13963,N_12713);
xnor U14401 (N_14401,N_13403,N_12331);
xnor U14402 (N_14402,N_12980,N_13845);
xnor U14403 (N_14403,N_12695,N_12237);
xnor U14404 (N_14404,N_13003,N_12146);
nand U14405 (N_14405,N_13844,N_12879);
or U14406 (N_14406,N_13391,N_13451);
nor U14407 (N_14407,N_13277,N_12193);
and U14408 (N_14408,N_13785,N_12612);
or U14409 (N_14409,N_12233,N_12600);
and U14410 (N_14410,N_12473,N_12866);
nand U14411 (N_14411,N_12101,N_13888);
or U14412 (N_14412,N_13632,N_12819);
nor U14413 (N_14413,N_12058,N_12742);
and U14414 (N_14414,N_13772,N_13550);
nor U14415 (N_14415,N_12130,N_12773);
xor U14416 (N_14416,N_13974,N_13043);
nor U14417 (N_14417,N_12602,N_13106);
or U14418 (N_14418,N_13151,N_13894);
and U14419 (N_14419,N_13371,N_13709);
xnor U14420 (N_14420,N_12298,N_13138);
nor U14421 (N_14421,N_13267,N_13738);
xor U14422 (N_14422,N_13367,N_12641);
and U14423 (N_14423,N_12490,N_13952);
xor U14424 (N_14424,N_12699,N_13862);
xnor U14425 (N_14425,N_13981,N_12888);
nor U14426 (N_14426,N_13569,N_12175);
nor U14427 (N_14427,N_12357,N_13340);
nand U14428 (N_14428,N_13831,N_13883);
nor U14429 (N_14429,N_13360,N_13825);
nand U14430 (N_14430,N_12911,N_12128);
and U14431 (N_14431,N_13586,N_13498);
xnor U14432 (N_14432,N_12420,N_13112);
nand U14433 (N_14433,N_13949,N_12625);
nor U14434 (N_14434,N_12090,N_13993);
nand U14435 (N_14435,N_12205,N_13641);
and U14436 (N_14436,N_13605,N_12771);
or U14437 (N_14437,N_13796,N_13935);
nor U14438 (N_14438,N_12841,N_13867);
and U14439 (N_14439,N_13467,N_12524);
nor U14440 (N_14440,N_12124,N_12132);
nor U14441 (N_14441,N_13642,N_13226);
nor U14442 (N_14442,N_12921,N_12384);
nor U14443 (N_14443,N_13292,N_13886);
and U14444 (N_14444,N_12038,N_13728);
xor U14445 (N_14445,N_13600,N_12736);
or U14446 (N_14446,N_12770,N_13101);
nor U14447 (N_14447,N_13024,N_12864);
or U14448 (N_14448,N_13356,N_12439);
nor U14449 (N_14449,N_13587,N_13909);
xor U14450 (N_14450,N_13861,N_12928);
xnor U14451 (N_14451,N_12084,N_13406);
xnor U14452 (N_14452,N_13390,N_13136);
nor U14453 (N_14453,N_12631,N_13685);
or U14454 (N_14454,N_12093,N_12192);
nand U14455 (N_14455,N_12375,N_13485);
nor U14456 (N_14456,N_12568,N_13473);
nor U14457 (N_14457,N_12348,N_13410);
nand U14458 (N_14458,N_12094,N_13967);
or U14459 (N_14459,N_12173,N_12171);
and U14460 (N_14460,N_13601,N_13735);
nand U14461 (N_14461,N_12720,N_12839);
nor U14462 (N_14462,N_12189,N_13178);
nand U14463 (N_14463,N_13965,N_13233);
and U14464 (N_14464,N_12943,N_12475);
or U14465 (N_14465,N_12099,N_13408);
or U14466 (N_14466,N_13094,N_12560);
or U14467 (N_14467,N_13911,N_13517);
nand U14468 (N_14468,N_13316,N_13165);
and U14469 (N_14469,N_12276,N_12039);
or U14470 (N_14470,N_12592,N_12707);
or U14471 (N_14471,N_12949,N_13354);
or U14472 (N_14472,N_13502,N_12884);
nand U14473 (N_14473,N_12299,N_12920);
and U14474 (N_14474,N_13052,N_12067);
or U14475 (N_14475,N_12555,N_13758);
and U14476 (N_14476,N_12703,N_13595);
nand U14477 (N_14477,N_13163,N_12528);
or U14478 (N_14478,N_12871,N_12836);
and U14479 (N_14479,N_13171,N_12005);
nand U14480 (N_14480,N_13017,N_12060);
and U14481 (N_14481,N_13676,N_12144);
xor U14482 (N_14482,N_13246,N_12050);
nor U14483 (N_14483,N_13955,N_13631);
nor U14484 (N_14484,N_13999,N_13836);
xor U14485 (N_14485,N_12614,N_13959);
or U14486 (N_14486,N_13004,N_12792);
and U14487 (N_14487,N_12526,N_13835);
xor U14488 (N_14488,N_12636,N_13592);
or U14489 (N_14489,N_13405,N_13333);
or U14490 (N_14490,N_12329,N_13068);
nor U14491 (N_14491,N_12334,N_13645);
or U14492 (N_14492,N_12958,N_13840);
and U14493 (N_14493,N_12458,N_13834);
or U14494 (N_14494,N_12380,N_13210);
nand U14495 (N_14495,N_12972,N_12100);
nor U14496 (N_14496,N_13044,N_13527);
or U14497 (N_14497,N_13418,N_13444);
and U14498 (N_14498,N_13432,N_12533);
xor U14499 (N_14499,N_13660,N_12107);
and U14500 (N_14500,N_13250,N_12654);
nor U14501 (N_14501,N_13706,N_12349);
and U14502 (N_14502,N_13013,N_13359);
or U14503 (N_14503,N_13705,N_13691);
xor U14504 (N_14504,N_13349,N_12578);
or U14505 (N_14505,N_12231,N_13639);
nor U14506 (N_14506,N_13006,N_13576);
nor U14507 (N_14507,N_12507,N_12489);
nand U14508 (N_14508,N_12414,N_12493);
and U14509 (N_14509,N_13189,N_12289);
xnor U14510 (N_14510,N_12529,N_12665);
xnor U14511 (N_14511,N_13819,N_13670);
and U14512 (N_14512,N_13726,N_12756);
nand U14513 (N_14513,N_13957,N_13217);
and U14514 (N_14514,N_13698,N_12969);
and U14515 (N_14515,N_12978,N_13008);
xnor U14516 (N_14516,N_12303,N_12106);
xor U14517 (N_14517,N_13442,N_13982);
xor U14518 (N_14518,N_13372,N_12737);
xnor U14519 (N_14519,N_13334,N_12001);
nor U14520 (N_14520,N_12433,N_12820);
nand U14521 (N_14521,N_12623,N_13220);
nand U14522 (N_14522,N_12547,N_13711);
nor U14523 (N_14523,N_12208,N_12946);
and U14524 (N_14524,N_12179,N_12912);
nand U14525 (N_14525,N_13073,N_13048);
nand U14526 (N_14526,N_13479,N_12523);
or U14527 (N_14527,N_12807,N_13928);
nor U14528 (N_14528,N_13588,N_13855);
or U14529 (N_14529,N_13425,N_13730);
xor U14530 (N_14530,N_12307,N_12422);
or U14531 (N_14531,N_12787,N_12408);
or U14532 (N_14532,N_13542,N_13780);
and U14533 (N_14533,N_12758,N_12136);
and U14534 (N_14534,N_13978,N_13615);
nand U14535 (N_14535,N_13975,N_13009);
and U14536 (N_14536,N_13537,N_12878);
xor U14537 (N_14537,N_13565,N_12009);
and U14538 (N_14538,N_12740,N_12455);
xor U14539 (N_14539,N_12317,N_12353);
nor U14540 (N_14540,N_13116,N_13038);
xnor U14541 (N_14541,N_12046,N_12858);
nor U14542 (N_14542,N_13771,N_13204);
or U14543 (N_14543,N_13077,N_13486);
xnor U14544 (N_14544,N_12708,N_13347);
or U14545 (N_14545,N_12661,N_12681);
nor U14546 (N_14546,N_12842,N_12121);
and U14547 (N_14547,N_12337,N_12240);
nor U14548 (N_14548,N_12915,N_12694);
and U14549 (N_14549,N_12874,N_13440);
nor U14550 (N_14550,N_13037,N_12715);
nor U14551 (N_14551,N_12627,N_12927);
nor U14552 (N_14552,N_12272,N_13464);
xor U14553 (N_14553,N_12405,N_13046);
and U14554 (N_14554,N_12615,N_12481);
and U14555 (N_14555,N_12488,N_13441);
nand U14556 (N_14556,N_12945,N_13330);
or U14557 (N_14557,N_13271,N_12531);
nor U14558 (N_14558,N_13203,N_13655);
xor U14559 (N_14559,N_13899,N_12120);
nand U14560 (N_14560,N_12082,N_13734);
nand U14561 (N_14561,N_12194,N_13117);
nor U14562 (N_14562,N_12108,N_12280);
nor U14563 (N_14563,N_13497,N_13484);
and U14564 (N_14564,N_12221,N_12019);
xor U14565 (N_14565,N_13428,N_13266);
xor U14566 (N_14566,N_13115,N_12254);
nand U14567 (N_14567,N_13881,N_12015);
and U14568 (N_14568,N_13696,N_13684);
xnor U14569 (N_14569,N_13688,N_12540);
nor U14570 (N_14570,N_13620,N_13144);
nand U14571 (N_14571,N_13652,N_13983);
xor U14572 (N_14572,N_13613,N_12962);
or U14573 (N_14573,N_13839,N_13232);
xnor U14574 (N_14574,N_13851,N_13708);
nor U14575 (N_14575,N_13858,N_12502);
or U14576 (N_14576,N_13187,N_12008);
nand U14577 (N_14577,N_12894,N_13830);
xor U14578 (N_14578,N_13841,N_12760);
or U14579 (N_14579,N_13874,N_13374);
nor U14580 (N_14580,N_13679,N_12453);
nor U14581 (N_14581,N_12595,N_12258);
nand U14582 (N_14582,N_13376,N_13298);
nor U14583 (N_14583,N_12432,N_13512);
nand U14584 (N_14584,N_12247,N_12761);
nor U14585 (N_14585,N_13154,N_13816);
and U14586 (N_14586,N_12482,N_13699);
or U14587 (N_14587,N_12153,N_12711);
xor U14588 (N_14588,N_12716,N_13108);
xnor U14589 (N_14589,N_12048,N_12245);
nor U14590 (N_14590,N_13849,N_12495);
nor U14591 (N_14591,N_12199,N_13335);
nand U14592 (N_14592,N_12242,N_13110);
nand U14593 (N_14593,N_13506,N_12103);
xor U14594 (N_14594,N_12796,N_12454);
xnor U14595 (N_14595,N_12520,N_12590);
nor U14596 (N_14596,N_13284,N_12982);
and U14597 (N_14597,N_12022,N_12834);
and U14598 (N_14598,N_13453,N_12352);
or U14599 (N_14599,N_12825,N_12400);
xor U14600 (N_14600,N_13563,N_13695);
or U14601 (N_14601,N_13582,N_12426);
and U14602 (N_14602,N_13986,N_13610);
or U14603 (N_14603,N_12591,N_13916);
and U14604 (N_14604,N_13581,N_12593);
nor U14605 (N_14605,N_12304,N_13030);
and U14606 (N_14606,N_12372,N_12151);
nor U14607 (N_14607,N_12786,N_13596);
xnor U14608 (N_14608,N_13083,N_13989);
nor U14609 (N_14609,N_12170,N_13938);
nor U14610 (N_14610,N_12463,N_12883);
or U14611 (N_14611,N_13873,N_13603);
nand U14612 (N_14612,N_12650,N_12333);
and U14613 (N_14613,N_13778,N_13257);
xnor U14614 (N_14614,N_12201,N_12662);
and U14615 (N_14615,N_12187,N_12332);
nand U14616 (N_14616,N_13891,N_13617);
nor U14617 (N_14617,N_12574,N_12356);
or U14618 (N_14618,N_12810,N_12955);
and U14619 (N_14619,N_13742,N_12212);
xnor U14620 (N_14620,N_12262,N_12183);
or U14621 (N_14621,N_13014,N_12163);
or U14622 (N_14622,N_12548,N_12550);
and U14623 (N_14623,N_13956,N_12198);
xnor U14624 (N_14624,N_13800,N_13507);
nand U14625 (N_14625,N_13754,N_13028);
nand U14626 (N_14626,N_12447,N_13141);
or U14627 (N_14627,N_13206,N_13703);
nand U14628 (N_14628,N_12335,N_12156);
nor U14629 (N_14629,N_12966,N_13104);
and U14630 (N_14630,N_13887,N_12068);
or U14631 (N_14631,N_13256,N_13251);
nand U14632 (N_14632,N_12049,N_12477);
or U14633 (N_14633,N_13918,N_12496);
nor U14634 (N_14634,N_13039,N_12363);
or U14635 (N_14635,N_12413,N_13061);
nor U14636 (N_14636,N_13319,N_13005);
xnor U14637 (N_14637,N_12564,N_12464);
and U14638 (N_14638,N_12012,N_12367);
or U14639 (N_14639,N_12211,N_12034);
nor U14640 (N_14640,N_12438,N_13128);
xnor U14641 (N_14641,N_12185,N_13126);
xnor U14642 (N_14642,N_13168,N_12394);
nand U14643 (N_14643,N_12462,N_13848);
xor U14644 (N_14644,N_13748,N_13188);
and U14645 (N_14645,N_12301,N_13001);
xor U14646 (N_14646,N_13091,N_13422);
nand U14647 (N_14647,N_13702,N_12975);
and U14648 (N_14648,N_13182,N_12345);
nand U14649 (N_14649,N_13944,N_12793);
nor U14650 (N_14650,N_13281,N_13519);
or U14651 (N_14651,N_13821,N_13770);
and U14652 (N_14652,N_12500,N_13012);
nor U14653 (N_14653,N_12308,N_12427);
or U14654 (N_14654,N_13773,N_12811);
and U14655 (N_14655,N_12109,N_13979);
nand U14656 (N_14656,N_13496,N_13471);
and U14657 (N_14657,N_13905,N_13122);
xor U14658 (N_14658,N_12610,N_12373);
nor U14659 (N_14659,N_13032,N_13692);
and U14660 (N_14660,N_13524,N_13491);
nand U14661 (N_14661,N_12785,N_13663);
nand U14662 (N_14662,N_12444,N_13133);
or U14663 (N_14663,N_12110,N_13207);
or U14664 (N_14664,N_13120,N_12010);
or U14665 (N_14665,N_13536,N_13757);
and U14666 (N_14666,N_12800,N_13420);
xnor U14667 (N_14667,N_12788,N_13931);
nand U14668 (N_14668,N_13876,N_12517);
nor U14669 (N_14669,N_12768,N_12314);
xor U14670 (N_14670,N_12580,N_13468);
or U14671 (N_14671,N_12534,N_13007);
nor U14672 (N_14672,N_13211,N_12095);
nor U14673 (N_14673,N_13010,N_13933);
nand U14674 (N_14674,N_12813,N_12611);
or U14675 (N_14675,N_13717,N_12117);
and U14676 (N_14676,N_12122,N_13123);
nand U14677 (N_14677,N_12129,N_12847);
xnor U14678 (N_14678,N_12232,N_13940);
xnor U14679 (N_14679,N_12374,N_13584);
xnor U14680 (N_14680,N_13205,N_13477);
nor U14681 (N_14681,N_13574,N_12096);
and U14682 (N_14682,N_13373,N_12145);
xnor U14683 (N_14683,N_13139,N_12619);
xnor U14684 (N_14684,N_12741,N_13954);
nor U14685 (N_14685,N_12930,N_13767);
and U14686 (N_14686,N_13363,N_12346);
xnor U14687 (N_14687,N_12350,N_13383);
xnor U14688 (N_14688,N_12284,N_12734);
and U14689 (N_14689,N_13622,N_12206);
xnor U14690 (N_14690,N_12248,N_12227);
or U14691 (N_14691,N_12976,N_13384);
nand U14692 (N_14692,N_12313,N_12721);
and U14693 (N_14693,N_13231,N_12586);
and U14694 (N_14694,N_12415,N_13490);
and U14695 (N_14695,N_13535,N_12343);
nand U14696 (N_14696,N_12166,N_12182);
nand U14697 (N_14697,N_12188,N_12965);
or U14698 (N_14698,N_13158,N_13332);
nand U14699 (N_14699,N_13326,N_12759);
nor U14700 (N_14700,N_13176,N_13086);
and U14701 (N_14701,N_13098,N_13306);
and U14702 (N_14702,N_13589,N_13134);
nand U14703 (N_14703,N_12948,N_13665);
and U14704 (N_14704,N_12535,N_12565);
and U14705 (N_14705,N_12638,N_13854);
or U14706 (N_14706,N_12895,N_13344);
nor U14707 (N_14707,N_12260,N_13560);
xnor U14708 (N_14708,N_13190,N_12494);
or U14709 (N_14709,N_13145,N_12797);
nand U14710 (N_14710,N_13016,N_12583);
nand U14711 (N_14711,N_13786,N_12476);
or U14712 (N_14712,N_13019,N_12549);
nor U14713 (N_14713,N_13930,N_12275);
or U14714 (N_14714,N_12562,N_12266);
nand U14715 (N_14715,N_12999,N_13675);
and U14716 (N_14716,N_13382,N_13964);
nand U14717 (N_14717,N_13343,N_12176);
or U14718 (N_14718,N_13258,N_13331);
nor U14719 (N_14719,N_13169,N_12941);
nand U14720 (N_14720,N_13866,N_12538);
and U14721 (N_14721,N_13463,N_13650);
xor U14722 (N_14722,N_13919,N_12857);
and U14723 (N_14723,N_13212,N_12177);
and U14724 (N_14724,N_13568,N_13355);
or U14725 (N_14725,N_12264,N_13791);
and U14726 (N_14726,N_13863,N_12430);
nor U14727 (N_14727,N_12828,N_13923);
and U14728 (N_14728,N_12377,N_12044);
or U14729 (N_14729,N_13985,N_12640);
and U14730 (N_14730,N_12907,N_13209);
xor U14731 (N_14731,N_12594,N_12799);
or U14732 (N_14732,N_13288,N_13980);
and U14733 (N_14733,N_13265,N_13328);
nand U14734 (N_14734,N_12351,N_12559);
nor U14735 (N_14735,N_13988,N_12274);
xnor U14736 (N_14736,N_13379,N_12666);
xnor U14737 (N_14737,N_13085,N_12831);
xor U14738 (N_14738,N_13345,N_12286);
xnor U14739 (N_14739,N_13059,N_13545);
and U14740 (N_14740,N_13365,N_12158);
nor U14741 (N_14741,N_13478,N_12755);
or U14742 (N_14742,N_13749,N_12362);
and U14743 (N_14743,N_13623,N_13236);
nor U14744 (N_14744,N_12294,N_12869);
xor U14745 (N_14745,N_13320,N_12499);
and U14746 (N_14746,N_13228,N_13294);
nor U14747 (N_14747,N_12047,N_13131);
and U14748 (N_14748,N_13913,N_12710);
or U14749 (N_14749,N_12582,N_12235);
or U14750 (N_14750,N_13915,N_12215);
nand U14751 (N_14751,N_12498,N_13179);
nand U14752 (N_14752,N_12062,N_13029);
nand U14753 (N_14753,N_12932,N_13608);
nor U14754 (N_14754,N_12442,N_13162);
or U14755 (N_14755,N_12532,N_12073);
and U14756 (N_14756,N_13227,N_13475);
nor U14757 (N_14757,N_13920,N_13636);
xor U14758 (N_14758,N_13058,N_13914);
and U14759 (N_14759,N_12909,N_12325);
and U14760 (N_14760,N_12769,N_12161);
nand U14761 (N_14761,N_13743,N_12717);
xnor U14762 (N_14762,N_12518,N_12577);
or U14763 (N_14763,N_13602,N_12604);
xnor U14764 (N_14764,N_13132,N_12781);
nor U14765 (N_14765,N_13947,N_12689);
nor U14766 (N_14766,N_13674,N_12006);
nor U14767 (N_14767,N_13454,N_12896);
and U14768 (N_14768,N_12868,N_13628);
nand U14769 (N_14769,N_12664,N_12541);
and U14770 (N_14770,N_12956,N_13953);
xor U14771 (N_14771,N_13649,N_13455);
xor U14772 (N_14772,N_12704,N_12506);
nand U14773 (N_14773,N_13252,N_12383);
nand U14774 (N_14774,N_13280,N_13556);
nand U14775 (N_14775,N_12390,N_12929);
and U14776 (N_14776,N_13245,N_12553);
and U14777 (N_14777,N_13075,N_13627);
xor U14778 (N_14778,N_13903,N_13064);
or U14779 (N_14779,N_12421,N_13712);
xnor U14780 (N_14780,N_12251,N_13875);
and U14781 (N_14781,N_12441,N_13714);
nand U14782 (N_14782,N_12270,N_12910);
nand U14783 (N_14783,N_13074,N_13625);
or U14784 (N_14784,N_13462,N_12746);
nor U14785 (N_14785,N_12354,N_12295);
nor U14786 (N_14786,N_12222,N_12994);
nand U14787 (N_14787,N_13523,N_12056);
xor U14788 (N_14788,N_12824,N_13105);
or U14789 (N_14789,N_13357,N_12744);
xnor U14790 (N_14790,N_12277,N_13842);
nand U14791 (N_14791,N_13968,N_13279);
or U14792 (N_14792,N_13718,N_12409);
nor U14793 (N_14793,N_13341,N_13580);
and U14794 (N_14794,N_12618,N_13370);
and U14795 (N_14795,N_13557,N_12668);
xnor U14796 (N_14796,N_13958,N_12634);
xnor U14797 (N_14797,N_13322,N_13142);
nor U14798 (N_14798,N_13927,N_12401);
and U14799 (N_14799,N_13810,N_13500);
and U14800 (N_14800,N_13417,N_13689);
xor U14801 (N_14801,N_12218,N_12905);
nand U14802 (N_14802,N_13249,N_12081);
and U14803 (N_14803,N_12923,N_12417);
xnor U14804 (N_14804,N_12754,N_13710);
nand U14805 (N_14805,N_13018,N_13526);
nand U14806 (N_14806,N_12263,N_12898);
or U14807 (N_14807,N_13912,N_12684);
nor U14808 (N_14808,N_13146,N_13518);
nand U14809 (N_14809,N_13807,N_12995);
nor U14810 (N_14810,N_13395,N_13885);
nor U14811 (N_14811,N_12750,N_12133);
or U14812 (N_14812,N_12403,N_13448);
nor U14813 (N_14813,N_13514,N_12452);
nand U14814 (N_14814,N_12244,N_13079);
nor U14815 (N_14815,N_12576,N_12725);
xor U14816 (N_14816,N_12279,N_13998);
nand U14817 (N_14817,N_12065,N_13693);
and U14818 (N_14818,N_12933,N_12446);
or U14819 (N_14819,N_13820,N_12846);
nor U14820 (N_14820,N_12378,N_13253);
nand U14821 (N_14821,N_12036,N_12953);
or U14822 (N_14822,N_12305,N_12902);
nand U14823 (N_14823,N_12224,N_12020);
or U14824 (N_14824,N_12471,N_13495);
nand U14825 (N_14825,N_12273,N_12971);
and U14826 (N_14826,N_12196,N_12687);
nand U14827 (N_14827,N_13604,N_12984);
nand U14828 (N_14828,N_13755,N_12190);
and U14829 (N_14829,N_13449,N_13314);
nor U14830 (N_14830,N_13977,N_13629);
xor U14831 (N_14831,N_12990,N_12645);
and U14832 (N_14832,N_12589,N_12989);
or U14833 (N_14833,N_13669,N_13540);
nor U14834 (N_14834,N_12938,N_12765);
and U14835 (N_14835,N_13529,N_12229);
xnor U14836 (N_14836,N_13824,N_12853);
or U14837 (N_14837,N_13716,N_12395);
nor U14838 (N_14838,N_13276,N_13409);
xor U14839 (N_14839,N_12098,N_12782);
xnor U14840 (N_14840,N_12478,N_13283);
xnor U14841 (N_14841,N_13583,N_13951);
xnor U14842 (N_14842,N_13301,N_13566);
nand U14843 (N_14843,N_13764,N_12997);
xnor U14844 (N_14844,N_13274,N_13080);
nand U14845 (N_14845,N_13488,N_12391);
or U14846 (N_14846,N_13397,N_13194);
and U14847 (N_14847,N_13678,N_13224);
xor U14848 (N_14848,N_12259,N_12748);
xor U14849 (N_14849,N_13161,N_13701);
nor U14850 (N_14850,N_13022,N_13525);
nand U14851 (N_14851,N_13720,N_12685);
or U14852 (N_14852,N_13042,N_13054);
or U14853 (N_14853,N_13031,N_13427);
or U14854 (N_14854,N_13111,N_13510);
xor U14855 (N_14855,N_12521,N_13843);
nand U14856 (N_14856,N_13946,N_12624);
xnor U14857 (N_14857,N_12566,N_12053);
or U14858 (N_14858,N_12829,N_13346);
xnor U14859 (N_14859,N_12674,N_12002);
and U14860 (N_14860,N_13538,N_12324);
nor U14861 (N_14861,N_12042,N_13289);
or U14862 (N_14862,N_12947,N_13530);
nand U14863 (N_14863,N_13658,N_12730);
or U14864 (N_14864,N_12818,N_12091);
and U14865 (N_14865,N_13838,N_12843);
xnor U14866 (N_14866,N_12598,N_12339);
or U14867 (N_14867,N_13248,N_13047);
and U14868 (N_14868,N_13681,N_12656);
nand U14869 (N_14869,N_12659,N_13015);
nor U14870 (N_14870,N_13991,N_13216);
xor U14871 (N_14871,N_13616,N_13736);
and U14872 (N_14872,N_12767,N_12282);
nand U14873 (N_14873,N_12216,N_12917);
or U14874 (N_14874,N_12077,N_13860);
or U14875 (N_14875,N_13638,N_12712);
and U14876 (N_14876,N_12801,N_12029);
nand U14877 (N_14877,N_13426,N_12658);
xnor U14878 (N_14878,N_12516,N_13969);
nor U14879 (N_14879,N_12783,N_13739);
and U14880 (N_14880,N_12398,N_13487);
xnor U14881 (N_14881,N_12358,N_13577);
nand U14882 (N_14882,N_13984,N_12004);
nand U14883 (N_14883,N_12316,N_13672);
nand U14884 (N_14884,N_12849,N_12724);
nor U14885 (N_14885,N_13159,N_13469);
and U14886 (N_14886,N_13878,N_13598);
nor U14887 (N_14887,N_13551,N_12766);
xnor U14888 (N_14888,N_12214,N_12657);
nor U14889 (N_14889,N_13071,N_13366);
and U14890 (N_14890,N_12472,N_12288);
nor U14891 (N_14891,N_12856,N_12900);
or U14892 (N_14892,N_13235,N_13214);
and U14893 (N_14893,N_12872,N_13192);
nor U14894 (N_14894,N_13318,N_12597);
nor U14895 (N_14895,N_12961,N_12043);
xnor U14896 (N_14896,N_13186,N_13150);
or U14897 (N_14897,N_13439,N_13429);
nand U14898 (N_14898,N_13368,N_12867);
or U14899 (N_14899,N_13766,N_12743);
nand U14900 (N_14900,N_12456,N_12739);
xnor U14901 (N_14901,N_12603,N_12539);
nor U14902 (N_14902,N_13661,N_12172);
xnor U14903 (N_14903,N_13609,N_12445);
nor U14904 (N_14904,N_13352,N_13089);
and U14905 (N_14905,N_12468,N_12794);
nand U14906 (N_14906,N_12676,N_13125);
nand U14907 (N_14907,N_12873,N_12569);
or U14908 (N_14908,N_13962,N_13597);
nor U14909 (N_14909,N_12697,N_12845);
nand U14910 (N_14910,N_12968,N_12607);
xnor U14911 (N_14911,N_12952,N_13483);
nor U14912 (N_14912,N_13520,N_13892);
nand U14913 (N_14913,N_12757,N_13697);
xnor U14914 (N_14914,N_12486,N_13337);
and U14915 (N_14915,N_13850,N_13025);
xnor U14916 (N_14916,N_12683,N_13445);
nand U14917 (N_14917,N_13087,N_13539);
or U14918 (N_14918,N_12512,N_12139);
or U14919 (N_14919,N_12423,N_12701);
or U14920 (N_14920,N_12881,N_13296);
and U14921 (N_14921,N_12429,N_12327);
nand U14922 (N_14922,N_13543,N_13732);
or U14923 (N_14923,N_12906,N_12184);
nand U14924 (N_14924,N_12223,N_13765);
xnor U14925 (N_14925,N_12018,N_13752);
and U14926 (N_14926,N_12297,N_12571);
or U14927 (N_14927,N_13465,N_13051);
or U14928 (N_14928,N_12063,N_12360);
nor U14929 (N_14929,N_13474,N_13503);
or U14930 (N_14930,N_12424,N_13388);
xnor U14931 (N_14931,N_12239,N_13901);
nor U14932 (N_14932,N_13884,N_12987);
and U14933 (N_14933,N_12479,N_13041);
xor U14934 (N_14934,N_12764,N_12342);
or U14935 (N_14935,N_13504,N_12652);
and U14936 (N_14936,N_13882,N_13994);
nand U14937 (N_14937,N_13090,N_12897);
nand U14938 (N_14938,N_13941,N_13313);
nand U14939 (N_14939,N_12870,N_13745);
xnor U14940 (N_14940,N_12366,N_12386);
and U14941 (N_14941,N_12207,N_12735);
xor U14942 (N_14942,N_12137,N_13939);
nor U14943 (N_14943,N_13443,N_13936);
xnor U14944 (N_14944,N_13799,N_13555);
nor U14945 (N_14945,N_12996,N_13431);
xor U14946 (N_14946,N_12112,N_13612);
xnor U14947 (N_14947,N_12964,N_13924);
and U14948 (N_14948,N_13303,N_13934);
nand U14949 (N_14949,N_12470,N_12364);
xor U14950 (N_14950,N_12637,N_13992);
and U14951 (N_14951,N_12138,N_13759);
and U14952 (N_14952,N_12527,N_12551);
nand U14953 (N_14953,N_13499,N_13547);
or U14954 (N_14954,N_13857,N_13411);
and U14955 (N_14955,N_13480,N_13865);
nand U14956 (N_14956,N_12967,N_13643);
or U14957 (N_14957,N_12862,N_12017);
and U14958 (N_14958,N_13868,N_12714);
and U14959 (N_14959,N_13237,N_13768);
nand U14960 (N_14960,N_13081,N_13459);
xnor U14961 (N_14961,N_12702,N_12379);
nand U14962 (N_14962,N_13651,N_13102);
nor U14963 (N_14963,N_13466,N_13247);
nand U14964 (N_14964,N_12525,N_13381);
nand U14965 (N_14965,N_13803,N_12164);
and U14966 (N_14966,N_12105,N_13553);
and U14967 (N_14967,N_12089,N_13902);
and U14968 (N_14968,N_13973,N_13591);
and U14969 (N_14969,N_13943,N_13482);
or U14970 (N_14970,N_13297,N_13291);
nand U14971 (N_14971,N_13430,N_13494);
and U14972 (N_14972,N_12887,N_12678);
nand U14973 (N_14973,N_12606,N_12672);
and U14974 (N_14974,N_12626,N_12480);
nand U14975 (N_14975,N_13401,N_12007);
and U14976 (N_14976,N_12733,N_13424);
or U14977 (N_14977,N_12457,N_13798);
nor U14978 (N_14978,N_13096,N_13143);
or U14979 (N_14979,N_12293,N_13635);
or U14980 (N_14980,N_12202,N_12209);
and U14981 (N_14981,N_12935,N_13348);
and U14982 (N_14982,N_12134,N_12686);
or U14983 (N_14983,N_12605,N_13932);
nand U14984 (N_14984,N_13872,N_13808);
or U14985 (N_14985,N_13195,N_13797);
or U14986 (N_14986,N_12630,N_12738);
xnor U14987 (N_14987,N_13997,N_13097);
xor U14988 (N_14988,N_12397,N_13970);
and U14989 (N_14989,N_12443,N_12848);
nor U14990 (N_14990,N_12054,N_12466);
nor U14991 (N_14991,N_13846,N_12885);
nand U14992 (N_14992,N_13446,N_13063);
nand U14993 (N_14993,N_13358,N_13321);
and U14994 (N_14994,N_12726,N_13668);
or U14995 (N_14995,N_12691,N_12826);
and U14996 (N_14996,N_12924,N_13634);
and U14997 (N_14997,N_12723,N_13413);
or U14998 (N_14998,N_13579,N_13364);
nor U14999 (N_14999,N_12281,N_12425);
xor U15000 (N_15000,N_12390,N_12605);
or U15001 (N_15001,N_12126,N_12181);
and U15002 (N_15002,N_12510,N_13047);
nand U15003 (N_15003,N_13252,N_13779);
and U15004 (N_15004,N_13540,N_12295);
or U15005 (N_15005,N_13895,N_13153);
and U15006 (N_15006,N_12577,N_13384);
nand U15007 (N_15007,N_12765,N_12550);
or U15008 (N_15008,N_13526,N_12476);
nor U15009 (N_15009,N_13622,N_13464);
or U15010 (N_15010,N_13323,N_13019);
or U15011 (N_15011,N_12651,N_13505);
or U15012 (N_15012,N_12804,N_13436);
and U15013 (N_15013,N_13114,N_13602);
nor U15014 (N_15014,N_13619,N_13448);
or U15015 (N_15015,N_13791,N_13784);
xor U15016 (N_15016,N_12212,N_12783);
nor U15017 (N_15017,N_12863,N_12735);
and U15018 (N_15018,N_13930,N_13872);
and U15019 (N_15019,N_12947,N_12199);
and U15020 (N_15020,N_12812,N_13126);
xnor U15021 (N_15021,N_13619,N_13095);
nor U15022 (N_15022,N_13276,N_13217);
and U15023 (N_15023,N_12380,N_13625);
nor U15024 (N_15024,N_13448,N_13999);
nor U15025 (N_15025,N_12314,N_13832);
xnor U15026 (N_15026,N_13523,N_13268);
xor U15027 (N_15027,N_13588,N_13053);
or U15028 (N_15028,N_13378,N_12694);
nand U15029 (N_15029,N_13538,N_12941);
or U15030 (N_15030,N_12604,N_12542);
or U15031 (N_15031,N_13473,N_12765);
or U15032 (N_15032,N_12813,N_12155);
xor U15033 (N_15033,N_12472,N_13935);
and U15034 (N_15034,N_12068,N_13144);
and U15035 (N_15035,N_13781,N_13898);
nand U15036 (N_15036,N_13752,N_12563);
or U15037 (N_15037,N_12762,N_12091);
and U15038 (N_15038,N_12423,N_13276);
or U15039 (N_15039,N_12649,N_13858);
nand U15040 (N_15040,N_12975,N_13545);
or U15041 (N_15041,N_12877,N_12011);
nand U15042 (N_15042,N_12267,N_12270);
nand U15043 (N_15043,N_13146,N_12443);
nor U15044 (N_15044,N_12076,N_12140);
or U15045 (N_15045,N_13028,N_12524);
nor U15046 (N_15046,N_12725,N_12852);
nor U15047 (N_15047,N_12505,N_13758);
xnor U15048 (N_15048,N_13152,N_13978);
nor U15049 (N_15049,N_13532,N_13800);
and U15050 (N_15050,N_13569,N_12746);
nor U15051 (N_15051,N_12574,N_12454);
or U15052 (N_15052,N_12579,N_13858);
and U15053 (N_15053,N_12185,N_13321);
nor U15054 (N_15054,N_12113,N_12109);
or U15055 (N_15055,N_13582,N_13806);
and U15056 (N_15056,N_12488,N_13147);
and U15057 (N_15057,N_12080,N_13075);
xor U15058 (N_15058,N_13775,N_13022);
nor U15059 (N_15059,N_12092,N_12084);
and U15060 (N_15060,N_13455,N_12175);
and U15061 (N_15061,N_13938,N_12768);
nand U15062 (N_15062,N_13968,N_12549);
and U15063 (N_15063,N_12799,N_12070);
xor U15064 (N_15064,N_12890,N_13301);
nand U15065 (N_15065,N_12239,N_13130);
xnor U15066 (N_15066,N_12818,N_13598);
or U15067 (N_15067,N_13743,N_13937);
nand U15068 (N_15068,N_13904,N_13629);
and U15069 (N_15069,N_13382,N_13074);
and U15070 (N_15070,N_13743,N_13705);
and U15071 (N_15071,N_12090,N_12387);
nand U15072 (N_15072,N_12569,N_13788);
nor U15073 (N_15073,N_13922,N_13323);
nor U15074 (N_15074,N_13239,N_13489);
xor U15075 (N_15075,N_13790,N_12966);
nand U15076 (N_15076,N_13905,N_13225);
and U15077 (N_15077,N_13484,N_13181);
and U15078 (N_15078,N_13044,N_12888);
xor U15079 (N_15079,N_13776,N_12706);
nand U15080 (N_15080,N_12807,N_12113);
xnor U15081 (N_15081,N_12308,N_12285);
nor U15082 (N_15082,N_13830,N_13301);
or U15083 (N_15083,N_13259,N_13310);
nor U15084 (N_15084,N_13107,N_13490);
nand U15085 (N_15085,N_12577,N_13666);
nand U15086 (N_15086,N_12188,N_12993);
nor U15087 (N_15087,N_12467,N_13891);
and U15088 (N_15088,N_13581,N_12474);
xor U15089 (N_15089,N_13348,N_12264);
and U15090 (N_15090,N_12734,N_12178);
or U15091 (N_15091,N_13543,N_12171);
xnor U15092 (N_15092,N_12284,N_13777);
or U15093 (N_15093,N_13236,N_12073);
xnor U15094 (N_15094,N_13528,N_13833);
nor U15095 (N_15095,N_12236,N_12256);
and U15096 (N_15096,N_13394,N_12438);
or U15097 (N_15097,N_13373,N_13123);
and U15098 (N_15098,N_12538,N_12773);
and U15099 (N_15099,N_12053,N_12949);
nand U15100 (N_15100,N_13052,N_13040);
nor U15101 (N_15101,N_12444,N_12887);
nor U15102 (N_15102,N_12820,N_13798);
or U15103 (N_15103,N_12543,N_13827);
and U15104 (N_15104,N_12641,N_12121);
or U15105 (N_15105,N_13563,N_12061);
or U15106 (N_15106,N_13949,N_13530);
and U15107 (N_15107,N_12457,N_12218);
xnor U15108 (N_15108,N_13259,N_12565);
or U15109 (N_15109,N_12697,N_12360);
and U15110 (N_15110,N_12828,N_13725);
xnor U15111 (N_15111,N_12482,N_12377);
and U15112 (N_15112,N_13215,N_13774);
or U15113 (N_15113,N_12110,N_13829);
or U15114 (N_15114,N_12668,N_13537);
nor U15115 (N_15115,N_13466,N_13499);
or U15116 (N_15116,N_13709,N_13625);
xnor U15117 (N_15117,N_13950,N_12651);
and U15118 (N_15118,N_12437,N_12220);
and U15119 (N_15119,N_12055,N_12328);
and U15120 (N_15120,N_12498,N_12263);
and U15121 (N_15121,N_13797,N_13975);
or U15122 (N_15122,N_13775,N_13831);
xor U15123 (N_15123,N_13168,N_13033);
nor U15124 (N_15124,N_12184,N_12413);
or U15125 (N_15125,N_13394,N_13693);
or U15126 (N_15126,N_13439,N_13495);
and U15127 (N_15127,N_13704,N_13190);
or U15128 (N_15128,N_12680,N_13311);
nor U15129 (N_15129,N_12759,N_12925);
and U15130 (N_15130,N_12856,N_12190);
nor U15131 (N_15131,N_12275,N_13634);
nand U15132 (N_15132,N_12026,N_12523);
nand U15133 (N_15133,N_13487,N_13169);
or U15134 (N_15134,N_13295,N_12045);
xnor U15135 (N_15135,N_12815,N_12881);
xnor U15136 (N_15136,N_12417,N_13575);
and U15137 (N_15137,N_12242,N_13734);
or U15138 (N_15138,N_12322,N_13443);
or U15139 (N_15139,N_13643,N_13179);
and U15140 (N_15140,N_13115,N_13361);
or U15141 (N_15141,N_12317,N_13365);
xnor U15142 (N_15142,N_12339,N_12612);
and U15143 (N_15143,N_13146,N_12146);
and U15144 (N_15144,N_13906,N_13135);
or U15145 (N_15145,N_13026,N_12810);
xor U15146 (N_15146,N_12526,N_12772);
nand U15147 (N_15147,N_12133,N_13207);
nor U15148 (N_15148,N_13244,N_12161);
or U15149 (N_15149,N_13546,N_13124);
nand U15150 (N_15150,N_12494,N_13914);
nor U15151 (N_15151,N_13633,N_12905);
or U15152 (N_15152,N_12439,N_12959);
nand U15153 (N_15153,N_13256,N_13778);
xor U15154 (N_15154,N_12080,N_12698);
xnor U15155 (N_15155,N_12635,N_12413);
xor U15156 (N_15156,N_12382,N_13932);
nand U15157 (N_15157,N_13458,N_12242);
or U15158 (N_15158,N_13116,N_13239);
nor U15159 (N_15159,N_13346,N_13567);
nand U15160 (N_15160,N_12196,N_13479);
nor U15161 (N_15161,N_13343,N_13934);
xnor U15162 (N_15162,N_13722,N_13787);
or U15163 (N_15163,N_12886,N_13358);
xor U15164 (N_15164,N_12130,N_13989);
xor U15165 (N_15165,N_13731,N_12237);
nor U15166 (N_15166,N_12377,N_12569);
xnor U15167 (N_15167,N_13099,N_12676);
xnor U15168 (N_15168,N_12814,N_12469);
or U15169 (N_15169,N_12229,N_13297);
xor U15170 (N_15170,N_12199,N_12527);
or U15171 (N_15171,N_13987,N_12082);
and U15172 (N_15172,N_12563,N_13021);
and U15173 (N_15173,N_13438,N_13183);
nand U15174 (N_15174,N_12570,N_12550);
or U15175 (N_15175,N_13517,N_12054);
and U15176 (N_15176,N_13623,N_12540);
xnor U15177 (N_15177,N_12536,N_12188);
xnor U15178 (N_15178,N_13138,N_13254);
nand U15179 (N_15179,N_13341,N_12616);
nor U15180 (N_15180,N_13993,N_13142);
xor U15181 (N_15181,N_13660,N_12513);
nand U15182 (N_15182,N_13964,N_12311);
nand U15183 (N_15183,N_13184,N_13265);
nor U15184 (N_15184,N_13190,N_13032);
xnor U15185 (N_15185,N_13134,N_13711);
nor U15186 (N_15186,N_12389,N_12556);
and U15187 (N_15187,N_13590,N_13120);
nand U15188 (N_15188,N_13484,N_13681);
nand U15189 (N_15189,N_13947,N_13953);
or U15190 (N_15190,N_12138,N_12945);
nand U15191 (N_15191,N_12393,N_13958);
or U15192 (N_15192,N_12419,N_12015);
and U15193 (N_15193,N_12475,N_12916);
and U15194 (N_15194,N_13173,N_12637);
nor U15195 (N_15195,N_13520,N_13248);
or U15196 (N_15196,N_13960,N_12900);
and U15197 (N_15197,N_13122,N_13897);
nor U15198 (N_15198,N_12774,N_12930);
nor U15199 (N_15199,N_12183,N_13101);
nor U15200 (N_15200,N_13952,N_12032);
or U15201 (N_15201,N_12075,N_12404);
xnor U15202 (N_15202,N_13614,N_12811);
xnor U15203 (N_15203,N_12158,N_12718);
and U15204 (N_15204,N_13678,N_13476);
and U15205 (N_15205,N_13411,N_12084);
xnor U15206 (N_15206,N_13550,N_13573);
or U15207 (N_15207,N_12099,N_12248);
xor U15208 (N_15208,N_12640,N_13155);
xor U15209 (N_15209,N_12752,N_13975);
or U15210 (N_15210,N_13972,N_13378);
and U15211 (N_15211,N_12267,N_13980);
nand U15212 (N_15212,N_12919,N_12057);
and U15213 (N_15213,N_12841,N_13011);
or U15214 (N_15214,N_13248,N_13952);
xor U15215 (N_15215,N_13476,N_12857);
nand U15216 (N_15216,N_12272,N_13578);
nor U15217 (N_15217,N_13191,N_13579);
xnor U15218 (N_15218,N_12129,N_12112);
nand U15219 (N_15219,N_13464,N_13327);
nand U15220 (N_15220,N_13995,N_12732);
nor U15221 (N_15221,N_12620,N_12200);
or U15222 (N_15222,N_12388,N_12803);
or U15223 (N_15223,N_12817,N_13090);
or U15224 (N_15224,N_12587,N_13094);
or U15225 (N_15225,N_12193,N_12472);
nand U15226 (N_15226,N_12820,N_13211);
xnor U15227 (N_15227,N_13992,N_12517);
or U15228 (N_15228,N_13613,N_12551);
nand U15229 (N_15229,N_13603,N_12659);
nor U15230 (N_15230,N_12045,N_12440);
xor U15231 (N_15231,N_12925,N_12203);
and U15232 (N_15232,N_13963,N_13298);
nor U15233 (N_15233,N_13591,N_12210);
nor U15234 (N_15234,N_12450,N_12548);
xor U15235 (N_15235,N_13034,N_13099);
nor U15236 (N_15236,N_13842,N_12962);
xor U15237 (N_15237,N_12681,N_12549);
nand U15238 (N_15238,N_13879,N_12120);
nor U15239 (N_15239,N_12831,N_12073);
nor U15240 (N_15240,N_13752,N_12150);
xor U15241 (N_15241,N_12445,N_12717);
or U15242 (N_15242,N_12753,N_13382);
xor U15243 (N_15243,N_13328,N_13847);
or U15244 (N_15244,N_13149,N_13311);
xor U15245 (N_15245,N_13631,N_13138);
and U15246 (N_15246,N_13937,N_13850);
or U15247 (N_15247,N_12682,N_12926);
or U15248 (N_15248,N_13419,N_13908);
xnor U15249 (N_15249,N_12415,N_12405);
nor U15250 (N_15250,N_12503,N_13605);
nand U15251 (N_15251,N_12878,N_12248);
nand U15252 (N_15252,N_13545,N_12645);
xnor U15253 (N_15253,N_13807,N_13327);
and U15254 (N_15254,N_13949,N_12438);
nor U15255 (N_15255,N_12442,N_12914);
nor U15256 (N_15256,N_13845,N_13836);
and U15257 (N_15257,N_12932,N_13839);
or U15258 (N_15258,N_13532,N_13144);
xnor U15259 (N_15259,N_13542,N_13485);
xor U15260 (N_15260,N_13555,N_12425);
nor U15261 (N_15261,N_12983,N_12501);
xor U15262 (N_15262,N_13302,N_13491);
nor U15263 (N_15263,N_12502,N_12921);
nor U15264 (N_15264,N_12148,N_12677);
or U15265 (N_15265,N_12001,N_12432);
nor U15266 (N_15266,N_12223,N_12890);
xnor U15267 (N_15267,N_12416,N_12439);
and U15268 (N_15268,N_12564,N_12103);
xnor U15269 (N_15269,N_13961,N_12925);
nand U15270 (N_15270,N_13583,N_13981);
xnor U15271 (N_15271,N_12702,N_13753);
nor U15272 (N_15272,N_12315,N_12312);
or U15273 (N_15273,N_13490,N_13840);
or U15274 (N_15274,N_12902,N_12592);
and U15275 (N_15275,N_12219,N_12300);
and U15276 (N_15276,N_13423,N_12193);
and U15277 (N_15277,N_12590,N_12533);
and U15278 (N_15278,N_13552,N_12392);
xnor U15279 (N_15279,N_13898,N_12133);
xor U15280 (N_15280,N_12954,N_12464);
nand U15281 (N_15281,N_12362,N_13134);
or U15282 (N_15282,N_12385,N_13255);
xnor U15283 (N_15283,N_12511,N_13234);
nor U15284 (N_15284,N_12499,N_12909);
or U15285 (N_15285,N_12274,N_12082);
nor U15286 (N_15286,N_13506,N_13255);
xnor U15287 (N_15287,N_12409,N_13603);
nor U15288 (N_15288,N_12886,N_12777);
xor U15289 (N_15289,N_12985,N_12118);
and U15290 (N_15290,N_13269,N_13388);
nor U15291 (N_15291,N_12673,N_12209);
and U15292 (N_15292,N_13093,N_13283);
and U15293 (N_15293,N_13841,N_12123);
xor U15294 (N_15294,N_12347,N_13893);
and U15295 (N_15295,N_13049,N_12236);
or U15296 (N_15296,N_13685,N_13724);
nor U15297 (N_15297,N_13088,N_13004);
nor U15298 (N_15298,N_12481,N_13660);
or U15299 (N_15299,N_13276,N_13043);
nor U15300 (N_15300,N_12568,N_12251);
and U15301 (N_15301,N_13694,N_13918);
and U15302 (N_15302,N_13559,N_13339);
or U15303 (N_15303,N_12587,N_12549);
or U15304 (N_15304,N_12246,N_13479);
xnor U15305 (N_15305,N_12064,N_13791);
nand U15306 (N_15306,N_12979,N_13485);
and U15307 (N_15307,N_12830,N_12704);
or U15308 (N_15308,N_12092,N_12994);
nor U15309 (N_15309,N_12607,N_13205);
and U15310 (N_15310,N_12173,N_13153);
and U15311 (N_15311,N_13027,N_12653);
and U15312 (N_15312,N_12256,N_13806);
or U15313 (N_15313,N_12181,N_12447);
and U15314 (N_15314,N_13020,N_12998);
and U15315 (N_15315,N_13373,N_12411);
or U15316 (N_15316,N_13154,N_13952);
nor U15317 (N_15317,N_13741,N_12306);
nor U15318 (N_15318,N_12938,N_12141);
xnor U15319 (N_15319,N_12209,N_12850);
nor U15320 (N_15320,N_12824,N_12312);
xnor U15321 (N_15321,N_12990,N_12960);
nand U15322 (N_15322,N_13315,N_12584);
or U15323 (N_15323,N_13918,N_13019);
and U15324 (N_15324,N_13708,N_13766);
and U15325 (N_15325,N_12093,N_13913);
xnor U15326 (N_15326,N_12762,N_12311);
or U15327 (N_15327,N_12458,N_13382);
and U15328 (N_15328,N_13304,N_12399);
nor U15329 (N_15329,N_12744,N_12082);
nand U15330 (N_15330,N_13782,N_12976);
nor U15331 (N_15331,N_12957,N_13169);
nor U15332 (N_15332,N_12469,N_13875);
or U15333 (N_15333,N_13014,N_12712);
and U15334 (N_15334,N_13470,N_13263);
and U15335 (N_15335,N_13129,N_13221);
or U15336 (N_15336,N_12495,N_13790);
nor U15337 (N_15337,N_12525,N_12489);
nand U15338 (N_15338,N_12546,N_12595);
or U15339 (N_15339,N_12265,N_12219);
and U15340 (N_15340,N_12967,N_13950);
nor U15341 (N_15341,N_13978,N_13168);
or U15342 (N_15342,N_13115,N_12650);
and U15343 (N_15343,N_12135,N_12391);
nand U15344 (N_15344,N_13638,N_12627);
xor U15345 (N_15345,N_13641,N_12339);
and U15346 (N_15346,N_13633,N_13292);
nand U15347 (N_15347,N_12320,N_12847);
nand U15348 (N_15348,N_12337,N_13256);
nor U15349 (N_15349,N_13891,N_13552);
nor U15350 (N_15350,N_13066,N_13624);
or U15351 (N_15351,N_12130,N_13027);
or U15352 (N_15352,N_12158,N_12482);
or U15353 (N_15353,N_13874,N_13090);
nor U15354 (N_15354,N_13504,N_13558);
and U15355 (N_15355,N_13878,N_13731);
and U15356 (N_15356,N_12323,N_13358);
xor U15357 (N_15357,N_13733,N_13734);
xnor U15358 (N_15358,N_12360,N_12677);
nand U15359 (N_15359,N_13381,N_12262);
nor U15360 (N_15360,N_12092,N_13615);
and U15361 (N_15361,N_12162,N_12677);
nand U15362 (N_15362,N_12565,N_12366);
or U15363 (N_15363,N_12361,N_12416);
nor U15364 (N_15364,N_13889,N_12652);
nor U15365 (N_15365,N_12187,N_13722);
nor U15366 (N_15366,N_12110,N_12925);
and U15367 (N_15367,N_13495,N_12074);
xnor U15368 (N_15368,N_12854,N_13495);
and U15369 (N_15369,N_12138,N_12376);
nor U15370 (N_15370,N_13301,N_12520);
nor U15371 (N_15371,N_12396,N_13447);
nor U15372 (N_15372,N_12895,N_13111);
nor U15373 (N_15373,N_12145,N_12845);
and U15374 (N_15374,N_12371,N_12855);
or U15375 (N_15375,N_13407,N_12689);
xor U15376 (N_15376,N_13657,N_12175);
xnor U15377 (N_15377,N_12265,N_13180);
and U15378 (N_15378,N_12935,N_13218);
nor U15379 (N_15379,N_13165,N_12205);
nand U15380 (N_15380,N_13523,N_12502);
nor U15381 (N_15381,N_13308,N_13400);
nand U15382 (N_15382,N_12997,N_13822);
or U15383 (N_15383,N_13168,N_13419);
nor U15384 (N_15384,N_13044,N_13015);
xnor U15385 (N_15385,N_12743,N_12351);
nand U15386 (N_15386,N_12309,N_13859);
and U15387 (N_15387,N_13936,N_12527);
or U15388 (N_15388,N_13120,N_13432);
or U15389 (N_15389,N_12632,N_13551);
and U15390 (N_15390,N_12814,N_13627);
nand U15391 (N_15391,N_13468,N_12770);
or U15392 (N_15392,N_13545,N_13935);
xor U15393 (N_15393,N_13747,N_12879);
nand U15394 (N_15394,N_13442,N_12502);
and U15395 (N_15395,N_12823,N_13692);
xor U15396 (N_15396,N_13272,N_13435);
or U15397 (N_15397,N_13388,N_12031);
or U15398 (N_15398,N_12098,N_13636);
xor U15399 (N_15399,N_12202,N_13668);
nor U15400 (N_15400,N_12313,N_13292);
xnor U15401 (N_15401,N_13654,N_13521);
nand U15402 (N_15402,N_13436,N_13130);
and U15403 (N_15403,N_13552,N_13654);
or U15404 (N_15404,N_12777,N_12696);
or U15405 (N_15405,N_12641,N_12287);
and U15406 (N_15406,N_12688,N_12217);
nor U15407 (N_15407,N_12257,N_13653);
and U15408 (N_15408,N_12531,N_12074);
or U15409 (N_15409,N_12595,N_13494);
or U15410 (N_15410,N_12126,N_12575);
nor U15411 (N_15411,N_13812,N_12539);
nor U15412 (N_15412,N_12965,N_13695);
or U15413 (N_15413,N_12910,N_13442);
and U15414 (N_15414,N_12782,N_13711);
nand U15415 (N_15415,N_12090,N_12533);
or U15416 (N_15416,N_13988,N_12962);
or U15417 (N_15417,N_13963,N_13807);
or U15418 (N_15418,N_12749,N_12985);
or U15419 (N_15419,N_12359,N_13323);
xnor U15420 (N_15420,N_12265,N_13896);
nor U15421 (N_15421,N_13802,N_13797);
or U15422 (N_15422,N_13063,N_12585);
nor U15423 (N_15423,N_13632,N_13113);
nand U15424 (N_15424,N_12016,N_12289);
nor U15425 (N_15425,N_13196,N_13751);
or U15426 (N_15426,N_13471,N_13080);
and U15427 (N_15427,N_13994,N_12096);
xnor U15428 (N_15428,N_13856,N_12914);
or U15429 (N_15429,N_13799,N_12340);
and U15430 (N_15430,N_13259,N_13547);
nand U15431 (N_15431,N_13743,N_13286);
nor U15432 (N_15432,N_12746,N_13135);
and U15433 (N_15433,N_13696,N_12460);
xnor U15434 (N_15434,N_12144,N_12843);
and U15435 (N_15435,N_12225,N_12027);
nand U15436 (N_15436,N_12660,N_12415);
or U15437 (N_15437,N_13693,N_12007);
nand U15438 (N_15438,N_13099,N_13860);
nand U15439 (N_15439,N_12732,N_13597);
nand U15440 (N_15440,N_13744,N_13423);
and U15441 (N_15441,N_13124,N_13578);
or U15442 (N_15442,N_13685,N_13947);
xor U15443 (N_15443,N_12209,N_13699);
and U15444 (N_15444,N_12378,N_13911);
and U15445 (N_15445,N_12262,N_13085);
nor U15446 (N_15446,N_13111,N_12091);
xor U15447 (N_15447,N_13071,N_13622);
nand U15448 (N_15448,N_13502,N_12129);
nand U15449 (N_15449,N_13589,N_13957);
or U15450 (N_15450,N_13538,N_12419);
and U15451 (N_15451,N_12567,N_12928);
and U15452 (N_15452,N_12880,N_12903);
nor U15453 (N_15453,N_12345,N_13036);
nand U15454 (N_15454,N_12118,N_13823);
or U15455 (N_15455,N_12733,N_13915);
or U15456 (N_15456,N_12903,N_13897);
nand U15457 (N_15457,N_12013,N_12608);
or U15458 (N_15458,N_13866,N_13491);
and U15459 (N_15459,N_13132,N_12511);
nor U15460 (N_15460,N_12631,N_12772);
xnor U15461 (N_15461,N_13253,N_12224);
nand U15462 (N_15462,N_13056,N_13085);
and U15463 (N_15463,N_13721,N_12449);
and U15464 (N_15464,N_13980,N_13423);
xor U15465 (N_15465,N_12996,N_13082);
nor U15466 (N_15466,N_13535,N_13414);
nand U15467 (N_15467,N_12850,N_13702);
or U15468 (N_15468,N_12749,N_12048);
and U15469 (N_15469,N_13502,N_13036);
nor U15470 (N_15470,N_12014,N_12716);
nand U15471 (N_15471,N_13513,N_13667);
or U15472 (N_15472,N_12077,N_12503);
nand U15473 (N_15473,N_12101,N_13417);
nand U15474 (N_15474,N_12723,N_13868);
nor U15475 (N_15475,N_13929,N_12652);
nand U15476 (N_15476,N_13649,N_13104);
xor U15477 (N_15477,N_12569,N_13640);
nand U15478 (N_15478,N_13918,N_13935);
or U15479 (N_15479,N_12015,N_13420);
and U15480 (N_15480,N_12492,N_13430);
xnor U15481 (N_15481,N_13753,N_12539);
xnor U15482 (N_15482,N_12827,N_12138);
xor U15483 (N_15483,N_13242,N_12901);
nand U15484 (N_15484,N_13236,N_13570);
and U15485 (N_15485,N_13527,N_13262);
or U15486 (N_15486,N_13258,N_12614);
nor U15487 (N_15487,N_12590,N_12618);
nor U15488 (N_15488,N_13503,N_13747);
or U15489 (N_15489,N_12550,N_13836);
nand U15490 (N_15490,N_13562,N_12285);
nand U15491 (N_15491,N_13976,N_12736);
and U15492 (N_15492,N_13481,N_12097);
or U15493 (N_15493,N_13441,N_12365);
nor U15494 (N_15494,N_12950,N_12591);
xnor U15495 (N_15495,N_13977,N_12541);
and U15496 (N_15496,N_13703,N_12735);
and U15497 (N_15497,N_13651,N_12376);
xnor U15498 (N_15498,N_12944,N_12484);
nand U15499 (N_15499,N_12571,N_12094);
or U15500 (N_15500,N_13569,N_13982);
xnor U15501 (N_15501,N_13694,N_13003);
or U15502 (N_15502,N_12812,N_12490);
and U15503 (N_15503,N_12641,N_12700);
nor U15504 (N_15504,N_12128,N_13432);
xor U15505 (N_15505,N_13399,N_13407);
and U15506 (N_15506,N_13875,N_13993);
or U15507 (N_15507,N_13790,N_13140);
nand U15508 (N_15508,N_12693,N_12109);
and U15509 (N_15509,N_13325,N_13760);
nand U15510 (N_15510,N_12991,N_13143);
nor U15511 (N_15511,N_12395,N_13884);
nand U15512 (N_15512,N_13297,N_12168);
xor U15513 (N_15513,N_12655,N_13910);
nand U15514 (N_15514,N_12542,N_12906);
nor U15515 (N_15515,N_13100,N_13783);
xnor U15516 (N_15516,N_13769,N_13064);
or U15517 (N_15517,N_13729,N_13117);
or U15518 (N_15518,N_13299,N_13000);
and U15519 (N_15519,N_12929,N_12788);
xor U15520 (N_15520,N_13602,N_13528);
and U15521 (N_15521,N_12585,N_12499);
nand U15522 (N_15522,N_12761,N_13854);
xnor U15523 (N_15523,N_12440,N_12724);
nor U15524 (N_15524,N_12030,N_13491);
xnor U15525 (N_15525,N_12214,N_12798);
xnor U15526 (N_15526,N_13675,N_12080);
xor U15527 (N_15527,N_12538,N_13978);
xnor U15528 (N_15528,N_13355,N_12602);
and U15529 (N_15529,N_12748,N_12281);
or U15530 (N_15530,N_12776,N_13669);
nand U15531 (N_15531,N_12545,N_12438);
or U15532 (N_15532,N_12380,N_12962);
or U15533 (N_15533,N_13898,N_12911);
nand U15534 (N_15534,N_12616,N_12089);
nor U15535 (N_15535,N_12226,N_12711);
nand U15536 (N_15536,N_13190,N_13116);
and U15537 (N_15537,N_12060,N_12352);
nand U15538 (N_15538,N_13839,N_12974);
and U15539 (N_15539,N_13632,N_12364);
nand U15540 (N_15540,N_12398,N_13231);
or U15541 (N_15541,N_12055,N_13005);
nand U15542 (N_15542,N_13413,N_13078);
nand U15543 (N_15543,N_13599,N_13097);
nor U15544 (N_15544,N_13706,N_12535);
or U15545 (N_15545,N_12996,N_13773);
or U15546 (N_15546,N_13854,N_12876);
nor U15547 (N_15547,N_13482,N_12877);
and U15548 (N_15548,N_12031,N_12002);
nand U15549 (N_15549,N_13022,N_12389);
or U15550 (N_15550,N_12166,N_12720);
or U15551 (N_15551,N_13634,N_13742);
and U15552 (N_15552,N_13060,N_12920);
nand U15553 (N_15553,N_12387,N_13431);
and U15554 (N_15554,N_13980,N_12409);
nand U15555 (N_15555,N_12511,N_13348);
and U15556 (N_15556,N_12116,N_12275);
and U15557 (N_15557,N_13779,N_13696);
or U15558 (N_15558,N_12534,N_13553);
nand U15559 (N_15559,N_12741,N_13321);
and U15560 (N_15560,N_13765,N_13667);
nor U15561 (N_15561,N_13957,N_12203);
xnor U15562 (N_15562,N_13231,N_12546);
xor U15563 (N_15563,N_13459,N_13315);
nand U15564 (N_15564,N_12125,N_13449);
nand U15565 (N_15565,N_13271,N_13504);
and U15566 (N_15566,N_12567,N_13886);
or U15567 (N_15567,N_13257,N_12088);
nand U15568 (N_15568,N_13127,N_12133);
xor U15569 (N_15569,N_13452,N_12458);
and U15570 (N_15570,N_13121,N_12642);
nand U15571 (N_15571,N_12208,N_12074);
xnor U15572 (N_15572,N_12022,N_13607);
nor U15573 (N_15573,N_12124,N_13888);
nand U15574 (N_15574,N_13481,N_12930);
xnor U15575 (N_15575,N_12289,N_13883);
and U15576 (N_15576,N_13957,N_13515);
or U15577 (N_15577,N_12007,N_13696);
nor U15578 (N_15578,N_12764,N_13466);
nor U15579 (N_15579,N_12728,N_12093);
xor U15580 (N_15580,N_12361,N_12135);
and U15581 (N_15581,N_13048,N_13737);
nand U15582 (N_15582,N_13873,N_12395);
xor U15583 (N_15583,N_13720,N_13145);
or U15584 (N_15584,N_13846,N_12953);
xor U15585 (N_15585,N_12025,N_12540);
xnor U15586 (N_15586,N_12779,N_12240);
or U15587 (N_15587,N_13666,N_13674);
nand U15588 (N_15588,N_13020,N_13159);
or U15589 (N_15589,N_13689,N_12683);
nor U15590 (N_15590,N_13654,N_12983);
xnor U15591 (N_15591,N_12202,N_13176);
nor U15592 (N_15592,N_12724,N_13392);
xnor U15593 (N_15593,N_13257,N_13982);
nor U15594 (N_15594,N_13693,N_12113);
nand U15595 (N_15595,N_12335,N_13759);
nor U15596 (N_15596,N_13388,N_13920);
nand U15597 (N_15597,N_12121,N_12470);
and U15598 (N_15598,N_12475,N_12975);
nand U15599 (N_15599,N_12872,N_12816);
nand U15600 (N_15600,N_12951,N_13251);
nand U15601 (N_15601,N_12135,N_12515);
nor U15602 (N_15602,N_13144,N_13070);
xor U15603 (N_15603,N_13615,N_13043);
nand U15604 (N_15604,N_12232,N_13572);
and U15605 (N_15605,N_13355,N_12258);
nor U15606 (N_15606,N_13266,N_12744);
nor U15607 (N_15607,N_13401,N_13478);
or U15608 (N_15608,N_13120,N_13111);
nor U15609 (N_15609,N_13649,N_12066);
xnor U15610 (N_15610,N_13094,N_13552);
nand U15611 (N_15611,N_13118,N_13980);
xor U15612 (N_15612,N_12185,N_12205);
nor U15613 (N_15613,N_12507,N_13122);
or U15614 (N_15614,N_12281,N_12360);
xor U15615 (N_15615,N_13525,N_13668);
and U15616 (N_15616,N_13043,N_13847);
and U15617 (N_15617,N_12855,N_12909);
or U15618 (N_15618,N_13788,N_13525);
and U15619 (N_15619,N_12422,N_12134);
xor U15620 (N_15620,N_12412,N_13217);
xor U15621 (N_15621,N_13012,N_13582);
nand U15622 (N_15622,N_13206,N_13519);
or U15623 (N_15623,N_13478,N_13684);
xnor U15624 (N_15624,N_12066,N_12555);
nor U15625 (N_15625,N_13687,N_13603);
nor U15626 (N_15626,N_12007,N_12096);
nor U15627 (N_15627,N_12561,N_12800);
xor U15628 (N_15628,N_13649,N_13466);
nand U15629 (N_15629,N_13301,N_12095);
or U15630 (N_15630,N_13953,N_12918);
nor U15631 (N_15631,N_12176,N_13477);
or U15632 (N_15632,N_12889,N_12178);
nor U15633 (N_15633,N_13531,N_12118);
and U15634 (N_15634,N_12241,N_13182);
and U15635 (N_15635,N_12190,N_13989);
xor U15636 (N_15636,N_13268,N_13686);
and U15637 (N_15637,N_13340,N_12542);
and U15638 (N_15638,N_13735,N_13386);
or U15639 (N_15639,N_12182,N_13484);
and U15640 (N_15640,N_13977,N_13987);
xor U15641 (N_15641,N_13909,N_12615);
or U15642 (N_15642,N_12194,N_12531);
or U15643 (N_15643,N_13949,N_13664);
and U15644 (N_15644,N_12684,N_13964);
xor U15645 (N_15645,N_12979,N_13684);
and U15646 (N_15646,N_12404,N_13233);
nand U15647 (N_15647,N_13980,N_12637);
and U15648 (N_15648,N_13483,N_12712);
and U15649 (N_15649,N_13288,N_12412);
or U15650 (N_15650,N_13479,N_12104);
nand U15651 (N_15651,N_13080,N_12897);
xor U15652 (N_15652,N_13074,N_12842);
nor U15653 (N_15653,N_12214,N_13847);
and U15654 (N_15654,N_13814,N_13385);
xnor U15655 (N_15655,N_12366,N_13167);
nand U15656 (N_15656,N_13125,N_13779);
nor U15657 (N_15657,N_13477,N_13533);
and U15658 (N_15658,N_13186,N_12529);
xor U15659 (N_15659,N_12723,N_13294);
or U15660 (N_15660,N_12386,N_12371);
xnor U15661 (N_15661,N_12070,N_13584);
xor U15662 (N_15662,N_12276,N_13221);
xnor U15663 (N_15663,N_13777,N_12856);
and U15664 (N_15664,N_12231,N_13759);
nand U15665 (N_15665,N_12465,N_12906);
and U15666 (N_15666,N_12487,N_12524);
xnor U15667 (N_15667,N_12364,N_13193);
and U15668 (N_15668,N_12132,N_13677);
nor U15669 (N_15669,N_12687,N_12662);
nand U15670 (N_15670,N_13848,N_12398);
or U15671 (N_15671,N_12824,N_13947);
nand U15672 (N_15672,N_12772,N_13024);
and U15673 (N_15673,N_13190,N_12477);
xnor U15674 (N_15674,N_12076,N_12784);
or U15675 (N_15675,N_12882,N_13738);
nor U15676 (N_15676,N_13379,N_12401);
nand U15677 (N_15677,N_12148,N_12040);
nor U15678 (N_15678,N_13795,N_12676);
or U15679 (N_15679,N_12414,N_12128);
and U15680 (N_15680,N_12992,N_13879);
and U15681 (N_15681,N_12577,N_13794);
or U15682 (N_15682,N_13254,N_13774);
nor U15683 (N_15683,N_12715,N_12409);
xnor U15684 (N_15684,N_13412,N_13503);
and U15685 (N_15685,N_12348,N_13964);
nand U15686 (N_15686,N_12175,N_12273);
nor U15687 (N_15687,N_13651,N_12919);
and U15688 (N_15688,N_12464,N_13542);
nand U15689 (N_15689,N_12354,N_13297);
nand U15690 (N_15690,N_12863,N_13410);
xor U15691 (N_15691,N_12062,N_13252);
nand U15692 (N_15692,N_12232,N_13936);
or U15693 (N_15693,N_13247,N_12060);
xnor U15694 (N_15694,N_13562,N_13064);
and U15695 (N_15695,N_12422,N_13467);
and U15696 (N_15696,N_13586,N_13475);
or U15697 (N_15697,N_13218,N_13398);
or U15698 (N_15698,N_13142,N_13850);
xor U15699 (N_15699,N_13791,N_13887);
or U15700 (N_15700,N_12663,N_12961);
and U15701 (N_15701,N_13091,N_13566);
or U15702 (N_15702,N_12600,N_13111);
xor U15703 (N_15703,N_12477,N_13383);
nor U15704 (N_15704,N_13295,N_13606);
or U15705 (N_15705,N_12181,N_13296);
or U15706 (N_15706,N_12205,N_12310);
and U15707 (N_15707,N_12371,N_13061);
xnor U15708 (N_15708,N_12474,N_13736);
xor U15709 (N_15709,N_13370,N_13204);
nand U15710 (N_15710,N_13824,N_13910);
nand U15711 (N_15711,N_13114,N_13006);
nand U15712 (N_15712,N_13717,N_13425);
nor U15713 (N_15713,N_13095,N_12985);
nand U15714 (N_15714,N_12132,N_13877);
or U15715 (N_15715,N_12257,N_13230);
xor U15716 (N_15716,N_13363,N_13881);
xnor U15717 (N_15717,N_12157,N_12852);
nor U15718 (N_15718,N_12809,N_12775);
nand U15719 (N_15719,N_13201,N_12258);
xor U15720 (N_15720,N_12072,N_13263);
nand U15721 (N_15721,N_13298,N_12729);
and U15722 (N_15722,N_12471,N_12428);
nand U15723 (N_15723,N_12663,N_13267);
or U15724 (N_15724,N_13473,N_12619);
nand U15725 (N_15725,N_12630,N_12890);
and U15726 (N_15726,N_12334,N_13269);
xor U15727 (N_15727,N_13280,N_13323);
nor U15728 (N_15728,N_12605,N_12481);
nand U15729 (N_15729,N_13268,N_12959);
xnor U15730 (N_15730,N_13716,N_12771);
xnor U15731 (N_15731,N_13982,N_13801);
xor U15732 (N_15732,N_12110,N_12011);
and U15733 (N_15733,N_12038,N_13820);
and U15734 (N_15734,N_13292,N_12870);
nand U15735 (N_15735,N_13535,N_13123);
xor U15736 (N_15736,N_12146,N_12799);
nand U15737 (N_15737,N_12213,N_13536);
nand U15738 (N_15738,N_13236,N_12989);
or U15739 (N_15739,N_13548,N_12301);
nand U15740 (N_15740,N_13920,N_12651);
or U15741 (N_15741,N_13673,N_13241);
nand U15742 (N_15742,N_12586,N_13324);
nor U15743 (N_15743,N_13930,N_12853);
or U15744 (N_15744,N_12466,N_12201);
or U15745 (N_15745,N_12670,N_13035);
xor U15746 (N_15746,N_13766,N_13347);
nor U15747 (N_15747,N_12000,N_12559);
and U15748 (N_15748,N_12947,N_13371);
nand U15749 (N_15749,N_13089,N_12733);
or U15750 (N_15750,N_12285,N_12340);
or U15751 (N_15751,N_12267,N_13666);
or U15752 (N_15752,N_12264,N_12027);
nor U15753 (N_15753,N_13535,N_12720);
and U15754 (N_15754,N_12437,N_13342);
and U15755 (N_15755,N_13942,N_12281);
nand U15756 (N_15756,N_12374,N_13081);
xor U15757 (N_15757,N_13338,N_13252);
nand U15758 (N_15758,N_13973,N_12765);
and U15759 (N_15759,N_12646,N_13512);
and U15760 (N_15760,N_13563,N_12899);
or U15761 (N_15761,N_12460,N_12296);
nand U15762 (N_15762,N_13818,N_12883);
nor U15763 (N_15763,N_13723,N_12932);
and U15764 (N_15764,N_12215,N_12560);
and U15765 (N_15765,N_13638,N_12512);
xnor U15766 (N_15766,N_13359,N_13197);
xnor U15767 (N_15767,N_13359,N_12659);
nor U15768 (N_15768,N_12033,N_12719);
nor U15769 (N_15769,N_13997,N_13022);
or U15770 (N_15770,N_13582,N_13973);
xnor U15771 (N_15771,N_12681,N_12618);
nand U15772 (N_15772,N_13709,N_12677);
or U15773 (N_15773,N_13205,N_13618);
or U15774 (N_15774,N_12374,N_12044);
nor U15775 (N_15775,N_13231,N_13555);
xnor U15776 (N_15776,N_13353,N_13664);
nand U15777 (N_15777,N_12201,N_12050);
nor U15778 (N_15778,N_12449,N_12777);
xnor U15779 (N_15779,N_13516,N_12233);
and U15780 (N_15780,N_12664,N_13161);
nor U15781 (N_15781,N_12342,N_12839);
or U15782 (N_15782,N_12668,N_13905);
xnor U15783 (N_15783,N_12314,N_13418);
nand U15784 (N_15784,N_13917,N_12260);
nor U15785 (N_15785,N_13423,N_13430);
and U15786 (N_15786,N_12365,N_12046);
nor U15787 (N_15787,N_13190,N_13072);
or U15788 (N_15788,N_12489,N_12666);
nand U15789 (N_15789,N_12939,N_12810);
nand U15790 (N_15790,N_13710,N_13943);
and U15791 (N_15791,N_13210,N_12129);
and U15792 (N_15792,N_13272,N_12032);
and U15793 (N_15793,N_13768,N_13367);
and U15794 (N_15794,N_13037,N_13049);
and U15795 (N_15795,N_12659,N_12162);
nor U15796 (N_15796,N_12624,N_13137);
and U15797 (N_15797,N_12541,N_13303);
xor U15798 (N_15798,N_13222,N_12846);
and U15799 (N_15799,N_13520,N_12925);
and U15800 (N_15800,N_13705,N_13247);
nor U15801 (N_15801,N_12631,N_12548);
xor U15802 (N_15802,N_12657,N_12254);
and U15803 (N_15803,N_12962,N_13953);
and U15804 (N_15804,N_12427,N_13799);
or U15805 (N_15805,N_12405,N_12812);
nor U15806 (N_15806,N_13661,N_12118);
nand U15807 (N_15807,N_12260,N_13850);
and U15808 (N_15808,N_12445,N_13031);
or U15809 (N_15809,N_13845,N_12731);
or U15810 (N_15810,N_13774,N_12398);
nand U15811 (N_15811,N_12938,N_13228);
or U15812 (N_15812,N_12567,N_13745);
and U15813 (N_15813,N_12449,N_12710);
and U15814 (N_15814,N_13066,N_12045);
or U15815 (N_15815,N_13070,N_13222);
or U15816 (N_15816,N_13866,N_13074);
and U15817 (N_15817,N_13966,N_13921);
xnor U15818 (N_15818,N_12568,N_13000);
or U15819 (N_15819,N_12010,N_13594);
or U15820 (N_15820,N_13779,N_12915);
and U15821 (N_15821,N_12265,N_13327);
and U15822 (N_15822,N_12006,N_13562);
or U15823 (N_15823,N_13680,N_13050);
and U15824 (N_15824,N_12943,N_12702);
and U15825 (N_15825,N_12465,N_13160);
xor U15826 (N_15826,N_13802,N_13427);
nor U15827 (N_15827,N_12853,N_13539);
and U15828 (N_15828,N_13568,N_13085);
or U15829 (N_15829,N_12891,N_13018);
and U15830 (N_15830,N_12054,N_12349);
or U15831 (N_15831,N_12148,N_12285);
or U15832 (N_15832,N_13801,N_12777);
and U15833 (N_15833,N_12194,N_12817);
or U15834 (N_15834,N_13296,N_12240);
or U15835 (N_15835,N_12060,N_13432);
or U15836 (N_15836,N_12438,N_12433);
xnor U15837 (N_15837,N_13046,N_12385);
or U15838 (N_15838,N_13329,N_12654);
nand U15839 (N_15839,N_12270,N_13198);
and U15840 (N_15840,N_12790,N_12691);
nor U15841 (N_15841,N_12172,N_12641);
or U15842 (N_15842,N_13419,N_12788);
xnor U15843 (N_15843,N_12318,N_12611);
or U15844 (N_15844,N_13915,N_13454);
and U15845 (N_15845,N_12956,N_12998);
nand U15846 (N_15846,N_13418,N_12879);
or U15847 (N_15847,N_13776,N_12868);
or U15848 (N_15848,N_12566,N_12326);
nor U15849 (N_15849,N_13753,N_12642);
nor U15850 (N_15850,N_12712,N_13935);
and U15851 (N_15851,N_13436,N_13084);
or U15852 (N_15852,N_13730,N_13402);
nor U15853 (N_15853,N_12773,N_13768);
nand U15854 (N_15854,N_12382,N_13983);
and U15855 (N_15855,N_12449,N_13526);
nand U15856 (N_15856,N_12913,N_13099);
nand U15857 (N_15857,N_12051,N_13710);
xnor U15858 (N_15858,N_13618,N_12543);
nand U15859 (N_15859,N_13637,N_12596);
nor U15860 (N_15860,N_12536,N_12555);
or U15861 (N_15861,N_13864,N_13526);
xnor U15862 (N_15862,N_13489,N_12897);
nand U15863 (N_15863,N_13119,N_12123);
nor U15864 (N_15864,N_13042,N_12437);
nand U15865 (N_15865,N_12566,N_13840);
and U15866 (N_15866,N_13816,N_12692);
nand U15867 (N_15867,N_12926,N_12024);
nor U15868 (N_15868,N_12498,N_13153);
and U15869 (N_15869,N_12874,N_12482);
or U15870 (N_15870,N_13188,N_12950);
xnor U15871 (N_15871,N_13478,N_12382);
or U15872 (N_15872,N_13621,N_12345);
xnor U15873 (N_15873,N_12003,N_13992);
nor U15874 (N_15874,N_12096,N_12562);
nand U15875 (N_15875,N_13930,N_12012);
or U15876 (N_15876,N_12174,N_13803);
or U15877 (N_15877,N_12172,N_13458);
and U15878 (N_15878,N_12690,N_13704);
nand U15879 (N_15879,N_12638,N_13815);
xnor U15880 (N_15880,N_13370,N_13536);
nand U15881 (N_15881,N_13811,N_13636);
and U15882 (N_15882,N_13611,N_13526);
or U15883 (N_15883,N_13821,N_12998);
nor U15884 (N_15884,N_13171,N_13888);
or U15885 (N_15885,N_12763,N_13020);
and U15886 (N_15886,N_13224,N_13779);
xnor U15887 (N_15887,N_12859,N_13919);
nand U15888 (N_15888,N_12616,N_12794);
nand U15889 (N_15889,N_13390,N_12479);
xor U15890 (N_15890,N_13606,N_13047);
xor U15891 (N_15891,N_13847,N_13496);
xor U15892 (N_15892,N_12910,N_13672);
xor U15893 (N_15893,N_13176,N_12920);
and U15894 (N_15894,N_12170,N_12670);
xnor U15895 (N_15895,N_13635,N_13607);
xor U15896 (N_15896,N_12466,N_12115);
nand U15897 (N_15897,N_13472,N_12298);
nand U15898 (N_15898,N_13710,N_13356);
or U15899 (N_15899,N_12718,N_13439);
xnor U15900 (N_15900,N_13008,N_13543);
xnor U15901 (N_15901,N_13710,N_12264);
and U15902 (N_15902,N_13947,N_12989);
nor U15903 (N_15903,N_13260,N_13560);
xnor U15904 (N_15904,N_12604,N_12349);
nor U15905 (N_15905,N_13375,N_12490);
or U15906 (N_15906,N_12191,N_12461);
nand U15907 (N_15907,N_12941,N_12234);
xor U15908 (N_15908,N_12397,N_13934);
and U15909 (N_15909,N_13077,N_12500);
nand U15910 (N_15910,N_13793,N_12484);
nor U15911 (N_15911,N_13578,N_13860);
and U15912 (N_15912,N_13781,N_13199);
nor U15913 (N_15913,N_13617,N_12389);
xor U15914 (N_15914,N_12672,N_13877);
nor U15915 (N_15915,N_13312,N_12568);
or U15916 (N_15916,N_12144,N_13360);
xor U15917 (N_15917,N_13562,N_12392);
or U15918 (N_15918,N_13742,N_12470);
or U15919 (N_15919,N_13050,N_12288);
and U15920 (N_15920,N_12147,N_12971);
or U15921 (N_15921,N_12567,N_12866);
nor U15922 (N_15922,N_12175,N_12991);
and U15923 (N_15923,N_12441,N_12286);
nand U15924 (N_15924,N_13305,N_13559);
nor U15925 (N_15925,N_13551,N_13456);
nand U15926 (N_15926,N_13211,N_13330);
or U15927 (N_15927,N_12820,N_12610);
or U15928 (N_15928,N_12505,N_12514);
xor U15929 (N_15929,N_13304,N_13971);
nor U15930 (N_15930,N_13785,N_13330);
and U15931 (N_15931,N_13205,N_12297);
nand U15932 (N_15932,N_13584,N_13303);
xor U15933 (N_15933,N_13505,N_13976);
nand U15934 (N_15934,N_13739,N_12830);
xnor U15935 (N_15935,N_13490,N_13536);
xnor U15936 (N_15936,N_13155,N_12778);
and U15937 (N_15937,N_12914,N_13048);
or U15938 (N_15938,N_12947,N_12745);
and U15939 (N_15939,N_12287,N_13617);
xnor U15940 (N_15940,N_12985,N_13002);
and U15941 (N_15941,N_13381,N_13693);
xnor U15942 (N_15942,N_12961,N_13116);
xnor U15943 (N_15943,N_13433,N_12662);
xor U15944 (N_15944,N_12378,N_13570);
nor U15945 (N_15945,N_12403,N_12532);
xor U15946 (N_15946,N_13877,N_12108);
xnor U15947 (N_15947,N_12201,N_13660);
and U15948 (N_15948,N_12947,N_13590);
or U15949 (N_15949,N_13825,N_13149);
or U15950 (N_15950,N_13057,N_13816);
nor U15951 (N_15951,N_13140,N_13123);
xor U15952 (N_15952,N_12701,N_12716);
and U15953 (N_15953,N_13061,N_13085);
or U15954 (N_15954,N_13319,N_12783);
nand U15955 (N_15955,N_13761,N_12915);
nor U15956 (N_15956,N_12257,N_12899);
and U15957 (N_15957,N_12584,N_13232);
or U15958 (N_15958,N_12527,N_13134);
nor U15959 (N_15959,N_13289,N_13761);
nor U15960 (N_15960,N_13728,N_13486);
xnor U15961 (N_15961,N_12628,N_12108);
nor U15962 (N_15962,N_13625,N_13405);
nand U15963 (N_15963,N_13919,N_13392);
or U15964 (N_15964,N_12140,N_12953);
nand U15965 (N_15965,N_12123,N_13370);
nand U15966 (N_15966,N_13038,N_13538);
xor U15967 (N_15967,N_13352,N_12724);
nand U15968 (N_15968,N_12880,N_12186);
nand U15969 (N_15969,N_13123,N_12121);
xor U15970 (N_15970,N_13032,N_12055);
and U15971 (N_15971,N_13915,N_12441);
or U15972 (N_15972,N_13931,N_13722);
and U15973 (N_15973,N_12136,N_12010);
nand U15974 (N_15974,N_12374,N_13909);
nand U15975 (N_15975,N_12091,N_13508);
xor U15976 (N_15976,N_12916,N_12103);
and U15977 (N_15977,N_13988,N_12059);
xor U15978 (N_15978,N_13909,N_12675);
nand U15979 (N_15979,N_12615,N_13013);
nor U15980 (N_15980,N_12653,N_13514);
or U15981 (N_15981,N_12031,N_12378);
xor U15982 (N_15982,N_12661,N_12479);
or U15983 (N_15983,N_12847,N_13749);
nand U15984 (N_15984,N_12787,N_13793);
and U15985 (N_15985,N_12874,N_12672);
or U15986 (N_15986,N_12170,N_12751);
and U15987 (N_15987,N_13010,N_12127);
or U15988 (N_15988,N_12049,N_13880);
or U15989 (N_15989,N_13754,N_12794);
nand U15990 (N_15990,N_12990,N_13974);
xnor U15991 (N_15991,N_12369,N_13288);
nand U15992 (N_15992,N_12913,N_12072);
and U15993 (N_15993,N_12747,N_12065);
or U15994 (N_15994,N_13410,N_13863);
or U15995 (N_15995,N_12096,N_13418);
nand U15996 (N_15996,N_12280,N_13640);
nor U15997 (N_15997,N_13767,N_13635);
xnor U15998 (N_15998,N_13396,N_12461);
or U15999 (N_15999,N_12610,N_13189);
and U16000 (N_16000,N_14867,N_15515);
or U16001 (N_16001,N_14132,N_14432);
nand U16002 (N_16002,N_15086,N_15546);
and U16003 (N_16003,N_15732,N_15933);
or U16004 (N_16004,N_14954,N_14176);
xor U16005 (N_16005,N_15590,N_14767);
and U16006 (N_16006,N_15765,N_15301);
nand U16007 (N_16007,N_14527,N_15180);
nand U16008 (N_16008,N_15893,N_15943);
nand U16009 (N_16009,N_14801,N_15811);
and U16010 (N_16010,N_15840,N_14962);
and U16011 (N_16011,N_14862,N_15179);
xnor U16012 (N_16012,N_15800,N_14378);
nand U16013 (N_16013,N_15278,N_15461);
nor U16014 (N_16014,N_15297,N_15453);
nor U16015 (N_16015,N_15136,N_15206);
nor U16016 (N_16016,N_15166,N_14911);
xnor U16017 (N_16017,N_14001,N_15958);
nand U16018 (N_16018,N_15176,N_14853);
or U16019 (N_16019,N_15776,N_14854);
xor U16020 (N_16020,N_14311,N_14893);
and U16021 (N_16021,N_14879,N_15754);
and U16022 (N_16022,N_14721,N_15409);
xnor U16023 (N_16023,N_15350,N_14929);
or U16024 (N_16024,N_15020,N_14582);
or U16025 (N_16025,N_14430,N_14446);
nand U16026 (N_16026,N_15427,N_14461);
xnor U16027 (N_16027,N_15940,N_14116);
nor U16028 (N_16028,N_14160,N_14612);
xnor U16029 (N_16029,N_14847,N_15869);
nor U16030 (N_16030,N_14591,N_15762);
xor U16031 (N_16031,N_15088,N_15486);
nor U16032 (N_16032,N_14387,N_15612);
or U16033 (N_16033,N_15045,N_14966);
nor U16034 (N_16034,N_15311,N_15859);
xnor U16035 (N_16035,N_15932,N_14683);
xor U16036 (N_16036,N_15817,N_15529);
xor U16037 (N_16037,N_14053,N_14921);
nor U16038 (N_16038,N_14778,N_15906);
nand U16039 (N_16039,N_14687,N_14354);
and U16040 (N_16040,N_15900,N_15568);
xor U16041 (N_16041,N_14498,N_15067);
nand U16042 (N_16042,N_14309,N_15174);
xnor U16043 (N_16043,N_14057,N_14535);
nor U16044 (N_16044,N_15693,N_14769);
or U16045 (N_16045,N_15234,N_15008);
nor U16046 (N_16046,N_15905,N_15489);
xor U16047 (N_16047,N_15471,N_15962);
nor U16048 (N_16048,N_14804,N_14232);
and U16049 (N_16049,N_14197,N_14363);
nand U16050 (N_16050,N_15858,N_14965);
xnor U16051 (N_16051,N_14956,N_15246);
and U16052 (N_16052,N_14062,N_14883);
nand U16053 (N_16053,N_15410,N_15043);
nand U16054 (N_16054,N_14168,N_15785);
xor U16055 (N_16055,N_14194,N_15218);
xnor U16056 (N_16056,N_15458,N_15294);
nor U16057 (N_16057,N_14216,N_14831);
and U16058 (N_16058,N_14188,N_14142);
nand U16059 (N_16059,N_14764,N_14816);
nor U16060 (N_16060,N_14439,N_15359);
and U16061 (N_16061,N_14749,N_15347);
nand U16062 (N_16062,N_15126,N_14551);
xor U16063 (N_16063,N_15065,N_15099);
nand U16064 (N_16064,N_14166,N_14085);
and U16065 (N_16065,N_15185,N_14340);
xor U16066 (N_16066,N_14127,N_15436);
and U16067 (N_16067,N_14915,N_14359);
xor U16068 (N_16068,N_15702,N_15030);
or U16069 (N_16069,N_15193,N_15782);
nor U16070 (N_16070,N_15059,N_14871);
or U16071 (N_16071,N_15672,N_15364);
nand U16072 (N_16072,N_15343,N_15586);
nand U16073 (N_16073,N_14468,N_14788);
nand U16074 (N_16074,N_15739,N_15678);
or U16075 (N_16075,N_15983,N_15325);
nand U16076 (N_16076,N_14914,N_14193);
or U16077 (N_16077,N_14576,N_15526);
and U16078 (N_16078,N_15330,N_15571);
xor U16079 (N_16079,N_14088,N_14652);
nor U16080 (N_16080,N_15087,N_15588);
nand U16081 (N_16081,N_14411,N_14138);
and U16082 (N_16082,N_14528,N_15930);
and U16083 (N_16083,N_15259,N_15315);
nand U16084 (N_16084,N_15505,N_15605);
nor U16085 (N_16085,N_15798,N_14248);
nand U16086 (N_16086,N_14348,N_14290);
xnor U16087 (N_16087,N_14316,N_14592);
nor U16088 (N_16088,N_14351,N_15477);
nand U16089 (N_16089,N_15456,N_14492);
xnor U16090 (N_16090,N_15894,N_15549);
xor U16091 (N_16091,N_14964,N_15808);
and U16092 (N_16092,N_15847,N_14648);
nor U16093 (N_16093,N_14917,N_15953);
xnor U16094 (N_16094,N_14018,N_14392);
nand U16095 (N_16095,N_14375,N_15552);
or U16096 (N_16096,N_15873,N_14995);
nor U16097 (N_16097,N_14136,N_15274);
xnor U16098 (N_16098,N_15169,N_15592);
nor U16099 (N_16099,N_15281,N_15215);
xor U16100 (N_16100,N_14066,N_14044);
xnor U16101 (N_16101,N_15133,N_14355);
and U16102 (N_16102,N_14611,N_15837);
or U16103 (N_16103,N_14310,N_14201);
nor U16104 (N_16104,N_14460,N_15767);
or U16105 (N_16105,N_14891,N_14296);
xor U16106 (N_16106,N_15202,N_15826);
nor U16107 (N_16107,N_15466,N_14656);
or U16108 (N_16108,N_14347,N_14990);
nor U16109 (N_16109,N_14986,N_15205);
nor U16110 (N_16110,N_15282,N_14972);
nor U16111 (N_16111,N_14101,N_15679);
nor U16112 (N_16112,N_15334,N_14901);
and U16113 (N_16113,N_15642,N_14613);
nor U16114 (N_16114,N_14462,N_14420);
nand U16115 (N_16115,N_15368,N_14561);
xor U16116 (N_16116,N_15751,N_14164);
or U16117 (N_16117,N_14813,N_14982);
and U16118 (N_16118,N_14930,N_14823);
nor U16119 (N_16119,N_15029,N_15690);
nand U16120 (N_16120,N_15286,N_14448);
nand U16121 (N_16121,N_15665,N_15794);
or U16122 (N_16122,N_14320,N_14558);
xor U16123 (N_16123,N_15077,N_15558);
xor U16124 (N_16124,N_15945,N_14607);
xor U16125 (N_16125,N_15777,N_14293);
or U16126 (N_16126,N_14330,N_14125);
nor U16127 (N_16127,N_14731,N_15769);
nor U16128 (N_16128,N_15952,N_15394);
nand U16129 (N_16129,N_15580,N_15251);
nand U16130 (N_16130,N_15581,N_14413);
and U16131 (N_16131,N_14510,N_14058);
xor U16132 (N_16132,N_14978,N_14619);
or U16133 (N_16133,N_15383,N_14659);
xor U16134 (N_16134,N_15390,N_15531);
nand U16135 (N_16135,N_15539,N_15031);
nand U16136 (N_16136,N_14685,N_15197);
nor U16137 (N_16137,N_14726,N_14999);
or U16138 (N_16138,N_15556,N_14897);
and U16139 (N_16139,N_15071,N_15125);
and U16140 (N_16140,N_14506,N_15670);
and U16141 (N_16141,N_14682,N_14512);
xor U16142 (N_16142,N_15896,N_14442);
nor U16143 (N_16143,N_15803,N_15622);
xnor U16144 (N_16144,N_15727,N_15012);
nand U16145 (N_16145,N_15457,N_14580);
and U16146 (N_16146,N_14383,N_14806);
or U16147 (N_16147,N_14514,N_14428);
nand U16148 (N_16148,N_15663,N_14519);
nor U16149 (N_16149,N_15058,N_15101);
or U16150 (N_16150,N_14975,N_15446);
nand U16151 (N_16151,N_14054,N_15788);
nor U16152 (N_16152,N_14758,N_15113);
xnor U16153 (N_16153,N_15685,N_15599);
xnor U16154 (N_16154,N_15870,N_15435);
nand U16155 (N_16155,N_14111,N_14278);
or U16156 (N_16156,N_14761,N_15097);
nand U16157 (N_16157,N_14313,N_15988);
xnor U16158 (N_16158,N_14333,N_15778);
nand U16159 (N_16159,N_15319,N_15810);
nand U16160 (N_16160,N_15167,N_15979);
and U16161 (N_16161,N_14665,N_14676);
nand U16162 (N_16162,N_15575,N_15011);
and U16163 (N_16163,N_15018,N_14770);
or U16164 (N_16164,N_14186,N_14467);
nor U16165 (N_16165,N_14302,N_15976);
or U16166 (N_16166,N_15266,N_14635);
nor U16167 (N_16167,N_15070,N_15492);
and U16168 (N_16168,N_14908,N_15037);
nand U16169 (N_16169,N_15992,N_14484);
nand U16170 (N_16170,N_14191,N_14239);
xor U16171 (N_16171,N_14745,N_14559);
nor U16172 (N_16172,N_14275,N_15540);
nand U16173 (N_16173,N_14071,N_15152);
nor U16174 (N_16174,N_14546,N_14390);
xor U16175 (N_16175,N_15559,N_14824);
nand U16176 (N_16176,N_15720,N_14729);
nor U16177 (N_16177,N_15861,N_14789);
nor U16178 (N_16178,N_14055,N_14502);
or U16179 (N_16179,N_15696,N_14171);
nand U16180 (N_16180,N_14896,N_15078);
xnor U16181 (N_16181,N_14748,N_14698);
or U16182 (N_16182,N_14977,N_15066);
or U16183 (N_16183,N_14589,N_15824);
and U16184 (N_16184,N_15822,N_14444);
or U16185 (N_16185,N_14950,N_15224);
or U16186 (N_16186,N_14096,N_15151);
and U16187 (N_16187,N_15463,N_15683);
and U16188 (N_16188,N_15853,N_15542);
xnor U16189 (N_16189,N_14543,N_15707);
nor U16190 (N_16190,N_14456,N_14155);
or U16191 (N_16191,N_14765,N_15809);
nand U16192 (N_16192,N_15912,N_15414);
xnor U16193 (N_16193,N_15230,N_15432);
nor U16194 (N_16194,N_15576,N_14918);
or U16195 (N_16195,N_15138,N_15996);
nor U16196 (N_16196,N_15638,N_14518);
nor U16197 (N_16197,N_15632,N_15265);
nor U16198 (N_16198,N_15789,N_15122);
nand U16199 (N_16199,N_14276,N_14606);
xnor U16200 (N_16200,N_14282,N_15922);
xnor U16201 (N_16201,N_15212,N_15271);
xnor U16202 (N_16202,N_14634,N_15474);
nor U16203 (N_16203,N_15135,N_15519);
or U16204 (N_16204,N_14259,N_15594);
or U16205 (N_16205,N_14401,N_14272);
xnor U16206 (N_16206,N_15304,N_14660);
xor U16207 (N_16207,N_14618,N_14567);
and U16208 (N_16208,N_14148,N_15225);
and U16209 (N_16209,N_15154,N_14455);
or U16210 (N_16210,N_15927,N_14107);
or U16211 (N_16211,N_15079,N_15621);
or U16212 (N_16212,N_15960,N_14041);
nand U16213 (N_16213,N_14773,N_15835);
xor U16214 (N_16214,N_14839,N_15157);
nor U16215 (N_16215,N_15986,N_15756);
nand U16216 (N_16216,N_15378,N_14605);
nor U16217 (N_16217,N_14489,N_14089);
or U16218 (N_16218,N_14882,N_14285);
nand U16219 (N_16219,N_15616,N_14126);
and U16220 (N_16220,N_15502,N_14959);
or U16221 (N_16221,N_14860,N_14938);
nand U16222 (N_16222,N_14775,N_15786);
nand U16223 (N_16223,N_15314,N_15994);
nand U16224 (N_16224,N_15273,N_14560);
nor U16225 (N_16225,N_14934,N_15182);
or U16226 (N_16226,N_14905,N_15573);
or U16227 (N_16227,N_15639,N_15236);
xor U16228 (N_16228,N_15761,N_14873);
and U16229 (N_16229,N_14204,N_14403);
and U16230 (N_16230,N_15721,N_15270);
and U16231 (N_16231,N_14398,N_14048);
nor U16232 (N_16232,N_15747,N_14260);
nand U16233 (N_16233,N_14723,N_15421);
nand U16234 (N_16234,N_14991,N_14212);
nor U16235 (N_16235,N_14206,N_15583);
nor U16236 (N_16236,N_15289,N_14124);
and U16237 (N_16237,N_15608,N_14301);
nand U16238 (N_16238,N_15998,N_14158);
and U16239 (N_16239,N_14620,N_15228);
nor U16240 (N_16240,N_14998,N_15134);
or U16241 (N_16241,N_15557,N_15802);
or U16242 (N_16242,N_15454,N_14415);
and U16243 (N_16243,N_15321,N_15082);
or U16244 (N_16244,N_14499,N_15444);
nor U16245 (N_16245,N_15541,N_14324);
or U16246 (N_16246,N_14199,N_14681);
nand U16247 (N_16247,N_14213,N_14440);
xor U16248 (N_16248,N_14488,N_15016);
and U16249 (N_16249,N_14641,N_15668);
nand U16250 (N_16250,N_14261,N_14562);
or U16251 (N_16251,N_15591,N_15401);
and U16252 (N_16252,N_14969,N_15719);
nor U16253 (N_16253,N_15641,N_14690);
nor U16254 (N_16254,N_15513,N_15797);
or U16255 (N_16255,N_14877,N_15628);
and U16256 (N_16256,N_14080,N_14530);
nor U16257 (N_16257,N_14081,N_15833);
nand U16258 (N_16258,N_14757,N_14548);
nand U16259 (N_16259,N_15969,N_15843);
nand U16260 (N_16260,N_14416,N_14183);
xor U16261 (N_16261,N_14247,N_15001);
nor U16262 (N_16262,N_14588,N_14570);
xnor U16263 (N_16263,N_15267,N_15323);
nand U16264 (N_16264,N_15970,N_15300);
nor U16265 (N_16265,N_14856,N_14246);
xor U16266 (N_16266,N_15886,N_15686);
nand U16267 (N_16267,N_14750,N_15563);
nor U16268 (N_16268,N_15380,N_15673);
and U16269 (N_16269,N_15269,N_15340);
nand U16270 (N_16270,N_15164,N_14625);
or U16271 (N_16271,N_14251,N_14815);
nor U16272 (N_16272,N_14190,N_15387);
nand U16273 (N_16273,N_14122,N_15977);
nor U16274 (N_16274,N_15199,N_14574);
nor U16275 (N_16275,N_14350,N_14549);
and U16276 (N_16276,N_14841,N_14357);
nor U16277 (N_16277,N_15033,N_15589);
or U16278 (N_16278,N_14875,N_15650);
xor U16279 (N_16279,N_15815,N_14167);
nor U16280 (N_16280,N_14807,N_14182);
or U16281 (N_16281,N_14257,N_15849);
nand U16282 (N_16282,N_14457,N_14668);
nor U16283 (N_16283,N_14389,N_15714);
and U16284 (N_16284,N_15851,N_15203);
nand U16285 (N_16285,N_14907,N_15255);
and U16286 (N_16286,N_14381,N_14894);
nor U16287 (N_16287,N_14139,N_15377);
and U16288 (N_16288,N_14242,N_15298);
nand U16289 (N_16289,N_14511,N_15419);
nand U16290 (N_16290,N_14289,N_15495);
nand U16291 (N_16291,N_14476,N_15533);
or U16292 (N_16292,N_14798,N_15290);
nor U16293 (N_16293,N_15299,N_15956);
and U16294 (N_16294,N_14819,N_14688);
or U16295 (N_16295,N_15691,N_14590);
xor U16296 (N_16296,N_14103,N_14932);
and U16297 (N_16297,N_14579,N_15076);
nor U16298 (N_16298,N_14105,N_15928);
nand U16299 (N_16299,N_14996,N_15991);
xor U16300 (N_16300,N_15659,N_14377);
and U16301 (N_16301,N_14400,N_14542);
or U16302 (N_16302,N_14827,N_15155);
xor U16303 (N_16303,N_14481,N_14855);
xnor U16304 (N_16304,N_15854,N_15000);
and U16305 (N_16305,N_15990,N_15327);
nor U16306 (N_16306,N_14739,N_15072);
nand U16307 (N_16307,N_14106,N_15468);
and U16308 (N_16308,N_14025,N_14933);
or U16309 (N_16309,N_14624,N_14743);
nor U16310 (N_16310,N_14060,N_15342);
nand U16311 (N_16311,N_14009,N_15884);
nor U16312 (N_16312,N_14077,N_14321);
or U16313 (N_16313,N_14633,N_15832);
and U16314 (N_16314,N_14100,N_15338);
nand U16315 (N_16315,N_15752,N_14727);
nand U16316 (N_16316,N_14779,N_15277);
xor U16317 (N_16317,N_15150,N_14144);
nor U16318 (N_16318,N_15827,N_14870);
or U16319 (N_16319,N_14545,N_15931);
or U16320 (N_16320,N_15115,N_14926);
or U16321 (N_16321,N_15656,N_15060);
xnor U16322 (N_16322,N_14180,N_15369);
xor U16323 (N_16323,N_14864,N_15561);
nor U16324 (N_16324,N_15324,N_14466);
and U16325 (N_16325,N_14479,N_14254);
nand U16326 (N_16326,N_14866,N_15287);
or U16327 (N_16327,N_14751,N_15475);
or U16328 (N_16328,N_14238,N_14117);
or U16329 (N_16329,N_15333,N_14184);
xor U16330 (N_16330,N_14037,N_14046);
or U16331 (N_16331,N_15061,N_14913);
nand U16332 (N_16332,N_14082,N_15820);
and U16333 (N_16333,N_14863,N_15569);
xnor U16334 (N_16334,N_14837,N_15636);
and U16335 (N_16335,N_15521,N_15784);
nor U16336 (N_16336,N_14715,N_15645);
nor U16337 (N_16337,N_15982,N_14300);
nor U16338 (N_16338,N_15613,N_14337);
nor U16339 (N_16339,N_15093,N_15307);
nor U16340 (N_16340,N_15089,N_14507);
xnor U16341 (N_16341,N_15276,N_14920);
or U16342 (N_16342,N_14544,N_14012);
xnor U16343 (N_16343,N_14435,N_14780);
nor U16344 (N_16344,N_14885,N_14419);
or U16345 (N_16345,N_14903,N_14657);
and U16346 (N_16346,N_14332,N_15528);
or U16347 (N_16347,N_15902,N_15339);
and U16348 (N_16348,N_15856,N_15838);
or U16349 (N_16349,N_15503,N_14042);
nor U16350 (N_16350,N_15074,N_15316);
and U16351 (N_16351,N_14280,N_15755);
xor U16352 (N_16352,N_14526,N_15158);
or U16353 (N_16353,N_15288,N_14553);
nor U16354 (N_16354,N_14240,N_14900);
nand U16355 (N_16355,N_14295,N_15178);
xor U16356 (N_16356,N_15211,N_14084);
xnor U16357 (N_16357,N_15795,N_15978);
or U16358 (N_16358,N_15149,N_14335);
or U16359 (N_16359,N_15724,N_15110);
and U16360 (N_16360,N_14137,N_15188);
nor U16361 (N_16361,N_15476,N_15302);
or U16362 (N_16362,N_14341,N_15891);
nor U16363 (N_16363,N_14224,N_15941);
nor U16364 (N_16364,N_15964,N_14755);
and U16365 (N_16365,N_14696,N_15925);
xnor U16366 (N_16366,N_14326,N_15834);
nand U16367 (N_16367,N_14454,N_15127);
nand U16368 (N_16368,N_14671,N_14402);
xor U16369 (N_16369,N_15213,N_14616);
xor U16370 (N_16370,N_15951,N_15601);
and U16371 (N_16371,N_15680,N_15883);
nor U16372 (N_16372,N_15047,N_15508);
and U16373 (N_16373,N_14872,N_14878);
xor U16374 (N_16374,N_14754,N_14369);
nand U16375 (N_16375,N_15014,N_14790);
nor U16376 (N_16376,N_14425,N_15517);
or U16377 (N_16377,N_15470,N_15602);
or U16378 (N_16378,N_14952,N_14365);
and U16379 (N_16379,N_15388,N_14346);
or U16380 (N_16380,N_15625,N_15365);
nand U16381 (N_16381,N_15184,N_15412);
xnor U16382 (N_16382,N_15312,N_15280);
nor U16383 (N_16383,N_14732,N_14145);
nand U16384 (N_16384,N_15813,N_14691);
or U16385 (N_16385,N_14610,N_15918);
nand U16386 (N_16386,N_15313,N_14987);
nor U16387 (N_16387,N_15780,N_15749);
nor U16388 (N_16388,N_14992,N_15416);
xor U16389 (N_16389,N_15177,N_15039);
nor U16390 (N_16390,N_14970,N_14361);
and U16391 (N_16391,N_15864,N_15880);
xnor U16392 (N_16392,N_15748,N_15863);
or U16393 (N_16393,N_15574,N_14079);
and U16394 (N_16394,N_14869,N_14264);
or U16395 (N_16395,N_15562,N_15356);
and U16396 (N_16396,N_15726,N_14857);
xnor U16397 (N_16397,N_15216,N_14904);
and U16398 (N_16398,N_15524,N_14207);
nor U16399 (N_16399,N_15181,N_15128);
nand U16400 (N_16400,N_14976,N_14584);
xnor U16401 (N_16401,N_15091,N_15688);
xor U16402 (N_16402,N_14233,N_15637);
or U16403 (N_16403,N_15243,N_14621);
nor U16404 (N_16404,N_15391,N_15148);
and U16405 (N_16405,N_14159,N_14536);
nand U16406 (N_16406,N_15279,N_15109);
nor U16407 (N_16407,N_15257,N_14636);
and U16408 (N_16408,N_15514,N_15430);
nor U16409 (N_16409,N_15825,N_15868);
nor U16410 (N_16410,N_14304,N_15923);
and U16411 (N_16411,N_15335,N_15386);
and U16412 (N_16412,N_14577,N_14215);
or U16413 (N_16413,N_14477,N_14802);
xor U16414 (N_16414,N_14465,N_15051);
or U16415 (N_16415,N_14703,N_15370);
and U16416 (N_16416,N_15210,N_15015);
nand U16417 (N_16417,N_14019,N_14922);
xor U16418 (N_16418,N_14794,N_15852);
nand U16419 (N_16419,N_15914,N_15735);
nand U16420 (N_16420,N_14931,N_15200);
xnor U16421 (N_16421,N_14781,N_14892);
xor U16422 (N_16422,N_15025,N_15232);
and U16423 (N_16423,N_14287,N_15305);
xor U16424 (N_16424,N_15111,N_14600);
or U16425 (N_16425,N_14031,N_14509);
or U16426 (N_16426,N_14388,N_14662);
and U16427 (N_16427,N_15003,N_15460);
or U16428 (N_16428,N_14719,N_15129);
nand U16429 (N_16429,N_15296,N_15793);
or U16430 (N_16430,N_14021,N_14140);
or U16431 (N_16431,N_14980,N_15063);
xor U16432 (N_16432,N_14017,N_15161);
or U16433 (N_16433,N_15283,N_15219);
nor U16434 (N_16434,N_14850,N_14935);
nor U16435 (N_16435,N_14459,N_14464);
and U16436 (N_16436,N_14851,N_14494);
nor U16437 (N_16437,N_15934,N_14473);
nand U16438 (N_16438,N_14412,N_14424);
and U16439 (N_16439,N_14585,N_15374);
nor U16440 (N_16440,N_14861,N_15473);
nor U16441 (N_16441,N_15395,N_15245);
or U16442 (N_16442,N_15908,N_15306);
nand U16443 (N_16443,N_14814,N_15242);
xnor U16444 (N_16444,N_15183,N_15026);
xor U16445 (N_16445,N_15472,N_14263);
and U16446 (N_16446,N_14886,N_14684);
and U16447 (N_16447,N_14177,N_15879);
nand U16448 (N_16448,N_14472,N_15704);
and U16449 (N_16449,N_14968,N_15587);
nor U16450 (N_16450,N_15814,N_15048);
nor U16451 (N_16451,N_14028,N_14581);
and U16452 (N_16452,N_15450,N_15173);
xnor U16453 (N_16453,N_14485,N_14327);
and U16454 (N_16454,N_14563,N_15949);
xnor U16455 (N_16455,N_14805,N_15346);
nand U16456 (N_16456,N_14989,N_15939);
nand U16457 (N_16457,N_15830,N_14768);
or U16458 (N_16458,N_15360,N_14895);
or U16459 (N_16459,N_15791,N_15146);
or U16460 (N_16460,N_15080,N_15081);
and U16461 (N_16461,N_14586,N_14973);
nand U16462 (N_16462,N_14051,N_15712);
nand U16463 (N_16463,N_14738,N_14228);
and U16464 (N_16464,N_15757,N_14393);
or U16465 (N_16465,N_15980,N_15439);
xnor U16466 (N_16466,N_14937,N_15331);
nor U16467 (N_16467,N_14003,N_15816);
nor U16468 (N_16468,N_14115,N_14035);
or U16469 (N_16469,N_14706,N_15805);
and U16470 (N_16470,N_15938,N_14076);
xor U16471 (N_16471,N_14294,N_15384);
and U16472 (N_16472,N_14078,N_15711);
nand U16473 (N_16473,N_14531,N_14414);
nor U16474 (N_16474,N_15405,N_15536);
and U16475 (N_16475,N_15872,N_14714);
nand U16476 (N_16476,N_14220,N_14550);
xnor U16477 (N_16477,N_14399,N_15829);
nand U16478 (N_16478,N_15090,N_15010);
and U16479 (N_16479,N_14318,N_14385);
and U16480 (N_16480,N_15194,N_14603);
and U16481 (N_16481,N_14705,N_15462);
or U16482 (N_16482,N_14445,N_14523);
nand U16483 (N_16483,N_15411,N_15841);
nand U16484 (N_16484,N_15915,N_15393);
or U16485 (N_16485,N_15677,N_15231);
or U16486 (N_16486,N_15104,N_15046);
xnor U16487 (N_16487,N_15196,N_14249);
nand U16488 (N_16488,N_14376,N_14408);
nor U16489 (N_16489,N_15112,N_14087);
or U16490 (N_16490,N_15885,N_15681);
nor U16491 (N_16491,N_14766,N_14532);
or U16492 (N_16492,N_15709,N_14626);
nor U16493 (N_16493,N_14349,N_15328);
nor U16494 (N_16494,N_14859,N_15911);
nand U16495 (N_16495,N_15443,N_14834);
or U16496 (N_16496,N_15781,N_15248);
nand U16497 (N_16497,N_14284,N_15332);
or U16498 (N_16498,N_15942,N_14840);
or U16499 (N_16499,N_14153,N_14949);
nor U16500 (N_16500,N_14104,N_15839);
nor U16501 (N_16501,N_15131,N_14014);
xor U16502 (N_16502,N_14410,N_15651);
nand U16503 (N_16503,N_15392,N_14899);
and U16504 (N_16504,N_15973,N_15222);
and U16505 (N_16505,N_15653,N_15907);
or U16506 (N_16506,N_14063,N_14373);
xnor U16507 (N_16507,N_14540,N_15376);
nor U16508 (N_16508,N_14593,N_15268);
xor U16509 (N_16509,N_15779,N_15320);
nand U16510 (N_16510,N_14520,N_15828);
and U16511 (N_16511,N_14846,N_15034);
nand U16512 (N_16512,N_15023,N_14267);
and U16513 (N_16513,N_14525,N_14024);
and U16514 (N_16514,N_14130,N_14967);
or U16515 (N_16515,N_14842,N_15867);
or U16516 (N_16516,N_15763,N_15551);
and U16517 (N_16517,N_15362,N_14418);
nand U16518 (N_16518,N_14615,N_14279);
nand U16519 (N_16519,N_14223,N_15351);
and U16520 (N_16520,N_15449,N_15961);
or U16521 (N_16521,N_15165,N_14010);
xnor U16522 (N_16522,N_14067,N_15052);
xnor U16523 (N_16523,N_15195,N_15611);
nor U16524 (N_16524,N_14537,N_15819);
and U16525 (N_16525,N_15692,N_15469);
nor U16526 (N_16526,N_15459,N_14843);
or U16527 (N_16527,N_14308,N_15806);
xnor U16528 (N_16528,N_14214,N_15488);
or U16529 (N_16529,N_15792,N_14747);
or U16530 (N_16530,N_14630,N_14627);
nor U16531 (N_16531,N_14874,N_15094);
nand U16532 (N_16532,N_15487,N_14953);
nor U16533 (N_16533,N_15674,N_15221);
and U16534 (N_16534,N_15027,N_15664);
nor U16535 (N_16535,N_15523,N_14034);
nand U16536 (N_16536,N_14097,N_15959);
and U16537 (N_16537,N_14655,N_15249);
or U16538 (N_16538,N_14849,N_15705);
nor U16539 (N_16539,N_14292,N_14380);
or U16540 (N_16540,N_15028,N_14759);
nand U16541 (N_16541,N_15937,N_15429);
nand U16542 (N_16542,N_15237,N_14368);
or U16543 (N_16543,N_15204,N_15233);
and U16544 (N_16544,N_14491,N_14200);
xnor U16545 (N_16545,N_15096,N_14452);
xnor U16546 (N_16546,N_14269,N_14644);
nand U16547 (N_16547,N_14594,N_14043);
nand U16548 (N_16548,N_15916,N_14713);
and U16549 (N_16549,N_15640,N_14753);
nor U16550 (N_16550,N_14678,N_15038);
nand U16551 (N_16551,N_14198,N_15660);
nand U16552 (N_16552,N_14480,N_14005);
and U16553 (N_16553,N_14945,N_14829);
and U16554 (N_16554,N_14787,N_14784);
nor U16555 (N_16555,N_14833,N_14396);
or U16556 (N_16556,N_15878,N_15263);
nor U16557 (N_16557,N_14640,N_14504);
or U16558 (N_16558,N_14679,N_14651);
xor U16559 (N_16559,N_14673,N_14912);
nor U16560 (N_16560,N_14812,N_15687);
nor U16561 (N_16561,N_14674,N_14564);
or U16562 (N_16562,N_15055,N_15002);
xnor U16563 (N_16563,N_14940,N_14209);
xor U16564 (N_16564,N_15669,N_15371);
and U16565 (N_16565,N_14370,N_14072);
xor U16566 (N_16566,N_15812,N_15550);
nand U16567 (N_16567,N_14822,N_14374);
or U16568 (N_16568,N_15764,N_14203);
and U16569 (N_16569,N_15715,N_15610);
and U16570 (N_16570,N_15217,N_15963);
or U16571 (N_16571,N_15572,N_15141);
xnor U16572 (N_16572,N_15609,N_15142);
nand U16573 (N_16573,N_14360,N_14407);
or U16574 (N_16574,N_14059,N_15506);
or U16575 (N_16575,N_14218,N_14047);
xor U16576 (N_16576,N_14270,N_14487);
nand U16577 (N_16577,N_14538,N_14033);
xor U16578 (N_16578,N_15153,N_15322);
nor U16579 (N_16579,N_14529,N_14925);
or U16580 (N_16580,N_15901,N_14032);
and U16581 (N_16581,N_15666,N_15972);
nand U16582 (N_16582,N_15100,N_14666);
nand U16583 (N_16583,N_15207,N_14686);
nor U16584 (N_16584,N_15760,N_15258);
nand U16585 (N_16585,N_14623,N_14803);
nand U16586 (N_16586,N_15095,N_15262);
or U16587 (N_16587,N_14702,N_14810);
or U16588 (N_16588,N_14181,N_15438);
nor U16589 (N_16589,N_14852,N_15584);
nor U16590 (N_16590,N_14016,N_14150);
nor U16591 (N_16591,N_14098,N_14312);
nand U16592 (N_16592,N_14742,N_14515);
and U16593 (N_16593,N_15718,N_15160);
nand U16594 (N_16594,N_15124,N_15745);
xnor U16595 (N_16595,N_14417,N_14169);
or U16596 (N_16596,N_14948,N_14828);
nand U16597 (N_16597,N_14221,N_14944);
and U16598 (N_16598,N_15498,N_15736);
and U16599 (N_16599,N_15818,N_14910);
and U16600 (N_16600,N_15223,N_14675);
xor U16601 (N_16601,N_15633,N_14314);
and U16602 (N_16602,N_15807,N_15981);
nor U16603 (N_16603,N_14984,N_15684);
nor U16604 (N_16604,N_15848,N_14818);
xnor U16605 (N_16605,N_14008,N_15054);
or U16606 (N_16606,N_15415,N_15787);
and U16607 (N_16607,N_14960,N_15566);
nor U16608 (N_16608,N_14916,N_14273);
xnor U16609 (N_16609,N_14881,N_14353);
nand U16610 (N_16610,N_15921,N_14128);
nor U16611 (N_16611,N_14717,N_14565);
or U16612 (N_16612,N_15534,N_14099);
and U16613 (N_16613,N_14013,N_15192);
or U16614 (N_16614,N_15264,N_15285);
nor U16615 (N_16615,N_15888,N_15750);
and U16616 (N_16616,N_14202,N_14095);
nand U16617 (N_16617,N_14074,N_15860);
nor U16618 (N_16618,N_14250,N_14928);
nand U16619 (N_16619,N_15247,N_14730);
nor U16620 (N_16620,N_14919,N_15984);
or U16621 (N_16621,N_14133,N_14572);
nand U16622 (N_16622,N_15974,N_15578);
or U16623 (N_16623,N_14578,N_14704);
nor U16624 (N_16624,N_15241,N_15518);
nand U16625 (N_16625,N_14252,N_15189);
nor U16626 (N_16626,N_15363,N_14756);
or U16627 (N_16627,N_14746,N_14170);
and U16628 (N_16628,N_14639,N_15701);
xnor U16629 (N_16629,N_15772,N_14596);
and U16630 (N_16630,N_15871,N_15021);
or U16631 (N_16631,N_14146,N_14994);
xnor U16632 (N_16632,N_15897,N_14614);
xor U16633 (N_16633,N_14006,N_15968);
nor U16634 (N_16634,N_15041,N_14352);
or U16635 (N_16635,N_14026,N_15451);
and U16636 (N_16636,N_14174,N_15293);
nand U16637 (N_16637,N_15596,N_14391);
nor U16638 (N_16638,N_15630,N_15455);
nand U16639 (N_16639,N_14771,N_14173);
xor U16640 (N_16640,N_14195,N_15543);
nor U16641 (N_16641,N_14858,N_14236);
and U16642 (N_16642,N_15308,N_15220);
nand U16643 (N_16643,N_15344,N_15117);
or U16644 (N_16644,N_15318,N_15538);
xnor U16645 (N_16645,N_14443,N_14331);
xnor U16646 (N_16646,N_14735,N_14384);
or U16647 (N_16647,N_15053,N_15337);
nor U16648 (N_16648,N_14064,N_15947);
xor U16649 (N_16649,N_14760,N_15032);
xor U16650 (N_16650,N_15865,N_14049);
or U16651 (N_16651,N_15646,N_14604);
and U16652 (N_16652,N_14211,N_14909);
nand U16653 (N_16653,N_15626,N_14923);
or U16654 (N_16654,N_15006,N_15585);
and U16655 (N_16655,N_14587,N_14052);
and U16656 (N_16656,N_14724,N_14149);
or U16657 (N_16657,N_14497,N_15068);
nor U16658 (N_16658,N_14172,N_15671);
xor U16659 (N_16659,N_15103,N_15620);
or U16660 (N_16660,N_15049,N_15105);
and U16661 (N_16661,N_15209,N_14483);
or U16662 (N_16662,N_14073,N_15108);
nor U16663 (N_16663,N_15478,N_15275);
xnor U16664 (N_16664,N_14740,N_14069);
and U16665 (N_16665,N_14880,N_14004);
xnor U16666 (N_16666,N_14832,N_14782);
xor U16667 (N_16667,N_15062,N_14123);
xnor U16668 (N_16668,N_14161,N_14557);
and U16669 (N_16669,N_14000,N_15083);
nand U16670 (N_16670,N_14927,N_15667);
or U16671 (N_16671,N_14256,N_14436);
and U16672 (N_16672,N_15682,N_15846);
and U16673 (N_16673,N_15102,N_14235);
xnor U16674 (N_16674,N_15579,N_15565);
and U16675 (N_16675,N_14939,N_15766);
nand U16676 (N_16676,N_15909,N_15214);
nor U16677 (N_16677,N_14135,N_14573);
xor U16678 (N_16678,N_15437,N_14119);
or U16679 (N_16679,N_14358,N_14608);
xor U16680 (N_16680,N_15892,N_14286);
xor U16681 (N_16681,N_14045,N_14902);
and U16682 (N_16682,N_15967,N_15510);
xnor U16683 (N_16683,N_15137,N_15500);
nor U16684 (N_16684,N_14040,N_15413);
and U16685 (N_16685,N_15433,N_15399);
nor U16686 (N_16686,N_15734,N_15771);
nor U16687 (N_16687,N_14151,N_14291);
and U16688 (N_16688,N_14338,N_14437);
nand U16689 (N_16689,N_14255,N_14065);
and U16690 (N_16690,N_15790,N_15163);
or U16691 (N_16691,N_14664,N_14555);
or U16692 (N_16692,N_14642,N_14029);
xor U16693 (N_16693,N_14471,N_15404);
or U16694 (N_16694,N_14793,N_14208);
and U16695 (N_16695,N_15836,N_15452);
nand U16696 (N_16696,N_15716,N_14441);
or U16697 (N_16697,N_14217,N_15250);
or U16698 (N_16698,N_15208,N_14056);
nor U16699 (N_16699,N_14669,N_15604);
nand U16700 (N_16700,N_14672,N_14786);
and U16701 (N_16701,N_14653,N_14092);
nand U16702 (N_16702,N_15920,N_15995);
or U16703 (N_16703,N_15139,N_15317);
or U16704 (N_16704,N_14617,N_15823);
nand U16705 (N_16705,N_15850,N_15801);
or U16706 (N_16706,N_15567,N_14297);
or U16707 (N_16707,N_15903,N_15198);
nor U16708 (N_16708,N_15501,N_15661);
xnor U16709 (N_16709,N_15844,N_15512);
and U16710 (N_16710,N_15357,N_14595);
xnor U16711 (N_16711,N_14783,N_14241);
and U16712 (N_16712,N_15689,N_15753);
or U16713 (N_16713,N_15698,N_14887);
or U16714 (N_16714,N_15326,N_15485);
or U16715 (N_16715,N_14112,N_15904);
and U16716 (N_16716,N_14482,N_15603);
nor U16717 (N_16717,N_14951,N_15162);
or U16718 (N_16718,N_14234,N_14737);
and U16719 (N_16719,N_14237,N_15845);
nand U16720 (N_16720,N_15073,N_14315);
or U16721 (N_16721,N_15491,N_14889);
xor U16722 (N_16722,N_15227,N_15168);
and U16723 (N_16723,N_15442,N_15773);
xnor U16724 (N_16724,N_14942,N_15582);
nor U16725 (N_16725,N_14156,N_15373);
xor U16726 (N_16726,N_14495,N_15658);
nand U16727 (N_16727,N_14113,N_15635);
nor U16728 (N_16728,N_15950,N_15496);
nand U16729 (N_16729,N_15554,N_15017);
xnor U16730 (N_16730,N_14277,N_14157);
or U16731 (N_16731,N_14710,N_15075);
nand U16732 (N_16732,N_15434,N_15548);
or U16733 (N_16733,N_14838,N_14797);
and U16734 (N_16734,N_15004,N_15783);
nand U16735 (N_16735,N_15560,N_14371);
nand U16736 (N_16736,N_15482,N_14426);
or U16737 (N_16737,N_15121,N_15532);
nand U16738 (N_16738,N_15064,N_15525);
and U16739 (N_16739,N_15403,N_15372);
nor U16740 (N_16740,N_15345,N_15098);
xnor U16741 (N_16741,N_14094,N_15624);
and U16742 (N_16742,N_15627,N_15367);
nand U16743 (N_16743,N_15120,N_15349);
or U16744 (N_16744,N_14697,N_15140);
or U16745 (N_16745,N_15522,N_14429);
or U16746 (N_16746,N_15647,N_15190);
xnor U16747 (N_16747,N_14667,N_15428);
and U16748 (N_16748,N_14453,N_14539);
or U16749 (N_16749,N_14638,N_15957);
xnor U16750 (N_16750,N_15379,N_15527);
nor U16751 (N_16751,N_14187,N_15040);
and U16752 (N_16752,N_14356,N_14274);
and U16753 (N_16753,N_14433,N_15382);
nand U16754 (N_16754,N_15424,N_15309);
nor U16755 (N_16755,N_15971,N_15465);
xnor U16756 (N_16756,N_15744,N_15553);
and U16757 (N_16757,N_15648,N_14533);
and U16758 (N_16758,N_14192,N_14712);
or U16759 (N_16759,N_14936,N_15145);
and U16760 (N_16760,N_14988,N_15713);
xnor U16761 (N_16761,N_14470,N_14458);
nor U16762 (N_16762,N_15240,N_15499);
xor U16763 (N_16763,N_15116,N_15044);
nand U16764 (N_16764,N_14266,N_15186);
nand U16765 (N_16765,N_14205,N_15831);
or U16766 (N_16766,N_15341,N_14646);
and U16767 (N_16767,N_15481,N_14711);
and U16768 (N_16768,N_14825,N_14725);
xnor U16769 (N_16769,N_14118,N_15606);
nand U16770 (N_16770,N_14792,N_15924);
and U16771 (N_16771,N_14830,N_15170);
or U16772 (N_16772,N_14722,N_15728);
nand U16773 (N_16773,N_15544,N_15700);
and U16774 (N_16774,N_15631,N_15036);
or U16775 (N_16775,N_14061,N_15022);
nor U16776 (N_16776,N_14141,N_15402);
nand U16777 (N_16777,N_14162,N_14070);
xnor U16778 (N_16778,N_14961,N_14974);
nor U16779 (N_16779,N_14406,N_15123);
nor U16780 (N_16780,N_15629,N_14486);
xnor U16781 (N_16781,N_15774,N_15857);
nand U16782 (N_16782,N_15643,N_14336);
nand U16783 (N_16783,N_15955,N_15497);
nand U16784 (N_16784,N_14463,N_14299);
nand U16785 (N_16785,N_15397,N_14508);
nand U16786 (N_16786,N_15490,N_15447);
or U16787 (N_16787,N_15598,N_14102);
and U16788 (N_16788,N_15730,N_14253);
or U16789 (N_16789,N_14317,N_15987);
nand U16790 (N_16790,N_15050,N_15600);
or U16791 (N_16791,N_15272,N_15799);
or U16792 (N_16792,N_14307,N_15303);
xor U16793 (N_16793,N_15775,N_14689);
xor U16794 (N_16794,N_14752,N_14776);
or U16795 (N_16795,N_15448,N_15729);
xnor U16796 (N_16796,N_14362,N_14680);
nand U16797 (N_16797,N_14075,N_15398);
or U16798 (N_16798,N_14134,N_14022);
xor U16799 (N_16799,N_14643,N_14645);
and U16800 (N_16800,N_15238,N_15355);
nand U16801 (N_16801,N_15483,N_14556);
or U16802 (N_16802,N_15024,N_14131);
nor U16803 (N_16803,N_15143,N_15975);
xor U16804 (N_16804,N_15440,N_14728);
nor U16805 (N_16805,N_14334,N_14298);
or U16806 (N_16806,N_14015,N_14552);
nor U16807 (N_16807,N_14303,N_14496);
nor U16808 (N_16808,N_14693,N_15917);
or U16809 (N_16809,N_15069,N_14541);
xnor U16810 (N_16810,N_14083,N_15348);
or U16811 (N_16811,N_14774,N_14554);
nor U16812 (N_16812,N_15467,N_15866);
nand U16813 (N_16813,N_14632,N_14971);
or U16814 (N_16814,N_15876,N_14597);
and U16815 (N_16815,N_14245,N_14178);
nor U16816 (N_16816,N_15577,N_14647);
or U16817 (N_16817,N_14888,N_15172);
nand U16818 (N_16818,N_15310,N_14720);
and U16819 (N_16819,N_14475,N_15119);
nand U16820 (N_16820,N_14890,N_14733);
xor U16821 (N_16821,N_14826,N_15898);
xor U16822 (N_16822,N_15644,N_14007);
or U16823 (N_16823,N_15175,N_14800);
and U16824 (N_16824,N_15375,N_15855);
and U16825 (N_16825,N_15889,N_15520);
nor U16826 (N_16826,N_15005,N_14997);
and U16827 (N_16827,N_14328,N_14175);
or U16828 (N_16828,N_14598,N_15910);
nand U16829 (N_16829,N_14744,N_15743);
xnor U16830 (N_16830,N_14050,N_15929);
xor U16831 (N_16831,N_15229,N_15366);
nand U16832 (N_16832,N_14658,N_14981);
or U16833 (N_16833,N_15875,N_14522);
nor U16834 (N_16834,N_14395,N_15420);
and U16835 (N_16835,N_15423,N_14707);
xor U16836 (N_16836,N_15731,N_15738);
xor U16837 (N_16837,N_14367,N_15407);
nor U16838 (N_16838,N_15881,N_15662);
nor U16839 (N_16839,N_14505,N_15329);
xnor U16840 (N_16840,N_15042,N_14898);
nor U16841 (N_16841,N_14086,N_14329);
or U16842 (N_16842,N_14163,N_15422);
nand U16843 (N_16843,N_14709,N_15919);
nand U16844 (N_16844,N_15913,N_15759);
xor U16845 (N_16845,N_15997,N_15895);
xor U16846 (N_16846,N_14517,N_14795);
or U16847 (N_16847,N_14694,N_14093);
xnor U16848 (N_16848,N_14503,N_14583);
and U16849 (N_16849,N_15768,N_15985);
nand U16850 (N_16850,N_14002,N_15400);
nor U16851 (N_16851,N_15593,N_15703);
nor U16852 (N_16852,N_15821,N_14229);
xnor U16853 (N_16853,N_15999,N_14884);
and U16854 (N_16854,N_15899,N_14474);
and U16855 (N_16855,N_14372,N_14397);
or U16856 (N_16856,N_15292,N_15226);
and U16857 (N_16857,N_15295,N_15699);
nor U16858 (N_16858,N_15418,N_15187);
or U16859 (N_16859,N_15597,N_14575);
nor U16860 (N_16860,N_14631,N_14629);
xnor U16861 (N_16861,N_15114,N_15634);
nand U16862 (N_16862,N_15954,N_14121);
or U16863 (N_16863,N_14262,N_15570);
nor U16864 (N_16864,N_15737,N_14421);
and U16865 (N_16865,N_15742,N_14179);
nand U16866 (N_16866,N_14379,N_14993);
xor U16867 (N_16867,N_15619,N_14811);
nor U16868 (N_16868,N_14342,N_14271);
or U16869 (N_16869,N_14152,N_14038);
nor U16870 (N_16870,N_15107,N_15291);
nand U16871 (N_16871,N_15842,N_15352);
and U16872 (N_16872,N_14493,N_14244);
nor U16873 (N_16873,N_15882,N_15710);
or U16874 (N_16874,N_14844,N_14513);
or U16875 (N_16875,N_15717,N_15516);
nand U16876 (N_16876,N_15676,N_14845);
nand U16877 (N_16877,N_14023,N_14670);
or U16878 (N_16878,N_14196,N_14547);
and U16879 (N_16879,N_15935,N_15353);
xor U16880 (N_16880,N_14985,N_15617);
nor U16881 (N_16881,N_14027,N_14692);
or U16882 (N_16882,N_15675,N_15201);
or U16883 (N_16883,N_15989,N_14109);
xor U16884 (N_16884,N_15746,N_14386);
nor U16885 (N_16885,N_14906,N_14030);
nor U16886 (N_16886,N_14020,N_14650);
nand U16887 (N_16887,N_15695,N_14957);
nor U16888 (N_16888,N_15697,N_14677);
and U16889 (N_16889,N_15007,N_14405);
nor U16890 (N_16890,N_14225,N_15804);
xor U16891 (N_16891,N_15965,N_15396);
or U16892 (N_16892,N_15504,N_14501);
xor U16893 (N_16893,N_14868,N_14129);
nand U16894 (N_16894,N_14305,N_15618);
nand U16895 (N_16895,N_15595,N_15657);
and U16896 (N_16896,N_15118,N_15130);
nand U16897 (N_16897,N_15708,N_15741);
and U16898 (N_16898,N_15946,N_14431);
nor U16899 (N_16899,N_14382,N_14323);
or U16900 (N_16900,N_14011,N_14258);
or U16901 (N_16901,N_14404,N_14319);
and U16902 (N_16902,N_15256,N_15555);
nor U16903 (N_16903,N_14409,N_14571);
and U16904 (N_16904,N_15147,N_14422);
and U16905 (N_16905,N_15132,N_14772);
nand U16906 (N_16906,N_14516,N_15085);
and U16907 (N_16907,N_14566,N_15649);
nor U16908 (N_16908,N_14339,N_14451);
nand U16909 (N_16909,N_14039,N_14762);
and U16910 (N_16910,N_14700,N_14345);
nor U16911 (N_16911,N_14343,N_15144);
and U16912 (N_16912,N_15084,N_14654);
and U16913 (N_16913,N_14268,N_14322);
xor U16914 (N_16914,N_14983,N_14243);
xor U16915 (N_16915,N_15009,N_14958);
nand U16916 (N_16916,N_14817,N_15426);
nand U16917 (N_16917,N_14438,N_14568);
nand U16918 (N_16918,N_15926,N_14068);
or U16919 (N_16919,N_15244,N_14701);
and U16920 (N_16920,N_15623,N_14924);
nand U16921 (N_16921,N_15171,N_15253);
and U16922 (N_16922,N_14943,N_15484);
nor U16923 (N_16923,N_15235,N_14091);
xor U16924 (N_16924,N_15694,N_15389);
xnor U16925 (N_16925,N_14478,N_14108);
nand U16926 (N_16926,N_15159,N_14820);
xor U16927 (N_16927,N_14423,N_14699);
and U16928 (N_16928,N_14521,N_15479);
xnor U16929 (N_16929,N_14796,N_14946);
nand U16930 (N_16930,N_15966,N_14785);
nand U16931 (N_16931,N_14306,N_14649);
or U16932 (N_16932,N_14808,N_14821);
or U16933 (N_16933,N_15723,N_15654);
xnor U16934 (N_16934,N_15740,N_14222);
and U16935 (N_16935,N_15261,N_15545);
nor U16936 (N_16936,N_15358,N_15615);
and U16937 (N_16937,N_14364,N_14227);
nor U16938 (N_16938,N_14708,N_14836);
and U16939 (N_16939,N_14344,N_14718);
xor U16940 (N_16940,N_14230,N_14325);
nor U16941 (N_16941,N_15796,N_14791);
or U16942 (N_16942,N_15890,N_14120);
nand U16943 (N_16943,N_14955,N_15417);
nand U16944 (N_16944,N_15381,N_15254);
and U16945 (N_16945,N_15862,N_15239);
nand U16946 (N_16946,N_15252,N_15509);
nand U16947 (N_16947,N_15877,N_15013);
nor U16948 (N_16948,N_14427,N_14143);
nor U16949 (N_16949,N_14449,N_14569);
and U16950 (N_16950,N_15464,N_15408);
or U16951 (N_16951,N_15948,N_14809);
nand U16952 (N_16952,N_15092,N_14663);
or U16953 (N_16953,N_14979,N_14628);
and U16954 (N_16954,N_14450,N_14226);
and U16955 (N_16955,N_15056,N_14524);
nor U16956 (N_16956,N_14876,N_14219);
and U16957 (N_16957,N_14661,N_14490);
nor U16958 (N_16958,N_14154,N_15655);
or U16959 (N_16959,N_14185,N_14941);
xor U16960 (N_16960,N_15057,N_14777);
and U16961 (N_16961,N_14637,N_15480);
xnor U16962 (N_16962,N_15511,N_15993);
nand U16963 (N_16963,N_14394,N_15944);
or U16964 (N_16964,N_15336,N_15564);
xor U16965 (N_16965,N_14599,N_15445);
xor U16966 (N_16966,N_14865,N_14283);
nand U16967 (N_16967,N_14799,N_15758);
nor U16968 (N_16968,N_14695,N_14189);
nor U16969 (N_16969,N_14622,N_14231);
or U16970 (N_16970,N_14210,N_14716);
xnor U16971 (N_16971,N_15035,N_14741);
nand U16972 (N_16972,N_14963,N_15493);
nor U16973 (N_16973,N_15725,N_14763);
xor U16974 (N_16974,N_15361,N_14602);
xnor U16975 (N_16975,N_15874,N_14288);
nand U16976 (N_16976,N_14036,N_14434);
nor U16977 (N_16977,N_15607,N_15530);
nor U16978 (N_16978,N_14147,N_15260);
nand U16979 (N_16979,N_14114,N_15614);
or U16980 (N_16980,N_14534,N_15706);
xor U16981 (N_16981,N_14601,N_15156);
and U16982 (N_16982,N_14110,N_14736);
and U16983 (N_16983,N_15652,N_14848);
and U16984 (N_16984,N_15494,N_15106);
or U16985 (N_16985,N_15936,N_14947);
nor U16986 (N_16986,N_14734,N_14447);
nor U16987 (N_16987,N_15354,N_15770);
and U16988 (N_16988,N_14165,N_15385);
or U16989 (N_16989,N_15547,N_14265);
xnor U16990 (N_16990,N_14835,N_14469);
and U16991 (N_16991,N_14609,N_14500);
nand U16992 (N_16992,N_14090,N_15722);
xnor U16993 (N_16993,N_15406,N_14366);
or U16994 (N_16994,N_15507,N_15191);
nand U16995 (N_16995,N_15431,N_15887);
and U16996 (N_16996,N_15425,N_14281);
and U16997 (N_16997,N_15441,N_15019);
nor U16998 (N_16998,N_15535,N_15284);
xor U16999 (N_16999,N_15733,N_15537);
nor U17000 (N_17000,N_15793,N_14329);
nand U17001 (N_17001,N_14997,N_15617);
nand U17002 (N_17002,N_14974,N_15061);
and U17003 (N_17003,N_14746,N_15503);
and U17004 (N_17004,N_14405,N_14128);
nand U17005 (N_17005,N_15462,N_15833);
and U17006 (N_17006,N_15324,N_15190);
xor U17007 (N_17007,N_15629,N_15244);
nor U17008 (N_17008,N_15233,N_15724);
xnor U17009 (N_17009,N_14638,N_15524);
nand U17010 (N_17010,N_14845,N_14991);
nand U17011 (N_17011,N_15058,N_15900);
and U17012 (N_17012,N_15575,N_14207);
or U17013 (N_17013,N_15723,N_15187);
nor U17014 (N_17014,N_15091,N_14246);
xnor U17015 (N_17015,N_14223,N_14600);
nand U17016 (N_17016,N_15098,N_15034);
xor U17017 (N_17017,N_14800,N_14976);
or U17018 (N_17018,N_14433,N_15158);
nor U17019 (N_17019,N_15052,N_14605);
and U17020 (N_17020,N_15767,N_14995);
or U17021 (N_17021,N_14661,N_15276);
or U17022 (N_17022,N_14233,N_14925);
nor U17023 (N_17023,N_15296,N_14175);
nor U17024 (N_17024,N_14660,N_15956);
xnor U17025 (N_17025,N_15016,N_15571);
nand U17026 (N_17026,N_14831,N_14303);
or U17027 (N_17027,N_15478,N_14510);
nand U17028 (N_17028,N_15235,N_14919);
nor U17029 (N_17029,N_14094,N_15299);
or U17030 (N_17030,N_14909,N_14313);
or U17031 (N_17031,N_15138,N_14631);
nand U17032 (N_17032,N_14815,N_15529);
or U17033 (N_17033,N_14415,N_14298);
nand U17034 (N_17034,N_14525,N_14686);
and U17035 (N_17035,N_14138,N_14141);
and U17036 (N_17036,N_14284,N_14465);
nor U17037 (N_17037,N_15478,N_14712);
and U17038 (N_17038,N_14407,N_14689);
nor U17039 (N_17039,N_14399,N_15160);
or U17040 (N_17040,N_14061,N_15818);
xnor U17041 (N_17041,N_15058,N_14177);
nor U17042 (N_17042,N_14728,N_15712);
nor U17043 (N_17043,N_14048,N_15145);
nand U17044 (N_17044,N_15592,N_15653);
nor U17045 (N_17045,N_15191,N_15416);
and U17046 (N_17046,N_14529,N_14135);
nor U17047 (N_17047,N_14810,N_14600);
or U17048 (N_17048,N_14146,N_14837);
or U17049 (N_17049,N_15281,N_14280);
and U17050 (N_17050,N_15772,N_15700);
nor U17051 (N_17051,N_14888,N_14889);
or U17052 (N_17052,N_15450,N_14634);
and U17053 (N_17053,N_14427,N_15598);
nand U17054 (N_17054,N_14569,N_14319);
or U17055 (N_17055,N_15369,N_14812);
xnor U17056 (N_17056,N_14581,N_14463);
and U17057 (N_17057,N_15309,N_15008);
nand U17058 (N_17058,N_15783,N_15357);
nand U17059 (N_17059,N_15058,N_15392);
nor U17060 (N_17060,N_14419,N_14967);
or U17061 (N_17061,N_14964,N_15860);
nand U17062 (N_17062,N_14428,N_15410);
and U17063 (N_17063,N_14345,N_15053);
nand U17064 (N_17064,N_15841,N_14994);
or U17065 (N_17065,N_14850,N_15445);
or U17066 (N_17066,N_14784,N_14619);
or U17067 (N_17067,N_15047,N_14111);
or U17068 (N_17068,N_14891,N_14965);
nand U17069 (N_17069,N_14253,N_14366);
xor U17070 (N_17070,N_14284,N_14268);
xor U17071 (N_17071,N_14975,N_15749);
nand U17072 (N_17072,N_14019,N_15350);
and U17073 (N_17073,N_15532,N_15079);
or U17074 (N_17074,N_14693,N_14657);
nor U17075 (N_17075,N_15343,N_15130);
and U17076 (N_17076,N_15498,N_14874);
or U17077 (N_17077,N_14974,N_14793);
nand U17078 (N_17078,N_14911,N_14688);
and U17079 (N_17079,N_15004,N_14660);
and U17080 (N_17080,N_15312,N_14535);
xor U17081 (N_17081,N_15531,N_14936);
and U17082 (N_17082,N_15935,N_15905);
nand U17083 (N_17083,N_14448,N_15451);
or U17084 (N_17084,N_14343,N_15447);
or U17085 (N_17085,N_14920,N_14510);
nand U17086 (N_17086,N_14860,N_15035);
nand U17087 (N_17087,N_15113,N_15640);
nand U17088 (N_17088,N_15239,N_14332);
nor U17089 (N_17089,N_14709,N_14158);
nand U17090 (N_17090,N_15859,N_15567);
or U17091 (N_17091,N_15873,N_14363);
or U17092 (N_17092,N_15824,N_14163);
and U17093 (N_17093,N_14301,N_14129);
nor U17094 (N_17094,N_14109,N_15844);
or U17095 (N_17095,N_15204,N_14524);
or U17096 (N_17096,N_14579,N_14909);
nor U17097 (N_17097,N_14577,N_14894);
nor U17098 (N_17098,N_15441,N_15875);
or U17099 (N_17099,N_15062,N_15055);
nor U17100 (N_17100,N_15205,N_15541);
nor U17101 (N_17101,N_14265,N_14655);
nor U17102 (N_17102,N_15269,N_14991);
nand U17103 (N_17103,N_15421,N_15967);
and U17104 (N_17104,N_15071,N_15573);
and U17105 (N_17105,N_15121,N_15488);
nor U17106 (N_17106,N_15793,N_14193);
xor U17107 (N_17107,N_14567,N_15520);
nand U17108 (N_17108,N_14078,N_15239);
nor U17109 (N_17109,N_14324,N_15621);
xnor U17110 (N_17110,N_15392,N_15343);
nand U17111 (N_17111,N_15108,N_14660);
nand U17112 (N_17112,N_14718,N_14004);
or U17113 (N_17113,N_14696,N_15167);
nor U17114 (N_17114,N_15008,N_14982);
nor U17115 (N_17115,N_14965,N_15078);
xor U17116 (N_17116,N_15751,N_14550);
nor U17117 (N_17117,N_15041,N_15244);
and U17118 (N_17118,N_14144,N_14375);
nand U17119 (N_17119,N_14629,N_14839);
or U17120 (N_17120,N_15304,N_15000);
xnor U17121 (N_17121,N_14006,N_14585);
or U17122 (N_17122,N_14068,N_15688);
or U17123 (N_17123,N_15193,N_14713);
nand U17124 (N_17124,N_14133,N_14829);
nand U17125 (N_17125,N_15250,N_15939);
nand U17126 (N_17126,N_15526,N_14249);
nor U17127 (N_17127,N_14372,N_15631);
and U17128 (N_17128,N_15042,N_14401);
xnor U17129 (N_17129,N_14687,N_15838);
nand U17130 (N_17130,N_15454,N_14712);
and U17131 (N_17131,N_15199,N_14158);
nand U17132 (N_17132,N_15436,N_14485);
xor U17133 (N_17133,N_15542,N_14219);
and U17134 (N_17134,N_15769,N_14234);
or U17135 (N_17135,N_15780,N_14065);
nand U17136 (N_17136,N_15369,N_14890);
xnor U17137 (N_17137,N_15858,N_14629);
or U17138 (N_17138,N_15698,N_15497);
xnor U17139 (N_17139,N_14498,N_14260);
nand U17140 (N_17140,N_15395,N_15690);
nand U17141 (N_17141,N_14946,N_15617);
nand U17142 (N_17142,N_15892,N_14345);
nor U17143 (N_17143,N_15888,N_14224);
xnor U17144 (N_17144,N_14455,N_15679);
nor U17145 (N_17145,N_14998,N_14179);
xnor U17146 (N_17146,N_15742,N_15691);
and U17147 (N_17147,N_14170,N_15524);
nor U17148 (N_17148,N_14661,N_15182);
xnor U17149 (N_17149,N_14683,N_14731);
or U17150 (N_17150,N_15525,N_14365);
nor U17151 (N_17151,N_15061,N_15602);
xor U17152 (N_17152,N_14729,N_14710);
xnor U17153 (N_17153,N_14056,N_14209);
and U17154 (N_17154,N_15693,N_14410);
nor U17155 (N_17155,N_14946,N_14479);
nand U17156 (N_17156,N_15159,N_14888);
nor U17157 (N_17157,N_15882,N_15948);
xor U17158 (N_17158,N_14332,N_14772);
xnor U17159 (N_17159,N_15214,N_15314);
nor U17160 (N_17160,N_14132,N_14104);
nand U17161 (N_17161,N_14831,N_15346);
nand U17162 (N_17162,N_15960,N_14346);
nand U17163 (N_17163,N_14726,N_15417);
xor U17164 (N_17164,N_15099,N_14529);
nor U17165 (N_17165,N_15496,N_14265);
and U17166 (N_17166,N_15378,N_15295);
xnor U17167 (N_17167,N_14366,N_15892);
and U17168 (N_17168,N_14381,N_14339);
xor U17169 (N_17169,N_15829,N_14548);
nand U17170 (N_17170,N_15423,N_14206);
xnor U17171 (N_17171,N_14904,N_15377);
nor U17172 (N_17172,N_15359,N_14720);
or U17173 (N_17173,N_15987,N_15701);
xnor U17174 (N_17174,N_14221,N_15509);
nand U17175 (N_17175,N_14878,N_15007);
xor U17176 (N_17176,N_14879,N_15465);
or U17177 (N_17177,N_15639,N_14379);
and U17178 (N_17178,N_14095,N_15984);
xnor U17179 (N_17179,N_14256,N_15850);
nand U17180 (N_17180,N_15272,N_15132);
and U17181 (N_17181,N_15630,N_14312);
or U17182 (N_17182,N_15931,N_14418);
and U17183 (N_17183,N_15515,N_14858);
nand U17184 (N_17184,N_14486,N_15612);
or U17185 (N_17185,N_14506,N_15231);
nor U17186 (N_17186,N_15245,N_15135);
nor U17187 (N_17187,N_14562,N_15097);
or U17188 (N_17188,N_14644,N_15262);
or U17189 (N_17189,N_14846,N_15691);
and U17190 (N_17190,N_14181,N_15653);
and U17191 (N_17191,N_15598,N_15919);
and U17192 (N_17192,N_14100,N_14237);
nor U17193 (N_17193,N_14964,N_14912);
nor U17194 (N_17194,N_15544,N_15048);
nand U17195 (N_17195,N_15052,N_15264);
and U17196 (N_17196,N_14986,N_14946);
nand U17197 (N_17197,N_15824,N_15866);
xnor U17198 (N_17198,N_15501,N_15214);
nor U17199 (N_17199,N_14819,N_15892);
xnor U17200 (N_17200,N_15513,N_15589);
nand U17201 (N_17201,N_15017,N_14360);
and U17202 (N_17202,N_15819,N_15304);
xnor U17203 (N_17203,N_15594,N_15701);
or U17204 (N_17204,N_14882,N_14670);
and U17205 (N_17205,N_15036,N_15890);
or U17206 (N_17206,N_14930,N_15427);
nor U17207 (N_17207,N_15073,N_15112);
nor U17208 (N_17208,N_15591,N_15220);
and U17209 (N_17209,N_15817,N_15763);
nand U17210 (N_17210,N_14013,N_15990);
nor U17211 (N_17211,N_15009,N_14684);
or U17212 (N_17212,N_15375,N_15195);
nand U17213 (N_17213,N_14579,N_14199);
xor U17214 (N_17214,N_15441,N_14127);
or U17215 (N_17215,N_15158,N_15442);
xnor U17216 (N_17216,N_15023,N_14929);
and U17217 (N_17217,N_15637,N_14889);
xnor U17218 (N_17218,N_14006,N_14287);
xnor U17219 (N_17219,N_14347,N_15130);
nor U17220 (N_17220,N_15129,N_14986);
xor U17221 (N_17221,N_15666,N_15805);
and U17222 (N_17222,N_15743,N_15909);
or U17223 (N_17223,N_14121,N_15008);
nand U17224 (N_17224,N_14280,N_14700);
nor U17225 (N_17225,N_15983,N_14954);
nor U17226 (N_17226,N_14753,N_14027);
and U17227 (N_17227,N_15773,N_15696);
nor U17228 (N_17228,N_14125,N_14716);
xor U17229 (N_17229,N_14807,N_15108);
xnor U17230 (N_17230,N_14287,N_15404);
nand U17231 (N_17231,N_15626,N_15181);
and U17232 (N_17232,N_14270,N_14317);
or U17233 (N_17233,N_14336,N_14440);
xor U17234 (N_17234,N_14181,N_15251);
and U17235 (N_17235,N_15317,N_14230);
and U17236 (N_17236,N_14578,N_14347);
xor U17237 (N_17237,N_14504,N_15253);
xnor U17238 (N_17238,N_14062,N_14491);
nor U17239 (N_17239,N_15069,N_15399);
or U17240 (N_17240,N_14152,N_15638);
nor U17241 (N_17241,N_15352,N_14858);
nor U17242 (N_17242,N_14619,N_14137);
xnor U17243 (N_17243,N_14888,N_14817);
and U17244 (N_17244,N_15393,N_15291);
or U17245 (N_17245,N_15764,N_15540);
or U17246 (N_17246,N_14086,N_14863);
or U17247 (N_17247,N_14744,N_15562);
xnor U17248 (N_17248,N_15284,N_15005);
nand U17249 (N_17249,N_15454,N_15960);
and U17250 (N_17250,N_14643,N_15171);
nor U17251 (N_17251,N_15935,N_15417);
or U17252 (N_17252,N_14010,N_14431);
nand U17253 (N_17253,N_15024,N_15454);
nor U17254 (N_17254,N_14245,N_14704);
xnor U17255 (N_17255,N_15719,N_14543);
xor U17256 (N_17256,N_14744,N_15363);
xor U17257 (N_17257,N_15324,N_15723);
and U17258 (N_17258,N_15240,N_15988);
or U17259 (N_17259,N_14108,N_15193);
nor U17260 (N_17260,N_15869,N_15603);
xor U17261 (N_17261,N_15039,N_14163);
or U17262 (N_17262,N_15940,N_15499);
and U17263 (N_17263,N_14788,N_14462);
or U17264 (N_17264,N_15850,N_15183);
nor U17265 (N_17265,N_14602,N_15112);
nand U17266 (N_17266,N_14384,N_14879);
and U17267 (N_17267,N_15523,N_14075);
nand U17268 (N_17268,N_15319,N_14746);
nand U17269 (N_17269,N_14087,N_15325);
and U17270 (N_17270,N_14833,N_15373);
or U17271 (N_17271,N_14414,N_14536);
nor U17272 (N_17272,N_14485,N_15371);
nor U17273 (N_17273,N_14682,N_15566);
nor U17274 (N_17274,N_15854,N_14563);
or U17275 (N_17275,N_14749,N_15254);
or U17276 (N_17276,N_15012,N_15170);
nor U17277 (N_17277,N_15142,N_15687);
and U17278 (N_17278,N_15963,N_14716);
and U17279 (N_17279,N_14823,N_15634);
nor U17280 (N_17280,N_14387,N_14986);
xor U17281 (N_17281,N_15170,N_15222);
and U17282 (N_17282,N_14230,N_14920);
nor U17283 (N_17283,N_14671,N_15721);
nand U17284 (N_17284,N_15592,N_14566);
and U17285 (N_17285,N_15922,N_15603);
and U17286 (N_17286,N_15002,N_15684);
xnor U17287 (N_17287,N_14457,N_14615);
xnor U17288 (N_17288,N_15077,N_15944);
nor U17289 (N_17289,N_15221,N_14852);
xnor U17290 (N_17290,N_14385,N_15670);
or U17291 (N_17291,N_15959,N_14399);
nor U17292 (N_17292,N_14785,N_14765);
nand U17293 (N_17293,N_14736,N_15749);
nand U17294 (N_17294,N_15712,N_14066);
nor U17295 (N_17295,N_14651,N_14992);
nor U17296 (N_17296,N_15642,N_14050);
or U17297 (N_17297,N_14210,N_14125);
nand U17298 (N_17298,N_15142,N_14377);
or U17299 (N_17299,N_15691,N_14535);
nor U17300 (N_17300,N_15777,N_15513);
nor U17301 (N_17301,N_14455,N_15956);
xor U17302 (N_17302,N_14492,N_14713);
xnor U17303 (N_17303,N_15621,N_14853);
xnor U17304 (N_17304,N_15490,N_15330);
xor U17305 (N_17305,N_14957,N_14682);
and U17306 (N_17306,N_14580,N_14620);
nand U17307 (N_17307,N_14677,N_15653);
nor U17308 (N_17308,N_15254,N_15417);
or U17309 (N_17309,N_14903,N_15160);
nor U17310 (N_17310,N_14975,N_14876);
and U17311 (N_17311,N_15430,N_14313);
nor U17312 (N_17312,N_15185,N_14414);
and U17313 (N_17313,N_15660,N_15982);
nand U17314 (N_17314,N_15874,N_14342);
nand U17315 (N_17315,N_14281,N_14580);
xnor U17316 (N_17316,N_15570,N_15522);
xor U17317 (N_17317,N_15658,N_15190);
nand U17318 (N_17318,N_15793,N_15439);
xor U17319 (N_17319,N_14474,N_15921);
nor U17320 (N_17320,N_15340,N_14451);
xor U17321 (N_17321,N_14250,N_14869);
and U17322 (N_17322,N_15309,N_14255);
nor U17323 (N_17323,N_14659,N_15407);
nand U17324 (N_17324,N_15142,N_14665);
or U17325 (N_17325,N_15642,N_15060);
xnor U17326 (N_17326,N_15476,N_14269);
nand U17327 (N_17327,N_15108,N_14259);
xor U17328 (N_17328,N_14099,N_15451);
and U17329 (N_17329,N_14094,N_15017);
and U17330 (N_17330,N_14639,N_14152);
nor U17331 (N_17331,N_14515,N_15031);
and U17332 (N_17332,N_15947,N_14405);
xnor U17333 (N_17333,N_14180,N_14772);
or U17334 (N_17334,N_14658,N_15093);
nor U17335 (N_17335,N_14877,N_14340);
nor U17336 (N_17336,N_15170,N_15705);
xnor U17337 (N_17337,N_15688,N_15615);
or U17338 (N_17338,N_14981,N_14848);
xor U17339 (N_17339,N_15887,N_15109);
nor U17340 (N_17340,N_14188,N_14682);
xor U17341 (N_17341,N_14959,N_15937);
nor U17342 (N_17342,N_15027,N_14305);
and U17343 (N_17343,N_14506,N_15313);
nor U17344 (N_17344,N_15077,N_14126);
or U17345 (N_17345,N_14159,N_14120);
xnor U17346 (N_17346,N_15675,N_15167);
nor U17347 (N_17347,N_14804,N_15545);
xor U17348 (N_17348,N_14608,N_15458);
or U17349 (N_17349,N_14289,N_15447);
nand U17350 (N_17350,N_14931,N_14887);
and U17351 (N_17351,N_15846,N_14682);
nand U17352 (N_17352,N_14154,N_14786);
nor U17353 (N_17353,N_15224,N_15693);
nand U17354 (N_17354,N_14311,N_15720);
nand U17355 (N_17355,N_15864,N_15807);
and U17356 (N_17356,N_15933,N_14938);
nor U17357 (N_17357,N_14578,N_15460);
xor U17358 (N_17358,N_15356,N_14773);
nor U17359 (N_17359,N_15618,N_15868);
nand U17360 (N_17360,N_14349,N_15273);
and U17361 (N_17361,N_15839,N_14577);
nand U17362 (N_17362,N_15216,N_14763);
nand U17363 (N_17363,N_15418,N_15429);
or U17364 (N_17364,N_15400,N_14958);
xnor U17365 (N_17365,N_14188,N_15762);
xnor U17366 (N_17366,N_15840,N_14653);
nor U17367 (N_17367,N_14325,N_15732);
or U17368 (N_17368,N_14936,N_14552);
or U17369 (N_17369,N_14944,N_14883);
nand U17370 (N_17370,N_15611,N_15584);
and U17371 (N_17371,N_14462,N_15351);
xor U17372 (N_17372,N_15758,N_15136);
xor U17373 (N_17373,N_14630,N_14431);
and U17374 (N_17374,N_14873,N_15775);
nand U17375 (N_17375,N_14952,N_15099);
nor U17376 (N_17376,N_14235,N_15028);
or U17377 (N_17377,N_15630,N_15777);
nor U17378 (N_17378,N_15007,N_14836);
and U17379 (N_17379,N_15802,N_15736);
or U17380 (N_17380,N_15832,N_14471);
xnor U17381 (N_17381,N_14192,N_15493);
nand U17382 (N_17382,N_14166,N_15160);
and U17383 (N_17383,N_14041,N_14507);
or U17384 (N_17384,N_14409,N_15590);
and U17385 (N_17385,N_14774,N_15797);
or U17386 (N_17386,N_14455,N_15307);
nor U17387 (N_17387,N_14440,N_14884);
or U17388 (N_17388,N_14796,N_14870);
nor U17389 (N_17389,N_14718,N_15521);
nand U17390 (N_17390,N_15515,N_15695);
and U17391 (N_17391,N_15833,N_14664);
xor U17392 (N_17392,N_14532,N_15860);
or U17393 (N_17393,N_14011,N_14472);
and U17394 (N_17394,N_15105,N_15477);
and U17395 (N_17395,N_15840,N_15127);
and U17396 (N_17396,N_14506,N_14511);
nor U17397 (N_17397,N_14319,N_14210);
xnor U17398 (N_17398,N_15781,N_15694);
xor U17399 (N_17399,N_14403,N_14000);
nand U17400 (N_17400,N_14241,N_14756);
xor U17401 (N_17401,N_14269,N_14962);
xnor U17402 (N_17402,N_14072,N_14514);
xnor U17403 (N_17403,N_14700,N_15119);
xor U17404 (N_17404,N_14164,N_15822);
or U17405 (N_17405,N_14804,N_14858);
xnor U17406 (N_17406,N_15011,N_14529);
and U17407 (N_17407,N_15696,N_14774);
and U17408 (N_17408,N_14395,N_14845);
and U17409 (N_17409,N_14179,N_15016);
nor U17410 (N_17410,N_15445,N_15648);
and U17411 (N_17411,N_15174,N_14580);
xor U17412 (N_17412,N_15475,N_14230);
xnor U17413 (N_17413,N_14541,N_14272);
xnor U17414 (N_17414,N_15547,N_14825);
nor U17415 (N_17415,N_15590,N_15756);
nor U17416 (N_17416,N_15337,N_15043);
nor U17417 (N_17417,N_15814,N_14617);
xor U17418 (N_17418,N_14859,N_14632);
or U17419 (N_17419,N_15802,N_14068);
nor U17420 (N_17420,N_14698,N_14164);
and U17421 (N_17421,N_15586,N_14670);
and U17422 (N_17422,N_15990,N_14655);
and U17423 (N_17423,N_14740,N_15854);
or U17424 (N_17424,N_15080,N_14830);
and U17425 (N_17425,N_14278,N_15426);
xnor U17426 (N_17426,N_15444,N_15762);
xnor U17427 (N_17427,N_14317,N_14472);
and U17428 (N_17428,N_15457,N_14447);
xor U17429 (N_17429,N_15713,N_15630);
nor U17430 (N_17430,N_15815,N_15272);
or U17431 (N_17431,N_14117,N_15576);
nand U17432 (N_17432,N_15963,N_14562);
nand U17433 (N_17433,N_15624,N_14575);
nand U17434 (N_17434,N_15585,N_14644);
or U17435 (N_17435,N_14121,N_15741);
xor U17436 (N_17436,N_15743,N_15883);
xnor U17437 (N_17437,N_14918,N_14354);
nor U17438 (N_17438,N_14845,N_15720);
and U17439 (N_17439,N_14761,N_14121);
and U17440 (N_17440,N_14338,N_14111);
nor U17441 (N_17441,N_14462,N_14533);
and U17442 (N_17442,N_15478,N_14864);
nor U17443 (N_17443,N_15844,N_14218);
nand U17444 (N_17444,N_15323,N_14043);
xor U17445 (N_17445,N_15783,N_15698);
and U17446 (N_17446,N_15563,N_15187);
and U17447 (N_17447,N_14217,N_14490);
and U17448 (N_17448,N_15938,N_15721);
xnor U17449 (N_17449,N_15861,N_15242);
or U17450 (N_17450,N_15729,N_15211);
nand U17451 (N_17451,N_15289,N_14633);
or U17452 (N_17452,N_15393,N_15649);
xnor U17453 (N_17453,N_15711,N_14416);
and U17454 (N_17454,N_14803,N_15461);
nor U17455 (N_17455,N_14728,N_15628);
and U17456 (N_17456,N_15681,N_15647);
nor U17457 (N_17457,N_15211,N_15194);
nor U17458 (N_17458,N_14298,N_14295);
nand U17459 (N_17459,N_15311,N_15478);
nor U17460 (N_17460,N_14297,N_14977);
and U17461 (N_17461,N_15050,N_15395);
xnor U17462 (N_17462,N_14169,N_14277);
xor U17463 (N_17463,N_15813,N_15670);
nand U17464 (N_17464,N_14716,N_14430);
or U17465 (N_17465,N_15918,N_14158);
and U17466 (N_17466,N_15455,N_15565);
or U17467 (N_17467,N_15850,N_14340);
or U17468 (N_17468,N_14135,N_14475);
and U17469 (N_17469,N_15680,N_15059);
xor U17470 (N_17470,N_15619,N_14458);
or U17471 (N_17471,N_14149,N_14253);
xnor U17472 (N_17472,N_14635,N_14123);
nand U17473 (N_17473,N_14169,N_14579);
nand U17474 (N_17474,N_15887,N_14010);
or U17475 (N_17475,N_15556,N_15403);
xor U17476 (N_17476,N_15878,N_14087);
or U17477 (N_17477,N_15472,N_15515);
and U17478 (N_17478,N_14482,N_14384);
or U17479 (N_17479,N_14594,N_15308);
nor U17480 (N_17480,N_15371,N_15693);
xor U17481 (N_17481,N_14956,N_14020);
nand U17482 (N_17482,N_14331,N_14465);
nand U17483 (N_17483,N_15963,N_15806);
nand U17484 (N_17484,N_14715,N_15422);
xor U17485 (N_17485,N_15446,N_15331);
and U17486 (N_17486,N_14444,N_15006);
nor U17487 (N_17487,N_14234,N_14850);
xor U17488 (N_17488,N_15420,N_14896);
nor U17489 (N_17489,N_14300,N_14945);
and U17490 (N_17490,N_14219,N_15431);
nor U17491 (N_17491,N_15618,N_14900);
or U17492 (N_17492,N_14252,N_15317);
and U17493 (N_17493,N_14046,N_14117);
nor U17494 (N_17494,N_14150,N_14600);
nor U17495 (N_17495,N_15273,N_15582);
nand U17496 (N_17496,N_14527,N_15283);
xor U17497 (N_17497,N_14042,N_15301);
or U17498 (N_17498,N_15434,N_15502);
or U17499 (N_17499,N_15845,N_14940);
and U17500 (N_17500,N_14001,N_15987);
nor U17501 (N_17501,N_15850,N_15060);
nor U17502 (N_17502,N_14756,N_15930);
and U17503 (N_17503,N_15466,N_15337);
and U17504 (N_17504,N_15296,N_14869);
or U17505 (N_17505,N_15902,N_14344);
nor U17506 (N_17506,N_15971,N_15369);
or U17507 (N_17507,N_14118,N_15853);
nand U17508 (N_17508,N_15450,N_14705);
or U17509 (N_17509,N_15232,N_15886);
nor U17510 (N_17510,N_14482,N_15249);
nor U17511 (N_17511,N_14090,N_15753);
xor U17512 (N_17512,N_15197,N_15424);
nor U17513 (N_17513,N_15175,N_14012);
or U17514 (N_17514,N_14259,N_15417);
xor U17515 (N_17515,N_14603,N_14794);
nor U17516 (N_17516,N_14649,N_14715);
and U17517 (N_17517,N_15610,N_15804);
or U17518 (N_17518,N_14201,N_14712);
and U17519 (N_17519,N_14582,N_15126);
nor U17520 (N_17520,N_15740,N_14027);
and U17521 (N_17521,N_14682,N_14903);
nor U17522 (N_17522,N_15936,N_15356);
and U17523 (N_17523,N_15768,N_15949);
xor U17524 (N_17524,N_15318,N_15705);
and U17525 (N_17525,N_14393,N_14080);
or U17526 (N_17526,N_15567,N_14869);
and U17527 (N_17527,N_15768,N_14011);
nand U17528 (N_17528,N_14665,N_14125);
nor U17529 (N_17529,N_14431,N_14328);
or U17530 (N_17530,N_14153,N_15259);
xor U17531 (N_17531,N_14906,N_15287);
xor U17532 (N_17532,N_15047,N_15569);
nor U17533 (N_17533,N_14987,N_15276);
and U17534 (N_17534,N_15617,N_15428);
nand U17535 (N_17535,N_15456,N_14057);
xnor U17536 (N_17536,N_15000,N_14423);
and U17537 (N_17537,N_14632,N_15786);
nor U17538 (N_17538,N_15646,N_15025);
nand U17539 (N_17539,N_14456,N_14778);
nand U17540 (N_17540,N_14755,N_15705);
or U17541 (N_17541,N_15169,N_15527);
or U17542 (N_17542,N_14391,N_15237);
xor U17543 (N_17543,N_14246,N_14649);
or U17544 (N_17544,N_15681,N_15377);
nor U17545 (N_17545,N_14012,N_14316);
and U17546 (N_17546,N_14036,N_15237);
and U17547 (N_17547,N_15846,N_14931);
xnor U17548 (N_17548,N_15637,N_14205);
or U17549 (N_17549,N_14145,N_14675);
nand U17550 (N_17550,N_14569,N_15635);
xor U17551 (N_17551,N_15399,N_14053);
nand U17552 (N_17552,N_15696,N_15014);
xor U17553 (N_17553,N_15917,N_15267);
nand U17554 (N_17554,N_14360,N_14973);
nor U17555 (N_17555,N_15968,N_15447);
nand U17556 (N_17556,N_15594,N_14486);
nand U17557 (N_17557,N_14724,N_14472);
nor U17558 (N_17558,N_15706,N_14416);
xor U17559 (N_17559,N_14641,N_15416);
nor U17560 (N_17560,N_14787,N_15663);
xor U17561 (N_17561,N_14127,N_14207);
xnor U17562 (N_17562,N_14908,N_14986);
and U17563 (N_17563,N_15644,N_15112);
or U17564 (N_17564,N_14293,N_14691);
and U17565 (N_17565,N_15372,N_15000);
or U17566 (N_17566,N_15851,N_15584);
and U17567 (N_17567,N_15072,N_14280);
nor U17568 (N_17568,N_14978,N_15574);
xnor U17569 (N_17569,N_14316,N_14947);
xor U17570 (N_17570,N_14340,N_15340);
nand U17571 (N_17571,N_14770,N_14120);
xor U17572 (N_17572,N_15799,N_14922);
and U17573 (N_17573,N_14149,N_14110);
nand U17574 (N_17574,N_14827,N_15151);
nand U17575 (N_17575,N_14860,N_14504);
or U17576 (N_17576,N_14273,N_14103);
xnor U17577 (N_17577,N_15653,N_15546);
and U17578 (N_17578,N_14235,N_14482);
nor U17579 (N_17579,N_15320,N_14144);
and U17580 (N_17580,N_15902,N_14320);
nor U17581 (N_17581,N_15620,N_14265);
or U17582 (N_17582,N_14220,N_15112);
and U17583 (N_17583,N_14189,N_14576);
xor U17584 (N_17584,N_14568,N_15554);
xor U17585 (N_17585,N_15554,N_15918);
nor U17586 (N_17586,N_14294,N_14664);
xor U17587 (N_17587,N_15011,N_15758);
and U17588 (N_17588,N_15731,N_15989);
xnor U17589 (N_17589,N_15740,N_15232);
or U17590 (N_17590,N_15160,N_14345);
or U17591 (N_17591,N_15168,N_14986);
and U17592 (N_17592,N_14659,N_15078);
xnor U17593 (N_17593,N_15374,N_15978);
or U17594 (N_17594,N_15419,N_15795);
or U17595 (N_17595,N_15877,N_15303);
or U17596 (N_17596,N_14371,N_15426);
nand U17597 (N_17597,N_15257,N_14460);
xor U17598 (N_17598,N_15340,N_15726);
and U17599 (N_17599,N_15669,N_15525);
nor U17600 (N_17600,N_15712,N_14191);
nor U17601 (N_17601,N_14658,N_14435);
and U17602 (N_17602,N_14333,N_14706);
xor U17603 (N_17603,N_15419,N_14957);
nand U17604 (N_17604,N_14089,N_15362);
xor U17605 (N_17605,N_14110,N_14488);
nor U17606 (N_17606,N_14745,N_15628);
and U17607 (N_17607,N_15688,N_15058);
nor U17608 (N_17608,N_14283,N_14037);
nand U17609 (N_17609,N_15873,N_14922);
and U17610 (N_17610,N_15998,N_15278);
and U17611 (N_17611,N_14349,N_14379);
and U17612 (N_17612,N_14579,N_14417);
xor U17613 (N_17613,N_15455,N_15577);
and U17614 (N_17614,N_14769,N_15226);
or U17615 (N_17615,N_14612,N_15988);
xor U17616 (N_17616,N_15427,N_15184);
nor U17617 (N_17617,N_14007,N_14215);
or U17618 (N_17618,N_15792,N_14011);
or U17619 (N_17619,N_14765,N_14306);
nor U17620 (N_17620,N_14685,N_15966);
and U17621 (N_17621,N_15857,N_15790);
xor U17622 (N_17622,N_14028,N_14478);
and U17623 (N_17623,N_14470,N_15893);
or U17624 (N_17624,N_15904,N_15435);
nor U17625 (N_17625,N_14171,N_15896);
nand U17626 (N_17626,N_14466,N_14713);
nand U17627 (N_17627,N_15211,N_14176);
nand U17628 (N_17628,N_15318,N_15765);
nor U17629 (N_17629,N_15520,N_14477);
or U17630 (N_17630,N_15532,N_14604);
xor U17631 (N_17631,N_14873,N_15921);
nor U17632 (N_17632,N_14789,N_14447);
xor U17633 (N_17633,N_15476,N_15960);
or U17634 (N_17634,N_14229,N_14848);
or U17635 (N_17635,N_15869,N_14899);
or U17636 (N_17636,N_14232,N_14163);
or U17637 (N_17637,N_15436,N_15097);
nor U17638 (N_17638,N_15862,N_15518);
xor U17639 (N_17639,N_14719,N_15399);
nor U17640 (N_17640,N_14642,N_15255);
nand U17641 (N_17641,N_14632,N_14440);
nor U17642 (N_17642,N_14691,N_14115);
and U17643 (N_17643,N_15975,N_15725);
xnor U17644 (N_17644,N_15354,N_15930);
or U17645 (N_17645,N_14749,N_15030);
xnor U17646 (N_17646,N_15119,N_15217);
nand U17647 (N_17647,N_15112,N_15721);
nand U17648 (N_17648,N_14927,N_15827);
nor U17649 (N_17649,N_14766,N_14207);
or U17650 (N_17650,N_15821,N_14167);
and U17651 (N_17651,N_15443,N_14931);
xor U17652 (N_17652,N_14126,N_14960);
and U17653 (N_17653,N_15804,N_14486);
and U17654 (N_17654,N_15969,N_14207);
nand U17655 (N_17655,N_14069,N_15908);
and U17656 (N_17656,N_14166,N_15587);
xor U17657 (N_17657,N_15268,N_14541);
nor U17658 (N_17658,N_14917,N_15613);
xnor U17659 (N_17659,N_15911,N_14598);
nor U17660 (N_17660,N_15876,N_14850);
xor U17661 (N_17661,N_14298,N_14950);
xor U17662 (N_17662,N_14028,N_15290);
and U17663 (N_17663,N_14411,N_14232);
xor U17664 (N_17664,N_14451,N_15085);
or U17665 (N_17665,N_15940,N_15745);
nand U17666 (N_17666,N_14541,N_15972);
nor U17667 (N_17667,N_14064,N_14960);
nand U17668 (N_17668,N_15448,N_15124);
or U17669 (N_17669,N_15523,N_15297);
and U17670 (N_17670,N_15551,N_14333);
or U17671 (N_17671,N_14417,N_14050);
or U17672 (N_17672,N_15502,N_14157);
nor U17673 (N_17673,N_14285,N_15040);
nand U17674 (N_17674,N_15582,N_15461);
or U17675 (N_17675,N_15599,N_15421);
and U17676 (N_17676,N_14821,N_15431);
xor U17677 (N_17677,N_14740,N_14080);
xnor U17678 (N_17678,N_14364,N_15943);
nand U17679 (N_17679,N_14236,N_14347);
nand U17680 (N_17680,N_14090,N_14826);
xor U17681 (N_17681,N_15211,N_14304);
or U17682 (N_17682,N_14526,N_14951);
nor U17683 (N_17683,N_14670,N_14141);
nor U17684 (N_17684,N_15908,N_14028);
nand U17685 (N_17685,N_15505,N_15448);
xnor U17686 (N_17686,N_15366,N_15894);
xnor U17687 (N_17687,N_15084,N_15925);
xor U17688 (N_17688,N_14517,N_15290);
xor U17689 (N_17689,N_15995,N_15806);
nand U17690 (N_17690,N_15088,N_14885);
xnor U17691 (N_17691,N_14417,N_14975);
nor U17692 (N_17692,N_14114,N_15753);
xnor U17693 (N_17693,N_15509,N_14021);
nand U17694 (N_17694,N_15278,N_15746);
and U17695 (N_17695,N_14417,N_15645);
nand U17696 (N_17696,N_15774,N_14271);
and U17697 (N_17697,N_14638,N_15372);
or U17698 (N_17698,N_15020,N_14231);
nand U17699 (N_17699,N_15633,N_15519);
and U17700 (N_17700,N_14129,N_14383);
nand U17701 (N_17701,N_15653,N_14392);
nand U17702 (N_17702,N_15478,N_14362);
or U17703 (N_17703,N_14167,N_15491);
nor U17704 (N_17704,N_14684,N_15146);
or U17705 (N_17705,N_15352,N_14318);
and U17706 (N_17706,N_14676,N_14470);
nand U17707 (N_17707,N_15398,N_14016);
nor U17708 (N_17708,N_15294,N_14095);
nand U17709 (N_17709,N_15350,N_14177);
and U17710 (N_17710,N_15939,N_14937);
or U17711 (N_17711,N_14368,N_15989);
xnor U17712 (N_17712,N_15483,N_14193);
nand U17713 (N_17713,N_15164,N_15598);
or U17714 (N_17714,N_14602,N_14320);
xor U17715 (N_17715,N_14199,N_14656);
nor U17716 (N_17716,N_15662,N_15930);
or U17717 (N_17717,N_15993,N_15702);
and U17718 (N_17718,N_15225,N_15577);
xnor U17719 (N_17719,N_15581,N_14961);
and U17720 (N_17720,N_14432,N_14874);
xnor U17721 (N_17721,N_15541,N_15041);
xor U17722 (N_17722,N_15019,N_15170);
nand U17723 (N_17723,N_15855,N_14159);
nor U17724 (N_17724,N_15727,N_15031);
nor U17725 (N_17725,N_15704,N_15458);
xnor U17726 (N_17726,N_14952,N_14411);
or U17727 (N_17727,N_14127,N_14049);
or U17728 (N_17728,N_15392,N_14114);
nand U17729 (N_17729,N_15437,N_15710);
or U17730 (N_17730,N_15770,N_14371);
nor U17731 (N_17731,N_14442,N_15720);
and U17732 (N_17732,N_15255,N_15426);
nor U17733 (N_17733,N_15692,N_14217);
xnor U17734 (N_17734,N_14424,N_14026);
or U17735 (N_17735,N_14898,N_15130);
xor U17736 (N_17736,N_14927,N_15356);
xnor U17737 (N_17737,N_14265,N_14140);
or U17738 (N_17738,N_14847,N_14922);
xor U17739 (N_17739,N_15433,N_14405);
xnor U17740 (N_17740,N_14266,N_15617);
nor U17741 (N_17741,N_15061,N_14473);
nor U17742 (N_17742,N_14193,N_14132);
nor U17743 (N_17743,N_14374,N_15542);
xor U17744 (N_17744,N_15784,N_14793);
or U17745 (N_17745,N_14398,N_14420);
xnor U17746 (N_17746,N_14031,N_14627);
nor U17747 (N_17747,N_15259,N_14159);
or U17748 (N_17748,N_15578,N_15594);
nand U17749 (N_17749,N_14659,N_15479);
xor U17750 (N_17750,N_15511,N_14656);
and U17751 (N_17751,N_14498,N_15588);
nor U17752 (N_17752,N_15912,N_15670);
nand U17753 (N_17753,N_15411,N_14659);
xor U17754 (N_17754,N_15310,N_15491);
or U17755 (N_17755,N_15789,N_14792);
nand U17756 (N_17756,N_15926,N_14197);
and U17757 (N_17757,N_15243,N_14920);
nand U17758 (N_17758,N_15518,N_15694);
and U17759 (N_17759,N_15077,N_14906);
or U17760 (N_17760,N_14821,N_15860);
nor U17761 (N_17761,N_14979,N_15091);
nor U17762 (N_17762,N_15462,N_14372);
xor U17763 (N_17763,N_14245,N_15767);
or U17764 (N_17764,N_14855,N_14207);
or U17765 (N_17765,N_15801,N_15142);
or U17766 (N_17766,N_15331,N_14766);
or U17767 (N_17767,N_14044,N_15014);
nand U17768 (N_17768,N_15764,N_15298);
or U17769 (N_17769,N_14481,N_15387);
nand U17770 (N_17770,N_15252,N_15432);
nand U17771 (N_17771,N_15658,N_15371);
nand U17772 (N_17772,N_15389,N_14772);
nor U17773 (N_17773,N_15322,N_15348);
nor U17774 (N_17774,N_15659,N_14782);
and U17775 (N_17775,N_15363,N_14387);
or U17776 (N_17776,N_14142,N_14711);
nand U17777 (N_17777,N_14220,N_14665);
xor U17778 (N_17778,N_14103,N_15932);
nor U17779 (N_17779,N_15220,N_15916);
xor U17780 (N_17780,N_15736,N_14817);
nand U17781 (N_17781,N_14189,N_14713);
xnor U17782 (N_17782,N_15249,N_15343);
nand U17783 (N_17783,N_15211,N_15042);
and U17784 (N_17784,N_15011,N_14895);
and U17785 (N_17785,N_14028,N_14052);
and U17786 (N_17786,N_15958,N_14431);
nor U17787 (N_17787,N_14354,N_14757);
xor U17788 (N_17788,N_14387,N_14811);
and U17789 (N_17789,N_15185,N_15658);
nor U17790 (N_17790,N_14028,N_14815);
and U17791 (N_17791,N_14247,N_14835);
nand U17792 (N_17792,N_15879,N_14083);
or U17793 (N_17793,N_14856,N_15343);
or U17794 (N_17794,N_14923,N_15023);
nor U17795 (N_17795,N_15517,N_14147);
nand U17796 (N_17796,N_15972,N_14344);
xor U17797 (N_17797,N_15567,N_15791);
and U17798 (N_17798,N_15589,N_15096);
or U17799 (N_17799,N_14255,N_14932);
or U17800 (N_17800,N_14134,N_14032);
nand U17801 (N_17801,N_14382,N_15244);
xnor U17802 (N_17802,N_15872,N_15354);
or U17803 (N_17803,N_15242,N_15536);
nor U17804 (N_17804,N_14582,N_14272);
nor U17805 (N_17805,N_14807,N_15930);
xnor U17806 (N_17806,N_15724,N_14393);
and U17807 (N_17807,N_15511,N_14104);
and U17808 (N_17808,N_15159,N_15678);
and U17809 (N_17809,N_14814,N_14678);
and U17810 (N_17810,N_14058,N_15348);
nor U17811 (N_17811,N_14375,N_14494);
nor U17812 (N_17812,N_14248,N_14168);
and U17813 (N_17813,N_15711,N_14410);
xor U17814 (N_17814,N_14622,N_15186);
and U17815 (N_17815,N_14300,N_14295);
nand U17816 (N_17816,N_15182,N_14641);
or U17817 (N_17817,N_15825,N_15258);
nor U17818 (N_17818,N_14387,N_14152);
or U17819 (N_17819,N_14300,N_14343);
nor U17820 (N_17820,N_15062,N_14903);
and U17821 (N_17821,N_14285,N_15025);
and U17822 (N_17822,N_14179,N_14326);
nand U17823 (N_17823,N_14132,N_14699);
or U17824 (N_17824,N_15078,N_14714);
nor U17825 (N_17825,N_14474,N_14698);
xnor U17826 (N_17826,N_14757,N_15146);
or U17827 (N_17827,N_14560,N_15624);
and U17828 (N_17828,N_15129,N_14631);
or U17829 (N_17829,N_14110,N_14659);
nand U17830 (N_17830,N_15509,N_14549);
and U17831 (N_17831,N_14819,N_14417);
and U17832 (N_17832,N_15624,N_15466);
xnor U17833 (N_17833,N_14914,N_15330);
xor U17834 (N_17834,N_15393,N_15587);
and U17835 (N_17835,N_15550,N_15864);
nor U17836 (N_17836,N_15948,N_15199);
nor U17837 (N_17837,N_14178,N_14206);
nor U17838 (N_17838,N_14593,N_15774);
and U17839 (N_17839,N_14580,N_14297);
and U17840 (N_17840,N_14603,N_15006);
and U17841 (N_17841,N_15679,N_14122);
xnor U17842 (N_17842,N_15021,N_14807);
and U17843 (N_17843,N_15689,N_14308);
and U17844 (N_17844,N_15340,N_15385);
nor U17845 (N_17845,N_15641,N_14508);
and U17846 (N_17846,N_15887,N_15372);
nand U17847 (N_17847,N_15490,N_14906);
or U17848 (N_17848,N_14850,N_15534);
xnor U17849 (N_17849,N_15751,N_15378);
nand U17850 (N_17850,N_15643,N_14718);
nand U17851 (N_17851,N_14305,N_14594);
and U17852 (N_17852,N_14801,N_15261);
and U17853 (N_17853,N_15777,N_15317);
xor U17854 (N_17854,N_14086,N_14043);
nor U17855 (N_17855,N_14171,N_15040);
and U17856 (N_17856,N_14359,N_14293);
xnor U17857 (N_17857,N_14408,N_14891);
nand U17858 (N_17858,N_15322,N_14914);
or U17859 (N_17859,N_14710,N_14187);
xnor U17860 (N_17860,N_15674,N_15801);
and U17861 (N_17861,N_15614,N_15346);
nand U17862 (N_17862,N_14545,N_15454);
xor U17863 (N_17863,N_15526,N_14053);
nor U17864 (N_17864,N_14871,N_14591);
and U17865 (N_17865,N_14859,N_15484);
nand U17866 (N_17866,N_14535,N_14162);
and U17867 (N_17867,N_15720,N_15592);
xnor U17868 (N_17868,N_15057,N_15610);
nor U17869 (N_17869,N_14715,N_15551);
xor U17870 (N_17870,N_14141,N_14000);
nand U17871 (N_17871,N_14747,N_15895);
and U17872 (N_17872,N_14632,N_15413);
or U17873 (N_17873,N_14655,N_14371);
nor U17874 (N_17874,N_15425,N_15202);
and U17875 (N_17875,N_15592,N_15388);
nor U17876 (N_17876,N_14670,N_15188);
and U17877 (N_17877,N_14818,N_15173);
or U17878 (N_17878,N_15425,N_15760);
nor U17879 (N_17879,N_14849,N_15029);
or U17880 (N_17880,N_14938,N_15165);
and U17881 (N_17881,N_14004,N_15283);
nor U17882 (N_17882,N_14494,N_14737);
xor U17883 (N_17883,N_15341,N_14749);
xnor U17884 (N_17884,N_14876,N_15823);
or U17885 (N_17885,N_14109,N_15980);
nand U17886 (N_17886,N_14879,N_15173);
xor U17887 (N_17887,N_15666,N_14901);
and U17888 (N_17888,N_15130,N_15944);
xnor U17889 (N_17889,N_15018,N_14432);
xnor U17890 (N_17890,N_15528,N_15949);
nor U17891 (N_17891,N_15538,N_14525);
nor U17892 (N_17892,N_14010,N_15912);
xor U17893 (N_17893,N_14916,N_14882);
and U17894 (N_17894,N_15223,N_14067);
xor U17895 (N_17895,N_15147,N_15121);
and U17896 (N_17896,N_15179,N_15440);
and U17897 (N_17897,N_14475,N_15730);
nor U17898 (N_17898,N_15604,N_14574);
and U17899 (N_17899,N_14747,N_15165);
xnor U17900 (N_17900,N_15535,N_14661);
nand U17901 (N_17901,N_15479,N_15278);
and U17902 (N_17902,N_14931,N_15738);
or U17903 (N_17903,N_15378,N_15226);
or U17904 (N_17904,N_15521,N_14183);
and U17905 (N_17905,N_15927,N_14328);
or U17906 (N_17906,N_15866,N_14493);
or U17907 (N_17907,N_15492,N_14929);
and U17908 (N_17908,N_14683,N_15280);
xor U17909 (N_17909,N_14261,N_14423);
nor U17910 (N_17910,N_15873,N_14619);
and U17911 (N_17911,N_14468,N_14957);
nand U17912 (N_17912,N_15158,N_15718);
nand U17913 (N_17913,N_15834,N_15191);
nand U17914 (N_17914,N_14098,N_15707);
or U17915 (N_17915,N_14368,N_15756);
nor U17916 (N_17916,N_14042,N_15285);
or U17917 (N_17917,N_15675,N_15264);
nand U17918 (N_17918,N_15467,N_14886);
xor U17919 (N_17919,N_14591,N_14919);
nand U17920 (N_17920,N_14163,N_14030);
xor U17921 (N_17921,N_15775,N_14640);
and U17922 (N_17922,N_15946,N_14389);
and U17923 (N_17923,N_14028,N_15000);
xnor U17924 (N_17924,N_14919,N_15034);
nor U17925 (N_17925,N_14620,N_15895);
nor U17926 (N_17926,N_15772,N_15425);
xor U17927 (N_17927,N_14017,N_14664);
or U17928 (N_17928,N_14325,N_15634);
or U17929 (N_17929,N_15129,N_14184);
nor U17930 (N_17930,N_14131,N_14678);
xor U17931 (N_17931,N_14207,N_15904);
or U17932 (N_17932,N_15135,N_15666);
and U17933 (N_17933,N_14614,N_14398);
nand U17934 (N_17934,N_15066,N_14948);
nor U17935 (N_17935,N_15497,N_14906);
or U17936 (N_17936,N_14865,N_14964);
nor U17937 (N_17937,N_15687,N_14397);
or U17938 (N_17938,N_14993,N_14151);
nand U17939 (N_17939,N_15969,N_15000);
xor U17940 (N_17940,N_14005,N_15418);
xor U17941 (N_17941,N_15718,N_14262);
and U17942 (N_17942,N_15881,N_14397);
and U17943 (N_17943,N_15203,N_15634);
nor U17944 (N_17944,N_14555,N_14464);
nor U17945 (N_17945,N_15703,N_15931);
nand U17946 (N_17946,N_14321,N_14679);
nand U17947 (N_17947,N_15734,N_14046);
nor U17948 (N_17948,N_15643,N_14759);
nor U17949 (N_17949,N_14404,N_15801);
nand U17950 (N_17950,N_14458,N_15099);
or U17951 (N_17951,N_15674,N_15691);
or U17952 (N_17952,N_15419,N_14845);
and U17953 (N_17953,N_14113,N_15219);
nor U17954 (N_17954,N_14625,N_15134);
xnor U17955 (N_17955,N_15362,N_14420);
or U17956 (N_17956,N_14551,N_15992);
and U17957 (N_17957,N_15483,N_15305);
xnor U17958 (N_17958,N_15018,N_15641);
nand U17959 (N_17959,N_15645,N_14497);
or U17960 (N_17960,N_14079,N_14437);
nand U17961 (N_17961,N_14492,N_14962);
nand U17962 (N_17962,N_15382,N_14535);
or U17963 (N_17963,N_15241,N_14984);
nand U17964 (N_17964,N_14716,N_15936);
nor U17965 (N_17965,N_14285,N_14910);
nor U17966 (N_17966,N_14266,N_14370);
nor U17967 (N_17967,N_14678,N_15811);
or U17968 (N_17968,N_15557,N_15806);
or U17969 (N_17969,N_15254,N_14151);
nand U17970 (N_17970,N_14526,N_15680);
xor U17971 (N_17971,N_14323,N_14831);
xnor U17972 (N_17972,N_15922,N_15008);
or U17973 (N_17973,N_14351,N_14254);
or U17974 (N_17974,N_14645,N_14302);
xor U17975 (N_17975,N_15811,N_15091);
nand U17976 (N_17976,N_15981,N_15322);
xor U17977 (N_17977,N_15130,N_15016);
xor U17978 (N_17978,N_15327,N_14714);
or U17979 (N_17979,N_14607,N_15721);
or U17980 (N_17980,N_15984,N_14159);
or U17981 (N_17981,N_15024,N_15865);
or U17982 (N_17982,N_15573,N_14066);
and U17983 (N_17983,N_14405,N_14108);
or U17984 (N_17984,N_15307,N_15673);
and U17985 (N_17985,N_14944,N_14394);
nor U17986 (N_17986,N_14996,N_14457);
and U17987 (N_17987,N_15376,N_15922);
xor U17988 (N_17988,N_14071,N_14092);
nand U17989 (N_17989,N_15225,N_15560);
or U17990 (N_17990,N_15207,N_14261);
xnor U17991 (N_17991,N_15284,N_14541);
and U17992 (N_17992,N_14364,N_14623);
and U17993 (N_17993,N_14992,N_14876);
nand U17994 (N_17994,N_14135,N_14545);
nand U17995 (N_17995,N_14550,N_14956);
nor U17996 (N_17996,N_14488,N_15772);
xnor U17997 (N_17997,N_14696,N_15054);
and U17998 (N_17998,N_15152,N_15940);
and U17999 (N_17999,N_14911,N_15624);
nand U18000 (N_18000,N_16054,N_16400);
nand U18001 (N_18001,N_16607,N_16250);
nand U18002 (N_18002,N_16806,N_17094);
nand U18003 (N_18003,N_17737,N_17066);
nand U18004 (N_18004,N_16677,N_17008);
xnor U18005 (N_18005,N_17051,N_17881);
and U18006 (N_18006,N_16302,N_16043);
or U18007 (N_18007,N_16570,N_16547);
and U18008 (N_18008,N_16784,N_17560);
nand U18009 (N_18009,N_17417,N_17508);
nor U18010 (N_18010,N_17766,N_17072);
nand U18011 (N_18011,N_17432,N_16123);
nand U18012 (N_18012,N_16863,N_16275);
or U18013 (N_18013,N_17116,N_17514);
or U18014 (N_18014,N_16617,N_16800);
xnor U18015 (N_18015,N_16826,N_17654);
and U18016 (N_18016,N_16445,N_16025);
xor U18017 (N_18017,N_16239,N_17976);
nor U18018 (N_18018,N_16814,N_17305);
nor U18019 (N_18019,N_17418,N_16538);
xnor U18020 (N_18020,N_16725,N_16364);
and U18021 (N_18021,N_16961,N_16565);
or U18022 (N_18022,N_17838,N_16212);
xnor U18023 (N_18023,N_17894,N_17637);
or U18024 (N_18024,N_16661,N_16980);
or U18025 (N_18025,N_16414,N_16830);
xnor U18026 (N_18026,N_16542,N_17071);
xor U18027 (N_18027,N_17190,N_17425);
nor U18028 (N_18028,N_16341,N_17668);
and U18029 (N_18029,N_17558,N_17678);
nand U18030 (N_18030,N_16890,N_16796);
and U18031 (N_18031,N_16096,N_17500);
xor U18032 (N_18032,N_17109,N_17424);
nand U18033 (N_18033,N_17696,N_17487);
and U18034 (N_18034,N_17315,N_16995);
nand U18035 (N_18035,N_17047,N_16129);
nand U18036 (N_18036,N_16573,N_17414);
xnor U18037 (N_18037,N_17216,N_17805);
nand U18038 (N_18038,N_16376,N_17741);
nand U18039 (N_18039,N_17307,N_16606);
xor U18040 (N_18040,N_16425,N_17588);
nor U18041 (N_18041,N_16184,N_16583);
or U18042 (N_18042,N_16769,N_17222);
and U18043 (N_18043,N_17773,N_17889);
or U18044 (N_18044,N_17409,N_17785);
xnor U18045 (N_18045,N_17614,N_16053);
nand U18046 (N_18046,N_17381,N_16066);
or U18047 (N_18047,N_16355,N_17384);
nor U18048 (N_18048,N_16549,N_17787);
nand U18049 (N_18049,N_17304,N_16517);
or U18050 (N_18050,N_16035,N_17437);
nand U18051 (N_18051,N_16094,N_16602);
or U18052 (N_18052,N_17306,N_17546);
nand U18053 (N_18053,N_16640,N_16442);
and U18054 (N_18054,N_17535,N_17471);
nor U18055 (N_18055,N_17082,N_16013);
nor U18056 (N_18056,N_17323,N_17795);
and U18057 (N_18057,N_16943,N_16306);
nor U18058 (N_18058,N_17853,N_16923);
xnor U18059 (N_18059,N_17857,N_16829);
xor U18060 (N_18060,N_16393,N_17803);
nor U18061 (N_18061,N_16969,N_17922);
xnor U18062 (N_18062,N_16344,N_16865);
or U18063 (N_18063,N_16213,N_17025);
nand U18064 (N_18064,N_16145,N_17444);
nor U18065 (N_18065,N_16703,N_17911);
nor U18066 (N_18066,N_16256,N_17412);
or U18067 (N_18067,N_16480,N_16642);
or U18068 (N_18068,N_16273,N_17530);
and U18069 (N_18069,N_16597,N_17156);
nor U18070 (N_18070,N_17322,N_16497);
and U18071 (N_18071,N_17955,N_16821);
nor U18072 (N_18072,N_16085,N_17801);
and U18073 (N_18073,N_16656,N_16698);
or U18074 (N_18074,N_17860,N_17617);
nand U18075 (N_18075,N_16496,N_17090);
or U18076 (N_18076,N_16699,N_17867);
or U18077 (N_18077,N_17137,N_17790);
and U18078 (N_18078,N_17781,N_16180);
or U18079 (N_18079,N_17849,N_16763);
and U18080 (N_18080,N_17028,N_16336);
and U18081 (N_18081,N_17632,N_16433);
nor U18082 (N_18082,N_16415,N_16343);
and U18083 (N_18083,N_17296,N_17117);
xor U18084 (N_18084,N_17233,N_17415);
or U18085 (N_18085,N_16713,N_17083);
and U18086 (N_18086,N_16790,N_16081);
and U18087 (N_18087,N_16323,N_17300);
xor U18088 (N_18088,N_17239,N_17764);
and U18089 (N_18089,N_16333,N_17148);
nand U18090 (N_18090,N_17526,N_17018);
nand U18091 (N_18091,N_16188,N_17348);
or U18092 (N_18092,N_16807,N_16742);
or U18093 (N_18093,N_16566,N_16799);
nand U18094 (N_18094,N_16113,N_16981);
nor U18095 (N_18095,N_16849,N_16115);
nand U18096 (N_18096,N_16100,N_17747);
or U18097 (N_18097,N_17224,N_16190);
nor U18098 (N_18098,N_16416,N_17200);
or U18099 (N_18099,N_17055,N_16310);
xnor U18100 (N_18100,N_16417,N_16105);
or U18101 (N_18101,N_16166,N_16637);
xor U18102 (N_18102,N_16901,N_17354);
and U18103 (N_18103,N_17511,N_17796);
and U18104 (N_18104,N_17554,N_16560);
xor U18105 (N_18105,N_16241,N_16752);
xnor U18106 (N_18106,N_16216,N_16282);
and U18107 (N_18107,N_17506,N_17212);
or U18108 (N_18108,N_16244,N_16689);
or U18109 (N_18109,N_16346,N_16397);
xor U18110 (N_18110,N_16057,N_17524);
nor U18111 (N_18111,N_17847,N_16682);
and U18112 (N_18112,N_17005,N_17081);
xor U18113 (N_18113,N_16011,N_16071);
or U18114 (N_18114,N_16338,N_17121);
or U18115 (N_18115,N_17177,N_16840);
nand U18116 (N_18116,N_17656,N_16972);
nand U18117 (N_18117,N_17149,N_17006);
and U18118 (N_18118,N_17325,N_17531);
nor U18119 (N_18119,N_17794,N_16394);
nand U18120 (N_18120,N_16571,N_16381);
or U18121 (N_18121,N_17097,N_17693);
or U18122 (N_18122,N_16756,N_16975);
nand U18123 (N_18123,N_16644,N_17247);
xnor U18124 (N_18124,N_16802,N_16041);
nand U18125 (N_18125,N_17447,N_17062);
nor U18126 (N_18126,N_16002,N_17906);
or U18127 (N_18127,N_16974,N_17126);
xor U18128 (N_18128,N_17229,N_16019);
and U18129 (N_18129,N_16657,N_16751);
or U18130 (N_18130,N_17218,N_16716);
or U18131 (N_18131,N_17251,N_16858);
or U18132 (N_18132,N_16843,N_16628);
xor U18133 (N_18133,N_17744,N_16842);
nand U18134 (N_18134,N_16245,N_17618);
and U18135 (N_18135,N_16342,N_17485);
and U18136 (N_18136,N_17427,N_17862);
xnor U18137 (N_18137,N_16569,N_16490);
and U18138 (N_18138,N_16423,N_16045);
nand U18139 (N_18139,N_17966,N_16813);
xor U18140 (N_18140,N_16676,N_16841);
or U18141 (N_18141,N_16287,N_17463);
xnor U18142 (N_18142,N_16691,N_16420);
and U18143 (N_18143,N_17024,N_17320);
xor U18144 (N_18144,N_16726,N_16407);
nor U18145 (N_18145,N_17114,N_17780);
or U18146 (N_18146,N_17184,N_16238);
nand U18147 (N_18147,N_17395,N_16237);
and U18148 (N_18148,N_16776,N_17026);
and U18149 (N_18149,N_16966,N_16353);
or U18150 (N_18150,N_17878,N_17194);
xor U18151 (N_18151,N_17909,N_16697);
xnor U18152 (N_18152,N_16064,N_17002);
and U18153 (N_18153,N_17711,N_16782);
nand U18154 (N_18154,N_16902,N_17575);
or U18155 (N_18155,N_16312,N_17421);
nand U18156 (N_18156,N_17192,N_16647);
nand U18157 (N_18157,N_16383,N_17905);
nand U18158 (N_18158,N_16819,N_17646);
and U18159 (N_18159,N_17816,N_17640);
and U18160 (N_18160,N_16350,N_17494);
nand U18161 (N_18161,N_17074,N_16382);
and U18162 (N_18162,N_17830,N_17677);
or U18163 (N_18163,N_16304,N_16429);
xnor U18164 (N_18164,N_16200,N_17826);
or U18165 (N_18165,N_16828,N_16872);
or U18166 (N_18166,N_17783,N_16097);
xor U18167 (N_18167,N_17951,N_16599);
nor U18168 (N_18168,N_17918,N_17515);
nor U18169 (N_18169,N_17331,N_16040);
nand U18170 (N_18170,N_17868,N_17161);
nand U18171 (N_18171,N_17621,N_16459);
xnor U18172 (N_18172,N_16046,N_17792);
or U18173 (N_18173,N_16329,N_17267);
nor U18174 (N_18174,N_17133,N_16309);
nand U18175 (N_18175,N_17250,N_16314);
nand U18176 (N_18176,N_17666,N_17954);
and U18177 (N_18177,N_17403,N_16463);
or U18178 (N_18178,N_16673,N_16932);
nand U18179 (N_18179,N_17393,N_16210);
nor U18180 (N_18180,N_16662,N_16130);
or U18181 (N_18181,N_17579,N_17863);
nor U18182 (N_18182,N_17214,N_17478);
nand U18183 (N_18183,N_17871,N_17459);
or U18184 (N_18184,N_17410,N_17316);
nor U18185 (N_18185,N_16267,N_16369);
xnor U18186 (N_18186,N_17705,N_16598);
nor U18187 (N_18187,N_17197,N_17465);
xor U18188 (N_18188,N_17844,N_16075);
xnor U18189 (N_18189,N_17848,N_16681);
and U18190 (N_18190,N_17532,N_16715);
or U18191 (N_18191,N_16331,N_16492);
or U18192 (N_18192,N_17277,N_16710);
xor U18193 (N_18193,N_16925,N_16551);
or U18194 (N_18194,N_17353,N_16553);
and U18195 (N_18195,N_17620,N_17015);
or U18196 (N_18196,N_17908,N_17633);
nor U18197 (N_18197,N_17891,N_17750);
nand U18198 (N_18198,N_17413,N_16455);
or U18199 (N_18199,N_17399,N_16375);
xor U18200 (N_18200,N_17866,N_16162);
nand U18201 (N_18201,N_17406,N_16095);
or U18202 (N_18202,N_17897,N_17635);
nor U18203 (N_18203,N_16540,N_17347);
xnor U18204 (N_18204,N_16793,N_17574);
xnor U18205 (N_18205,N_16176,N_17375);
nor U18206 (N_18206,N_16092,N_16387);
nor U18207 (N_18207,N_17439,N_17103);
and U18208 (N_18208,N_16984,N_16852);
nand U18209 (N_18209,N_17552,N_16125);
xnor U18210 (N_18210,N_16700,N_16265);
nand U18211 (N_18211,N_17992,N_16593);
or U18212 (N_18212,N_17970,N_17742);
and U18213 (N_18213,N_16029,N_16144);
or U18214 (N_18214,N_17333,N_17130);
xor U18215 (N_18215,N_16143,N_16630);
or U18216 (N_18216,N_16724,N_17400);
nand U18217 (N_18217,N_17509,N_17598);
nor U18218 (N_18218,N_16501,N_17179);
and U18219 (N_18219,N_17964,N_17941);
and U18220 (N_18220,N_17884,N_16308);
nor U18221 (N_18221,N_16987,N_17690);
and U18222 (N_18222,N_17850,N_16937);
nand U18223 (N_18223,N_17145,N_16615);
and U18224 (N_18224,N_16514,N_17110);
xnor U18225 (N_18225,N_16515,N_16426);
nor U18226 (N_18226,N_16701,N_16744);
nor U18227 (N_18227,N_16106,N_17521);
nor U18228 (N_18228,N_17398,N_17356);
nor U18229 (N_18229,N_17920,N_17310);
nand U18230 (N_18230,N_17584,N_17147);
nor U18231 (N_18231,N_17688,N_16218);
xor U18232 (N_18232,N_16939,N_16208);
xnor U18233 (N_18233,N_17450,N_17448);
nor U18234 (N_18234,N_16935,N_17158);
or U18235 (N_18235,N_17729,N_16623);
nor U18236 (N_18236,N_16114,N_17292);
xnor U18237 (N_18237,N_17928,N_16068);
nand U18238 (N_18238,N_17469,N_16295);
xnor U18239 (N_18239,N_16665,N_17397);
or U18240 (N_18240,N_17674,N_16619);
and U18241 (N_18241,N_17776,N_17100);
xor U18242 (N_18242,N_17673,N_17800);
and U18243 (N_18243,N_17276,N_17483);
nand U18244 (N_18244,N_17502,N_17893);
nand U18245 (N_18245,N_17163,N_17237);
and U18246 (N_18246,N_16797,N_17470);
xnor U18247 (N_18247,N_16452,N_16518);
and U18248 (N_18248,N_16942,N_16652);
nand U18249 (N_18249,N_17252,N_17468);
or U18250 (N_18250,N_16528,N_16122);
xor U18251 (N_18251,N_17176,N_17030);
and U18252 (N_18252,N_17504,N_17942);
nand U18253 (N_18253,N_17544,N_16946);
nor U18254 (N_18254,N_17359,N_17767);
nor U18255 (N_18255,N_17203,N_16436);
nor U18256 (N_18256,N_17570,N_17022);
or U18257 (N_18257,N_17289,N_16608);
and U18258 (N_18258,N_16891,N_16734);
and U18259 (N_18259,N_16042,N_16610);
and U18260 (N_18260,N_16747,N_16368);
or U18261 (N_18261,N_16303,N_17645);
nor U18262 (N_18262,N_17698,N_17856);
or U18263 (N_18263,N_16795,N_16307);
nor U18264 (N_18264,N_17726,N_16757);
nor U18265 (N_18265,N_16945,N_17076);
xor U18266 (N_18266,N_17340,N_17533);
or U18267 (N_18267,N_17612,N_16531);
nor U18268 (N_18268,N_16242,N_16067);
and U18269 (N_18269,N_17983,N_16773);
nand U18270 (N_18270,N_17473,N_17971);
xnor U18271 (N_18271,N_17091,N_16552);
or U18272 (N_18272,N_17428,N_17843);
or U18273 (N_18273,N_17754,N_17536);
xor U18274 (N_18274,N_17105,N_17311);
or U18275 (N_18275,N_17935,N_16908);
or U18276 (N_18276,N_17590,N_17609);
nor U18277 (N_18277,N_17649,N_17129);
xor U18278 (N_18278,N_16198,N_16627);
nand U18279 (N_18279,N_16709,N_17962);
nor U18280 (N_18280,N_17073,N_17832);
or U18281 (N_18281,N_16228,N_17016);
nand U18282 (N_18282,N_17700,N_16207);
and U18283 (N_18283,N_17321,N_17038);
or U18284 (N_18284,N_17260,N_16900);
nor U18285 (N_18285,N_16008,N_16133);
nand U18286 (N_18286,N_16386,N_16181);
and U18287 (N_18287,N_16476,N_16823);
nor U18288 (N_18288,N_16648,N_17128);
nor U18289 (N_18289,N_16495,N_17762);
and U18290 (N_18290,N_16360,N_17630);
or U18291 (N_18291,N_17628,N_16033);
and U18292 (N_18292,N_17739,N_16913);
xnor U18293 (N_18293,N_17175,N_17749);
or U18294 (N_18294,N_17341,N_16246);
nand U18295 (N_18295,N_16579,N_16958);
or U18296 (N_18296,N_17288,N_17572);
xor U18297 (N_18297,N_17926,N_16948);
and U18298 (N_18298,N_17594,N_16158);
nand U18299 (N_18299,N_16880,N_16535);
xnor U18300 (N_18300,N_16846,N_17733);
xnor U18301 (N_18301,N_17360,N_16051);
nor U18302 (N_18302,N_17576,N_16587);
nand U18303 (N_18303,N_17188,N_16848);
and U18304 (N_18304,N_17187,N_16151);
or U18305 (N_18305,N_17170,N_17591);
xnor U18306 (N_18306,N_16674,N_16050);
nand U18307 (N_18307,N_16996,N_16283);
or U18308 (N_18308,N_17706,N_16301);
nor U18309 (N_18309,N_16924,N_16613);
or U18310 (N_18310,N_16477,N_17346);
nand U18311 (N_18311,N_17461,N_16847);
or U18312 (N_18312,N_16855,N_17061);
xor U18313 (N_18313,N_16403,N_17405);
and U18314 (N_18314,N_16487,N_17058);
or U18315 (N_18315,N_16581,N_16157);
nor U18316 (N_18316,N_17160,N_16297);
xnor U18317 (N_18317,N_17065,N_17443);
xnor U18318 (N_18318,N_17938,N_17627);
nor U18319 (N_18319,N_17556,N_16159);
and U18320 (N_18320,N_16233,N_17817);
xnor U18321 (N_18321,N_17391,N_17522);
nor U18322 (N_18322,N_17139,N_17720);
nand U18323 (N_18323,N_17261,N_16534);
xnor U18324 (N_18324,N_17709,N_16230);
or U18325 (N_18325,N_16780,N_16419);
xor U18326 (N_18326,N_16907,N_16470);
and U18327 (N_18327,N_17355,N_16499);
xor U18328 (N_18328,N_16277,N_16424);
nor U18329 (N_18329,N_16690,N_17581);
xnor U18330 (N_18330,N_17045,N_17144);
nor U18331 (N_18331,N_16018,N_16833);
xor U18332 (N_18332,N_16010,N_17802);
nand U18333 (N_18333,N_17312,N_17387);
nor U18334 (N_18334,N_16554,N_17264);
and U18335 (N_18335,N_16785,N_16917);
nor U18336 (N_18336,N_16577,N_16664);
xor U18337 (N_18337,N_16851,N_17265);
xor U18338 (N_18338,N_16137,N_16529);
nand U18339 (N_18339,N_17269,N_16441);
or U18340 (N_18340,N_17087,N_17917);
xnor U18341 (N_18341,N_16997,N_17249);
nor U18342 (N_18342,N_16491,N_16928);
and U18343 (N_18343,N_17350,N_17510);
nor U18344 (N_18344,N_16748,N_17472);
nand U18345 (N_18345,N_17191,N_16136);
nand U18346 (N_18346,N_16895,N_16107);
nor U18347 (N_18347,N_16149,N_17299);
xor U18348 (N_18348,N_16559,N_16992);
xor U18349 (N_18349,N_17131,N_17394);
xor U18350 (N_18350,N_16027,N_16395);
xor U18351 (N_18351,N_17845,N_17303);
nor U18352 (N_18352,N_16867,N_17728);
or U18353 (N_18353,N_17807,N_17063);
nor U18354 (N_18354,N_17118,N_16270);
xor U18355 (N_18355,N_17344,N_17692);
and U18356 (N_18356,N_17186,N_17883);
or U18357 (N_18357,N_16197,N_17842);
nor U18358 (N_18358,N_16767,N_16586);
or U18359 (N_18359,N_16740,N_16600);
or U18360 (N_18360,N_16285,N_17697);
nand U18361 (N_18361,N_17771,N_16380);
and U18362 (N_18362,N_17257,N_17349);
xnor U18363 (N_18363,N_17112,N_17124);
nand U18364 (N_18364,N_17841,N_17080);
or U18365 (N_18365,N_17565,N_17263);
and U18366 (N_18366,N_17752,N_17501);
nor U18367 (N_18367,N_16435,N_17481);
nand U18368 (N_18368,N_17758,N_17230);
or U18369 (N_18369,N_17279,N_17774);
nor U18370 (N_18370,N_17583,N_16206);
or U18371 (N_18371,N_17159,N_17503);
nand U18372 (N_18372,N_16810,N_17965);
xor U18373 (N_18373,N_17235,N_17205);
nor U18374 (N_18374,N_17716,N_16370);
and U18375 (N_18375,N_17031,N_17695);
and U18376 (N_18376,N_17507,N_16649);
xnor U18377 (N_18377,N_17474,N_16469);
and U18378 (N_18378,N_17702,N_17527);
and U18379 (N_18379,N_17939,N_16111);
nand U18380 (N_18380,N_17498,N_16221);
nand U18381 (N_18381,N_17610,N_16930);
nand U18382 (N_18382,N_17580,N_17366);
or U18383 (N_18383,N_16004,N_17636);
xor U18384 (N_18384,N_16766,N_17597);
xnor U18385 (N_18385,N_17753,N_16635);
or U18386 (N_18386,N_16335,N_16142);
xor U18387 (N_18387,N_16174,N_16076);
nor U18388 (N_18388,N_17256,N_16318);
xnor U18389 (N_18389,N_17834,N_16227);
nand U18390 (N_18390,N_16163,N_16967);
nand U18391 (N_18391,N_17993,N_17095);
nor U18392 (N_18392,N_17738,N_17262);
xor U18393 (N_18393,N_16406,N_16103);
or U18394 (N_18394,N_17870,N_16585);
and U18395 (N_18395,N_16862,N_16402);
nand U18396 (N_18396,N_16127,N_16288);
or U18397 (N_18397,N_17812,N_16031);
xor U18398 (N_18398,N_16325,N_16222);
or U18399 (N_18399,N_16888,N_17388);
or U18400 (N_18400,N_16220,N_16711);
and U18401 (N_18401,N_17445,N_17440);
and U18402 (N_18402,N_17534,N_17687);
nor U18403 (N_18403,N_17547,N_16352);
or U18404 (N_18404,N_16705,N_17596);
nor U18405 (N_18405,N_17223,N_16121);
or U18406 (N_18406,N_16794,N_16390);
nor U18407 (N_18407,N_17295,N_16367);
and U18408 (N_18408,N_17266,N_17180);
or U18409 (N_18409,N_17611,N_17352);
and U18410 (N_18410,N_16328,N_17746);
or U18411 (N_18411,N_17479,N_17512);
nor U18412 (N_18412,N_16831,N_17784);
nor U18413 (N_18413,N_17995,N_17806);
and U18414 (N_18414,N_17763,N_17357);
or U18415 (N_18415,N_16410,N_17625);
nor U18416 (N_18416,N_17157,N_17972);
nor U18417 (N_18417,N_16885,N_17958);
nor U18418 (N_18418,N_16110,N_16882);
xnor U18419 (N_18419,N_17220,N_17648);
or U18420 (N_18420,N_16461,N_16749);
and U18421 (N_18421,N_16440,N_16186);
nand U18422 (N_18422,N_17495,N_16211);
nor U18423 (N_18423,N_17172,N_17833);
and U18424 (N_18424,N_16601,N_17587);
or U18425 (N_18425,N_17595,N_17258);
xnor U18426 (N_18426,N_17014,N_16595);
or U18427 (N_18427,N_16680,N_16761);
nor U18428 (N_18428,N_16527,N_17936);
and U18429 (N_18429,N_16922,N_17107);
xnor U18430 (N_18430,N_17336,N_17890);
nand U18431 (N_18431,N_16804,N_16209);
or U18432 (N_18432,N_16983,N_17290);
nor U18433 (N_18433,N_16266,N_16788);
nor U18434 (N_18434,N_16519,N_17327);
nor U18435 (N_18435,N_16253,N_17111);
nand U18436 (N_18436,N_17345,N_16837);
or U18437 (N_18437,N_16413,N_16399);
nand U18438 (N_18438,N_17189,N_17974);
and U18439 (N_18439,N_17438,N_16605);
or U18440 (N_18440,N_16853,N_17064);
and U18441 (N_18441,N_16478,N_17734);
xor U18442 (N_18442,N_16927,N_16696);
or U18443 (N_18443,N_16152,N_17482);
nand U18444 (N_18444,N_16060,N_16772);
and U18445 (N_18445,N_16348,N_16356);
or U18446 (N_18446,N_16032,N_16117);
and U18447 (N_18447,N_16576,N_16723);
and U18448 (N_18448,N_17386,N_17904);
nor U18449 (N_18449,N_16779,N_17318);
or U18450 (N_18450,N_17671,N_16909);
nand U18451 (N_18451,N_17944,N_16953);
or U18452 (N_18452,N_17858,N_17644);
nand U18453 (N_18453,N_16450,N_17564);
xor U18454 (N_18454,N_17271,N_17846);
xnor U18455 (N_18455,N_16305,N_17799);
and U18456 (N_18456,N_17167,N_16427);
or U18457 (N_18457,N_17641,N_17919);
xor U18458 (N_18458,N_16667,N_16327);
nor U18459 (N_18459,N_16998,N_17012);
xor U18460 (N_18460,N_16373,N_16363);
or U18461 (N_18461,N_16372,N_16062);
nor U18462 (N_18462,N_17770,N_16692);
or U18463 (N_18463,N_17255,N_17286);
nor U18464 (N_18464,N_16481,N_17067);
xnor U18465 (N_18465,N_17985,N_16977);
nor U18466 (N_18466,N_16116,N_17411);
nor U18467 (N_18467,N_16488,N_16090);
nor U18468 (N_18468,N_17537,N_16666);
xnor U18469 (N_18469,N_17589,N_16976);
or U18470 (N_18470,N_16507,N_17722);
nand U18471 (N_18471,N_16622,N_16339);
nand U18472 (N_18472,N_17712,N_17689);
and U18473 (N_18473,N_17562,N_17810);
nor U18474 (N_18474,N_16679,N_17924);
xnor U18475 (N_18475,N_17077,N_17616);
or U18476 (N_18476,N_16291,N_16038);
and U18477 (N_18477,N_16252,N_17046);
or U18478 (N_18478,N_16758,N_17125);
xnor U18479 (N_18479,N_17086,N_17070);
xnor U18480 (N_18480,N_17735,N_16345);
or U18481 (N_18481,N_17135,N_16962);
nand U18482 (N_18482,N_17268,N_17108);
nand U18483 (N_18483,N_16857,N_17401);
nor U18484 (N_18484,N_17134,N_16484);
nand U18485 (N_18485,N_16860,N_17244);
nor U18486 (N_18486,N_17123,N_16330);
nor U18487 (N_18487,N_16052,N_17392);
nor U18488 (N_18488,N_16418,N_16432);
nand U18489 (N_18489,N_17851,N_16707);
nor U18490 (N_18490,N_17777,N_17786);
nand U18491 (N_18491,N_17466,N_17308);
nand U18492 (N_18492,N_16434,N_17281);
and U18493 (N_18493,N_16284,N_17140);
nor U18494 (N_18494,N_16119,N_17896);
or U18495 (N_18495,N_17284,N_17342);
and U18496 (N_18496,N_16508,N_17036);
nor U18497 (N_18497,N_17793,N_16947);
and U18498 (N_18498,N_17068,N_17907);
nor U18499 (N_18499,N_17615,N_17910);
nor U18500 (N_18500,N_17782,N_16278);
or U18501 (N_18501,N_17199,N_17193);
and U18502 (N_18502,N_16687,N_17980);
xnor U18503 (N_18503,N_17676,N_16899);
or U18504 (N_18504,N_16192,N_17748);
nand U18505 (N_18505,N_17836,N_16590);
and U18506 (N_18506,N_16546,N_17768);
nand U18507 (N_18507,N_16839,N_17569);
nor U18508 (N_18508,N_17246,N_16171);
and U18509 (N_18509,N_17961,N_16544);
xor U18510 (N_18510,N_17339,N_17788);
and U18511 (N_18511,N_16164,N_16866);
or U18512 (N_18512,N_17694,N_17946);
nor U18513 (N_18513,N_16485,N_16678);
and U18514 (N_18514,N_17945,N_17458);
nand U18515 (N_18515,N_17960,N_16412);
nand U18516 (N_18516,N_16494,N_17740);
nand U18517 (N_18517,N_16545,N_17196);
and U18518 (N_18518,N_17548,N_16086);
nand U18519 (N_18519,N_17379,N_17765);
and U18520 (N_18520,N_16746,N_17529);
xor U18521 (N_18521,N_16777,N_16362);
nand U18522 (N_18522,N_16466,N_16204);
and U18523 (N_18523,N_16109,N_16388);
and U18524 (N_18524,N_17819,N_16694);
and U18525 (N_18525,N_17714,N_16850);
and U18526 (N_18526,N_16896,N_16592);
nor U18527 (N_18527,N_17213,N_16525);
and U18528 (N_18528,N_17060,N_17981);
nand U18529 (N_18529,N_16988,N_16202);
nor U18530 (N_18530,N_17736,N_17099);
xor U18531 (N_18531,N_16065,N_16183);
nor U18532 (N_18532,N_17152,N_17903);
and U18533 (N_18533,N_17811,N_17377);
and U18534 (N_18534,N_17389,N_16447);
and U18535 (N_18535,N_16124,N_16512);
or U18536 (N_18536,N_17234,N_16258);
nor U18537 (N_18537,N_17142,N_16486);
nand U18538 (N_18538,N_17376,N_17566);
and U18539 (N_18539,N_16347,N_17183);
nand U18540 (N_18540,N_16675,N_16322);
or U18541 (N_18541,N_16684,N_17650);
or U18542 (N_18542,N_16695,N_16884);
xor U18543 (N_18543,N_16869,N_16168);
and U18544 (N_18544,N_16179,N_16620);
or U18545 (N_18545,N_16582,N_16530);
and U18546 (N_18546,N_17998,N_16730);
and U18547 (N_18547,N_17426,N_16941);
and U18548 (N_18548,N_17997,N_17839);
or U18549 (N_18549,N_17019,N_16836);
nor U18550 (N_18550,N_17975,N_17000);
and U18551 (N_18551,N_16520,N_17453);
nor U18552 (N_18552,N_17039,N_16626);
nor U18553 (N_18553,N_16089,N_16185);
nor U18554 (N_18554,N_16787,N_17488);
or U18555 (N_18555,N_16989,N_17240);
nand U18556 (N_18556,N_16378,N_16879);
and U18557 (N_18557,N_16396,N_16555);
nand U18558 (N_18558,N_16543,N_16016);
and U18559 (N_18559,N_16493,N_16811);
xor U18560 (N_18560,N_17451,N_17563);
nand U18561 (N_18561,N_16154,N_17642);
xor U18562 (N_18562,N_17452,N_17248);
and U18563 (N_18563,N_16704,N_17165);
xnor U18564 (N_18564,N_16589,N_16257);
and U18565 (N_18565,N_16580,N_17899);
xnor U18566 (N_18566,N_17837,N_17808);
nor U18567 (N_18567,N_16876,N_17827);
nand U18568 (N_18568,N_16357,N_16856);
and U18569 (N_18569,N_16861,N_16156);
nand U18570 (N_18570,N_16101,N_16351);
and U18571 (N_18571,N_16082,N_17298);
or U18572 (N_18572,N_17048,N_16120);
and U18573 (N_18573,N_16561,N_17682);
or U18574 (N_18574,N_17371,N_16498);
and U18575 (N_18575,N_17651,N_16140);
and U18576 (N_18576,N_17150,N_16658);
nor U18577 (N_18577,N_16574,N_17923);
and U18578 (N_18578,N_17979,N_17162);
nand U18579 (N_18579,N_16229,N_17042);
or U18580 (N_18580,N_17542,N_16138);
nor U18581 (N_18581,N_16832,N_16177);
xor U18582 (N_18582,N_16039,N_16219);
and U18583 (N_18583,N_16059,N_17829);
xnor U18584 (N_18584,N_17491,N_17994);
nand U18585 (N_18585,N_16017,N_16645);
xnor U18586 (N_18586,N_16371,N_17680);
and U18587 (N_18587,N_16558,N_16037);
nand U18588 (N_18588,N_17719,N_16319);
xnor U18589 (N_18589,N_17929,N_17390);
xor U18590 (N_18590,N_17053,N_17730);
xor U18591 (N_18591,N_17865,N_17855);
or U18592 (N_18592,N_17013,N_16077);
nor U18593 (N_18593,N_17551,N_17713);
nor U18594 (N_18594,N_17422,N_17755);
xnor U18595 (N_18595,N_17593,N_16718);
or U18596 (N_18596,N_17075,N_17324);
xnor U18597 (N_18597,N_17599,N_17294);
or U18598 (N_18598,N_17343,N_17034);
and U18599 (N_18599,N_16482,N_16260);
or U18600 (N_18600,N_16654,N_17681);
and U18601 (N_18601,N_17335,N_16063);
xor U18602 (N_18602,N_16439,N_16651);
nand U18603 (N_18603,N_17404,N_16955);
and U18604 (N_18604,N_17210,N_16232);
nand U18605 (N_18605,N_17420,N_17854);
and U18606 (N_18606,N_16564,N_17442);
and U18607 (N_18607,N_17631,N_17416);
and U18608 (N_18608,N_16759,N_16078);
nand U18609 (N_18609,N_16007,N_16296);
nor U18610 (N_18610,N_17555,N_17185);
or U18611 (N_18611,N_17701,N_16148);
or U18612 (N_18612,N_17959,N_16134);
nand U18613 (N_18613,N_17332,N_16624);
xor U18614 (N_18614,N_17102,N_16870);
and U18615 (N_18615,N_17996,N_17809);
nor U18616 (N_18616,N_16669,N_16894);
or U18617 (N_18617,N_17798,N_16240);
xor U18618 (N_18618,N_17634,N_16003);
nor U18619 (N_18619,N_17543,N_16816);
xnor U18620 (N_18620,N_17933,N_16683);
xnor U18621 (N_18621,N_16178,N_17363);
and U18622 (N_18622,N_16337,N_16391);
xnor U18623 (N_18623,N_17900,N_16074);
and U18624 (N_18624,N_17052,N_17873);
and U18625 (N_18625,N_17079,N_17429);
or U18626 (N_18626,N_17146,N_16999);
or U18627 (N_18627,N_16093,N_17605);
nor U18628 (N_18628,N_16877,N_16791);
or U18629 (N_18629,N_16072,N_17603);
or U18630 (N_18630,N_17302,N_16311);
nand U18631 (N_18631,N_17567,N_16950);
nand U18632 (N_18632,N_16286,N_17760);
xnor U18633 (N_18633,N_16887,N_17358);
or U18634 (N_18634,N_16886,N_16170);
and U18635 (N_18635,N_16921,N_16934);
nand U18636 (N_18636,N_16276,N_16778);
and U18637 (N_18637,N_16020,N_16903);
xor U18638 (N_18638,N_16128,N_16712);
nor U18639 (N_18639,N_16910,N_16548);
xnor U18640 (N_18640,N_16611,N_17513);
nand U18641 (N_18641,N_16889,N_17493);
and U18642 (N_18642,N_16803,N_16005);
nand U18643 (N_18643,N_17672,N_17761);
nor U18644 (N_18644,N_16073,N_16625);
xor U18645 (N_18645,N_17285,N_17882);
or U18646 (N_18646,N_17820,N_17601);
nand U18647 (N_18647,N_17989,N_16006);
or U18648 (N_18648,N_17549,N_17049);
xor U18649 (N_18649,N_17280,N_17622);
nor U18650 (N_18650,N_16451,N_16224);
xnor U18651 (N_18651,N_16822,N_16167);
nor U18652 (N_18652,N_16268,N_16034);
nor U18653 (N_18653,N_16956,N_16916);
nor U18654 (N_18654,N_16083,N_17916);
xnor U18655 (N_18655,N_16182,N_16516);
or U18656 (N_18656,N_16141,N_17242);
xor U18657 (N_18657,N_16022,N_17545);
nand U18658 (N_18658,N_17202,N_17977);
and U18659 (N_18659,N_17119,N_16147);
xor U18660 (N_18660,N_17151,N_17791);
nor U18661 (N_18661,N_17927,N_17953);
nor U18662 (N_18662,N_16289,N_16805);
and U18663 (N_18663,N_17113,N_17362);
nor U18664 (N_18664,N_17085,N_16783);
or U18665 (N_18665,N_17221,N_17999);
or U18666 (N_18666,N_16398,N_17492);
and U18667 (N_18667,N_17898,N_17559);
and U18668 (N_18668,N_17824,N_17041);
nor U18669 (N_18669,N_17624,N_16474);
and U18670 (N_18670,N_16438,N_16568);
nor U18671 (N_18671,N_17950,N_17745);
xor U18672 (N_18672,N_17943,N_16374);
nand U18673 (N_18673,N_17454,N_17523);
and U18674 (N_18674,N_16428,N_16280);
nor U18675 (N_18675,N_17462,N_16693);
xnor U18676 (N_18676,N_16506,N_16235);
or U18677 (N_18677,N_16150,N_17115);
nand U18678 (N_18678,N_16437,N_17001);
xor U18679 (N_18679,N_16655,N_17540);
nor U18680 (N_18680,N_17840,N_17921);
nand U18681 (N_18681,N_17021,N_17455);
nand U18682 (N_18682,N_17707,N_17607);
nand U18683 (N_18683,N_16949,N_16524);
and U18684 (N_18684,N_17699,N_16897);
or U18685 (N_18685,N_16905,N_17779);
or U18686 (N_18686,N_16706,N_17023);
xnor U18687 (N_18687,N_16798,N_16951);
nor U18688 (N_18688,N_16446,N_17499);
nand U18689 (N_18689,N_17330,N_17956);
or U18690 (N_18690,N_17477,N_17775);
nand U18691 (N_18691,N_17769,N_16971);
and U18692 (N_18692,N_17708,N_16931);
or U18693 (N_18693,N_17326,N_17657);
nor U18694 (N_18694,N_17667,N_16389);
xnor U18695 (N_18695,N_16026,N_17169);
nor U18696 (N_18696,N_16727,N_17154);
and U18697 (N_18697,N_16604,N_17984);
nand U18698 (N_18698,N_17164,N_17132);
nor U18699 (N_18699,N_17664,N_17623);
xor U18700 (N_18700,N_16153,N_17228);
xor U18701 (N_18701,N_16919,N_17940);
nand U18702 (N_18702,N_17035,N_16271);
nand U18703 (N_18703,N_17772,N_17143);
xnor U18704 (N_18704,N_17717,N_16668);
nor U18705 (N_18705,N_16024,N_16789);
xor U18706 (N_18706,N_17516,N_16194);
xnor U18707 (N_18707,N_16904,N_16313);
or U18708 (N_18708,N_16774,N_16631);
nand U18709 (N_18709,N_16702,N_17902);
and U18710 (N_18710,N_17004,N_16960);
nor U18711 (N_18711,N_17329,N_16044);
and U18712 (N_18712,N_16261,N_17818);
or U18713 (N_18713,N_17020,N_17822);
nand U18714 (N_18714,N_17480,N_17852);
nor U18715 (N_18715,N_16933,N_17592);
or U18716 (N_18716,N_17659,N_16911);
or U18717 (N_18717,N_16878,N_16621);
nand U18718 (N_18718,N_17319,N_17155);
xor U18719 (N_18719,N_17457,N_17382);
xnor U18720 (N_18720,N_16165,N_17178);
and U18721 (N_18721,N_16557,N_16957);
xnor U18722 (N_18722,N_16537,N_17338);
nor U18723 (N_18723,N_16379,N_16729);
nor U18724 (N_18724,N_17050,N_16079);
nand U18725 (N_18725,N_17721,N_16358);
nand U18726 (N_18726,N_17029,N_16898);
nor U18727 (N_18727,N_16279,N_17578);
nor U18728 (N_18728,N_17054,N_17369);
xor U18729 (N_18729,N_17639,N_16575);
or U18730 (N_18730,N_16112,N_16963);
and U18731 (N_18731,N_17270,N_16483);
or U18732 (N_18732,N_16883,N_17517);
xor U18733 (N_18733,N_16926,N_16646);
nor U18734 (N_18734,N_16912,N_16236);
nor U18735 (N_18735,N_16108,N_16365);
nor U18736 (N_18736,N_16146,N_17638);
or U18737 (N_18737,N_17434,N_17602);
and U18738 (N_18738,N_16259,N_16618);
or U18739 (N_18739,N_16952,N_16201);
and U18740 (N_18740,N_16098,N_17520);
xnor U18741 (N_18741,N_17831,N_16722);
nand U18742 (N_18742,N_16249,N_17287);
nor U18743 (N_18743,N_16510,N_16199);
and U18744 (N_18744,N_16986,N_16196);
or U18745 (N_18745,N_17912,N_17647);
nand U18746 (N_18746,N_16061,N_16728);
xor U18747 (N_18747,N_17003,N_17915);
nand U18748 (N_18748,N_17553,N_17497);
or U18749 (N_18749,N_17098,N_17686);
nor U18750 (N_18750,N_17561,N_16001);
xnor U18751 (N_18751,N_16731,N_17278);
nor U18752 (N_18752,N_17778,N_17059);
or U18753 (N_18753,N_16191,N_16844);
or U18754 (N_18754,N_16293,N_17875);
xor U18755 (N_18755,N_17253,N_16070);
or U18756 (N_18756,N_16104,N_16868);
nor U18757 (N_18757,N_17460,N_16299);
or U18758 (N_18758,N_17374,N_17365);
nor U18759 (N_18759,N_17092,N_17027);
and U18760 (N_18760,N_16028,N_16047);
xor U18761 (N_18761,N_17604,N_16444);
nand U18762 (N_18762,N_17227,N_17914);
nor U18763 (N_18763,N_16012,N_16753);
nor U18764 (N_18764,N_16503,N_16349);
and U18765 (N_18765,N_16929,N_17880);
nand U18766 (N_18766,N_16809,N_17679);
or U18767 (N_18767,N_16422,N_16055);
or U18768 (N_18768,N_17814,N_16361);
and U18769 (N_18769,N_16768,N_17813);
nor U18770 (N_18770,N_16556,N_16578);
nand U18771 (N_18771,N_16762,N_17367);
xor U18772 (N_18772,N_16824,N_16504);
nand U18773 (N_18773,N_16641,N_17613);
or U18774 (N_18774,N_16755,N_16173);
xnor U18775 (N_18775,N_16985,N_17166);
and U18776 (N_18776,N_17724,N_16464);
and U18777 (N_18777,N_16603,N_17539);
xnor U18778 (N_18778,N_16460,N_16859);
nand U18779 (N_18779,N_16650,N_17009);
or U18780 (N_18780,N_17869,N_17877);
or U18781 (N_18781,N_17982,N_16775);
nand U18782 (N_18782,N_17888,N_16225);
xnor U18783 (N_18783,N_17282,N_17084);
nand U18784 (N_18784,N_17757,N_17173);
nand U18785 (N_18785,N_17093,N_16736);
or U18786 (N_18786,N_17691,N_16502);
nand U18787 (N_18787,N_16473,N_17370);
or U18788 (N_18788,N_17913,N_16263);
and U18789 (N_18789,N_16745,N_16854);
nor U18790 (N_18790,N_16801,N_17407);
nor U18791 (N_18791,N_16835,N_17226);
nor U18792 (N_18792,N_17204,N_16596);
and U18793 (N_18793,N_16255,N_16562);
or U18794 (N_18794,N_16454,N_17949);
nor U18795 (N_18795,N_17309,N_17328);
or U18796 (N_18796,N_16195,N_16764);
xor U18797 (N_18797,N_16226,N_16080);
and U18798 (N_18798,N_17823,N_16511);
nor U18799 (N_18799,N_17120,N_17449);
or U18800 (N_18800,N_16915,N_17484);
nand U18801 (N_18801,N_17274,N_16993);
nor U18802 (N_18802,N_16978,N_17585);
nand U18803 (N_18803,N_16354,N_17600);
xor U18804 (N_18804,N_16523,N_16223);
nand U18805 (N_18805,N_16737,N_16771);
nor U18806 (N_18806,N_17419,N_17732);
nor U18807 (N_18807,N_17496,N_16214);
nand U18808 (N_18808,N_16522,N_17219);
and U18809 (N_18809,N_17127,N_17608);
xor U18810 (N_18810,N_16084,N_17987);
nand U18811 (N_18811,N_17653,N_16126);
xor U18812 (N_18812,N_17476,N_16315);
nor U18813 (N_18813,N_17797,N_16274);
nand U18814 (N_18814,N_16954,N_17937);
nand U18815 (N_18815,N_16721,N_16462);
xor U18816 (N_18816,N_16688,N_16738);
and U18817 (N_18817,N_16091,N_17241);
xnor U18818 (N_18818,N_17577,N_17423);
and U18819 (N_18819,N_17104,N_16049);
nand U18820 (N_18820,N_17619,N_16262);
xor U18821 (N_18821,N_16968,N_16172);
xnor U18822 (N_18822,N_16614,N_17859);
nand U18823 (N_18823,N_16979,N_17206);
xor U18824 (N_18824,N_16633,N_16155);
nor U18825 (N_18825,N_16663,N_17901);
xor U18826 (N_18826,N_17106,N_16409);
xnor U18827 (N_18827,N_16475,N_17259);
and U18828 (N_18828,N_16591,N_16918);
nand U18829 (N_18829,N_17337,N_16743);
nand U18830 (N_18830,N_16818,N_16189);
and U18831 (N_18831,N_17582,N_16489);
and U18832 (N_18832,N_16205,N_16264);
nand U18833 (N_18833,N_16500,N_16634);
xnor U18834 (N_18834,N_16965,N_17887);
or U18835 (N_18835,N_17138,N_16940);
xor U18836 (N_18836,N_17723,N_17528);
xor U18837 (N_18837,N_16944,N_17430);
nor U18838 (N_18838,N_17895,N_17886);
nor U18839 (N_18839,N_16326,N_17931);
nor U18840 (N_18840,N_17665,N_16448);
nor U18841 (N_18841,N_17243,N_16000);
and U18842 (N_18842,N_16893,N_16099);
or U18843 (N_18843,N_16735,N_16838);
and U18844 (N_18844,N_16739,N_17505);
xnor U18845 (N_18845,N_17978,N_16864);
nor U18846 (N_18846,N_16294,N_16638);
and U18847 (N_18847,N_17275,N_16732);
xor U18848 (N_18848,N_17892,N_16056);
nand U18849 (N_18849,N_17334,N_17372);
nand U18850 (N_18850,N_17433,N_17731);
xor U18851 (N_18851,N_16563,N_16340);
nand U18852 (N_18852,N_17885,N_17663);
nor U18853 (N_18853,N_16708,N_16892);
nor U18854 (N_18854,N_16750,N_17096);
and U18855 (N_18855,N_17402,N_17408);
xnor U18856 (N_18856,N_16873,N_16914);
xor U18857 (N_18857,N_16938,N_17670);
nor U18858 (N_18858,N_17789,N_17626);
nor U18859 (N_18859,N_17436,N_16405);
and U18860 (N_18860,N_17101,N_16431);
nand U18861 (N_18861,N_16401,N_16653);
nor U18862 (N_18862,N_16269,N_17217);
and U18863 (N_18863,N_17238,N_16449);
xnor U18864 (N_18864,N_17211,N_16765);
nor U18865 (N_18865,N_16272,N_16572);
xnor U18866 (N_18866,N_16251,N_16281);
xnor U18867 (N_18867,N_16404,N_16139);
nand U18868 (N_18868,N_17368,N_17373);
xnor U18869 (N_18869,N_16521,N_17586);
xor U18870 (N_18870,N_17141,N_17317);
nor U18871 (N_18871,N_17969,N_17879);
or U18872 (N_18872,N_17182,N_17467);
or U18873 (N_18873,N_16458,N_17464);
nor U18874 (N_18874,N_17456,N_17727);
nand U18875 (N_18875,N_16871,N_17446);
nor U18876 (N_18876,N_17568,N_17704);
nor U18877 (N_18877,N_17519,N_17057);
and U18878 (N_18878,N_16817,N_17864);
and U18879 (N_18879,N_17032,N_17435);
xnor U18880 (N_18880,N_17171,N_17685);
and U18881 (N_18881,N_17661,N_16471);
xor U18882 (N_18882,N_17815,N_17088);
or U18883 (N_18883,N_17872,N_16421);
xnor U18884 (N_18884,N_16643,N_17396);
nor U18885 (N_18885,N_17181,N_17010);
nor U18886 (N_18886,N_17301,N_17541);
or U18887 (N_18887,N_16671,N_17518);
and U18888 (N_18888,N_16612,N_17198);
nor U18889 (N_18889,N_16714,N_16820);
or U18890 (N_18890,N_17441,N_17153);
nor U18891 (N_18891,N_16754,N_17040);
xor U18892 (N_18892,N_16660,N_17475);
nor U18893 (N_18893,N_17174,N_17489);
and U18894 (N_18894,N_17056,N_16023);
or U18895 (N_18895,N_17122,N_16541);
nor U18896 (N_18896,N_17743,N_16584);
or U18897 (N_18897,N_16479,N_16187);
nor U18898 (N_18898,N_17874,N_16457);
nand U18899 (N_18899,N_17947,N_16014);
nand U18900 (N_18900,N_16670,N_17759);
xnor U18901 (N_18901,N_17380,N_16467);
nand U18902 (N_18902,N_17232,N_16973);
and U18903 (N_18903,N_16248,N_17017);
and U18904 (N_18904,N_16719,N_17606);
xnor U18905 (N_18905,N_16720,N_17684);
or U18906 (N_18906,N_16169,N_17573);
xor U18907 (N_18907,N_17660,N_17703);
nor U18908 (N_18908,N_16550,N_17254);
xor U18909 (N_18909,N_17683,N_17313);
and U18910 (N_18910,N_16030,N_17876);
nand U18911 (N_18911,N_17751,N_17293);
nand U18912 (N_18912,N_17209,N_16135);
or U18913 (N_18913,N_17225,N_16131);
nor U18914 (N_18914,N_17078,N_16786);
nor U18915 (N_18915,N_17486,N_17208);
nor U18916 (N_18916,N_16875,N_16132);
or U18917 (N_18917,N_17934,N_16874);
or U18918 (N_18918,N_17089,N_16609);
nand U18919 (N_18919,N_16290,N_16320);
nor U18920 (N_18920,N_16513,N_16321);
nor U18921 (N_18921,N_16385,N_16430);
and U18922 (N_18922,N_17925,N_16526);
nand U18923 (N_18923,N_16629,N_16594);
nand U18924 (N_18924,N_17378,N_17988);
nor U18925 (N_18925,N_16539,N_17986);
and U18926 (N_18926,N_17383,N_16231);
or U18927 (N_18927,N_17168,N_17957);
and U18928 (N_18928,N_17364,N_17710);
xor U18929 (N_18929,N_16472,N_16324);
xor U18930 (N_18930,N_16659,N_17037);
or U18931 (N_18931,N_16036,N_17990);
xor U18932 (N_18932,N_16058,N_17231);
and U18933 (N_18933,N_17291,N_16254);
nor U18934 (N_18934,N_17351,N_16392);
or U18935 (N_18935,N_17932,N_17973);
or U18936 (N_18936,N_17550,N_16443);
and U18937 (N_18937,N_16243,N_17033);
nand U18938 (N_18938,N_17669,N_17629);
xnor U18939 (N_18939,N_16685,N_17272);
or U18940 (N_18940,N_17725,N_17655);
nor U18941 (N_18941,N_16102,N_16505);
nor U18942 (N_18942,N_16812,N_17297);
and U18943 (N_18943,N_16834,N_16686);
nand U18944 (N_18944,N_16827,N_17136);
nor U18945 (N_18945,N_16359,N_17314);
and U18946 (N_18946,N_16298,N_16247);
and U18947 (N_18947,N_16815,N_16377);
nor U18948 (N_18948,N_16741,N_16292);
or U18949 (N_18949,N_17662,N_17007);
or U18950 (N_18950,N_16384,N_17968);
nand U18951 (N_18951,N_16468,N_17652);
and U18952 (N_18952,N_16964,N_16453);
nor U18953 (N_18953,N_16792,N_17715);
nand U18954 (N_18954,N_16015,N_17557);
nand U18955 (N_18955,N_17490,N_17930);
nand U18956 (N_18956,N_16632,N_17948);
nand U18957 (N_18957,N_17675,N_16994);
nand U18958 (N_18958,N_17215,N_17963);
xnor U18959 (N_18959,N_16088,N_16317);
nor U18960 (N_18960,N_16533,N_17361);
nor U18961 (N_18961,N_16087,N_16781);
nand U18962 (N_18962,N_17991,N_16334);
xnor U18963 (N_18963,N_17571,N_17431);
nand U18964 (N_18964,N_17525,N_16845);
or U18965 (N_18965,N_17952,N_16733);
nand U18966 (N_18966,N_17821,N_17825);
xor U18967 (N_18967,N_16408,N_16175);
nand U18968 (N_18968,N_17043,N_17069);
nand U18969 (N_18969,N_17207,N_16332);
nor U18970 (N_18970,N_16672,N_16808);
and U18971 (N_18971,N_17756,N_16717);
or U18972 (N_18972,N_16316,N_17835);
xor U18973 (N_18973,N_16970,N_16509);
and U18974 (N_18974,N_16203,N_16536);
nand U18975 (N_18975,N_17283,N_17044);
nand U18976 (N_18976,N_16300,N_16048);
xor U18977 (N_18977,N_17967,N_16588);
nor U18978 (N_18978,N_16636,N_17385);
nand U18979 (N_18979,N_16411,N_17828);
xnor U18980 (N_18980,N_17245,N_16920);
nand U18981 (N_18981,N_16456,N_17804);
xnor U18982 (N_18982,N_16936,N_16118);
and U18983 (N_18983,N_16770,N_17643);
nor U18984 (N_18984,N_16193,N_16161);
nand U18985 (N_18985,N_16639,N_17011);
and U18986 (N_18986,N_17538,N_16021);
nor U18987 (N_18987,N_16009,N_16465);
or U18988 (N_18988,N_16760,N_16982);
or U18989 (N_18989,N_16234,N_16991);
nand U18990 (N_18990,N_17273,N_16616);
and U18991 (N_18991,N_17718,N_16160);
and U18992 (N_18992,N_17658,N_17236);
and U18993 (N_18993,N_17195,N_17861);
and U18994 (N_18994,N_16567,N_16990);
nor U18995 (N_18995,N_16881,N_16906);
or U18996 (N_18996,N_16215,N_16532);
xnor U18997 (N_18997,N_16825,N_16217);
xnor U18998 (N_18998,N_16959,N_17201);
and U18999 (N_18999,N_16366,N_16069);
xor U19000 (N_19000,N_17739,N_17937);
xnor U19001 (N_19001,N_16719,N_16302);
and U19002 (N_19002,N_17764,N_17781);
and U19003 (N_19003,N_17801,N_16557);
xnor U19004 (N_19004,N_16258,N_17921);
or U19005 (N_19005,N_17846,N_16734);
nor U19006 (N_19006,N_16708,N_17938);
nor U19007 (N_19007,N_16125,N_17890);
nand U19008 (N_19008,N_16395,N_17416);
nor U19009 (N_19009,N_17843,N_17021);
xor U19010 (N_19010,N_16549,N_17315);
or U19011 (N_19011,N_17387,N_16362);
and U19012 (N_19012,N_17055,N_17353);
and U19013 (N_19013,N_16408,N_17576);
or U19014 (N_19014,N_16120,N_17109);
nand U19015 (N_19015,N_17941,N_17883);
or U19016 (N_19016,N_17293,N_16335);
nand U19017 (N_19017,N_16468,N_16723);
or U19018 (N_19018,N_17562,N_16302);
and U19019 (N_19019,N_16529,N_16316);
or U19020 (N_19020,N_17696,N_16609);
xnor U19021 (N_19021,N_17442,N_16141);
nand U19022 (N_19022,N_17522,N_16359);
xor U19023 (N_19023,N_16024,N_16119);
nand U19024 (N_19024,N_17126,N_16323);
nand U19025 (N_19025,N_17799,N_16431);
or U19026 (N_19026,N_17183,N_17264);
and U19027 (N_19027,N_16528,N_16198);
nor U19028 (N_19028,N_16502,N_16440);
and U19029 (N_19029,N_17179,N_16541);
and U19030 (N_19030,N_16202,N_17058);
nor U19031 (N_19031,N_17682,N_16525);
or U19032 (N_19032,N_16346,N_16272);
or U19033 (N_19033,N_17209,N_17172);
and U19034 (N_19034,N_17358,N_17490);
nor U19035 (N_19035,N_16291,N_16169);
nor U19036 (N_19036,N_16079,N_16348);
xor U19037 (N_19037,N_16099,N_16115);
xor U19038 (N_19038,N_17066,N_17265);
xnor U19039 (N_19039,N_16749,N_17649);
and U19040 (N_19040,N_17490,N_16642);
or U19041 (N_19041,N_16890,N_17997);
nand U19042 (N_19042,N_17980,N_16291);
and U19043 (N_19043,N_16030,N_17441);
and U19044 (N_19044,N_16435,N_16267);
or U19045 (N_19045,N_17973,N_17918);
xor U19046 (N_19046,N_17903,N_17898);
xnor U19047 (N_19047,N_16335,N_17503);
or U19048 (N_19048,N_16142,N_16036);
nor U19049 (N_19049,N_17656,N_16218);
nor U19050 (N_19050,N_17157,N_16992);
xnor U19051 (N_19051,N_16462,N_16502);
or U19052 (N_19052,N_17122,N_17796);
nand U19053 (N_19053,N_16765,N_17277);
or U19054 (N_19054,N_17284,N_17529);
or U19055 (N_19055,N_17603,N_17751);
or U19056 (N_19056,N_16511,N_17435);
or U19057 (N_19057,N_16273,N_16402);
nor U19058 (N_19058,N_17848,N_17308);
and U19059 (N_19059,N_16571,N_17864);
nor U19060 (N_19060,N_16306,N_16956);
or U19061 (N_19061,N_16258,N_17305);
and U19062 (N_19062,N_17743,N_17182);
nor U19063 (N_19063,N_17589,N_17382);
and U19064 (N_19064,N_17842,N_17748);
nand U19065 (N_19065,N_16556,N_17237);
nand U19066 (N_19066,N_16758,N_17957);
nor U19067 (N_19067,N_17910,N_16004);
or U19068 (N_19068,N_16968,N_17716);
nand U19069 (N_19069,N_17180,N_17035);
xnor U19070 (N_19070,N_17418,N_16948);
and U19071 (N_19071,N_16577,N_17915);
nand U19072 (N_19072,N_16068,N_16618);
xor U19073 (N_19073,N_17391,N_16672);
and U19074 (N_19074,N_17375,N_16696);
nand U19075 (N_19075,N_17472,N_17784);
nor U19076 (N_19076,N_16915,N_16633);
xnor U19077 (N_19077,N_16572,N_16635);
nor U19078 (N_19078,N_16188,N_17383);
xnor U19079 (N_19079,N_17113,N_17408);
nor U19080 (N_19080,N_16225,N_17439);
nor U19081 (N_19081,N_17245,N_17158);
nor U19082 (N_19082,N_17085,N_17106);
and U19083 (N_19083,N_16141,N_16431);
or U19084 (N_19084,N_16900,N_16640);
nor U19085 (N_19085,N_17676,N_17276);
nand U19086 (N_19086,N_17451,N_16505);
nand U19087 (N_19087,N_17106,N_17283);
and U19088 (N_19088,N_17080,N_16765);
nor U19089 (N_19089,N_17892,N_17572);
and U19090 (N_19090,N_17996,N_17825);
nor U19091 (N_19091,N_16834,N_16008);
or U19092 (N_19092,N_16932,N_16374);
or U19093 (N_19093,N_17568,N_16008);
or U19094 (N_19094,N_17808,N_16184);
xor U19095 (N_19095,N_16043,N_17339);
nor U19096 (N_19096,N_17609,N_17748);
or U19097 (N_19097,N_17428,N_16769);
xnor U19098 (N_19098,N_17476,N_17139);
or U19099 (N_19099,N_17661,N_16898);
nor U19100 (N_19100,N_16564,N_17832);
nor U19101 (N_19101,N_17242,N_16993);
nor U19102 (N_19102,N_16114,N_17062);
xnor U19103 (N_19103,N_17530,N_16502);
nor U19104 (N_19104,N_17262,N_17329);
or U19105 (N_19105,N_17557,N_17660);
or U19106 (N_19106,N_17519,N_16478);
or U19107 (N_19107,N_17776,N_17667);
nor U19108 (N_19108,N_17114,N_16184);
nand U19109 (N_19109,N_17166,N_17363);
nand U19110 (N_19110,N_17420,N_17058);
nor U19111 (N_19111,N_17920,N_16566);
xor U19112 (N_19112,N_16272,N_16233);
xnor U19113 (N_19113,N_16617,N_17256);
xor U19114 (N_19114,N_16368,N_16016);
xor U19115 (N_19115,N_16127,N_16844);
or U19116 (N_19116,N_17521,N_17317);
and U19117 (N_19117,N_17795,N_17579);
nand U19118 (N_19118,N_17351,N_17551);
xnor U19119 (N_19119,N_17950,N_17288);
or U19120 (N_19120,N_16805,N_16904);
nand U19121 (N_19121,N_16774,N_17187);
and U19122 (N_19122,N_17430,N_17292);
nand U19123 (N_19123,N_17217,N_17004);
nand U19124 (N_19124,N_17387,N_16460);
xor U19125 (N_19125,N_16071,N_17935);
and U19126 (N_19126,N_17285,N_16892);
xnor U19127 (N_19127,N_17684,N_16879);
nor U19128 (N_19128,N_17748,N_16858);
nand U19129 (N_19129,N_16774,N_16816);
or U19130 (N_19130,N_16268,N_17909);
nor U19131 (N_19131,N_16211,N_17765);
or U19132 (N_19132,N_17568,N_16197);
or U19133 (N_19133,N_17260,N_17411);
nand U19134 (N_19134,N_17141,N_16160);
and U19135 (N_19135,N_17887,N_16330);
and U19136 (N_19136,N_16959,N_17144);
nand U19137 (N_19137,N_17913,N_16952);
nor U19138 (N_19138,N_17588,N_17524);
and U19139 (N_19139,N_16780,N_17133);
and U19140 (N_19140,N_16854,N_17910);
nor U19141 (N_19141,N_16353,N_16218);
or U19142 (N_19142,N_16405,N_17384);
and U19143 (N_19143,N_17124,N_16817);
or U19144 (N_19144,N_16321,N_17607);
nand U19145 (N_19145,N_17875,N_16910);
or U19146 (N_19146,N_17978,N_16970);
or U19147 (N_19147,N_17855,N_17885);
xor U19148 (N_19148,N_17892,N_17389);
and U19149 (N_19149,N_16504,N_16707);
or U19150 (N_19150,N_16316,N_17806);
nand U19151 (N_19151,N_17713,N_16456);
or U19152 (N_19152,N_16965,N_17097);
nor U19153 (N_19153,N_16366,N_16149);
xnor U19154 (N_19154,N_17139,N_17589);
nor U19155 (N_19155,N_17805,N_16621);
nor U19156 (N_19156,N_17481,N_17074);
nor U19157 (N_19157,N_17219,N_16599);
or U19158 (N_19158,N_17539,N_16940);
or U19159 (N_19159,N_17848,N_17068);
xnor U19160 (N_19160,N_16662,N_16676);
nor U19161 (N_19161,N_16901,N_17157);
or U19162 (N_19162,N_17960,N_17820);
nor U19163 (N_19163,N_16633,N_17551);
xor U19164 (N_19164,N_17323,N_17051);
xnor U19165 (N_19165,N_17856,N_16373);
nor U19166 (N_19166,N_17886,N_17933);
nand U19167 (N_19167,N_17893,N_17787);
xor U19168 (N_19168,N_17319,N_17805);
or U19169 (N_19169,N_17722,N_16723);
nor U19170 (N_19170,N_16837,N_17455);
xor U19171 (N_19171,N_17773,N_16513);
xnor U19172 (N_19172,N_17011,N_17428);
or U19173 (N_19173,N_17079,N_17684);
and U19174 (N_19174,N_17360,N_16089);
xnor U19175 (N_19175,N_17608,N_17235);
nor U19176 (N_19176,N_17159,N_16994);
and U19177 (N_19177,N_17268,N_16681);
xor U19178 (N_19178,N_16394,N_16891);
nand U19179 (N_19179,N_17301,N_16359);
nand U19180 (N_19180,N_16043,N_17549);
or U19181 (N_19181,N_16211,N_17736);
or U19182 (N_19182,N_17908,N_17512);
or U19183 (N_19183,N_17148,N_17622);
xor U19184 (N_19184,N_17102,N_16181);
nand U19185 (N_19185,N_17407,N_16785);
nor U19186 (N_19186,N_17166,N_16925);
nor U19187 (N_19187,N_16162,N_17923);
nor U19188 (N_19188,N_16047,N_17830);
nand U19189 (N_19189,N_16476,N_16328);
or U19190 (N_19190,N_17112,N_17352);
xor U19191 (N_19191,N_17184,N_17108);
nand U19192 (N_19192,N_16888,N_16267);
or U19193 (N_19193,N_16952,N_16783);
and U19194 (N_19194,N_17008,N_17740);
nor U19195 (N_19195,N_17628,N_16563);
nand U19196 (N_19196,N_16944,N_17030);
xor U19197 (N_19197,N_16200,N_16903);
nand U19198 (N_19198,N_16787,N_16562);
xor U19199 (N_19199,N_16680,N_17762);
nor U19200 (N_19200,N_16044,N_17271);
and U19201 (N_19201,N_16189,N_16575);
nor U19202 (N_19202,N_16499,N_16106);
nor U19203 (N_19203,N_17386,N_17040);
and U19204 (N_19204,N_17995,N_17410);
and U19205 (N_19205,N_16282,N_16618);
nand U19206 (N_19206,N_16764,N_16783);
nor U19207 (N_19207,N_16485,N_17062);
xor U19208 (N_19208,N_17711,N_17570);
nand U19209 (N_19209,N_16140,N_17367);
nand U19210 (N_19210,N_16446,N_17296);
xor U19211 (N_19211,N_17104,N_16517);
and U19212 (N_19212,N_17274,N_17121);
nand U19213 (N_19213,N_16719,N_17438);
and U19214 (N_19214,N_16996,N_17184);
xor U19215 (N_19215,N_17427,N_17000);
xnor U19216 (N_19216,N_16264,N_16890);
nor U19217 (N_19217,N_17557,N_17260);
xor U19218 (N_19218,N_16658,N_17132);
or U19219 (N_19219,N_17098,N_16723);
and U19220 (N_19220,N_17667,N_17116);
or U19221 (N_19221,N_16117,N_17623);
and U19222 (N_19222,N_16385,N_16368);
xnor U19223 (N_19223,N_17251,N_17931);
nor U19224 (N_19224,N_16299,N_17012);
and U19225 (N_19225,N_17471,N_16487);
or U19226 (N_19226,N_17673,N_16098);
or U19227 (N_19227,N_17083,N_17260);
xor U19228 (N_19228,N_16336,N_16220);
nor U19229 (N_19229,N_17118,N_17598);
nor U19230 (N_19230,N_17811,N_16076);
nor U19231 (N_19231,N_17175,N_17689);
nand U19232 (N_19232,N_16284,N_16872);
nor U19233 (N_19233,N_17798,N_16074);
or U19234 (N_19234,N_16561,N_17125);
nor U19235 (N_19235,N_17039,N_16851);
xor U19236 (N_19236,N_17765,N_17411);
or U19237 (N_19237,N_17735,N_16138);
or U19238 (N_19238,N_16895,N_16769);
nand U19239 (N_19239,N_17261,N_17573);
and U19240 (N_19240,N_16764,N_17010);
nand U19241 (N_19241,N_17195,N_17495);
xor U19242 (N_19242,N_16718,N_17318);
nand U19243 (N_19243,N_16432,N_17613);
nand U19244 (N_19244,N_16171,N_16846);
nor U19245 (N_19245,N_17414,N_17732);
and U19246 (N_19246,N_17387,N_17995);
nand U19247 (N_19247,N_16368,N_16806);
or U19248 (N_19248,N_16462,N_16787);
xnor U19249 (N_19249,N_16677,N_17648);
nand U19250 (N_19250,N_16451,N_17398);
and U19251 (N_19251,N_16097,N_16680);
nor U19252 (N_19252,N_17488,N_16927);
and U19253 (N_19253,N_16157,N_17252);
nor U19254 (N_19254,N_16888,N_17682);
nand U19255 (N_19255,N_16836,N_17014);
nor U19256 (N_19256,N_16667,N_16759);
or U19257 (N_19257,N_16183,N_17181);
nand U19258 (N_19258,N_16166,N_17405);
nor U19259 (N_19259,N_16269,N_17312);
nor U19260 (N_19260,N_16449,N_17435);
and U19261 (N_19261,N_16339,N_17977);
and U19262 (N_19262,N_16701,N_17878);
or U19263 (N_19263,N_16387,N_16999);
and U19264 (N_19264,N_16024,N_17283);
or U19265 (N_19265,N_16254,N_17781);
or U19266 (N_19266,N_16176,N_17476);
nand U19267 (N_19267,N_17240,N_17939);
and U19268 (N_19268,N_16859,N_16881);
and U19269 (N_19269,N_17272,N_17906);
nor U19270 (N_19270,N_17931,N_17841);
or U19271 (N_19271,N_16012,N_17625);
nand U19272 (N_19272,N_17434,N_17216);
and U19273 (N_19273,N_16778,N_17257);
nor U19274 (N_19274,N_16172,N_17228);
nand U19275 (N_19275,N_16926,N_17754);
xor U19276 (N_19276,N_17818,N_17396);
or U19277 (N_19277,N_16365,N_16227);
xor U19278 (N_19278,N_17548,N_16851);
nor U19279 (N_19279,N_17552,N_17508);
or U19280 (N_19280,N_16811,N_17760);
and U19281 (N_19281,N_16106,N_17538);
nand U19282 (N_19282,N_17354,N_17084);
nor U19283 (N_19283,N_17324,N_16238);
nand U19284 (N_19284,N_17898,N_17631);
or U19285 (N_19285,N_17506,N_17868);
nor U19286 (N_19286,N_17811,N_16386);
or U19287 (N_19287,N_17528,N_16715);
xnor U19288 (N_19288,N_17653,N_17176);
nand U19289 (N_19289,N_17675,N_17485);
xor U19290 (N_19290,N_16824,N_16968);
xor U19291 (N_19291,N_17707,N_17937);
or U19292 (N_19292,N_17771,N_17187);
and U19293 (N_19293,N_16243,N_16533);
nor U19294 (N_19294,N_17374,N_16313);
and U19295 (N_19295,N_17206,N_17401);
nand U19296 (N_19296,N_17883,N_17444);
or U19297 (N_19297,N_16451,N_17235);
xor U19298 (N_19298,N_16493,N_16242);
nor U19299 (N_19299,N_17367,N_16824);
and U19300 (N_19300,N_17157,N_17022);
or U19301 (N_19301,N_16332,N_16729);
nor U19302 (N_19302,N_17508,N_17418);
xnor U19303 (N_19303,N_16161,N_16642);
nor U19304 (N_19304,N_16619,N_17672);
nor U19305 (N_19305,N_17380,N_17723);
nand U19306 (N_19306,N_17471,N_16526);
nor U19307 (N_19307,N_17513,N_16339);
or U19308 (N_19308,N_17206,N_16934);
and U19309 (N_19309,N_16446,N_16714);
and U19310 (N_19310,N_16151,N_17479);
or U19311 (N_19311,N_17771,N_17386);
nand U19312 (N_19312,N_17870,N_16238);
nand U19313 (N_19313,N_16562,N_17916);
nor U19314 (N_19314,N_16018,N_17549);
or U19315 (N_19315,N_16690,N_17304);
or U19316 (N_19316,N_16652,N_16265);
or U19317 (N_19317,N_17186,N_16393);
nand U19318 (N_19318,N_16958,N_17631);
and U19319 (N_19319,N_16019,N_17077);
and U19320 (N_19320,N_16228,N_16209);
nand U19321 (N_19321,N_16169,N_17477);
xnor U19322 (N_19322,N_16646,N_17342);
or U19323 (N_19323,N_16122,N_16491);
nor U19324 (N_19324,N_17123,N_16159);
and U19325 (N_19325,N_16315,N_17973);
nand U19326 (N_19326,N_16968,N_17346);
nor U19327 (N_19327,N_17044,N_17269);
xor U19328 (N_19328,N_16299,N_17635);
xor U19329 (N_19329,N_16358,N_17122);
nand U19330 (N_19330,N_17747,N_16754);
or U19331 (N_19331,N_16975,N_16776);
nor U19332 (N_19332,N_17897,N_16116);
and U19333 (N_19333,N_17578,N_16686);
or U19334 (N_19334,N_16177,N_17623);
nor U19335 (N_19335,N_16292,N_16491);
nor U19336 (N_19336,N_16416,N_17460);
nor U19337 (N_19337,N_16874,N_16131);
nor U19338 (N_19338,N_16317,N_16923);
nor U19339 (N_19339,N_16648,N_16126);
xnor U19340 (N_19340,N_16731,N_17698);
and U19341 (N_19341,N_16351,N_17159);
nand U19342 (N_19342,N_17447,N_16755);
xor U19343 (N_19343,N_16167,N_16392);
nor U19344 (N_19344,N_16875,N_17244);
or U19345 (N_19345,N_17093,N_16925);
xnor U19346 (N_19346,N_16388,N_17949);
xnor U19347 (N_19347,N_17307,N_16404);
nor U19348 (N_19348,N_16326,N_16393);
nand U19349 (N_19349,N_16011,N_17359);
xnor U19350 (N_19350,N_17832,N_16793);
nand U19351 (N_19351,N_16485,N_17696);
and U19352 (N_19352,N_16790,N_16628);
nand U19353 (N_19353,N_17001,N_16527);
and U19354 (N_19354,N_17071,N_16465);
or U19355 (N_19355,N_17343,N_17315);
nand U19356 (N_19356,N_16275,N_16200);
and U19357 (N_19357,N_17954,N_17358);
or U19358 (N_19358,N_17279,N_17586);
nor U19359 (N_19359,N_16904,N_16351);
xnor U19360 (N_19360,N_17611,N_17836);
xnor U19361 (N_19361,N_17204,N_17452);
xor U19362 (N_19362,N_17225,N_16749);
nor U19363 (N_19363,N_16074,N_17545);
nor U19364 (N_19364,N_17956,N_16775);
xor U19365 (N_19365,N_17999,N_17230);
and U19366 (N_19366,N_17497,N_17842);
and U19367 (N_19367,N_17281,N_16098);
nor U19368 (N_19368,N_16508,N_16161);
nor U19369 (N_19369,N_16500,N_16708);
and U19370 (N_19370,N_17506,N_17196);
nor U19371 (N_19371,N_17182,N_17560);
nor U19372 (N_19372,N_16498,N_16196);
xor U19373 (N_19373,N_16759,N_16652);
or U19374 (N_19374,N_16960,N_16105);
nand U19375 (N_19375,N_16643,N_17725);
nand U19376 (N_19376,N_16936,N_17508);
and U19377 (N_19377,N_17394,N_16154);
and U19378 (N_19378,N_17370,N_17692);
nand U19379 (N_19379,N_17945,N_16909);
nor U19380 (N_19380,N_17877,N_17099);
nand U19381 (N_19381,N_16359,N_16695);
and U19382 (N_19382,N_16120,N_17056);
nand U19383 (N_19383,N_16419,N_17995);
nor U19384 (N_19384,N_16840,N_17674);
and U19385 (N_19385,N_17526,N_17229);
or U19386 (N_19386,N_16794,N_17012);
xnor U19387 (N_19387,N_16852,N_16589);
or U19388 (N_19388,N_17778,N_17830);
or U19389 (N_19389,N_16798,N_17843);
and U19390 (N_19390,N_17334,N_17030);
or U19391 (N_19391,N_16931,N_17688);
nor U19392 (N_19392,N_17984,N_16105);
xor U19393 (N_19393,N_16649,N_16964);
nand U19394 (N_19394,N_16637,N_16079);
and U19395 (N_19395,N_17553,N_17203);
nor U19396 (N_19396,N_16873,N_16763);
nand U19397 (N_19397,N_17377,N_17275);
xor U19398 (N_19398,N_16211,N_17125);
nor U19399 (N_19399,N_16117,N_17121);
xnor U19400 (N_19400,N_17462,N_16231);
or U19401 (N_19401,N_17638,N_17916);
nor U19402 (N_19402,N_16292,N_16507);
and U19403 (N_19403,N_16080,N_17099);
nand U19404 (N_19404,N_17833,N_16979);
nor U19405 (N_19405,N_17927,N_16004);
nor U19406 (N_19406,N_16512,N_16618);
nor U19407 (N_19407,N_16437,N_17680);
nor U19408 (N_19408,N_17863,N_16660);
nand U19409 (N_19409,N_16613,N_17655);
nor U19410 (N_19410,N_17159,N_16411);
nor U19411 (N_19411,N_17548,N_16120);
or U19412 (N_19412,N_16217,N_17190);
xnor U19413 (N_19413,N_17740,N_17728);
xnor U19414 (N_19414,N_17157,N_17172);
nand U19415 (N_19415,N_16159,N_16698);
or U19416 (N_19416,N_17988,N_16854);
nor U19417 (N_19417,N_17825,N_16373);
xnor U19418 (N_19418,N_17000,N_16987);
xnor U19419 (N_19419,N_16953,N_17840);
nor U19420 (N_19420,N_16627,N_16632);
nor U19421 (N_19421,N_16486,N_17556);
xor U19422 (N_19422,N_16484,N_16651);
xnor U19423 (N_19423,N_16423,N_17584);
xor U19424 (N_19424,N_16639,N_17631);
xor U19425 (N_19425,N_16152,N_16440);
nor U19426 (N_19426,N_16899,N_17279);
or U19427 (N_19427,N_17692,N_17110);
xor U19428 (N_19428,N_17999,N_17362);
or U19429 (N_19429,N_16930,N_17581);
or U19430 (N_19430,N_16669,N_16832);
nand U19431 (N_19431,N_16864,N_16463);
or U19432 (N_19432,N_17280,N_16466);
nand U19433 (N_19433,N_17154,N_17723);
nor U19434 (N_19434,N_16181,N_17099);
nor U19435 (N_19435,N_16351,N_17792);
or U19436 (N_19436,N_17371,N_16222);
and U19437 (N_19437,N_17492,N_17508);
or U19438 (N_19438,N_17818,N_17268);
nand U19439 (N_19439,N_17085,N_17286);
nor U19440 (N_19440,N_17286,N_16132);
nand U19441 (N_19441,N_17203,N_16007);
nor U19442 (N_19442,N_16311,N_17843);
nand U19443 (N_19443,N_17632,N_17765);
xnor U19444 (N_19444,N_17464,N_17712);
and U19445 (N_19445,N_16228,N_17288);
nand U19446 (N_19446,N_16583,N_17100);
or U19447 (N_19447,N_17337,N_16961);
xor U19448 (N_19448,N_17385,N_17490);
nor U19449 (N_19449,N_16794,N_16490);
and U19450 (N_19450,N_17483,N_17105);
nand U19451 (N_19451,N_17188,N_16380);
or U19452 (N_19452,N_16972,N_17536);
nor U19453 (N_19453,N_16661,N_16852);
nand U19454 (N_19454,N_16600,N_17334);
nor U19455 (N_19455,N_17863,N_17902);
and U19456 (N_19456,N_16667,N_17244);
nor U19457 (N_19457,N_16853,N_17651);
xnor U19458 (N_19458,N_17111,N_16690);
xnor U19459 (N_19459,N_17753,N_16981);
nor U19460 (N_19460,N_16156,N_17233);
nand U19461 (N_19461,N_17732,N_17492);
or U19462 (N_19462,N_17184,N_16731);
xor U19463 (N_19463,N_16983,N_16875);
xor U19464 (N_19464,N_16539,N_17909);
nand U19465 (N_19465,N_16859,N_16482);
xor U19466 (N_19466,N_16292,N_16718);
xnor U19467 (N_19467,N_17293,N_17660);
nand U19468 (N_19468,N_16695,N_16685);
or U19469 (N_19469,N_16566,N_16170);
xnor U19470 (N_19470,N_16670,N_16581);
nand U19471 (N_19471,N_17574,N_17485);
or U19472 (N_19472,N_16009,N_16735);
or U19473 (N_19473,N_17394,N_17780);
nand U19474 (N_19474,N_17023,N_16292);
xor U19475 (N_19475,N_16637,N_17872);
nor U19476 (N_19476,N_17568,N_16024);
nor U19477 (N_19477,N_16305,N_16797);
nand U19478 (N_19478,N_16772,N_17785);
nor U19479 (N_19479,N_16222,N_16236);
xnor U19480 (N_19480,N_17898,N_16057);
nor U19481 (N_19481,N_16082,N_17619);
nand U19482 (N_19482,N_16282,N_16790);
nor U19483 (N_19483,N_17226,N_17972);
nand U19484 (N_19484,N_16609,N_16937);
nand U19485 (N_19485,N_16402,N_17238);
nand U19486 (N_19486,N_17770,N_17873);
nor U19487 (N_19487,N_16504,N_16181);
and U19488 (N_19488,N_17642,N_17528);
or U19489 (N_19489,N_17466,N_17829);
nor U19490 (N_19490,N_17309,N_16842);
and U19491 (N_19491,N_17344,N_16265);
nand U19492 (N_19492,N_16031,N_17388);
nor U19493 (N_19493,N_17557,N_17742);
nor U19494 (N_19494,N_17380,N_16852);
nor U19495 (N_19495,N_17780,N_17523);
nor U19496 (N_19496,N_17026,N_17308);
nand U19497 (N_19497,N_16457,N_16581);
nor U19498 (N_19498,N_16943,N_16393);
nand U19499 (N_19499,N_16181,N_17182);
or U19500 (N_19500,N_17205,N_17729);
xnor U19501 (N_19501,N_17559,N_17424);
or U19502 (N_19502,N_17284,N_17859);
nor U19503 (N_19503,N_16980,N_16879);
or U19504 (N_19504,N_16976,N_17612);
nand U19505 (N_19505,N_17636,N_17245);
and U19506 (N_19506,N_16972,N_16533);
or U19507 (N_19507,N_16741,N_17111);
xor U19508 (N_19508,N_16965,N_17909);
xor U19509 (N_19509,N_16371,N_16764);
and U19510 (N_19510,N_16667,N_17047);
and U19511 (N_19511,N_17643,N_16444);
or U19512 (N_19512,N_16962,N_16034);
xnor U19513 (N_19513,N_17796,N_17622);
and U19514 (N_19514,N_16289,N_16039);
nor U19515 (N_19515,N_17445,N_17104);
nand U19516 (N_19516,N_17156,N_17897);
nand U19517 (N_19517,N_17425,N_17340);
and U19518 (N_19518,N_16669,N_17100);
nor U19519 (N_19519,N_17798,N_17499);
nand U19520 (N_19520,N_17418,N_17723);
nor U19521 (N_19521,N_17762,N_17670);
nand U19522 (N_19522,N_17057,N_16299);
nor U19523 (N_19523,N_16467,N_16848);
xor U19524 (N_19524,N_17878,N_16747);
nor U19525 (N_19525,N_17222,N_17389);
or U19526 (N_19526,N_16432,N_16387);
or U19527 (N_19527,N_17955,N_17553);
or U19528 (N_19528,N_17905,N_16908);
and U19529 (N_19529,N_16657,N_17830);
xor U19530 (N_19530,N_17723,N_17651);
xnor U19531 (N_19531,N_17857,N_16552);
and U19532 (N_19532,N_16188,N_17667);
and U19533 (N_19533,N_17044,N_17398);
xor U19534 (N_19534,N_16288,N_17013);
or U19535 (N_19535,N_16609,N_16841);
xnor U19536 (N_19536,N_17897,N_16179);
nand U19537 (N_19537,N_17531,N_17316);
xnor U19538 (N_19538,N_17794,N_16528);
nor U19539 (N_19539,N_16766,N_16075);
xnor U19540 (N_19540,N_17346,N_17904);
nor U19541 (N_19541,N_16274,N_17545);
and U19542 (N_19542,N_16540,N_16884);
nor U19543 (N_19543,N_17343,N_16861);
xor U19544 (N_19544,N_16702,N_16947);
and U19545 (N_19545,N_17450,N_16850);
xor U19546 (N_19546,N_17830,N_17581);
xor U19547 (N_19547,N_17402,N_17173);
or U19548 (N_19548,N_17275,N_16807);
xor U19549 (N_19549,N_17368,N_17078);
nand U19550 (N_19550,N_16117,N_16842);
or U19551 (N_19551,N_16844,N_17767);
nor U19552 (N_19552,N_16048,N_17610);
nand U19553 (N_19553,N_16357,N_17443);
nor U19554 (N_19554,N_16680,N_17810);
and U19555 (N_19555,N_17508,N_16492);
nand U19556 (N_19556,N_16101,N_16198);
or U19557 (N_19557,N_17893,N_16244);
xnor U19558 (N_19558,N_16275,N_16534);
and U19559 (N_19559,N_16082,N_17712);
and U19560 (N_19560,N_16198,N_16688);
nand U19561 (N_19561,N_17317,N_16588);
and U19562 (N_19562,N_17037,N_16960);
nor U19563 (N_19563,N_17509,N_16912);
nand U19564 (N_19564,N_17740,N_17736);
and U19565 (N_19565,N_17592,N_16014);
xnor U19566 (N_19566,N_17604,N_16864);
or U19567 (N_19567,N_16237,N_16255);
or U19568 (N_19568,N_17762,N_16776);
nand U19569 (N_19569,N_17891,N_16811);
nor U19570 (N_19570,N_17809,N_17922);
nand U19571 (N_19571,N_17104,N_16465);
and U19572 (N_19572,N_16294,N_17026);
xnor U19573 (N_19573,N_16216,N_16381);
xnor U19574 (N_19574,N_16309,N_17517);
or U19575 (N_19575,N_16807,N_16918);
and U19576 (N_19576,N_17291,N_17444);
nor U19577 (N_19577,N_17432,N_17201);
nor U19578 (N_19578,N_17348,N_16053);
or U19579 (N_19579,N_16689,N_17076);
and U19580 (N_19580,N_16218,N_16635);
nand U19581 (N_19581,N_16865,N_16660);
and U19582 (N_19582,N_17756,N_16129);
xor U19583 (N_19583,N_17664,N_17597);
nor U19584 (N_19584,N_16446,N_16145);
xnor U19585 (N_19585,N_17529,N_17891);
xor U19586 (N_19586,N_16462,N_16645);
nand U19587 (N_19587,N_17449,N_17298);
nand U19588 (N_19588,N_17220,N_16744);
or U19589 (N_19589,N_17129,N_17617);
nor U19590 (N_19590,N_17466,N_16637);
or U19591 (N_19591,N_16061,N_16379);
nor U19592 (N_19592,N_17334,N_16403);
and U19593 (N_19593,N_16268,N_16647);
xnor U19594 (N_19594,N_17258,N_17945);
or U19595 (N_19595,N_16443,N_16015);
xor U19596 (N_19596,N_16292,N_17684);
nand U19597 (N_19597,N_17314,N_17356);
or U19598 (N_19598,N_16544,N_17221);
nor U19599 (N_19599,N_17395,N_17383);
and U19600 (N_19600,N_17274,N_17955);
xor U19601 (N_19601,N_17153,N_17690);
xor U19602 (N_19602,N_17541,N_16958);
xnor U19603 (N_19603,N_16517,N_17105);
xnor U19604 (N_19604,N_16567,N_16269);
nand U19605 (N_19605,N_17519,N_17401);
nand U19606 (N_19606,N_17176,N_17633);
xnor U19607 (N_19607,N_17374,N_16629);
nand U19608 (N_19608,N_16201,N_16179);
or U19609 (N_19609,N_16740,N_16782);
nand U19610 (N_19610,N_16977,N_17216);
and U19611 (N_19611,N_16842,N_16824);
and U19612 (N_19612,N_16490,N_17243);
xnor U19613 (N_19613,N_16564,N_16502);
nor U19614 (N_19614,N_16453,N_16638);
and U19615 (N_19615,N_16136,N_17438);
and U19616 (N_19616,N_16395,N_17109);
and U19617 (N_19617,N_17325,N_16401);
or U19618 (N_19618,N_17985,N_16835);
and U19619 (N_19619,N_17980,N_17134);
nor U19620 (N_19620,N_17100,N_17492);
nor U19621 (N_19621,N_16608,N_16190);
and U19622 (N_19622,N_17700,N_17927);
or U19623 (N_19623,N_17155,N_17301);
or U19624 (N_19624,N_17448,N_17589);
and U19625 (N_19625,N_16977,N_17025);
nand U19626 (N_19626,N_16799,N_16417);
and U19627 (N_19627,N_17682,N_17533);
nand U19628 (N_19628,N_17634,N_17664);
or U19629 (N_19629,N_16847,N_17493);
xnor U19630 (N_19630,N_17920,N_17988);
or U19631 (N_19631,N_16426,N_16801);
and U19632 (N_19632,N_17285,N_16836);
xnor U19633 (N_19633,N_17098,N_16380);
nand U19634 (N_19634,N_17712,N_16790);
or U19635 (N_19635,N_17801,N_16770);
or U19636 (N_19636,N_17868,N_16883);
or U19637 (N_19637,N_17181,N_17855);
and U19638 (N_19638,N_17801,N_16927);
xnor U19639 (N_19639,N_17127,N_16764);
or U19640 (N_19640,N_16430,N_17103);
or U19641 (N_19641,N_17547,N_17828);
nor U19642 (N_19642,N_17497,N_17605);
nor U19643 (N_19643,N_16115,N_16961);
or U19644 (N_19644,N_17247,N_17690);
and U19645 (N_19645,N_16354,N_17780);
xor U19646 (N_19646,N_16483,N_17559);
nor U19647 (N_19647,N_16388,N_16393);
nor U19648 (N_19648,N_16387,N_16515);
nor U19649 (N_19649,N_16533,N_17587);
xnor U19650 (N_19650,N_17599,N_17771);
or U19651 (N_19651,N_17125,N_17599);
nand U19652 (N_19652,N_16669,N_17555);
and U19653 (N_19653,N_17930,N_16121);
nand U19654 (N_19654,N_17534,N_17507);
and U19655 (N_19655,N_16856,N_16864);
or U19656 (N_19656,N_16890,N_16400);
and U19657 (N_19657,N_16353,N_17963);
nor U19658 (N_19658,N_17011,N_17640);
or U19659 (N_19659,N_16561,N_17782);
nand U19660 (N_19660,N_16422,N_16552);
nor U19661 (N_19661,N_16621,N_16723);
nor U19662 (N_19662,N_16175,N_16810);
or U19663 (N_19663,N_16970,N_17999);
xor U19664 (N_19664,N_16065,N_16326);
nor U19665 (N_19665,N_17074,N_17884);
or U19666 (N_19666,N_16402,N_17815);
nand U19667 (N_19667,N_17060,N_17093);
xnor U19668 (N_19668,N_16265,N_16826);
or U19669 (N_19669,N_17007,N_16029);
xnor U19670 (N_19670,N_16392,N_16188);
or U19671 (N_19671,N_17822,N_16222);
nand U19672 (N_19672,N_16910,N_17008);
and U19673 (N_19673,N_17554,N_17994);
xnor U19674 (N_19674,N_17963,N_16334);
and U19675 (N_19675,N_17955,N_16430);
xor U19676 (N_19676,N_16785,N_17046);
and U19677 (N_19677,N_16852,N_16946);
nand U19678 (N_19678,N_17215,N_16930);
and U19679 (N_19679,N_17801,N_16971);
or U19680 (N_19680,N_16412,N_16576);
or U19681 (N_19681,N_16550,N_16453);
or U19682 (N_19682,N_16253,N_16415);
xor U19683 (N_19683,N_16739,N_16765);
nor U19684 (N_19684,N_17011,N_17665);
nor U19685 (N_19685,N_16440,N_17081);
or U19686 (N_19686,N_17670,N_16831);
nand U19687 (N_19687,N_17227,N_16172);
nand U19688 (N_19688,N_16092,N_16475);
xnor U19689 (N_19689,N_17162,N_17378);
or U19690 (N_19690,N_17860,N_17498);
nor U19691 (N_19691,N_16508,N_17683);
and U19692 (N_19692,N_16522,N_16626);
and U19693 (N_19693,N_17689,N_17595);
nor U19694 (N_19694,N_17129,N_16409);
xor U19695 (N_19695,N_16847,N_16967);
or U19696 (N_19696,N_17837,N_16257);
or U19697 (N_19697,N_16188,N_17011);
nand U19698 (N_19698,N_17962,N_16732);
and U19699 (N_19699,N_16000,N_16582);
nor U19700 (N_19700,N_17620,N_17344);
xor U19701 (N_19701,N_16034,N_17857);
nand U19702 (N_19702,N_16171,N_17788);
xnor U19703 (N_19703,N_17304,N_17132);
and U19704 (N_19704,N_17201,N_17159);
nand U19705 (N_19705,N_16063,N_16738);
nand U19706 (N_19706,N_17918,N_17318);
xnor U19707 (N_19707,N_17616,N_16024);
nand U19708 (N_19708,N_17612,N_16357);
xor U19709 (N_19709,N_17315,N_17169);
nand U19710 (N_19710,N_16710,N_16198);
xor U19711 (N_19711,N_16191,N_17785);
or U19712 (N_19712,N_16359,N_16445);
nor U19713 (N_19713,N_16198,N_16112);
nand U19714 (N_19714,N_16307,N_16150);
nand U19715 (N_19715,N_16768,N_17847);
nor U19716 (N_19716,N_16883,N_16132);
xor U19717 (N_19717,N_17760,N_17973);
and U19718 (N_19718,N_17025,N_16523);
xnor U19719 (N_19719,N_17632,N_16760);
and U19720 (N_19720,N_17418,N_17833);
nor U19721 (N_19721,N_16636,N_17898);
and U19722 (N_19722,N_16627,N_17330);
nor U19723 (N_19723,N_16829,N_17513);
and U19724 (N_19724,N_16461,N_17560);
or U19725 (N_19725,N_17590,N_16384);
nor U19726 (N_19726,N_16145,N_17115);
or U19727 (N_19727,N_16819,N_16875);
and U19728 (N_19728,N_17514,N_16120);
xor U19729 (N_19729,N_16313,N_17836);
or U19730 (N_19730,N_17674,N_16475);
xnor U19731 (N_19731,N_17335,N_16004);
nand U19732 (N_19732,N_16221,N_17122);
and U19733 (N_19733,N_16447,N_16851);
nand U19734 (N_19734,N_17906,N_17592);
nand U19735 (N_19735,N_16029,N_17998);
or U19736 (N_19736,N_17993,N_16792);
or U19737 (N_19737,N_17511,N_17178);
or U19738 (N_19738,N_17168,N_16408);
or U19739 (N_19739,N_17038,N_17018);
nor U19740 (N_19740,N_17016,N_17708);
xor U19741 (N_19741,N_16195,N_16848);
nor U19742 (N_19742,N_17973,N_16550);
xor U19743 (N_19743,N_16404,N_16186);
and U19744 (N_19744,N_17104,N_17927);
nand U19745 (N_19745,N_16396,N_16110);
nand U19746 (N_19746,N_16428,N_17125);
xnor U19747 (N_19747,N_17298,N_17193);
and U19748 (N_19748,N_16611,N_16589);
nand U19749 (N_19749,N_16497,N_17306);
nand U19750 (N_19750,N_16683,N_16762);
and U19751 (N_19751,N_16828,N_17086);
nor U19752 (N_19752,N_16298,N_16916);
xor U19753 (N_19753,N_17364,N_17708);
nor U19754 (N_19754,N_17210,N_17484);
or U19755 (N_19755,N_17285,N_17481);
and U19756 (N_19756,N_17994,N_16439);
xor U19757 (N_19757,N_16227,N_16031);
or U19758 (N_19758,N_17995,N_16664);
nand U19759 (N_19759,N_16601,N_17522);
or U19760 (N_19760,N_17261,N_17880);
nor U19761 (N_19761,N_16086,N_17847);
nor U19762 (N_19762,N_17263,N_17591);
nor U19763 (N_19763,N_17673,N_16827);
xnor U19764 (N_19764,N_16645,N_16648);
and U19765 (N_19765,N_16741,N_16870);
nor U19766 (N_19766,N_17228,N_17912);
and U19767 (N_19767,N_17530,N_16622);
nand U19768 (N_19768,N_16102,N_16064);
nand U19769 (N_19769,N_17688,N_16610);
xnor U19770 (N_19770,N_17149,N_17793);
xor U19771 (N_19771,N_17937,N_16445);
nand U19772 (N_19772,N_17109,N_17344);
xor U19773 (N_19773,N_17879,N_17934);
nand U19774 (N_19774,N_17587,N_17004);
nor U19775 (N_19775,N_17055,N_16856);
or U19776 (N_19776,N_16335,N_16236);
or U19777 (N_19777,N_16563,N_17921);
xor U19778 (N_19778,N_17330,N_16324);
and U19779 (N_19779,N_16273,N_16993);
or U19780 (N_19780,N_17613,N_16830);
nand U19781 (N_19781,N_16705,N_17570);
xnor U19782 (N_19782,N_17456,N_16561);
or U19783 (N_19783,N_17527,N_17886);
and U19784 (N_19784,N_16996,N_16473);
and U19785 (N_19785,N_17750,N_17312);
xnor U19786 (N_19786,N_17866,N_16011);
nor U19787 (N_19787,N_17476,N_17068);
nand U19788 (N_19788,N_17704,N_17610);
nor U19789 (N_19789,N_17510,N_16853);
and U19790 (N_19790,N_16114,N_16187);
and U19791 (N_19791,N_17897,N_17693);
nand U19792 (N_19792,N_16834,N_17761);
nor U19793 (N_19793,N_16151,N_16004);
nand U19794 (N_19794,N_16702,N_17575);
or U19795 (N_19795,N_17608,N_16883);
nor U19796 (N_19796,N_16998,N_17471);
and U19797 (N_19797,N_16123,N_16291);
xnor U19798 (N_19798,N_17316,N_17427);
or U19799 (N_19799,N_16358,N_16285);
or U19800 (N_19800,N_17701,N_16080);
nor U19801 (N_19801,N_17458,N_16307);
xnor U19802 (N_19802,N_17301,N_17504);
and U19803 (N_19803,N_17995,N_17187);
or U19804 (N_19804,N_17797,N_16377);
and U19805 (N_19805,N_16108,N_17549);
nor U19806 (N_19806,N_17544,N_17011);
or U19807 (N_19807,N_17026,N_17091);
and U19808 (N_19808,N_17376,N_17807);
or U19809 (N_19809,N_17431,N_17196);
or U19810 (N_19810,N_17922,N_16017);
nand U19811 (N_19811,N_16735,N_17228);
nor U19812 (N_19812,N_16292,N_16220);
nor U19813 (N_19813,N_16617,N_17730);
nand U19814 (N_19814,N_16766,N_17008);
and U19815 (N_19815,N_16895,N_16065);
xor U19816 (N_19816,N_16558,N_17793);
nand U19817 (N_19817,N_17970,N_16460);
xor U19818 (N_19818,N_16845,N_17718);
or U19819 (N_19819,N_16767,N_16259);
nor U19820 (N_19820,N_16208,N_16302);
nor U19821 (N_19821,N_16691,N_17681);
xor U19822 (N_19822,N_17630,N_16876);
nand U19823 (N_19823,N_16238,N_17495);
and U19824 (N_19824,N_17539,N_17327);
xor U19825 (N_19825,N_16931,N_16068);
nand U19826 (N_19826,N_17943,N_16803);
or U19827 (N_19827,N_16376,N_16103);
nand U19828 (N_19828,N_16485,N_17887);
xor U19829 (N_19829,N_17128,N_17116);
nor U19830 (N_19830,N_16150,N_16385);
nand U19831 (N_19831,N_16041,N_16328);
or U19832 (N_19832,N_17933,N_16993);
and U19833 (N_19833,N_17446,N_16418);
nand U19834 (N_19834,N_16379,N_16845);
and U19835 (N_19835,N_16446,N_16625);
and U19836 (N_19836,N_16706,N_17460);
nor U19837 (N_19837,N_17243,N_16528);
or U19838 (N_19838,N_17916,N_17902);
or U19839 (N_19839,N_16612,N_16424);
nor U19840 (N_19840,N_17567,N_16790);
xor U19841 (N_19841,N_17497,N_16930);
xor U19842 (N_19842,N_16518,N_16654);
xnor U19843 (N_19843,N_16891,N_16031);
or U19844 (N_19844,N_17633,N_17427);
nand U19845 (N_19845,N_16845,N_17764);
and U19846 (N_19846,N_16773,N_17291);
or U19847 (N_19847,N_17044,N_16654);
nor U19848 (N_19848,N_16220,N_16259);
nor U19849 (N_19849,N_16436,N_16947);
xor U19850 (N_19850,N_17389,N_17531);
xor U19851 (N_19851,N_17341,N_16721);
or U19852 (N_19852,N_16548,N_16303);
xor U19853 (N_19853,N_16727,N_17041);
and U19854 (N_19854,N_16858,N_16554);
nor U19855 (N_19855,N_16389,N_17942);
or U19856 (N_19856,N_16545,N_16553);
nand U19857 (N_19857,N_16755,N_16442);
xor U19858 (N_19858,N_16180,N_16380);
or U19859 (N_19859,N_16394,N_16696);
nand U19860 (N_19860,N_17086,N_17024);
nor U19861 (N_19861,N_16623,N_17927);
xnor U19862 (N_19862,N_16005,N_17840);
nand U19863 (N_19863,N_16440,N_16945);
and U19864 (N_19864,N_17747,N_16958);
and U19865 (N_19865,N_17643,N_16284);
nor U19866 (N_19866,N_17466,N_17024);
or U19867 (N_19867,N_17792,N_17169);
and U19868 (N_19868,N_16092,N_16488);
nor U19869 (N_19869,N_16411,N_17896);
and U19870 (N_19870,N_16480,N_17480);
xor U19871 (N_19871,N_16697,N_17234);
xnor U19872 (N_19872,N_17084,N_16354);
xor U19873 (N_19873,N_16862,N_17651);
nor U19874 (N_19874,N_17681,N_16825);
or U19875 (N_19875,N_16931,N_16752);
or U19876 (N_19876,N_17604,N_17451);
xor U19877 (N_19877,N_17738,N_16226);
or U19878 (N_19878,N_17614,N_17058);
and U19879 (N_19879,N_17619,N_17869);
nand U19880 (N_19880,N_16198,N_16159);
or U19881 (N_19881,N_16234,N_16075);
or U19882 (N_19882,N_16348,N_16622);
or U19883 (N_19883,N_16280,N_17883);
nand U19884 (N_19884,N_17571,N_16302);
and U19885 (N_19885,N_16224,N_16020);
and U19886 (N_19886,N_16625,N_16179);
xor U19887 (N_19887,N_16666,N_16820);
or U19888 (N_19888,N_17019,N_16336);
xor U19889 (N_19889,N_17710,N_16932);
xnor U19890 (N_19890,N_16440,N_16023);
or U19891 (N_19891,N_16762,N_17864);
nor U19892 (N_19892,N_16650,N_17806);
and U19893 (N_19893,N_17451,N_17631);
nand U19894 (N_19894,N_17666,N_17216);
xnor U19895 (N_19895,N_17036,N_17354);
and U19896 (N_19896,N_16315,N_17401);
nor U19897 (N_19897,N_16197,N_17282);
nand U19898 (N_19898,N_16179,N_17507);
nor U19899 (N_19899,N_16655,N_17699);
nor U19900 (N_19900,N_17613,N_16446);
xnor U19901 (N_19901,N_17434,N_16056);
or U19902 (N_19902,N_17213,N_16298);
xnor U19903 (N_19903,N_16076,N_17722);
xnor U19904 (N_19904,N_17714,N_17160);
nand U19905 (N_19905,N_16092,N_16612);
xor U19906 (N_19906,N_16721,N_17304);
nor U19907 (N_19907,N_16908,N_17676);
or U19908 (N_19908,N_17821,N_17312);
nand U19909 (N_19909,N_16803,N_17793);
xor U19910 (N_19910,N_16418,N_17944);
and U19911 (N_19911,N_16235,N_16470);
nor U19912 (N_19912,N_16476,N_16965);
and U19913 (N_19913,N_16135,N_16085);
nand U19914 (N_19914,N_16944,N_17941);
xnor U19915 (N_19915,N_16372,N_16665);
xnor U19916 (N_19916,N_16872,N_16464);
nor U19917 (N_19917,N_16003,N_17165);
nor U19918 (N_19918,N_17360,N_17567);
nor U19919 (N_19919,N_17924,N_16343);
or U19920 (N_19920,N_17667,N_17783);
nand U19921 (N_19921,N_17415,N_16764);
or U19922 (N_19922,N_17854,N_17041);
and U19923 (N_19923,N_16293,N_16371);
and U19924 (N_19924,N_16919,N_16152);
nor U19925 (N_19925,N_17181,N_17996);
nor U19926 (N_19926,N_16538,N_16056);
or U19927 (N_19927,N_16412,N_16477);
xor U19928 (N_19928,N_16365,N_16313);
nor U19929 (N_19929,N_17305,N_17814);
xnor U19930 (N_19930,N_16430,N_17273);
or U19931 (N_19931,N_17147,N_16348);
nand U19932 (N_19932,N_16033,N_17038);
and U19933 (N_19933,N_16355,N_16283);
or U19934 (N_19934,N_16299,N_16406);
nand U19935 (N_19935,N_16160,N_17659);
or U19936 (N_19936,N_16713,N_17018);
or U19937 (N_19937,N_17306,N_16870);
nor U19938 (N_19938,N_16528,N_16553);
nand U19939 (N_19939,N_17078,N_16968);
and U19940 (N_19940,N_17970,N_16730);
or U19941 (N_19941,N_16622,N_16097);
and U19942 (N_19942,N_17065,N_17023);
nand U19943 (N_19943,N_17542,N_17389);
and U19944 (N_19944,N_16279,N_17663);
and U19945 (N_19945,N_17356,N_16189);
nor U19946 (N_19946,N_16246,N_17295);
nor U19947 (N_19947,N_16492,N_17865);
xor U19948 (N_19948,N_16272,N_17299);
xor U19949 (N_19949,N_16471,N_17027);
or U19950 (N_19950,N_16301,N_16962);
or U19951 (N_19951,N_17965,N_16868);
nor U19952 (N_19952,N_16540,N_16457);
or U19953 (N_19953,N_16952,N_16869);
nor U19954 (N_19954,N_17088,N_16167);
nor U19955 (N_19955,N_17465,N_16555);
nand U19956 (N_19956,N_17385,N_16577);
xor U19957 (N_19957,N_17602,N_16946);
and U19958 (N_19958,N_16162,N_17350);
nand U19959 (N_19959,N_16098,N_17688);
nor U19960 (N_19960,N_17638,N_16960);
xnor U19961 (N_19961,N_16819,N_16641);
or U19962 (N_19962,N_17182,N_16783);
or U19963 (N_19963,N_16109,N_16089);
nor U19964 (N_19964,N_16806,N_17377);
and U19965 (N_19965,N_16880,N_16343);
xor U19966 (N_19966,N_16788,N_16463);
or U19967 (N_19967,N_16055,N_17895);
xnor U19968 (N_19968,N_16665,N_17913);
xnor U19969 (N_19969,N_16902,N_17932);
nor U19970 (N_19970,N_17363,N_17993);
or U19971 (N_19971,N_16640,N_16409);
nor U19972 (N_19972,N_16320,N_17427);
nand U19973 (N_19973,N_17411,N_16445);
or U19974 (N_19974,N_17724,N_17602);
and U19975 (N_19975,N_16376,N_17427);
xor U19976 (N_19976,N_17730,N_16990);
nand U19977 (N_19977,N_17434,N_16067);
nand U19978 (N_19978,N_17100,N_17382);
and U19979 (N_19979,N_17447,N_16818);
or U19980 (N_19980,N_17215,N_17867);
and U19981 (N_19981,N_17223,N_17856);
nor U19982 (N_19982,N_16758,N_16886);
or U19983 (N_19983,N_17482,N_17978);
nor U19984 (N_19984,N_16478,N_16963);
and U19985 (N_19985,N_17928,N_17383);
and U19986 (N_19986,N_16452,N_16952);
nand U19987 (N_19987,N_17645,N_17465);
nor U19988 (N_19988,N_16612,N_17598);
xor U19989 (N_19989,N_16783,N_17563);
or U19990 (N_19990,N_16945,N_16737);
and U19991 (N_19991,N_17828,N_16785);
and U19992 (N_19992,N_17971,N_17890);
nor U19993 (N_19993,N_16844,N_17020);
or U19994 (N_19994,N_17523,N_17409);
nor U19995 (N_19995,N_17047,N_16412);
or U19996 (N_19996,N_17030,N_17338);
xor U19997 (N_19997,N_17393,N_17374);
xor U19998 (N_19998,N_16911,N_16948);
and U19999 (N_19999,N_17459,N_16737);
nand U20000 (N_20000,N_18452,N_18700);
xor U20001 (N_20001,N_18492,N_19184);
nor U20002 (N_20002,N_19227,N_19755);
nand U20003 (N_20003,N_18319,N_19158);
nor U20004 (N_20004,N_18054,N_19068);
and U20005 (N_20005,N_19396,N_18393);
and U20006 (N_20006,N_19077,N_18638);
nand U20007 (N_20007,N_18411,N_18625);
nand U20008 (N_20008,N_19290,N_18973);
nand U20009 (N_20009,N_19766,N_18690);
nand U20010 (N_20010,N_19540,N_19357);
and U20011 (N_20011,N_19023,N_18056);
and U20012 (N_20012,N_19124,N_18738);
and U20013 (N_20013,N_19033,N_19499);
and U20014 (N_20014,N_18962,N_18339);
xor U20015 (N_20015,N_18156,N_19727);
xnor U20016 (N_20016,N_18821,N_18155);
nand U20017 (N_20017,N_18385,N_18554);
nand U20018 (N_20018,N_18015,N_18640);
nor U20019 (N_20019,N_18489,N_18151);
xor U20020 (N_20020,N_19716,N_19643);
nor U20021 (N_20021,N_19853,N_18753);
nand U20022 (N_20022,N_18429,N_18143);
or U20023 (N_20023,N_19194,N_18482);
and U20024 (N_20024,N_19329,N_18943);
or U20025 (N_20025,N_19059,N_19537);
nand U20026 (N_20026,N_18849,N_18032);
and U20027 (N_20027,N_19423,N_19425);
nand U20028 (N_20028,N_18951,N_19688);
nor U20029 (N_20029,N_19260,N_19702);
xnor U20030 (N_20030,N_19620,N_19377);
or U20031 (N_20031,N_19681,N_19833);
nor U20032 (N_20032,N_18696,N_18689);
and U20033 (N_20033,N_18179,N_18108);
or U20034 (N_20034,N_18802,N_19299);
and U20035 (N_20035,N_18290,N_18342);
nor U20036 (N_20036,N_19690,N_18978);
and U20037 (N_20037,N_18534,N_18910);
or U20038 (N_20038,N_19141,N_18722);
and U20039 (N_20039,N_19202,N_18016);
and U20040 (N_20040,N_19579,N_19862);
and U20041 (N_20041,N_18217,N_18855);
nor U20042 (N_20042,N_18386,N_18782);
nor U20043 (N_20043,N_19957,N_19349);
nand U20044 (N_20044,N_18323,N_18642);
nor U20045 (N_20045,N_19952,N_18355);
xnor U20046 (N_20046,N_18245,N_19713);
nor U20047 (N_20047,N_19895,N_19315);
or U20048 (N_20048,N_19422,N_18511);
and U20049 (N_20049,N_19750,N_19719);
and U20050 (N_20050,N_19804,N_19117);
or U20051 (N_20051,N_18714,N_18878);
and U20052 (N_20052,N_18925,N_19032);
nand U20053 (N_20053,N_19872,N_19510);
nor U20054 (N_20054,N_19498,N_18706);
nand U20055 (N_20055,N_19138,N_19506);
nor U20056 (N_20056,N_18189,N_19283);
or U20057 (N_20057,N_19372,N_19896);
and U20058 (N_20058,N_19263,N_18129);
nor U20059 (N_20059,N_18516,N_18705);
and U20060 (N_20060,N_19293,N_18093);
and U20061 (N_20061,N_19947,N_19687);
and U20062 (N_20062,N_19663,N_18409);
or U20063 (N_20063,N_19777,N_18546);
xor U20064 (N_20064,N_19522,N_19883);
nor U20065 (N_20065,N_19708,N_18278);
and U20066 (N_20066,N_18915,N_18646);
xnor U20067 (N_20067,N_18345,N_19876);
and U20068 (N_20068,N_18947,N_19289);
xor U20069 (N_20069,N_18993,N_18987);
and U20070 (N_20070,N_18160,N_18281);
nor U20071 (N_20071,N_18203,N_19135);
or U20072 (N_20072,N_18034,N_19346);
and U20073 (N_20073,N_18443,N_19507);
xnor U20074 (N_20074,N_19359,N_18930);
nand U20075 (N_20075,N_19277,N_19519);
or U20076 (N_20076,N_19917,N_18515);
nor U20077 (N_20077,N_19257,N_18748);
xnor U20078 (N_20078,N_18717,N_18576);
and U20079 (N_20079,N_19742,N_18966);
or U20080 (N_20080,N_18436,N_19776);
and U20081 (N_20081,N_18922,N_19902);
and U20082 (N_20082,N_19928,N_18502);
nand U20083 (N_20083,N_19144,N_18266);
and U20084 (N_20084,N_18424,N_19993);
or U20085 (N_20085,N_19903,N_19464);
or U20086 (N_20086,N_18289,N_19893);
nand U20087 (N_20087,N_19218,N_19488);
nand U20088 (N_20088,N_18138,N_19604);
and U20089 (N_20089,N_18604,N_18383);
nand U20090 (N_20090,N_19764,N_19255);
xnor U20091 (N_20091,N_19955,N_19948);
nor U20092 (N_20092,N_18685,N_19244);
nor U20093 (N_20093,N_18663,N_18486);
xor U20094 (N_20094,N_18288,N_18140);
nand U20095 (N_20095,N_19236,N_19775);
nand U20096 (N_20096,N_19840,N_18859);
and U20097 (N_20097,N_18553,N_19075);
nand U20098 (N_20098,N_18841,N_19094);
and U20099 (N_20099,N_19841,N_18454);
xor U20100 (N_20100,N_19502,N_19565);
and U20101 (N_20101,N_18114,N_19516);
or U20102 (N_20102,N_19961,N_19102);
or U20103 (N_20103,N_18484,N_19668);
xnor U20104 (N_20104,N_19941,N_18602);
xnor U20105 (N_20105,N_18072,N_18536);
or U20106 (N_20106,N_19044,N_19868);
or U20107 (N_20107,N_18039,N_18719);
or U20108 (N_20108,N_19992,N_18809);
or U20109 (N_20109,N_19615,N_19524);
nand U20110 (N_20110,N_18976,N_18335);
or U20111 (N_20111,N_19570,N_19991);
nor U20112 (N_20112,N_19793,N_18621);
and U20113 (N_20113,N_18358,N_18656);
and U20114 (N_20114,N_18927,N_19539);
or U20115 (N_20115,N_18344,N_19401);
nor U20116 (N_20116,N_18329,N_18626);
and U20117 (N_20117,N_19168,N_18500);
xnor U20118 (N_20118,N_19374,N_18250);
and U20119 (N_20119,N_19944,N_19419);
xnor U20120 (N_20120,N_19462,N_19945);
nand U20121 (N_20121,N_18771,N_18899);
or U20122 (N_20122,N_18767,N_19292);
and U20123 (N_20123,N_18012,N_18134);
nand U20124 (N_20124,N_18397,N_19030);
and U20125 (N_20125,N_18092,N_19455);
xor U20126 (N_20126,N_19307,N_18121);
xor U20127 (N_20127,N_19005,N_18029);
or U20128 (N_20128,N_18606,N_19380);
nand U20129 (N_20129,N_18081,N_18875);
and U20130 (N_20130,N_18333,N_19787);
and U20131 (N_20131,N_18061,N_18028);
xnor U20132 (N_20132,N_18382,N_19305);
xnor U20133 (N_20133,N_19136,N_18330);
or U20134 (N_20134,N_19974,N_19458);
nand U20135 (N_20135,N_18362,N_18472);
or U20136 (N_20136,N_19616,N_18159);
and U20137 (N_20137,N_18400,N_19686);
xnor U20138 (N_20138,N_19376,N_19015);
or U20139 (N_20139,N_19723,N_19870);
xnor U20140 (N_20140,N_19205,N_19778);
nor U20141 (N_20141,N_18870,N_18543);
and U20142 (N_20142,N_18622,N_18227);
and U20143 (N_20143,N_18014,N_18456);
nand U20144 (N_20144,N_18157,N_19363);
xor U20145 (N_20145,N_19816,N_19536);
xnor U20146 (N_20146,N_18508,N_19371);
xor U20147 (N_20147,N_19020,N_19397);
nand U20148 (N_20148,N_18221,N_19467);
or U20149 (N_20149,N_18783,N_18242);
and U20150 (N_20150,N_19210,N_18119);
xnor U20151 (N_20151,N_19421,N_18449);
and U20152 (N_20152,N_18905,N_19933);
xnor U20153 (N_20153,N_18125,N_18439);
nand U20154 (N_20154,N_18810,N_19009);
nand U20155 (N_20155,N_19268,N_19989);
or U20156 (N_20156,N_18024,N_18800);
xor U20157 (N_20157,N_19406,N_19905);
nand U20158 (N_20158,N_19103,N_19395);
xnor U20159 (N_20159,N_19348,N_18805);
or U20160 (N_20160,N_18846,N_19695);
or U20161 (N_20161,N_18234,N_19389);
and U20162 (N_20162,N_18582,N_18201);
nor U20163 (N_20163,N_19879,N_18297);
xor U20164 (N_20164,N_19771,N_19826);
nor U20165 (N_20165,N_18139,N_18438);
or U20166 (N_20166,N_18331,N_19275);
nand U20167 (N_20167,N_19373,N_18924);
and U20168 (N_20168,N_18527,N_19797);
or U20169 (N_20169,N_19664,N_18737);
or U20170 (N_20170,N_18294,N_18914);
nor U20171 (N_20171,N_19980,N_18908);
xnor U20172 (N_20172,N_19854,N_18723);
xor U20173 (N_20173,N_18801,N_19909);
and U20174 (N_20174,N_18760,N_18078);
nand U20175 (N_20175,N_19112,N_19682);
nand U20176 (N_20176,N_19962,N_19317);
and U20177 (N_20177,N_19514,N_18420);
nor U20178 (N_20178,N_18146,N_19556);
or U20179 (N_20179,N_19466,N_18929);
xor U20180 (N_20180,N_19106,N_19786);
or U20181 (N_20181,N_19320,N_19067);
and U20182 (N_20182,N_19589,N_18059);
nand U20183 (N_20183,N_18967,N_19429);
and U20184 (N_20184,N_19433,N_18698);
nand U20185 (N_20185,N_18148,N_19544);
or U20186 (N_20186,N_18003,N_18388);
and U20187 (N_20187,N_19801,N_19898);
xnor U20188 (N_20188,N_18555,N_19935);
nand U20189 (N_20189,N_18799,N_18475);
and U20190 (N_20190,N_18752,N_18701);
or U20191 (N_20191,N_18883,N_19864);
and U20192 (N_20192,N_18528,N_18237);
nor U20193 (N_20193,N_18675,N_18444);
and U20194 (N_20194,N_18795,N_18468);
nor U20195 (N_20195,N_19200,N_19762);
nand U20196 (N_20196,N_18983,N_19774);
or U20197 (N_20197,N_19937,N_18540);
nor U20198 (N_20198,N_18441,N_19621);
nor U20199 (N_20199,N_19865,N_19652);
nor U20200 (N_20200,N_18650,N_18267);
nor U20201 (N_20201,N_19733,N_19956);
nor U20202 (N_20202,N_18046,N_18187);
xnor U20203 (N_20203,N_19875,N_18601);
and U20204 (N_20204,N_19129,N_18969);
nand U20205 (N_20205,N_18285,N_19157);
and U20206 (N_20206,N_18097,N_18594);
nor U20207 (N_20207,N_19079,N_18241);
and U20208 (N_20208,N_18586,N_19789);
xor U20209 (N_20209,N_19704,N_18863);
nand U20210 (N_20210,N_18755,N_18797);
nand U20211 (N_20211,N_18686,N_18431);
and U20212 (N_20212,N_19390,N_18403);
xnor U20213 (N_20213,N_19926,N_18616);
nor U20214 (N_20214,N_18746,N_19580);
nand U20215 (N_20215,N_19356,N_18506);
nor U20216 (N_20216,N_18986,N_19585);
nor U20217 (N_20217,N_18270,N_19553);
or U20218 (N_20218,N_19193,N_18259);
and U20219 (N_20219,N_18233,N_18624);
xor U20220 (N_20220,N_18643,N_18340);
nand U20221 (N_20221,N_18142,N_19309);
and U20222 (N_20222,N_18672,N_18171);
nor U20223 (N_20223,N_19831,N_19179);
nor U20224 (N_20224,N_19147,N_19700);
nor U20225 (N_20225,N_18440,N_18896);
and U20226 (N_20226,N_18186,N_18775);
and U20227 (N_20227,N_18396,N_19583);
or U20228 (N_20228,N_18652,N_18090);
nor U20229 (N_20229,N_19345,N_19927);
nand U20230 (N_20230,N_19527,N_19784);
nand U20231 (N_20231,N_18036,N_19832);
or U20232 (N_20232,N_18745,N_19542);
or U20233 (N_20233,N_19567,N_19680);
xnor U20234 (N_20234,N_19427,N_19358);
nor U20235 (N_20235,N_19163,N_18094);
xor U20236 (N_20236,N_19873,N_18796);
nor U20237 (N_20237,N_19963,N_18079);
nor U20238 (N_20238,N_19858,N_19754);
and U20239 (N_20239,N_18113,N_19245);
nor U20240 (N_20240,N_19976,N_19326);
nand U20241 (N_20241,N_18618,N_19319);
or U20242 (N_20242,N_19874,N_19468);
nor U20243 (N_20243,N_19986,N_18903);
and U20244 (N_20244,N_19773,N_18052);
xor U20245 (N_20245,N_19611,N_19648);
or U20246 (N_20246,N_18517,N_18944);
and U20247 (N_20247,N_19642,N_18038);
and U20248 (N_20248,N_19535,N_19714);
xnor U20249 (N_20249,N_18100,N_18595);
nor U20250 (N_20250,N_18501,N_19384);
nor U20251 (N_20251,N_18699,N_18984);
xnor U20252 (N_20252,N_18276,N_18430);
nor U20253 (N_20253,N_19501,N_18713);
or U20254 (N_20254,N_18286,N_19850);
and U20255 (N_20255,N_19772,N_18960);
xor U20256 (N_20256,N_19867,N_18000);
xor U20257 (N_20257,N_19125,N_18940);
nor U20258 (N_20258,N_19369,N_18450);
nor U20259 (N_20259,N_19685,N_18434);
or U20260 (N_20260,N_18902,N_19981);
and U20261 (N_20261,N_18483,N_18426);
or U20262 (N_20262,N_19949,N_18488);
or U20263 (N_20263,N_19448,N_19053);
and U20264 (N_20264,N_18295,N_19222);
and U20265 (N_20265,N_18510,N_19391);
nand U20266 (N_20266,N_19054,N_19285);
nor U20267 (N_20267,N_18402,N_18998);
xor U20268 (N_20268,N_19813,N_18349);
xnor U20269 (N_20269,N_18739,N_18123);
nor U20270 (N_20270,N_19444,N_18551);
nand U20271 (N_20271,N_18812,N_18145);
xor U20272 (N_20272,N_19609,N_18715);
and U20273 (N_20273,N_19192,N_18682);
nand U20274 (N_20274,N_18044,N_18939);
nor U20275 (N_20275,N_18088,N_18677);
nand U20276 (N_20276,N_18222,N_19119);
nand U20277 (N_20277,N_18704,N_18631);
nand U20278 (N_20278,N_18872,N_19294);
nor U20279 (N_20279,N_18893,N_19650);
nand U20280 (N_20280,N_18418,N_19159);
nor U20281 (N_20281,N_18126,N_19296);
xnor U20282 (N_20282,N_18164,N_19509);
nand U20283 (N_20283,N_19148,N_18619);
or U20284 (N_20284,N_19970,N_19493);
nor U20285 (N_20285,N_19953,N_18136);
nand U20286 (N_20286,N_18152,N_19212);
and U20287 (N_20287,N_18918,N_18740);
or U20288 (N_20288,N_19794,N_18684);
and U20289 (N_20289,N_19906,N_18758);
nand U20290 (N_20290,N_19631,N_19249);
or U20291 (N_20291,N_18098,N_19213);
nor U20292 (N_20292,N_18592,N_18596);
xor U20293 (N_20293,N_19730,N_19080);
or U20294 (N_20294,N_19582,N_19569);
nor U20295 (N_20295,N_19900,N_19392);
and U20296 (N_20296,N_19798,N_18963);
xor U20297 (N_20297,N_18292,N_19386);
nor U20298 (N_20298,N_18769,N_18082);
xor U20299 (N_20299,N_19880,N_19388);
or U20300 (N_20300,N_19201,N_19821);
nand U20301 (N_20301,N_19368,N_19495);
nand U20302 (N_20302,N_18253,N_18741);
nand U20303 (N_20303,N_18135,N_18694);
nor U20304 (N_20304,N_19247,N_18254);
and U20305 (N_20305,N_18542,N_18847);
nand U20306 (N_20306,N_19634,N_19671);
xnor U20307 (N_20307,N_19143,N_19693);
xor U20308 (N_20308,N_19532,N_18577);
and U20309 (N_20309,N_18585,N_19046);
and U20310 (N_20310,N_18336,N_19526);
nor U20311 (N_20311,N_18005,N_18026);
xor U20312 (N_20312,N_19060,N_19871);
or U20313 (N_20313,N_19341,N_18830);
or U20314 (N_20314,N_18283,N_18009);
nand U20315 (N_20315,N_19325,N_19712);
and U20316 (N_20316,N_19844,N_19554);
nor U20317 (N_20317,N_19123,N_18556);
nor U20318 (N_20318,N_19441,N_19779);
and U20319 (N_20319,N_18230,N_19960);
and U20320 (N_20320,N_19132,N_18369);
xnor U20321 (N_20321,N_19781,N_18166);
or U20322 (N_20322,N_18572,N_18188);
nor U20323 (N_20323,N_18632,N_18666);
nor U20324 (N_20324,N_19515,N_18563);
nor U20325 (N_20325,N_19050,N_19039);
or U20326 (N_20326,N_19920,N_19450);
xor U20327 (N_20327,N_18916,N_18047);
or U20328 (N_20328,N_18174,N_18900);
and U20329 (N_20329,N_18321,N_18371);
nor U20330 (N_20330,N_19977,N_19415);
or U20331 (N_20331,N_18310,N_19291);
and U20332 (N_20332,N_18569,N_19313);
xor U20333 (N_20333,N_19199,N_19601);
and U20334 (N_20334,N_18568,N_19156);
or U20335 (N_20335,N_19658,N_19412);
nand U20336 (N_20336,N_19560,N_19281);
or U20337 (N_20337,N_18433,N_19280);
and U20338 (N_20338,N_18163,N_19521);
xnor U20339 (N_20339,N_18573,N_18062);
nor U20340 (N_20340,N_18118,N_18854);
nand U20341 (N_20341,N_19810,N_19936);
nor U20342 (N_20342,N_18101,N_18392);
or U20343 (N_20343,N_19724,N_18832);
nor U20344 (N_20344,N_19983,N_18469);
and U20345 (N_20345,N_18653,N_19796);
and U20346 (N_20346,N_18819,N_18466);
xor U20347 (N_20347,N_18067,N_19253);
nand U20348 (N_20348,N_18001,N_19154);
nor U20349 (N_20349,N_18202,N_18181);
xor U20350 (N_20350,N_18584,N_18476);
and U20351 (N_20351,N_18603,N_19916);
nor U20352 (N_20352,N_19606,N_18949);
and U20353 (N_20353,N_18974,N_18971);
or U20354 (N_20354,N_18647,N_18491);
nor U20355 (N_20355,N_19891,N_19932);
nand U20356 (N_20356,N_18890,N_19968);
nor U20357 (N_20357,N_19500,N_19021);
nand U20358 (N_20358,N_18935,N_18932);
or U20359 (N_20359,N_18793,N_18977);
nor U20360 (N_20360,N_19508,N_18887);
or U20361 (N_20361,N_19645,N_19321);
and U20362 (N_20362,N_18884,N_18185);
nor U20363 (N_20363,N_18025,N_19463);
xnor U20364 (N_20364,N_18509,N_19528);
nand U20365 (N_20365,N_18002,N_19165);
and U20366 (N_20366,N_19114,N_18375);
nor U20367 (N_20367,N_18610,N_19476);
or U20368 (N_20368,N_18228,N_18892);
and U20369 (N_20369,N_19988,N_19452);
nand U20370 (N_20370,N_19910,N_18667);
nand U20371 (N_20371,N_19474,N_19003);
and U20372 (N_20372,N_18050,N_19950);
nor U20373 (N_20373,N_18351,N_18838);
and U20374 (N_20374,N_18301,N_19061);
and U20375 (N_20375,N_19849,N_19577);
nor U20376 (N_20376,N_18504,N_18346);
nand U20377 (N_20377,N_19545,N_18116);
and U20378 (N_20378,N_18258,N_19259);
and U20379 (N_20379,N_18850,N_19482);
xnor U20380 (N_20380,N_19940,N_19739);
nor U20381 (N_20381,N_18693,N_19994);
xnor U20382 (N_20382,N_18879,N_18395);
nor U20383 (N_20383,N_18590,N_19698);
or U20384 (N_20384,N_18498,N_19166);
nor U20385 (N_20385,N_18750,N_18525);
and U20386 (N_20386,N_18165,N_18379);
or U20387 (N_20387,N_19622,N_19034);
xnor U20388 (N_20388,N_19791,N_18593);
xor U20389 (N_20389,N_19214,N_19770);
xor U20390 (N_20390,N_18235,N_19109);
and U20391 (N_20391,N_19057,N_19711);
or U20392 (N_20392,N_18209,N_19603);
or U20393 (N_20393,N_18814,N_19265);
or U20394 (N_20394,N_19904,N_19161);
and U20395 (N_20395,N_19487,N_18353);
or U20396 (N_20396,N_18337,N_18298);
nand U20397 (N_20397,N_19365,N_19261);
xor U20398 (N_20398,N_18309,N_18749);
xor U20399 (N_20399,N_18792,N_19279);
nand U20400 (N_20400,N_18754,N_19518);
or U20401 (N_20401,N_19149,N_18881);
nor U20402 (N_20402,N_18315,N_19566);
and U20403 (N_20403,N_18304,N_19598);
xor U20404 (N_20404,N_19602,N_19099);
or U20405 (N_20405,N_19113,N_18579);
nand U20406 (N_20406,N_19899,N_18788);
and U20407 (N_20407,N_19056,N_18711);
xor U20408 (N_20408,N_19885,N_18284);
or U20409 (N_20409,N_18414,N_19651);
and U20410 (N_20410,N_18807,N_18535);
xor U20411 (N_20411,N_18183,N_18858);
nand U20412 (N_20412,N_19803,N_19531);
and U20413 (N_20413,N_18589,N_19845);
xnor U20414 (N_20414,N_19613,N_18913);
nand U20415 (N_20415,N_19997,N_18687);
xor U20416 (N_20416,N_19869,N_18751);
or U20417 (N_20417,N_18708,N_18886);
nor U20418 (N_20418,N_18182,N_18548);
and U20419 (N_20419,N_19111,N_19298);
xnor U20420 (N_20420,N_18175,N_18053);
and U20421 (N_20421,N_19923,N_19633);
nand U20422 (N_20422,N_18607,N_18495);
nand U20423 (N_20423,N_19599,N_18609);
nor U20424 (N_20424,N_19207,N_18505);
and U20425 (N_20425,N_18410,N_18419);
nand U20426 (N_20426,N_19878,N_19763);
xor U20427 (N_20427,N_18566,N_18280);
xor U20428 (N_20428,N_19048,N_19297);
or U20429 (N_20429,N_18075,N_18868);
nand U20430 (N_20430,N_18720,N_19353);
nand U20431 (N_20431,N_18432,N_18343);
nor U20432 (N_20432,N_18764,N_18023);
nor U20433 (N_20433,N_18654,N_18096);
xnor U20434 (N_20434,N_19262,N_18831);
and U20435 (N_20435,N_18367,N_18318);
or U20436 (N_20436,N_19133,N_18122);
nor U20437 (N_20437,N_18459,N_18218);
and U20438 (N_20438,N_18839,N_18011);
or U20439 (N_20439,N_18030,N_18137);
and U20440 (N_20440,N_18453,N_18599);
or U20441 (N_20441,N_18487,N_19115);
or U20442 (N_20442,N_18707,N_18086);
nand U20443 (N_20443,N_19817,N_19459);
and U20444 (N_20444,N_18837,N_19335);
or U20445 (N_20445,N_18635,N_18390);
nand U20446 (N_20446,N_18354,N_19336);
nand U20447 (N_20447,N_18637,N_19830);
and U20448 (N_20448,N_18808,N_19533);
xor U20449 (N_20449,N_19503,N_19035);
nor U20450 (N_20450,N_19756,N_19672);
nand U20451 (N_20451,N_18048,N_19145);
nand U20452 (N_20452,N_19120,N_19211);
or U20453 (N_20453,N_18184,N_18574);
xor U20454 (N_20454,N_18778,N_19209);
nand U20455 (N_20455,N_19027,N_19834);
or U20456 (N_20456,N_19065,N_18945);
and U20457 (N_20457,N_18350,N_18785);
and U20458 (N_20458,N_19715,N_19839);
and U20459 (N_20459,N_18981,N_18827);
xor U20460 (N_20460,N_19654,N_19894);
xor U20461 (N_20461,N_19022,N_18065);
nand U20462 (N_20462,N_18676,N_19096);
and U20463 (N_20463,N_19918,N_18168);
or U20464 (N_20464,N_18368,N_18085);
or U20465 (N_20465,N_18926,N_19759);
or U20466 (N_20466,N_18198,N_18702);
nor U20467 (N_20467,N_19130,N_18912);
nand U20468 (N_20468,N_18730,N_18144);
nor U20469 (N_20469,N_18172,N_18133);
nor U20470 (N_20470,N_18147,N_18757);
nor U20471 (N_20471,N_18774,N_19965);
xor U20472 (N_20472,N_18732,N_19568);
nand U20473 (N_20473,N_19859,N_18532);
xor U20474 (N_20474,N_18669,N_18091);
xor U20475 (N_20475,N_18364,N_19819);
xor U20476 (N_20476,N_18398,N_19188);
nor U20477 (N_20477,N_19699,N_18107);
or U20478 (N_20478,N_19001,N_18493);
and U20479 (N_20479,N_18851,N_18010);
xnor U20480 (N_20480,N_19990,N_19855);
nand U20481 (N_20481,N_19355,N_19344);
and U20482 (N_20482,N_18102,N_18867);
nand U20483 (N_20483,N_19558,N_19354);
nor U20484 (N_20484,N_18816,N_18404);
or U20485 (N_20485,N_18953,N_19753);
nand U20486 (N_20486,N_19471,N_18683);
nor U20487 (N_20487,N_18220,N_18461);
xnor U20488 (N_20488,N_19825,N_19352);
or U20489 (N_20489,N_19413,N_18246);
xnor U20490 (N_20490,N_18756,N_18733);
nor U20491 (N_20491,N_19971,N_18215);
nor U20492 (N_20492,N_18539,N_19541);
and U20493 (N_20493,N_18997,N_19480);
or U20494 (N_20494,N_18964,N_19447);
nand U20495 (N_20495,N_19311,N_19042);
or U20496 (N_20496,N_18972,N_19543);
xor U20497 (N_20497,N_19812,N_18710);
or U20498 (N_20498,N_19641,N_18547);
or U20499 (N_20499,N_18176,N_19958);
xor U20500 (N_20500,N_18597,N_18600);
nor U20501 (N_20501,N_18192,N_19972);
nor U20502 (N_20502,N_19451,N_18485);
nand U20503 (N_20503,N_19860,N_18679);
nor U20504 (N_20504,N_19176,N_19638);
nand U20505 (N_20505,N_19607,N_18781);
xor U20506 (N_20506,N_19827,N_19593);
or U20507 (N_20507,N_18381,N_19547);
nand U20508 (N_20508,N_19551,N_18040);
nor U20509 (N_20509,N_18734,N_19187);
or U20510 (N_20510,N_19729,N_18214);
xor U20511 (N_20511,N_18243,N_19721);
nor U20512 (N_20512,N_19943,N_18264);
nand U20513 (N_20513,N_18938,N_19036);
and U20514 (N_20514,N_18538,N_18762);
nand U20515 (N_20515,N_19497,N_18520);
or U20516 (N_20516,N_19456,N_18503);
or U20517 (N_20517,N_19019,N_19982);
and U20518 (N_20518,N_19924,N_19726);
nor U20519 (N_20519,N_19457,N_19489);
xor U20520 (N_20520,N_18992,N_19673);
and U20521 (N_20521,N_19382,N_18019);
nor U20522 (N_20522,N_18356,N_18692);
xnor U20523 (N_20523,N_18985,N_19795);
nand U20524 (N_20524,N_18691,N_19024);
or U20525 (N_20525,N_19747,N_19866);
nand U20526 (N_20526,N_18999,N_18833);
nor U20527 (N_20527,N_19186,N_19150);
nand U20528 (N_20528,N_18885,N_18623);
and U20529 (N_20529,N_19954,N_19220);
or U20530 (N_20530,N_19520,N_18366);
xor U20531 (N_20531,N_18968,N_18399);
xnor U20532 (N_20532,N_18614,N_19446);
nor U20533 (N_20533,N_18815,N_19481);
nor U20534 (N_20534,N_18408,N_18413);
and U20535 (N_20535,N_19381,N_18864);
xnor U20536 (N_20536,N_19807,N_18423);
nor U20537 (N_20537,N_19512,N_19863);
nand U20538 (N_20538,N_18260,N_18127);
or U20539 (N_20539,N_19829,N_18583);
nand U20540 (N_20540,N_19725,N_19635);
and U20541 (N_20541,N_19235,N_18817);
xor U20542 (N_20542,N_19752,N_19555);
nor U20543 (N_20543,N_19818,N_19461);
or U20544 (N_20544,N_18124,N_19256);
xor U20545 (N_20545,N_19851,N_18961);
xor U20546 (N_20546,N_18236,N_18877);
and U20547 (N_20547,N_19434,N_18575);
xor U20548 (N_20548,N_18213,N_19107);
or U20549 (N_20549,N_19511,N_18777);
and U20550 (N_20550,N_18249,N_19271);
nor U20551 (N_20551,N_19575,N_19930);
and U20552 (N_20552,N_19669,N_19189);
or U20553 (N_20553,N_18013,N_19814);
xor U20554 (N_20554,N_18636,N_19529);
nand U20555 (N_20555,N_18149,N_19999);
nor U20556 (N_20556,N_18045,N_19969);
xnor U20557 (N_20557,N_19911,N_18306);
and U20558 (N_20558,N_19314,N_18822);
or U20559 (N_20559,N_19004,N_19240);
nor U20560 (N_20560,N_19612,N_19473);
nand U20561 (N_20561,N_19063,N_18518);
nor U20562 (N_20562,N_18223,N_19626);
nand U20563 (N_20563,N_19697,N_19966);
nand U20564 (N_20564,N_19137,N_19677);
nor U20565 (N_20565,N_18161,N_18244);
and U20566 (N_20566,N_18020,N_19780);
or U20567 (N_20567,N_18980,N_19435);
xor U20568 (N_20568,N_18587,N_19744);
or U20569 (N_20569,N_19403,N_19361);
xnor U20570 (N_20570,N_19416,N_19710);
nand U20571 (N_20571,N_18735,N_19226);
nand U20572 (N_20572,N_19696,N_19548);
xnor U20573 (N_20573,N_18041,N_19884);
xor U20574 (N_20574,N_19140,N_18588);
or U20575 (N_20575,N_19173,N_18191);
nor U20576 (N_20576,N_18070,N_19234);
nand U20577 (N_20577,N_19996,N_19219);
and U20578 (N_20578,N_18282,N_19040);
xor U20579 (N_20579,N_19597,N_19206);
xnor U20580 (N_20580,N_19026,N_19939);
nor U20581 (N_20581,N_18848,N_19978);
and U20582 (N_20582,N_18768,N_18727);
nand U20583 (N_20583,N_18763,N_18557);
and U20584 (N_20584,N_18917,N_19300);
nand U20585 (N_20585,N_18678,N_18377);
nand U20586 (N_20586,N_18018,N_18004);
xor U20587 (N_20587,N_19636,N_18391);
or U20588 (N_20588,N_19494,N_19233);
and U20589 (N_20589,N_18671,N_19089);
nor U20590 (N_20590,N_19995,N_18743);
nor U20591 (N_20591,N_19504,N_19066);
and U20592 (N_20592,N_19139,N_18950);
nand U20593 (N_20593,N_18376,N_18314);
nor U20594 (N_20594,N_18957,N_19153);
nor U20595 (N_20595,N_18860,N_18296);
and U20596 (N_20596,N_19128,N_19052);
nand U20597 (N_20597,N_19470,N_19946);
xor U20598 (N_20598,N_19180,N_19237);
nor U20599 (N_20599,N_19045,N_18316);
nor U20600 (N_20600,N_18639,N_19393);
xor U20601 (N_20601,N_19334,N_18869);
and U20602 (N_20602,N_19857,N_19550);
nand U20603 (N_20603,N_18513,N_19717);
xor U20604 (N_20604,N_18370,N_18158);
or U20605 (N_20605,N_19666,N_18611);
xor U20606 (N_20606,N_18729,N_19006);
xnor U20607 (N_20607,N_19670,N_19479);
xor U20608 (N_20608,N_19823,N_19267);
nand U20609 (N_20609,N_18455,N_19404);
and U20610 (N_20610,N_19323,N_19769);
or U20611 (N_20611,N_18111,N_19047);
or U20612 (N_20612,N_19284,N_19190);
nand U20613 (N_20613,N_18578,N_18591);
and U20614 (N_20614,N_19546,N_19731);
and U20615 (N_20615,N_19984,N_18412);
nand U20616 (N_20616,N_18728,N_18338);
nor U20617 (N_20617,N_19908,N_19692);
xor U20618 (N_20618,N_19892,N_19258);
nor U20619 (N_20619,N_18109,N_18470);
and U20620 (N_20620,N_19925,N_19847);
nand U20621 (N_20621,N_18066,N_19571);
or U20622 (N_20622,N_18840,N_18897);
nor U20623 (N_20623,N_19485,N_18042);
xor U20624 (N_20624,N_18263,N_19092);
and U20625 (N_20625,N_19318,N_19007);
or U20626 (N_20626,N_18332,N_18826);
nand U20627 (N_20627,N_18919,N_18552);
xor U20628 (N_20628,N_18975,N_18630);
or U20629 (N_20629,N_18153,N_18959);
nor U20630 (N_20630,N_19785,N_18255);
and U20631 (N_20631,N_19322,N_18571);
nor U20632 (N_20632,N_18965,N_18105);
xnor U20633 (N_20633,N_19351,N_19152);
or U20634 (N_20634,N_19276,N_19064);
nand U20635 (N_20635,N_18804,N_19242);
and U20636 (N_20636,N_18979,N_18507);
nand U20637 (N_20637,N_19738,N_19088);
nand U20638 (N_20638,N_18194,N_18196);
and U20639 (N_20639,N_19805,N_19661);
and U20640 (N_20640,N_18565,N_18894);
or U20641 (N_20641,N_19225,N_19815);
nor U20642 (N_20642,N_18084,N_18064);
nor U20643 (N_20643,N_19216,N_19557);
nor U20644 (N_20644,N_19749,N_19385);
and U20645 (N_20645,N_18790,N_18843);
nor U20646 (N_20646,N_19848,N_18891);
nor U20647 (N_20647,N_19660,N_19217);
xor U20648 (N_20648,N_19587,N_19572);
nand U20649 (N_20649,N_18617,N_19239);
or U20650 (N_20650,N_19185,N_19160);
nor U20651 (N_20651,N_18560,N_19655);
nand U20652 (N_20652,N_18931,N_18406);
nor U20653 (N_20653,N_19734,N_19198);
nand U20654 (N_20654,N_19248,N_18644);
nand U20655 (N_20655,N_19405,N_19073);
nand U20656 (N_20656,N_19414,N_18776);
nand U20657 (N_20657,N_19667,N_18888);
nor U20658 (N_20658,N_18417,N_18681);
and U20659 (N_20659,N_18995,N_19178);
nor U20660 (N_20660,N_19410,N_18856);
nor U20661 (N_20661,N_18274,N_18862);
nand U20662 (N_20662,N_18526,N_19312);
nor U20663 (N_20663,N_19306,N_19424);
nor U20664 (N_20664,N_19630,N_19720);
and U20665 (N_20665,N_18256,N_19408);
nand U20666 (N_20666,N_19656,N_18268);
xnor U20667 (N_20667,N_18718,N_18580);
nor U20668 (N_20668,N_18389,N_18197);
nand U20669 (N_20669,N_19229,N_19486);
or U20670 (N_20670,N_19090,N_19496);
nor U20671 (N_20671,N_18920,N_19093);
xnor U20672 (N_20672,N_19843,N_19295);
nand U20673 (N_20673,N_18641,N_19460);
or U20674 (N_20674,N_19912,N_18811);
xnor U20675 (N_20675,N_19523,N_18320);
and U20676 (N_20676,N_18287,N_19806);
or U20677 (N_20677,N_18195,N_18180);
nand U20678 (N_20678,N_18035,N_19562);
nand U20679 (N_20679,N_19728,N_18844);
xnor U20680 (N_20680,N_18823,N_18357);
and U20681 (N_20681,N_18205,N_19888);
or U20682 (N_20682,N_18224,N_18523);
nor U20683 (N_20683,N_19398,N_19084);
or U20684 (N_20684,N_19316,N_19907);
xor U20685 (N_20685,N_18372,N_19431);
or U20686 (N_20686,N_19366,N_19653);
and U20687 (N_20687,N_18232,N_18057);
or U20688 (N_20688,N_19768,N_19967);
or U20689 (N_20689,N_18017,N_19915);
and U20690 (N_20690,N_19131,N_18829);
nand U20691 (N_20691,N_18060,N_18921);
xnor U20692 (N_20692,N_18464,N_18269);
xor U20693 (N_20693,N_19877,N_18519);
and U20694 (N_20694,N_18080,N_18334);
xor U20695 (N_20695,N_19505,N_19931);
or U20696 (N_20696,N_19921,N_19250);
or U20697 (N_20697,N_19407,N_18341);
nand U20698 (N_20698,N_18360,N_18697);
xor U20699 (N_20699,N_18303,N_19574);
nand U20700 (N_20700,N_18514,N_19707);
nor U20701 (N_20701,N_19087,N_19679);
or U20702 (N_20702,N_18231,N_19765);
nor U20703 (N_20703,N_19627,N_19913);
nand U20704 (N_20704,N_19674,N_19304);
and U20705 (N_20705,N_18291,N_18445);
xor U20706 (N_20706,N_18533,N_18348);
nor U20707 (N_20707,N_19155,N_18825);
and U20708 (N_20708,N_18428,N_19328);
xor U20709 (N_20709,N_18008,N_19342);
nand U20710 (N_20710,N_19951,N_18836);
xnor U20711 (N_20711,N_18907,N_18895);
xnor U20712 (N_20712,N_19938,N_18293);
nor U20713 (N_20713,N_19287,N_18873);
and U20714 (N_20714,N_19998,N_19432);
and U20715 (N_20715,N_18212,N_18721);
xor U20716 (N_20716,N_19478,N_18261);
or U20717 (N_20717,N_18661,N_19303);
or U20718 (N_20718,N_19332,N_19104);
and U20719 (N_20719,N_19031,N_19083);
and U20720 (N_20720,N_18007,N_19167);
or U20721 (N_20721,N_19118,N_18933);
xor U20722 (N_20722,N_18435,N_19333);
nor U20723 (N_20723,N_18076,N_18649);
xnor U20724 (N_20724,N_18544,N_19657);
and U20725 (N_20725,N_18628,N_19243);
xor U20726 (N_20726,N_19151,N_19628);
nand U20727 (N_20727,N_19676,N_18529);
xor U20728 (N_20728,N_18629,N_19097);
nor U20729 (N_20729,N_19171,N_19426);
and U20730 (N_20730,N_18657,N_19861);
or U20731 (N_20731,N_18112,N_19889);
nor U20732 (N_20732,N_18955,N_19563);
nand U20733 (N_20733,N_19230,N_18904);
nand U20734 (N_20734,N_19324,N_19055);
and U20735 (N_20735,N_19449,N_19782);
and U20736 (N_20736,N_18736,N_19362);
xor U20737 (N_20737,N_19985,N_19596);
nand U20738 (N_20738,N_19051,N_18906);
or U20739 (N_20739,N_18021,N_18211);
or U20740 (N_20740,N_18324,N_19746);
xor U20741 (N_20741,N_19223,N_19379);
nor U20742 (N_20742,N_19231,N_19709);
and U20743 (N_20743,N_18499,N_18407);
nor U20744 (N_20744,N_18608,N_18141);
nand U20745 (N_20745,N_19605,N_18068);
xnor U20746 (N_20746,N_19922,N_19204);
nand U20747 (N_20747,N_18462,N_18150);
and U20748 (N_20748,N_18522,N_18901);
xor U20749 (N_20749,N_19331,N_18813);
xnor U20750 (N_20750,N_19975,N_18006);
or U20751 (N_20751,N_18446,N_19987);
xnor U20752 (N_20752,N_18865,N_18347);
nand U20753 (N_20753,N_19691,N_18668);
nand U20754 (N_20754,N_18199,N_18058);
or U20755 (N_20755,N_19110,N_19792);
or U20756 (N_20756,N_18219,N_19164);
and U20757 (N_20757,N_19174,N_18680);
xor U20758 (N_20758,N_18828,N_18273);
xor U20759 (N_20759,N_19367,N_19684);
xnor U20760 (N_20760,N_19043,N_18857);
nor U20761 (N_20761,N_18087,N_18173);
and U20762 (N_20762,N_18633,N_19745);
or U20763 (N_20763,N_18770,N_19347);
and U20764 (N_20764,N_19808,N_19000);
nor U20765 (N_20765,N_19586,N_18442);
xor U20766 (N_20766,N_18530,N_18322);
xnor U20767 (N_20767,N_18447,N_18251);
nor U20768 (N_20768,N_18069,N_18982);
xnor U20769 (N_20769,N_19513,N_18063);
nor U20770 (N_20770,N_19881,N_18465);
and U20771 (N_20771,N_19683,N_19735);
and U20772 (N_20772,N_19282,N_18882);
nor U20773 (N_20773,N_19454,N_18991);
or U20774 (N_20774,N_19302,N_18724);
xnor U20775 (N_20775,N_19886,N_18787);
nand U20776 (N_20776,N_18747,N_18238);
nand U20777 (N_20777,N_19678,N_19538);
xor U20778 (N_20778,N_19802,N_18272);
or U20779 (N_20779,N_18695,N_18167);
nand U20780 (N_20780,N_18759,N_18128);
or U20781 (N_20781,N_19012,N_18786);
xnor U20782 (N_20782,N_18037,N_18541);
nor U20783 (N_20783,N_19890,N_18662);
xnor U20784 (N_20784,N_18989,N_18558);
xnor U20785 (N_20785,N_18262,N_19062);
nand U20786 (N_20786,N_19477,N_18073);
or U20787 (N_20787,N_18549,N_19014);
or U20788 (N_20788,N_19625,N_19028);
nand U20789 (N_20789,N_19269,N_19278);
or U20790 (N_20790,N_18110,N_19041);
or U20791 (N_20791,N_19162,N_19581);
or U20792 (N_20792,N_19594,N_19049);
and U20793 (N_20793,N_18473,N_19440);
nor U20794 (N_20794,N_19608,N_19732);
or U20795 (N_20795,N_18784,N_18421);
xnor U20796 (N_20796,N_19838,N_18803);
nor U20797 (N_20797,N_18467,N_18210);
nand U20798 (N_20798,N_18031,N_19264);
or U20799 (N_20799,N_18562,N_19288);
and U20800 (N_20800,N_19409,N_18206);
and U20801 (N_20801,N_19172,N_19887);
nand U20802 (N_20802,N_19360,N_19038);
nand U20803 (N_20803,N_18361,N_19127);
nor U20804 (N_20804,N_19286,N_18022);
and U20805 (N_20805,N_19375,N_18422);
and U20806 (N_20806,N_18634,N_19629);
nand U20807 (N_20807,N_18326,N_18425);
nor U20808 (N_20808,N_18673,N_19343);
xnor U20809 (N_20809,N_19430,N_19082);
nor U20810 (N_20810,N_18302,N_19108);
or U20811 (N_20811,N_19134,N_19246);
or U20812 (N_20812,N_19105,N_18871);
nor U20813 (N_20813,N_19018,N_18852);
nor U20814 (N_20814,N_18394,N_18937);
nand U20815 (N_20815,N_19646,N_18478);
nor U20816 (N_20816,N_19301,N_19919);
xor U20817 (N_20817,N_19703,N_19475);
or U20818 (N_20818,N_18889,N_18325);
or U20819 (N_20819,N_19330,N_18311);
xnor U20820 (N_20820,N_19100,N_18190);
xor U20821 (N_20821,N_19272,N_18208);
or U20822 (N_20822,N_18275,N_19252);
nand U20823 (N_20823,N_19400,N_19071);
and U20824 (N_20824,N_18909,N_19078);
nor U20825 (N_20825,N_18178,N_19126);
and U20826 (N_20826,N_19091,N_19758);
nand U20827 (N_20827,N_18103,N_19689);
nor U20828 (N_20828,N_19069,N_18615);
nand U20829 (N_20829,N_18531,N_18089);
or U20830 (N_20830,N_18359,N_18561);
xnor U20831 (N_20831,N_19116,N_18416);
and U20832 (N_20832,N_19420,N_19525);
or U20833 (N_20833,N_18162,N_19530);
and U20834 (N_20834,N_19013,N_18570);
xor U20835 (N_20835,N_18193,N_18928);
and U20836 (N_20836,N_19142,N_19722);
nand U20837 (N_20837,N_19701,N_18384);
nor U20838 (N_20838,N_18365,N_19169);
or U20839 (N_20839,N_19370,N_19751);
nor U20840 (N_20840,N_18427,N_18780);
nand U20841 (N_20841,N_18380,N_19350);
nand U20842 (N_20842,N_19076,N_18225);
nor U20843 (N_20843,N_19241,N_19934);
xor U20844 (N_20844,N_18709,N_18794);
and U20845 (N_20845,N_18378,N_18327);
nand U20846 (N_20846,N_19649,N_18725);
nor U20847 (N_20847,N_18537,N_19761);
or U20848 (N_20848,N_19614,N_18798);
xor U20849 (N_20849,N_19428,N_19469);
or U20850 (N_20850,N_19492,N_19964);
nor U20851 (N_20851,N_18490,N_18806);
and U20852 (N_20852,N_19095,N_18083);
nand U20853 (N_20853,N_18744,N_18437);
nand U20854 (N_20854,N_18132,N_18373);
xor U20855 (N_20855,N_19647,N_18954);
xor U20856 (N_20856,N_19842,N_18941);
or U20857 (N_20857,N_18824,N_19820);
nor U20858 (N_20858,N_18387,N_19016);
nor U20859 (N_20859,N_18471,N_18791);
nand U20860 (N_20860,N_19183,N_18648);
or U20861 (N_20861,N_19327,N_18117);
nor U20862 (N_20862,N_19659,N_19266);
and U20863 (N_20863,N_18257,N_18934);
nor U20864 (N_20864,N_18313,N_18567);
nor U20865 (N_20865,N_18789,N_18613);
nand U20866 (N_20866,N_19442,N_18460);
nor U20867 (N_20867,N_18106,N_18761);
and U20868 (N_20868,N_18405,N_19783);
nor U20869 (N_20869,N_19718,N_18550);
or U20870 (N_20870,N_19578,N_19914);
nor U20871 (N_20871,N_19453,N_19979);
or U20872 (N_20872,N_19058,N_19617);
nand U20873 (N_20873,N_19836,N_19098);
and U20874 (N_20874,N_18994,N_19025);
and U20875 (N_20875,N_19228,N_18835);
xor U20876 (N_20876,N_18481,N_18512);
nand U20877 (N_20877,N_18317,N_19472);
xor U20878 (N_20878,N_19181,N_19743);
nor U20879 (N_20879,N_19491,N_18095);
or U20880 (N_20880,N_18773,N_19074);
nand U20881 (N_20881,N_19196,N_19736);
nand U20882 (N_20882,N_19008,N_18027);
nor U20883 (N_20883,N_18071,N_19101);
or U20884 (N_20884,N_18670,N_18277);
nor U20885 (N_20885,N_18077,N_18598);
nand U20886 (N_20886,N_19828,N_19639);
nand U20887 (N_20887,N_19364,N_19484);
or U20888 (N_20888,N_19706,N_19215);
and U20889 (N_20889,N_19595,N_19195);
or U20890 (N_20890,N_19443,N_18265);
nand U20891 (N_20891,N_18946,N_19017);
or U20892 (N_20892,N_18074,N_19897);
or U20893 (N_20893,N_19445,N_18866);
and U20894 (N_20894,N_19573,N_18120);
nor U20895 (N_20895,N_18252,N_19224);
or U20896 (N_20896,N_18307,N_19610);
xor U20897 (N_20897,N_18612,N_18229);
xnor U20898 (N_20898,N_18651,N_19846);
xor U20899 (N_20899,N_19121,N_19418);
and U20900 (N_20900,N_18876,N_18474);
xor U20901 (N_20901,N_19788,N_18952);
nor U20902 (N_20902,N_18415,N_19640);
xnor U20903 (N_20903,N_18772,N_19308);
and U20904 (N_20904,N_19588,N_18328);
nor U20905 (N_20905,N_18239,N_18818);
and U20906 (N_20906,N_18479,N_19387);
and U20907 (N_20907,N_18521,N_19394);
and U20908 (N_20908,N_18299,N_19081);
nand U20909 (N_20909,N_19600,N_19085);
nor U20910 (N_20910,N_18559,N_18842);
and U20911 (N_20911,N_19852,N_19824);
and U20912 (N_20912,N_19799,N_19208);
nand U20913 (N_20913,N_18055,N_18463);
nand U20914 (N_20914,N_18627,N_19675);
and U20915 (N_20915,N_19942,N_19010);
or U20916 (N_20916,N_19632,N_18765);
and U20917 (N_20917,N_19191,N_19694);
nor U20918 (N_20918,N_18674,N_18308);
or U20919 (N_20919,N_18305,N_19837);
xor U20920 (N_20920,N_18448,N_18564);
nor U20921 (N_20921,N_19254,N_18312);
nor U20922 (N_20922,N_19177,N_19238);
nand U20923 (N_20923,N_19439,N_19559);
xnor U20924 (N_20924,N_19624,N_18115);
xnor U20925 (N_20925,N_18911,N_19809);
or U20926 (N_20926,N_18726,N_19882);
or U20927 (N_20927,N_19175,N_19790);
and U20928 (N_20928,N_18874,N_18898);
xor U20929 (N_20929,N_19002,N_19182);
xnor U20930 (N_20930,N_19465,N_18861);
nor U20931 (N_20931,N_18820,N_19378);
or U20932 (N_20932,N_18401,N_19576);
xnor U20933 (N_20933,N_19760,N_18104);
or U20934 (N_20934,N_18169,N_18279);
nand U20935 (N_20935,N_19619,N_19561);
nand U20936 (N_20936,N_18154,N_19383);
nor U20937 (N_20937,N_18996,N_18942);
xnor U20938 (N_20938,N_18688,N_18300);
and U20939 (N_20939,N_18271,N_18581);
and U20940 (N_20940,N_18496,N_18216);
and U20941 (N_20941,N_19835,N_18936);
or U20942 (N_20942,N_19122,N_19662);
nor U20943 (N_20943,N_18451,N_18545);
xnor U20944 (N_20944,N_19534,N_19310);
and U20945 (N_20945,N_18779,N_18655);
nor U20946 (N_20946,N_18645,N_19436);
nand U20947 (N_20947,N_19221,N_18880);
xor U20948 (N_20948,N_19623,N_19973);
nand U20949 (N_20949,N_18363,N_19417);
xor U20950 (N_20950,N_19438,N_19665);
and U20951 (N_20951,N_18988,N_18956);
nand U20952 (N_20952,N_19197,N_19767);
and U20953 (N_20953,N_19929,N_18620);
and U20954 (N_20954,N_18480,N_18494);
and U20955 (N_20955,N_18170,N_19270);
and U20956 (N_20956,N_19340,N_19399);
or U20957 (N_20957,N_18970,N_18524);
and U20958 (N_20958,N_19800,N_18712);
xor U20959 (N_20959,N_18605,N_19549);
xnor U20960 (N_20960,N_19705,N_18477);
and U20961 (N_20961,N_18659,N_18204);
and U20962 (N_20962,N_18703,N_19901);
and U20963 (N_20963,N_18948,N_19070);
xor U20964 (N_20964,N_19490,N_19584);
nand U20965 (N_20965,N_19637,N_19273);
xnor U20966 (N_20966,N_19592,N_19741);
and U20967 (N_20967,N_18990,N_19011);
xor U20968 (N_20968,N_19146,N_18051);
nand U20969 (N_20969,N_19072,N_19552);
or U20970 (N_20970,N_18240,N_19618);
nor U20971 (N_20971,N_19811,N_19822);
nor U20972 (N_20972,N_19338,N_19644);
and U20973 (N_20973,N_19170,N_18834);
nand U20974 (N_20974,N_18845,N_18177);
or U20975 (N_20975,N_19856,N_18958);
nor U20976 (N_20976,N_19339,N_18664);
nand U20977 (N_20977,N_19402,N_19029);
or U20978 (N_20978,N_18716,N_19564);
nor U20979 (N_20979,N_19959,N_19251);
xor U20980 (N_20980,N_18043,N_18131);
or U20981 (N_20981,N_18200,N_19337);
nand U20982 (N_20982,N_18033,N_19517);
nand U20983 (N_20983,N_18352,N_19437);
nand U20984 (N_20984,N_19037,N_18665);
xor U20985 (N_20985,N_19086,N_18457);
or U20986 (N_20986,N_19483,N_19203);
nor U20987 (N_20987,N_19590,N_18497);
xnor U20988 (N_20988,N_18658,N_19274);
nor U20989 (N_20989,N_19740,N_19748);
xor U20990 (N_20990,N_18049,N_18207);
xor U20991 (N_20991,N_19757,N_18374);
and U20992 (N_20992,N_19411,N_18766);
nor U20993 (N_20993,N_19591,N_18247);
or U20994 (N_20994,N_18731,N_18248);
and U20995 (N_20995,N_18226,N_18130);
and U20996 (N_20996,N_18923,N_18853);
and U20997 (N_20997,N_18099,N_18742);
nand U20998 (N_20998,N_19232,N_19737);
nor U20999 (N_20999,N_18660,N_18458);
nand U21000 (N_21000,N_19730,N_19217);
and U21001 (N_21001,N_18132,N_18656);
xor U21002 (N_21002,N_19544,N_19509);
nand U21003 (N_21003,N_18176,N_19395);
xor U21004 (N_21004,N_19601,N_18352);
nor U21005 (N_21005,N_18517,N_18931);
and U21006 (N_21006,N_19793,N_18144);
xnor U21007 (N_21007,N_18114,N_19822);
or U21008 (N_21008,N_19619,N_18383);
nor U21009 (N_21009,N_18858,N_19887);
nand U21010 (N_21010,N_18543,N_18052);
xor U21011 (N_21011,N_18774,N_18814);
and U21012 (N_21012,N_18101,N_19839);
nor U21013 (N_21013,N_19260,N_18875);
xnor U21014 (N_21014,N_18553,N_19302);
or U21015 (N_21015,N_19330,N_18486);
xor U21016 (N_21016,N_19588,N_19697);
xor U21017 (N_21017,N_19764,N_18299);
or U21018 (N_21018,N_18426,N_18493);
nor U21019 (N_21019,N_18899,N_19419);
nor U21020 (N_21020,N_19398,N_19023);
nand U21021 (N_21021,N_19193,N_19934);
or U21022 (N_21022,N_19015,N_18875);
or U21023 (N_21023,N_18403,N_18940);
nor U21024 (N_21024,N_19995,N_18469);
xor U21025 (N_21025,N_19281,N_18339);
nand U21026 (N_21026,N_18054,N_18702);
xnor U21027 (N_21027,N_18405,N_19834);
and U21028 (N_21028,N_18834,N_18430);
and U21029 (N_21029,N_18173,N_19196);
and U21030 (N_21030,N_18534,N_18301);
xnor U21031 (N_21031,N_19063,N_18379);
xnor U21032 (N_21032,N_19069,N_18596);
nor U21033 (N_21033,N_18891,N_18900);
nor U21034 (N_21034,N_18374,N_19749);
and U21035 (N_21035,N_18795,N_19446);
and U21036 (N_21036,N_19149,N_19477);
nand U21037 (N_21037,N_18099,N_19733);
nand U21038 (N_21038,N_19741,N_19916);
nor U21039 (N_21039,N_19210,N_19350);
nor U21040 (N_21040,N_18883,N_18114);
nor U21041 (N_21041,N_18387,N_18576);
nand U21042 (N_21042,N_18787,N_19517);
xnor U21043 (N_21043,N_18211,N_19621);
nor U21044 (N_21044,N_19145,N_18404);
and U21045 (N_21045,N_19459,N_19366);
and U21046 (N_21046,N_19604,N_18595);
xnor U21047 (N_21047,N_19357,N_18985);
xnor U21048 (N_21048,N_19091,N_19621);
xnor U21049 (N_21049,N_19514,N_18264);
xor U21050 (N_21050,N_18487,N_18747);
nor U21051 (N_21051,N_18863,N_18823);
nand U21052 (N_21052,N_19050,N_19381);
nor U21053 (N_21053,N_18798,N_18805);
nand U21054 (N_21054,N_18207,N_18822);
nor U21055 (N_21055,N_18378,N_18180);
nand U21056 (N_21056,N_19967,N_19556);
xor U21057 (N_21057,N_18760,N_19856);
xor U21058 (N_21058,N_19135,N_19993);
or U21059 (N_21059,N_18319,N_19143);
or U21060 (N_21060,N_19855,N_19684);
nor U21061 (N_21061,N_18869,N_19444);
nand U21062 (N_21062,N_19190,N_18580);
nand U21063 (N_21063,N_19103,N_19043);
xnor U21064 (N_21064,N_18202,N_18267);
nor U21065 (N_21065,N_18798,N_18797);
and U21066 (N_21066,N_18006,N_18912);
xnor U21067 (N_21067,N_18645,N_18052);
nor U21068 (N_21068,N_18709,N_19349);
nor U21069 (N_21069,N_18582,N_19170);
and U21070 (N_21070,N_18728,N_18816);
nor U21071 (N_21071,N_18387,N_18820);
or U21072 (N_21072,N_19475,N_19054);
and U21073 (N_21073,N_18542,N_18938);
nand U21074 (N_21074,N_19533,N_18061);
nor U21075 (N_21075,N_19262,N_19199);
xnor U21076 (N_21076,N_18645,N_18330);
xor U21077 (N_21077,N_18649,N_19319);
and U21078 (N_21078,N_18772,N_18607);
or U21079 (N_21079,N_19683,N_18268);
xor U21080 (N_21080,N_18354,N_18328);
xor U21081 (N_21081,N_19562,N_18271);
and U21082 (N_21082,N_18940,N_19599);
nor U21083 (N_21083,N_18653,N_18926);
nor U21084 (N_21084,N_19896,N_18069);
and U21085 (N_21085,N_19012,N_18696);
or U21086 (N_21086,N_19758,N_18081);
and U21087 (N_21087,N_19087,N_19152);
and U21088 (N_21088,N_18093,N_19861);
or U21089 (N_21089,N_19418,N_18102);
nor U21090 (N_21090,N_19775,N_18233);
or U21091 (N_21091,N_18843,N_18868);
xnor U21092 (N_21092,N_19542,N_18945);
or U21093 (N_21093,N_18431,N_19462);
xor U21094 (N_21094,N_19381,N_19127);
nand U21095 (N_21095,N_18332,N_18463);
or U21096 (N_21096,N_19997,N_19450);
xnor U21097 (N_21097,N_18865,N_18111);
nand U21098 (N_21098,N_19585,N_18102);
or U21099 (N_21099,N_18550,N_19407);
and U21100 (N_21100,N_19292,N_18729);
and U21101 (N_21101,N_19869,N_18498);
or U21102 (N_21102,N_19285,N_18308);
nor U21103 (N_21103,N_19177,N_18899);
nand U21104 (N_21104,N_18573,N_19010);
nor U21105 (N_21105,N_19711,N_18385);
nand U21106 (N_21106,N_18634,N_19318);
xnor U21107 (N_21107,N_18772,N_19485);
nor U21108 (N_21108,N_19304,N_18248);
nor U21109 (N_21109,N_19793,N_18498);
xnor U21110 (N_21110,N_19345,N_19396);
xnor U21111 (N_21111,N_18072,N_19714);
and U21112 (N_21112,N_18021,N_19792);
and U21113 (N_21113,N_19123,N_19793);
and U21114 (N_21114,N_19006,N_19120);
and U21115 (N_21115,N_19984,N_19066);
nor U21116 (N_21116,N_18360,N_18673);
nand U21117 (N_21117,N_19991,N_18019);
nand U21118 (N_21118,N_19030,N_19430);
nand U21119 (N_21119,N_18600,N_19006);
and U21120 (N_21120,N_19982,N_19092);
and U21121 (N_21121,N_18073,N_19474);
nand U21122 (N_21122,N_18741,N_18135);
and U21123 (N_21123,N_18174,N_18314);
nor U21124 (N_21124,N_19122,N_18326);
xnor U21125 (N_21125,N_19678,N_19580);
or U21126 (N_21126,N_19462,N_18029);
nand U21127 (N_21127,N_18916,N_19217);
nor U21128 (N_21128,N_19077,N_19876);
xnor U21129 (N_21129,N_18864,N_18574);
or U21130 (N_21130,N_18462,N_18950);
xnor U21131 (N_21131,N_18308,N_19731);
or U21132 (N_21132,N_18414,N_18506);
xnor U21133 (N_21133,N_18510,N_18640);
nand U21134 (N_21134,N_18916,N_18141);
or U21135 (N_21135,N_19284,N_19741);
or U21136 (N_21136,N_19297,N_18306);
or U21137 (N_21137,N_18170,N_18138);
and U21138 (N_21138,N_19425,N_18606);
xnor U21139 (N_21139,N_18787,N_18297);
nor U21140 (N_21140,N_18880,N_18236);
or U21141 (N_21141,N_18098,N_18390);
nor U21142 (N_21142,N_19015,N_19521);
nor U21143 (N_21143,N_19164,N_19472);
nor U21144 (N_21144,N_18025,N_18494);
xor U21145 (N_21145,N_18482,N_19846);
and U21146 (N_21146,N_19976,N_18941);
nor U21147 (N_21147,N_19238,N_19635);
and U21148 (N_21148,N_19353,N_19608);
nand U21149 (N_21149,N_19024,N_18913);
or U21150 (N_21150,N_18710,N_19963);
nand U21151 (N_21151,N_18069,N_18539);
nand U21152 (N_21152,N_19623,N_19899);
and U21153 (N_21153,N_19637,N_18702);
and U21154 (N_21154,N_19334,N_18802);
xor U21155 (N_21155,N_18751,N_19466);
nand U21156 (N_21156,N_18550,N_18854);
and U21157 (N_21157,N_19491,N_19498);
or U21158 (N_21158,N_18821,N_18219);
nor U21159 (N_21159,N_18630,N_19375);
or U21160 (N_21160,N_18007,N_19106);
xor U21161 (N_21161,N_19372,N_19184);
xor U21162 (N_21162,N_18653,N_18482);
nand U21163 (N_21163,N_18576,N_18920);
and U21164 (N_21164,N_19678,N_18365);
and U21165 (N_21165,N_18059,N_19510);
nor U21166 (N_21166,N_18489,N_18395);
nand U21167 (N_21167,N_18290,N_18163);
nor U21168 (N_21168,N_18325,N_18695);
xor U21169 (N_21169,N_19121,N_19596);
or U21170 (N_21170,N_19577,N_18680);
nand U21171 (N_21171,N_19980,N_19413);
nor U21172 (N_21172,N_19616,N_18986);
and U21173 (N_21173,N_19706,N_18411);
xor U21174 (N_21174,N_18869,N_18498);
xnor U21175 (N_21175,N_19378,N_19740);
and U21176 (N_21176,N_19051,N_19035);
nor U21177 (N_21177,N_18829,N_18679);
nand U21178 (N_21178,N_18621,N_19157);
nand U21179 (N_21179,N_19221,N_19069);
or U21180 (N_21180,N_19127,N_18534);
nand U21181 (N_21181,N_18294,N_18999);
xor U21182 (N_21182,N_18000,N_19588);
and U21183 (N_21183,N_18275,N_19383);
xor U21184 (N_21184,N_18277,N_18736);
and U21185 (N_21185,N_19491,N_18456);
and U21186 (N_21186,N_19517,N_19314);
or U21187 (N_21187,N_19524,N_18563);
or U21188 (N_21188,N_19928,N_18213);
or U21189 (N_21189,N_18933,N_19299);
nor U21190 (N_21190,N_18485,N_19158);
or U21191 (N_21191,N_19720,N_18068);
xor U21192 (N_21192,N_18133,N_19755);
and U21193 (N_21193,N_18995,N_18986);
nor U21194 (N_21194,N_19285,N_18591);
or U21195 (N_21195,N_18609,N_18886);
and U21196 (N_21196,N_18988,N_19257);
or U21197 (N_21197,N_18176,N_19340);
nor U21198 (N_21198,N_19021,N_18463);
nand U21199 (N_21199,N_19909,N_18820);
nor U21200 (N_21200,N_19265,N_19472);
nor U21201 (N_21201,N_18115,N_19584);
or U21202 (N_21202,N_19974,N_18570);
xnor U21203 (N_21203,N_19172,N_19692);
xor U21204 (N_21204,N_19960,N_18424);
nor U21205 (N_21205,N_19869,N_19581);
xnor U21206 (N_21206,N_19117,N_18718);
and U21207 (N_21207,N_18545,N_18317);
xor U21208 (N_21208,N_18132,N_18708);
and U21209 (N_21209,N_18894,N_19168);
and U21210 (N_21210,N_19304,N_18885);
and U21211 (N_21211,N_18409,N_18321);
and U21212 (N_21212,N_19883,N_18513);
and U21213 (N_21213,N_18918,N_18646);
nand U21214 (N_21214,N_19273,N_19839);
and U21215 (N_21215,N_18831,N_19789);
nand U21216 (N_21216,N_18251,N_19359);
nand U21217 (N_21217,N_18302,N_19298);
nand U21218 (N_21218,N_19412,N_19132);
nor U21219 (N_21219,N_19817,N_19423);
and U21220 (N_21220,N_18638,N_18430);
nand U21221 (N_21221,N_18383,N_19377);
nand U21222 (N_21222,N_18346,N_18720);
and U21223 (N_21223,N_18719,N_18367);
nor U21224 (N_21224,N_18347,N_18897);
xnor U21225 (N_21225,N_18359,N_18929);
xnor U21226 (N_21226,N_19893,N_18923);
or U21227 (N_21227,N_18851,N_19400);
xor U21228 (N_21228,N_18404,N_18619);
and U21229 (N_21229,N_18088,N_18163);
or U21230 (N_21230,N_18606,N_19157);
and U21231 (N_21231,N_18676,N_18810);
or U21232 (N_21232,N_19812,N_18939);
xnor U21233 (N_21233,N_18898,N_19395);
nor U21234 (N_21234,N_18458,N_18197);
nand U21235 (N_21235,N_18747,N_18457);
or U21236 (N_21236,N_19211,N_19839);
xor U21237 (N_21237,N_19148,N_18097);
and U21238 (N_21238,N_18864,N_18241);
or U21239 (N_21239,N_19156,N_18657);
and U21240 (N_21240,N_18072,N_19277);
nor U21241 (N_21241,N_19656,N_19686);
or U21242 (N_21242,N_19626,N_19439);
and U21243 (N_21243,N_18099,N_18485);
nor U21244 (N_21244,N_18007,N_18103);
xor U21245 (N_21245,N_19988,N_18456);
and U21246 (N_21246,N_19817,N_18955);
or U21247 (N_21247,N_18154,N_19337);
or U21248 (N_21248,N_18252,N_19388);
nand U21249 (N_21249,N_19247,N_19731);
nand U21250 (N_21250,N_19840,N_19924);
and U21251 (N_21251,N_18629,N_19644);
and U21252 (N_21252,N_18544,N_19148);
nand U21253 (N_21253,N_19471,N_18936);
xor U21254 (N_21254,N_18050,N_19627);
or U21255 (N_21255,N_18816,N_19702);
and U21256 (N_21256,N_18222,N_18286);
and U21257 (N_21257,N_19203,N_18126);
nor U21258 (N_21258,N_18187,N_18540);
nand U21259 (N_21259,N_18316,N_18026);
or U21260 (N_21260,N_18714,N_19678);
and U21261 (N_21261,N_18596,N_19671);
xor U21262 (N_21262,N_19842,N_18745);
or U21263 (N_21263,N_18491,N_19069);
nor U21264 (N_21264,N_18319,N_19500);
and U21265 (N_21265,N_18179,N_19908);
or U21266 (N_21266,N_18215,N_18307);
xnor U21267 (N_21267,N_18477,N_19637);
nor U21268 (N_21268,N_18812,N_19319);
and U21269 (N_21269,N_18768,N_18399);
and U21270 (N_21270,N_18998,N_19832);
xnor U21271 (N_21271,N_19862,N_19611);
xnor U21272 (N_21272,N_18983,N_19548);
nand U21273 (N_21273,N_19768,N_18287);
xnor U21274 (N_21274,N_18224,N_18741);
xnor U21275 (N_21275,N_19150,N_19009);
xor U21276 (N_21276,N_18435,N_18966);
nand U21277 (N_21277,N_18109,N_18089);
nor U21278 (N_21278,N_18434,N_18916);
or U21279 (N_21279,N_18623,N_19477);
and U21280 (N_21280,N_19239,N_19759);
nand U21281 (N_21281,N_18211,N_19992);
or U21282 (N_21282,N_18183,N_18280);
xor U21283 (N_21283,N_19515,N_19586);
nand U21284 (N_21284,N_19919,N_18779);
and U21285 (N_21285,N_19709,N_19042);
xnor U21286 (N_21286,N_19681,N_19032);
nor U21287 (N_21287,N_18636,N_19942);
nand U21288 (N_21288,N_19693,N_18307);
or U21289 (N_21289,N_19407,N_19483);
and U21290 (N_21290,N_18796,N_19520);
nand U21291 (N_21291,N_18402,N_18893);
or U21292 (N_21292,N_19969,N_19053);
and U21293 (N_21293,N_18928,N_19074);
nor U21294 (N_21294,N_19396,N_18050);
xnor U21295 (N_21295,N_18160,N_19255);
xor U21296 (N_21296,N_18652,N_18187);
nor U21297 (N_21297,N_19407,N_18307);
and U21298 (N_21298,N_18849,N_18794);
xnor U21299 (N_21299,N_18059,N_19036);
and U21300 (N_21300,N_18836,N_18913);
and U21301 (N_21301,N_18219,N_18276);
nand U21302 (N_21302,N_18389,N_18894);
nor U21303 (N_21303,N_18061,N_18087);
nor U21304 (N_21304,N_19843,N_19189);
xor U21305 (N_21305,N_19909,N_18196);
or U21306 (N_21306,N_18793,N_18695);
or U21307 (N_21307,N_19952,N_18475);
xor U21308 (N_21308,N_18586,N_19308);
and U21309 (N_21309,N_19968,N_18850);
xnor U21310 (N_21310,N_19076,N_18980);
or U21311 (N_21311,N_19164,N_19526);
nand U21312 (N_21312,N_18338,N_18363);
and U21313 (N_21313,N_19849,N_19706);
xnor U21314 (N_21314,N_18246,N_19591);
xnor U21315 (N_21315,N_18954,N_18432);
xnor U21316 (N_21316,N_18115,N_18240);
or U21317 (N_21317,N_19639,N_19740);
xnor U21318 (N_21318,N_18409,N_18145);
nor U21319 (N_21319,N_19302,N_18914);
and U21320 (N_21320,N_18715,N_18905);
and U21321 (N_21321,N_19311,N_19822);
or U21322 (N_21322,N_19866,N_18018);
nor U21323 (N_21323,N_18541,N_19855);
and U21324 (N_21324,N_19383,N_19666);
nor U21325 (N_21325,N_18150,N_18943);
nand U21326 (N_21326,N_18110,N_18201);
and U21327 (N_21327,N_18247,N_18697);
nor U21328 (N_21328,N_18860,N_18578);
and U21329 (N_21329,N_18499,N_19112);
xnor U21330 (N_21330,N_18669,N_19378);
and U21331 (N_21331,N_19592,N_18873);
or U21332 (N_21332,N_18905,N_19102);
or U21333 (N_21333,N_19611,N_19913);
or U21334 (N_21334,N_18745,N_18659);
nor U21335 (N_21335,N_19647,N_18423);
and U21336 (N_21336,N_18123,N_19273);
nand U21337 (N_21337,N_19992,N_18367);
nor U21338 (N_21338,N_19546,N_19549);
nor U21339 (N_21339,N_19961,N_18442);
nor U21340 (N_21340,N_18320,N_19988);
xor U21341 (N_21341,N_19465,N_18516);
nor U21342 (N_21342,N_18253,N_18857);
or U21343 (N_21343,N_19930,N_18350);
or U21344 (N_21344,N_19059,N_18634);
nand U21345 (N_21345,N_18099,N_19002);
xor U21346 (N_21346,N_18597,N_18408);
nand U21347 (N_21347,N_18527,N_18335);
and U21348 (N_21348,N_19851,N_19040);
or U21349 (N_21349,N_18973,N_18060);
or U21350 (N_21350,N_18560,N_19155);
xor U21351 (N_21351,N_19515,N_18235);
or U21352 (N_21352,N_18798,N_18956);
nor U21353 (N_21353,N_19538,N_19432);
xor U21354 (N_21354,N_18912,N_18569);
nand U21355 (N_21355,N_18374,N_19021);
and U21356 (N_21356,N_18755,N_19000);
nor U21357 (N_21357,N_18563,N_19136);
or U21358 (N_21358,N_18367,N_19153);
or U21359 (N_21359,N_19156,N_18391);
xor U21360 (N_21360,N_18949,N_18070);
or U21361 (N_21361,N_18967,N_18128);
xnor U21362 (N_21362,N_19836,N_18232);
nor U21363 (N_21363,N_18908,N_19266);
nor U21364 (N_21364,N_19909,N_18448);
and U21365 (N_21365,N_18250,N_19581);
or U21366 (N_21366,N_19317,N_18561);
nor U21367 (N_21367,N_19430,N_18710);
or U21368 (N_21368,N_18913,N_19169);
nand U21369 (N_21369,N_18701,N_18929);
and U21370 (N_21370,N_18800,N_19167);
or U21371 (N_21371,N_19230,N_18163);
or U21372 (N_21372,N_18601,N_18657);
and U21373 (N_21373,N_19450,N_19405);
nor U21374 (N_21374,N_19137,N_19247);
and U21375 (N_21375,N_19625,N_19692);
xnor U21376 (N_21376,N_19794,N_19428);
nor U21377 (N_21377,N_19478,N_19324);
xor U21378 (N_21378,N_18284,N_19213);
or U21379 (N_21379,N_19171,N_18574);
nor U21380 (N_21380,N_19718,N_18471);
nand U21381 (N_21381,N_18515,N_19413);
xor U21382 (N_21382,N_18437,N_18599);
nor U21383 (N_21383,N_19365,N_19318);
nor U21384 (N_21384,N_19354,N_19396);
xnor U21385 (N_21385,N_19455,N_18847);
nor U21386 (N_21386,N_19521,N_18696);
xnor U21387 (N_21387,N_19475,N_18112);
or U21388 (N_21388,N_19921,N_18408);
xor U21389 (N_21389,N_18717,N_18864);
and U21390 (N_21390,N_18050,N_19504);
and U21391 (N_21391,N_19022,N_19068);
nand U21392 (N_21392,N_19766,N_18719);
nand U21393 (N_21393,N_19840,N_19799);
or U21394 (N_21394,N_19608,N_18784);
or U21395 (N_21395,N_19387,N_18506);
and U21396 (N_21396,N_19495,N_19315);
or U21397 (N_21397,N_18085,N_19293);
nand U21398 (N_21398,N_18089,N_19030);
nand U21399 (N_21399,N_19257,N_18799);
nand U21400 (N_21400,N_19664,N_18904);
nor U21401 (N_21401,N_18851,N_19018);
nor U21402 (N_21402,N_19214,N_19702);
nor U21403 (N_21403,N_19505,N_18514);
and U21404 (N_21404,N_19078,N_19750);
or U21405 (N_21405,N_18742,N_18985);
or U21406 (N_21406,N_18373,N_19749);
or U21407 (N_21407,N_18828,N_18576);
or U21408 (N_21408,N_19589,N_18348);
nand U21409 (N_21409,N_19514,N_19684);
nor U21410 (N_21410,N_19524,N_19782);
and U21411 (N_21411,N_19119,N_19620);
nor U21412 (N_21412,N_18755,N_19966);
and U21413 (N_21413,N_19423,N_18706);
nor U21414 (N_21414,N_19399,N_18106);
or U21415 (N_21415,N_19583,N_19412);
xnor U21416 (N_21416,N_19679,N_19154);
or U21417 (N_21417,N_19007,N_19862);
and U21418 (N_21418,N_18421,N_18636);
xor U21419 (N_21419,N_18860,N_19693);
nand U21420 (N_21420,N_18675,N_19450);
and U21421 (N_21421,N_19134,N_18229);
xor U21422 (N_21422,N_19362,N_18516);
nand U21423 (N_21423,N_19396,N_18332);
or U21424 (N_21424,N_19680,N_18676);
or U21425 (N_21425,N_19093,N_19102);
or U21426 (N_21426,N_18144,N_18924);
nand U21427 (N_21427,N_18934,N_18691);
nor U21428 (N_21428,N_19878,N_19700);
xnor U21429 (N_21429,N_19137,N_19179);
nand U21430 (N_21430,N_19372,N_19082);
or U21431 (N_21431,N_18445,N_19806);
xnor U21432 (N_21432,N_18811,N_19548);
or U21433 (N_21433,N_19282,N_19027);
nand U21434 (N_21434,N_19750,N_19377);
or U21435 (N_21435,N_19147,N_18273);
nand U21436 (N_21436,N_19117,N_19782);
or U21437 (N_21437,N_18054,N_18373);
nand U21438 (N_21438,N_18175,N_18255);
nor U21439 (N_21439,N_19543,N_19429);
and U21440 (N_21440,N_19484,N_19620);
or U21441 (N_21441,N_18379,N_18997);
or U21442 (N_21442,N_18671,N_19003);
and U21443 (N_21443,N_18913,N_19436);
or U21444 (N_21444,N_18008,N_19666);
nor U21445 (N_21445,N_18148,N_18441);
or U21446 (N_21446,N_18618,N_19437);
nor U21447 (N_21447,N_19536,N_18711);
nor U21448 (N_21448,N_18302,N_18729);
or U21449 (N_21449,N_19231,N_18799);
or U21450 (N_21450,N_19895,N_19090);
nor U21451 (N_21451,N_19573,N_19050);
nand U21452 (N_21452,N_18890,N_18053);
and U21453 (N_21453,N_18719,N_18838);
and U21454 (N_21454,N_18013,N_18774);
and U21455 (N_21455,N_18228,N_19523);
nand U21456 (N_21456,N_18367,N_18609);
nand U21457 (N_21457,N_19238,N_18421);
xor U21458 (N_21458,N_19970,N_19251);
and U21459 (N_21459,N_19293,N_18740);
and U21460 (N_21460,N_19909,N_19972);
xnor U21461 (N_21461,N_19533,N_18982);
xnor U21462 (N_21462,N_18339,N_19759);
or U21463 (N_21463,N_18653,N_19262);
nand U21464 (N_21464,N_18571,N_18009);
nor U21465 (N_21465,N_18291,N_18138);
nand U21466 (N_21466,N_18613,N_18564);
nand U21467 (N_21467,N_18322,N_19468);
nor U21468 (N_21468,N_19487,N_18045);
nor U21469 (N_21469,N_18962,N_19446);
or U21470 (N_21470,N_19438,N_19660);
or U21471 (N_21471,N_19273,N_19471);
xnor U21472 (N_21472,N_19241,N_19953);
nor U21473 (N_21473,N_19937,N_18099);
and U21474 (N_21474,N_18902,N_18284);
or U21475 (N_21475,N_19982,N_19271);
nor U21476 (N_21476,N_19144,N_19535);
or U21477 (N_21477,N_18636,N_18757);
xor U21478 (N_21478,N_19845,N_19857);
nor U21479 (N_21479,N_18555,N_19101);
nand U21480 (N_21480,N_19835,N_19402);
xor U21481 (N_21481,N_18811,N_19824);
xor U21482 (N_21482,N_18569,N_19150);
xor U21483 (N_21483,N_18325,N_18409);
or U21484 (N_21484,N_19813,N_19892);
nor U21485 (N_21485,N_19071,N_18797);
or U21486 (N_21486,N_18384,N_18827);
xnor U21487 (N_21487,N_19464,N_18227);
and U21488 (N_21488,N_19198,N_19688);
nor U21489 (N_21489,N_18453,N_19520);
or U21490 (N_21490,N_18203,N_18961);
xnor U21491 (N_21491,N_19037,N_19924);
or U21492 (N_21492,N_18493,N_19101);
xor U21493 (N_21493,N_19467,N_19390);
and U21494 (N_21494,N_19421,N_18509);
nand U21495 (N_21495,N_18722,N_19576);
or U21496 (N_21496,N_18713,N_19371);
nor U21497 (N_21497,N_18033,N_18249);
nand U21498 (N_21498,N_19989,N_18495);
or U21499 (N_21499,N_19834,N_18232);
nand U21500 (N_21500,N_18313,N_19260);
nor U21501 (N_21501,N_18074,N_18417);
xnor U21502 (N_21502,N_18009,N_19004);
nand U21503 (N_21503,N_19127,N_19238);
nand U21504 (N_21504,N_19923,N_19095);
xor U21505 (N_21505,N_18183,N_19913);
or U21506 (N_21506,N_19442,N_19331);
nor U21507 (N_21507,N_18823,N_19357);
nor U21508 (N_21508,N_18458,N_18893);
or U21509 (N_21509,N_19948,N_18384);
nor U21510 (N_21510,N_18034,N_19631);
nor U21511 (N_21511,N_18657,N_18043);
and U21512 (N_21512,N_19812,N_19540);
and U21513 (N_21513,N_18344,N_19921);
and U21514 (N_21514,N_18522,N_19207);
and U21515 (N_21515,N_18228,N_18151);
and U21516 (N_21516,N_18797,N_19427);
xor U21517 (N_21517,N_18578,N_18341);
or U21518 (N_21518,N_19936,N_18248);
nor U21519 (N_21519,N_19749,N_19467);
or U21520 (N_21520,N_18115,N_18004);
and U21521 (N_21521,N_18271,N_19048);
nand U21522 (N_21522,N_19307,N_18940);
and U21523 (N_21523,N_19519,N_18301);
nor U21524 (N_21524,N_18542,N_19459);
and U21525 (N_21525,N_18832,N_18112);
nand U21526 (N_21526,N_18522,N_19545);
and U21527 (N_21527,N_19484,N_18266);
nor U21528 (N_21528,N_18341,N_18403);
xor U21529 (N_21529,N_19037,N_18605);
nand U21530 (N_21530,N_18815,N_19246);
nor U21531 (N_21531,N_18796,N_18976);
or U21532 (N_21532,N_18848,N_18413);
and U21533 (N_21533,N_18451,N_19666);
and U21534 (N_21534,N_18473,N_18894);
and U21535 (N_21535,N_18704,N_19388);
and U21536 (N_21536,N_18156,N_19832);
nor U21537 (N_21537,N_18558,N_19231);
xor U21538 (N_21538,N_19796,N_19590);
nand U21539 (N_21539,N_18556,N_18712);
xnor U21540 (N_21540,N_19751,N_19894);
nand U21541 (N_21541,N_19509,N_18543);
xor U21542 (N_21542,N_18947,N_18419);
xor U21543 (N_21543,N_18838,N_18152);
and U21544 (N_21544,N_18008,N_19098);
nor U21545 (N_21545,N_19051,N_19832);
and U21546 (N_21546,N_18303,N_18592);
or U21547 (N_21547,N_18816,N_18906);
and U21548 (N_21548,N_19131,N_18111);
or U21549 (N_21549,N_19146,N_18018);
or U21550 (N_21550,N_19063,N_18403);
nor U21551 (N_21551,N_18735,N_19980);
xnor U21552 (N_21552,N_18559,N_19716);
or U21553 (N_21553,N_18186,N_18617);
xor U21554 (N_21554,N_19200,N_18906);
nand U21555 (N_21555,N_18994,N_19190);
xnor U21556 (N_21556,N_19747,N_18460);
and U21557 (N_21557,N_19131,N_18029);
nand U21558 (N_21558,N_19221,N_18878);
nand U21559 (N_21559,N_18190,N_19359);
nand U21560 (N_21560,N_19530,N_18397);
xor U21561 (N_21561,N_19404,N_19176);
nand U21562 (N_21562,N_18640,N_18934);
xnor U21563 (N_21563,N_18736,N_18356);
and U21564 (N_21564,N_18733,N_18730);
nand U21565 (N_21565,N_19305,N_18195);
xnor U21566 (N_21566,N_19241,N_18672);
xnor U21567 (N_21567,N_19696,N_18294);
xor U21568 (N_21568,N_18846,N_18827);
and U21569 (N_21569,N_18376,N_19727);
xnor U21570 (N_21570,N_18576,N_19207);
nand U21571 (N_21571,N_18182,N_19370);
nor U21572 (N_21572,N_19737,N_19066);
or U21573 (N_21573,N_19506,N_19246);
nand U21574 (N_21574,N_19628,N_18152);
and U21575 (N_21575,N_19606,N_19098);
or U21576 (N_21576,N_19468,N_19542);
xor U21577 (N_21577,N_18129,N_19716);
or U21578 (N_21578,N_19276,N_19675);
nor U21579 (N_21579,N_19761,N_18666);
or U21580 (N_21580,N_18421,N_19397);
or U21581 (N_21581,N_18268,N_18161);
xor U21582 (N_21582,N_18687,N_19774);
nand U21583 (N_21583,N_18268,N_18688);
nand U21584 (N_21584,N_19921,N_19162);
or U21585 (N_21585,N_19803,N_18504);
nand U21586 (N_21586,N_18175,N_18408);
xor U21587 (N_21587,N_18821,N_19448);
nand U21588 (N_21588,N_19373,N_19194);
nor U21589 (N_21589,N_19005,N_18637);
xnor U21590 (N_21590,N_19958,N_18157);
nor U21591 (N_21591,N_18136,N_18838);
and U21592 (N_21592,N_19760,N_19429);
nand U21593 (N_21593,N_19539,N_19304);
nand U21594 (N_21594,N_19702,N_19146);
nor U21595 (N_21595,N_19722,N_18881);
xnor U21596 (N_21596,N_19834,N_19303);
nor U21597 (N_21597,N_19657,N_18892);
nor U21598 (N_21598,N_18453,N_18077);
nand U21599 (N_21599,N_18870,N_18321);
xnor U21600 (N_21600,N_18370,N_18350);
or U21601 (N_21601,N_18853,N_18778);
and U21602 (N_21602,N_19895,N_18619);
or U21603 (N_21603,N_19204,N_19849);
nor U21604 (N_21604,N_19345,N_19923);
nand U21605 (N_21605,N_18168,N_18330);
and U21606 (N_21606,N_19915,N_19044);
or U21607 (N_21607,N_18390,N_19565);
nand U21608 (N_21608,N_19762,N_19401);
xnor U21609 (N_21609,N_19126,N_19049);
nand U21610 (N_21610,N_19078,N_18457);
xnor U21611 (N_21611,N_18523,N_18084);
and U21612 (N_21612,N_18025,N_18882);
nor U21613 (N_21613,N_19166,N_18409);
xor U21614 (N_21614,N_18465,N_18822);
and U21615 (N_21615,N_18499,N_19106);
and U21616 (N_21616,N_18660,N_19885);
nand U21617 (N_21617,N_18949,N_19600);
xor U21618 (N_21618,N_19250,N_19428);
nand U21619 (N_21619,N_19926,N_18990);
and U21620 (N_21620,N_18418,N_19484);
or U21621 (N_21621,N_19369,N_18388);
xnor U21622 (N_21622,N_18779,N_18153);
nand U21623 (N_21623,N_18459,N_18137);
xnor U21624 (N_21624,N_18190,N_18725);
or U21625 (N_21625,N_18929,N_19882);
and U21626 (N_21626,N_19004,N_19028);
nand U21627 (N_21627,N_18639,N_18042);
nand U21628 (N_21628,N_19263,N_19300);
or U21629 (N_21629,N_18894,N_18935);
nand U21630 (N_21630,N_18468,N_18899);
nor U21631 (N_21631,N_19610,N_19128);
xnor U21632 (N_21632,N_18016,N_19295);
or U21633 (N_21633,N_19371,N_18259);
and U21634 (N_21634,N_19537,N_19357);
nand U21635 (N_21635,N_18044,N_18572);
xnor U21636 (N_21636,N_19526,N_18418);
and U21637 (N_21637,N_19148,N_18181);
and U21638 (N_21638,N_18905,N_18171);
nand U21639 (N_21639,N_18174,N_18005);
nor U21640 (N_21640,N_18915,N_18880);
and U21641 (N_21641,N_19704,N_19332);
and U21642 (N_21642,N_19719,N_19765);
and U21643 (N_21643,N_18987,N_19100);
or U21644 (N_21644,N_19249,N_19229);
and U21645 (N_21645,N_18056,N_19781);
xor U21646 (N_21646,N_18784,N_18098);
and U21647 (N_21647,N_19540,N_18185);
nand U21648 (N_21648,N_19661,N_18115);
nand U21649 (N_21649,N_19124,N_19386);
xnor U21650 (N_21650,N_18027,N_18024);
xnor U21651 (N_21651,N_18019,N_19169);
nor U21652 (N_21652,N_19393,N_19975);
or U21653 (N_21653,N_18377,N_19547);
and U21654 (N_21654,N_18945,N_19237);
and U21655 (N_21655,N_18595,N_18273);
or U21656 (N_21656,N_18512,N_18936);
xor U21657 (N_21657,N_19279,N_18040);
and U21658 (N_21658,N_18428,N_19678);
and U21659 (N_21659,N_18571,N_18196);
nand U21660 (N_21660,N_19076,N_18671);
nand U21661 (N_21661,N_19560,N_18206);
xor U21662 (N_21662,N_19286,N_19075);
and U21663 (N_21663,N_19549,N_18024);
xor U21664 (N_21664,N_18001,N_18883);
nand U21665 (N_21665,N_19033,N_18434);
xor U21666 (N_21666,N_18893,N_19805);
xor U21667 (N_21667,N_18076,N_19559);
nand U21668 (N_21668,N_18965,N_18269);
nand U21669 (N_21669,N_19418,N_19109);
xor U21670 (N_21670,N_19412,N_19397);
and U21671 (N_21671,N_18376,N_19824);
or U21672 (N_21672,N_18628,N_19997);
nor U21673 (N_21673,N_18841,N_18701);
nand U21674 (N_21674,N_18435,N_18513);
xor U21675 (N_21675,N_18401,N_18134);
nor U21676 (N_21676,N_19562,N_19333);
xor U21677 (N_21677,N_18989,N_19185);
and U21678 (N_21678,N_19432,N_18811);
xnor U21679 (N_21679,N_18872,N_18449);
nand U21680 (N_21680,N_19152,N_19031);
and U21681 (N_21681,N_18108,N_19836);
nand U21682 (N_21682,N_19478,N_19756);
xnor U21683 (N_21683,N_18473,N_19434);
nand U21684 (N_21684,N_19411,N_18980);
nor U21685 (N_21685,N_18578,N_18921);
or U21686 (N_21686,N_18751,N_19807);
nand U21687 (N_21687,N_19654,N_18279);
or U21688 (N_21688,N_18295,N_19352);
nand U21689 (N_21689,N_19065,N_18432);
and U21690 (N_21690,N_18073,N_18956);
or U21691 (N_21691,N_18129,N_18046);
or U21692 (N_21692,N_18691,N_19627);
nor U21693 (N_21693,N_19089,N_18230);
nor U21694 (N_21694,N_18851,N_18202);
xor U21695 (N_21695,N_19269,N_19995);
and U21696 (N_21696,N_19033,N_18686);
nand U21697 (N_21697,N_18843,N_18104);
and U21698 (N_21698,N_18840,N_19265);
nand U21699 (N_21699,N_19562,N_19173);
nand U21700 (N_21700,N_18273,N_19068);
and U21701 (N_21701,N_19140,N_19714);
xor U21702 (N_21702,N_18120,N_19236);
xor U21703 (N_21703,N_18575,N_19662);
and U21704 (N_21704,N_19503,N_18640);
nand U21705 (N_21705,N_19456,N_19624);
and U21706 (N_21706,N_19122,N_19255);
nand U21707 (N_21707,N_19112,N_19748);
nor U21708 (N_21708,N_19918,N_19677);
nand U21709 (N_21709,N_19030,N_19155);
xor U21710 (N_21710,N_19001,N_19542);
nand U21711 (N_21711,N_18191,N_18613);
nor U21712 (N_21712,N_19203,N_18536);
or U21713 (N_21713,N_19544,N_18507);
or U21714 (N_21714,N_19358,N_19018);
xnor U21715 (N_21715,N_18019,N_18751);
xnor U21716 (N_21716,N_18152,N_19629);
and U21717 (N_21717,N_18261,N_19398);
nand U21718 (N_21718,N_19901,N_19966);
xnor U21719 (N_21719,N_18371,N_18635);
xor U21720 (N_21720,N_19660,N_18820);
or U21721 (N_21721,N_19694,N_18184);
and U21722 (N_21722,N_19500,N_18783);
or U21723 (N_21723,N_19012,N_19930);
and U21724 (N_21724,N_18006,N_19877);
xor U21725 (N_21725,N_19936,N_18013);
and U21726 (N_21726,N_18863,N_19767);
xnor U21727 (N_21727,N_18949,N_18765);
nor U21728 (N_21728,N_18518,N_19678);
nor U21729 (N_21729,N_18075,N_19598);
nor U21730 (N_21730,N_18186,N_19905);
xnor U21731 (N_21731,N_18401,N_18903);
nand U21732 (N_21732,N_19913,N_18294);
xnor U21733 (N_21733,N_18894,N_19444);
xor U21734 (N_21734,N_18912,N_18653);
nor U21735 (N_21735,N_19875,N_19712);
nor U21736 (N_21736,N_18429,N_19487);
or U21737 (N_21737,N_18190,N_18458);
xor U21738 (N_21738,N_18541,N_18353);
and U21739 (N_21739,N_19342,N_19457);
and U21740 (N_21740,N_18865,N_18194);
xor U21741 (N_21741,N_18404,N_19725);
or U21742 (N_21742,N_19277,N_18076);
or U21743 (N_21743,N_19363,N_18265);
or U21744 (N_21744,N_19207,N_18783);
nor U21745 (N_21745,N_18758,N_18206);
xnor U21746 (N_21746,N_18886,N_19620);
and U21747 (N_21747,N_19257,N_19935);
nor U21748 (N_21748,N_18299,N_19848);
xor U21749 (N_21749,N_19114,N_19888);
nor U21750 (N_21750,N_19410,N_18944);
nand U21751 (N_21751,N_19296,N_19989);
nand U21752 (N_21752,N_19648,N_18142);
and U21753 (N_21753,N_18124,N_19961);
xor U21754 (N_21754,N_18286,N_19408);
and U21755 (N_21755,N_18255,N_18742);
nor U21756 (N_21756,N_18429,N_18224);
xnor U21757 (N_21757,N_19907,N_18339);
xor U21758 (N_21758,N_19077,N_19794);
nand U21759 (N_21759,N_19248,N_19857);
nand U21760 (N_21760,N_18347,N_19503);
nor U21761 (N_21761,N_19068,N_18140);
or U21762 (N_21762,N_19614,N_19616);
or U21763 (N_21763,N_19488,N_19046);
nand U21764 (N_21764,N_18047,N_18093);
or U21765 (N_21765,N_19272,N_18384);
or U21766 (N_21766,N_18108,N_18682);
xor U21767 (N_21767,N_18068,N_19521);
and U21768 (N_21768,N_19862,N_19375);
xnor U21769 (N_21769,N_18330,N_19921);
and U21770 (N_21770,N_19827,N_19747);
xor U21771 (N_21771,N_19993,N_19600);
or U21772 (N_21772,N_19943,N_18246);
nand U21773 (N_21773,N_18216,N_18922);
nand U21774 (N_21774,N_19919,N_19383);
nand U21775 (N_21775,N_18059,N_19832);
nand U21776 (N_21776,N_19551,N_19814);
or U21777 (N_21777,N_18351,N_18397);
or U21778 (N_21778,N_18372,N_18806);
xor U21779 (N_21779,N_18361,N_19577);
nor U21780 (N_21780,N_19629,N_19004);
nor U21781 (N_21781,N_18180,N_18945);
and U21782 (N_21782,N_18358,N_19040);
or U21783 (N_21783,N_19982,N_18094);
nor U21784 (N_21784,N_19074,N_18831);
nand U21785 (N_21785,N_19906,N_18546);
nor U21786 (N_21786,N_18523,N_19127);
or U21787 (N_21787,N_18152,N_19882);
or U21788 (N_21788,N_18535,N_19611);
nor U21789 (N_21789,N_19650,N_18616);
xnor U21790 (N_21790,N_18875,N_18730);
nand U21791 (N_21791,N_19745,N_19341);
nor U21792 (N_21792,N_18552,N_18379);
xor U21793 (N_21793,N_19400,N_18855);
xnor U21794 (N_21794,N_18068,N_18338);
xnor U21795 (N_21795,N_19621,N_18772);
or U21796 (N_21796,N_19188,N_18568);
or U21797 (N_21797,N_19610,N_19165);
or U21798 (N_21798,N_18197,N_18274);
xnor U21799 (N_21799,N_18702,N_19523);
or U21800 (N_21800,N_19308,N_18910);
xnor U21801 (N_21801,N_19549,N_18641);
xnor U21802 (N_21802,N_18453,N_18358);
xor U21803 (N_21803,N_19190,N_19354);
or U21804 (N_21804,N_18822,N_19725);
nand U21805 (N_21805,N_18213,N_18586);
and U21806 (N_21806,N_19963,N_19254);
nand U21807 (N_21807,N_19849,N_18495);
and U21808 (N_21808,N_19549,N_18986);
xnor U21809 (N_21809,N_18287,N_18228);
nor U21810 (N_21810,N_19247,N_19889);
and U21811 (N_21811,N_18734,N_19512);
xor U21812 (N_21812,N_19473,N_19078);
nor U21813 (N_21813,N_19537,N_19714);
or U21814 (N_21814,N_19232,N_19274);
and U21815 (N_21815,N_18299,N_18982);
and U21816 (N_21816,N_19329,N_18840);
xor U21817 (N_21817,N_19309,N_18140);
nor U21818 (N_21818,N_18444,N_19802);
xor U21819 (N_21819,N_19019,N_19467);
or U21820 (N_21820,N_18991,N_18681);
nand U21821 (N_21821,N_18593,N_19928);
nand U21822 (N_21822,N_19261,N_18525);
xnor U21823 (N_21823,N_19473,N_19407);
nor U21824 (N_21824,N_18093,N_18451);
and U21825 (N_21825,N_19795,N_19740);
and U21826 (N_21826,N_19371,N_19382);
and U21827 (N_21827,N_19910,N_18586);
nor U21828 (N_21828,N_18442,N_19109);
nor U21829 (N_21829,N_19149,N_19753);
xor U21830 (N_21830,N_19443,N_19430);
xor U21831 (N_21831,N_18739,N_19635);
or U21832 (N_21832,N_19257,N_19869);
nor U21833 (N_21833,N_19388,N_19307);
nand U21834 (N_21834,N_19748,N_19675);
or U21835 (N_21835,N_19732,N_18730);
nand U21836 (N_21836,N_19076,N_19083);
xnor U21837 (N_21837,N_18317,N_19325);
nor U21838 (N_21838,N_18267,N_18170);
xor U21839 (N_21839,N_19851,N_18737);
nor U21840 (N_21840,N_19357,N_19994);
nand U21841 (N_21841,N_19746,N_19467);
and U21842 (N_21842,N_19309,N_18314);
nand U21843 (N_21843,N_19922,N_18032);
nor U21844 (N_21844,N_19593,N_19449);
and U21845 (N_21845,N_19712,N_18741);
nor U21846 (N_21846,N_18954,N_19209);
or U21847 (N_21847,N_19502,N_19380);
nor U21848 (N_21848,N_19129,N_19313);
xor U21849 (N_21849,N_18638,N_19200);
or U21850 (N_21850,N_19687,N_19109);
and U21851 (N_21851,N_18097,N_18190);
or U21852 (N_21852,N_19344,N_19484);
or U21853 (N_21853,N_19602,N_19661);
nand U21854 (N_21854,N_18581,N_18511);
or U21855 (N_21855,N_19977,N_18372);
nor U21856 (N_21856,N_18892,N_18353);
and U21857 (N_21857,N_18402,N_19667);
nand U21858 (N_21858,N_19844,N_19701);
xor U21859 (N_21859,N_18763,N_18646);
and U21860 (N_21860,N_19764,N_18612);
xor U21861 (N_21861,N_18505,N_19933);
xnor U21862 (N_21862,N_18865,N_19038);
or U21863 (N_21863,N_19610,N_19845);
nor U21864 (N_21864,N_18541,N_18800);
xor U21865 (N_21865,N_18844,N_18032);
nor U21866 (N_21866,N_18186,N_19255);
and U21867 (N_21867,N_19062,N_19299);
nor U21868 (N_21868,N_19298,N_19349);
xnor U21869 (N_21869,N_19768,N_18964);
nand U21870 (N_21870,N_18782,N_19191);
nor U21871 (N_21871,N_19145,N_19880);
nand U21872 (N_21872,N_19924,N_19317);
and U21873 (N_21873,N_18354,N_19469);
and U21874 (N_21874,N_18066,N_18736);
xnor U21875 (N_21875,N_19021,N_18348);
xor U21876 (N_21876,N_18267,N_19742);
nand U21877 (N_21877,N_19269,N_19340);
nor U21878 (N_21878,N_18626,N_19811);
nor U21879 (N_21879,N_19188,N_18684);
nor U21880 (N_21880,N_18386,N_18787);
or U21881 (N_21881,N_18858,N_19004);
or U21882 (N_21882,N_19361,N_18949);
nand U21883 (N_21883,N_19976,N_19044);
and U21884 (N_21884,N_19598,N_19286);
xnor U21885 (N_21885,N_18057,N_18685);
and U21886 (N_21886,N_19862,N_18522);
nand U21887 (N_21887,N_19768,N_18877);
nor U21888 (N_21888,N_19263,N_19220);
and U21889 (N_21889,N_19708,N_18366);
and U21890 (N_21890,N_18301,N_19053);
xnor U21891 (N_21891,N_18623,N_18864);
nor U21892 (N_21892,N_19883,N_18610);
xor U21893 (N_21893,N_18855,N_18933);
and U21894 (N_21894,N_18604,N_18386);
and U21895 (N_21895,N_19510,N_18296);
nand U21896 (N_21896,N_18567,N_19392);
and U21897 (N_21897,N_18520,N_19209);
and U21898 (N_21898,N_18725,N_19292);
or U21899 (N_21899,N_19266,N_18624);
or U21900 (N_21900,N_19251,N_18274);
and U21901 (N_21901,N_19293,N_19902);
and U21902 (N_21902,N_19556,N_19592);
nand U21903 (N_21903,N_19717,N_19099);
nor U21904 (N_21904,N_19979,N_18981);
nor U21905 (N_21905,N_19833,N_19105);
and U21906 (N_21906,N_18794,N_18632);
or U21907 (N_21907,N_19286,N_19070);
or U21908 (N_21908,N_19582,N_19499);
nand U21909 (N_21909,N_18158,N_18172);
or U21910 (N_21910,N_19057,N_19657);
nor U21911 (N_21911,N_19655,N_19724);
xnor U21912 (N_21912,N_19231,N_18814);
and U21913 (N_21913,N_18669,N_19023);
or U21914 (N_21914,N_19502,N_19847);
or U21915 (N_21915,N_18196,N_18260);
nor U21916 (N_21916,N_18149,N_18933);
xnor U21917 (N_21917,N_18233,N_18773);
nand U21918 (N_21918,N_19789,N_19241);
nand U21919 (N_21919,N_19102,N_18422);
nand U21920 (N_21920,N_18220,N_19644);
and U21921 (N_21921,N_18412,N_19926);
and U21922 (N_21922,N_18698,N_18558);
nand U21923 (N_21923,N_19243,N_18589);
xnor U21924 (N_21924,N_19777,N_19693);
and U21925 (N_21925,N_18911,N_19340);
or U21926 (N_21926,N_19581,N_18973);
nand U21927 (N_21927,N_19541,N_19543);
xor U21928 (N_21928,N_19402,N_18999);
xnor U21929 (N_21929,N_19262,N_19693);
or U21930 (N_21930,N_18227,N_19198);
or U21931 (N_21931,N_18267,N_18673);
nand U21932 (N_21932,N_18923,N_18998);
xor U21933 (N_21933,N_18823,N_19987);
xnor U21934 (N_21934,N_19065,N_18270);
nor U21935 (N_21935,N_19705,N_18932);
and U21936 (N_21936,N_19790,N_18524);
and U21937 (N_21937,N_19477,N_19306);
and U21938 (N_21938,N_18015,N_19435);
nand U21939 (N_21939,N_18515,N_19351);
nor U21940 (N_21940,N_19842,N_19330);
and U21941 (N_21941,N_19474,N_18311);
and U21942 (N_21942,N_19813,N_18541);
xnor U21943 (N_21943,N_18959,N_19442);
nor U21944 (N_21944,N_19759,N_19233);
nor U21945 (N_21945,N_19147,N_19157);
nand U21946 (N_21946,N_19355,N_18355);
nor U21947 (N_21947,N_18859,N_19003);
or U21948 (N_21948,N_18579,N_19893);
nor U21949 (N_21949,N_19275,N_18890);
nand U21950 (N_21950,N_19634,N_18564);
nand U21951 (N_21951,N_18959,N_19609);
and U21952 (N_21952,N_18744,N_18419);
nor U21953 (N_21953,N_19570,N_18331);
nor U21954 (N_21954,N_19905,N_19034);
nand U21955 (N_21955,N_19910,N_18464);
or U21956 (N_21956,N_19654,N_18000);
xor U21957 (N_21957,N_19037,N_19705);
xnor U21958 (N_21958,N_19494,N_19601);
nand U21959 (N_21959,N_18978,N_18300);
nor U21960 (N_21960,N_18937,N_19493);
or U21961 (N_21961,N_18922,N_19246);
nor U21962 (N_21962,N_19647,N_18645);
nand U21963 (N_21963,N_19567,N_18995);
or U21964 (N_21964,N_18202,N_19986);
nor U21965 (N_21965,N_19861,N_19167);
nand U21966 (N_21966,N_18596,N_19960);
or U21967 (N_21967,N_18375,N_19446);
nor U21968 (N_21968,N_19397,N_19745);
xor U21969 (N_21969,N_18576,N_18032);
nor U21970 (N_21970,N_19356,N_19449);
nor U21971 (N_21971,N_19267,N_18250);
nor U21972 (N_21972,N_18137,N_19819);
nand U21973 (N_21973,N_19561,N_18806);
or U21974 (N_21974,N_19166,N_19912);
nand U21975 (N_21975,N_19443,N_19227);
nor U21976 (N_21976,N_18262,N_19155);
or U21977 (N_21977,N_19560,N_18245);
and U21978 (N_21978,N_18240,N_19215);
and U21979 (N_21979,N_18816,N_19430);
or U21980 (N_21980,N_18642,N_19716);
nor U21981 (N_21981,N_18796,N_19256);
or U21982 (N_21982,N_18587,N_18716);
nor U21983 (N_21983,N_19061,N_19472);
xor U21984 (N_21984,N_18380,N_19093);
or U21985 (N_21985,N_19987,N_18217);
and U21986 (N_21986,N_18081,N_19409);
nand U21987 (N_21987,N_19598,N_18898);
xnor U21988 (N_21988,N_19582,N_18954);
nand U21989 (N_21989,N_19819,N_18727);
and U21990 (N_21990,N_19551,N_19798);
and U21991 (N_21991,N_18994,N_18785);
xor U21992 (N_21992,N_19029,N_18101);
and U21993 (N_21993,N_19148,N_18212);
nand U21994 (N_21994,N_19381,N_18877);
xor U21995 (N_21995,N_19046,N_19974);
xor U21996 (N_21996,N_18194,N_18074);
or U21997 (N_21997,N_18922,N_18976);
nor U21998 (N_21998,N_18012,N_19213);
nor U21999 (N_21999,N_18352,N_19305);
or U22000 (N_22000,N_20498,N_20304);
nor U22001 (N_22001,N_21501,N_21992);
xor U22002 (N_22002,N_20683,N_21449);
and U22003 (N_22003,N_20710,N_20042);
and U22004 (N_22004,N_20962,N_21628);
nand U22005 (N_22005,N_20605,N_20456);
nor U22006 (N_22006,N_21728,N_20355);
or U22007 (N_22007,N_21503,N_20813);
or U22008 (N_22008,N_20977,N_20271);
xor U22009 (N_22009,N_21465,N_21004);
nor U22010 (N_22010,N_21622,N_21869);
or U22011 (N_22011,N_20628,N_20237);
nand U22012 (N_22012,N_20442,N_20814);
xnor U22013 (N_22013,N_21643,N_21597);
nor U22014 (N_22014,N_21020,N_20365);
or U22015 (N_22015,N_21419,N_20689);
nand U22016 (N_22016,N_21873,N_21408);
xor U22017 (N_22017,N_21448,N_21749);
and U22018 (N_22018,N_21730,N_20255);
nor U22019 (N_22019,N_20286,N_20380);
or U22020 (N_22020,N_21743,N_20172);
or U22021 (N_22021,N_20862,N_21195);
xnor U22022 (N_22022,N_20161,N_21192);
or U22023 (N_22023,N_21005,N_21126);
or U22024 (N_22024,N_21470,N_21634);
nor U22025 (N_22025,N_20815,N_20030);
and U22026 (N_22026,N_21085,N_21674);
nor U22027 (N_22027,N_20972,N_20690);
or U22028 (N_22028,N_21318,N_20546);
or U22029 (N_22029,N_21473,N_21074);
and U22030 (N_22030,N_20553,N_21003);
or U22031 (N_22031,N_21496,N_21573);
nand U22032 (N_22032,N_21920,N_20795);
xnor U22033 (N_22033,N_21861,N_21185);
xnor U22034 (N_22034,N_20412,N_21064);
or U22035 (N_22035,N_20706,N_20408);
xnor U22036 (N_22036,N_21859,N_21351);
and U22037 (N_22037,N_20336,N_20407);
nor U22038 (N_22038,N_20115,N_21407);
or U22039 (N_22039,N_21245,N_20671);
and U22040 (N_22040,N_20673,N_20726);
nand U22041 (N_22041,N_21693,N_20481);
nor U22042 (N_22042,N_20718,N_21598);
nand U22043 (N_22043,N_20174,N_21355);
and U22044 (N_22044,N_20419,N_21427);
and U22045 (N_22045,N_21441,N_21250);
xnor U22046 (N_22046,N_21849,N_20214);
or U22047 (N_22047,N_21309,N_20542);
nand U22048 (N_22048,N_21812,N_21115);
nand U22049 (N_22049,N_20005,N_21369);
nor U22050 (N_22050,N_21517,N_21008);
nand U22051 (N_22051,N_21667,N_20952);
or U22052 (N_22052,N_21048,N_21977);
or U22053 (N_22053,N_20845,N_21684);
nor U22054 (N_22054,N_21118,N_21970);
nand U22055 (N_22055,N_21746,N_20200);
or U22056 (N_22056,N_21392,N_20154);
or U22057 (N_22057,N_20538,N_21299);
nand U22058 (N_22058,N_20675,N_21376);
nand U22059 (N_22059,N_21854,N_21153);
nand U22060 (N_22060,N_21577,N_20289);
and U22061 (N_22061,N_21941,N_21343);
or U22062 (N_22062,N_21090,N_20729);
or U22063 (N_22063,N_21150,N_21719);
nand U22064 (N_22064,N_20034,N_21574);
nor U22065 (N_22065,N_21155,N_21949);
xnor U22066 (N_22066,N_20211,N_20253);
nor U22067 (N_22067,N_20478,N_21404);
or U22068 (N_22068,N_20556,N_21214);
and U22069 (N_22069,N_21362,N_21616);
or U22070 (N_22070,N_20668,N_21678);
or U22071 (N_22071,N_20396,N_20300);
or U22072 (N_22072,N_21895,N_21896);
nor U22073 (N_22073,N_21261,N_21219);
nor U22074 (N_22074,N_21872,N_21151);
nor U22075 (N_22075,N_20804,N_21946);
nand U22076 (N_22076,N_21224,N_20399);
nor U22077 (N_22077,N_20133,N_20522);
xnor U22078 (N_22078,N_20111,N_21035);
xor U22079 (N_22079,N_21805,N_20132);
or U22080 (N_22080,N_21971,N_21531);
and U22081 (N_22081,N_20341,N_21753);
xnor U22082 (N_22082,N_20142,N_20618);
or U22083 (N_22083,N_21511,N_21609);
nor U22084 (N_22084,N_20947,N_20185);
or U22085 (N_22085,N_21852,N_20513);
and U22086 (N_22086,N_20526,N_21669);
or U22087 (N_22087,N_21129,N_20489);
or U22088 (N_22088,N_21336,N_20642);
nor U22089 (N_22089,N_21714,N_21402);
or U22090 (N_22090,N_20505,N_20598);
or U22091 (N_22091,N_20896,N_20960);
nor U22092 (N_22092,N_20811,N_21038);
or U22093 (N_22093,N_20359,N_20208);
nor U22094 (N_22094,N_21122,N_21468);
or U22095 (N_22095,N_20997,N_21477);
nor U22096 (N_22096,N_20181,N_20721);
nor U22097 (N_22097,N_20741,N_20917);
nor U22098 (N_22098,N_21796,N_20897);
nor U22099 (N_22099,N_21989,N_21611);
nor U22100 (N_22100,N_20469,N_21990);
xnor U22101 (N_22101,N_20383,N_21530);
and U22102 (N_22102,N_21256,N_20901);
xor U22103 (N_22103,N_20892,N_21056);
or U22104 (N_22104,N_20207,N_21641);
nand U22105 (N_22105,N_20096,N_20603);
and U22106 (N_22106,N_21579,N_21799);
nor U22107 (N_22107,N_20939,N_21043);
and U22108 (N_22108,N_20557,N_21152);
nand U22109 (N_22109,N_21067,N_20371);
xnor U22110 (N_22110,N_21569,N_20678);
nand U22111 (N_22111,N_20338,N_20606);
nand U22112 (N_22112,N_21270,N_21361);
xnor U22113 (N_22113,N_20998,N_20390);
xor U22114 (N_22114,N_21509,N_20744);
and U22115 (N_22115,N_20982,N_20504);
and U22116 (N_22116,N_21222,N_21752);
nand U22117 (N_22117,N_20309,N_21167);
nand U22118 (N_22118,N_20876,N_21472);
xor U22119 (N_22119,N_21385,N_21239);
xnor U22120 (N_22120,N_20477,N_20078);
nor U22121 (N_22121,N_21527,N_21938);
or U22122 (N_22122,N_20613,N_20331);
nand U22123 (N_22123,N_21398,N_21191);
or U22124 (N_22124,N_21238,N_21211);
nor U22125 (N_22125,N_20316,N_21323);
nor U22126 (N_22126,N_20523,N_20107);
nor U22127 (N_22127,N_20621,N_21864);
xnor U22128 (N_22128,N_20296,N_20311);
nand U22129 (N_22129,N_20994,N_20752);
nor U22130 (N_22130,N_21958,N_20209);
or U22131 (N_22131,N_21105,N_20910);
nand U22132 (N_22132,N_21025,N_21367);
or U22133 (N_22133,N_20785,N_20935);
nor U22134 (N_22134,N_20828,N_21178);
nor U22135 (N_22135,N_21237,N_20632);
or U22136 (N_22136,N_20017,N_20413);
and U22137 (N_22137,N_20362,N_20554);
or U22138 (N_22138,N_21965,N_20758);
or U22139 (N_22139,N_20152,N_21866);
and U22140 (N_22140,N_20946,N_21042);
and U22141 (N_22141,N_21326,N_21246);
nor U22142 (N_22142,N_20568,N_20567);
nor U22143 (N_22143,N_21306,N_20048);
nand U22144 (N_22144,N_21533,N_21773);
xnor U22145 (N_22145,N_21443,N_21140);
or U22146 (N_22146,N_21423,N_20130);
xor U22147 (N_22147,N_21974,N_20833);
and U22148 (N_22148,N_20225,N_20645);
and U22149 (N_22149,N_20558,N_21280);
nand U22150 (N_22150,N_21430,N_21750);
nand U22151 (N_22151,N_21633,N_21350);
xor U22152 (N_22152,N_21547,N_20178);
or U22153 (N_22153,N_20416,N_20528);
nor U22154 (N_22154,N_20614,N_20855);
and U22155 (N_22155,N_21613,N_21006);
and U22156 (N_22156,N_20691,N_21127);
nor U22157 (N_22157,N_20076,N_20491);
or U22158 (N_22158,N_20285,N_20870);
and U22159 (N_22159,N_21851,N_21329);
nor U22160 (N_22160,N_20943,N_20024);
xnor U22161 (N_22161,N_20850,N_20375);
nand U22162 (N_22162,N_21998,N_20669);
nand U22163 (N_22163,N_20098,N_21434);
or U22164 (N_22164,N_21291,N_20584);
nor U22165 (N_22165,N_21128,N_20025);
nor U22166 (N_22166,N_20288,N_21037);
nand U22167 (N_22167,N_21662,N_21297);
and U22168 (N_22168,N_21903,N_20484);
or U22169 (N_22169,N_20890,N_20422);
and U22170 (N_22170,N_21700,N_20630);
nand U22171 (N_22171,N_20770,N_20596);
nor U22172 (N_22172,N_21725,N_21591);
xnor U22173 (N_22173,N_21007,N_20378);
and U22174 (N_22174,N_21391,N_21097);
nand U22175 (N_22175,N_20431,N_20873);
xnor U22176 (N_22176,N_20908,N_21695);
and U22177 (N_22177,N_20751,N_21396);
and U22178 (N_22178,N_20266,N_21439);
or U22179 (N_22179,N_21934,N_21915);
and U22180 (N_22180,N_21411,N_20747);
and U22181 (N_22181,N_20900,N_21196);
or U22182 (N_22182,N_20806,N_21108);
or U22183 (N_22183,N_21138,N_20435);
nor U22184 (N_22184,N_20434,N_21790);
or U22185 (N_22185,N_20641,N_21926);
or U22186 (N_22186,N_20506,N_21855);
or U22187 (N_22187,N_21368,N_20019);
xor U22188 (N_22188,N_20634,N_20427);
nor U22189 (N_22189,N_21401,N_20291);
or U22190 (N_22190,N_20129,N_20622);
or U22191 (N_22191,N_21156,N_21959);
nor U22192 (N_22192,N_20525,N_20376);
or U22193 (N_22193,N_20458,N_20916);
nand U22194 (N_22194,N_20791,N_21844);
nand U22195 (N_22195,N_21980,N_20457);
nand U22196 (N_22196,N_21254,N_20953);
nand U22197 (N_22197,N_20032,N_21302);
xnor U22198 (N_22198,N_21703,N_21400);
or U22199 (N_22199,N_20439,N_20945);
nor U22200 (N_22200,N_20308,N_21635);
xnor U22201 (N_22201,N_20186,N_20961);
or U22202 (N_22202,N_20466,N_20921);
nand U22203 (N_22203,N_20570,N_20905);
xor U22204 (N_22204,N_21739,N_21661);
or U22205 (N_22205,N_21491,N_20595);
nor U22206 (N_22206,N_21751,N_21894);
or U22207 (N_22207,N_21241,N_20702);
or U22208 (N_22208,N_21555,N_21819);
nand U22209 (N_22209,N_21966,N_21943);
xnor U22210 (N_22210,N_20500,N_20834);
and U22211 (N_22211,N_20305,N_20841);
or U22212 (N_22212,N_20049,N_21672);
xnor U22213 (N_22213,N_21809,N_21850);
xor U22214 (N_22214,N_21708,N_21077);
nor U22215 (N_22215,N_21079,N_20600);
nor U22216 (N_22216,N_21808,N_21865);
nand U22217 (N_22217,N_20112,N_20609);
xor U22218 (N_22218,N_21409,N_21642);
xnor U22219 (N_22219,N_21467,N_20821);
nand U22220 (N_22220,N_21699,N_20263);
nor U22221 (N_22221,N_20650,N_20432);
and U22222 (N_22222,N_21052,N_20626);
xor U22223 (N_22223,N_20927,N_21029);
and U22224 (N_22224,N_21879,N_20170);
nand U22225 (N_22225,N_20321,N_20313);
xnor U22226 (N_22226,N_20347,N_20382);
or U22227 (N_22227,N_20050,N_20459);
or U22228 (N_22228,N_20965,N_21871);
or U22229 (N_22229,N_20087,N_21081);
nor U22230 (N_22230,N_20323,N_20242);
and U22231 (N_22231,N_20144,N_20307);
and U22232 (N_22232,N_21164,N_20410);
nand U22233 (N_22233,N_20685,N_20543);
and U22234 (N_22234,N_21015,N_21050);
and U22235 (N_22235,N_20631,N_20837);
xnor U22236 (N_22236,N_21310,N_21701);
or U22237 (N_22237,N_20232,N_20889);
nand U22238 (N_22238,N_20276,N_21656);
or U22239 (N_22239,N_20386,N_21471);
and U22240 (N_22240,N_21294,N_21199);
nand U22241 (N_22241,N_21390,N_21353);
nand U22242 (N_22242,N_20428,N_21110);
xnor U22243 (N_22243,N_20056,N_20635);
and U22244 (N_22244,N_21774,N_20665);
and U22245 (N_22245,N_21452,N_20333);
and U22246 (N_22246,N_21308,N_21464);
xor U22247 (N_22247,N_20501,N_20817);
and U22248 (N_22248,N_20773,N_20495);
or U22249 (N_22249,N_21093,N_21381);
or U22250 (N_22250,N_21540,N_21180);
xnor U22251 (N_22251,N_21515,N_21431);
and U22252 (N_22252,N_21826,N_20767);
nor U22253 (N_22253,N_21242,N_20353);
xor U22254 (N_22254,N_21157,N_21829);
nand U22255 (N_22255,N_20951,N_21897);
nand U22256 (N_22256,N_21820,N_20166);
or U22257 (N_22257,N_20497,N_21220);
or U22258 (N_22258,N_20586,N_21145);
nand U22259 (N_22259,N_20394,N_20853);
and U22260 (N_22260,N_21546,N_20964);
nor U22261 (N_22261,N_21276,N_20616);
and U22262 (N_22262,N_20881,N_20444);
xnor U22263 (N_22263,N_20448,N_20120);
nand U22264 (N_22264,N_21717,N_21010);
or U22265 (N_22265,N_21779,N_21262);
nor U22266 (N_22266,N_21541,N_21818);
and U22267 (N_22267,N_20589,N_20282);
or U22268 (N_22268,N_20737,N_21679);
and U22269 (N_22269,N_21715,N_20661);
xnor U22270 (N_22270,N_21558,N_20297);
or U22271 (N_22271,N_20933,N_20083);
nand U22272 (N_22272,N_21563,N_21560);
nor U22273 (N_22273,N_20023,N_21993);
and U22274 (N_22274,N_21047,N_20093);
or U22275 (N_22275,N_20011,N_20337);
xnor U22276 (N_22276,N_20617,N_20189);
and U22277 (N_22277,N_20854,N_20453);
nand U22278 (N_22278,N_20753,N_21620);
and U22279 (N_22279,N_20342,N_20080);
or U22280 (N_22280,N_21028,N_20016);
nand U22281 (N_22281,N_20026,N_21756);
nor U22282 (N_22282,N_20660,N_21916);
and U22283 (N_22283,N_20540,N_20739);
nand U22284 (N_22284,N_21320,N_21566);
and U22285 (N_22285,N_21552,N_21098);
nor U22286 (N_22286,N_21636,N_20438);
nand U22287 (N_22287,N_21416,N_21522);
and U22288 (N_22288,N_21482,N_21032);
xnor U22289 (N_22289,N_21133,N_21960);
and U22290 (N_22290,N_21248,N_20891);
xnor U22291 (N_22291,N_20638,N_21782);
and U22292 (N_22292,N_20217,N_20867);
and U22293 (N_22293,N_20693,N_20629);
nor U22294 (N_22294,N_21836,N_20437);
nand U22295 (N_22295,N_20141,N_21041);
xor U22296 (N_22296,N_21065,N_20510);
and U22297 (N_22297,N_20984,N_20717);
nand U22298 (N_22298,N_21957,N_20145);
nor U22299 (N_22299,N_21272,N_20680);
or U22300 (N_22300,N_20421,N_20010);
and U22301 (N_22301,N_20919,N_21901);
or U22302 (N_22302,N_21251,N_20797);
nand U22303 (N_22303,N_21979,N_21475);
nor U22304 (N_22304,N_21424,N_21617);
xnor U22305 (N_22305,N_21741,N_21762);
and U22306 (N_22306,N_21914,N_21824);
nor U22307 (N_22307,N_20480,N_21596);
and U22308 (N_22308,N_20351,N_20732);
nand U22309 (N_22309,N_20712,N_20159);
nand U22310 (N_22310,N_21189,N_20681);
xor U22311 (N_22311,N_20201,N_21557);
nor U22312 (N_22312,N_20820,N_20877);
nor U22313 (N_22313,N_21217,N_20708);
xor U22314 (N_22314,N_20793,N_20155);
xor U22315 (N_22315,N_21313,N_21520);
or U22316 (N_22316,N_21426,N_21040);
nand U22317 (N_22317,N_20511,N_20515);
nand U22318 (N_22318,N_21259,N_20268);
nor U22319 (N_22319,N_21581,N_20358);
nor U22320 (N_22320,N_21228,N_21322);
or U22321 (N_22321,N_21660,N_21583);
nand U22322 (N_22322,N_20167,N_20473);
and U22323 (N_22323,N_21521,N_21646);
xnor U22324 (N_22324,N_20949,N_21462);
nand U22325 (N_22325,N_20195,N_20700);
nand U22326 (N_22326,N_20045,N_21456);
and U22327 (N_22327,N_21794,N_21691);
and U22328 (N_22328,N_20157,N_21778);
nor U22329 (N_22329,N_20688,N_21139);
xnor U22330 (N_22330,N_20588,N_20925);
nand U22331 (N_22331,N_20139,N_20607);
nor U22332 (N_22332,N_20969,N_20583);
nand U22333 (N_22333,N_20363,N_21011);
xnor U22334 (N_22334,N_21882,N_20047);
and U22335 (N_22335,N_20381,N_20138);
xnor U22336 (N_22336,N_21365,N_21627);
nor U22337 (N_22337,N_20411,N_21344);
and U22338 (N_22338,N_21223,N_20251);
or U22339 (N_22339,N_20649,N_20731);
xor U22340 (N_22340,N_21083,N_21201);
xnor U22341 (N_22341,N_21648,N_20991);
or U22342 (N_22342,N_21594,N_21202);
nand U22343 (N_22343,N_20875,N_20981);
and U22344 (N_22344,N_20475,N_21921);
xnor U22345 (N_22345,N_21379,N_21688);
nand U22346 (N_22346,N_20198,N_21184);
nor U22347 (N_22347,N_21208,N_20488);
nor U22348 (N_22348,N_20109,N_20103);
and U22349 (N_22349,N_21564,N_20587);
nand U22350 (N_22350,N_20401,N_21630);
xor U22351 (N_22351,N_20524,N_20020);
and U22352 (N_22352,N_20999,N_20552);
xnor U22353 (N_22353,N_20277,N_20403);
and U22354 (N_22354,N_21961,N_21162);
xor U22355 (N_22355,N_21789,N_20108);
and U22356 (N_22356,N_20822,N_20959);
and U22357 (N_22357,N_21282,N_21828);
nand U22358 (N_22358,N_21289,N_21726);
nand U22359 (N_22359,N_21504,N_21802);
or U22360 (N_22360,N_20090,N_21166);
nand U22361 (N_22361,N_20633,N_21822);
nand U22362 (N_22362,N_21233,N_20377);
or U22363 (N_22363,N_21252,N_20116);
nor U22364 (N_22364,N_20188,N_21625);
xor U22365 (N_22365,N_21507,N_21094);
nand U22366 (N_22366,N_21922,N_20101);
xnor U22367 (N_22367,N_20924,N_20212);
and U22368 (N_22368,N_20730,N_20406);
or U22369 (N_22369,N_21158,N_21478);
xor U22370 (N_22370,N_20716,N_21523);
nand U22371 (N_22371,N_20865,N_20840);
nor U22372 (N_22372,N_21994,N_20073);
and U22373 (N_22373,N_21638,N_21623);
or U22374 (N_22374,N_20923,N_20836);
xor U22375 (N_22375,N_21243,N_21445);
nand U22376 (N_22376,N_21493,N_20465);
nor U22377 (N_22377,N_21497,N_20179);
and U22378 (N_22378,N_20888,N_20886);
nand U22379 (N_22379,N_21375,N_20696);
nor U22380 (N_22380,N_20171,N_20199);
nand U22381 (N_22381,N_20637,N_21709);
nor U22382 (N_22382,N_20222,N_20252);
nand U22383 (N_22383,N_20372,N_20326);
nor U22384 (N_22384,N_21516,N_21944);
or U22385 (N_22385,N_20162,N_20483);
and U22386 (N_22386,N_20679,N_21919);
nor U22387 (N_22387,N_21374,N_20978);
and U22388 (N_22388,N_21706,N_20128);
nor U22389 (N_22389,N_20593,N_21486);
and U22390 (N_22390,N_21455,N_21311);
or U22391 (N_22391,N_20423,N_21053);
nor U22392 (N_22392,N_20127,N_20029);
nand U22393 (N_22393,N_20125,N_21589);
xnor U22394 (N_22394,N_20560,N_21413);
or U22395 (N_22395,N_21466,N_20364);
or U22396 (N_22396,N_21345,N_21877);
xnor U22397 (N_22397,N_21784,N_20234);
and U22398 (N_22398,N_21543,N_20893);
xor U22399 (N_22399,N_20153,N_21529);
nor U22400 (N_22400,N_21595,N_20749);
or U22401 (N_22401,N_21724,N_21176);
nand U22402 (N_22402,N_20829,N_21489);
xor U22403 (N_22403,N_20223,N_21287);
nand U22404 (N_22404,N_21666,N_20393);
nor U22405 (N_22405,N_20137,N_20265);
or U22406 (N_22406,N_21410,N_20878);
xnor U22407 (N_22407,N_21207,N_21985);
and U22408 (N_22408,N_20779,N_20656);
xnor U22409 (N_22409,N_20714,N_21347);
and U22410 (N_22410,N_20544,N_20824);
xnor U22411 (N_22411,N_20314,N_20248);
xor U22412 (N_22412,N_21858,N_21403);
nor U22413 (N_22413,N_20985,N_21745);
nand U22414 (N_22414,N_21227,N_21874);
nand U22415 (N_22415,N_21253,N_20180);
nand U22416 (N_22416,N_21783,N_20738);
nand U22417 (N_22417,N_20537,N_21435);
xor U22418 (N_22418,N_20452,N_20963);
or U22419 (N_22419,N_21317,N_20135);
and U22420 (N_22420,N_20264,N_20988);
nor U22421 (N_22421,N_21476,N_21490);
or U22422 (N_22422,N_20869,N_20445);
nand U22423 (N_22423,N_21049,N_21170);
nand U22424 (N_22424,N_21316,N_20119);
xor U22425 (N_22425,N_20451,N_20204);
and U22426 (N_22426,N_21168,N_20727);
and U22427 (N_22427,N_21969,N_20315);
and U22428 (N_22428,N_20864,N_20360);
and U22429 (N_22429,N_21837,N_20312);
xor U22430 (N_22430,N_21101,N_21652);
and U22431 (N_22431,N_20194,N_20227);
xnor U22432 (N_22432,N_21319,N_20259);
or U22433 (N_22433,N_20858,N_20646);
xnor U22434 (N_22434,N_21740,N_21687);
or U22435 (N_22435,N_21061,N_21017);
nor U22436 (N_22436,N_20851,N_21981);
or U22437 (N_22437,N_21335,N_20958);
nand U22438 (N_22438,N_21880,N_20446);
xor U22439 (N_22439,N_20470,N_21770);
nand U22440 (N_22440,N_21767,N_21247);
nor U22441 (N_22441,N_20404,N_20398);
or U22442 (N_22442,N_20368,N_21255);
nand U22443 (N_22443,N_20832,N_20503);
and U22444 (N_22444,N_20932,N_20165);
and U22445 (N_22445,N_20579,N_20374);
nor U22446 (N_22446,N_20856,N_20018);
and U22447 (N_22447,N_21014,N_21172);
nand U22448 (N_22448,N_20694,N_20907);
nand U22449 (N_22449,N_21288,N_20941);
and U22450 (N_22450,N_20574,N_20027);
nand U22451 (N_22451,N_20561,N_20490);
nand U22452 (N_22452,N_21063,N_20676);
xor U22453 (N_22453,N_21279,N_21103);
or U22454 (N_22454,N_20105,N_20303);
and U22455 (N_22455,N_21442,N_20361);
xnor U22456 (N_22456,N_21481,N_20789);
or U22457 (N_22457,N_20827,N_20149);
and U22458 (N_22458,N_21117,N_20415);
and U22459 (N_22459,N_20966,N_20530);
nor U22460 (N_22460,N_21425,N_21328);
nand U22461 (N_22461,N_21833,N_21022);
xor U22462 (N_22462,N_20674,N_20043);
and U22463 (N_22463,N_20722,N_20549);
xor U22464 (N_22464,N_21976,N_21120);
and U22465 (N_22465,N_20648,N_20755);
nor U22466 (N_22466,N_21235,N_21967);
xnor U22467 (N_22467,N_21664,N_21163);
nor U22468 (N_22468,N_21058,N_20102);
or U22469 (N_22469,N_21654,N_20550);
and U22470 (N_22470,N_21078,N_20601);
or U22471 (N_22471,N_20254,N_20033);
nor U22472 (N_22472,N_21888,N_20736);
and U22473 (N_22473,N_21856,N_20474);
nand U22474 (N_22474,N_21825,N_20912);
nand U22475 (N_22475,N_20909,N_21806);
and U22476 (N_22476,N_20514,N_21811);
nor U22477 (N_22477,N_21173,N_21898);
or U22478 (N_22478,N_20104,N_20492);
or U22479 (N_22479,N_20136,N_21334);
nor U22480 (N_22480,N_21187,N_21668);
nor U22481 (N_22481,N_21514,N_20006);
xor U22482 (N_22482,N_21137,N_20838);
nor U22483 (N_22483,N_20147,N_20521);
or U22484 (N_22484,N_20914,N_21354);
nor U22485 (N_22485,N_20723,N_21612);
nor U22486 (N_22486,N_20610,N_20564);
or U22487 (N_22487,N_20482,N_21054);
nand U22488 (N_22488,N_20110,N_21030);
and U22489 (N_22489,N_21146,N_20748);
nand U22490 (N_22490,N_20235,N_21876);
or U22491 (N_22491,N_20742,N_20258);
nor U22492 (N_22492,N_21937,N_20662);
nand U22493 (N_22493,N_21188,N_21136);
or U22494 (N_22494,N_20322,N_21846);
or U22495 (N_22495,N_21565,N_20059);
nor U22496 (N_22496,N_21084,N_20290);
nor U22497 (N_22497,N_20384,N_20468);
nor U22498 (N_22498,N_21996,N_21653);
nor U22499 (N_22499,N_21075,N_21154);
nand U22500 (N_22500,N_20247,N_21225);
nor U22501 (N_22501,N_20215,N_20783);
and U22502 (N_22502,N_21119,N_20895);
nor U22503 (N_22503,N_21382,N_20839);
nand U22504 (N_22504,N_20983,N_20913);
and U22505 (N_22505,N_21265,N_21575);
xor U22506 (N_22506,N_20654,N_21983);
nand U22507 (N_22507,N_21099,N_21907);
nor U22508 (N_22508,N_20395,N_20069);
nor U22509 (N_22509,N_20343,N_21925);
and U22510 (N_22510,N_20099,N_20539);
or U22511 (N_22511,N_21776,N_21890);
xnor U22512 (N_22512,N_21655,N_20046);
and U22513 (N_22513,N_21458,N_21621);
and U22514 (N_22514,N_21102,N_21795);
nor U22515 (N_22515,N_21206,N_20619);
nor U22516 (N_22516,N_21436,N_21518);
or U22517 (N_22517,N_21830,N_20799);
nand U22518 (N_22518,N_20863,N_20257);
nand U22519 (N_22519,N_21305,N_20666);
xor U22520 (N_22520,N_20267,N_20778);
or U22521 (N_22521,N_20699,N_21912);
or U22522 (N_22522,N_21087,N_20318);
nand U22523 (N_22523,N_20812,N_20192);
nor U22524 (N_22524,N_21232,N_21902);
xnor U22525 (N_22525,N_20819,N_21132);
and U22526 (N_22526,N_20191,N_21339);
nor U22527 (N_22527,N_21013,N_21694);
nor U22528 (N_22528,N_20464,N_21685);
and U22529 (N_22529,N_20868,N_20986);
nand U22530 (N_22530,N_21096,N_20274);
or U22531 (N_22531,N_21720,N_20885);
nand U22532 (N_22532,N_21624,N_21578);
nand U22533 (N_22533,N_20571,N_21731);
xor U22534 (N_22534,N_20509,N_21973);
or U22535 (N_22535,N_21421,N_20807);
xnor U22536 (N_22536,N_21759,N_21815);
nor U22537 (N_22537,N_20805,N_21771);
nand U22538 (N_22538,N_20565,N_21198);
xor U22539 (N_22539,N_20231,N_21590);
and U22540 (N_22540,N_21657,N_21019);
and U22541 (N_22541,N_20085,N_21349);
nor U22542 (N_22542,N_20756,N_20803);
xnor U22543 (N_22543,N_21307,N_21352);
nand U22544 (N_22544,N_21733,N_21927);
or U22545 (N_22545,N_20894,N_20930);
xnor U22546 (N_22546,N_21904,N_21519);
and U22547 (N_22547,N_21658,N_21502);
xnor U22548 (N_22548,N_20038,N_21716);
and U22549 (N_22549,N_20599,N_21459);
xnor U22550 (N_22550,N_20608,N_21513);
nand U22551 (N_22551,N_21619,N_20954);
nor U22552 (N_22552,N_20580,N_21269);
nor U22553 (N_22553,N_20123,N_21559);
nor U22554 (N_22554,N_20008,N_21463);
nor U22555 (N_22555,N_20777,N_20725);
nor U22556 (N_22556,N_21860,N_21281);
or U22557 (N_22557,N_20652,N_21364);
nand U22558 (N_22558,N_20884,N_20385);
nand U22559 (N_22559,N_21542,N_21545);
xnor U22560 (N_22560,N_20664,N_20711);
xor U22561 (N_22561,N_20672,N_21814);
and U22562 (N_22562,N_20246,N_20074);
xnor U22563 (N_22563,N_21359,N_21076);
and U22564 (N_22564,N_20117,N_20429);
and U22565 (N_22565,N_20317,N_21457);
nor U22566 (N_22566,N_21236,N_21342);
nand U22567 (N_22567,N_20091,N_20066);
nand U22568 (N_22568,N_20417,N_21234);
nand U22569 (N_22569,N_21614,N_20230);
or U22570 (N_22570,N_20575,N_21905);
or U22571 (N_22571,N_21062,N_20114);
nand U22572 (N_22572,N_20531,N_21690);
xnor U22573 (N_22573,N_21605,N_20425);
and U22574 (N_22574,N_21092,N_20971);
and U22575 (N_22575,N_21692,N_20463);
and U22576 (N_22576,N_20126,N_20433);
nor U22577 (N_22577,N_21209,N_21748);
xor U22578 (N_22578,N_20306,N_20883);
or U22579 (N_22579,N_21356,N_21060);
or U22580 (N_22580,N_21303,N_20857);
nand U22581 (N_22581,N_21689,N_20887);
and U22582 (N_22582,N_21875,N_21505);
or U22583 (N_22583,N_20790,N_21383);
nor U22584 (N_22584,N_21568,N_20944);
nand U22585 (N_22585,N_20535,N_20788);
nor U22586 (N_22586,N_20146,N_20197);
nor U22587 (N_22587,N_21673,N_21816);
and U22588 (N_22588,N_20763,N_20443);
nor U22589 (N_22589,N_21982,N_20657);
nand U22590 (N_22590,N_20182,N_20370);
nand U22591 (N_22591,N_21863,N_21378);
xnor U22592 (N_22592,N_20866,N_20345);
and U22593 (N_22593,N_21870,N_21044);
or U22594 (N_22594,N_20658,N_21592);
nor U22595 (N_22595,N_21911,N_21582);
nor U22596 (N_22596,N_20298,N_20990);
xnor U22597 (N_22597,N_20084,N_20319);
nand U22598 (N_22598,N_21567,N_21397);
xor U22599 (N_22599,N_20387,N_21488);
nand U22600 (N_22600,N_21432,N_20871);
nand U22601 (N_22601,N_20957,N_21125);
nand U22602 (N_22602,N_20004,N_21524);
nand U22603 (N_22603,N_20639,N_20344);
xor U22604 (N_22604,N_21412,N_21499);
nor U22605 (N_22605,N_21862,N_20077);
nand U22606 (N_22606,N_20229,N_20121);
and U22607 (N_22607,N_21018,N_21538);
or U22608 (N_22608,N_21535,N_21663);
and U22609 (N_22609,N_21572,N_21479);
and U22610 (N_22610,N_21615,N_20728);
xor U22611 (N_22611,N_20349,N_21988);
xor U22612 (N_22612,N_20063,N_21377);
nand U22613 (N_22613,N_20566,N_21104);
nand U22614 (N_22614,N_20151,N_20007);
xor U22615 (N_22615,N_20620,N_20054);
and U22616 (N_22616,N_20279,N_21800);
nand U22617 (N_22617,N_21405,N_21267);
and U22618 (N_22618,N_21840,N_21112);
xor U22619 (N_22619,N_21600,N_20447);
nor U22620 (N_22620,N_21460,N_21797);
nor U22621 (N_22621,N_20243,N_21696);
and U22622 (N_22622,N_21357,N_20771);
nor U22623 (N_22623,N_21955,N_20496);
nor U22624 (N_22624,N_21675,N_21024);
nor U22625 (N_22625,N_20031,N_20594);
nand U22626 (N_22626,N_21599,N_20081);
and U22627 (N_22627,N_20354,N_20843);
nand U22628 (N_22628,N_20768,N_21842);
nor U22629 (N_22629,N_21394,N_20734);
nand U22630 (N_22630,N_21372,N_21286);
nor U22631 (N_22631,N_21705,N_21031);
or U22632 (N_22632,N_20436,N_20774);
nand U22633 (N_22633,N_21544,N_21141);
or U22634 (N_22634,N_21106,N_20118);
nand U22635 (N_22635,N_20670,N_21952);
and U22636 (N_22636,N_21012,N_20562);
nor U22637 (N_22637,N_21230,N_20060);
nand U22638 (N_22638,N_20938,N_21754);
nand U22639 (N_22639,N_21179,N_20720);
xor U22640 (N_22640,N_21330,N_20541);
and U22641 (N_22641,N_21086,N_21144);
or U22642 (N_22642,N_21315,N_21414);
nand U22643 (N_22643,N_20880,N_21512);
xnor U22644 (N_22644,N_20955,N_21175);
nand U22645 (N_22645,N_21429,N_21148);
xor U22646 (N_22646,N_20213,N_20636);
xor U22647 (N_22647,N_21454,N_20070);
nor U22648 (N_22648,N_21834,N_21968);
and U22649 (N_22649,N_21525,N_21827);
nand U22650 (N_22650,N_21761,N_20825);
xnor U22651 (N_22651,N_21556,N_20507);
and U22652 (N_22652,N_20329,N_20330);
xnor U22653 (N_22653,N_20392,N_20224);
nor U22654 (N_22654,N_20992,N_21213);
xnor U22655 (N_22655,N_21301,N_21174);
nand U22656 (N_22656,N_20775,N_20373);
and U22657 (N_22657,N_20970,N_20547);
xnor U22658 (N_22658,N_21821,N_20183);
nor U22659 (N_22659,N_20177,N_20022);
nand U22660 (N_22660,N_20709,N_20461);
or U22661 (N_22661,N_20239,N_21312);
xnor U22662 (N_22662,N_20735,N_20559);
and U22663 (N_22663,N_21987,N_20061);
nor U22664 (N_22664,N_20527,N_20071);
xnor U22665 (N_22665,N_20898,N_20615);
nor U22666 (N_22666,N_21082,N_20784);
or U22667 (N_22667,N_21736,N_20611);
xor U22668 (N_22668,N_21244,N_21451);
nor U22669 (N_22669,N_20228,N_20572);
xnor U22670 (N_22670,N_21803,N_20764);
or U22671 (N_22671,N_21986,N_21755);
nand U22672 (N_22672,N_21450,N_21645);
nand U22673 (N_22673,N_21494,N_20350);
and U22674 (N_22674,N_20089,N_20519);
and U22675 (N_22675,N_21659,N_21266);
xor U22676 (N_22676,N_21857,N_20518);
nand U22677 (N_22677,N_20929,N_20980);
xor U22678 (N_22678,N_21924,N_20190);
nand U22679 (N_22679,N_21707,N_21324);
or U22680 (N_22680,N_20703,N_21216);
nor U22681 (N_22681,N_21747,N_20512);
xnor U22682 (N_22682,N_21780,N_20926);
and U22683 (N_22683,N_21147,N_20335);
nor U22684 (N_22684,N_20001,N_20906);
nor U22685 (N_22685,N_20426,N_21777);
and U22686 (N_22686,N_20339,N_21480);
or U22687 (N_22687,N_20798,N_20987);
xnor U22688 (N_22688,N_20206,N_21055);
and U22689 (N_22689,N_20454,N_21918);
nand U22690 (N_22690,N_20623,N_21721);
xnor U22691 (N_22691,N_21951,N_21212);
or U22692 (N_22692,N_20879,N_20294);
xor U22693 (N_22693,N_20036,N_20692);
and U22694 (N_22694,N_21813,N_21215);
nor U22695 (N_22695,N_21009,N_20169);
or U22696 (N_22696,N_21554,N_21095);
or U22697 (N_22697,N_20801,N_21292);
and U22698 (N_22698,N_20455,N_20830);
and U22699 (N_22699,N_21295,N_20782);
or U22700 (N_22700,N_21580,N_21991);
nor U22701 (N_22701,N_21534,N_21070);
or U22702 (N_22702,N_20920,N_20293);
or U22703 (N_22703,N_21999,N_20272);
or U22704 (N_22704,N_21210,N_20441);
or U22705 (N_22705,N_20573,N_21051);
xor U22706 (N_22706,N_20389,N_21604);
nor U22707 (N_22707,N_21964,N_21704);
or U22708 (N_22708,N_21149,N_21399);
or U22709 (N_22709,N_20140,N_21629);
xnor U22710 (N_22710,N_21893,N_20193);
nand U22711 (N_22711,N_20563,N_21562);
or U22712 (N_22712,N_20551,N_21537);
xor U22713 (N_22713,N_21735,N_21881);
and U22714 (N_22714,N_20499,N_20903);
or U22715 (N_22715,N_20122,N_20766);
and U22716 (N_22716,N_20516,N_21586);
nor U22717 (N_22717,N_21603,N_20327);
or U22718 (N_22718,N_20203,N_20948);
and U22719 (N_22719,N_20405,N_20245);
nand U22720 (N_22720,N_20578,N_20904);
and U22721 (N_22721,N_21193,N_20450);
nor U22722 (N_22722,N_21422,N_21171);
and U22723 (N_22723,N_21433,N_21792);
nand U22724 (N_22724,N_21665,N_20979);
nand U22725 (N_22725,N_21950,N_20440);
nand U22726 (N_22726,N_21742,N_21495);
or U22727 (N_22727,N_20086,N_20379);
nand U22728 (N_22728,N_20928,N_21333);
xnor U22729 (N_22729,N_20148,N_21878);
xnor U22730 (N_22730,N_21626,N_21057);
or U22731 (N_22731,N_20874,N_21899);
nor U22732 (N_22732,N_21338,N_21712);
xor U22733 (N_22733,N_20705,N_21325);
or U22734 (N_22734,N_21204,N_20075);
and U22735 (N_22735,N_21930,N_21197);
or U22736 (N_22736,N_21738,N_20647);
and U22737 (N_22737,N_20826,N_21884);
nor U22738 (N_22738,N_20035,N_21134);
nand U22739 (N_22739,N_20052,N_21929);
and U22740 (N_22740,N_21539,N_21346);
xor U22741 (N_22741,N_21231,N_20357);
nor U22742 (N_22742,N_20460,N_20911);
or U22743 (N_22743,N_21296,N_20462);
nor U22744 (N_22744,N_20719,N_21650);
nor U22745 (N_22745,N_21190,N_21034);
nand U22746 (N_22746,N_21177,N_20210);
or U22747 (N_22747,N_21670,N_20655);
nand U22748 (N_22748,N_21002,N_21393);
nand U22749 (N_22749,N_20430,N_21764);
and U22750 (N_22750,N_20967,N_20015);
and U22751 (N_22751,N_21718,N_20485);
xnor U22752 (N_22752,N_21737,N_20733);
xor U22753 (N_22753,N_20226,N_20202);
and U22754 (N_22754,N_21080,N_20695);
xnor U22755 (N_22755,N_20976,N_21159);
nor U22756 (N_22756,N_20366,N_21415);
or U22757 (N_22757,N_21606,N_21327);
and U22758 (N_22758,N_20143,N_20302);
or U22759 (N_22759,N_21887,N_21181);
or U22760 (N_22760,N_20860,N_21283);
nor U22761 (N_22761,N_21380,N_20467);
nand U22762 (N_22762,N_20014,N_20160);
xor U22763 (N_22763,N_20934,N_21066);
xnor U22764 (N_22764,N_20508,N_21440);
nor U22765 (N_22765,N_20794,N_21284);
nor U22766 (N_22766,N_20942,N_21766);
xor U22767 (N_22767,N_20013,N_21387);
nand U22768 (N_22768,N_20219,N_20156);
nand U22769 (N_22769,N_20057,N_20240);
nor U22770 (N_22770,N_21249,N_21823);
nand U22771 (N_22771,N_20769,N_21277);
or U22772 (N_22772,N_21781,N_21948);
nor U22773 (N_22773,N_20479,N_21218);
or U22774 (N_22774,N_20847,N_20848);
and U22775 (N_22775,N_20677,N_21229);
or U22776 (N_22776,N_21702,N_21910);
xor U22777 (N_22777,N_21713,N_21804);
and U22778 (N_22778,N_21576,N_21161);
nor U22779 (N_22779,N_21791,N_21113);
and U22780 (N_22780,N_21059,N_21071);
xnor U22781 (N_22781,N_21723,N_20545);
nand U22782 (N_22782,N_21274,N_20555);
nand U22783 (N_22783,N_20082,N_20659);
or U22784 (N_22784,N_21570,N_20068);
and U22785 (N_22785,N_20835,N_20707);
xor U22786 (N_22786,N_21917,N_21293);
and U22787 (N_22787,N_21632,N_21386);
nor U22788 (N_22788,N_21046,N_21226);
xnor U22789 (N_22789,N_20534,N_21532);
and U22790 (N_22790,N_21639,N_20899);
nor U22791 (N_22791,N_20597,N_20249);
or U22792 (N_22792,N_20761,N_20859);
nand U22793 (N_22793,N_21886,N_21200);
nor U22794 (N_22794,N_20260,N_20786);
and U22795 (N_22795,N_21945,N_21610);
or U22796 (N_22796,N_20088,N_20989);
nand U22797 (N_22797,N_20846,N_21817);
nor U22798 (N_22798,N_20028,N_21469);
or U22799 (N_22799,N_20241,N_20810);
xor U22800 (N_22800,N_21021,N_21848);
xor U22801 (N_22801,N_20536,N_21109);
nand U22802 (N_22802,N_20644,N_20287);
and U22803 (N_22803,N_21727,N_21258);
and U22804 (N_22804,N_21366,N_21722);
nand U22805 (N_22805,N_20802,N_20292);
or U22806 (N_22806,N_20280,N_20762);
nand U22807 (N_22807,N_20262,N_20471);
or U22808 (N_22808,N_20414,N_20486);
and U22809 (N_22809,N_20698,N_20334);
and U22810 (N_22810,N_20062,N_21314);
xnor U22811 (N_22811,N_20348,N_20950);
nor U22812 (N_22812,N_20218,N_20687);
and U22813 (N_22813,N_21549,N_21909);
or U22814 (N_22814,N_20612,N_21832);
xor U22815 (N_22815,N_21487,N_20759);
nand U22816 (N_22816,N_21954,N_20236);
xnor U22817 (N_22817,N_20332,N_21785);
nor U22818 (N_22818,N_21913,N_20882);
and U22819 (N_22819,N_20809,N_20150);
nor U22820 (N_22820,N_21121,N_20765);
xor U22821 (N_22821,N_20569,N_20533);
nor U22822 (N_22822,N_21975,N_20624);
or U22823 (N_22823,N_21143,N_20651);
nand U22824 (N_22824,N_20915,N_21417);
and U22825 (N_22825,N_21935,N_20367);
xnor U22826 (N_22826,N_21984,N_20284);
and U22827 (N_22827,N_21073,N_20502);
nand U22828 (N_22828,N_21384,N_21483);
xor U22829 (N_22829,N_21835,N_20922);
nand U22830 (N_22830,N_21373,N_21278);
nand U22831 (N_22831,N_20973,N_21775);
and U22832 (N_22832,N_21337,N_21165);
xor U22833 (N_22833,N_21275,N_20816);
or U22834 (N_22834,N_21788,N_20936);
or U22835 (N_22835,N_21710,N_20667);
or U22836 (N_22836,N_21942,N_20346);
nand U22837 (N_22837,N_20682,N_21257);
and U22838 (N_22838,N_21978,N_21682);
nor U22839 (N_22839,N_20487,N_21300);
or U22840 (N_22840,N_20055,N_21587);
or U22841 (N_22841,N_20301,N_21900);
and U22842 (N_22842,N_20772,N_21972);
xor U22843 (N_22843,N_20697,N_21221);
or U22844 (N_22844,N_21584,N_20577);
nand U22845 (N_22845,N_21111,N_20233);
and U22846 (N_22846,N_21928,N_21729);
xnor U22847 (N_22847,N_20039,N_21963);
and U22848 (N_22848,N_21602,N_21550);
and U22849 (N_22849,N_20823,N_20995);
xor U22850 (N_22850,N_21388,N_21711);
nor U22851 (N_22851,N_21114,N_20472);
nand U22852 (N_22852,N_21268,N_20548);
nand U22853 (N_22853,N_20591,N_20184);
or U22854 (N_22854,N_21885,N_21183);
nand U22855 (N_22855,N_21647,N_20106);
and U22856 (N_22856,N_20072,N_20627);
or U22857 (N_22857,N_21395,N_21169);
xor U22858 (N_22858,N_20051,N_20704);
xor U22859 (N_22859,N_20164,N_20244);
nand U22860 (N_22860,N_21528,N_21551);
xnor U22861 (N_22861,N_21607,N_20205);
and U22862 (N_22862,N_21838,N_21786);
nor U22863 (N_22863,N_21601,N_20931);
nor U22864 (N_22864,N_20064,N_21757);
nor U22865 (N_22865,N_20872,N_20173);
nand U22866 (N_22866,N_21847,N_21810);
or U22867 (N_22867,N_21765,N_20324);
or U22868 (N_22868,N_21506,N_20940);
or U22869 (N_22869,N_21360,N_21045);
nand U22870 (N_22870,N_20065,N_20269);
nand U22871 (N_22871,N_21260,N_20849);
and U22872 (N_22872,N_20400,N_20176);
xor U22873 (N_22873,N_20974,N_20079);
nand U22874 (N_22874,N_21677,N_21039);
or U22875 (N_22875,N_21906,N_21418);
and U22876 (N_22876,N_21263,N_20750);
nand U22877 (N_22877,N_20021,N_20653);
and U22878 (N_22878,N_20310,N_21160);
xor U22879 (N_22879,N_21194,N_21406);
xor U22880 (N_22880,N_21068,N_20094);
nor U22881 (N_22881,N_20808,N_21131);
nor U22882 (N_22882,N_21036,N_20067);
nor U22883 (N_22883,N_21000,N_21371);
or U22884 (N_22884,N_21732,N_20585);
xnor U22885 (N_22885,N_20602,N_20175);
nor U22886 (N_22886,N_20113,N_20746);
nor U22887 (N_22887,N_20724,N_21526);
xnor U22888 (N_22888,N_21608,N_21321);
xnor U22889 (N_22889,N_21331,N_21298);
or U22890 (N_22890,N_21023,N_20684);
or U22891 (N_22891,N_20818,N_21453);
nand U22892 (N_22892,N_20740,N_20449);
nor U22893 (N_22893,N_21348,N_20281);
xnor U22894 (N_22894,N_21588,N_20134);
or U22895 (N_22895,N_21116,N_21843);
nor U22896 (N_22896,N_21358,N_20743);
and U22897 (N_22897,N_20757,N_21908);
and U22898 (N_22898,N_21680,N_20409);
nor U22899 (N_22899,N_21088,N_21264);
or U22900 (N_22900,N_21428,N_21763);
nand U22901 (N_22901,N_21676,N_20299);
xor U22902 (N_22902,N_20273,N_20643);
xor U22903 (N_22903,N_20861,N_20012);
xnor U22904 (N_22904,N_20003,N_20275);
nand U22905 (N_22905,N_21485,N_20041);
nor U22906 (N_22906,N_20800,N_21853);
nor U22907 (N_22907,N_21548,N_20009);
and U22908 (N_22908,N_20494,N_20037);
xnor U22909 (N_22909,N_21130,N_20424);
nand U22910 (N_22910,N_20745,N_21484);
nor U22911 (N_22911,N_21341,N_21304);
nand U22912 (N_22912,N_20529,N_21768);
nand U22913 (N_22913,N_20792,N_20590);
and U22914 (N_22914,N_21123,N_20968);
nor U22915 (N_22915,N_20095,N_21363);
xor U22916 (N_22916,N_20356,N_21686);
and U22917 (N_22917,N_20221,N_20369);
nand U22918 (N_22918,N_21698,N_21923);
or U22919 (N_22919,N_21697,N_20216);
or U22920 (N_22920,N_20780,N_21240);
nor U22921 (N_22921,N_21940,N_21671);
nand U22922 (N_22922,N_21026,N_20760);
and U22923 (N_22923,N_20391,N_21135);
xor U22924 (N_22924,N_20713,N_21142);
and U22925 (N_22925,N_20975,N_20270);
xnor U22926 (N_22926,N_20781,N_20604);
nor U22927 (N_22927,N_21500,N_21585);
xor U22928 (N_22928,N_20402,N_21883);
and U22929 (N_22929,N_20196,N_21933);
nand U22930 (N_22930,N_21271,N_20776);
or U22931 (N_22931,N_20163,N_21536);
nor U22932 (N_22932,N_20100,N_20238);
nand U22933 (N_22933,N_20576,N_20295);
and U22934 (N_22934,N_21553,N_21845);
nor U22935 (N_22935,N_20397,N_20532);
nor U22936 (N_22936,N_21389,N_21498);
xnor U22937 (N_22937,N_20250,N_21340);
or U22938 (N_22938,N_21618,N_21461);
nand U22939 (N_22939,N_20993,N_20996);
nor U22940 (N_22940,N_20256,N_21124);
and U22941 (N_22941,N_21787,N_20418);
or U22942 (N_22942,N_21995,N_21793);
nor U22943 (N_22943,N_21290,N_20625);
xor U22944 (N_22944,N_21203,N_20053);
and U22945 (N_22945,N_20261,N_20352);
xor U22946 (N_22946,N_20581,N_20283);
or U22947 (N_22947,N_20320,N_21273);
nand U22948 (N_22948,N_21734,N_20918);
nor U22949 (N_22949,N_20842,N_20000);
xnor U22950 (N_22950,N_21953,N_20325);
xnor U22951 (N_22951,N_20754,N_20058);
nand U22952 (N_22952,N_20044,N_21939);
nor U22953 (N_22953,N_21892,N_21644);
or U22954 (N_22954,N_21437,N_20592);
nor U22955 (N_22955,N_20131,N_20902);
or U22956 (N_22956,N_21744,N_20517);
or U22957 (N_22957,N_21798,N_21016);
and U22958 (N_22958,N_20663,N_21839);
xor U22959 (N_22959,N_21182,N_21420);
and U22960 (N_22960,N_21069,N_21947);
and U22961 (N_22961,N_21867,N_20340);
or U22962 (N_22962,N_21593,N_20278);
nand U22963 (N_22963,N_21107,N_21956);
nand U22964 (N_22964,N_21571,N_21100);
xor U22965 (N_22965,N_21649,N_21438);
and U22966 (N_22966,N_20582,N_20388);
xnor U22967 (N_22967,N_20701,N_20640);
xnor U22968 (N_22968,N_21651,N_20844);
or U22969 (N_22969,N_21492,N_20168);
and U22970 (N_22970,N_21683,N_21332);
xnor U22971 (N_22971,N_21474,N_20040);
xnor U22972 (N_22972,N_21962,N_21033);
nor U22973 (N_22973,N_21001,N_21637);
nand U22974 (N_22974,N_20158,N_20328);
or U22975 (N_22975,N_21072,N_21801);
nand U22976 (N_22976,N_21891,N_21758);
nand U22977 (N_22977,N_21997,N_21186);
nand U22978 (N_22978,N_20187,N_21089);
xnor U22979 (N_22979,N_20493,N_20097);
nor U22980 (N_22980,N_21027,N_21841);
or U22981 (N_22981,N_21640,N_21510);
nand U22982 (N_22982,N_21561,N_21769);
and U22983 (N_22983,N_21444,N_21508);
or U22984 (N_22984,N_20852,N_21868);
or U22985 (N_22985,N_21931,N_20092);
nor U22986 (N_22986,N_20476,N_21205);
xnor U22987 (N_22987,N_20796,N_21446);
and U22988 (N_22988,N_20787,N_20686);
or U22989 (N_22989,N_21889,N_21807);
and U22990 (N_22990,N_21932,N_21091);
nand U22991 (N_22991,N_21936,N_21831);
or U22992 (N_22992,N_20220,N_21285);
nor U22993 (N_22993,N_20124,N_21681);
nor U22994 (N_22994,N_21447,N_20520);
nor U22995 (N_22995,N_20831,N_20715);
nand U22996 (N_22996,N_21772,N_21370);
nor U22997 (N_22997,N_20937,N_20956);
or U22998 (N_22998,N_20420,N_21760);
and U22999 (N_22999,N_20002,N_21631);
nor U23000 (N_23000,N_20492,N_21894);
nand U23001 (N_23001,N_20518,N_20867);
nand U23002 (N_23002,N_21527,N_20393);
nand U23003 (N_23003,N_21746,N_21255);
nand U23004 (N_23004,N_21125,N_21217);
nor U23005 (N_23005,N_21709,N_21152);
nand U23006 (N_23006,N_20097,N_21162);
and U23007 (N_23007,N_20148,N_20544);
nor U23008 (N_23008,N_20876,N_21791);
and U23009 (N_23009,N_20077,N_20570);
and U23010 (N_23010,N_21369,N_20109);
or U23011 (N_23011,N_21617,N_21655);
nor U23012 (N_23012,N_20679,N_21378);
nand U23013 (N_23013,N_20838,N_21334);
or U23014 (N_23014,N_20557,N_20182);
and U23015 (N_23015,N_21708,N_20564);
xnor U23016 (N_23016,N_20464,N_20636);
or U23017 (N_23017,N_20898,N_20383);
nand U23018 (N_23018,N_20615,N_20933);
or U23019 (N_23019,N_20974,N_21260);
or U23020 (N_23020,N_21369,N_20646);
nor U23021 (N_23021,N_20724,N_20234);
xnor U23022 (N_23022,N_21995,N_21231);
nand U23023 (N_23023,N_21133,N_20998);
nand U23024 (N_23024,N_20210,N_20717);
or U23025 (N_23025,N_20650,N_20835);
xnor U23026 (N_23026,N_21137,N_21574);
xor U23027 (N_23027,N_21604,N_21121);
and U23028 (N_23028,N_21356,N_21703);
nand U23029 (N_23029,N_21018,N_20622);
nand U23030 (N_23030,N_21020,N_20021);
xnor U23031 (N_23031,N_21783,N_20242);
or U23032 (N_23032,N_21740,N_21297);
or U23033 (N_23033,N_20421,N_21351);
nor U23034 (N_23034,N_21719,N_20039);
or U23035 (N_23035,N_21741,N_21031);
or U23036 (N_23036,N_20019,N_21175);
or U23037 (N_23037,N_21532,N_21733);
xnor U23038 (N_23038,N_20130,N_20362);
xnor U23039 (N_23039,N_20569,N_20089);
or U23040 (N_23040,N_20065,N_20880);
or U23041 (N_23041,N_20989,N_21124);
or U23042 (N_23042,N_20254,N_20294);
nand U23043 (N_23043,N_21596,N_21383);
nor U23044 (N_23044,N_21250,N_21816);
and U23045 (N_23045,N_20377,N_20192);
xor U23046 (N_23046,N_21651,N_21086);
xnor U23047 (N_23047,N_20114,N_20119);
and U23048 (N_23048,N_20027,N_20757);
nand U23049 (N_23049,N_20792,N_21684);
nor U23050 (N_23050,N_20724,N_20867);
and U23051 (N_23051,N_20496,N_20871);
or U23052 (N_23052,N_20157,N_21212);
nand U23053 (N_23053,N_20282,N_21395);
or U23054 (N_23054,N_21445,N_21032);
or U23055 (N_23055,N_21079,N_21475);
xor U23056 (N_23056,N_21838,N_21078);
nor U23057 (N_23057,N_20077,N_21129);
nand U23058 (N_23058,N_21470,N_21718);
nand U23059 (N_23059,N_21061,N_20609);
and U23060 (N_23060,N_20172,N_20191);
nor U23061 (N_23061,N_21034,N_20124);
nand U23062 (N_23062,N_20309,N_21937);
nand U23063 (N_23063,N_20314,N_21076);
xor U23064 (N_23064,N_20246,N_20175);
xor U23065 (N_23065,N_20542,N_20157);
nand U23066 (N_23066,N_21044,N_20515);
nor U23067 (N_23067,N_20322,N_20708);
and U23068 (N_23068,N_21108,N_20961);
or U23069 (N_23069,N_20617,N_20713);
xor U23070 (N_23070,N_21708,N_20853);
or U23071 (N_23071,N_21504,N_20746);
nand U23072 (N_23072,N_20253,N_20831);
or U23073 (N_23073,N_20413,N_21550);
nor U23074 (N_23074,N_21288,N_20656);
or U23075 (N_23075,N_21530,N_21469);
nand U23076 (N_23076,N_20951,N_20154);
or U23077 (N_23077,N_20374,N_20767);
nor U23078 (N_23078,N_21183,N_21053);
xor U23079 (N_23079,N_20282,N_20659);
nand U23080 (N_23080,N_21727,N_20657);
nor U23081 (N_23081,N_20568,N_20717);
nand U23082 (N_23082,N_20811,N_20469);
or U23083 (N_23083,N_21541,N_20585);
or U23084 (N_23084,N_20601,N_21011);
and U23085 (N_23085,N_20359,N_21558);
and U23086 (N_23086,N_20420,N_20243);
or U23087 (N_23087,N_20533,N_20188);
or U23088 (N_23088,N_21948,N_21425);
and U23089 (N_23089,N_21065,N_21214);
nand U23090 (N_23090,N_20848,N_20911);
xor U23091 (N_23091,N_20274,N_21665);
nand U23092 (N_23092,N_20192,N_20228);
and U23093 (N_23093,N_21809,N_20891);
xor U23094 (N_23094,N_21718,N_20664);
and U23095 (N_23095,N_20931,N_20451);
xnor U23096 (N_23096,N_20858,N_20573);
and U23097 (N_23097,N_20486,N_21874);
nor U23098 (N_23098,N_20224,N_21412);
and U23099 (N_23099,N_20675,N_20951);
and U23100 (N_23100,N_20575,N_21733);
and U23101 (N_23101,N_20742,N_21363);
or U23102 (N_23102,N_20516,N_21881);
nand U23103 (N_23103,N_21256,N_20323);
nor U23104 (N_23104,N_21464,N_21436);
xnor U23105 (N_23105,N_21624,N_20217);
nand U23106 (N_23106,N_21776,N_21754);
xor U23107 (N_23107,N_20997,N_21288);
or U23108 (N_23108,N_21695,N_20240);
nand U23109 (N_23109,N_21680,N_21574);
and U23110 (N_23110,N_21411,N_20191);
or U23111 (N_23111,N_20774,N_21414);
and U23112 (N_23112,N_21560,N_20815);
nor U23113 (N_23113,N_20557,N_20424);
nand U23114 (N_23114,N_21556,N_20837);
and U23115 (N_23115,N_21734,N_21771);
and U23116 (N_23116,N_21966,N_20375);
nand U23117 (N_23117,N_20340,N_21734);
nor U23118 (N_23118,N_20231,N_21402);
xor U23119 (N_23119,N_20474,N_21914);
or U23120 (N_23120,N_21842,N_20758);
and U23121 (N_23121,N_21051,N_20526);
nand U23122 (N_23122,N_21212,N_20936);
xnor U23123 (N_23123,N_21537,N_21067);
nor U23124 (N_23124,N_20184,N_21209);
nor U23125 (N_23125,N_20434,N_21321);
nand U23126 (N_23126,N_20956,N_20863);
xnor U23127 (N_23127,N_21001,N_21004);
and U23128 (N_23128,N_20921,N_20359);
nor U23129 (N_23129,N_21924,N_21818);
or U23130 (N_23130,N_21846,N_21333);
nor U23131 (N_23131,N_20118,N_21610);
nand U23132 (N_23132,N_20156,N_21602);
nor U23133 (N_23133,N_20250,N_21968);
or U23134 (N_23134,N_20905,N_20162);
or U23135 (N_23135,N_21053,N_21054);
and U23136 (N_23136,N_20345,N_21169);
and U23137 (N_23137,N_21779,N_20610);
nor U23138 (N_23138,N_21551,N_20849);
nand U23139 (N_23139,N_20850,N_20201);
xor U23140 (N_23140,N_21645,N_20084);
xor U23141 (N_23141,N_20103,N_21685);
and U23142 (N_23142,N_20004,N_20234);
or U23143 (N_23143,N_21587,N_21954);
nand U23144 (N_23144,N_20011,N_20192);
or U23145 (N_23145,N_21045,N_21396);
nor U23146 (N_23146,N_21784,N_21497);
or U23147 (N_23147,N_21460,N_20271);
nor U23148 (N_23148,N_20344,N_20678);
nand U23149 (N_23149,N_21521,N_20556);
or U23150 (N_23150,N_20649,N_21969);
or U23151 (N_23151,N_20611,N_20229);
nor U23152 (N_23152,N_20576,N_20440);
nand U23153 (N_23153,N_21897,N_21896);
xnor U23154 (N_23154,N_21463,N_20795);
nand U23155 (N_23155,N_21804,N_20670);
xnor U23156 (N_23156,N_20858,N_20323);
xor U23157 (N_23157,N_21108,N_20708);
or U23158 (N_23158,N_21906,N_21981);
or U23159 (N_23159,N_20291,N_21566);
nor U23160 (N_23160,N_20793,N_20601);
nand U23161 (N_23161,N_21443,N_21489);
xor U23162 (N_23162,N_21524,N_20794);
xor U23163 (N_23163,N_21692,N_20037);
nor U23164 (N_23164,N_20817,N_21322);
nor U23165 (N_23165,N_21734,N_20445);
nor U23166 (N_23166,N_20518,N_20324);
nand U23167 (N_23167,N_21986,N_21904);
nand U23168 (N_23168,N_21007,N_20151);
or U23169 (N_23169,N_20372,N_20502);
nand U23170 (N_23170,N_20348,N_20959);
and U23171 (N_23171,N_20124,N_20186);
nand U23172 (N_23172,N_20857,N_21978);
nor U23173 (N_23173,N_21009,N_20458);
and U23174 (N_23174,N_20370,N_20857);
and U23175 (N_23175,N_20880,N_20119);
or U23176 (N_23176,N_21604,N_20485);
or U23177 (N_23177,N_21859,N_20141);
nor U23178 (N_23178,N_21501,N_21869);
or U23179 (N_23179,N_21620,N_21684);
nand U23180 (N_23180,N_21088,N_20994);
xor U23181 (N_23181,N_21027,N_20813);
nand U23182 (N_23182,N_20929,N_20793);
xor U23183 (N_23183,N_20515,N_21911);
xnor U23184 (N_23184,N_20802,N_20123);
or U23185 (N_23185,N_21558,N_20794);
nor U23186 (N_23186,N_21492,N_21221);
and U23187 (N_23187,N_20071,N_20231);
nor U23188 (N_23188,N_21965,N_21267);
nand U23189 (N_23189,N_21358,N_20659);
nor U23190 (N_23190,N_21446,N_20564);
nand U23191 (N_23191,N_20854,N_20881);
or U23192 (N_23192,N_20708,N_20531);
or U23193 (N_23193,N_21448,N_21426);
or U23194 (N_23194,N_20555,N_21701);
or U23195 (N_23195,N_20408,N_21778);
xor U23196 (N_23196,N_20921,N_20767);
nor U23197 (N_23197,N_21085,N_21178);
xnor U23198 (N_23198,N_20785,N_20903);
nand U23199 (N_23199,N_21477,N_21210);
nor U23200 (N_23200,N_21238,N_21666);
or U23201 (N_23201,N_20900,N_21460);
and U23202 (N_23202,N_20796,N_20757);
xor U23203 (N_23203,N_20166,N_20405);
xor U23204 (N_23204,N_21462,N_20389);
nand U23205 (N_23205,N_21995,N_21525);
or U23206 (N_23206,N_21439,N_20394);
nor U23207 (N_23207,N_20539,N_21998);
nor U23208 (N_23208,N_20676,N_21478);
nor U23209 (N_23209,N_20601,N_20479);
and U23210 (N_23210,N_21188,N_21218);
xnor U23211 (N_23211,N_21060,N_21268);
nor U23212 (N_23212,N_21297,N_21028);
or U23213 (N_23213,N_20677,N_20912);
nand U23214 (N_23214,N_21354,N_21999);
and U23215 (N_23215,N_21188,N_21225);
nor U23216 (N_23216,N_20098,N_21813);
or U23217 (N_23217,N_21467,N_21205);
or U23218 (N_23218,N_20477,N_21739);
xor U23219 (N_23219,N_20163,N_21761);
nor U23220 (N_23220,N_21081,N_21409);
nand U23221 (N_23221,N_20670,N_21487);
nor U23222 (N_23222,N_20347,N_21362);
nand U23223 (N_23223,N_21802,N_20403);
nand U23224 (N_23224,N_21510,N_21986);
xor U23225 (N_23225,N_20655,N_21718);
nand U23226 (N_23226,N_20489,N_20524);
nand U23227 (N_23227,N_20155,N_21524);
xnor U23228 (N_23228,N_20389,N_21999);
or U23229 (N_23229,N_21321,N_20553);
or U23230 (N_23230,N_21493,N_20397);
nand U23231 (N_23231,N_21438,N_21964);
nand U23232 (N_23232,N_20630,N_20566);
or U23233 (N_23233,N_20170,N_21498);
xor U23234 (N_23234,N_20907,N_20885);
and U23235 (N_23235,N_20387,N_21859);
xor U23236 (N_23236,N_21913,N_20223);
nand U23237 (N_23237,N_20663,N_21265);
and U23238 (N_23238,N_21357,N_21485);
and U23239 (N_23239,N_21152,N_20948);
nor U23240 (N_23240,N_21216,N_21077);
and U23241 (N_23241,N_20627,N_21302);
nand U23242 (N_23242,N_20119,N_21977);
or U23243 (N_23243,N_21235,N_21498);
or U23244 (N_23244,N_21041,N_21384);
xor U23245 (N_23245,N_21915,N_21550);
and U23246 (N_23246,N_21074,N_21787);
nand U23247 (N_23247,N_20171,N_21018);
or U23248 (N_23248,N_21277,N_20235);
nand U23249 (N_23249,N_20067,N_20042);
or U23250 (N_23250,N_20697,N_20299);
xor U23251 (N_23251,N_20014,N_21563);
nor U23252 (N_23252,N_20205,N_21523);
xor U23253 (N_23253,N_20926,N_21947);
nand U23254 (N_23254,N_20617,N_20755);
nand U23255 (N_23255,N_20786,N_20891);
xor U23256 (N_23256,N_20514,N_21776);
nor U23257 (N_23257,N_21460,N_20179);
nand U23258 (N_23258,N_20886,N_21752);
or U23259 (N_23259,N_21239,N_21217);
and U23260 (N_23260,N_21436,N_20560);
xnor U23261 (N_23261,N_21996,N_21176);
xor U23262 (N_23262,N_20068,N_20578);
or U23263 (N_23263,N_20976,N_20760);
nand U23264 (N_23264,N_21203,N_20571);
nand U23265 (N_23265,N_20567,N_20688);
nand U23266 (N_23266,N_21466,N_21755);
nor U23267 (N_23267,N_21630,N_21323);
xnor U23268 (N_23268,N_20182,N_20827);
nand U23269 (N_23269,N_20040,N_21434);
and U23270 (N_23270,N_20077,N_21371);
nor U23271 (N_23271,N_21012,N_21270);
nor U23272 (N_23272,N_20265,N_20244);
xor U23273 (N_23273,N_21729,N_20332);
nand U23274 (N_23274,N_20522,N_21547);
or U23275 (N_23275,N_21968,N_20809);
or U23276 (N_23276,N_21502,N_21699);
nor U23277 (N_23277,N_20741,N_21741);
nor U23278 (N_23278,N_21097,N_21123);
nand U23279 (N_23279,N_20974,N_20480);
nor U23280 (N_23280,N_20690,N_20821);
nand U23281 (N_23281,N_20989,N_21802);
or U23282 (N_23282,N_20254,N_20653);
xnor U23283 (N_23283,N_20326,N_20880);
nor U23284 (N_23284,N_21057,N_21903);
nor U23285 (N_23285,N_20635,N_21008);
xnor U23286 (N_23286,N_21479,N_20723);
and U23287 (N_23287,N_21775,N_21454);
or U23288 (N_23288,N_20385,N_21577);
or U23289 (N_23289,N_21035,N_20524);
and U23290 (N_23290,N_20327,N_20195);
nand U23291 (N_23291,N_21719,N_21192);
and U23292 (N_23292,N_20468,N_20352);
or U23293 (N_23293,N_20194,N_20843);
nor U23294 (N_23294,N_21230,N_20242);
xnor U23295 (N_23295,N_20462,N_21751);
or U23296 (N_23296,N_21288,N_21677);
or U23297 (N_23297,N_21773,N_20208);
or U23298 (N_23298,N_21782,N_21078);
or U23299 (N_23299,N_21774,N_20337);
xor U23300 (N_23300,N_20649,N_20406);
and U23301 (N_23301,N_21705,N_21773);
or U23302 (N_23302,N_20591,N_21896);
or U23303 (N_23303,N_21815,N_21043);
and U23304 (N_23304,N_20308,N_20114);
nor U23305 (N_23305,N_20473,N_20679);
or U23306 (N_23306,N_21576,N_20834);
nand U23307 (N_23307,N_21555,N_21141);
xnor U23308 (N_23308,N_20934,N_21794);
xor U23309 (N_23309,N_21114,N_20439);
nand U23310 (N_23310,N_21903,N_21193);
nand U23311 (N_23311,N_21500,N_20169);
nor U23312 (N_23312,N_21703,N_21046);
nor U23313 (N_23313,N_20950,N_21396);
nand U23314 (N_23314,N_21278,N_20039);
or U23315 (N_23315,N_21149,N_20272);
or U23316 (N_23316,N_20727,N_21790);
nand U23317 (N_23317,N_20504,N_20560);
or U23318 (N_23318,N_21756,N_21150);
and U23319 (N_23319,N_20000,N_20935);
or U23320 (N_23320,N_20654,N_20447);
nor U23321 (N_23321,N_21268,N_20606);
and U23322 (N_23322,N_20503,N_21558);
or U23323 (N_23323,N_21120,N_21994);
xnor U23324 (N_23324,N_21514,N_21810);
xnor U23325 (N_23325,N_20652,N_20767);
or U23326 (N_23326,N_20730,N_21596);
and U23327 (N_23327,N_21928,N_20225);
nor U23328 (N_23328,N_21197,N_20903);
nor U23329 (N_23329,N_20661,N_20514);
nor U23330 (N_23330,N_20203,N_20504);
xnor U23331 (N_23331,N_20556,N_21553);
nand U23332 (N_23332,N_20684,N_21008);
or U23333 (N_23333,N_21421,N_21505);
xor U23334 (N_23334,N_21667,N_20014);
nand U23335 (N_23335,N_21426,N_21207);
nor U23336 (N_23336,N_21972,N_21820);
or U23337 (N_23337,N_21802,N_21510);
nand U23338 (N_23338,N_21832,N_21550);
nand U23339 (N_23339,N_21456,N_21751);
xnor U23340 (N_23340,N_21233,N_21908);
and U23341 (N_23341,N_21016,N_20766);
or U23342 (N_23342,N_21343,N_21615);
xnor U23343 (N_23343,N_20250,N_21250);
nor U23344 (N_23344,N_20215,N_20324);
or U23345 (N_23345,N_20485,N_20942);
nor U23346 (N_23346,N_20617,N_21972);
and U23347 (N_23347,N_21974,N_21903);
nand U23348 (N_23348,N_20571,N_20858);
xnor U23349 (N_23349,N_21026,N_21360);
and U23350 (N_23350,N_20497,N_21699);
or U23351 (N_23351,N_21421,N_20074);
or U23352 (N_23352,N_21866,N_20988);
nor U23353 (N_23353,N_21430,N_21601);
xor U23354 (N_23354,N_21479,N_21626);
and U23355 (N_23355,N_20707,N_21277);
or U23356 (N_23356,N_20685,N_20745);
xnor U23357 (N_23357,N_20862,N_21220);
and U23358 (N_23358,N_21986,N_20636);
nand U23359 (N_23359,N_20411,N_20053);
xnor U23360 (N_23360,N_21913,N_20467);
and U23361 (N_23361,N_21471,N_21343);
xor U23362 (N_23362,N_20269,N_20311);
nand U23363 (N_23363,N_20990,N_21785);
nor U23364 (N_23364,N_21781,N_21313);
nor U23365 (N_23365,N_21120,N_20080);
or U23366 (N_23366,N_20267,N_20097);
and U23367 (N_23367,N_20810,N_20761);
and U23368 (N_23368,N_21811,N_21253);
and U23369 (N_23369,N_21644,N_20924);
xnor U23370 (N_23370,N_20886,N_20182);
nor U23371 (N_23371,N_21687,N_21754);
nand U23372 (N_23372,N_21991,N_20327);
xor U23373 (N_23373,N_20534,N_21053);
xnor U23374 (N_23374,N_21233,N_20952);
and U23375 (N_23375,N_20323,N_20820);
nand U23376 (N_23376,N_21368,N_20049);
nand U23377 (N_23377,N_20893,N_21897);
nor U23378 (N_23378,N_20317,N_21769);
or U23379 (N_23379,N_21823,N_21511);
nand U23380 (N_23380,N_20069,N_20808);
nor U23381 (N_23381,N_20391,N_20638);
nand U23382 (N_23382,N_20435,N_21628);
xnor U23383 (N_23383,N_20846,N_20360);
and U23384 (N_23384,N_20810,N_21412);
nand U23385 (N_23385,N_20961,N_21098);
nand U23386 (N_23386,N_21415,N_21117);
nor U23387 (N_23387,N_21914,N_21255);
xor U23388 (N_23388,N_20713,N_21336);
nor U23389 (N_23389,N_21185,N_21377);
xnor U23390 (N_23390,N_21598,N_20121);
or U23391 (N_23391,N_21719,N_20389);
nand U23392 (N_23392,N_20828,N_20774);
or U23393 (N_23393,N_20765,N_21443);
and U23394 (N_23394,N_21144,N_20761);
xnor U23395 (N_23395,N_21459,N_21711);
xor U23396 (N_23396,N_21750,N_21176);
and U23397 (N_23397,N_20539,N_21588);
nor U23398 (N_23398,N_21959,N_20620);
and U23399 (N_23399,N_20511,N_20604);
nand U23400 (N_23400,N_20853,N_20669);
or U23401 (N_23401,N_21245,N_20535);
nor U23402 (N_23402,N_21441,N_20739);
nand U23403 (N_23403,N_20278,N_21620);
and U23404 (N_23404,N_21397,N_21904);
and U23405 (N_23405,N_20050,N_20819);
or U23406 (N_23406,N_21802,N_21039);
xnor U23407 (N_23407,N_20442,N_20115);
nor U23408 (N_23408,N_20605,N_21922);
nor U23409 (N_23409,N_21715,N_21013);
and U23410 (N_23410,N_20525,N_20442);
xor U23411 (N_23411,N_20865,N_21516);
and U23412 (N_23412,N_20163,N_21677);
nor U23413 (N_23413,N_21971,N_21670);
nand U23414 (N_23414,N_20852,N_21606);
nor U23415 (N_23415,N_21844,N_20844);
nand U23416 (N_23416,N_20975,N_21458);
xnor U23417 (N_23417,N_20340,N_21637);
nand U23418 (N_23418,N_20503,N_20662);
nand U23419 (N_23419,N_21132,N_21444);
nor U23420 (N_23420,N_21922,N_21419);
and U23421 (N_23421,N_20574,N_21473);
xnor U23422 (N_23422,N_20490,N_20457);
xor U23423 (N_23423,N_21596,N_21791);
nor U23424 (N_23424,N_21936,N_21917);
nor U23425 (N_23425,N_20701,N_21028);
xor U23426 (N_23426,N_20884,N_21397);
nor U23427 (N_23427,N_20509,N_21688);
nor U23428 (N_23428,N_21191,N_21350);
and U23429 (N_23429,N_20221,N_21483);
and U23430 (N_23430,N_20682,N_21677);
nor U23431 (N_23431,N_20336,N_20162);
nor U23432 (N_23432,N_20907,N_21544);
or U23433 (N_23433,N_20240,N_20719);
xnor U23434 (N_23434,N_21081,N_21534);
and U23435 (N_23435,N_20773,N_21358);
xor U23436 (N_23436,N_20259,N_21210);
nor U23437 (N_23437,N_21507,N_20276);
and U23438 (N_23438,N_20410,N_21126);
xor U23439 (N_23439,N_21978,N_21138);
xor U23440 (N_23440,N_21437,N_20311);
xor U23441 (N_23441,N_20914,N_20587);
xnor U23442 (N_23442,N_20298,N_20153);
xor U23443 (N_23443,N_20645,N_21699);
and U23444 (N_23444,N_20533,N_20789);
nor U23445 (N_23445,N_20537,N_21891);
nand U23446 (N_23446,N_21764,N_21698);
nor U23447 (N_23447,N_21798,N_21815);
nor U23448 (N_23448,N_21623,N_21821);
nand U23449 (N_23449,N_21114,N_20467);
and U23450 (N_23450,N_20575,N_20425);
xor U23451 (N_23451,N_21187,N_20745);
or U23452 (N_23452,N_20169,N_20030);
or U23453 (N_23453,N_21516,N_21527);
nand U23454 (N_23454,N_21204,N_21526);
or U23455 (N_23455,N_21000,N_21318);
and U23456 (N_23456,N_21468,N_21324);
nand U23457 (N_23457,N_20380,N_20689);
nor U23458 (N_23458,N_21129,N_20679);
and U23459 (N_23459,N_21456,N_21341);
xor U23460 (N_23460,N_20916,N_21961);
nand U23461 (N_23461,N_20391,N_21003);
or U23462 (N_23462,N_20651,N_20074);
or U23463 (N_23463,N_21649,N_20299);
or U23464 (N_23464,N_21903,N_20449);
xor U23465 (N_23465,N_21201,N_21047);
and U23466 (N_23466,N_20790,N_21362);
and U23467 (N_23467,N_20579,N_21122);
nor U23468 (N_23468,N_21009,N_20775);
or U23469 (N_23469,N_21029,N_20368);
and U23470 (N_23470,N_21396,N_21119);
and U23471 (N_23471,N_21122,N_21632);
xnor U23472 (N_23472,N_20235,N_20152);
nor U23473 (N_23473,N_21975,N_20836);
nor U23474 (N_23474,N_20218,N_20940);
nand U23475 (N_23475,N_21377,N_20161);
or U23476 (N_23476,N_21726,N_20307);
xnor U23477 (N_23477,N_21418,N_21369);
or U23478 (N_23478,N_21670,N_21236);
nor U23479 (N_23479,N_20899,N_21928);
xnor U23480 (N_23480,N_21934,N_21194);
and U23481 (N_23481,N_20619,N_21014);
nor U23482 (N_23482,N_21843,N_20257);
nor U23483 (N_23483,N_21176,N_20224);
nor U23484 (N_23484,N_21506,N_20244);
xor U23485 (N_23485,N_20786,N_21871);
and U23486 (N_23486,N_21207,N_20468);
xnor U23487 (N_23487,N_21063,N_20322);
and U23488 (N_23488,N_20241,N_21446);
nand U23489 (N_23489,N_20217,N_20647);
and U23490 (N_23490,N_20664,N_21789);
xor U23491 (N_23491,N_21820,N_21507);
and U23492 (N_23492,N_21657,N_20180);
or U23493 (N_23493,N_20664,N_21234);
and U23494 (N_23494,N_21343,N_20778);
nor U23495 (N_23495,N_20533,N_20365);
and U23496 (N_23496,N_21777,N_20776);
xnor U23497 (N_23497,N_20398,N_20189);
and U23498 (N_23498,N_20007,N_20364);
nand U23499 (N_23499,N_20640,N_20537);
or U23500 (N_23500,N_20968,N_20598);
xor U23501 (N_23501,N_20566,N_20944);
or U23502 (N_23502,N_20067,N_20361);
xor U23503 (N_23503,N_21606,N_20563);
nor U23504 (N_23504,N_20995,N_20722);
or U23505 (N_23505,N_21920,N_20469);
or U23506 (N_23506,N_21777,N_20861);
nor U23507 (N_23507,N_20112,N_20656);
nor U23508 (N_23508,N_20319,N_21229);
or U23509 (N_23509,N_21683,N_21674);
or U23510 (N_23510,N_21363,N_20814);
nor U23511 (N_23511,N_20437,N_20560);
and U23512 (N_23512,N_20628,N_20713);
nand U23513 (N_23513,N_20903,N_20110);
xor U23514 (N_23514,N_21583,N_20111);
or U23515 (N_23515,N_20627,N_21793);
or U23516 (N_23516,N_20785,N_20886);
and U23517 (N_23517,N_21139,N_21438);
nor U23518 (N_23518,N_21356,N_20357);
and U23519 (N_23519,N_21572,N_20628);
or U23520 (N_23520,N_20589,N_20513);
nand U23521 (N_23521,N_21498,N_21786);
and U23522 (N_23522,N_20573,N_21194);
nand U23523 (N_23523,N_20453,N_21191);
nor U23524 (N_23524,N_21673,N_20122);
nand U23525 (N_23525,N_20004,N_21141);
xnor U23526 (N_23526,N_21718,N_20841);
or U23527 (N_23527,N_21660,N_21095);
and U23528 (N_23528,N_21598,N_20010);
xor U23529 (N_23529,N_21185,N_20379);
nor U23530 (N_23530,N_20433,N_20440);
nor U23531 (N_23531,N_20791,N_21818);
nor U23532 (N_23532,N_21361,N_21537);
nor U23533 (N_23533,N_20060,N_21689);
nand U23534 (N_23534,N_20595,N_21300);
nand U23535 (N_23535,N_21339,N_21563);
or U23536 (N_23536,N_20505,N_20843);
or U23537 (N_23537,N_21464,N_21201);
nor U23538 (N_23538,N_21747,N_21969);
nor U23539 (N_23539,N_20930,N_20763);
xnor U23540 (N_23540,N_21214,N_20816);
and U23541 (N_23541,N_20329,N_21209);
nand U23542 (N_23542,N_20254,N_21420);
and U23543 (N_23543,N_20292,N_21758);
nor U23544 (N_23544,N_20303,N_20506);
xnor U23545 (N_23545,N_21104,N_21575);
nor U23546 (N_23546,N_20977,N_20544);
and U23547 (N_23547,N_20462,N_20614);
xor U23548 (N_23548,N_21917,N_21343);
xnor U23549 (N_23549,N_20069,N_21522);
or U23550 (N_23550,N_21480,N_20996);
nor U23551 (N_23551,N_21228,N_20366);
nand U23552 (N_23552,N_20829,N_20169);
nand U23553 (N_23553,N_21094,N_20584);
and U23554 (N_23554,N_21227,N_20552);
xnor U23555 (N_23555,N_21275,N_21817);
and U23556 (N_23556,N_21040,N_20200);
nand U23557 (N_23557,N_20147,N_20802);
or U23558 (N_23558,N_21484,N_21182);
nand U23559 (N_23559,N_21427,N_21570);
and U23560 (N_23560,N_20094,N_21562);
xor U23561 (N_23561,N_20657,N_21784);
nor U23562 (N_23562,N_21341,N_20373);
nand U23563 (N_23563,N_20944,N_20862);
xor U23564 (N_23564,N_20921,N_20897);
nor U23565 (N_23565,N_20142,N_20060);
xnor U23566 (N_23566,N_20154,N_20293);
nand U23567 (N_23567,N_20531,N_21988);
nor U23568 (N_23568,N_21581,N_20276);
and U23569 (N_23569,N_20352,N_20060);
xor U23570 (N_23570,N_21568,N_21052);
nor U23571 (N_23571,N_21726,N_21775);
xnor U23572 (N_23572,N_20660,N_21796);
and U23573 (N_23573,N_20394,N_21441);
and U23574 (N_23574,N_21402,N_20541);
nand U23575 (N_23575,N_21102,N_20004);
or U23576 (N_23576,N_21820,N_20623);
and U23577 (N_23577,N_20318,N_20142);
xor U23578 (N_23578,N_20212,N_21235);
nand U23579 (N_23579,N_20505,N_20415);
nand U23580 (N_23580,N_20535,N_21569);
nor U23581 (N_23581,N_20961,N_20943);
nand U23582 (N_23582,N_21554,N_20083);
nor U23583 (N_23583,N_20071,N_21778);
or U23584 (N_23584,N_21528,N_20363);
nand U23585 (N_23585,N_20142,N_20660);
or U23586 (N_23586,N_20254,N_20365);
or U23587 (N_23587,N_20365,N_20484);
or U23588 (N_23588,N_20062,N_21718);
nand U23589 (N_23589,N_21348,N_20161);
and U23590 (N_23590,N_21426,N_21368);
xor U23591 (N_23591,N_21967,N_21202);
or U23592 (N_23592,N_21698,N_20299);
nor U23593 (N_23593,N_20884,N_20997);
nand U23594 (N_23594,N_21011,N_20701);
and U23595 (N_23595,N_20874,N_20166);
xnor U23596 (N_23596,N_21604,N_20095);
and U23597 (N_23597,N_21808,N_20729);
and U23598 (N_23598,N_20589,N_21049);
and U23599 (N_23599,N_21077,N_20512);
nand U23600 (N_23600,N_21494,N_21208);
xor U23601 (N_23601,N_20006,N_21452);
and U23602 (N_23602,N_21261,N_21553);
nand U23603 (N_23603,N_20357,N_20939);
nand U23604 (N_23604,N_20373,N_21668);
and U23605 (N_23605,N_20403,N_20734);
and U23606 (N_23606,N_20515,N_20891);
xnor U23607 (N_23607,N_20327,N_20563);
nor U23608 (N_23608,N_21607,N_21042);
and U23609 (N_23609,N_21193,N_21291);
nor U23610 (N_23610,N_20964,N_20838);
and U23611 (N_23611,N_21922,N_21861);
nor U23612 (N_23612,N_21140,N_20569);
and U23613 (N_23613,N_20540,N_20516);
xor U23614 (N_23614,N_20579,N_21691);
and U23615 (N_23615,N_20662,N_20742);
nor U23616 (N_23616,N_20966,N_20562);
xor U23617 (N_23617,N_20398,N_20205);
and U23618 (N_23618,N_20723,N_20287);
nor U23619 (N_23619,N_21802,N_20652);
and U23620 (N_23620,N_20211,N_20852);
and U23621 (N_23621,N_20809,N_21732);
and U23622 (N_23622,N_21029,N_20121);
nor U23623 (N_23623,N_20055,N_21420);
nand U23624 (N_23624,N_20623,N_21203);
nand U23625 (N_23625,N_21536,N_20033);
nor U23626 (N_23626,N_21787,N_20302);
nand U23627 (N_23627,N_20520,N_21897);
nand U23628 (N_23628,N_21218,N_21897);
nor U23629 (N_23629,N_21446,N_21226);
and U23630 (N_23630,N_20184,N_21766);
nand U23631 (N_23631,N_20693,N_20103);
nand U23632 (N_23632,N_21544,N_21755);
nor U23633 (N_23633,N_20752,N_20999);
and U23634 (N_23634,N_21224,N_20734);
xor U23635 (N_23635,N_21911,N_21797);
and U23636 (N_23636,N_20972,N_21765);
and U23637 (N_23637,N_20775,N_20640);
and U23638 (N_23638,N_20414,N_21561);
and U23639 (N_23639,N_21498,N_21507);
xor U23640 (N_23640,N_21364,N_20243);
nor U23641 (N_23641,N_20829,N_20168);
nor U23642 (N_23642,N_21731,N_20348);
nand U23643 (N_23643,N_21998,N_21812);
and U23644 (N_23644,N_20675,N_20047);
nand U23645 (N_23645,N_20145,N_20967);
nand U23646 (N_23646,N_21982,N_20342);
or U23647 (N_23647,N_21804,N_20641);
nor U23648 (N_23648,N_21045,N_20517);
xor U23649 (N_23649,N_20459,N_20754);
nor U23650 (N_23650,N_20148,N_21514);
nand U23651 (N_23651,N_20546,N_21425);
xor U23652 (N_23652,N_20162,N_20748);
or U23653 (N_23653,N_20426,N_21438);
nand U23654 (N_23654,N_20498,N_20409);
xnor U23655 (N_23655,N_20621,N_21973);
xor U23656 (N_23656,N_21157,N_20116);
nor U23657 (N_23657,N_20693,N_21443);
nor U23658 (N_23658,N_21046,N_20849);
nor U23659 (N_23659,N_20760,N_21324);
or U23660 (N_23660,N_20968,N_20319);
or U23661 (N_23661,N_21329,N_21676);
nor U23662 (N_23662,N_20723,N_20629);
nand U23663 (N_23663,N_20910,N_20205);
nand U23664 (N_23664,N_20223,N_21679);
nor U23665 (N_23665,N_20676,N_20486);
nor U23666 (N_23666,N_20172,N_21382);
and U23667 (N_23667,N_20699,N_20426);
xnor U23668 (N_23668,N_20317,N_21309);
nand U23669 (N_23669,N_21165,N_20883);
xnor U23670 (N_23670,N_20410,N_21786);
or U23671 (N_23671,N_21352,N_21388);
xnor U23672 (N_23672,N_21126,N_20720);
nor U23673 (N_23673,N_20494,N_20002);
xor U23674 (N_23674,N_21306,N_20582);
and U23675 (N_23675,N_21598,N_21068);
and U23676 (N_23676,N_20575,N_20324);
nand U23677 (N_23677,N_20578,N_20664);
nand U23678 (N_23678,N_20320,N_21748);
nand U23679 (N_23679,N_21497,N_21805);
xnor U23680 (N_23680,N_20214,N_20799);
nor U23681 (N_23681,N_20065,N_21157);
nor U23682 (N_23682,N_20572,N_20561);
or U23683 (N_23683,N_20052,N_21548);
xnor U23684 (N_23684,N_21001,N_20196);
xor U23685 (N_23685,N_21865,N_20106);
xor U23686 (N_23686,N_21152,N_20016);
nand U23687 (N_23687,N_20396,N_20502);
and U23688 (N_23688,N_20392,N_21266);
nand U23689 (N_23689,N_20189,N_21022);
or U23690 (N_23690,N_20358,N_20095);
nand U23691 (N_23691,N_20881,N_21968);
nor U23692 (N_23692,N_21096,N_21353);
and U23693 (N_23693,N_21767,N_21655);
or U23694 (N_23694,N_21381,N_20493);
nor U23695 (N_23695,N_20459,N_21865);
and U23696 (N_23696,N_21755,N_21037);
xor U23697 (N_23697,N_21649,N_21874);
nand U23698 (N_23698,N_20612,N_21976);
xnor U23699 (N_23699,N_21654,N_20790);
nor U23700 (N_23700,N_21548,N_21205);
or U23701 (N_23701,N_21155,N_20971);
nor U23702 (N_23702,N_20399,N_20426);
xnor U23703 (N_23703,N_21938,N_20139);
nand U23704 (N_23704,N_20225,N_21245);
and U23705 (N_23705,N_21801,N_20582);
and U23706 (N_23706,N_20755,N_20689);
nor U23707 (N_23707,N_20922,N_20759);
xor U23708 (N_23708,N_21104,N_21904);
and U23709 (N_23709,N_20165,N_20078);
and U23710 (N_23710,N_20734,N_21280);
nor U23711 (N_23711,N_21606,N_21383);
nand U23712 (N_23712,N_20911,N_21581);
nand U23713 (N_23713,N_21983,N_20131);
nor U23714 (N_23714,N_20207,N_21428);
and U23715 (N_23715,N_21928,N_21622);
xnor U23716 (N_23716,N_20991,N_21751);
nand U23717 (N_23717,N_21881,N_20159);
nor U23718 (N_23718,N_21810,N_21239);
and U23719 (N_23719,N_20245,N_21475);
xor U23720 (N_23720,N_21646,N_21420);
or U23721 (N_23721,N_21571,N_21555);
nand U23722 (N_23722,N_20019,N_20884);
xnor U23723 (N_23723,N_20537,N_20873);
or U23724 (N_23724,N_20051,N_21726);
or U23725 (N_23725,N_21949,N_21528);
xor U23726 (N_23726,N_21544,N_21510);
nor U23727 (N_23727,N_20613,N_21195);
nor U23728 (N_23728,N_20341,N_21709);
xor U23729 (N_23729,N_21338,N_20990);
nor U23730 (N_23730,N_20986,N_20369);
xnor U23731 (N_23731,N_20562,N_20696);
nand U23732 (N_23732,N_21688,N_20236);
and U23733 (N_23733,N_21012,N_20219);
nand U23734 (N_23734,N_21350,N_20686);
nor U23735 (N_23735,N_21321,N_20230);
and U23736 (N_23736,N_21587,N_20571);
and U23737 (N_23737,N_20969,N_20473);
nor U23738 (N_23738,N_21609,N_20579);
xnor U23739 (N_23739,N_20688,N_20052);
nand U23740 (N_23740,N_20891,N_21936);
or U23741 (N_23741,N_21793,N_21124);
and U23742 (N_23742,N_20283,N_20205);
and U23743 (N_23743,N_20149,N_20707);
or U23744 (N_23744,N_20944,N_20214);
or U23745 (N_23745,N_20209,N_21973);
and U23746 (N_23746,N_21958,N_20417);
nor U23747 (N_23747,N_20661,N_20162);
and U23748 (N_23748,N_21954,N_20405);
and U23749 (N_23749,N_20178,N_20124);
nor U23750 (N_23750,N_21967,N_20414);
and U23751 (N_23751,N_21474,N_21930);
xor U23752 (N_23752,N_21418,N_21987);
nand U23753 (N_23753,N_20352,N_20691);
or U23754 (N_23754,N_21850,N_20610);
nor U23755 (N_23755,N_20421,N_21064);
or U23756 (N_23756,N_20970,N_21383);
xor U23757 (N_23757,N_20030,N_20443);
or U23758 (N_23758,N_20156,N_20290);
xnor U23759 (N_23759,N_21310,N_20386);
and U23760 (N_23760,N_21086,N_20291);
or U23761 (N_23761,N_20271,N_21114);
xnor U23762 (N_23762,N_20608,N_20153);
nand U23763 (N_23763,N_20301,N_20039);
xor U23764 (N_23764,N_21389,N_21603);
or U23765 (N_23765,N_21299,N_20671);
nand U23766 (N_23766,N_20648,N_21188);
nand U23767 (N_23767,N_20519,N_21109);
nand U23768 (N_23768,N_20787,N_20583);
and U23769 (N_23769,N_20796,N_21821);
or U23770 (N_23770,N_21117,N_20440);
and U23771 (N_23771,N_20916,N_21759);
or U23772 (N_23772,N_21569,N_20985);
nor U23773 (N_23773,N_21609,N_20302);
or U23774 (N_23774,N_20788,N_20981);
nand U23775 (N_23775,N_20196,N_21503);
or U23776 (N_23776,N_20034,N_21022);
nand U23777 (N_23777,N_20601,N_21836);
or U23778 (N_23778,N_20529,N_20655);
nor U23779 (N_23779,N_21433,N_21648);
xnor U23780 (N_23780,N_21585,N_21914);
or U23781 (N_23781,N_21507,N_21037);
nor U23782 (N_23782,N_21643,N_20567);
and U23783 (N_23783,N_20581,N_21434);
nor U23784 (N_23784,N_21368,N_21581);
or U23785 (N_23785,N_20135,N_21916);
nor U23786 (N_23786,N_21587,N_21502);
and U23787 (N_23787,N_21581,N_21331);
nor U23788 (N_23788,N_21385,N_21132);
nor U23789 (N_23789,N_21137,N_21400);
nor U23790 (N_23790,N_20117,N_20789);
xor U23791 (N_23791,N_20220,N_21086);
nor U23792 (N_23792,N_20124,N_21981);
xor U23793 (N_23793,N_21079,N_20640);
nor U23794 (N_23794,N_21357,N_21413);
xnor U23795 (N_23795,N_21738,N_21265);
xor U23796 (N_23796,N_21325,N_21309);
nor U23797 (N_23797,N_20963,N_21916);
and U23798 (N_23798,N_20330,N_20271);
nor U23799 (N_23799,N_20386,N_21189);
nor U23800 (N_23800,N_20031,N_21524);
or U23801 (N_23801,N_21454,N_21175);
nand U23802 (N_23802,N_20845,N_20401);
xnor U23803 (N_23803,N_20147,N_21450);
or U23804 (N_23804,N_21774,N_20360);
or U23805 (N_23805,N_20672,N_20099);
and U23806 (N_23806,N_21895,N_20124);
or U23807 (N_23807,N_21098,N_21943);
or U23808 (N_23808,N_20329,N_21690);
nor U23809 (N_23809,N_20394,N_21743);
nand U23810 (N_23810,N_21669,N_20723);
nor U23811 (N_23811,N_20828,N_20021);
xnor U23812 (N_23812,N_21685,N_20195);
nor U23813 (N_23813,N_21912,N_21863);
nor U23814 (N_23814,N_21928,N_20117);
xor U23815 (N_23815,N_20853,N_20415);
nand U23816 (N_23816,N_21417,N_20865);
xnor U23817 (N_23817,N_20498,N_20741);
or U23818 (N_23818,N_21727,N_20798);
or U23819 (N_23819,N_20258,N_20696);
or U23820 (N_23820,N_21148,N_21009);
nand U23821 (N_23821,N_20966,N_21932);
and U23822 (N_23822,N_20197,N_21025);
and U23823 (N_23823,N_21192,N_21563);
nand U23824 (N_23824,N_21649,N_20609);
or U23825 (N_23825,N_21801,N_21359);
nand U23826 (N_23826,N_21426,N_20237);
or U23827 (N_23827,N_20750,N_21837);
or U23828 (N_23828,N_21052,N_21233);
xor U23829 (N_23829,N_21202,N_20185);
nor U23830 (N_23830,N_20248,N_20272);
nor U23831 (N_23831,N_21284,N_20104);
or U23832 (N_23832,N_20445,N_21173);
nand U23833 (N_23833,N_21689,N_20424);
or U23834 (N_23834,N_21927,N_20121);
or U23835 (N_23835,N_21477,N_21155);
and U23836 (N_23836,N_21280,N_20955);
nor U23837 (N_23837,N_21793,N_21059);
xnor U23838 (N_23838,N_20089,N_21227);
xnor U23839 (N_23839,N_20703,N_21617);
or U23840 (N_23840,N_20693,N_21401);
or U23841 (N_23841,N_20481,N_20496);
xor U23842 (N_23842,N_21332,N_21402);
and U23843 (N_23843,N_21749,N_20921);
nand U23844 (N_23844,N_20358,N_21283);
nand U23845 (N_23845,N_21500,N_21632);
nand U23846 (N_23846,N_21060,N_20286);
and U23847 (N_23847,N_20512,N_20783);
or U23848 (N_23848,N_21629,N_20192);
xnor U23849 (N_23849,N_20644,N_21016);
xor U23850 (N_23850,N_20322,N_21056);
and U23851 (N_23851,N_21970,N_20981);
nor U23852 (N_23852,N_21379,N_21017);
nand U23853 (N_23853,N_20091,N_20692);
xor U23854 (N_23854,N_20115,N_21341);
and U23855 (N_23855,N_20428,N_20432);
or U23856 (N_23856,N_21167,N_21641);
nor U23857 (N_23857,N_20398,N_20523);
nand U23858 (N_23858,N_20415,N_21605);
nor U23859 (N_23859,N_21999,N_21583);
nand U23860 (N_23860,N_20916,N_20146);
xor U23861 (N_23861,N_20414,N_21884);
nor U23862 (N_23862,N_20955,N_20808);
nor U23863 (N_23863,N_21106,N_21175);
nor U23864 (N_23864,N_20309,N_21309);
xnor U23865 (N_23865,N_20196,N_21664);
or U23866 (N_23866,N_21012,N_20034);
xnor U23867 (N_23867,N_21768,N_20560);
or U23868 (N_23868,N_20649,N_20615);
nand U23869 (N_23869,N_21274,N_21020);
nor U23870 (N_23870,N_20430,N_21623);
and U23871 (N_23871,N_21631,N_21195);
xnor U23872 (N_23872,N_20972,N_21926);
and U23873 (N_23873,N_21153,N_20596);
xor U23874 (N_23874,N_21622,N_21961);
or U23875 (N_23875,N_21863,N_21034);
xor U23876 (N_23876,N_20595,N_20537);
and U23877 (N_23877,N_21101,N_21794);
and U23878 (N_23878,N_20033,N_20222);
nand U23879 (N_23879,N_21376,N_21458);
nand U23880 (N_23880,N_21506,N_21064);
xnor U23881 (N_23881,N_20026,N_20163);
nor U23882 (N_23882,N_20696,N_20533);
nor U23883 (N_23883,N_20450,N_20148);
or U23884 (N_23884,N_21229,N_20249);
nand U23885 (N_23885,N_21242,N_20917);
nand U23886 (N_23886,N_21238,N_21806);
or U23887 (N_23887,N_21659,N_21165);
nor U23888 (N_23888,N_20849,N_21024);
and U23889 (N_23889,N_20671,N_20460);
nor U23890 (N_23890,N_20855,N_20021);
nor U23891 (N_23891,N_21950,N_20717);
nand U23892 (N_23892,N_20915,N_21162);
nor U23893 (N_23893,N_20944,N_20361);
nor U23894 (N_23894,N_20686,N_21417);
xor U23895 (N_23895,N_20756,N_20381);
nand U23896 (N_23896,N_20807,N_21464);
or U23897 (N_23897,N_21411,N_20749);
or U23898 (N_23898,N_21480,N_21128);
nand U23899 (N_23899,N_20606,N_20442);
or U23900 (N_23900,N_20878,N_20264);
nor U23901 (N_23901,N_21078,N_21556);
nand U23902 (N_23902,N_21693,N_20352);
nand U23903 (N_23903,N_20071,N_20041);
or U23904 (N_23904,N_21980,N_21108);
xor U23905 (N_23905,N_20383,N_20325);
or U23906 (N_23906,N_20499,N_20926);
nor U23907 (N_23907,N_20775,N_21361);
and U23908 (N_23908,N_21030,N_21949);
nand U23909 (N_23909,N_20908,N_21623);
nand U23910 (N_23910,N_20141,N_21808);
nand U23911 (N_23911,N_20091,N_20993);
and U23912 (N_23912,N_21009,N_21489);
nor U23913 (N_23913,N_21274,N_21778);
nand U23914 (N_23914,N_21147,N_20572);
nor U23915 (N_23915,N_20753,N_20688);
or U23916 (N_23916,N_21584,N_20910);
and U23917 (N_23917,N_21710,N_21985);
nand U23918 (N_23918,N_20373,N_21724);
or U23919 (N_23919,N_21675,N_20780);
xor U23920 (N_23920,N_20294,N_20065);
nor U23921 (N_23921,N_20191,N_21130);
nand U23922 (N_23922,N_21015,N_21935);
xor U23923 (N_23923,N_20995,N_21560);
xnor U23924 (N_23924,N_20678,N_20754);
nor U23925 (N_23925,N_20257,N_21790);
and U23926 (N_23926,N_21778,N_20351);
nand U23927 (N_23927,N_21706,N_21874);
and U23928 (N_23928,N_21448,N_20168);
xnor U23929 (N_23929,N_20314,N_21290);
xnor U23930 (N_23930,N_21800,N_20714);
nand U23931 (N_23931,N_21859,N_21474);
nand U23932 (N_23932,N_21990,N_20254);
or U23933 (N_23933,N_21541,N_21813);
nand U23934 (N_23934,N_21878,N_20709);
and U23935 (N_23935,N_21758,N_20646);
or U23936 (N_23936,N_20621,N_20892);
nand U23937 (N_23937,N_21833,N_20558);
or U23938 (N_23938,N_21400,N_21640);
nand U23939 (N_23939,N_21541,N_20115);
nor U23940 (N_23940,N_21717,N_21997);
xnor U23941 (N_23941,N_21939,N_21352);
nand U23942 (N_23942,N_21888,N_20046);
nor U23943 (N_23943,N_20872,N_20854);
and U23944 (N_23944,N_20905,N_20629);
xor U23945 (N_23945,N_21201,N_21783);
or U23946 (N_23946,N_20550,N_20474);
nand U23947 (N_23947,N_20060,N_20173);
nand U23948 (N_23948,N_20883,N_20100);
or U23949 (N_23949,N_21598,N_21333);
nor U23950 (N_23950,N_20287,N_21805);
xnor U23951 (N_23951,N_20156,N_20743);
and U23952 (N_23952,N_20357,N_21340);
nor U23953 (N_23953,N_21066,N_21632);
xor U23954 (N_23954,N_20621,N_20371);
nand U23955 (N_23955,N_20462,N_20734);
nor U23956 (N_23956,N_20509,N_21995);
nand U23957 (N_23957,N_20368,N_20371);
nand U23958 (N_23958,N_21734,N_21610);
or U23959 (N_23959,N_21272,N_20475);
and U23960 (N_23960,N_21564,N_21882);
or U23961 (N_23961,N_21752,N_20569);
or U23962 (N_23962,N_20683,N_21578);
and U23963 (N_23963,N_20441,N_20585);
and U23964 (N_23964,N_21429,N_20162);
nand U23965 (N_23965,N_21612,N_20837);
or U23966 (N_23966,N_20383,N_20436);
nor U23967 (N_23967,N_20454,N_21797);
nand U23968 (N_23968,N_20482,N_20386);
nor U23969 (N_23969,N_20306,N_21817);
xor U23970 (N_23970,N_20392,N_20036);
and U23971 (N_23971,N_20618,N_20279);
and U23972 (N_23972,N_20728,N_20146);
nand U23973 (N_23973,N_20722,N_20526);
xor U23974 (N_23974,N_20388,N_20361);
nand U23975 (N_23975,N_21964,N_20722);
xor U23976 (N_23976,N_21297,N_20229);
and U23977 (N_23977,N_21213,N_20646);
xor U23978 (N_23978,N_21278,N_21131);
xor U23979 (N_23979,N_21189,N_20081);
xnor U23980 (N_23980,N_21658,N_20838);
nand U23981 (N_23981,N_20291,N_20376);
nand U23982 (N_23982,N_20268,N_20606);
and U23983 (N_23983,N_20831,N_21499);
and U23984 (N_23984,N_20034,N_21778);
and U23985 (N_23985,N_20925,N_20057);
nor U23986 (N_23986,N_20626,N_21813);
nand U23987 (N_23987,N_21520,N_20884);
or U23988 (N_23988,N_21680,N_21568);
nor U23989 (N_23989,N_20740,N_20639);
nand U23990 (N_23990,N_20918,N_20521);
or U23991 (N_23991,N_20740,N_21894);
or U23992 (N_23992,N_21755,N_20076);
and U23993 (N_23993,N_21229,N_20831);
nor U23994 (N_23994,N_20474,N_21018);
nand U23995 (N_23995,N_21128,N_20381);
nand U23996 (N_23996,N_21894,N_20738);
nor U23997 (N_23997,N_21884,N_20868);
nor U23998 (N_23998,N_21278,N_21649);
or U23999 (N_23999,N_20364,N_21341);
xnor U24000 (N_24000,N_23508,N_22017);
xnor U24001 (N_24001,N_22478,N_23721);
or U24002 (N_24002,N_23377,N_23396);
xnor U24003 (N_24003,N_22998,N_23639);
and U24004 (N_24004,N_23014,N_22952);
or U24005 (N_24005,N_23400,N_22908);
nand U24006 (N_24006,N_22672,N_23353);
or U24007 (N_24007,N_23903,N_23866);
nand U24008 (N_24008,N_22184,N_22535);
nor U24009 (N_24009,N_23781,N_22306);
or U24010 (N_24010,N_23130,N_22423);
nand U24011 (N_24011,N_23669,N_23934);
or U24012 (N_24012,N_23688,N_23730);
nand U24013 (N_24013,N_22863,N_22492);
or U24014 (N_24014,N_22240,N_23051);
and U24015 (N_24015,N_23239,N_23163);
xor U24016 (N_24016,N_22411,N_22586);
nand U24017 (N_24017,N_23324,N_22313);
nand U24018 (N_24018,N_22329,N_23339);
and U24019 (N_24019,N_23332,N_22805);
or U24020 (N_24020,N_22930,N_22500);
and U24021 (N_24021,N_22137,N_22747);
or U24022 (N_24022,N_23869,N_22258);
and U24023 (N_24023,N_22080,N_22364);
nor U24024 (N_24024,N_23712,N_22297);
and U24025 (N_24025,N_22657,N_23605);
or U24026 (N_24026,N_23567,N_23178);
and U24027 (N_24027,N_22516,N_22125);
nor U24028 (N_24028,N_23329,N_22558);
nor U24029 (N_24029,N_23804,N_22572);
and U24030 (N_24030,N_22565,N_23293);
nor U24031 (N_24031,N_22163,N_23547);
nand U24032 (N_24032,N_22990,N_22984);
and U24033 (N_24033,N_22269,N_23114);
or U24034 (N_24034,N_23938,N_23408);
xor U24035 (N_24035,N_22386,N_22161);
and U24036 (N_24036,N_22631,N_23728);
nor U24037 (N_24037,N_22376,N_23836);
nand U24038 (N_24038,N_22627,N_23162);
xnor U24039 (N_24039,N_22917,N_22488);
or U24040 (N_24040,N_23574,N_22911);
nand U24041 (N_24041,N_23224,N_23583);
and U24042 (N_24042,N_22771,N_22018);
or U24043 (N_24043,N_22206,N_23762);
nor U24044 (N_24044,N_22547,N_22868);
nand U24045 (N_24045,N_23538,N_23165);
xnor U24046 (N_24046,N_23283,N_22961);
or U24047 (N_24047,N_23455,N_23700);
nor U24048 (N_24048,N_23778,N_22044);
nor U24049 (N_24049,N_23169,N_22926);
xnor U24050 (N_24050,N_22587,N_23823);
or U24051 (N_24051,N_23735,N_22309);
or U24052 (N_24052,N_22997,N_22482);
or U24053 (N_24053,N_22605,N_23199);
and U24054 (N_24054,N_22864,N_22742);
and U24055 (N_24055,N_22877,N_23996);
nor U24056 (N_24056,N_23794,N_22828);
nand U24057 (N_24057,N_22344,N_23837);
or U24058 (N_24058,N_22729,N_22232);
nor U24059 (N_24059,N_23540,N_23173);
nand U24060 (N_24060,N_23141,N_22463);
or U24061 (N_24061,N_23854,N_23348);
nor U24062 (N_24062,N_23845,N_23280);
nand U24063 (N_24063,N_23187,N_23429);
nand U24064 (N_24064,N_23554,N_22429);
nor U24065 (N_24065,N_23608,N_22737);
xor U24066 (N_24066,N_23084,N_23120);
nor U24067 (N_24067,N_22455,N_23186);
and U24068 (N_24068,N_22073,N_23880);
nor U24069 (N_24069,N_23001,N_22860);
and U24070 (N_24070,N_23815,N_23589);
xnor U24071 (N_24071,N_22881,N_23537);
and U24072 (N_24072,N_22920,N_23419);
nand U24073 (N_24073,N_23058,N_23248);
xor U24074 (N_24074,N_22798,N_23358);
or U24075 (N_24075,N_23479,N_23500);
and U24076 (N_24076,N_22004,N_22359);
xnor U24077 (N_24077,N_23369,N_22584);
nand U24078 (N_24078,N_22788,N_22103);
xnor U24079 (N_24079,N_23595,N_23156);
or U24080 (N_24080,N_23963,N_23974);
nand U24081 (N_24081,N_23436,N_22902);
xor U24082 (N_24082,N_22635,N_22321);
nand U24083 (N_24083,N_22322,N_23428);
or U24084 (N_24084,N_22827,N_22424);
nand U24085 (N_24085,N_22611,N_23684);
nand U24086 (N_24086,N_22178,N_22343);
nand U24087 (N_24087,N_23502,N_22289);
or U24088 (N_24088,N_22550,N_22304);
xor U24089 (N_24089,N_22156,N_23264);
nor U24090 (N_24090,N_22314,N_22738);
nand U24091 (N_24091,N_23081,N_22569);
nor U24092 (N_24092,N_23300,N_23294);
or U24093 (N_24093,N_22140,N_23769);
or U24094 (N_24094,N_22234,N_23260);
and U24095 (N_24095,N_23102,N_22058);
nand U24096 (N_24096,N_23045,N_23009);
nor U24097 (N_24097,N_23219,N_22616);
and U24098 (N_24098,N_22981,N_23371);
and U24099 (N_24099,N_22172,N_23016);
nor U24100 (N_24100,N_23734,N_22277);
nand U24101 (N_24101,N_22882,N_22578);
or U24102 (N_24102,N_23343,N_22751);
nand U24103 (N_24103,N_23088,N_23074);
nand U24104 (N_24104,N_23747,N_22652);
nor U24105 (N_24105,N_22461,N_23126);
nor U24106 (N_24106,N_23720,N_22146);
nor U24107 (N_24107,N_23367,N_23862);
and U24108 (N_24108,N_22664,N_23767);
or U24109 (N_24109,N_22493,N_23690);
nor U24110 (N_24110,N_22727,N_23476);
nor U24111 (N_24111,N_22843,N_22370);
nand U24112 (N_24112,N_23237,N_22465);
nand U24113 (N_24113,N_22532,N_22462);
nand U24114 (N_24114,N_22392,N_23797);
nand U24115 (N_24115,N_22078,N_23822);
xnor U24116 (N_24116,N_23751,N_22119);
xor U24117 (N_24117,N_23898,N_23240);
xnor U24118 (N_24118,N_22399,N_23362);
and U24119 (N_24119,N_22043,N_23992);
and U24120 (N_24120,N_22921,N_23039);
xnor U24121 (N_24121,N_23401,N_23368);
xnor U24122 (N_24122,N_23327,N_23259);
nand U24123 (N_24123,N_22084,N_23139);
nand U24124 (N_24124,N_23775,N_22247);
xor U24125 (N_24125,N_22733,N_23023);
or U24126 (N_24126,N_23281,N_23956);
and U24127 (N_24127,N_23033,N_22754);
nand U24128 (N_24128,N_23653,N_23674);
xor U24129 (N_24129,N_22797,N_23415);
and U24130 (N_24130,N_22062,N_23939);
or U24131 (N_24131,N_22139,N_23911);
nand U24132 (N_24132,N_22000,N_23894);
and U24133 (N_24133,N_23168,N_22238);
and U24134 (N_24134,N_22342,N_23962);
nor U24135 (N_24135,N_22316,N_23179);
or U24136 (N_24136,N_23809,N_23873);
nor U24137 (N_24137,N_22481,N_23292);
nand U24138 (N_24138,N_23137,N_22046);
and U24139 (N_24139,N_22832,N_23662);
nor U24140 (N_24140,N_22900,N_22334);
nand U24141 (N_24141,N_22006,N_22336);
xor U24142 (N_24142,N_22702,N_22230);
nor U24143 (N_24143,N_22517,N_23525);
nand U24144 (N_24144,N_22726,N_23352);
or U24145 (N_24145,N_22677,N_22272);
xnor U24146 (N_24146,N_23454,N_22873);
nand U24147 (N_24147,N_22352,N_22113);
nand U24148 (N_24148,N_23875,N_22948);
nor U24149 (N_24149,N_22308,N_22590);
nor U24150 (N_24150,N_22714,N_23125);
nor U24151 (N_24151,N_22402,N_22824);
nor U24152 (N_24152,N_23807,N_22962);
nand U24153 (N_24153,N_22685,N_22955);
and U24154 (N_24154,N_22562,N_23780);
nor U24155 (N_24155,N_23610,N_23227);
nand U24156 (N_24156,N_22869,N_23622);
or U24157 (N_24157,N_23533,N_22471);
xor U24158 (N_24158,N_22118,N_23215);
nor U24159 (N_24159,N_23593,N_22435);
or U24160 (N_24160,N_23093,N_22668);
nand U24161 (N_24161,N_23979,N_23346);
xnor U24162 (N_24162,N_22709,N_23117);
xor U24163 (N_24163,N_23636,N_22872);
xor U24164 (N_24164,N_22225,N_23626);
and U24165 (N_24165,N_22151,N_23599);
or U24166 (N_24166,N_22212,N_22433);
nand U24167 (N_24167,N_23066,N_23450);
and U24168 (N_24168,N_23976,N_22169);
or U24169 (N_24169,N_23030,N_23201);
nand U24170 (N_24170,N_22598,N_23036);
xnor U24171 (N_24171,N_23810,N_23558);
xnor U24172 (N_24172,N_23695,N_22762);
nor U24173 (N_24173,N_22670,N_22106);
nand U24174 (N_24174,N_23407,N_22005);
or U24175 (N_24175,N_22434,N_23064);
xor U24176 (N_24176,N_22307,N_23548);
xor U24177 (N_24177,N_22905,N_23732);
or U24178 (N_24178,N_23801,N_22242);
or U24179 (N_24179,N_22656,N_22241);
nand U24180 (N_24180,N_22191,N_22899);
nand U24181 (N_24181,N_23038,N_22883);
xor U24182 (N_24182,N_23954,N_23345);
or U24183 (N_24183,N_23856,N_22780);
xnor U24184 (N_24184,N_23099,N_23303);
nand U24185 (N_24185,N_22394,N_23657);
nand U24186 (N_24186,N_22195,N_23266);
xor U24187 (N_24187,N_22730,N_22628);
nor U24188 (N_24188,N_23082,N_22270);
xor U24189 (N_24189,N_22132,N_22815);
or U24190 (N_24190,N_23889,N_23155);
nand U24191 (N_24191,N_22319,N_23258);
nor U24192 (N_24192,N_22085,N_22327);
and U24193 (N_24193,N_23566,N_23481);
and U24194 (N_24194,N_23390,N_22442);
nor U24195 (N_24195,N_23592,N_22328);
or U24196 (N_24196,N_23398,N_22875);
or U24197 (N_24197,N_23685,N_22126);
nand U24198 (N_24198,N_22444,N_22214);
or U24199 (N_24199,N_23793,N_23698);
nor U24200 (N_24200,N_23136,N_22404);
and U24201 (N_24201,N_23249,N_22360);
nand U24202 (N_24202,N_22735,N_22977);
and U24203 (N_24203,N_22989,N_22541);
and U24204 (N_24204,N_23406,N_23218);
nor U24205 (N_24205,N_23174,N_22077);
or U24206 (N_24206,N_22655,N_22796);
and U24207 (N_24207,N_22925,N_23032);
or U24208 (N_24208,N_23412,N_22661);
nor U24209 (N_24209,N_22032,N_22979);
nand U24210 (N_24210,N_23632,N_23262);
and U24211 (N_24211,N_23645,N_22098);
nand U24212 (N_24212,N_22676,N_23251);
xor U24213 (N_24213,N_23252,N_22378);
nand U24214 (N_24214,N_23555,N_23681);
nand U24215 (N_24215,N_23448,N_23531);
nor U24216 (N_24216,N_23587,N_23151);
xnor U24217 (N_24217,N_22120,N_22208);
nor U24218 (N_24218,N_22725,N_23335);
and U24219 (N_24219,N_22059,N_23005);
nand U24220 (N_24220,N_23637,N_22091);
and U24221 (N_24221,N_22207,N_23029);
xor U24222 (N_24222,N_22871,N_22839);
xor U24223 (N_24223,N_23946,N_22162);
and U24224 (N_24224,N_23590,N_23671);
nor U24225 (N_24225,N_23049,N_23176);
and U24226 (N_24226,N_23212,N_23432);
or U24227 (N_24227,N_22066,N_22333);
nand U24228 (N_24228,N_22781,N_23515);
xnor U24229 (N_24229,N_22669,N_23418);
nand U24230 (N_24230,N_22728,N_23693);
nor U24231 (N_24231,N_22255,N_22468);
nor U24232 (N_24232,N_22959,N_22422);
nor U24233 (N_24233,N_22681,N_22182);
and U24234 (N_24234,N_22494,N_23235);
and U24235 (N_24235,N_23598,N_22245);
nand U24236 (N_24236,N_23103,N_22618);
or U24237 (N_24237,N_22141,N_23988);
xnor U24238 (N_24238,N_23061,N_23675);
nor U24239 (N_24239,N_23146,N_22732);
xnor U24240 (N_24240,N_22713,N_22217);
xnor U24241 (N_24241,N_23184,N_22410);
nor U24242 (N_24242,N_22353,N_23276);
xor U24243 (N_24243,N_23618,N_22013);
or U24244 (N_24244,N_22564,N_23469);
or U24245 (N_24245,N_22001,N_22758);
nor U24246 (N_24246,N_23497,N_22679);
nand U24247 (N_24247,N_22480,N_22030);
or U24248 (N_24248,N_22470,N_22741);
nor U24249 (N_24249,N_23756,N_23376);
or U24250 (N_24250,N_22787,N_23982);
and U24251 (N_24251,N_23388,N_23763);
and U24252 (N_24252,N_22346,N_22160);
and U24253 (N_24253,N_23143,N_22008);
nor U24254 (N_24254,N_23973,N_22357);
and U24255 (N_24255,N_23314,N_22449);
xor U24256 (N_24256,N_23907,N_23070);
nand U24257 (N_24257,N_23511,N_23350);
nor U24258 (N_24258,N_22786,N_23777);
or U24259 (N_24259,N_23648,N_23483);
nand U24260 (N_24260,N_22074,N_23472);
nor U24261 (N_24261,N_22248,N_23792);
xor U24262 (N_24262,N_23062,N_22556);
xnor U24263 (N_24263,N_23572,N_22350);
nor U24264 (N_24264,N_23349,N_22042);
or U24265 (N_24265,N_23884,N_22348);
or U24266 (N_24266,N_23943,N_23167);
xor U24267 (N_24267,N_23286,N_22674);
and U24268 (N_24268,N_22094,N_22794);
or U24269 (N_24269,N_22266,N_22448);
xor U24270 (N_24270,N_22913,N_23312);
and U24271 (N_24271,N_23788,N_22064);
nand U24272 (N_24272,N_23409,N_23813);
nand U24273 (N_24273,N_23785,N_23570);
nor U24274 (N_24274,N_23449,N_22539);
or U24275 (N_24275,N_23468,N_23282);
xnor U24276 (N_24276,N_23296,N_22855);
xor U24277 (N_24277,N_23933,N_23319);
nor U24278 (N_24278,N_23516,N_22812);
nand U24279 (N_24279,N_23896,N_22823);
nor U24280 (N_24280,N_22789,N_23052);
and U24281 (N_24281,N_22703,N_22601);
nor U24282 (N_24282,N_22107,N_22596);
nand U24283 (N_24283,N_23656,N_22603);
xnor U24284 (N_24284,N_23112,N_23609);
nand U24285 (N_24285,N_22755,N_23098);
and U24286 (N_24286,N_22678,N_22756);
nand U24287 (N_24287,N_23037,N_22715);
and U24288 (N_24288,N_23440,N_22838);
or U24289 (N_24289,N_22570,N_22845);
nand U24290 (N_24290,N_23113,N_23274);
nor U24291 (N_24291,N_22957,N_22615);
and U24292 (N_24292,N_23147,N_22822);
xor U24293 (N_24293,N_22575,N_22560);
or U24294 (N_24294,N_23910,N_23275);
or U24295 (N_24295,N_22299,N_22439);
nand U24296 (N_24296,N_22581,N_22180);
nor U24297 (N_24297,N_22779,N_22190);
and U24298 (N_24298,N_22143,N_22278);
nand U24299 (N_24299,N_23999,N_23729);
nand U24300 (N_24300,N_22804,N_22858);
or U24301 (N_24301,N_22526,N_23160);
or U24302 (N_24302,N_23253,N_23509);
and U24303 (N_24303,N_23439,N_23072);
and U24304 (N_24304,N_23507,N_22183);
xor U24305 (N_24305,N_23825,N_23514);
nor U24306 (N_24306,N_22373,N_22795);
nor U24307 (N_24307,N_23188,N_22452);
nand U24308 (N_24308,N_22237,N_23024);
xor U24309 (N_24309,N_23007,N_22599);
and U24310 (N_24310,N_23978,N_22821);
xor U24311 (N_24311,N_22475,N_22358);
nor U24312 (N_24312,N_22573,N_22557);
xor U24313 (N_24313,N_23743,N_22450);
and U24314 (N_24314,N_23261,N_22019);
nor U24315 (N_24315,N_22415,N_22179);
nor U24316 (N_24316,N_23059,N_22813);
xor U24317 (N_24317,N_22852,N_22545);
nand U24318 (N_24318,N_23612,N_23389);
nor U24319 (N_24319,N_22923,N_23142);
nor U24320 (N_24320,N_23960,N_22110);
and U24321 (N_24321,N_22186,N_23847);
nor U24322 (N_24322,N_23620,N_23581);
or U24323 (N_24323,N_23707,N_23944);
or U24324 (N_24324,N_23647,N_22070);
nand U24325 (N_24325,N_22089,N_23393);
nor U24326 (N_24326,N_23158,N_22706);
and U24327 (N_24327,N_22651,N_23687);
nand U24328 (N_24328,N_22775,N_23272);
or U24329 (N_24329,N_23560,N_22721);
nor U24330 (N_24330,N_23927,N_22443);
and U24331 (N_24331,N_23307,N_23246);
or U24332 (N_24332,N_22673,N_22777);
nor U24333 (N_24333,N_23228,N_22338);
nor U24334 (N_24334,N_22458,N_22147);
nor U24335 (N_24335,N_23532,N_23107);
or U24336 (N_24336,N_23841,N_23949);
or U24337 (N_24337,N_22591,N_22181);
xnor U24338 (N_24338,N_23591,N_22885);
nor U24339 (N_24339,N_22226,N_23668);
xor U24340 (N_24340,N_22566,N_22381);
nand U24341 (N_24341,N_22551,N_22818);
nor U24342 (N_24342,N_23802,N_22039);
and U24343 (N_24343,N_23492,N_23364);
nand U24344 (N_24344,N_23263,N_22985);
xnor U24345 (N_24345,N_23488,N_22081);
nor U24346 (N_24346,N_23553,N_22154);
or U24347 (N_24347,N_23604,N_22014);
and U24348 (N_24348,N_23075,N_22649);
and U24349 (N_24349,N_23325,N_22093);
nor U24350 (N_24350,N_23152,N_22325);
nor U24351 (N_24351,N_23858,N_23421);
nor U24352 (N_24352,N_23706,N_22108);
and U24353 (N_24353,N_22159,N_23705);
xor U24354 (N_24354,N_23057,N_22960);
or U24355 (N_24355,N_23965,N_22451);
xor U24356 (N_24356,N_22896,N_22769);
or U24357 (N_24357,N_23185,N_23851);
nand U24358 (N_24358,N_22967,N_23597);
nand U24359 (N_24359,N_23341,N_22368);
nor U24360 (N_24360,N_23918,N_22809);
nor U24361 (N_24361,N_23676,N_22782);
nor U24362 (N_24362,N_22369,N_23855);
xnor U24363 (N_24363,N_22432,N_23213);
and U24364 (N_24364,N_22970,N_22683);
nand U24365 (N_24365,N_23122,N_22421);
or U24366 (N_24366,N_23824,N_22577);
xnor U24367 (N_24367,N_22974,N_22453);
xor U24368 (N_24368,N_22007,N_22192);
xor U24369 (N_24369,N_23857,N_23373);
and U24370 (N_24370,N_23530,N_22521);
nor U24371 (N_24371,N_22511,N_22665);
nor U24372 (N_24372,N_22700,N_22216);
nand U24373 (N_24373,N_22428,N_23050);
nand U24374 (N_24374,N_22847,N_22138);
and U24375 (N_24375,N_22175,N_23783);
xnor U24376 (N_24376,N_22221,N_22907);
nor U24377 (N_24377,N_23206,N_23926);
nor U24378 (N_24378,N_23990,N_22663);
and U24379 (N_24379,N_22764,N_22072);
and U24380 (N_24380,N_22354,N_23011);
nand U24381 (N_24381,N_22130,N_23026);
nor U24382 (N_24382,N_23055,N_23402);
nand U24383 (N_24383,N_22708,N_23629);
xnor U24384 (N_24384,N_23818,N_22994);
xnor U24385 (N_24385,N_23499,N_23193);
nor U24386 (N_24386,N_23754,N_22753);
nor U24387 (N_24387,N_23452,N_23053);
and U24388 (N_24388,N_22867,N_23733);
xnor U24389 (N_24389,N_22095,N_23475);
xor U24390 (N_24390,N_22928,N_23708);
nand U24391 (N_24391,N_22326,N_22637);
xnor U24392 (N_24392,N_23287,N_23717);
xnor U24393 (N_24393,N_22662,N_22318);
nand U24394 (N_24394,N_23094,N_22487);
and U24395 (N_24395,N_23427,N_23365);
nor U24396 (N_24396,N_23666,N_22379);
nor U24397 (N_24397,N_22459,N_22115);
and U24398 (N_24398,N_23607,N_23462);
nor U24399 (N_24399,N_22153,N_22534);
nand U24400 (N_24400,N_23195,N_22552);
nand U24401 (N_24401,N_22167,N_23087);
nand U24402 (N_24402,N_22978,N_23306);
or U24403 (N_24403,N_23265,N_22220);
or U24404 (N_24404,N_23196,N_22171);
nor U24405 (N_24405,N_22196,N_23344);
or U24406 (N_24406,N_23635,N_23380);
nand U24407 (N_24407,N_22740,N_22026);
or U24408 (N_24408,N_22231,N_22785);
nor U24409 (N_24409,N_23255,N_22529);
or U24410 (N_24410,N_23434,N_23812);
and U24411 (N_24411,N_23197,N_23640);
nand U24412 (N_24412,N_22667,N_23711);
nand U24413 (N_24413,N_23908,N_23441);
xor U24414 (N_24414,N_23459,N_23317);
nor U24415 (N_24415,N_23882,N_22071);
or U24416 (N_24416,N_22704,N_22722);
xnor U24417 (N_24417,N_23241,N_23715);
or U24418 (N_24418,N_23465,N_23897);
or U24419 (N_24419,N_22114,N_22388);
and U24420 (N_24420,N_23132,N_23017);
or U24421 (N_24421,N_22840,N_23776);
and U24422 (N_24422,N_22305,N_23138);
nor U24423 (N_24423,N_23998,N_23018);
nor U24424 (N_24424,N_22589,N_22718);
xnor U24425 (N_24425,N_23919,N_23904);
xnor U24426 (N_24426,N_22554,N_22976);
xnor U24427 (N_24427,N_23225,N_23646);
nor U24428 (N_24428,N_22609,N_23811);
xnor U24429 (N_24429,N_22524,N_23839);
or U24430 (N_24430,N_22880,N_22457);
nand U24431 (N_24431,N_23386,N_22284);
and U24432 (N_24432,N_23236,N_23972);
or U24433 (N_24433,N_22264,N_23539);
or U24434 (N_24434,N_23602,N_22879);
xnor U24435 (N_24435,N_23727,N_23411);
or U24436 (N_24436,N_23835,N_23105);
xnor U24437 (N_24437,N_23277,N_23526);
nand U24438 (N_24438,N_23931,N_22965);
and U24439 (N_24439,N_22472,N_23498);
and U24440 (N_24440,N_23370,N_23331);
and U24441 (N_24441,N_22279,N_22053);
xor U24442 (N_24442,N_22505,N_23718);
nand U24443 (N_24443,N_22810,N_22774);
or U24444 (N_24444,N_22011,N_22317);
xor U24445 (N_24445,N_22987,N_22111);
nor U24446 (N_24446,N_23920,N_23803);
or U24447 (N_24447,N_23496,N_23888);
or U24448 (N_24448,N_22536,N_22015);
or U24449 (N_24449,N_23861,N_22101);
nand U24450 (N_24450,N_23477,N_23381);
and U24451 (N_24451,N_22503,N_22403);
xor U24452 (N_24452,N_22105,N_22940);
nor U24453 (N_24453,N_23183,N_22945);
xnor U24454 (N_24454,N_22414,N_22134);
xor U24455 (N_24455,N_23063,N_22456);
and U24456 (N_24456,N_22016,N_23760);
and U24457 (N_24457,N_23773,N_23194);
nor U24458 (N_24458,N_23881,N_23003);
nor U24459 (N_24459,N_23028,N_23478);
nand U24460 (N_24460,N_23270,N_22265);
and U24461 (N_24461,N_23202,N_22387);
nor U24462 (N_24462,N_22744,N_23901);
xnor U24463 (N_24463,N_22128,N_22784);
xnor U24464 (N_24464,N_22276,N_22176);
nor U24465 (N_24465,N_22624,N_22501);
or U24466 (N_24466,N_22250,N_22363);
and U24467 (N_24467,N_23489,N_23971);
nor U24468 (N_24468,N_23772,N_22644);
nor U24469 (N_24469,N_22559,N_23546);
and U24470 (N_24470,N_23692,N_23221);
nor U24471 (N_24471,N_22502,N_23746);
nand U24472 (N_24472,N_22235,N_23615);
and U24473 (N_24473,N_23095,N_22097);
or U24474 (N_24474,N_23291,N_22942);
xnor U24475 (N_24475,N_22993,N_22604);
or U24476 (N_24476,N_23435,N_23031);
and U24477 (N_24477,N_22909,N_23921);
nor U24478 (N_24478,N_23359,N_23230);
xor U24479 (N_24479,N_22548,N_23131);
or U24480 (N_24480,N_23322,N_23736);
and U24481 (N_24481,N_22012,N_23046);
nand U24482 (N_24482,N_23594,N_22213);
nand U24483 (N_24483,N_23298,N_23832);
nor U24484 (N_24484,N_22983,N_22067);
and U24485 (N_24485,N_22876,N_23993);
nor U24486 (N_24486,N_23513,N_22968);
or U24487 (N_24487,N_23121,N_22853);
and U24488 (N_24488,N_23104,N_22254);
and U24489 (N_24489,N_23118,N_23153);
nor U24490 (N_24490,N_23820,N_23336);
or U24491 (N_24491,N_22198,N_22506);
nor U24492 (N_24492,N_22287,N_23422);
nand U24493 (N_24493,N_23086,N_23628);
or U24494 (N_24494,N_23437,N_22698);
xor U24495 (N_24495,N_23579,N_23947);
nand U24496 (N_24496,N_22746,N_23576);
or U24497 (N_24497,N_23774,N_22613);
or U24498 (N_24498,N_23784,N_22717);
and U24499 (N_24499,N_22129,N_22412);
nor U24500 (N_24500,N_23853,N_22922);
and U24501 (N_24501,N_23652,N_23724);
nor U24502 (N_24502,N_22303,N_23970);
and U24503 (N_24503,N_23744,N_22525);
nand U24504 (N_24504,N_22100,N_22766);
and U24505 (N_24505,N_22219,N_23796);
or U24506 (N_24506,N_23748,N_23892);
nor U24507 (N_24507,N_22311,N_23545);
xnor U24508 (N_24508,N_22020,N_23814);
xnor U24509 (N_24509,N_23768,N_22041);
nor U24510 (N_24510,N_22491,N_23269);
nand U24511 (N_24511,N_23234,N_22537);
and U24512 (N_24512,N_23713,N_22332);
nor U24513 (N_24513,N_22696,N_23577);
or U24514 (N_24514,N_22891,N_22654);
and U24515 (N_24515,N_22079,N_22750);
nor U24516 (N_24516,N_23582,N_23310);
xor U24517 (N_24517,N_23890,N_23200);
nand U24518 (N_24518,N_22104,N_23374);
nor U24519 (N_24519,N_22901,N_23683);
and U24520 (N_24520,N_22705,N_22933);
nor U24521 (N_24521,N_22692,N_22165);
or U24522 (N_24522,N_23651,N_23758);
nor U24523 (N_24523,N_22887,N_22800);
nor U24524 (N_24524,N_22257,N_22024);
nor U24525 (N_24525,N_23543,N_23115);
nand U24526 (N_24526,N_23643,N_23484);
nor U24527 (N_24527,N_23394,N_22324);
and U24528 (N_24528,N_22142,N_22793);
xor U24529 (N_24529,N_23827,N_22150);
nand U24530 (N_24530,N_23905,N_22274);
nor U24531 (N_24531,N_23969,N_23189);
or U24532 (N_24532,N_22215,N_22975);
or U24533 (N_24533,N_23642,N_23625);
xnor U24534 (N_24534,N_22916,N_23217);
nor U24535 (N_24535,N_22608,N_23416);
xor U24536 (N_24536,N_22477,N_22236);
and U24537 (N_24537,N_22931,N_22497);
nand U24538 (N_24538,N_23124,N_23865);
nor U24539 (N_24539,N_23127,N_23060);
xnor U24540 (N_24540,N_23667,N_22223);
nand U24541 (N_24541,N_22861,N_22966);
and U24542 (N_24542,N_22918,N_22919);
nand U24543 (N_24543,N_23504,N_23355);
nand U24544 (N_24544,N_23015,N_22910);
xnor U24545 (N_24545,N_22294,N_22894);
nand U24546 (N_24546,N_23925,N_22530);
xnor U24547 (N_24547,N_23968,N_23250);
xnor U24548 (N_24548,N_22496,N_23150);
nor U24549 (N_24549,N_22002,N_22914);
nand U24550 (N_24550,N_22602,N_22096);
xor U24551 (N_24551,N_22906,N_22383);
and U24552 (N_24552,N_22375,N_22009);
nor U24553 (N_24553,N_22341,N_23534);
xnor U24554 (N_24554,N_22136,N_22083);
nor U24555 (N_24555,N_22811,N_23425);
nand U24556 (N_24556,N_23523,N_23914);
nand U24557 (N_24557,N_23211,N_23782);
and U24558 (N_24558,N_22037,N_22723);
xor U24559 (N_24559,N_22831,N_22986);
or U24560 (N_24560,N_23922,N_23860);
or U24561 (N_24561,N_23940,N_22148);
and U24562 (N_24562,N_22281,N_22038);
nor U24563 (N_24563,N_23559,N_22124);
xor U24564 (N_24564,N_22406,N_22023);
nor U24565 (N_24565,N_23989,N_22082);
nor U24566 (N_24566,N_22340,N_23722);
nor U24567 (N_24567,N_23069,N_23012);
and U24568 (N_24568,N_22380,N_23691);
nor U24569 (N_24569,N_23334,N_22267);
xor U24570 (N_24570,N_23677,N_22050);
or U24571 (N_24571,N_22561,N_23229);
or U24572 (N_24572,N_23738,N_23673);
and U24573 (N_24573,N_22293,N_23297);
and U24574 (N_24574,N_22988,N_23661);
and U24575 (N_24575,N_22331,N_22634);
xor U24576 (N_24576,N_22301,N_22944);
nand U24577 (N_24577,N_22650,N_22315);
and U24578 (N_24578,N_22372,N_23220);
and U24579 (N_24579,N_23659,N_23458);
and U24580 (N_24580,N_23078,N_22389);
nor U24581 (N_24581,N_22620,N_22145);
nor U24582 (N_24582,N_23817,N_23315);
nand U24583 (N_24583,N_23385,N_23244);
xnor U24584 (N_24584,N_22036,N_23040);
nand U24585 (N_24585,N_23770,N_23843);
nand U24586 (N_24586,N_22991,N_23549);
nor U24587 (N_24587,N_23106,N_23544);
and U24588 (N_24588,N_22200,N_23161);
xor U24589 (N_24589,N_23603,N_23719);
nor U24590 (N_24590,N_22946,N_22850);
and U24591 (N_24591,N_23585,N_23065);
nand U24592 (N_24592,N_22320,N_22057);
nand U24593 (N_24593,N_23231,N_23703);
nand U24594 (N_24594,N_23709,N_23611);
nand U24595 (N_24595,N_22227,N_23453);
nor U24596 (N_24596,N_23360,N_23798);
nand U24597 (N_24597,N_23883,N_22210);
nor U24598 (N_24598,N_22187,N_23631);
nor U24599 (N_24599,N_23850,N_23980);
or U24600 (N_24600,N_22640,N_23948);
nor U24601 (N_24601,N_23140,N_22086);
or U24602 (N_24602,N_23906,N_23679);
or U24603 (N_24603,N_23575,N_23791);
or U24604 (N_24604,N_23382,N_23089);
and U24605 (N_24605,N_23446,N_22260);
and U24606 (N_24606,N_23305,N_23366);
and U24607 (N_24607,N_22772,N_23790);
nor U24608 (N_24608,N_22395,N_23493);
xnor U24609 (N_24609,N_22647,N_23828);
and U24610 (N_24610,N_23984,N_22606);
or U24611 (N_24611,N_23426,N_22710);
nor U24612 (N_24612,N_22712,N_22155);
nor U24613 (N_24613,N_23928,N_22298);
nor U24614 (N_24614,N_23096,N_22112);
nand U24615 (N_24615,N_22638,N_22574);
xnor U24616 (N_24616,N_23157,N_23145);
xnor U24617 (N_24617,N_23170,N_22523);
nor U24618 (N_24618,N_23830,N_23379);
or U24619 (N_24619,N_23417,N_22420);
nor U24620 (N_24620,N_22540,N_22518);
or U24621 (N_24621,N_22253,N_23243);
and U24622 (N_24622,N_22767,N_22865);
and U24623 (N_24623,N_22407,N_23464);
nor U24624 (N_24624,N_23986,N_23871);
xor U24625 (N_24625,N_22531,N_22801);
or U24626 (N_24626,N_23456,N_22312);
nor U24627 (N_24627,N_23073,N_23975);
xor U24628 (N_24628,N_23844,N_22438);
and U24629 (N_24629,N_23977,N_23356);
xor U24630 (N_24630,N_23682,N_22296);
xnor U24631 (N_24631,N_23311,N_23171);
xor U24632 (N_24632,N_22286,N_22202);
nor U24633 (N_24633,N_22642,N_23295);
nor U24634 (N_24634,N_23019,N_23872);
and U24635 (N_24635,N_23852,N_22460);
xnor U24636 (N_24636,N_23238,N_22870);
xor U24637 (N_24637,N_23868,N_22658);
xnor U24638 (N_24638,N_22413,N_23284);
nand U24639 (N_24639,N_23627,N_23342);
or U24640 (N_24640,N_23863,N_22636);
or U24641 (N_24641,N_23323,N_22251);
nand U24642 (N_24642,N_22109,N_22996);
xor U24643 (N_24643,N_23164,N_23689);
nor U24644 (N_24644,N_22600,N_23384);
or U24645 (N_24645,N_23564,N_22622);
nand U24646 (N_24646,N_22856,N_23787);
nor U24647 (N_24647,N_22648,N_23891);
nor U24648 (N_24648,N_22256,N_22205);
or U24649 (N_24649,N_23457,N_22844);
or U24650 (N_24650,N_22054,N_22123);
nor U24651 (N_24651,N_22623,N_23487);
and U24652 (N_24652,N_22859,N_23535);
nand U24653 (N_24653,N_22999,N_23877);
and U24654 (N_24654,N_22218,N_22197);
xnor U24655 (N_24655,N_22934,N_23375);
xor U24656 (N_24656,N_23936,N_23551);
xor U24657 (N_24657,N_23714,N_22739);
and U24658 (N_24658,N_22593,N_23886);
xnor U24659 (N_24659,N_23955,N_22133);
or U24660 (N_24660,N_23765,N_23867);
xor U24661 (N_24661,N_22047,N_22339);
xor U24662 (N_24662,N_23309,N_22228);
and U24663 (N_24663,N_22691,N_22897);
xnor U24664 (N_24664,N_23849,N_23829);
nor U24665 (N_24665,N_23461,N_22385);
or U24666 (N_24666,N_23759,N_23232);
and U24667 (N_24667,N_22833,N_23313);
xor U24668 (N_24668,N_23644,N_23299);
or U24669 (N_24669,N_22935,N_22031);
and U24670 (N_24670,N_22469,N_22483);
and U24671 (N_24671,N_22335,N_23964);
and U24672 (N_24672,N_22510,N_23166);
nand U24673 (N_24673,N_22610,N_22224);
and U24674 (N_24674,N_22173,N_22445);
or U24675 (N_24675,N_23083,N_23387);
or U24676 (N_24676,N_22088,N_22643);
nor U24677 (N_24677,N_23198,N_23207);
xnor U24678 (N_24678,N_23085,N_23601);
or U24679 (N_24679,N_23410,N_23725);
or U24680 (N_24680,N_22958,N_22612);
or U24681 (N_24681,N_22499,N_23068);
or U24682 (N_24682,N_23006,N_22268);
and U24683 (N_24683,N_22641,N_22862);
nand U24684 (N_24684,N_22121,N_23672);
nor U24685 (N_24685,N_22895,N_23789);
nand U24686 (N_24686,N_23347,N_23552);
nand U24687 (N_24687,N_22310,N_23800);
nand U24688 (N_24688,N_22356,N_22048);
xnor U24689 (N_24689,N_23318,N_23290);
or U24690 (N_24690,N_22440,N_22122);
nand U24691 (N_24691,N_22807,N_22166);
or U24692 (N_24692,N_22614,N_23893);
nor U24693 (N_24693,N_23354,N_22699);
nand U24694 (N_24694,N_23042,N_22087);
nor U24695 (N_24695,N_22446,N_23273);
or U24696 (N_24696,N_23361,N_23148);
nor U24697 (N_24697,N_23930,N_23338);
nor U24698 (N_24698,N_23431,N_22209);
nand U24699 (N_24699,N_23923,N_22571);
xor U24700 (N_24700,N_23204,N_22515);
nor U24701 (N_24701,N_22349,N_22969);
or U24702 (N_24702,N_22929,N_23180);
or U24703 (N_24703,N_23563,N_23519);
nor U24704 (N_24704,N_22936,N_23020);
and U24705 (N_24705,N_22052,N_22802);
nand U24706 (N_24706,N_22135,N_23779);
or U24707 (N_24707,N_23565,N_23233);
and U24708 (N_24708,N_23405,N_22816);
nand U24709 (N_24709,N_23753,N_22233);
and U24710 (N_24710,N_22203,N_23941);
and U24711 (N_24711,N_23080,N_23952);
nand U24712 (N_24712,N_23929,N_23378);
nand U24713 (N_24713,N_23092,N_22776);
or U24714 (N_24714,N_23430,N_22243);
nor U24715 (N_24715,N_22164,N_23002);
nand U24716 (N_24716,N_23494,N_22454);
nand U24717 (N_24717,N_23864,N_22904);
xor U24718 (N_24718,N_22585,N_22543);
or U24719 (N_24719,N_23466,N_23885);
xnor U24720 (N_24720,N_22690,N_23128);
or U24721 (N_24721,N_22127,N_22398);
xor U24722 (N_24722,N_23008,N_22393);
nor U24723 (N_24723,N_22061,N_23333);
nand U24724 (N_24724,N_22937,N_23924);
nand U24725 (N_24725,N_22711,N_22924);
xnor U24726 (N_24726,N_23247,N_22854);
and U24727 (N_24727,N_22849,N_22826);
and U24728 (N_24728,N_22367,N_23404);
nand U24729 (N_24729,N_23451,N_22416);
or U24730 (N_24730,N_22244,N_22168);
nor U24731 (N_24731,N_22594,N_23172);
or U24732 (N_24732,N_23134,N_23578);
and U24733 (N_24733,N_22639,N_23932);
xor U24734 (N_24734,N_22842,N_23686);
nor U24735 (N_24735,N_22527,N_23420);
xnor U24736 (N_24736,N_22973,N_23491);
nand U24737 (N_24737,N_22595,N_23702);
nand U24738 (N_24738,N_22426,N_23991);
nand U24739 (N_24739,N_22888,N_22437);
xnor U24740 (N_24740,N_23831,N_23022);
nor U24741 (N_24741,N_23848,N_23536);
xnor U24742 (N_24742,N_22028,N_23256);
xnor U24743 (N_24743,N_23222,N_23983);
xor U24744 (N_24744,N_22992,N_22629);
xor U24745 (N_24745,N_22719,N_22189);
nor U24746 (N_24746,N_23054,N_23226);
nand U24747 (N_24747,N_22157,N_23967);
xnor U24748 (N_24748,N_23288,N_23067);
nand U24749 (N_24749,N_22563,N_22544);
xnor U24750 (N_24750,N_23442,N_22273);
nor U24751 (N_24751,N_22972,N_23524);
and U24752 (N_24752,N_22391,N_23757);
or U24753 (N_24753,N_23895,N_22466);
and U24754 (N_24754,N_23522,N_22397);
xor U24755 (N_24755,N_22271,N_23761);
or U24756 (N_24756,N_23742,N_22886);
or U24757 (N_24757,N_23320,N_22889);
xnor U24758 (N_24758,N_23205,N_23580);
xor U24759 (N_24759,N_23289,N_22884);
nor U24760 (N_24760,N_23192,N_23665);
and U24761 (N_24761,N_22076,N_23528);
and U24762 (N_24762,N_22580,N_23208);
nor U24763 (N_24763,N_22659,N_23144);
nor U24764 (N_24764,N_22436,N_23953);
nor U24765 (N_24765,N_23878,N_22222);
xnor U24766 (N_24766,N_23859,N_22361);
or U24767 (N_24767,N_22418,N_22898);
or U24768 (N_24768,N_22366,N_22694);
xnor U24769 (N_24769,N_23047,N_23874);
nand U24770 (N_24770,N_22553,N_23606);
or U24771 (N_24771,N_23351,N_23985);
nand U24772 (N_24772,N_22430,N_22051);
nand U24773 (N_24773,N_22520,N_22878);
or U24774 (N_24774,N_22950,N_22029);
nand U24775 (N_24775,N_22743,N_23308);
and U24776 (N_24776,N_22249,N_22194);
nor U24777 (N_24777,N_23177,N_22390);
nand U24778 (N_24778,N_22408,N_23805);
or U24779 (N_24779,N_22857,N_23937);
nor U24780 (N_24780,N_23444,N_23808);
nor U24781 (N_24781,N_22300,N_22427);
nor U24782 (N_24782,N_22464,N_22405);
or U24783 (N_24783,N_23571,N_23614);
and U24784 (N_24784,N_22010,N_22174);
and U24785 (N_24785,N_23505,N_22964);
or U24786 (N_24786,N_22144,N_23749);
xnor U24787 (N_24787,N_23650,N_23994);
nand U24788 (N_24788,N_23301,N_22630);
xnor U24789 (N_24789,N_22090,N_23182);
nand U24790 (N_24790,N_22522,N_22045);
or U24791 (N_24791,N_22684,N_22971);
or U24792 (N_24792,N_22295,N_22396);
nor U24793 (N_24793,N_23541,N_22025);
nand U24794 (N_24794,N_22749,N_23586);
and U24795 (N_24795,N_22261,N_22285);
xor U24796 (N_24796,N_23027,N_22689);
nand U24797 (N_24797,N_22400,N_23658);
or U24798 (N_24798,N_22507,N_22830);
nor U24799 (N_24799,N_23568,N_22848);
and U24800 (N_24800,N_23490,N_23337);
nand U24801 (N_24801,N_23503,N_23694);
nor U24802 (N_24802,N_22660,N_22149);
xnor U24803 (N_24803,N_23518,N_23771);
nand U24804 (N_24804,N_23833,N_23048);
or U24805 (N_24805,N_22953,N_23834);
xor U24806 (N_24806,N_22290,N_23302);
and U24807 (N_24807,N_23501,N_22791);
or U24808 (N_24808,N_23819,N_22803);
nand U24809 (N_24809,N_23945,N_22778);
xnor U24810 (N_24810,N_22745,N_23223);
nor U24811 (N_24811,N_22204,N_23678);
nand U24812 (N_24812,N_23482,N_23271);
and U24813 (N_24813,N_23326,N_22377);
and U24814 (N_24814,N_23110,N_22263);
xnor U24815 (N_24815,N_23097,N_22687);
nor U24816 (N_24816,N_22890,N_23091);
nor U24817 (N_24817,N_23181,N_23654);
nor U24818 (N_24818,N_22474,N_23838);
nor U24819 (N_24819,N_22027,N_22542);
xor U24820 (N_24820,N_22695,N_23726);
nor U24821 (N_24821,N_23191,N_23701);
and U24822 (N_24822,N_22486,N_23902);
and U24823 (N_24823,N_23357,N_22504);
and U24824 (N_24824,N_22941,N_23795);
nor U24825 (N_24825,N_23704,N_23034);
and U24826 (N_24826,N_22567,N_23285);
or U24827 (N_24827,N_23013,N_23876);
nor U24828 (N_24828,N_23846,N_23995);
or U24829 (N_24829,N_23997,N_22763);
xnor U24830 (N_24830,N_23278,N_22382);
and U24831 (N_24831,N_23616,N_23447);
nand U24832 (N_24832,N_23633,N_22201);
nand U24833 (N_24833,N_23670,N_23664);
or U24834 (N_24834,N_22808,N_23395);
nand U24835 (N_24835,N_23573,N_22099);
and U24836 (N_24836,N_23000,N_22425);
nand U24837 (N_24837,N_22583,N_22302);
xnor U24838 (N_24838,N_23392,N_22773);
nand U24839 (N_24839,N_22371,N_22995);
nor U24840 (N_24840,N_22680,N_22597);
and U24841 (N_24841,N_23723,N_23043);
nor U24842 (N_24842,N_23279,N_23741);
nand U24843 (N_24843,N_22951,N_23619);
nor U24844 (N_24844,N_22549,N_22814);
or U24845 (N_24845,N_23242,N_22489);
and U24846 (N_24846,N_23363,N_22792);
or U24847 (N_24847,N_22579,N_23510);
or U24848 (N_24848,N_22607,N_23624);
nand U24849 (N_24849,N_22576,N_22193);
and U24850 (N_24850,N_22682,N_22055);
xnor U24851 (N_24851,N_22757,N_22441);
nand U24852 (N_24852,N_23630,N_22963);
or U24853 (N_24853,N_22765,N_23966);
and U24854 (N_24854,N_22783,N_23021);
and U24855 (N_24855,N_22943,N_23391);
nand U24856 (N_24856,N_22069,N_23542);
xor U24857 (N_24857,N_23879,N_23569);
or U24858 (N_24858,N_22799,N_23737);
nand U24859 (N_24859,N_23959,N_23842);
nor U24860 (N_24860,N_23981,N_22033);
xnor U24861 (N_24861,N_22513,N_23004);
xnor U24862 (N_24862,N_22075,N_23460);
and U24863 (N_24863,N_23413,N_23077);
or U24864 (N_24864,N_22282,N_22473);
and U24865 (N_24865,N_23950,N_23445);
and U24866 (N_24866,N_22927,N_23159);
and U24867 (N_24867,N_22841,N_23506);
nor U24868 (N_24868,N_22533,N_22035);
nand U24869 (N_24869,N_23399,N_23621);
xor U24870 (N_24870,N_23071,N_22065);
nor U24871 (N_24871,N_23100,N_23600);
and U24872 (N_24872,N_22625,N_22666);
nand U24873 (N_24873,N_23755,N_23699);
and U24874 (N_24874,N_23190,N_23584);
nor U24875 (N_24875,N_23101,N_22068);
nand U24876 (N_24876,N_22697,N_22485);
or U24877 (N_24877,N_22528,N_22021);
nand U24878 (N_24878,N_23520,N_22519);
or U24879 (N_24879,N_23696,N_23041);
nand U24880 (N_24880,N_22063,N_22806);
nand U24881 (N_24881,N_22056,N_22954);
nand U24882 (N_24882,N_23203,N_22819);
xnor U24883 (N_24883,N_22417,N_22748);
nor U24884 (N_24884,N_23438,N_23116);
nand U24885 (N_24885,N_23987,N_22246);
nor U24886 (N_24886,N_22323,N_22645);
and U24887 (N_24887,N_23245,N_22060);
or U24888 (N_24888,N_23557,N_22817);
or U24889 (N_24889,N_22626,N_22479);
nor U24890 (N_24890,N_23915,N_23916);
nor U24891 (N_24891,N_22419,N_22835);
xnor U24892 (N_24892,N_22834,N_22720);
or U24893 (N_24893,N_22003,N_22568);
nand U24894 (N_24894,N_23471,N_22837);
or U24895 (N_24895,N_23119,N_23517);
nor U24896 (N_24896,N_23254,N_22229);
and U24897 (N_24897,N_23467,N_22675);
nor U24898 (N_24898,N_23056,N_22467);
xnor U24899 (N_24899,N_22915,N_22939);
or U24900 (N_24900,N_23909,N_22337);
xnor U24901 (N_24901,N_23328,N_23826);
xor U24902 (N_24902,N_22736,N_23470);
xnor U24903 (N_24903,N_22384,N_22874);
nor U24904 (N_24904,N_23957,N_22932);
nand U24905 (N_24905,N_23216,N_23816);
nor U24906 (N_24906,N_23617,N_22508);
xor U24907 (N_24907,N_23806,N_22633);
and U24908 (N_24908,N_22707,N_23917);
nand U24909 (N_24909,N_23175,N_23655);
nand U24910 (N_24910,N_23316,N_23752);
xnor U24911 (N_24911,N_23840,N_23076);
nand U24912 (N_24912,N_22734,N_23958);
or U24913 (N_24913,N_22621,N_22825);
xnor U24914 (N_24914,N_22401,N_23821);
nand U24915 (N_24915,N_22912,N_23660);
nand U24916 (N_24916,N_22546,N_22022);
nand U24917 (N_24917,N_23268,N_23321);
or U24918 (N_24918,N_23330,N_22653);
and U24919 (N_24919,N_23766,N_22851);
or U24920 (N_24920,N_23154,N_23133);
or U24921 (N_24921,N_23550,N_23010);
and U24922 (N_24922,N_22538,N_23935);
nand U24923 (N_24923,N_22514,N_23870);
nor U24924 (N_24924,N_22351,N_23745);
xor U24925 (N_24925,N_22345,N_22283);
nor U24926 (N_24926,N_22355,N_22829);
nand U24927 (N_24927,N_23649,N_23799);
xor U24928 (N_24928,N_22582,N_23716);
and U24929 (N_24929,N_23111,N_23527);
and U24930 (N_24930,N_22291,N_22688);
or U24931 (N_24931,N_22761,N_22447);
nor U24932 (N_24932,N_23786,N_22770);
xor U24933 (N_24933,N_23562,N_22239);
or U24934 (N_24934,N_23641,N_22177);
nor U24935 (N_24935,N_23912,N_22131);
xnor U24936 (N_24936,N_22275,N_22555);
nor U24937 (N_24937,N_22724,N_23433);
nand U24938 (N_24938,N_22701,N_22512);
and U24939 (N_24939,N_22693,N_22619);
nand U24940 (N_24940,N_23556,N_22752);
xor U24941 (N_24941,N_23123,N_22185);
and U24942 (N_24942,N_22846,N_23596);
and U24943 (N_24943,N_22498,N_23521);
or U24944 (N_24944,N_23750,N_22956);
xnor U24945 (N_24945,N_22292,N_22431);
and U24946 (N_24946,N_23463,N_23423);
and U24947 (N_24947,N_22288,N_22040);
or U24948 (N_24948,N_22049,N_23109);
nor U24949 (N_24949,N_23529,N_23403);
and U24950 (N_24950,N_22892,N_22347);
nand U24951 (N_24951,N_23942,N_22409);
xor U24952 (N_24952,N_22982,N_23383);
or U24953 (N_24953,N_23340,N_23485);
or U24954 (N_24954,N_22117,N_22768);
and U24955 (N_24955,N_23414,N_22199);
or U24956 (N_24956,N_23913,N_23372);
xnor U24957 (N_24957,N_23588,N_23486);
and U24958 (N_24958,N_23561,N_22866);
and U24959 (N_24959,N_23900,N_22170);
and U24960 (N_24960,N_22790,N_23739);
or U24961 (N_24961,N_22759,N_23108);
nand U24962 (N_24962,N_22476,N_23638);
xnor U24963 (N_24963,N_23135,N_23025);
xnor U24964 (N_24964,N_22188,N_22592);
xor U24965 (N_24965,N_22820,N_23899);
xor U24966 (N_24966,N_22686,N_23397);
nor U24967 (N_24967,N_23512,N_23214);
nand U24968 (N_24968,N_22330,N_22484);
and U24969 (N_24969,N_22362,N_23035);
nor U24970 (N_24970,N_22116,N_23129);
xnor U24971 (N_24971,N_23663,N_22938);
xor U24972 (N_24972,N_22262,N_23079);
and U24973 (N_24973,N_22490,N_22980);
or U24974 (N_24974,N_22509,N_22646);
and U24975 (N_24975,N_23764,N_23210);
and U24976 (N_24976,N_22947,N_23887);
or U24977 (N_24977,N_22092,N_22259);
or U24978 (N_24978,N_23257,N_22034);
xor U24979 (N_24979,N_23443,N_23424);
nor U24980 (N_24980,N_22716,N_23480);
nor U24981 (N_24981,N_22365,N_22152);
nand U24982 (N_24982,N_23697,N_23680);
xnor U24983 (N_24983,N_23209,N_23495);
and U24984 (N_24984,N_23474,N_23710);
xor U24985 (N_24985,N_22903,N_23731);
or U24986 (N_24986,N_23044,N_22280);
nand U24987 (N_24987,N_23961,N_22588);
xor U24988 (N_24988,N_22760,N_22252);
xnor U24989 (N_24989,N_22731,N_22836);
nor U24990 (N_24990,N_22374,N_23613);
xor U24991 (N_24991,N_22102,N_22495);
or U24992 (N_24992,N_23267,N_22158);
xnor U24993 (N_24993,N_23090,N_23473);
and U24994 (N_24994,N_22893,N_23740);
or U24995 (N_24995,N_23149,N_22211);
and U24996 (N_24996,N_23634,N_23304);
nand U24997 (N_24997,N_23623,N_22632);
nand U24998 (N_24998,N_23951,N_22671);
and U24999 (N_24999,N_22949,N_22617);
xor U25000 (N_25000,N_22096,N_22949);
or U25001 (N_25001,N_22762,N_23275);
nor U25002 (N_25002,N_23951,N_23090);
nand U25003 (N_25003,N_23051,N_22410);
xnor U25004 (N_25004,N_23966,N_22750);
xnor U25005 (N_25005,N_22896,N_22159);
nor U25006 (N_25006,N_23799,N_23589);
and U25007 (N_25007,N_22429,N_23980);
xnor U25008 (N_25008,N_22048,N_22877);
nand U25009 (N_25009,N_22028,N_22481);
and U25010 (N_25010,N_23360,N_22834);
or U25011 (N_25011,N_23840,N_22971);
or U25012 (N_25012,N_23369,N_22985);
nand U25013 (N_25013,N_22236,N_23427);
and U25014 (N_25014,N_22065,N_22828);
xnor U25015 (N_25015,N_22443,N_22539);
xnor U25016 (N_25016,N_23372,N_22143);
nand U25017 (N_25017,N_22629,N_23163);
xor U25018 (N_25018,N_22711,N_23215);
nand U25019 (N_25019,N_23583,N_22862);
nor U25020 (N_25020,N_22036,N_22419);
nand U25021 (N_25021,N_22356,N_22711);
nor U25022 (N_25022,N_23030,N_23086);
or U25023 (N_25023,N_23238,N_22614);
or U25024 (N_25024,N_22125,N_22197);
xnor U25025 (N_25025,N_22427,N_22400);
or U25026 (N_25026,N_22057,N_23790);
and U25027 (N_25027,N_23042,N_23594);
nor U25028 (N_25028,N_22422,N_22033);
nand U25029 (N_25029,N_23295,N_23365);
and U25030 (N_25030,N_23536,N_23374);
and U25031 (N_25031,N_23954,N_23651);
and U25032 (N_25032,N_23159,N_22777);
and U25033 (N_25033,N_22819,N_22988);
and U25034 (N_25034,N_22541,N_23652);
and U25035 (N_25035,N_23455,N_22445);
nor U25036 (N_25036,N_22941,N_22166);
or U25037 (N_25037,N_22261,N_23629);
nor U25038 (N_25038,N_23690,N_23749);
xnor U25039 (N_25039,N_22005,N_22316);
and U25040 (N_25040,N_22425,N_23877);
nand U25041 (N_25041,N_22173,N_22203);
or U25042 (N_25042,N_23470,N_22080);
or U25043 (N_25043,N_23379,N_23473);
xor U25044 (N_25044,N_23357,N_22159);
nand U25045 (N_25045,N_23746,N_22864);
nand U25046 (N_25046,N_22361,N_23270);
xnor U25047 (N_25047,N_23693,N_22340);
nand U25048 (N_25048,N_23517,N_22339);
nand U25049 (N_25049,N_22975,N_23528);
nor U25050 (N_25050,N_23342,N_23811);
xor U25051 (N_25051,N_22334,N_22581);
xor U25052 (N_25052,N_22056,N_22895);
xor U25053 (N_25053,N_22262,N_22832);
or U25054 (N_25054,N_23383,N_23645);
or U25055 (N_25055,N_22656,N_23444);
nand U25056 (N_25056,N_23067,N_22001);
or U25057 (N_25057,N_22389,N_23973);
xnor U25058 (N_25058,N_22276,N_22477);
xor U25059 (N_25059,N_23615,N_22801);
or U25060 (N_25060,N_23198,N_22484);
nor U25061 (N_25061,N_22478,N_23383);
and U25062 (N_25062,N_22502,N_23379);
xor U25063 (N_25063,N_23159,N_22928);
nor U25064 (N_25064,N_23290,N_23001);
nor U25065 (N_25065,N_22893,N_23774);
or U25066 (N_25066,N_23499,N_23874);
or U25067 (N_25067,N_23881,N_23567);
nor U25068 (N_25068,N_22812,N_22017);
xnor U25069 (N_25069,N_23931,N_22948);
nor U25070 (N_25070,N_23796,N_23875);
nand U25071 (N_25071,N_23678,N_23111);
nor U25072 (N_25072,N_23614,N_23681);
xor U25073 (N_25073,N_22615,N_22911);
nor U25074 (N_25074,N_23028,N_22670);
nor U25075 (N_25075,N_23243,N_23441);
and U25076 (N_25076,N_23067,N_22890);
and U25077 (N_25077,N_23432,N_22874);
and U25078 (N_25078,N_22997,N_22208);
nand U25079 (N_25079,N_23092,N_22676);
nor U25080 (N_25080,N_22399,N_23317);
nand U25081 (N_25081,N_23583,N_23579);
nand U25082 (N_25082,N_22562,N_22842);
nor U25083 (N_25083,N_22045,N_23473);
and U25084 (N_25084,N_22046,N_23963);
or U25085 (N_25085,N_22877,N_22645);
nand U25086 (N_25086,N_22359,N_22876);
and U25087 (N_25087,N_22061,N_22660);
nor U25088 (N_25088,N_23251,N_23764);
and U25089 (N_25089,N_22128,N_22520);
or U25090 (N_25090,N_23972,N_22024);
nand U25091 (N_25091,N_22981,N_22099);
xor U25092 (N_25092,N_23843,N_23955);
or U25093 (N_25093,N_22622,N_22519);
nand U25094 (N_25094,N_22874,N_23630);
nor U25095 (N_25095,N_23165,N_23170);
or U25096 (N_25096,N_23328,N_22824);
or U25097 (N_25097,N_23079,N_23580);
nor U25098 (N_25098,N_23866,N_23209);
or U25099 (N_25099,N_22124,N_22089);
nand U25100 (N_25100,N_22469,N_23230);
and U25101 (N_25101,N_23405,N_23367);
xnor U25102 (N_25102,N_23705,N_23169);
or U25103 (N_25103,N_23075,N_23063);
nor U25104 (N_25104,N_22360,N_23264);
or U25105 (N_25105,N_22824,N_23547);
xor U25106 (N_25106,N_23870,N_22276);
xnor U25107 (N_25107,N_22547,N_22382);
xnor U25108 (N_25108,N_23564,N_23458);
or U25109 (N_25109,N_23209,N_22759);
and U25110 (N_25110,N_23185,N_22563);
xor U25111 (N_25111,N_23693,N_22540);
xor U25112 (N_25112,N_23358,N_22922);
and U25113 (N_25113,N_23732,N_23028);
or U25114 (N_25114,N_23268,N_22865);
and U25115 (N_25115,N_22027,N_22500);
nand U25116 (N_25116,N_23023,N_22366);
or U25117 (N_25117,N_23974,N_23866);
nor U25118 (N_25118,N_22521,N_23831);
nand U25119 (N_25119,N_23165,N_22462);
nand U25120 (N_25120,N_22711,N_23989);
nor U25121 (N_25121,N_23710,N_22989);
nand U25122 (N_25122,N_22966,N_23689);
xnor U25123 (N_25123,N_22328,N_23181);
and U25124 (N_25124,N_22814,N_22235);
nor U25125 (N_25125,N_22846,N_23291);
nand U25126 (N_25126,N_22364,N_22629);
xnor U25127 (N_25127,N_23162,N_23465);
or U25128 (N_25128,N_22527,N_22927);
and U25129 (N_25129,N_23579,N_23914);
or U25130 (N_25130,N_23506,N_22905);
nor U25131 (N_25131,N_23111,N_23900);
xor U25132 (N_25132,N_23287,N_22280);
and U25133 (N_25133,N_23071,N_22257);
xnor U25134 (N_25134,N_23383,N_23045);
nand U25135 (N_25135,N_22365,N_23304);
xor U25136 (N_25136,N_23721,N_23488);
nor U25137 (N_25137,N_22581,N_22870);
xnor U25138 (N_25138,N_22761,N_23725);
or U25139 (N_25139,N_22833,N_22001);
nand U25140 (N_25140,N_23832,N_22765);
nand U25141 (N_25141,N_23147,N_23405);
nor U25142 (N_25142,N_23688,N_22026);
or U25143 (N_25143,N_22408,N_22016);
xor U25144 (N_25144,N_23276,N_23147);
xnor U25145 (N_25145,N_22974,N_22506);
xnor U25146 (N_25146,N_22593,N_22010);
and U25147 (N_25147,N_23883,N_22816);
nand U25148 (N_25148,N_23529,N_22553);
and U25149 (N_25149,N_23213,N_22361);
and U25150 (N_25150,N_23770,N_23653);
nor U25151 (N_25151,N_22474,N_23392);
or U25152 (N_25152,N_22551,N_23470);
and U25153 (N_25153,N_23648,N_22637);
nand U25154 (N_25154,N_22662,N_22542);
or U25155 (N_25155,N_22233,N_22690);
nand U25156 (N_25156,N_23146,N_23181);
nand U25157 (N_25157,N_23857,N_22032);
nor U25158 (N_25158,N_23155,N_23286);
xnor U25159 (N_25159,N_23959,N_23856);
and U25160 (N_25160,N_23361,N_23225);
nand U25161 (N_25161,N_23105,N_23655);
nand U25162 (N_25162,N_23031,N_23628);
or U25163 (N_25163,N_22757,N_22587);
xnor U25164 (N_25164,N_22397,N_22665);
xnor U25165 (N_25165,N_23623,N_22062);
nor U25166 (N_25166,N_22991,N_23942);
nand U25167 (N_25167,N_22910,N_22112);
nand U25168 (N_25168,N_23562,N_22840);
and U25169 (N_25169,N_23412,N_22164);
or U25170 (N_25170,N_22399,N_22335);
nand U25171 (N_25171,N_23119,N_22044);
nand U25172 (N_25172,N_23392,N_22494);
or U25173 (N_25173,N_23609,N_22835);
or U25174 (N_25174,N_22241,N_22216);
xnor U25175 (N_25175,N_23925,N_22704);
and U25176 (N_25176,N_22889,N_23576);
or U25177 (N_25177,N_22393,N_22811);
nand U25178 (N_25178,N_23353,N_22446);
and U25179 (N_25179,N_22851,N_23077);
nand U25180 (N_25180,N_23138,N_23387);
and U25181 (N_25181,N_23739,N_22216);
nor U25182 (N_25182,N_22846,N_23961);
and U25183 (N_25183,N_23806,N_23841);
xor U25184 (N_25184,N_23170,N_22611);
nor U25185 (N_25185,N_22363,N_23183);
nand U25186 (N_25186,N_22608,N_23336);
nor U25187 (N_25187,N_23767,N_23903);
nor U25188 (N_25188,N_22368,N_22008);
and U25189 (N_25189,N_22766,N_22206);
nor U25190 (N_25190,N_22426,N_22763);
xor U25191 (N_25191,N_23318,N_22639);
xor U25192 (N_25192,N_22836,N_23793);
xnor U25193 (N_25193,N_22868,N_23452);
xor U25194 (N_25194,N_22732,N_22007);
xnor U25195 (N_25195,N_23921,N_23770);
or U25196 (N_25196,N_23641,N_22182);
nand U25197 (N_25197,N_23302,N_23567);
or U25198 (N_25198,N_23856,N_23098);
or U25199 (N_25199,N_22555,N_23303);
nor U25200 (N_25200,N_23933,N_23120);
xor U25201 (N_25201,N_22573,N_23612);
or U25202 (N_25202,N_23113,N_22751);
xnor U25203 (N_25203,N_23045,N_22695);
or U25204 (N_25204,N_23473,N_22431);
nor U25205 (N_25205,N_22124,N_22119);
nor U25206 (N_25206,N_22961,N_22580);
xor U25207 (N_25207,N_23799,N_23220);
and U25208 (N_25208,N_23317,N_22483);
nand U25209 (N_25209,N_22067,N_23668);
xnor U25210 (N_25210,N_23604,N_22506);
xor U25211 (N_25211,N_23614,N_22847);
and U25212 (N_25212,N_22681,N_22642);
xor U25213 (N_25213,N_22715,N_23499);
xor U25214 (N_25214,N_22402,N_22466);
or U25215 (N_25215,N_23550,N_23988);
or U25216 (N_25216,N_22010,N_22818);
or U25217 (N_25217,N_22783,N_22714);
xor U25218 (N_25218,N_23156,N_23663);
xnor U25219 (N_25219,N_22137,N_23991);
or U25220 (N_25220,N_22006,N_22286);
nor U25221 (N_25221,N_22309,N_23306);
xnor U25222 (N_25222,N_23269,N_23993);
or U25223 (N_25223,N_23195,N_22570);
or U25224 (N_25224,N_22823,N_23082);
or U25225 (N_25225,N_23921,N_22516);
xor U25226 (N_25226,N_22050,N_22569);
and U25227 (N_25227,N_23119,N_23714);
and U25228 (N_25228,N_23466,N_22029);
xor U25229 (N_25229,N_22120,N_23346);
nand U25230 (N_25230,N_23007,N_22530);
and U25231 (N_25231,N_23523,N_23387);
nand U25232 (N_25232,N_23761,N_23202);
xor U25233 (N_25233,N_22880,N_23095);
or U25234 (N_25234,N_22253,N_22866);
xor U25235 (N_25235,N_22762,N_22026);
and U25236 (N_25236,N_22159,N_23409);
or U25237 (N_25237,N_22245,N_23424);
and U25238 (N_25238,N_22157,N_23992);
xnor U25239 (N_25239,N_22659,N_23586);
or U25240 (N_25240,N_22107,N_23992);
xor U25241 (N_25241,N_22105,N_22089);
or U25242 (N_25242,N_23715,N_22064);
or U25243 (N_25243,N_23823,N_23640);
or U25244 (N_25244,N_23656,N_22437);
and U25245 (N_25245,N_22159,N_23788);
xor U25246 (N_25246,N_22691,N_23671);
or U25247 (N_25247,N_23625,N_23897);
xnor U25248 (N_25248,N_22483,N_23769);
nand U25249 (N_25249,N_22526,N_23212);
xnor U25250 (N_25250,N_23094,N_23510);
nor U25251 (N_25251,N_23331,N_22741);
or U25252 (N_25252,N_23411,N_23782);
nor U25253 (N_25253,N_23649,N_23829);
or U25254 (N_25254,N_22426,N_23266);
and U25255 (N_25255,N_23747,N_22791);
or U25256 (N_25256,N_23674,N_22841);
nor U25257 (N_25257,N_23532,N_23100);
xnor U25258 (N_25258,N_23315,N_23561);
or U25259 (N_25259,N_22745,N_22728);
and U25260 (N_25260,N_23642,N_23055);
nand U25261 (N_25261,N_23890,N_22478);
nor U25262 (N_25262,N_23967,N_23739);
xnor U25263 (N_25263,N_22304,N_22991);
and U25264 (N_25264,N_23949,N_22943);
and U25265 (N_25265,N_23287,N_22923);
nor U25266 (N_25266,N_23572,N_23062);
or U25267 (N_25267,N_23946,N_23752);
nor U25268 (N_25268,N_23228,N_23019);
nor U25269 (N_25269,N_22101,N_23765);
or U25270 (N_25270,N_23381,N_22027);
nand U25271 (N_25271,N_23155,N_22241);
nand U25272 (N_25272,N_22924,N_23641);
nor U25273 (N_25273,N_23788,N_22519);
or U25274 (N_25274,N_22499,N_23718);
nand U25275 (N_25275,N_23553,N_23783);
or U25276 (N_25276,N_23604,N_23127);
nand U25277 (N_25277,N_23984,N_23812);
xor U25278 (N_25278,N_23048,N_22655);
nor U25279 (N_25279,N_22952,N_23343);
nor U25280 (N_25280,N_23165,N_22951);
nor U25281 (N_25281,N_23865,N_22081);
nand U25282 (N_25282,N_22497,N_22734);
xnor U25283 (N_25283,N_22535,N_22029);
nor U25284 (N_25284,N_22825,N_23040);
nor U25285 (N_25285,N_22351,N_22051);
nor U25286 (N_25286,N_23110,N_23664);
nand U25287 (N_25287,N_22975,N_23688);
nand U25288 (N_25288,N_23344,N_22776);
nand U25289 (N_25289,N_23952,N_22049);
nand U25290 (N_25290,N_23876,N_22264);
or U25291 (N_25291,N_22280,N_22562);
and U25292 (N_25292,N_22921,N_22821);
or U25293 (N_25293,N_22801,N_23440);
nand U25294 (N_25294,N_23143,N_22136);
nand U25295 (N_25295,N_23781,N_22926);
or U25296 (N_25296,N_23559,N_22324);
and U25297 (N_25297,N_23853,N_22717);
xnor U25298 (N_25298,N_22204,N_22490);
and U25299 (N_25299,N_23669,N_23763);
xor U25300 (N_25300,N_22760,N_22410);
or U25301 (N_25301,N_22511,N_22763);
and U25302 (N_25302,N_23581,N_22951);
nand U25303 (N_25303,N_22393,N_23733);
and U25304 (N_25304,N_22936,N_23060);
nand U25305 (N_25305,N_22968,N_23165);
xnor U25306 (N_25306,N_23392,N_23932);
and U25307 (N_25307,N_23126,N_22435);
or U25308 (N_25308,N_22796,N_22928);
and U25309 (N_25309,N_23762,N_22025);
or U25310 (N_25310,N_22902,N_22338);
nand U25311 (N_25311,N_23937,N_22659);
nor U25312 (N_25312,N_23495,N_22125);
or U25313 (N_25313,N_22428,N_22972);
nand U25314 (N_25314,N_23082,N_23544);
nor U25315 (N_25315,N_22299,N_22062);
xor U25316 (N_25316,N_22002,N_23637);
and U25317 (N_25317,N_22800,N_23895);
nor U25318 (N_25318,N_22407,N_22402);
nand U25319 (N_25319,N_23617,N_23268);
nand U25320 (N_25320,N_22080,N_22943);
xnor U25321 (N_25321,N_23830,N_22829);
nor U25322 (N_25322,N_22698,N_22212);
xor U25323 (N_25323,N_22528,N_23816);
nand U25324 (N_25324,N_23899,N_22504);
xor U25325 (N_25325,N_22699,N_22566);
xnor U25326 (N_25326,N_23267,N_22538);
or U25327 (N_25327,N_22556,N_23317);
or U25328 (N_25328,N_23806,N_22191);
xor U25329 (N_25329,N_23065,N_23176);
xor U25330 (N_25330,N_22106,N_22703);
or U25331 (N_25331,N_23379,N_22004);
nor U25332 (N_25332,N_22072,N_22683);
nand U25333 (N_25333,N_23220,N_22681);
xnor U25334 (N_25334,N_22911,N_23674);
nor U25335 (N_25335,N_22384,N_22209);
nor U25336 (N_25336,N_22497,N_23043);
nand U25337 (N_25337,N_22781,N_23370);
nand U25338 (N_25338,N_23000,N_22228);
xor U25339 (N_25339,N_22201,N_22747);
and U25340 (N_25340,N_23323,N_22741);
nor U25341 (N_25341,N_23119,N_22793);
or U25342 (N_25342,N_22568,N_23240);
and U25343 (N_25343,N_22492,N_22663);
nor U25344 (N_25344,N_23675,N_23604);
and U25345 (N_25345,N_23530,N_23029);
or U25346 (N_25346,N_23848,N_23912);
nand U25347 (N_25347,N_22493,N_22082);
and U25348 (N_25348,N_23437,N_23106);
xnor U25349 (N_25349,N_23850,N_23450);
nor U25350 (N_25350,N_22053,N_23366);
or U25351 (N_25351,N_22251,N_23659);
and U25352 (N_25352,N_23254,N_23991);
and U25353 (N_25353,N_22480,N_22372);
nor U25354 (N_25354,N_22122,N_23073);
or U25355 (N_25355,N_22895,N_23463);
and U25356 (N_25356,N_23513,N_22297);
nor U25357 (N_25357,N_22786,N_23984);
or U25358 (N_25358,N_22951,N_22190);
nand U25359 (N_25359,N_22944,N_23507);
and U25360 (N_25360,N_22192,N_22117);
and U25361 (N_25361,N_22072,N_22895);
nor U25362 (N_25362,N_22428,N_22741);
xor U25363 (N_25363,N_22378,N_22949);
nor U25364 (N_25364,N_22289,N_23993);
xnor U25365 (N_25365,N_23218,N_22551);
nor U25366 (N_25366,N_23332,N_23585);
nor U25367 (N_25367,N_22532,N_23981);
and U25368 (N_25368,N_23428,N_22455);
nand U25369 (N_25369,N_23024,N_22205);
and U25370 (N_25370,N_22005,N_22649);
nand U25371 (N_25371,N_23407,N_22893);
nor U25372 (N_25372,N_22428,N_22167);
xor U25373 (N_25373,N_22535,N_23109);
xor U25374 (N_25374,N_23511,N_23697);
or U25375 (N_25375,N_22514,N_22323);
nor U25376 (N_25376,N_23639,N_22812);
or U25377 (N_25377,N_22930,N_23422);
or U25378 (N_25378,N_23737,N_23493);
or U25379 (N_25379,N_22647,N_22167);
or U25380 (N_25380,N_22859,N_23527);
nand U25381 (N_25381,N_23516,N_23850);
nand U25382 (N_25382,N_23089,N_22499);
or U25383 (N_25383,N_22507,N_22506);
nand U25384 (N_25384,N_22128,N_22545);
or U25385 (N_25385,N_23291,N_23149);
and U25386 (N_25386,N_22571,N_23075);
nand U25387 (N_25387,N_22989,N_22007);
or U25388 (N_25388,N_23477,N_23997);
nor U25389 (N_25389,N_22990,N_23317);
nand U25390 (N_25390,N_23285,N_22649);
and U25391 (N_25391,N_22417,N_23257);
nor U25392 (N_25392,N_23320,N_23281);
and U25393 (N_25393,N_22374,N_22798);
nor U25394 (N_25394,N_23967,N_23909);
nor U25395 (N_25395,N_22845,N_22378);
and U25396 (N_25396,N_23454,N_22893);
or U25397 (N_25397,N_22013,N_22382);
xnor U25398 (N_25398,N_22629,N_23560);
nor U25399 (N_25399,N_23736,N_22268);
and U25400 (N_25400,N_23969,N_22368);
or U25401 (N_25401,N_22560,N_22069);
xor U25402 (N_25402,N_22874,N_23961);
nand U25403 (N_25403,N_22299,N_23142);
xnor U25404 (N_25404,N_23702,N_22256);
xor U25405 (N_25405,N_23245,N_22405);
and U25406 (N_25406,N_23117,N_23770);
nand U25407 (N_25407,N_23853,N_22066);
nor U25408 (N_25408,N_23747,N_22801);
or U25409 (N_25409,N_22262,N_23718);
nor U25410 (N_25410,N_23046,N_23852);
xnor U25411 (N_25411,N_23529,N_22908);
or U25412 (N_25412,N_22895,N_23368);
or U25413 (N_25413,N_22948,N_22038);
and U25414 (N_25414,N_22756,N_22740);
and U25415 (N_25415,N_23780,N_22076);
xor U25416 (N_25416,N_23762,N_22269);
nor U25417 (N_25417,N_23023,N_22039);
xnor U25418 (N_25418,N_23075,N_23853);
xor U25419 (N_25419,N_23171,N_23667);
nand U25420 (N_25420,N_22684,N_23979);
nand U25421 (N_25421,N_23152,N_23118);
and U25422 (N_25422,N_23978,N_23737);
and U25423 (N_25423,N_22074,N_23551);
nor U25424 (N_25424,N_23702,N_23077);
xor U25425 (N_25425,N_23851,N_23705);
and U25426 (N_25426,N_23526,N_22577);
and U25427 (N_25427,N_23169,N_22610);
or U25428 (N_25428,N_22625,N_23841);
and U25429 (N_25429,N_23825,N_22826);
and U25430 (N_25430,N_22103,N_23335);
nor U25431 (N_25431,N_23362,N_23112);
nand U25432 (N_25432,N_23281,N_22844);
nor U25433 (N_25433,N_23067,N_23218);
nand U25434 (N_25434,N_22270,N_22856);
and U25435 (N_25435,N_23552,N_23581);
or U25436 (N_25436,N_23309,N_22722);
or U25437 (N_25437,N_23223,N_22225);
nor U25438 (N_25438,N_23273,N_22539);
xor U25439 (N_25439,N_23437,N_22955);
or U25440 (N_25440,N_22621,N_22549);
and U25441 (N_25441,N_22665,N_23828);
or U25442 (N_25442,N_22730,N_23494);
xnor U25443 (N_25443,N_22810,N_23970);
xnor U25444 (N_25444,N_23433,N_23094);
nand U25445 (N_25445,N_23048,N_22604);
nor U25446 (N_25446,N_22220,N_22434);
nand U25447 (N_25447,N_23851,N_23541);
xnor U25448 (N_25448,N_23305,N_22029);
xor U25449 (N_25449,N_22442,N_22632);
or U25450 (N_25450,N_22424,N_23706);
and U25451 (N_25451,N_22310,N_22935);
or U25452 (N_25452,N_22264,N_23042);
or U25453 (N_25453,N_22892,N_22799);
nand U25454 (N_25454,N_23396,N_23770);
or U25455 (N_25455,N_23715,N_22012);
and U25456 (N_25456,N_22999,N_23042);
and U25457 (N_25457,N_22499,N_23926);
and U25458 (N_25458,N_23931,N_23533);
and U25459 (N_25459,N_22016,N_23792);
nor U25460 (N_25460,N_23249,N_22589);
nor U25461 (N_25461,N_23536,N_22352);
nand U25462 (N_25462,N_22794,N_23151);
nand U25463 (N_25463,N_23177,N_22568);
and U25464 (N_25464,N_22527,N_23750);
and U25465 (N_25465,N_22171,N_23283);
xor U25466 (N_25466,N_22535,N_22414);
nand U25467 (N_25467,N_22132,N_22434);
nand U25468 (N_25468,N_22228,N_22971);
or U25469 (N_25469,N_22862,N_22087);
or U25470 (N_25470,N_22715,N_22374);
or U25471 (N_25471,N_22540,N_22508);
and U25472 (N_25472,N_22729,N_23180);
nand U25473 (N_25473,N_22795,N_23158);
and U25474 (N_25474,N_23286,N_23837);
xnor U25475 (N_25475,N_23541,N_23324);
or U25476 (N_25476,N_23188,N_22968);
or U25477 (N_25477,N_22504,N_23698);
xor U25478 (N_25478,N_23930,N_23487);
or U25479 (N_25479,N_22496,N_23788);
nor U25480 (N_25480,N_23554,N_22888);
and U25481 (N_25481,N_23386,N_23026);
and U25482 (N_25482,N_22487,N_22633);
xor U25483 (N_25483,N_23361,N_22473);
and U25484 (N_25484,N_22086,N_23161);
nand U25485 (N_25485,N_23856,N_23982);
nor U25486 (N_25486,N_23519,N_22982);
nand U25487 (N_25487,N_22821,N_22237);
and U25488 (N_25488,N_22040,N_23927);
xnor U25489 (N_25489,N_23027,N_22220);
nor U25490 (N_25490,N_22676,N_23135);
xor U25491 (N_25491,N_23658,N_23310);
and U25492 (N_25492,N_22455,N_22896);
nand U25493 (N_25493,N_22603,N_23376);
or U25494 (N_25494,N_22736,N_23069);
or U25495 (N_25495,N_23285,N_23148);
xor U25496 (N_25496,N_22904,N_23425);
nor U25497 (N_25497,N_23839,N_23168);
xor U25498 (N_25498,N_22530,N_23397);
xor U25499 (N_25499,N_22376,N_22984);
or U25500 (N_25500,N_22388,N_23716);
and U25501 (N_25501,N_23167,N_22260);
or U25502 (N_25502,N_23498,N_22382);
or U25503 (N_25503,N_22609,N_22289);
xor U25504 (N_25504,N_22848,N_22970);
nand U25505 (N_25505,N_23060,N_22167);
nor U25506 (N_25506,N_22362,N_23204);
nor U25507 (N_25507,N_23562,N_22372);
nand U25508 (N_25508,N_23137,N_23618);
nand U25509 (N_25509,N_23616,N_22105);
or U25510 (N_25510,N_23960,N_22248);
or U25511 (N_25511,N_23980,N_22482);
nor U25512 (N_25512,N_22480,N_22613);
or U25513 (N_25513,N_23126,N_23618);
xnor U25514 (N_25514,N_23612,N_23749);
xnor U25515 (N_25515,N_22979,N_23861);
nand U25516 (N_25516,N_23100,N_22752);
or U25517 (N_25517,N_23281,N_22486);
or U25518 (N_25518,N_22174,N_23502);
or U25519 (N_25519,N_22090,N_22664);
xnor U25520 (N_25520,N_22273,N_23226);
nor U25521 (N_25521,N_23576,N_22917);
xor U25522 (N_25522,N_23711,N_23633);
nor U25523 (N_25523,N_23971,N_22741);
xor U25524 (N_25524,N_22632,N_22252);
nor U25525 (N_25525,N_23237,N_22951);
xnor U25526 (N_25526,N_23853,N_22606);
or U25527 (N_25527,N_23589,N_22604);
xnor U25528 (N_25528,N_23395,N_23302);
nand U25529 (N_25529,N_22727,N_22569);
nor U25530 (N_25530,N_23583,N_22970);
nor U25531 (N_25531,N_23552,N_22647);
and U25532 (N_25532,N_22467,N_22928);
or U25533 (N_25533,N_23408,N_22199);
or U25534 (N_25534,N_22528,N_22523);
and U25535 (N_25535,N_22487,N_23657);
nor U25536 (N_25536,N_23524,N_23262);
xnor U25537 (N_25537,N_22586,N_23203);
nor U25538 (N_25538,N_23059,N_23219);
xor U25539 (N_25539,N_22392,N_22411);
nor U25540 (N_25540,N_22668,N_23606);
or U25541 (N_25541,N_22379,N_22473);
nor U25542 (N_25542,N_22350,N_22162);
or U25543 (N_25543,N_23204,N_23935);
nand U25544 (N_25544,N_22294,N_22020);
xnor U25545 (N_25545,N_22316,N_23067);
nand U25546 (N_25546,N_23478,N_22983);
nand U25547 (N_25547,N_22072,N_22252);
xnor U25548 (N_25548,N_22340,N_22294);
xor U25549 (N_25549,N_23643,N_22095);
or U25550 (N_25550,N_23396,N_23278);
nand U25551 (N_25551,N_23749,N_22378);
nand U25552 (N_25552,N_22557,N_22434);
xnor U25553 (N_25553,N_22764,N_23952);
and U25554 (N_25554,N_22065,N_22542);
or U25555 (N_25555,N_22955,N_23934);
and U25556 (N_25556,N_22646,N_22292);
and U25557 (N_25557,N_22912,N_23848);
nand U25558 (N_25558,N_23351,N_22484);
or U25559 (N_25559,N_22388,N_22781);
xnor U25560 (N_25560,N_22171,N_22235);
xnor U25561 (N_25561,N_23966,N_22834);
nand U25562 (N_25562,N_23922,N_23344);
xnor U25563 (N_25563,N_23773,N_22621);
xor U25564 (N_25564,N_22167,N_23856);
and U25565 (N_25565,N_22706,N_22897);
nand U25566 (N_25566,N_23653,N_23238);
or U25567 (N_25567,N_23113,N_23157);
xnor U25568 (N_25568,N_22922,N_22309);
nand U25569 (N_25569,N_22880,N_23700);
and U25570 (N_25570,N_22115,N_23774);
or U25571 (N_25571,N_23033,N_23155);
nand U25572 (N_25572,N_22109,N_23129);
or U25573 (N_25573,N_22398,N_22822);
nand U25574 (N_25574,N_23325,N_22300);
or U25575 (N_25575,N_23188,N_22268);
or U25576 (N_25576,N_23741,N_23045);
and U25577 (N_25577,N_22975,N_22565);
and U25578 (N_25578,N_23758,N_23047);
or U25579 (N_25579,N_23407,N_23813);
nor U25580 (N_25580,N_23676,N_23225);
nor U25581 (N_25581,N_23342,N_22262);
or U25582 (N_25582,N_22098,N_22862);
or U25583 (N_25583,N_22525,N_23896);
xnor U25584 (N_25584,N_23834,N_23724);
nor U25585 (N_25585,N_23559,N_23141);
nor U25586 (N_25586,N_22699,N_22980);
nand U25587 (N_25587,N_23835,N_23765);
xnor U25588 (N_25588,N_22443,N_23998);
and U25589 (N_25589,N_23934,N_22478);
or U25590 (N_25590,N_23765,N_23269);
and U25591 (N_25591,N_23855,N_22737);
and U25592 (N_25592,N_22615,N_23512);
and U25593 (N_25593,N_23915,N_22603);
nand U25594 (N_25594,N_23882,N_23260);
nor U25595 (N_25595,N_23550,N_22778);
or U25596 (N_25596,N_23628,N_23801);
xnor U25597 (N_25597,N_22643,N_23459);
or U25598 (N_25598,N_23036,N_23969);
xor U25599 (N_25599,N_22697,N_22561);
xor U25600 (N_25600,N_23360,N_23960);
xnor U25601 (N_25601,N_23571,N_22625);
or U25602 (N_25602,N_22536,N_22783);
nand U25603 (N_25603,N_22408,N_23311);
nor U25604 (N_25604,N_23283,N_22380);
or U25605 (N_25605,N_22809,N_23583);
or U25606 (N_25606,N_23402,N_23152);
and U25607 (N_25607,N_22976,N_22298);
or U25608 (N_25608,N_22465,N_23628);
nand U25609 (N_25609,N_23994,N_23631);
nor U25610 (N_25610,N_23936,N_22905);
nand U25611 (N_25611,N_23421,N_22491);
nor U25612 (N_25612,N_22359,N_23520);
or U25613 (N_25613,N_23519,N_23887);
or U25614 (N_25614,N_23157,N_22393);
nor U25615 (N_25615,N_23195,N_23230);
nand U25616 (N_25616,N_23049,N_23909);
nand U25617 (N_25617,N_22261,N_22061);
nand U25618 (N_25618,N_23008,N_23392);
or U25619 (N_25619,N_23165,N_22132);
xor U25620 (N_25620,N_23508,N_22135);
nand U25621 (N_25621,N_23276,N_23864);
or U25622 (N_25622,N_23025,N_22721);
xnor U25623 (N_25623,N_23900,N_22714);
and U25624 (N_25624,N_22556,N_22075);
nand U25625 (N_25625,N_22644,N_22548);
xor U25626 (N_25626,N_22229,N_22102);
and U25627 (N_25627,N_22982,N_22990);
or U25628 (N_25628,N_23361,N_22761);
nor U25629 (N_25629,N_23593,N_23805);
xor U25630 (N_25630,N_22603,N_23710);
and U25631 (N_25631,N_23545,N_22621);
nor U25632 (N_25632,N_23081,N_22856);
nor U25633 (N_25633,N_22926,N_22461);
nor U25634 (N_25634,N_23829,N_22685);
xor U25635 (N_25635,N_22303,N_23638);
or U25636 (N_25636,N_23096,N_23517);
xor U25637 (N_25637,N_22911,N_23020);
and U25638 (N_25638,N_23709,N_23092);
xnor U25639 (N_25639,N_22035,N_23495);
or U25640 (N_25640,N_23326,N_23671);
xnor U25641 (N_25641,N_22874,N_22994);
nor U25642 (N_25642,N_22693,N_23425);
nand U25643 (N_25643,N_23339,N_23199);
xnor U25644 (N_25644,N_23819,N_22748);
nand U25645 (N_25645,N_22066,N_22870);
and U25646 (N_25646,N_23798,N_22924);
xnor U25647 (N_25647,N_23243,N_22687);
nand U25648 (N_25648,N_22161,N_22393);
nand U25649 (N_25649,N_22541,N_22017);
nor U25650 (N_25650,N_22592,N_23404);
and U25651 (N_25651,N_23213,N_23792);
xor U25652 (N_25652,N_23629,N_23739);
and U25653 (N_25653,N_22647,N_23305);
nor U25654 (N_25654,N_22765,N_22649);
or U25655 (N_25655,N_22350,N_23442);
nand U25656 (N_25656,N_23580,N_22688);
or U25657 (N_25657,N_23701,N_23812);
and U25658 (N_25658,N_23091,N_22816);
xnor U25659 (N_25659,N_23322,N_22560);
nor U25660 (N_25660,N_22303,N_23407);
nand U25661 (N_25661,N_23640,N_22385);
nor U25662 (N_25662,N_23929,N_23524);
nand U25663 (N_25663,N_23317,N_22277);
xnor U25664 (N_25664,N_23503,N_22568);
xor U25665 (N_25665,N_23677,N_22802);
nor U25666 (N_25666,N_23131,N_22101);
or U25667 (N_25667,N_22785,N_23364);
nor U25668 (N_25668,N_22806,N_22293);
nor U25669 (N_25669,N_23644,N_23283);
and U25670 (N_25670,N_22468,N_22520);
nor U25671 (N_25671,N_23432,N_23423);
xor U25672 (N_25672,N_22309,N_22473);
nand U25673 (N_25673,N_22162,N_23334);
xor U25674 (N_25674,N_23372,N_23789);
nor U25675 (N_25675,N_23042,N_23280);
nor U25676 (N_25676,N_23283,N_23724);
or U25677 (N_25677,N_22209,N_22518);
xnor U25678 (N_25678,N_23524,N_23936);
or U25679 (N_25679,N_22508,N_22415);
or U25680 (N_25680,N_22109,N_22140);
nand U25681 (N_25681,N_22510,N_23841);
and U25682 (N_25682,N_23647,N_23920);
nand U25683 (N_25683,N_23546,N_23291);
and U25684 (N_25684,N_22817,N_23476);
or U25685 (N_25685,N_22803,N_23766);
nand U25686 (N_25686,N_23960,N_22373);
nand U25687 (N_25687,N_22274,N_22033);
xor U25688 (N_25688,N_23766,N_23525);
or U25689 (N_25689,N_23643,N_22291);
and U25690 (N_25690,N_22035,N_23566);
and U25691 (N_25691,N_22845,N_23982);
nor U25692 (N_25692,N_22203,N_22556);
or U25693 (N_25693,N_22903,N_23642);
and U25694 (N_25694,N_22905,N_22729);
nor U25695 (N_25695,N_23916,N_23993);
nand U25696 (N_25696,N_23370,N_22728);
and U25697 (N_25697,N_22811,N_22037);
or U25698 (N_25698,N_22250,N_23186);
and U25699 (N_25699,N_23245,N_22741);
xor U25700 (N_25700,N_23525,N_23310);
and U25701 (N_25701,N_23905,N_23345);
and U25702 (N_25702,N_23441,N_22060);
nand U25703 (N_25703,N_22031,N_22906);
nand U25704 (N_25704,N_22102,N_23067);
and U25705 (N_25705,N_22933,N_23213);
nand U25706 (N_25706,N_22366,N_23942);
nand U25707 (N_25707,N_22581,N_23725);
and U25708 (N_25708,N_23751,N_22558);
nor U25709 (N_25709,N_22680,N_23782);
or U25710 (N_25710,N_22066,N_23936);
xnor U25711 (N_25711,N_23660,N_23387);
or U25712 (N_25712,N_23167,N_23735);
xnor U25713 (N_25713,N_22232,N_23397);
or U25714 (N_25714,N_22076,N_23212);
or U25715 (N_25715,N_23163,N_22387);
nor U25716 (N_25716,N_22059,N_22917);
or U25717 (N_25717,N_22897,N_23991);
xnor U25718 (N_25718,N_22482,N_23927);
or U25719 (N_25719,N_22544,N_23553);
nand U25720 (N_25720,N_23708,N_23254);
xor U25721 (N_25721,N_22555,N_22286);
or U25722 (N_25722,N_23354,N_22207);
and U25723 (N_25723,N_22321,N_23368);
nor U25724 (N_25724,N_23381,N_23908);
nand U25725 (N_25725,N_22156,N_22902);
nand U25726 (N_25726,N_22410,N_22922);
nor U25727 (N_25727,N_23799,N_22250);
or U25728 (N_25728,N_22514,N_23615);
nand U25729 (N_25729,N_23088,N_23329);
xnor U25730 (N_25730,N_22959,N_22427);
or U25731 (N_25731,N_22250,N_22699);
or U25732 (N_25732,N_23417,N_23567);
nor U25733 (N_25733,N_22932,N_23145);
nand U25734 (N_25734,N_23015,N_23253);
nand U25735 (N_25735,N_22539,N_23302);
and U25736 (N_25736,N_23290,N_23730);
or U25737 (N_25737,N_22655,N_22286);
or U25738 (N_25738,N_23642,N_23897);
nor U25739 (N_25739,N_23616,N_22553);
or U25740 (N_25740,N_23716,N_23185);
nand U25741 (N_25741,N_22836,N_22263);
nor U25742 (N_25742,N_23435,N_22011);
and U25743 (N_25743,N_23020,N_22782);
or U25744 (N_25744,N_22144,N_23909);
or U25745 (N_25745,N_23283,N_23747);
nor U25746 (N_25746,N_22034,N_23699);
xor U25747 (N_25747,N_23911,N_22469);
xnor U25748 (N_25748,N_23034,N_22941);
nand U25749 (N_25749,N_22179,N_23690);
nor U25750 (N_25750,N_22138,N_23583);
and U25751 (N_25751,N_22284,N_23503);
nand U25752 (N_25752,N_22981,N_22566);
nand U25753 (N_25753,N_23562,N_23572);
nor U25754 (N_25754,N_22430,N_22470);
xnor U25755 (N_25755,N_22001,N_23652);
and U25756 (N_25756,N_22472,N_23487);
or U25757 (N_25757,N_22216,N_23098);
nor U25758 (N_25758,N_23067,N_22481);
or U25759 (N_25759,N_22764,N_22982);
nand U25760 (N_25760,N_23875,N_23793);
nor U25761 (N_25761,N_23716,N_23346);
nand U25762 (N_25762,N_22252,N_22478);
xnor U25763 (N_25763,N_23313,N_23595);
nand U25764 (N_25764,N_22259,N_22776);
or U25765 (N_25765,N_23717,N_23159);
or U25766 (N_25766,N_23677,N_23192);
and U25767 (N_25767,N_23790,N_22913);
or U25768 (N_25768,N_23575,N_23182);
xnor U25769 (N_25769,N_23406,N_23657);
and U25770 (N_25770,N_22166,N_22575);
nand U25771 (N_25771,N_22425,N_22979);
nand U25772 (N_25772,N_23559,N_23328);
xor U25773 (N_25773,N_22864,N_22713);
xor U25774 (N_25774,N_22997,N_22659);
nand U25775 (N_25775,N_22086,N_23151);
nor U25776 (N_25776,N_22476,N_23662);
nor U25777 (N_25777,N_22271,N_23730);
nor U25778 (N_25778,N_23882,N_23395);
nor U25779 (N_25779,N_23723,N_23154);
and U25780 (N_25780,N_22078,N_23595);
and U25781 (N_25781,N_22074,N_22187);
and U25782 (N_25782,N_22002,N_23219);
or U25783 (N_25783,N_22649,N_23141);
nor U25784 (N_25784,N_22349,N_23339);
nand U25785 (N_25785,N_22175,N_23330);
nand U25786 (N_25786,N_23107,N_23957);
nor U25787 (N_25787,N_23695,N_23169);
xnor U25788 (N_25788,N_23746,N_22392);
xor U25789 (N_25789,N_22627,N_23331);
and U25790 (N_25790,N_23422,N_23600);
and U25791 (N_25791,N_23640,N_22854);
nor U25792 (N_25792,N_23140,N_22363);
nor U25793 (N_25793,N_23499,N_23254);
or U25794 (N_25794,N_23748,N_22238);
or U25795 (N_25795,N_22486,N_23086);
nor U25796 (N_25796,N_23550,N_22812);
xor U25797 (N_25797,N_22188,N_22406);
nand U25798 (N_25798,N_22786,N_23524);
nor U25799 (N_25799,N_22897,N_23888);
xor U25800 (N_25800,N_23296,N_22970);
or U25801 (N_25801,N_22918,N_23275);
nand U25802 (N_25802,N_22004,N_22954);
and U25803 (N_25803,N_22838,N_23746);
xnor U25804 (N_25804,N_23530,N_22336);
or U25805 (N_25805,N_22774,N_23294);
or U25806 (N_25806,N_23699,N_23083);
nand U25807 (N_25807,N_23014,N_23397);
and U25808 (N_25808,N_23197,N_22586);
nand U25809 (N_25809,N_22008,N_22087);
nor U25810 (N_25810,N_22311,N_22854);
nor U25811 (N_25811,N_23970,N_22756);
xor U25812 (N_25812,N_22341,N_22111);
xnor U25813 (N_25813,N_22355,N_22791);
xor U25814 (N_25814,N_23349,N_23208);
xor U25815 (N_25815,N_22305,N_23689);
nor U25816 (N_25816,N_22543,N_23032);
or U25817 (N_25817,N_23962,N_23093);
nand U25818 (N_25818,N_22332,N_22898);
nor U25819 (N_25819,N_23755,N_23019);
nor U25820 (N_25820,N_22231,N_23056);
or U25821 (N_25821,N_23418,N_22372);
nor U25822 (N_25822,N_22510,N_23212);
xnor U25823 (N_25823,N_22035,N_23969);
and U25824 (N_25824,N_22680,N_22548);
nor U25825 (N_25825,N_23133,N_22634);
xnor U25826 (N_25826,N_22791,N_22845);
nand U25827 (N_25827,N_22471,N_23722);
nor U25828 (N_25828,N_23699,N_23750);
nor U25829 (N_25829,N_23610,N_23305);
nand U25830 (N_25830,N_22470,N_22172);
nor U25831 (N_25831,N_22921,N_22590);
or U25832 (N_25832,N_22619,N_22475);
or U25833 (N_25833,N_23270,N_22130);
xor U25834 (N_25834,N_22543,N_22476);
xor U25835 (N_25835,N_22765,N_23041);
xor U25836 (N_25836,N_23970,N_22528);
nor U25837 (N_25837,N_22985,N_22223);
or U25838 (N_25838,N_23909,N_22199);
or U25839 (N_25839,N_22317,N_23170);
and U25840 (N_25840,N_22815,N_22248);
xnor U25841 (N_25841,N_23596,N_22898);
or U25842 (N_25842,N_23274,N_23654);
nand U25843 (N_25843,N_22775,N_23201);
nor U25844 (N_25844,N_22427,N_22527);
nand U25845 (N_25845,N_23209,N_23034);
or U25846 (N_25846,N_22330,N_22682);
nand U25847 (N_25847,N_23104,N_22871);
and U25848 (N_25848,N_23298,N_22821);
and U25849 (N_25849,N_23073,N_22158);
xor U25850 (N_25850,N_23482,N_22827);
or U25851 (N_25851,N_23429,N_22594);
and U25852 (N_25852,N_22408,N_22414);
xor U25853 (N_25853,N_23426,N_22667);
xnor U25854 (N_25854,N_23772,N_23739);
and U25855 (N_25855,N_23925,N_22258);
nand U25856 (N_25856,N_22870,N_23880);
xor U25857 (N_25857,N_23618,N_23362);
nand U25858 (N_25858,N_22907,N_22269);
nand U25859 (N_25859,N_22203,N_22783);
nand U25860 (N_25860,N_23795,N_22048);
xor U25861 (N_25861,N_22149,N_22541);
or U25862 (N_25862,N_22785,N_22038);
xnor U25863 (N_25863,N_22079,N_23735);
and U25864 (N_25864,N_22875,N_22148);
nand U25865 (N_25865,N_22733,N_22127);
xnor U25866 (N_25866,N_23122,N_22830);
nor U25867 (N_25867,N_23730,N_23570);
xor U25868 (N_25868,N_23955,N_23500);
xnor U25869 (N_25869,N_22327,N_23932);
xor U25870 (N_25870,N_23535,N_23667);
or U25871 (N_25871,N_23756,N_23894);
xnor U25872 (N_25872,N_22012,N_23064);
nor U25873 (N_25873,N_22438,N_23872);
nor U25874 (N_25874,N_22031,N_22064);
nor U25875 (N_25875,N_23096,N_22951);
or U25876 (N_25876,N_22315,N_23035);
nor U25877 (N_25877,N_23021,N_22323);
nor U25878 (N_25878,N_22434,N_23520);
nand U25879 (N_25879,N_23689,N_22059);
and U25880 (N_25880,N_22650,N_22153);
or U25881 (N_25881,N_23183,N_23286);
xor U25882 (N_25882,N_22720,N_23664);
nand U25883 (N_25883,N_23284,N_23083);
nand U25884 (N_25884,N_22871,N_23177);
nor U25885 (N_25885,N_23801,N_22325);
nand U25886 (N_25886,N_22010,N_22347);
xnor U25887 (N_25887,N_22722,N_22813);
and U25888 (N_25888,N_22454,N_23228);
or U25889 (N_25889,N_23873,N_23921);
or U25890 (N_25890,N_23725,N_23563);
nand U25891 (N_25891,N_23920,N_22301);
nand U25892 (N_25892,N_22911,N_23459);
nand U25893 (N_25893,N_23138,N_23515);
nor U25894 (N_25894,N_22434,N_23915);
and U25895 (N_25895,N_23611,N_23601);
nor U25896 (N_25896,N_23223,N_23731);
and U25897 (N_25897,N_22638,N_22575);
nor U25898 (N_25898,N_22569,N_22391);
and U25899 (N_25899,N_22626,N_22604);
nand U25900 (N_25900,N_23035,N_22866);
or U25901 (N_25901,N_23471,N_22399);
or U25902 (N_25902,N_22302,N_22645);
and U25903 (N_25903,N_22287,N_22278);
xor U25904 (N_25904,N_23696,N_22613);
nor U25905 (N_25905,N_22861,N_23853);
and U25906 (N_25906,N_23335,N_22681);
nand U25907 (N_25907,N_23138,N_23316);
xnor U25908 (N_25908,N_23957,N_23863);
xor U25909 (N_25909,N_23772,N_22008);
xor U25910 (N_25910,N_23290,N_23657);
and U25911 (N_25911,N_23949,N_22119);
or U25912 (N_25912,N_22840,N_22629);
xor U25913 (N_25913,N_22931,N_23446);
nand U25914 (N_25914,N_22385,N_23153);
xor U25915 (N_25915,N_23416,N_23501);
nand U25916 (N_25916,N_22857,N_23224);
or U25917 (N_25917,N_23529,N_22487);
nand U25918 (N_25918,N_22721,N_23586);
nor U25919 (N_25919,N_22894,N_22828);
and U25920 (N_25920,N_23782,N_23421);
xnor U25921 (N_25921,N_22689,N_22104);
and U25922 (N_25922,N_22962,N_23104);
or U25923 (N_25923,N_22703,N_22594);
xnor U25924 (N_25924,N_22078,N_22971);
nand U25925 (N_25925,N_23131,N_23103);
xor U25926 (N_25926,N_23323,N_23562);
or U25927 (N_25927,N_22904,N_22238);
nor U25928 (N_25928,N_23333,N_23155);
nand U25929 (N_25929,N_23419,N_22131);
xnor U25930 (N_25930,N_22727,N_23251);
xor U25931 (N_25931,N_23417,N_22416);
or U25932 (N_25932,N_22693,N_23613);
and U25933 (N_25933,N_23130,N_22322);
xnor U25934 (N_25934,N_22326,N_23067);
xor U25935 (N_25935,N_23246,N_22424);
and U25936 (N_25936,N_22542,N_23690);
nor U25937 (N_25937,N_22591,N_23655);
and U25938 (N_25938,N_22564,N_23975);
nor U25939 (N_25939,N_22627,N_23726);
and U25940 (N_25940,N_23090,N_22758);
or U25941 (N_25941,N_22996,N_22204);
or U25942 (N_25942,N_22022,N_23227);
xor U25943 (N_25943,N_22181,N_23673);
nor U25944 (N_25944,N_22524,N_23687);
xor U25945 (N_25945,N_22547,N_23435);
or U25946 (N_25946,N_22735,N_23624);
nand U25947 (N_25947,N_23280,N_22479);
nor U25948 (N_25948,N_23209,N_23528);
xor U25949 (N_25949,N_23014,N_22518);
or U25950 (N_25950,N_23094,N_23046);
or U25951 (N_25951,N_22185,N_22403);
xor U25952 (N_25952,N_23186,N_22974);
and U25953 (N_25953,N_22196,N_23937);
xnor U25954 (N_25954,N_22857,N_22289);
xor U25955 (N_25955,N_23647,N_23994);
nand U25956 (N_25956,N_23811,N_23031);
xnor U25957 (N_25957,N_23391,N_22520);
nor U25958 (N_25958,N_23176,N_23478);
and U25959 (N_25959,N_22437,N_22467);
or U25960 (N_25960,N_22048,N_23952);
xor U25961 (N_25961,N_22705,N_23191);
or U25962 (N_25962,N_23305,N_22525);
or U25963 (N_25963,N_23397,N_22785);
nand U25964 (N_25964,N_22754,N_22476);
xor U25965 (N_25965,N_23343,N_23828);
nand U25966 (N_25966,N_22312,N_23092);
and U25967 (N_25967,N_23328,N_22395);
xnor U25968 (N_25968,N_22204,N_22413);
xor U25969 (N_25969,N_22814,N_23417);
xor U25970 (N_25970,N_23273,N_23398);
xor U25971 (N_25971,N_22382,N_22027);
or U25972 (N_25972,N_22909,N_22271);
nor U25973 (N_25973,N_23403,N_22698);
or U25974 (N_25974,N_23629,N_23252);
nor U25975 (N_25975,N_22303,N_23424);
xor U25976 (N_25976,N_23314,N_22466);
nand U25977 (N_25977,N_23205,N_22496);
nor U25978 (N_25978,N_22704,N_22655);
nor U25979 (N_25979,N_23392,N_23197);
or U25980 (N_25980,N_23087,N_23593);
and U25981 (N_25981,N_22779,N_23729);
and U25982 (N_25982,N_22156,N_23314);
and U25983 (N_25983,N_22871,N_22938);
or U25984 (N_25984,N_22800,N_22305);
or U25985 (N_25985,N_23097,N_22203);
xor U25986 (N_25986,N_22185,N_22454);
xor U25987 (N_25987,N_23941,N_23861);
or U25988 (N_25988,N_22198,N_23209);
and U25989 (N_25989,N_22148,N_22544);
nor U25990 (N_25990,N_22149,N_23468);
or U25991 (N_25991,N_23421,N_23251);
xor U25992 (N_25992,N_23524,N_22473);
nor U25993 (N_25993,N_22188,N_23058);
xor U25994 (N_25994,N_23564,N_23943);
xnor U25995 (N_25995,N_22839,N_23924);
or U25996 (N_25996,N_22971,N_22252);
xnor U25997 (N_25997,N_22930,N_23356);
nand U25998 (N_25998,N_22488,N_22749);
nand U25999 (N_25999,N_23542,N_23425);
nor U26000 (N_26000,N_24246,N_24534);
nor U26001 (N_26001,N_25098,N_24503);
and U26002 (N_26002,N_24376,N_25026);
nand U26003 (N_26003,N_25378,N_25107);
and U26004 (N_26004,N_24433,N_25917);
and U26005 (N_26005,N_25270,N_25096);
nand U26006 (N_26006,N_25703,N_25308);
nand U26007 (N_26007,N_25512,N_24483);
or U26008 (N_26008,N_24087,N_25733);
nand U26009 (N_26009,N_24167,N_24964);
nor U26010 (N_26010,N_25741,N_24439);
and U26011 (N_26011,N_24093,N_25545);
nor U26012 (N_26012,N_25236,N_24407);
or U26013 (N_26013,N_25557,N_24289);
nor U26014 (N_26014,N_25387,N_24787);
or U26015 (N_26015,N_25989,N_24318);
and U26016 (N_26016,N_25941,N_25625);
nand U26017 (N_26017,N_24430,N_25569);
and U26018 (N_26018,N_24987,N_25145);
or U26019 (N_26019,N_25413,N_24477);
or U26020 (N_26020,N_25393,N_24290);
and U26021 (N_26021,N_25597,N_25793);
xor U26022 (N_26022,N_24535,N_25876);
and U26023 (N_26023,N_25033,N_24123);
nand U26024 (N_26024,N_24938,N_24858);
xnor U26025 (N_26025,N_24736,N_25357);
or U26026 (N_26026,N_25209,N_24287);
and U26027 (N_26027,N_24546,N_24580);
or U26028 (N_26028,N_25503,N_24824);
or U26029 (N_26029,N_25656,N_25669);
nor U26030 (N_26030,N_24391,N_24868);
nor U26031 (N_26031,N_24423,N_24730);
xor U26032 (N_26032,N_24276,N_25037);
or U26033 (N_26033,N_25804,N_25817);
xor U26034 (N_26034,N_24993,N_24945);
xor U26035 (N_26035,N_25304,N_25662);
or U26036 (N_26036,N_24462,N_24136);
nand U26037 (N_26037,N_25577,N_25801);
or U26038 (N_26038,N_25161,N_25406);
nand U26039 (N_26039,N_24576,N_25551);
nand U26040 (N_26040,N_25836,N_24979);
nor U26041 (N_26041,N_24778,N_25157);
xor U26042 (N_26042,N_25115,N_24807);
or U26043 (N_26043,N_24811,N_25878);
or U26044 (N_26044,N_24268,N_24883);
xnor U26045 (N_26045,N_24659,N_24583);
nor U26046 (N_26046,N_25556,N_24822);
nand U26047 (N_26047,N_25409,N_25376);
and U26048 (N_26048,N_24022,N_25114);
or U26049 (N_26049,N_24984,N_25527);
xor U26050 (N_26050,N_24539,N_24080);
nor U26051 (N_26051,N_25666,N_24595);
nand U26052 (N_26052,N_25862,N_24820);
or U26053 (N_26053,N_24745,N_25663);
nand U26054 (N_26054,N_25926,N_25588);
nand U26055 (N_26055,N_24906,N_24602);
nor U26056 (N_26056,N_24163,N_25476);
nand U26057 (N_26057,N_25253,N_25701);
or U26058 (N_26058,N_24644,N_24085);
nand U26059 (N_26059,N_24177,N_24470);
and U26060 (N_26060,N_25920,N_25748);
or U26061 (N_26061,N_24734,N_25947);
xor U26062 (N_26062,N_24758,N_25453);
and U26063 (N_26063,N_24601,N_24058);
nor U26064 (N_26064,N_24670,N_24817);
nand U26065 (N_26065,N_25795,N_24489);
nor U26066 (N_26066,N_24281,N_24394);
xnor U26067 (N_26067,N_25097,N_24762);
or U26068 (N_26068,N_25062,N_24774);
or U26069 (N_26069,N_25080,N_25011);
nor U26070 (N_26070,N_25298,N_25574);
and U26071 (N_26071,N_24557,N_24231);
and U26072 (N_26072,N_24506,N_25605);
nor U26073 (N_26073,N_25398,N_24514);
or U26074 (N_26074,N_24213,N_24673);
xor U26075 (N_26075,N_24999,N_24755);
nor U26076 (N_26076,N_24959,N_25382);
and U26077 (N_26077,N_25294,N_24218);
or U26078 (N_26078,N_24666,N_25404);
xnor U26079 (N_26079,N_24860,N_25530);
nor U26080 (N_26080,N_25423,N_24401);
nand U26081 (N_26081,N_25054,N_24482);
nand U26082 (N_26082,N_25565,N_24299);
nor U26083 (N_26083,N_25699,N_25491);
and U26084 (N_26084,N_24886,N_25461);
xnor U26085 (N_26085,N_24083,N_25706);
nor U26086 (N_26086,N_25984,N_25639);
or U26087 (N_26087,N_24928,N_24708);
nand U26088 (N_26088,N_24063,N_25859);
nand U26089 (N_26089,N_25119,N_24252);
or U26090 (N_26090,N_25180,N_25620);
xor U26091 (N_26091,N_24584,N_25022);
nand U26092 (N_26092,N_25231,N_25071);
nand U26093 (N_26093,N_24799,N_24374);
or U26094 (N_26094,N_24074,N_24003);
nand U26095 (N_26095,N_25729,N_25192);
or U26096 (N_26096,N_25811,N_25002);
xnor U26097 (N_26097,N_25693,N_25200);
nor U26098 (N_26098,N_24371,N_25233);
xnor U26099 (N_26099,N_24570,N_25589);
nand U26100 (N_26100,N_24272,N_25865);
nor U26101 (N_26101,N_24419,N_25289);
or U26102 (N_26102,N_24235,N_25558);
xnor U26103 (N_26103,N_24622,N_25074);
xor U26104 (N_26104,N_24118,N_25609);
nor U26105 (N_26105,N_25221,N_25585);
xor U26106 (N_26106,N_24679,N_25362);
xnor U26107 (N_26107,N_24453,N_25228);
and U26108 (N_26108,N_25088,N_24322);
nor U26109 (N_26109,N_24922,N_25985);
nor U26110 (N_26110,N_24390,N_24344);
or U26111 (N_26111,N_24388,N_24712);
and U26112 (N_26112,N_24075,N_25126);
nand U26113 (N_26113,N_24171,N_25477);
or U26114 (N_26114,N_24264,N_25529);
xnor U26115 (N_26115,N_25894,N_24315);
and U26116 (N_26116,N_25132,N_24047);
nor U26117 (N_26117,N_24193,N_24400);
or U26118 (N_26118,N_25995,N_24744);
xor U26119 (N_26119,N_25861,N_25373);
nand U26120 (N_26120,N_24677,N_25389);
or U26121 (N_26121,N_24133,N_24809);
nor U26122 (N_26122,N_24802,N_25714);
xor U26123 (N_26123,N_24387,N_24784);
or U26124 (N_26124,N_24338,N_25388);
or U26125 (N_26125,N_25038,N_25246);
or U26126 (N_26126,N_24876,N_24782);
and U26127 (N_26127,N_25043,N_24366);
xnor U26128 (N_26128,N_25873,N_25055);
nor U26129 (N_26129,N_25903,N_24259);
xor U26130 (N_26130,N_25006,N_25945);
xnor U26131 (N_26131,N_25579,N_24950);
xnor U26132 (N_26132,N_25509,N_24944);
nor U26133 (N_26133,N_24530,N_25142);
nand U26134 (N_26134,N_24612,N_25902);
nor U26135 (N_26135,N_24236,N_25749);
or U26136 (N_26136,N_25268,N_25436);
xnor U26137 (N_26137,N_25705,N_25540);
or U26138 (N_26138,N_24362,N_24027);
nor U26139 (N_26139,N_24845,N_25069);
xor U26140 (N_26140,N_25694,N_25963);
nor U26141 (N_26141,N_25691,N_25980);
nor U26142 (N_26142,N_24375,N_24175);
or U26143 (N_26143,N_24096,N_25918);
nand U26144 (N_26144,N_24790,N_24020);
nand U26145 (N_26145,N_25602,N_25375);
or U26146 (N_26146,N_25300,N_25549);
nor U26147 (N_26147,N_25189,N_25201);
xor U26148 (N_26148,N_24701,N_25335);
nor U26149 (N_26149,N_25131,N_25879);
xnor U26150 (N_26150,N_24030,N_25784);
and U26151 (N_26151,N_24151,N_24088);
nand U26152 (N_26152,N_25402,N_25084);
nor U26153 (N_26153,N_25287,N_25970);
or U26154 (N_26154,N_24269,N_25892);
or U26155 (N_26155,N_24091,N_24705);
or U26156 (N_26156,N_25178,N_24295);
xnor U26157 (N_26157,N_25251,N_24494);
nor U26158 (N_26158,N_25356,N_24977);
nor U26159 (N_26159,N_25618,N_25645);
or U26160 (N_26160,N_25248,N_24207);
or U26161 (N_26161,N_25622,N_25773);
nor U26162 (N_26162,N_24053,N_25849);
nand U26163 (N_26163,N_25973,N_24351);
and U26164 (N_26164,N_24021,N_25360);
or U26165 (N_26165,N_25806,N_24927);
nor U26166 (N_26166,N_25944,N_24357);
nor U26167 (N_26167,N_24326,N_24940);
nor U26168 (N_26168,N_24077,N_24540);
nor U26169 (N_26169,N_24992,N_24880);
or U26170 (N_26170,N_25826,N_25151);
or U26171 (N_26171,N_25967,N_24198);
or U26172 (N_26172,N_25538,N_24324);
nor U26173 (N_26173,N_24909,N_25909);
nand U26174 (N_26174,N_25782,N_24455);
nand U26175 (N_26175,N_25722,N_25363);
xnor U26176 (N_26176,N_24352,N_24617);
or U26177 (N_26177,N_25257,N_25969);
or U26178 (N_26178,N_24104,N_25056);
nand U26179 (N_26179,N_25272,N_25981);
xnor U26180 (N_26180,N_25302,N_25689);
nor U26181 (N_26181,N_24624,N_24262);
xnor U26182 (N_26182,N_25658,N_24792);
and U26183 (N_26183,N_25156,N_24237);
xnor U26184 (N_26184,N_24835,N_24429);
nor U26185 (N_26185,N_24282,N_25960);
nand U26186 (N_26186,N_25939,N_25499);
nand U26187 (N_26187,N_25123,N_25634);
xnor U26188 (N_26188,N_24829,N_24998);
and U26189 (N_26189,N_24948,N_25717);
xor U26190 (N_26190,N_25174,N_25447);
or U26191 (N_26191,N_24628,N_25392);
and U26192 (N_26192,N_25290,N_25031);
nand U26193 (N_26193,N_24731,N_25009);
and U26194 (N_26194,N_24035,N_25803);
nand U26195 (N_26195,N_25050,N_24355);
and U26196 (N_26196,N_25737,N_24690);
and U26197 (N_26197,N_25396,N_24441);
and U26198 (N_26198,N_24051,N_24331);
nor U26199 (N_26199,N_25889,N_24187);
and U26200 (N_26200,N_24781,N_24191);
xor U26201 (N_26201,N_24941,N_25715);
and U26202 (N_26202,N_24816,N_25925);
and U26203 (N_26203,N_25815,N_25912);
or U26204 (N_26204,N_25866,N_24848);
and U26205 (N_26205,N_25188,N_24052);
and U26206 (N_26206,N_25172,N_25506);
xor U26207 (N_26207,N_25590,N_24660);
xnor U26208 (N_26208,N_24966,N_24891);
and U26209 (N_26209,N_24432,N_24188);
xor U26210 (N_26210,N_24159,N_25489);
nor U26211 (N_26211,N_24378,N_24751);
nor U26212 (N_26212,N_25800,N_24084);
xor U26213 (N_26213,N_25421,N_25948);
xor U26214 (N_26214,N_25510,N_24241);
or U26215 (N_26215,N_24367,N_25137);
nor U26216 (N_26216,N_25734,N_24898);
nand U26217 (N_26217,N_25553,N_25345);
or U26218 (N_26218,N_25845,N_25352);
or U26219 (N_26219,N_24438,N_24797);
nor U26220 (N_26220,N_24346,N_24460);
xnor U26221 (N_26221,N_24650,N_24105);
and U26222 (N_26222,N_25511,N_25853);
nand U26223 (N_26223,N_24431,N_24975);
nor U26224 (N_26224,N_25008,N_25343);
or U26225 (N_26225,N_25924,N_24386);
nor U26226 (N_26226,N_25518,N_24448);
or U26227 (N_26227,N_24568,N_25735);
nand U26228 (N_26228,N_25213,N_24435);
and U26229 (N_26229,N_24564,N_25668);
or U26230 (N_26230,N_25988,N_24109);
xnor U26231 (N_26231,N_25998,N_25014);
nand U26232 (N_26232,N_25887,N_24526);
nor U26233 (N_26233,N_24095,N_24541);
nand U26234 (N_26234,N_25670,N_25724);
or U26235 (N_26235,N_25064,N_25850);
nor U26236 (N_26236,N_24204,N_25768);
xor U26237 (N_26237,N_25643,N_24862);
or U26238 (N_26238,N_24960,N_25312);
nand U26239 (N_26239,N_24256,N_25697);
xnor U26240 (N_26240,N_24142,N_25567);
nor U26241 (N_26241,N_25316,N_25394);
xor U26242 (N_26242,N_25310,N_24900);
or U26243 (N_26243,N_25010,N_25792);
nand U26244 (N_26244,N_24559,N_25383);
nand U26245 (N_26245,N_25539,N_24878);
xor U26246 (N_26246,N_24416,N_24411);
and U26247 (N_26247,N_24072,N_25429);
and U26248 (N_26248,N_24094,N_24957);
and U26249 (N_26249,N_25032,N_24718);
nand U26250 (N_26250,N_24573,N_25802);
and U26251 (N_26251,N_24556,N_25323);
nand U26252 (N_26252,N_25730,N_25030);
nand U26253 (N_26253,N_24680,N_24059);
and U26254 (N_26254,N_24578,N_24041);
nor U26255 (N_26255,N_25437,N_25515);
or U26256 (N_26256,N_24565,N_25522);
and U26257 (N_26257,N_24582,N_25281);
xor U26258 (N_26258,N_25058,N_24552);
and U26259 (N_26259,N_24682,N_24464);
xor U26260 (N_26260,N_24491,N_25053);
or U26261 (N_26261,N_24261,N_24365);
nor U26262 (N_26262,N_25163,N_25752);
nand U26263 (N_26263,N_24769,N_24046);
xor U26264 (N_26264,N_25570,N_25355);
xnor U26265 (N_26265,N_25994,N_24476);
nor U26266 (N_26266,N_25872,N_24888);
or U26267 (N_26267,N_25600,N_25313);
xnor U26268 (N_26268,N_24078,N_25481);
nand U26269 (N_26269,N_25035,N_24457);
nor U26270 (N_26270,N_25883,N_24801);
and U26271 (N_26271,N_24152,N_24498);
xnor U26272 (N_26272,N_25259,N_25346);
and U26273 (N_26273,N_25440,N_24819);
and U26274 (N_26274,N_25915,N_25710);
nand U26275 (N_26275,N_25756,N_24990);
and U26276 (N_26276,N_24361,N_24120);
and U26277 (N_26277,N_24250,N_25168);
and U26278 (N_26278,N_24525,N_24651);
nor U26279 (N_26279,N_24134,N_24309);
or U26280 (N_26280,N_25068,N_24024);
nor U26281 (N_26281,N_25677,N_24590);
and U26282 (N_26282,N_24086,N_25432);
nand U26283 (N_26283,N_24840,N_24759);
xor U26284 (N_26284,N_25513,N_25454);
nand U26285 (N_26285,N_25934,N_25207);
nor U26286 (N_26286,N_24234,N_24638);
nor U26287 (N_26287,N_24861,N_25000);
or U26288 (N_26288,N_24469,N_24837);
xnor U26289 (N_26289,N_24828,N_25854);
nor U26290 (N_26290,N_24221,N_25573);
xor U26291 (N_26291,N_24995,N_25249);
nand U26292 (N_26292,N_25910,N_25520);
or U26293 (N_26293,N_25514,N_24872);
xnor U26294 (N_26294,N_25435,N_24722);
nor U26295 (N_26295,N_25542,N_25480);
nor U26296 (N_26296,N_24254,N_25780);
nor U26297 (N_26297,N_24776,N_24200);
nor U26298 (N_26298,N_25462,N_25630);
xnor U26299 (N_26299,N_24846,N_24292);
nand U26300 (N_26300,N_24709,N_24418);
or U26301 (N_26301,N_25239,N_24255);
nand U26302 (N_26302,N_25841,N_25566);
or U26303 (N_26303,N_25198,N_24173);
nor U26304 (N_26304,N_25834,N_24572);
and U26305 (N_26305,N_25875,N_25046);
nor U26306 (N_26306,N_25659,N_25606);
or U26307 (N_26307,N_25610,N_25400);
or U26308 (N_26308,N_25830,N_25505);
nand U26309 (N_26309,N_25870,N_24994);
nor U26310 (N_26310,N_24353,N_24753);
and U26311 (N_26311,N_24288,N_25017);
and U26312 (N_26312,N_24678,N_25087);
nor U26313 (N_26313,N_25134,N_25066);
xnor U26314 (N_26314,N_24521,N_24903);
and U26315 (N_26315,N_24851,N_25607);
nand U26316 (N_26316,N_25457,N_25391);
nor U26317 (N_26317,N_25837,N_24267);
nor U26318 (N_26318,N_25208,N_25637);
and U26319 (N_26319,N_25018,N_25472);
or U26320 (N_26320,N_24038,N_24935);
nand U26321 (N_26321,N_25500,N_25040);
nor U26322 (N_26322,N_25334,N_24114);
nor U26323 (N_26323,N_24836,N_25293);
or U26324 (N_26324,N_24519,N_24695);
xnor U26325 (N_26325,N_25578,N_25379);
or U26326 (N_26326,N_25229,N_25195);
nor U26327 (N_26327,N_24765,N_24833);
nand U26328 (N_26328,N_24146,N_25349);
nor U26329 (N_26329,N_24686,N_24547);
nor U26330 (N_26330,N_24757,N_25593);
or U26331 (N_26331,N_25633,N_25754);
or U26332 (N_26332,N_25237,N_24796);
nor U26333 (N_26333,N_24025,N_24749);
nor U26334 (N_26334,N_24916,N_24517);
and U26335 (N_26335,N_24283,N_24581);
xor U26336 (N_26336,N_25561,N_24332);
nor U26337 (N_26337,N_25446,N_24982);
nor U26338 (N_26338,N_24766,N_25616);
nor U26339 (N_26339,N_24634,N_24536);
xor U26340 (N_26340,N_24485,N_24885);
nand U26341 (N_26341,N_24504,N_25952);
nor U26342 (N_26342,N_24911,N_25015);
nand U26343 (N_26343,N_24877,N_25159);
xor U26344 (N_26344,N_24158,N_24258);
or U26345 (N_26345,N_25533,N_24791);
nand U26346 (N_26346,N_24415,N_24426);
and U26347 (N_26347,N_25916,N_25718);
nor U26348 (N_26348,N_25665,N_24773);
nand U26349 (N_26349,N_25888,N_25885);
xor U26350 (N_26350,N_25671,N_25956);
xor U26351 (N_26351,N_25230,N_25318);
or U26352 (N_26352,N_24103,N_24026);
or U26353 (N_26353,N_24185,N_25488);
and U26354 (N_26354,N_24915,N_25354);
and U26355 (N_26355,N_24490,N_24111);
xor U26356 (N_26356,N_25740,N_24296);
nand U26357 (N_26357,N_25100,N_24649);
or U26358 (N_26358,N_24545,N_25791);
nor U26359 (N_26359,N_25342,N_24681);
or U26360 (N_26360,N_25012,N_25441);
or U26361 (N_26361,N_24838,N_24724);
nand U26362 (N_26362,N_24277,N_24991);
or U26363 (N_26363,N_24859,N_25678);
xnor U26364 (N_26364,N_25285,N_24825);
nor U26365 (N_26365,N_24520,N_25232);
nor U26366 (N_26366,N_25431,N_25417);
or U26367 (N_26367,N_25775,N_25218);
and U26368 (N_26368,N_25824,N_25914);
or U26369 (N_26369,N_24920,N_24067);
xnor U26370 (N_26370,N_25004,N_24076);
xnor U26371 (N_26371,N_24897,N_24337);
nand U26372 (N_26372,N_24939,N_25743);
and U26373 (N_26373,N_25559,N_24770);
xnor U26374 (N_26374,N_24425,N_25786);
or U26375 (N_26375,N_24537,N_25138);
nand U26376 (N_26376,N_25470,N_25992);
nor U26377 (N_26377,N_25771,N_25747);
nand U26378 (N_26378,N_24713,N_25858);
or U26379 (N_26379,N_24031,N_25485);
or U26380 (N_26380,N_25466,N_25993);
nor U26381 (N_26381,N_25629,N_24449);
or U26382 (N_26382,N_24106,N_24140);
xor U26383 (N_26383,N_25449,N_25274);
nand U26384 (N_26384,N_25199,N_25519);
and U26385 (N_26385,N_25372,N_25158);
nand U26386 (N_26386,N_24980,N_24392);
nand U26387 (N_26387,N_25351,N_24314);
xor U26388 (N_26388,N_25077,N_25864);
or U26389 (N_26389,N_24308,N_24481);
or U26390 (N_26390,N_25089,N_24414);
and U26391 (N_26391,N_24124,N_24719);
or U26392 (N_26392,N_24865,N_24399);
nor U26393 (N_26393,N_25664,N_24502);
and U26394 (N_26394,N_24779,N_24976);
nand U26395 (N_26395,N_24451,N_25419);
nand U26396 (N_26396,N_24126,N_24369);
or U26397 (N_26397,N_25370,N_24182);
nand U26398 (N_26398,N_24579,N_25537);
xor U26399 (N_26399,N_25091,N_25269);
or U26400 (N_26400,N_25193,N_25202);
and U26401 (N_26401,N_25555,N_24248);
xor U26402 (N_26402,N_25899,N_24450);
or U26403 (N_26403,N_25082,N_24139);
nand U26404 (N_26404,N_25884,N_25978);
or U26405 (N_26405,N_25309,N_25972);
xnor U26406 (N_26406,N_25908,N_24669);
xor U26407 (N_26407,N_24280,N_24863);
or U26408 (N_26408,N_25296,N_24456);
xor U26409 (N_26409,N_24715,N_25594);
nand U26410 (N_26410,N_24630,N_25962);
nor U26411 (N_26411,N_25847,N_25852);
and U26412 (N_26412,N_24653,N_24150);
nor U26413 (N_26413,N_25166,N_25688);
or U26414 (N_26414,N_24699,N_25968);
nor U26415 (N_26415,N_24434,N_25681);
nand U26416 (N_26416,N_25072,N_24341);
or U26417 (N_26417,N_24065,N_25911);
nor U26418 (N_26418,N_24223,N_24488);
or U26419 (N_26419,N_24968,N_25240);
and U26420 (N_26420,N_25328,N_25769);
and U26421 (N_26421,N_25479,N_24529);
and U26422 (N_26422,N_24997,N_25680);
nand U26423 (N_26423,N_25860,N_25214);
and U26424 (N_26424,N_24403,N_25626);
nand U26425 (N_26425,N_25154,N_24036);
and U26426 (N_26426,N_24070,N_25721);
and U26427 (N_26427,N_25109,N_25987);
or U26428 (N_26428,N_24002,N_25807);
nor U26429 (N_26429,N_24217,N_25319);
nor U26430 (N_26430,N_25874,N_25112);
or U26431 (N_26431,N_25546,N_24238);
xor U26432 (N_26432,N_25245,N_25619);
nor U26433 (N_26433,N_25086,N_24339);
and U26434 (N_26434,N_25045,N_24293);
or U26435 (N_26435,N_25350,N_25983);
xor U26436 (N_26436,N_25247,N_25337);
or U26437 (N_26437,N_24926,N_24108);
nor U26438 (N_26438,N_25164,N_25595);
nor U26439 (N_26439,N_24060,N_24301);
nor U26440 (N_26440,N_25212,N_25763);
nor U26441 (N_26441,N_25919,N_24604);
nand U26442 (N_26442,N_25636,N_24014);
nand U26443 (N_26443,N_24222,N_25320);
xnor U26444 (N_26444,N_25139,N_25906);
xnor U26445 (N_26445,N_24607,N_25957);
or U26446 (N_26446,N_25332,N_24297);
and U26447 (N_26447,N_24113,N_24015);
or U26448 (N_26448,N_25152,N_24009);
and U26449 (N_26449,N_24727,N_24623);
and U26450 (N_26450,N_24179,N_25591);
nor U26451 (N_26451,N_24733,N_25867);
xnor U26452 (N_26452,N_25073,N_25943);
or U26453 (N_26453,N_24228,N_24599);
or U26454 (N_26454,N_25708,N_24597);
or U26455 (N_26455,N_25592,N_24100);
nor U26456 (N_26456,N_24062,N_24963);
or U26457 (N_26457,N_24227,N_25484);
nand U26458 (N_26458,N_24793,N_25617);
or U26459 (N_26459,N_24923,N_24588);
nand U26460 (N_26460,N_25661,N_24513);
and U26461 (N_26461,N_25772,N_25848);
nor U26462 (N_26462,N_24054,N_24122);
nand U26463 (N_26463,N_25525,N_24592);
and U26464 (N_26464,N_25965,N_24571);
nand U26465 (N_26465,N_25898,N_24841);
xnor U26466 (N_26466,N_25223,N_24463);
xor U26467 (N_26467,N_25621,N_24081);
nor U26468 (N_26468,N_24631,N_24635);
and U26469 (N_26469,N_24741,N_25424);
and U26470 (N_26470,N_24655,N_25125);
nor U26471 (N_26471,N_24129,N_24609);
nand U26472 (N_26472,N_24676,N_24274);
nand U26473 (N_26473,N_25966,N_24064);
nand U26474 (N_26474,N_24808,N_24107);
or U26475 (N_26475,N_24925,N_25608);
nor U26476 (N_26476,N_24726,N_25061);
nand U26477 (N_26477,N_24484,N_24697);
nor U26478 (N_26478,N_24311,N_25408);
and U26479 (N_26479,N_24884,N_25322);
and U26480 (N_26480,N_24600,N_24988);
or U26481 (N_26481,N_25374,N_25492);
and U26482 (N_26482,N_25448,N_25809);
or U26483 (N_26483,N_24099,N_25203);
nand U26484 (N_26484,N_25067,N_25410);
xor U26485 (N_26485,N_25751,N_24098);
or U26486 (N_26486,N_24763,N_25971);
and U26487 (N_26487,N_24402,N_25059);
and U26488 (N_26488,N_24278,N_24814);
nor U26489 (N_26489,N_25843,N_24379);
and U26490 (N_26490,N_25065,N_25444);
nand U26491 (N_26491,N_25921,N_25458);
and U26492 (N_26492,N_24382,N_24852);
nor U26493 (N_26493,N_25439,N_25467);
nor U26494 (N_26494,N_24577,N_24616);
nand U26495 (N_26495,N_25990,N_24700);
nand U26496 (N_26496,N_25105,N_25927);
or U26497 (N_26497,N_24424,N_24788);
xnor U26498 (N_26498,N_24466,N_25483);
nand U26499 (N_26499,N_25425,N_24034);
and U26500 (N_26500,N_24698,N_24443);
nand U26501 (N_26501,N_25936,N_24196);
and U26502 (N_26502,N_25907,N_24006);
nor U26503 (N_26503,N_24023,N_25020);
or U26504 (N_26504,N_25133,N_24893);
or U26505 (N_26505,N_24750,N_25130);
nor U26506 (N_26506,N_24397,N_24398);
and U26507 (N_26507,N_24180,N_24875);
or U26508 (N_26508,N_24347,N_25871);
nor U26509 (N_26509,N_24986,N_25655);
or U26510 (N_26510,N_24610,N_24042);
and U26511 (N_26511,N_25991,N_25816);
or U26512 (N_26512,N_25738,N_25880);
and U26513 (N_26513,N_25486,N_24683);
nor U26514 (N_26514,N_25104,N_25092);
nand U26515 (N_26515,N_25767,N_25788);
and U26516 (N_26516,N_24170,N_24772);
xor U26517 (N_26517,N_24226,N_24795);
nor U26518 (N_26518,N_24203,N_24973);
xor U26519 (N_26519,N_24161,N_24831);
or U26520 (N_26520,N_25753,N_25380);
nor U26521 (N_26521,N_25601,N_24854);
and U26522 (N_26522,N_25958,N_25401);
or U26523 (N_26523,N_24496,N_24794);
xnor U26524 (N_26524,N_24115,N_25224);
nor U26525 (N_26525,N_25583,N_25177);
nor U26526 (N_26526,N_25079,N_24147);
and U26527 (N_26527,N_25007,N_25280);
or U26528 (N_26528,N_25535,N_24890);
nand U26529 (N_26529,N_25122,N_24327);
and U26530 (N_26530,N_25819,N_25922);
or U26531 (N_26531,N_24866,N_24028);
or U26532 (N_26532,N_24404,N_24654);
nand U26533 (N_26533,N_25377,N_25368);
xor U26534 (N_26534,N_24704,N_24055);
or U26535 (N_26535,N_25675,N_24786);
nand U26536 (N_26536,N_25442,N_25758);
nor U26537 (N_26537,N_24743,N_25810);
nor U26538 (N_26538,N_24497,N_24384);
xor U26539 (N_26539,N_24279,N_24330);
xor U26540 (N_26540,N_25982,N_25599);
or U26541 (N_26541,N_24145,N_24864);
nor U26542 (N_26542,N_24810,N_24372);
and U26543 (N_26543,N_25365,N_25366);
or U26544 (N_26544,N_25361,N_24454);
nand U26545 (N_26545,N_24544,N_25955);
xor U26546 (N_26546,N_25162,N_25183);
nand U26547 (N_26547,N_25828,N_24285);
nor U26548 (N_26548,N_25612,N_25961);
nor U26549 (N_26549,N_24505,N_25475);
nor U26550 (N_26550,N_24620,N_25986);
nor U26551 (N_26551,N_25823,N_24567);
xor U26552 (N_26552,N_24527,N_24001);
nor U26553 (N_26553,N_24220,N_24186);
xnor U26554 (N_26554,N_25371,N_24575);
xnor U26555 (N_26555,N_24933,N_25584);
nand U26556 (N_26556,N_24818,N_24422);
or U26557 (N_26557,N_25463,N_24148);
nor U26558 (N_26558,N_24317,N_25576);
nand U26559 (N_26559,N_25465,N_24127);
and U26560 (N_26560,N_24714,N_24551);
or U26561 (N_26561,N_25672,N_24232);
xnor U26562 (N_26562,N_24073,N_25938);
nand U26563 (N_26563,N_24370,N_24629);
xnor U26564 (N_26564,N_24621,N_24197);
nor U26565 (N_26565,N_24017,N_25039);
or U26566 (N_26566,N_24178,N_25727);
or U26567 (N_26567,N_24815,N_25265);
nand U26568 (N_26568,N_24472,N_25036);
and U26569 (N_26569,N_24032,N_24413);
nor U26570 (N_26570,N_24195,N_24594);
or U26571 (N_26571,N_25390,N_24230);
and U26572 (N_26572,N_25326,N_25790);
nor U26573 (N_26573,N_24789,N_24249);
nand U26574 (N_26574,N_25167,N_24889);
or U26575 (N_26575,N_24389,N_25856);
nor U26576 (N_26576,N_25403,N_24048);
or U26577 (N_26577,N_25282,N_25324);
and U26578 (N_26578,N_25950,N_25103);
nor U26579 (N_26579,N_25384,N_25660);
xor U26580 (N_26580,N_24137,N_25745);
nor U26581 (N_26581,N_24639,N_24442);
xor U26582 (N_26582,N_25455,N_24154);
xnor U26583 (N_26583,N_25759,N_24420);
nor U26584 (N_26584,N_24040,N_25459);
nor U26585 (N_26585,N_25855,N_24247);
nand U26586 (N_26586,N_25684,N_25438);
xnor U26587 (N_26587,N_24857,N_24192);
nor U26588 (N_26588,N_25615,N_25238);
and U26589 (N_26589,N_24242,N_24518);
or U26590 (N_26590,N_24615,N_24043);
and U26591 (N_26591,N_25502,N_25244);
xnor U26592 (N_26592,N_25528,N_24847);
xor U26593 (N_26593,N_24068,N_24626);
nor U26594 (N_26594,N_25698,N_24842);
or U26595 (N_26595,N_25284,N_24661);
and U26596 (N_26596,N_25882,N_25877);
xnor U26597 (N_26597,N_25869,N_24335);
nor U26598 (N_26598,N_24918,N_24029);
nand U26599 (N_26599,N_25341,N_24981);
nand U26600 (N_26600,N_24542,N_25124);
nor U26601 (N_26601,N_25445,N_24771);
nor U26602 (N_26602,N_25785,N_24155);
and U26603 (N_26603,N_25742,N_25153);
and U26604 (N_26604,N_25624,N_24942);
and U26605 (N_26605,N_24495,N_24598);
nor U26606 (N_26606,N_24516,N_24487);
xnor U26607 (N_26607,N_25649,N_24509);
nor U26608 (N_26608,N_25418,N_25227);
nor U26609 (N_26609,N_24962,N_24510);
xor U26610 (N_26610,N_25179,N_25932);
nand U26611 (N_26611,N_25562,N_24160);
and U26612 (N_26612,N_25381,N_24619);
xor U26613 (N_26613,N_24149,N_24548);
or U26614 (N_26614,N_24627,N_25674);
xor U26615 (N_26615,N_25532,N_24354);
or U26616 (N_26616,N_25306,N_24381);
nand U26617 (N_26617,N_25507,N_25813);
and U26618 (N_26618,N_24209,N_24066);
nor U26619 (N_26619,N_25331,N_24904);
nand U26620 (N_26620,N_24486,N_24316);
nor U26621 (N_26621,N_25094,N_24408);
nor U26622 (N_26622,N_25611,N_25964);
and U26623 (N_26623,N_24947,N_24711);
nor U26624 (N_26624,N_24587,N_24493);
or U26625 (N_26625,N_25818,N_25271);
and U26626 (N_26626,N_24069,N_24672);
and U26627 (N_26627,N_25327,N_25060);
or U26628 (N_26628,N_25534,N_25667);
or U26629 (N_26629,N_24586,N_25129);
and U26630 (N_26630,N_24614,N_25420);
or U26631 (N_26631,N_24368,N_25709);
nand U26632 (N_26632,N_25187,N_24409);
nor U26633 (N_26633,N_24320,N_25789);
and U26634 (N_26634,N_25333,N_24881);
nor U26635 (N_26635,N_25640,N_24202);
or U26636 (N_26636,N_25170,N_24194);
or U26637 (N_26637,N_24869,N_24325);
and U26638 (N_26638,N_25147,N_24625);
and U26639 (N_26639,N_25541,N_25582);
or U26640 (N_26640,N_25547,N_24174);
xnor U26641 (N_26641,N_25252,N_25923);
or U26642 (N_26642,N_25731,N_25501);
nand U26643 (N_26643,N_25977,N_24970);
nand U26644 (N_26644,N_24303,N_24300);
or U26645 (N_26645,N_24912,N_25568);
nor U26646 (N_26646,N_25305,N_24856);
xor U26647 (N_26647,N_24471,N_25185);
or U26648 (N_26648,N_25078,N_25580);
xnor U26649 (N_26649,N_24164,N_25140);
xor U26650 (N_26650,N_25278,N_25256);
xor U26651 (N_26651,N_24780,N_25422);
nand U26652 (N_26652,N_25732,N_24560);
nor U26653 (N_26653,N_24319,N_24931);
or U26654 (N_26654,N_24729,N_25155);
xor U26655 (N_26655,N_25234,N_25353);
or U26656 (N_26656,N_25891,N_24742);
and U26657 (N_26657,N_24532,N_24645);
xor U26658 (N_26658,N_25543,N_24333);
nand U26659 (N_26659,N_24039,N_24685);
nor U26660 (N_26660,N_24637,N_25497);
or U26661 (N_26661,N_24983,N_25707);
nand U26662 (N_26662,N_25777,N_24692);
or U26663 (N_26663,N_24910,N_25799);
nand U26664 (N_26664,N_25711,N_25241);
or U26665 (N_26665,N_25364,N_24728);
or U26666 (N_26666,N_24225,N_25034);
and U26667 (N_26667,N_24266,N_24874);
and U26668 (N_26668,N_24951,N_24735);
nor U26669 (N_26669,N_24008,N_24907);
or U26670 (N_26670,N_24646,N_25719);
nor U26671 (N_26671,N_24596,N_24343);
nor U26672 (N_26672,N_24648,N_24128);
or U26673 (N_26673,N_24130,N_24452);
nand U26674 (N_26674,N_25473,N_24323);
xor U26675 (N_26675,N_25474,N_25254);
or U26676 (N_26676,N_24363,N_25148);
xor U26677 (N_26677,N_25106,N_25831);
nand U26678 (N_26678,N_24508,N_25893);
xor U26679 (N_26679,N_24512,N_25638);
nor U26680 (N_26680,N_25653,N_25716);
nor U26681 (N_26681,N_24633,N_25575);
xor U26682 (N_26682,N_25196,N_24143);
nand U26683 (N_26683,N_24298,N_25650);
nor U26684 (N_26684,N_24566,N_24641);
xnor U26685 (N_26685,N_24589,N_24385);
or U26686 (N_26686,N_25013,N_25564);
nor U26687 (N_26687,N_24929,N_25654);
nand U26688 (N_26688,N_25211,N_24636);
and U26689 (N_26689,N_24675,N_24050);
or U26690 (N_26690,N_24834,N_24005);
nor U26691 (N_26691,N_25222,N_25083);
and U26692 (N_26692,N_25314,N_25524);
nor U26693 (N_26693,N_25979,N_25242);
or U26694 (N_26694,N_25226,N_25160);
nor U26695 (N_26695,N_25635,N_24932);
or U26696 (N_26696,N_24492,N_24377);
or U26697 (N_26697,N_24224,N_24783);
nand U26698 (N_26698,N_25812,N_25704);
and U26699 (N_26699,N_25048,N_25508);
and U26700 (N_26700,N_25464,N_25598);
and U26701 (N_26701,N_24967,N_24761);
nor U26702 (N_26702,N_25286,N_25135);
xor U26703 (N_26703,N_24844,N_25250);
or U26704 (N_26704,N_24183,N_25329);
nor U26705 (N_26705,N_25623,N_24243);
or U26706 (N_26706,N_25641,N_24827);
nand U26707 (N_26707,N_25165,N_24412);
xnor U26708 (N_26708,N_25210,N_25128);
xor U26709 (N_26709,N_25794,N_25217);
or U26710 (N_26710,N_25261,N_24427);
or U26711 (N_26711,N_25760,N_25359);
xor U26712 (N_26712,N_25243,N_25095);
or U26713 (N_26713,N_24349,N_25821);
or U26714 (N_26714,N_25205,N_25063);
xnor U26715 (N_26715,N_25110,N_25136);
nor U26716 (N_26716,N_25490,N_24908);
nor U26717 (N_26717,N_25750,N_24380);
nand U26718 (N_26718,N_24674,N_25487);
xor U26719 (N_26719,N_25456,N_25468);
and U26720 (N_26720,N_24373,N_25186);
xnor U26721 (N_26721,N_24887,N_25798);
nand U26722 (N_26722,N_24899,N_25118);
and U26723 (N_26723,N_24461,N_25820);
nor U26724 (N_26724,N_25171,N_24740);
xnor U26725 (N_26725,N_25604,N_24144);
xor U26726 (N_26726,N_25832,N_24116);
nor U26727 (N_26727,N_24364,N_24955);
nor U26728 (N_26728,N_24201,N_25288);
or U26729 (N_26729,N_24181,N_25264);
nand U26730 (N_26730,N_25690,N_24166);
and U26731 (N_26731,N_24215,N_24647);
nor U26732 (N_26732,N_24668,N_25929);
and U26733 (N_26733,N_24538,N_24767);
nand U26734 (N_26734,N_25028,N_25258);
or U26735 (N_26735,N_25450,N_25504);
nand U26736 (N_26736,N_25093,N_25301);
or U26737 (N_26737,N_25197,N_24359);
nand U26738 (N_26738,N_25339,N_24919);
nand U26739 (N_26739,N_24805,N_25778);
nor U26740 (N_26740,N_25516,N_25808);
nor U26741 (N_26741,N_24632,N_24131);
and U26742 (N_26742,N_25041,N_24417);
and U26743 (N_26743,N_25712,N_25839);
xnor U26744 (N_26744,N_24090,N_24849);
nor U26745 (N_26745,N_24605,N_24141);
nor U26746 (N_26746,N_25651,N_24251);
and U26747 (N_26747,N_24169,N_24480);
nor U26748 (N_26748,N_25949,N_25412);
nand U26749 (N_26749,N_24689,N_24777);
nor U26750 (N_26750,N_25603,N_25552);
xnor U26751 (N_26751,N_24664,N_24310);
and U26752 (N_26752,N_24405,N_25796);
xnor U26753 (N_26753,N_24383,N_25206);
or U26754 (N_26754,N_25397,N_24618);
nor U26755 (N_26755,N_24229,N_25495);
and U26756 (N_26756,N_25434,N_24800);
nor U26757 (N_26757,N_24937,N_25550);
or U26758 (N_26758,N_25176,N_24306);
and U26759 (N_26759,N_24737,N_24985);
xnor U26760 (N_26760,N_25307,N_25779);
and U26761 (N_26761,N_24305,N_24000);
or U26762 (N_26762,N_24395,N_25702);
nand U26763 (N_26763,N_24593,N_24803);
and U26764 (N_26764,N_24826,N_24717);
xor U26765 (N_26765,N_25686,N_25628);
and U26766 (N_26766,N_25696,N_25070);
xnor U26767 (N_26767,N_25027,N_25311);
nor U26768 (N_26768,N_24853,N_24117);
xnor U26769 (N_26769,N_24212,N_25024);
nand U26770 (N_26770,N_24190,N_25143);
or U26771 (N_26771,N_25739,N_25896);
nor U26772 (N_26772,N_25498,N_24930);
xor U26773 (N_26773,N_24393,N_25255);
nor U26774 (N_26774,N_24216,N_25216);
xnor U26775 (N_26775,N_25219,N_25407);
nand U26776 (N_26776,N_24253,N_24265);
nand U26777 (N_26777,N_24662,N_25627);
and U26778 (N_26778,N_25913,N_25220);
nand U26779 (N_26779,N_24989,N_25348);
or U26780 (N_26780,N_25725,N_24156);
or U26781 (N_26781,N_25728,N_25648);
and U26782 (N_26782,N_24307,N_25976);
and U26783 (N_26783,N_24798,N_25586);
or U26784 (N_26784,N_25121,N_25029);
or U26785 (N_26785,N_24895,N_24396);
nand U26786 (N_26786,N_25005,N_24721);
and U26787 (N_26787,N_25652,N_24421);
or U26788 (N_26788,N_24694,N_24304);
and U26789 (N_26789,N_24092,N_24892);
and U26790 (N_26790,N_24468,N_24153);
nand U26791 (N_26791,N_24061,N_25101);
nor U26792 (N_26792,N_24943,N_24458);
nand U26793 (N_26793,N_24696,N_24302);
or U26794 (N_26794,N_24873,N_25695);
xnor U26795 (N_26795,N_25426,N_24562);
nor U26796 (N_26796,N_25042,N_25838);
nor U26797 (N_26797,N_24953,N_24756);
xnor U26798 (N_26798,N_24334,N_25781);
xnor U26799 (N_26799,N_24554,N_25774);
and U26800 (N_26800,N_25761,N_25416);
or U26801 (N_26801,N_24444,N_24356);
and U26802 (N_26802,N_24291,N_25614);
nand U26803 (N_26803,N_24257,N_24703);
or U26804 (N_26804,N_24561,N_25478);
xnor U26805 (N_26805,N_25996,N_24667);
or U26806 (N_26806,N_24049,N_25683);
and U26807 (N_26807,N_24522,N_24119);
and U26808 (N_26808,N_25521,N_25291);
nand U26809 (N_26809,N_25146,N_25358);
nor U26810 (N_26810,N_24642,N_25405);
nand U26811 (N_26811,N_25975,N_25016);
or U26812 (N_26812,N_25942,N_25496);
nand U26813 (N_26813,N_25764,N_24958);
nand U26814 (N_26814,N_25325,N_25881);
nand U26815 (N_26815,N_24011,N_24172);
xor U26816 (N_26816,N_25825,N_24286);
and U26817 (N_26817,N_25277,N_25632);
xnor U26818 (N_26818,N_24125,N_25260);
or U26819 (N_26819,N_24138,N_24440);
and U26820 (N_26820,N_24913,N_25414);
or U26821 (N_26821,N_24921,N_25940);
nand U26822 (N_26822,N_25347,N_25023);
or U26823 (N_26823,N_24132,N_24747);
xnor U26824 (N_26824,N_25517,N_24606);
nand U26825 (N_26825,N_24056,N_25685);
and U26826 (N_26826,N_24240,N_24785);
nor U26827 (N_26827,N_25399,N_25317);
nor U26828 (N_26828,N_24342,N_25266);
nor U26829 (N_26829,N_24723,N_24531);
nor U26830 (N_26830,N_24446,N_24467);
or U26831 (N_26831,N_25842,N_25108);
xor U26832 (N_26832,N_24523,N_24739);
or U26833 (N_26833,N_25299,N_24507);
nor U26834 (N_26834,N_24436,N_25868);
and U26835 (N_26835,N_24211,N_24839);
xnor U26836 (N_26836,N_25194,N_24652);
nand U26837 (N_26837,N_24263,N_25340);
nand U26838 (N_26838,N_24553,N_24273);
nor U26839 (N_26839,N_25003,N_25523);
nand U26840 (N_26840,N_25482,N_24867);
and U26841 (N_26841,N_24350,N_25111);
or U26842 (N_26842,N_25085,N_25757);
nor U26843 (N_26843,N_24823,N_24754);
xor U26844 (N_26844,N_24210,N_24687);
xor U26845 (N_26845,N_24033,N_25113);
and U26846 (N_26846,N_25762,N_24524);
and U26847 (N_26847,N_24406,N_25181);
and U26848 (N_26848,N_25267,N_25933);
and U26849 (N_26849,N_24804,N_25726);
nor U26850 (N_26850,N_24569,N_25644);
nand U26851 (N_26851,N_24720,N_25275);
and U26852 (N_26852,N_24019,N_25587);
and U26853 (N_26853,N_24738,N_24345);
xnor U26854 (N_26854,N_24214,N_24312);
or U26855 (N_26855,N_25746,N_25297);
xnor U26856 (N_26856,N_24707,N_24245);
or U26857 (N_26857,N_24208,N_24437);
xor U26858 (N_26858,N_25755,N_25321);
nand U26859 (N_26859,N_25931,N_24275);
nor U26860 (N_26860,N_25844,N_24640);
nor U26861 (N_26861,N_24870,N_25904);
and U26862 (N_26862,N_24089,N_25631);
nand U26863 (N_26863,N_25263,N_25338);
xnor U26864 (N_26864,N_25531,N_25827);
nand U26865 (N_26865,N_25857,N_25385);
xnor U26866 (N_26866,N_25736,N_24896);
or U26867 (N_26867,N_25204,N_24732);
and U26868 (N_26868,N_25897,N_25025);
and U26869 (N_26869,N_25150,N_24135);
xor U26870 (N_26870,N_25262,N_24206);
and U26871 (N_26871,N_25596,N_25215);
and U26872 (N_26872,N_24013,N_25766);
or U26873 (N_26873,N_24428,N_24321);
or U26874 (N_26874,N_25191,N_24474);
nand U26875 (N_26875,N_24882,N_25427);
or U26876 (N_26876,N_24157,N_24558);
nand U26877 (N_26877,N_25283,N_25544);
or U26878 (N_26878,N_24974,N_25692);
nand U26879 (N_26879,N_25292,N_25713);
nor U26880 (N_26880,N_24045,N_24112);
and U26881 (N_26881,N_24260,N_25930);
nor U26882 (N_26882,N_24832,N_24764);
nand U26883 (N_26883,N_24097,N_25560);
and U26884 (N_26884,N_24611,N_24550);
xnor U26885 (N_26885,N_25526,N_25049);
or U26886 (N_26886,N_24924,N_25905);
xnor U26887 (N_26887,N_24165,N_24010);
or U26888 (N_26888,N_24746,N_25493);
or U26889 (N_26889,N_25840,N_24971);
xor U26890 (N_26890,N_25044,N_25369);
xor U26891 (N_26891,N_25581,N_24965);
nor U26892 (N_26892,N_25851,N_24549);
and U26893 (N_26893,N_25169,N_24037);
nor U26894 (N_26894,N_24244,N_24360);
nor U26895 (N_26895,N_24294,N_24189);
or U26896 (N_26896,N_24949,N_24946);
or U26897 (N_26897,N_25344,N_24219);
nand U26898 (N_26898,N_25117,N_24271);
nand U26899 (N_26899,N_25120,N_25471);
nand U26900 (N_26900,N_24716,N_24914);
or U26901 (N_26901,N_25075,N_24905);
xor U26902 (N_26902,N_24855,N_24879);
and U26903 (N_26903,N_25494,N_24358);
or U26904 (N_26904,N_24479,N_25935);
or U26905 (N_26905,N_24563,N_24813);
xor U26906 (N_26906,N_24725,N_24447);
xor U26907 (N_26907,N_24656,N_24079);
nand U26908 (N_26908,N_24004,N_25829);
and U26909 (N_26909,N_25336,N_25900);
xnor U26910 (N_26910,N_24533,N_24688);
xor U26911 (N_26911,N_24684,N_24121);
xor U26912 (N_26912,N_24168,N_25700);
nand U26913 (N_26913,N_24665,N_25116);
nand U26914 (N_26914,N_25647,N_25279);
xnor U26915 (N_26915,N_24917,N_24603);
xnor U26916 (N_26916,N_25235,N_24894);
and U26917 (N_26917,N_24830,N_25175);
nand U26918 (N_26918,N_25822,N_24543);
and U26919 (N_26919,N_24936,N_24710);
xnor U26920 (N_26920,N_24233,N_25273);
nand U26921 (N_26921,N_24806,N_24768);
nand U26922 (N_26922,N_25814,N_24702);
nor U26923 (N_26923,N_24329,N_24657);
xor U26924 (N_26924,N_24956,N_25846);
or U26925 (N_26925,N_25430,N_25051);
xnor U26926 (N_26926,N_25057,N_25657);
nor U26927 (N_26927,N_24671,N_24902);
xnor U26928 (N_26928,N_24328,N_25997);
nor U26929 (N_26929,N_24663,N_24465);
or U26930 (N_26930,N_24515,N_25787);
xnor U26931 (N_26931,N_25548,N_25951);
and U26932 (N_26932,N_25295,N_24591);
xnor U26933 (N_26933,N_25090,N_24961);
or U26934 (N_26934,N_24528,N_25076);
and U26935 (N_26935,N_25954,N_25443);
or U26936 (N_26936,N_24284,N_24199);
nand U26937 (N_26937,N_25928,N_24340);
nor U26938 (N_26938,N_24574,N_24016);
nor U26939 (N_26939,N_25646,N_24110);
and U26940 (N_26940,N_25460,N_25613);
nor U26941 (N_26941,N_24954,N_25330);
nand U26942 (N_26942,N_25863,N_25433);
or U26943 (N_26943,N_25001,N_25127);
nand U26944 (N_26944,N_25974,N_24057);
or U26945 (N_26945,N_24752,N_25411);
xnor U26946 (N_26946,N_24969,N_25047);
nor U26947 (N_26947,N_25999,N_25776);
or U26948 (N_26948,N_24205,N_25184);
nand U26949 (N_26949,N_25687,N_25744);
and U26950 (N_26950,N_25571,N_24850);
nand U26951 (N_26951,N_25081,N_25890);
or U26952 (N_26952,N_25386,N_24184);
and U26953 (N_26953,N_25303,N_24613);
and U26954 (N_26954,N_24706,N_25173);
nor U26955 (N_26955,N_25783,N_24176);
xnor U26956 (N_26956,N_24007,N_24812);
xnor U26957 (N_26957,N_24643,N_24511);
nand U26958 (N_26958,N_24934,N_25099);
or U26959 (N_26959,N_25959,N_25052);
xnor U26960 (N_26960,N_25835,N_24585);
or U26961 (N_26961,N_24555,N_24410);
or U26962 (N_26962,N_24071,N_25225);
nand U26963 (N_26963,N_25451,N_25395);
nand U26964 (N_26964,N_24473,N_25901);
and U26965 (N_26965,N_24996,N_25469);
nand U26966 (N_26966,N_25019,N_24478);
xnor U26967 (N_26967,N_24952,N_25021);
and U26968 (N_26968,N_24978,N_24693);
xor U26969 (N_26969,N_24475,N_25953);
xnor U26970 (N_26970,N_25102,N_25937);
and U26971 (N_26971,N_24748,N_24044);
or U26972 (N_26972,N_24972,N_25682);
xnor U26973 (N_26973,N_25833,N_24459);
xnor U26974 (N_26974,N_24348,N_24445);
nand U26975 (N_26975,N_25144,N_25428);
nand U26976 (N_26976,N_25770,N_25190);
or U26977 (N_26977,N_25367,N_25946);
nand U26978 (N_26978,N_25723,N_24012);
or U26979 (N_26979,N_24843,N_24101);
xnor U26980 (N_26980,N_24239,N_25679);
nand U26981 (N_26981,N_25886,N_25315);
and U26982 (N_26982,N_24775,N_25720);
nand U26983 (N_26983,N_25554,N_24018);
and U26984 (N_26984,N_24270,N_25563);
and U26985 (N_26985,N_24760,N_25536);
nor U26986 (N_26986,N_25415,N_25149);
xor U26987 (N_26987,N_24082,N_25676);
and U26988 (N_26988,N_24608,N_25572);
nor U26989 (N_26989,N_24162,N_25141);
nor U26990 (N_26990,N_25182,N_24658);
nor U26991 (N_26991,N_25765,N_25895);
nand U26992 (N_26992,N_24501,N_25797);
nor U26993 (N_26993,N_24102,N_24691);
or U26994 (N_26994,N_24500,N_24336);
or U26995 (N_26995,N_24313,N_25642);
xnor U26996 (N_26996,N_24901,N_25276);
or U26997 (N_26997,N_25452,N_25805);
and U26998 (N_26998,N_24821,N_25673);
nand U26999 (N_26999,N_24871,N_24499);
xnor U27000 (N_27000,N_24088,N_25796);
nor U27001 (N_27001,N_24688,N_25135);
nor U27002 (N_27002,N_25213,N_25708);
and U27003 (N_27003,N_25087,N_24501);
and U27004 (N_27004,N_25809,N_24114);
and U27005 (N_27005,N_25421,N_24696);
and U27006 (N_27006,N_25986,N_25635);
or U27007 (N_27007,N_25883,N_25440);
or U27008 (N_27008,N_25389,N_24856);
nand U27009 (N_27009,N_24620,N_25813);
xor U27010 (N_27010,N_25723,N_24740);
xnor U27011 (N_27011,N_24373,N_24844);
or U27012 (N_27012,N_24904,N_25590);
nor U27013 (N_27013,N_24827,N_24461);
xnor U27014 (N_27014,N_25874,N_25492);
and U27015 (N_27015,N_24898,N_25188);
xnor U27016 (N_27016,N_24968,N_25013);
xnor U27017 (N_27017,N_24474,N_24313);
xnor U27018 (N_27018,N_24130,N_25316);
and U27019 (N_27019,N_25836,N_24723);
nor U27020 (N_27020,N_24154,N_25016);
nand U27021 (N_27021,N_25125,N_25737);
or U27022 (N_27022,N_25833,N_25323);
nand U27023 (N_27023,N_25251,N_24648);
xnor U27024 (N_27024,N_24692,N_25648);
nor U27025 (N_27025,N_24940,N_25441);
and U27026 (N_27026,N_25021,N_24445);
nand U27027 (N_27027,N_25394,N_24066);
xnor U27028 (N_27028,N_25736,N_24395);
nor U27029 (N_27029,N_24204,N_24303);
nand U27030 (N_27030,N_25090,N_25010);
or U27031 (N_27031,N_25572,N_24941);
and U27032 (N_27032,N_24845,N_24320);
xnor U27033 (N_27033,N_25779,N_24543);
or U27034 (N_27034,N_24257,N_24212);
or U27035 (N_27035,N_24741,N_25144);
and U27036 (N_27036,N_24096,N_24442);
or U27037 (N_27037,N_24052,N_24396);
xor U27038 (N_27038,N_24403,N_24779);
and U27039 (N_27039,N_24932,N_25007);
and U27040 (N_27040,N_24535,N_24033);
and U27041 (N_27041,N_24794,N_25661);
or U27042 (N_27042,N_24369,N_25826);
and U27043 (N_27043,N_24089,N_25657);
and U27044 (N_27044,N_24513,N_25187);
and U27045 (N_27045,N_24955,N_24123);
or U27046 (N_27046,N_24371,N_24899);
xor U27047 (N_27047,N_24790,N_24310);
or U27048 (N_27048,N_25063,N_24915);
or U27049 (N_27049,N_25812,N_25548);
and U27050 (N_27050,N_25406,N_24844);
and U27051 (N_27051,N_25433,N_25353);
nor U27052 (N_27052,N_25792,N_25922);
xnor U27053 (N_27053,N_25560,N_24176);
xnor U27054 (N_27054,N_25808,N_24835);
and U27055 (N_27055,N_24319,N_25400);
xnor U27056 (N_27056,N_24861,N_24909);
or U27057 (N_27057,N_25481,N_25712);
nand U27058 (N_27058,N_25440,N_25280);
or U27059 (N_27059,N_25915,N_25438);
xor U27060 (N_27060,N_24899,N_25668);
xnor U27061 (N_27061,N_24882,N_25140);
or U27062 (N_27062,N_24860,N_24182);
or U27063 (N_27063,N_25460,N_25425);
nor U27064 (N_27064,N_24740,N_25038);
nand U27065 (N_27065,N_25965,N_24659);
or U27066 (N_27066,N_25482,N_24700);
nor U27067 (N_27067,N_25673,N_25116);
xor U27068 (N_27068,N_24980,N_25598);
or U27069 (N_27069,N_25281,N_25292);
xor U27070 (N_27070,N_24933,N_24641);
nand U27071 (N_27071,N_24360,N_24987);
or U27072 (N_27072,N_24820,N_25812);
and U27073 (N_27073,N_25321,N_25872);
and U27074 (N_27074,N_24231,N_25129);
nand U27075 (N_27075,N_24860,N_25829);
nor U27076 (N_27076,N_24625,N_24955);
xor U27077 (N_27077,N_24567,N_25727);
and U27078 (N_27078,N_25014,N_25259);
and U27079 (N_27079,N_24208,N_25507);
nand U27080 (N_27080,N_25030,N_24575);
and U27081 (N_27081,N_24739,N_24018);
nor U27082 (N_27082,N_25653,N_25027);
nand U27083 (N_27083,N_25032,N_25475);
nor U27084 (N_27084,N_25858,N_25617);
xor U27085 (N_27085,N_24924,N_25349);
and U27086 (N_27086,N_24730,N_24993);
xor U27087 (N_27087,N_25486,N_25195);
nand U27088 (N_27088,N_25225,N_24722);
nor U27089 (N_27089,N_24255,N_25705);
nand U27090 (N_27090,N_25909,N_24426);
or U27091 (N_27091,N_25084,N_25660);
xor U27092 (N_27092,N_24428,N_25974);
nand U27093 (N_27093,N_25303,N_24366);
or U27094 (N_27094,N_24554,N_24606);
nand U27095 (N_27095,N_24216,N_24696);
xnor U27096 (N_27096,N_24219,N_25577);
nand U27097 (N_27097,N_24826,N_24757);
nor U27098 (N_27098,N_25161,N_24374);
or U27099 (N_27099,N_25269,N_24810);
nor U27100 (N_27100,N_24337,N_24847);
or U27101 (N_27101,N_25608,N_24555);
nand U27102 (N_27102,N_24723,N_24889);
and U27103 (N_27103,N_25409,N_25959);
and U27104 (N_27104,N_24017,N_24814);
nor U27105 (N_27105,N_25702,N_25494);
nand U27106 (N_27106,N_25774,N_24817);
and U27107 (N_27107,N_25048,N_24616);
xnor U27108 (N_27108,N_25877,N_25978);
xnor U27109 (N_27109,N_24424,N_24310);
and U27110 (N_27110,N_24527,N_24821);
nor U27111 (N_27111,N_25846,N_25722);
xor U27112 (N_27112,N_25778,N_24702);
and U27113 (N_27113,N_25665,N_25482);
or U27114 (N_27114,N_24200,N_25715);
xor U27115 (N_27115,N_25749,N_24040);
and U27116 (N_27116,N_25032,N_25472);
xor U27117 (N_27117,N_25985,N_24035);
xnor U27118 (N_27118,N_24458,N_25804);
nor U27119 (N_27119,N_24822,N_24477);
xnor U27120 (N_27120,N_25899,N_24621);
nand U27121 (N_27121,N_24557,N_24773);
or U27122 (N_27122,N_25420,N_24944);
nor U27123 (N_27123,N_25464,N_24604);
nor U27124 (N_27124,N_24103,N_24822);
nand U27125 (N_27125,N_24715,N_25876);
and U27126 (N_27126,N_24404,N_25833);
or U27127 (N_27127,N_25325,N_25638);
nand U27128 (N_27128,N_24567,N_24958);
or U27129 (N_27129,N_25610,N_24426);
xor U27130 (N_27130,N_24769,N_24651);
xor U27131 (N_27131,N_25344,N_25719);
and U27132 (N_27132,N_24027,N_24926);
and U27133 (N_27133,N_25852,N_25255);
or U27134 (N_27134,N_25113,N_25669);
nand U27135 (N_27135,N_25296,N_24176);
and U27136 (N_27136,N_24664,N_24382);
xnor U27137 (N_27137,N_24086,N_24013);
xor U27138 (N_27138,N_25140,N_25945);
or U27139 (N_27139,N_25231,N_24878);
or U27140 (N_27140,N_24815,N_24009);
xor U27141 (N_27141,N_24653,N_25887);
nor U27142 (N_27142,N_25035,N_24952);
nor U27143 (N_27143,N_24869,N_25183);
nand U27144 (N_27144,N_24663,N_25128);
or U27145 (N_27145,N_25532,N_25333);
xor U27146 (N_27146,N_24447,N_25126);
xor U27147 (N_27147,N_25404,N_25033);
xnor U27148 (N_27148,N_24143,N_24813);
or U27149 (N_27149,N_24025,N_24977);
xor U27150 (N_27150,N_25709,N_24674);
xnor U27151 (N_27151,N_25441,N_24915);
nor U27152 (N_27152,N_25208,N_25895);
or U27153 (N_27153,N_24199,N_24090);
xor U27154 (N_27154,N_24757,N_24515);
nand U27155 (N_27155,N_25050,N_24079);
xor U27156 (N_27156,N_25493,N_25705);
and U27157 (N_27157,N_24299,N_24090);
and U27158 (N_27158,N_25717,N_25090);
or U27159 (N_27159,N_24256,N_24910);
and U27160 (N_27160,N_25284,N_24232);
and U27161 (N_27161,N_25745,N_25974);
nand U27162 (N_27162,N_24327,N_24314);
or U27163 (N_27163,N_25284,N_25619);
and U27164 (N_27164,N_25610,N_25379);
or U27165 (N_27165,N_24399,N_24976);
or U27166 (N_27166,N_25549,N_25712);
and U27167 (N_27167,N_24513,N_24362);
xnor U27168 (N_27168,N_25129,N_24253);
nand U27169 (N_27169,N_24808,N_24368);
nor U27170 (N_27170,N_25294,N_25867);
xnor U27171 (N_27171,N_25114,N_25098);
nor U27172 (N_27172,N_25712,N_25339);
or U27173 (N_27173,N_24702,N_25891);
or U27174 (N_27174,N_24773,N_24750);
xnor U27175 (N_27175,N_24771,N_24368);
or U27176 (N_27176,N_24093,N_24531);
and U27177 (N_27177,N_25111,N_25284);
and U27178 (N_27178,N_25676,N_25855);
xor U27179 (N_27179,N_25227,N_25763);
nand U27180 (N_27180,N_25243,N_25553);
xnor U27181 (N_27181,N_25037,N_24294);
xnor U27182 (N_27182,N_24079,N_24190);
or U27183 (N_27183,N_25157,N_25040);
nand U27184 (N_27184,N_25431,N_24475);
xor U27185 (N_27185,N_24126,N_24816);
nor U27186 (N_27186,N_24951,N_24830);
nor U27187 (N_27187,N_25979,N_25894);
xnor U27188 (N_27188,N_24208,N_25608);
and U27189 (N_27189,N_25399,N_24883);
xor U27190 (N_27190,N_25426,N_25578);
and U27191 (N_27191,N_25675,N_25186);
nor U27192 (N_27192,N_24474,N_24364);
or U27193 (N_27193,N_25691,N_24204);
nor U27194 (N_27194,N_24065,N_24588);
and U27195 (N_27195,N_24139,N_24685);
nand U27196 (N_27196,N_24388,N_24885);
xnor U27197 (N_27197,N_25748,N_25087);
nor U27198 (N_27198,N_24828,N_24710);
or U27199 (N_27199,N_25355,N_24240);
or U27200 (N_27200,N_24995,N_25145);
xor U27201 (N_27201,N_25703,N_25142);
or U27202 (N_27202,N_25461,N_25925);
and U27203 (N_27203,N_24756,N_25675);
nand U27204 (N_27204,N_24593,N_25674);
nand U27205 (N_27205,N_24543,N_25186);
nand U27206 (N_27206,N_25457,N_24032);
and U27207 (N_27207,N_24098,N_24903);
and U27208 (N_27208,N_24581,N_24831);
nand U27209 (N_27209,N_24834,N_24335);
xnor U27210 (N_27210,N_24549,N_24447);
nand U27211 (N_27211,N_25804,N_25983);
nor U27212 (N_27212,N_24270,N_25046);
xor U27213 (N_27213,N_24617,N_24337);
xor U27214 (N_27214,N_25875,N_24868);
nand U27215 (N_27215,N_24309,N_25615);
or U27216 (N_27216,N_24914,N_24457);
or U27217 (N_27217,N_24331,N_24783);
nand U27218 (N_27218,N_25772,N_25829);
nor U27219 (N_27219,N_24730,N_25747);
or U27220 (N_27220,N_25899,N_24059);
xor U27221 (N_27221,N_25942,N_24567);
nor U27222 (N_27222,N_25337,N_25286);
nand U27223 (N_27223,N_25873,N_25335);
nand U27224 (N_27224,N_24969,N_25700);
nand U27225 (N_27225,N_25924,N_24165);
nand U27226 (N_27226,N_25331,N_24471);
or U27227 (N_27227,N_24716,N_24115);
nand U27228 (N_27228,N_25410,N_24380);
nor U27229 (N_27229,N_25072,N_24365);
or U27230 (N_27230,N_25295,N_25926);
nor U27231 (N_27231,N_25532,N_24710);
and U27232 (N_27232,N_25267,N_25386);
nor U27233 (N_27233,N_25145,N_25536);
nor U27234 (N_27234,N_24721,N_25923);
nand U27235 (N_27235,N_24108,N_24662);
and U27236 (N_27236,N_24155,N_25246);
and U27237 (N_27237,N_25989,N_25164);
or U27238 (N_27238,N_25550,N_25111);
or U27239 (N_27239,N_25908,N_24478);
xnor U27240 (N_27240,N_25682,N_24177);
and U27241 (N_27241,N_24541,N_25212);
and U27242 (N_27242,N_24750,N_25228);
or U27243 (N_27243,N_25118,N_25802);
or U27244 (N_27244,N_25413,N_25802);
nor U27245 (N_27245,N_24256,N_24856);
xnor U27246 (N_27246,N_25236,N_24562);
nor U27247 (N_27247,N_25765,N_25263);
or U27248 (N_27248,N_24172,N_24883);
or U27249 (N_27249,N_25469,N_24257);
or U27250 (N_27250,N_24532,N_25919);
xor U27251 (N_27251,N_24244,N_25941);
or U27252 (N_27252,N_24169,N_25402);
xor U27253 (N_27253,N_25589,N_24952);
nand U27254 (N_27254,N_25211,N_24682);
or U27255 (N_27255,N_25810,N_24676);
nor U27256 (N_27256,N_24213,N_24763);
nand U27257 (N_27257,N_24275,N_25044);
xnor U27258 (N_27258,N_24113,N_25988);
nor U27259 (N_27259,N_25723,N_25579);
nor U27260 (N_27260,N_25946,N_25783);
or U27261 (N_27261,N_25436,N_24855);
nand U27262 (N_27262,N_24941,N_25898);
and U27263 (N_27263,N_24470,N_24233);
nand U27264 (N_27264,N_24229,N_25580);
xnor U27265 (N_27265,N_24388,N_25424);
nand U27266 (N_27266,N_25760,N_25252);
and U27267 (N_27267,N_25753,N_25980);
nor U27268 (N_27268,N_24753,N_24534);
and U27269 (N_27269,N_24805,N_24537);
xnor U27270 (N_27270,N_24822,N_25646);
nor U27271 (N_27271,N_24822,N_24505);
and U27272 (N_27272,N_25918,N_25646);
nor U27273 (N_27273,N_24809,N_25996);
nor U27274 (N_27274,N_25662,N_25717);
and U27275 (N_27275,N_24351,N_25932);
nor U27276 (N_27276,N_24978,N_25384);
and U27277 (N_27277,N_25634,N_25831);
nor U27278 (N_27278,N_24551,N_25538);
or U27279 (N_27279,N_25071,N_25762);
xnor U27280 (N_27280,N_24027,N_25206);
xnor U27281 (N_27281,N_25783,N_24583);
or U27282 (N_27282,N_24384,N_25590);
nand U27283 (N_27283,N_25409,N_24642);
xnor U27284 (N_27284,N_24320,N_25406);
nor U27285 (N_27285,N_24139,N_25684);
or U27286 (N_27286,N_24140,N_24998);
or U27287 (N_27287,N_25427,N_24703);
xor U27288 (N_27288,N_25362,N_25532);
and U27289 (N_27289,N_25863,N_24450);
and U27290 (N_27290,N_25058,N_24283);
nor U27291 (N_27291,N_25860,N_24711);
nor U27292 (N_27292,N_25215,N_25653);
nor U27293 (N_27293,N_24863,N_25391);
or U27294 (N_27294,N_24047,N_25539);
or U27295 (N_27295,N_25881,N_24093);
nand U27296 (N_27296,N_25688,N_25262);
nor U27297 (N_27297,N_25924,N_24767);
or U27298 (N_27298,N_25832,N_25890);
xnor U27299 (N_27299,N_24109,N_24962);
nand U27300 (N_27300,N_24618,N_24179);
or U27301 (N_27301,N_24860,N_25957);
xor U27302 (N_27302,N_25128,N_24501);
xor U27303 (N_27303,N_24286,N_25419);
nor U27304 (N_27304,N_25159,N_24262);
nand U27305 (N_27305,N_25170,N_24599);
nand U27306 (N_27306,N_25696,N_25716);
or U27307 (N_27307,N_25758,N_24741);
and U27308 (N_27308,N_24594,N_25526);
and U27309 (N_27309,N_25236,N_24891);
or U27310 (N_27310,N_25937,N_25825);
nor U27311 (N_27311,N_24262,N_24647);
nor U27312 (N_27312,N_25623,N_25406);
and U27313 (N_27313,N_25766,N_25819);
xnor U27314 (N_27314,N_24887,N_24638);
xnor U27315 (N_27315,N_25460,N_25343);
nor U27316 (N_27316,N_25280,N_24795);
nor U27317 (N_27317,N_25446,N_24183);
nand U27318 (N_27318,N_25627,N_25933);
nand U27319 (N_27319,N_25692,N_25918);
and U27320 (N_27320,N_25172,N_24455);
nor U27321 (N_27321,N_24814,N_25086);
nand U27322 (N_27322,N_25762,N_24293);
nor U27323 (N_27323,N_25198,N_25439);
nand U27324 (N_27324,N_24498,N_25209);
or U27325 (N_27325,N_25174,N_24282);
xnor U27326 (N_27326,N_25124,N_24618);
xor U27327 (N_27327,N_24412,N_24490);
or U27328 (N_27328,N_24770,N_25058);
nand U27329 (N_27329,N_24647,N_25170);
and U27330 (N_27330,N_24279,N_24157);
and U27331 (N_27331,N_24874,N_24765);
or U27332 (N_27332,N_25568,N_25046);
or U27333 (N_27333,N_25782,N_24425);
and U27334 (N_27334,N_25253,N_24937);
and U27335 (N_27335,N_25166,N_25627);
and U27336 (N_27336,N_25679,N_24700);
nor U27337 (N_27337,N_24946,N_25365);
nor U27338 (N_27338,N_24671,N_24315);
nand U27339 (N_27339,N_25453,N_25636);
or U27340 (N_27340,N_24115,N_24407);
nand U27341 (N_27341,N_25546,N_25788);
nand U27342 (N_27342,N_25641,N_24068);
or U27343 (N_27343,N_25879,N_25434);
nand U27344 (N_27344,N_25190,N_24290);
nor U27345 (N_27345,N_24416,N_25469);
xor U27346 (N_27346,N_25471,N_25418);
nor U27347 (N_27347,N_25132,N_24479);
or U27348 (N_27348,N_25689,N_25028);
nor U27349 (N_27349,N_24194,N_24489);
nor U27350 (N_27350,N_24434,N_24140);
nand U27351 (N_27351,N_25343,N_25862);
nand U27352 (N_27352,N_25870,N_25107);
nand U27353 (N_27353,N_24486,N_25382);
xnor U27354 (N_27354,N_24440,N_25004);
or U27355 (N_27355,N_24654,N_24732);
or U27356 (N_27356,N_24803,N_25118);
or U27357 (N_27357,N_24662,N_24132);
nand U27358 (N_27358,N_25001,N_25258);
xnor U27359 (N_27359,N_25653,N_25328);
nor U27360 (N_27360,N_24236,N_25161);
nand U27361 (N_27361,N_25619,N_24067);
or U27362 (N_27362,N_25788,N_24520);
xor U27363 (N_27363,N_24738,N_24152);
nand U27364 (N_27364,N_25588,N_24169);
nor U27365 (N_27365,N_24106,N_24622);
nor U27366 (N_27366,N_24155,N_25650);
or U27367 (N_27367,N_24996,N_24896);
or U27368 (N_27368,N_24050,N_25102);
nand U27369 (N_27369,N_24033,N_25849);
or U27370 (N_27370,N_25459,N_25831);
or U27371 (N_27371,N_24265,N_24524);
and U27372 (N_27372,N_24635,N_25409);
or U27373 (N_27373,N_25117,N_24236);
nor U27374 (N_27374,N_25116,N_25572);
nor U27375 (N_27375,N_25119,N_24622);
nand U27376 (N_27376,N_24736,N_25072);
or U27377 (N_27377,N_24094,N_24088);
nor U27378 (N_27378,N_24862,N_25157);
or U27379 (N_27379,N_24582,N_24942);
nand U27380 (N_27380,N_25327,N_24610);
xor U27381 (N_27381,N_24784,N_24506);
or U27382 (N_27382,N_24563,N_24539);
xor U27383 (N_27383,N_25133,N_24786);
or U27384 (N_27384,N_24482,N_25984);
or U27385 (N_27385,N_24451,N_24537);
nor U27386 (N_27386,N_25606,N_25137);
and U27387 (N_27387,N_24690,N_24574);
or U27388 (N_27388,N_24566,N_25631);
and U27389 (N_27389,N_24109,N_24418);
and U27390 (N_27390,N_25887,N_24061);
nand U27391 (N_27391,N_25988,N_24901);
nand U27392 (N_27392,N_24390,N_25286);
or U27393 (N_27393,N_25519,N_24134);
nor U27394 (N_27394,N_25720,N_25885);
nand U27395 (N_27395,N_24520,N_24537);
nand U27396 (N_27396,N_25817,N_24351);
nor U27397 (N_27397,N_25378,N_25114);
or U27398 (N_27398,N_24085,N_24210);
nor U27399 (N_27399,N_25153,N_24534);
nand U27400 (N_27400,N_24447,N_24230);
and U27401 (N_27401,N_24685,N_25003);
xor U27402 (N_27402,N_24581,N_24587);
or U27403 (N_27403,N_25249,N_24688);
nand U27404 (N_27404,N_24817,N_25600);
or U27405 (N_27405,N_25833,N_24524);
xor U27406 (N_27406,N_24809,N_24896);
and U27407 (N_27407,N_24606,N_25333);
nor U27408 (N_27408,N_24877,N_25192);
and U27409 (N_27409,N_24335,N_25165);
xnor U27410 (N_27410,N_24370,N_24251);
or U27411 (N_27411,N_24842,N_25150);
nor U27412 (N_27412,N_25481,N_24084);
nor U27413 (N_27413,N_25572,N_25926);
nor U27414 (N_27414,N_25781,N_24302);
nor U27415 (N_27415,N_24718,N_24369);
xor U27416 (N_27416,N_24356,N_24776);
xnor U27417 (N_27417,N_24981,N_25064);
xor U27418 (N_27418,N_25275,N_24397);
xor U27419 (N_27419,N_24806,N_25240);
xor U27420 (N_27420,N_25238,N_25830);
and U27421 (N_27421,N_25350,N_25956);
nand U27422 (N_27422,N_25691,N_24218);
nand U27423 (N_27423,N_24315,N_25024);
or U27424 (N_27424,N_24210,N_25223);
or U27425 (N_27425,N_25907,N_25468);
xnor U27426 (N_27426,N_24948,N_24928);
xnor U27427 (N_27427,N_24699,N_25620);
and U27428 (N_27428,N_25769,N_25644);
xnor U27429 (N_27429,N_25627,N_25958);
xor U27430 (N_27430,N_24367,N_25827);
nor U27431 (N_27431,N_25788,N_25864);
nor U27432 (N_27432,N_24588,N_24468);
xnor U27433 (N_27433,N_24809,N_24138);
nor U27434 (N_27434,N_24737,N_25559);
nand U27435 (N_27435,N_25710,N_24480);
or U27436 (N_27436,N_25637,N_25461);
nor U27437 (N_27437,N_25666,N_24069);
xnor U27438 (N_27438,N_25683,N_24220);
nand U27439 (N_27439,N_25963,N_24435);
or U27440 (N_27440,N_24632,N_24682);
nand U27441 (N_27441,N_24549,N_25760);
xnor U27442 (N_27442,N_24955,N_25344);
xnor U27443 (N_27443,N_25216,N_25852);
xnor U27444 (N_27444,N_25070,N_24290);
nor U27445 (N_27445,N_25327,N_24732);
or U27446 (N_27446,N_24166,N_25843);
or U27447 (N_27447,N_24385,N_24606);
nor U27448 (N_27448,N_24346,N_24958);
and U27449 (N_27449,N_25380,N_24373);
or U27450 (N_27450,N_25433,N_24020);
and U27451 (N_27451,N_24351,N_25079);
and U27452 (N_27452,N_24280,N_25273);
or U27453 (N_27453,N_25516,N_24692);
nand U27454 (N_27454,N_24803,N_25619);
and U27455 (N_27455,N_24285,N_25465);
or U27456 (N_27456,N_25207,N_24736);
and U27457 (N_27457,N_24583,N_25736);
nand U27458 (N_27458,N_25224,N_24978);
nand U27459 (N_27459,N_25679,N_24317);
and U27460 (N_27460,N_25005,N_25616);
and U27461 (N_27461,N_25323,N_25620);
nand U27462 (N_27462,N_25146,N_24947);
or U27463 (N_27463,N_24563,N_24850);
xor U27464 (N_27464,N_24458,N_24003);
nor U27465 (N_27465,N_25533,N_24378);
xor U27466 (N_27466,N_25548,N_24355);
nor U27467 (N_27467,N_24765,N_25018);
and U27468 (N_27468,N_24260,N_24250);
xor U27469 (N_27469,N_24909,N_24497);
nand U27470 (N_27470,N_24156,N_24900);
and U27471 (N_27471,N_24289,N_24679);
nand U27472 (N_27472,N_24693,N_25299);
nand U27473 (N_27473,N_25019,N_24208);
and U27474 (N_27474,N_24767,N_25813);
nor U27475 (N_27475,N_25085,N_25012);
and U27476 (N_27476,N_25344,N_24690);
nor U27477 (N_27477,N_25435,N_25025);
and U27478 (N_27478,N_24237,N_25846);
xor U27479 (N_27479,N_25663,N_24552);
or U27480 (N_27480,N_25883,N_24652);
xor U27481 (N_27481,N_24150,N_25163);
and U27482 (N_27482,N_24109,N_24789);
nor U27483 (N_27483,N_25315,N_24104);
or U27484 (N_27484,N_24680,N_24886);
xnor U27485 (N_27485,N_25909,N_24482);
or U27486 (N_27486,N_24829,N_24033);
nor U27487 (N_27487,N_25979,N_24829);
nand U27488 (N_27488,N_24337,N_24612);
or U27489 (N_27489,N_24823,N_25138);
xnor U27490 (N_27490,N_25631,N_25623);
nand U27491 (N_27491,N_25068,N_25233);
xnor U27492 (N_27492,N_24127,N_25561);
nand U27493 (N_27493,N_25184,N_25507);
nor U27494 (N_27494,N_25361,N_24818);
xor U27495 (N_27495,N_25109,N_25500);
or U27496 (N_27496,N_24904,N_24212);
nor U27497 (N_27497,N_24557,N_25869);
nor U27498 (N_27498,N_25842,N_24653);
xnor U27499 (N_27499,N_25822,N_25590);
nand U27500 (N_27500,N_25831,N_24146);
nor U27501 (N_27501,N_25374,N_25500);
xnor U27502 (N_27502,N_24126,N_25230);
nand U27503 (N_27503,N_24513,N_25405);
and U27504 (N_27504,N_24816,N_25603);
and U27505 (N_27505,N_24938,N_24466);
xor U27506 (N_27506,N_25767,N_24681);
or U27507 (N_27507,N_25106,N_24247);
xor U27508 (N_27508,N_24646,N_25349);
or U27509 (N_27509,N_24257,N_24947);
nand U27510 (N_27510,N_24708,N_24799);
or U27511 (N_27511,N_25905,N_24154);
and U27512 (N_27512,N_24378,N_24984);
and U27513 (N_27513,N_24026,N_24344);
nor U27514 (N_27514,N_24749,N_25950);
nor U27515 (N_27515,N_25630,N_24093);
nor U27516 (N_27516,N_24305,N_25931);
and U27517 (N_27517,N_25150,N_25511);
and U27518 (N_27518,N_25793,N_24853);
nand U27519 (N_27519,N_25841,N_24063);
nor U27520 (N_27520,N_25892,N_25246);
or U27521 (N_27521,N_24739,N_25108);
or U27522 (N_27522,N_25147,N_25544);
nor U27523 (N_27523,N_25122,N_25045);
nand U27524 (N_27524,N_25257,N_24957);
or U27525 (N_27525,N_25122,N_25504);
and U27526 (N_27526,N_25871,N_24415);
nor U27527 (N_27527,N_25905,N_24890);
nand U27528 (N_27528,N_24547,N_25159);
nor U27529 (N_27529,N_25145,N_25576);
nor U27530 (N_27530,N_25563,N_25207);
nor U27531 (N_27531,N_24832,N_25533);
and U27532 (N_27532,N_24056,N_25870);
and U27533 (N_27533,N_25095,N_24559);
nand U27534 (N_27534,N_25306,N_25343);
xnor U27535 (N_27535,N_25061,N_24187);
or U27536 (N_27536,N_24055,N_24862);
nor U27537 (N_27537,N_25352,N_24205);
nor U27538 (N_27538,N_24347,N_25139);
nor U27539 (N_27539,N_25980,N_25587);
nor U27540 (N_27540,N_25559,N_24249);
or U27541 (N_27541,N_24139,N_24966);
or U27542 (N_27542,N_25983,N_24242);
nand U27543 (N_27543,N_24326,N_24551);
and U27544 (N_27544,N_25614,N_24498);
xor U27545 (N_27545,N_24753,N_25348);
or U27546 (N_27546,N_24565,N_25285);
nand U27547 (N_27547,N_24318,N_24789);
nand U27548 (N_27548,N_24772,N_24607);
xor U27549 (N_27549,N_25993,N_24945);
or U27550 (N_27550,N_24383,N_25356);
nand U27551 (N_27551,N_24412,N_25522);
or U27552 (N_27552,N_24234,N_24845);
and U27553 (N_27553,N_24073,N_24199);
and U27554 (N_27554,N_25512,N_25540);
xnor U27555 (N_27555,N_25117,N_25431);
nand U27556 (N_27556,N_25973,N_24966);
or U27557 (N_27557,N_25410,N_25403);
and U27558 (N_27558,N_25212,N_25327);
nand U27559 (N_27559,N_24132,N_24876);
nor U27560 (N_27560,N_25382,N_25001);
nand U27561 (N_27561,N_25330,N_25251);
or U27562 (N_27562,N_24696,N_24189);
nand U27563 (N_27563,N_25149,N_25115);
nor U27564 (N_27564,N_25715,N_25174);
nand U27565 (N_27565,N_24194,N_25069);
and U27566 (N_27566,N_24828,N_25616);
nand U27567 (N_27567,N_24446,N_25322);
nand U27568 (N_27568,N_25516,N_25492);
or U27569 (N_27569,N_24119,N_24408);
and U27570 (N_27570,N_24840,N_24961);
or U27571 (N_27571,N_25807,N_25466);
xnor U27572 (N_27572,N_24755,N_25366);
and U27573 (N_27573,N_24852,N_25845);
and U27574 (N_27574,N_25414,N_24837);
nor U27575 (N_27575,N_25189,N_24029);
or U27576 (N_27576,N_25087,N_25523);
and U27577 (N_27577,N_25015,N_25837);
nor U27578 (N_27578,N_24043,N_24136);
and U27579 (N_27579,N_24550,N_24861);
xor U27580 (N_27580,N_24558,N_24916);
nor U27581 (N_27581,N_25302,N_24116);
and U27582 (N_27582,N_25858,N_24184);
xor U27583 (N_27583,N_24827,N_24255);
nand U27584 (N_27584,N_24475,N_24010);
nor U27585 (N_27585,N_24783,N_24334);
xnor U27586 (N_27586,N_25745,N_25068);
and U27587 (N_27587,N_25445,N_24640);
and U27588 (N_27588,N_24524,N_25136);
xor U27589 (N_27589,N_24550,N_25688);
xnor U27590 (N_27590,N_24120,N_25625);
nand U27591 (N_27591,N_24363,N_25951);
nand U27592 (N_27592,N_24539,N_24176);
nand U27593 (N_27593,N_25577,N_24153);
and U27594 (N_27594,N_24902,N_25728);
and U27595 (N_27595,N_24648,N_24241);
xnor U27596 (N_27596,N_24159,N_25684);
or U27597 (N_27597,N_24442,N_25999);
xor U27598 (N_27598,N_24570,N_25285);
or U27599 (N_27599,N_25788,N_24121);
nand U27600 (N_27600,N_24684,N_24795);
and U27601 (N_27601,N_24448,N_24004);
xnor U27602 (N_27602,N_24073,N_25337);
and U27603 (N_27603,N_24359,N_24558);
or U27604 (N_27604,N_24183,N_25956);
nor U27605 (N_27605,N_24319,N_24162);
xor U27606 (N_27606,N_25409,N_25261);
nor U27607 (N_27607,N_25716,N_24873);
xnor U27608 (N_27608,N_24545,N_24493);
nor U27609 (N_27609,N_25333,N_25114);
nand U27610 (N_27610,N_24115,N_24194);
nand U27611 (N_27611,N_24357,N_24934);
nand U27612 (N_27612,N_24565,N_24492);
nand U27613 (N_27613,N_25235,N_24676);
or U27614 (N_27614,N_25824,N_25072);
nand U27615 (N_27615,N_25724,N_24012);
nand U27616 (N_27616,N_24864,N_25717);
xnor U27617 (N_27617,N_24759,N_25981);
nor U27618 (N_27618,N_25714,N_24935);
xnor U27619 (N_27619,N_24524,N_25428);
nor U27620 (N_27620,N_24926,N_24310);
xor U27621 (N_27621,N_25332,N_25141);
nor U27622 (N_27622,N_24446,N_24805);
and U27623 (N_27623,N_24373,N_24389);
and U27624 (N_27624,N_25865,N_25204);
or U27625 (N_27625,N_25056,N_25794);
and U27626 (N_27626,N_24532,N_25953);
nand U27627 (N_27627,N_24424,N_25389);
nand U27628 (N_27628,N_25413,N_25631);
nor U27629 (N_27629,N_25111,N_24885);
xor U27630 (N_27630,N_24456,N_24092);
or U27631 (N_27631,N_24807,N_24220);
or U27632 (N_27632,N_25700,N_25005);
or U27633 (N_27633,N_24975,N_24869);
xor U27634 (N_27634,N_25679,N_25943);
nand U27635 (N_27635,N_24287,N_24998);
xnor U27636 (N_27636,N_24613,N_24205);
xnor U27637 (N_27637,N_25129,N_24101);
xor U27638 (N_27638,N_25153,N_25294);
and U27639 (N_27639,N_25133,N_24198);
and U27640 (N_27640,N_25538,N_24680);
nor U27641 (N_27641,N_25407,N_25851);
nor U27642 (N_27642,N_24238,N_24893);
xnor U27643 (N_27643,N_25580,N_24505);
nor U27644 (N_27644,N_24822,N_25793);
nor U27645 (N_27645,N_25383,N_25037);
and U27646 (N_27646,N_24679,N_24143);
and U27647 (N_27647,N_25135,N_25282);
or U27648 (N_27648,N_24765,N_25434);
and U27649 (N_27649,N_24888,N_24055);
and U27650 (N_27650,N_25345,N_25291);
nand U27651 (N_27651,N_25899,N_25283);
xnor U27652 (N_27652,N_24123,N_24683);
nand U27653 (N_27653,N_24063,N_24578);
xor U27654 (N_27654,N_24755,N_24935);
nor U27655 (N_27655,N_24335,N_24981);
or U27656 (N_27656,N_25745,N_25603);
or U27657 (N_27657,N_24755,N_24277);
and U27658 (N_27658,N_25164,N_24628);
or U27659 (N_27659,N_25965,N_25057);
nand U27660 (N_27660,N_24293,N_25885);
xnor U27661 (N_27661,N_25629,N_25714);
nor U27662 (N_27662,N_24843,N_25205);
or U27663 (N_27663,N_24083,N_24501);
or U27664 (N_27664,N_24819,N_24214);
or U27665 (N_27665,N_24403,N_25154);
xor U27666 (N_27666,N_24202,N_25619);
or U27667 (N_27667,N_25209,N_25728);
nand U27668 (N_27668,N_25471,N_24919);
xor U27669 (N_27669,N_25624,N_25249);
or U27670 (N_27670,N_25827,N_24386);
nor U27671 (N_27671,N_24164,N_24676);
xor U27672 (N_27672,N_25580,N_25256);
nand U27673 (N_27673,N_24849,N_24871);
nand U27674 (N_27674,N_24555,N_24243);
nor U27675 (N_27675,N_24055,N_24300);
nor U27676 (N_27676,N_25341,N_24284);
nand U27677 (N_27677,N_24278,N_24797);
or U27678 (N_27678,N_24181,N_24481);
and U27679 (N_27679,N_24924,N_24138);
or U27680 (N_27680,N_24880,N_24621);
nor U27681 (N_27681,N_25913,N_25904);
xor U27682 (N_27682,N_25839,N_25411);
xnor U27683 (N_27683,N_24820,N_25084);
xor U27684 (N_27684,N_24576,N_25072);
xor U27685 (N_27685,N_24633,N_25962);
or U27686 (N_27686,N_25236,N_25709);
nand U27687 (N_27687,N_25164,N_25048);
xor U27688 (N_27688,N_24471,N_24970);
xor U27689 (N_27689,N_24823,N_24267);
and U27690 (N_27690,N_24803,N_25057);
xnor U27691 (N_27691,N_24887,N_25299);
or U27692 (N_27692,N_24983,N_24245);
or U27693 (N_27693,N_25031,N_25856);
xor U27694 (N_27694,N_24120,N_24633);
or U27695 (N_27695,N_25787,N_25206);
nor U27696 (N_27696,N_25045,N_24545);
or U27697 (N_27697,N_25045,N_24106);
or U27698 (N_27698,N_25512,N_25754);
and U27699 (N_27699,N_25631,N_25370);
nand U27700 (N_27700,N_24906,N_24311);
nand U27701 (N_27701,N_25496,N_24696);
xnor U27702 (N_27702,N_25426,N_24080);
xor U27703 (N_27703,N_25115,N_25356);
and U27704 (N_27704,N_24483,N_24924);
nor U27705 (N_27705,N_24961,N_25097);
nand U27706 (N_27706,N_24000,N_24242);
xnor U27707 (N_27707,N_25363,N_24732);
xnor U27708 (N_27708,N_25785,N_25463);
and U27709 (N_27709,N_25984,N_25107);
or U27710 (N_27710,N_24756,N_25191);
or U27711 (N_27711,N_24072,N_25421);
and U27712 (N_27712,N_24226,N_25615);
and U27713 (N_27713,N_24972,N_25987);
nor U27714 (N_27714,N_24039,N_24476);
xnor U27715 (N_27715,N_25214,N_24428);
nor U27716 (N_27716,N_24520,N_24482);
or U27717 (N_27717,N_24278,N_24821);
nor U27718 (N_27718,N_24929,N_24578);
and U27719 (N_27719,N_25622,N_25749);
nor U27720 (N_27720,N_24995,N_24496);
or U27721 (N_27721,N_24263,N_25739);
nand U27722 (N_27722,N_24309,N_24477);
nand U27723 (N_27723,N_24897,N_25003);
or U27724 (N_27724,N_25454,N_24267);
and U27725 (N_27725,N_25170,N_25582);
or U27726 (N_27726,N_25810,N_25608);
xor U27727 (N_27727,N_25612,N_25365);
nor U27728 (N_27728,N_24487,N_25902);
nor U27729 (N_27729,N_24350,N_24056);
nor U27730 (N_27730,N_25272,N_24543);
nor U27731 (N_27731,N_25938,N_24387);
nor U27732 (N_27732,N_24075,N_24401);
nand U27733 (N_27733,N_25483,N_25544);
and U27734 (N_27734,N_25342,N_25068);
or U27735 (N_27735,N_24813,N_24106);
xnor U27736 (N_27736,N_24047,N_25207);
xnor U27737 (N_27737,N_25119,N_24973);
and U27738 (N_27738,N_25668,N_25624);
nand U27739 (N_27739,N_25167,N_24456);
and U27740 (N_27740,N_24264,N_25194);
nand U27741 (N_27741,N_25876,N_25385);
and U27742 (N_27742,N_25659,N_25385);
or U27743 (N_27743,N_25071,N_25533);
nand U27744 (N_27744,N_25408,N_25817);
or U27745 (N_27745,N_25264,N_25845);
or U27746 (N_27746,N_25906,N_24681);
or U27747 (N_27747,N_25006,N_25226);
nand U27748 (N_27748,N_24599,N_24883);
xnor U27749 (N_27749,N_24322,N_25005);
or U27750 (N_27750,N_24107,N_24072);
xnor U27751 (N_27751,N_25698,N_24580);
or U27752 (N_27752,N_25810,N_24586);
or U27753 (N_27753,N_25005,N_24581);
nor U27754 (N_27754,N_25753,N_25510);
nand U27755 (N_27755,N_24316,N_24274);
and U27756 (N_27756,N_25585,N_25533);
nand U27757 (N_27757,N_24008,N_24361);
or U27758 (N_27758,N_25192,N_25558);
or U27759 (N_27759,N_25532,N_24932);
and U27760 (N_27760,N_25876,N_24832);
and U27761 (N_27761,N_24938,N_24796);
nor U27762 (N_27762,N_24985,N_25812);
and U27763 (N_27763,N_24647,N_25127);
or U27764 (N_27764,N_25390,N_25807);
nor U27765 (N_27765,N_24061,N_24348);
xor U27766 (N_27766,N_25910,N_24952);
and U27767 (N_27767,N_25911,N_24772);
xor U27768 (N_27768,N_24793,N_25817);
xor U27769 (N_27769,N_25179,N_24126);
nand U27770 (N_27770,N_24914,N_24394);
and U27771 (N_27771,N_25930,N_24062);
or U27772 (N_27772,N_25080,N_24896);
nor U27773 (N_27773,N_24742,N_24860);
and U27774 (N_27774,N_24557,N_25749);
xnor U27775 (N_27775,N_25993,N_24589);
and U27776 (N_27776,N_24190,N_24153);
nor U27777 (N_27777,N_24104,N_24875);
nand U27778 (N_27778,N_24022,N_24065);
xnor U27779 (N_27779,N_24881,N_24130);
or U27780 (N_27780,N_24303,N_25557);
nor U27781 (N_27781,N_24987,N_25065);
nor U27782 (N_27782,N_24703,N_25101);
nand U27783 (N_27783,N_25735,N_25849);
or U27784 (N_27784,N_25332,N_25266);
or U27785 (N_27785,N_24389,N_24661);
or U27786 (N_27786,N_24553,N_25244);
or U27787 (N_27787,N_25154,N_24480);
nand U27788 (N_27788,N_24301,N_24132);
or U27789 (N_27789,N_25254,N_24348);
or U27790 (N_27790,N_24924,N_24645);
xor U27791 (N_27791,N_24117,N_24346);
or U27792 (N_27792,N_25712,N_24970);
xnor U27793 (N_27793,N_24067,N_24238);
xnor U27794 (N_27794,N_24562,N_25874);
xor U27795 (N_27795,N_25834,N_24833);
nand U27796 (N_27796,N_25364,N_25296);
xor U27797 (N_27797,N_24345,N_25634);
and U27798 (N_27798,N_24636,N_25422);
xnor U27799 (N_27799,N_25265,N_25570);
nor U27800 (N_27800,N_25263,N_24914);
nor U27801 (N_27801,N_25371,N_25083);
xor U27802 (N_27802,N_25792,N_24595);
and U27803 (N_27803,N_25750,N_25567);
xnor U27804 (N_27804,N_24929,N_25257);
nor U27805 (N_27805,N_25022,N_25555);
and U27806 (N_27806,N_24686,N_24307);
nand U27807 (N_27807,N_24321,N_25478);
xor U27808 (N_27808,N_25348,N_24621);
nor U27809 (N_27809,N_24312,N_25668);
nor U27810 (N_27810,N_24741,N_24929);
nor U27811 (N_27811,N_25205,N_24247);
nor U27812 (N_27812,N_25453,N_24237);
or U27813 (N_27813,N_25871,N_24001);
nand U27814 (N_27814,N_24699,N_24528);
or U27815 (N_27815,N_25778,N_24228);
nor U27816 (N_27816,N_24843,N_25133);
xor U27817 (N_27817,N_25514,N_24876);
nand U27818 (N_27818,N_25435,N_24626);
and U27819 (N_27819,N_25041,N_25947);
xnor U27820 (N_27820,N_25593,N_24006);
and U27821 (N_27821,N_24469,N_24417);
and U27822 (N_27822,N_24640,N_25478);
nor U27823 (N_27823,N_25136,N_24077);
nor U27824 (N_27824,N_24340,N_25582);
xnor U27825 (N_27825,N_25000,N_24860);
or U27826 (N_27826,N_25025,N_25966);
or U27827 (N_27827,N_24185,N_25049);
and U27828 (N_27828,N_25031,N_24148);
or U27829 (N_27829,N_25903,N_24792);
or U27830 (N_27830,N_24100,N_24309);
nand U27831 (N_27831,N_25372,N_24182);
and U27832 (N_27832,N_24607,N_24055);
xor U27833 (N_27833,N_24864,N_25776);
nor U27834 (N_27834,N_25337,N_24808);
nor U27835 (N_27835,N_25928,N_25288);
or U27836 (N_27836,N_25656,N_24098);
nor U27837 (N_27837,N_24359,N_24037);
xor U27838 (N_27838,N_25202,N_24723);
or U27839 (N_27839,N_25606,N_24765);
nand U27840 (N_27840,N_25325,N_24953);
nor U27841 (N_27841,N_24249,N_25762);
xnor U27842 (N_27842,N_24295,N_25333);
xor U27843 (N_27843,N_25125,N_24643);
and U27844 (N_27844,N_25760,N_25929);
and U27845 (N_27845,N_24629,N_24278);
xnor U27846 (N_27846,N_24114,N_25234);
nand U27847 (N_27847,N_25908,N_24544);
xnor U27848 (N_27848,N_24537,N_24542);
or U27849 (N_27849,N_24636,N_24358);
xor U27850 (N_27850,N_25510,N_24293);
nand U27851 (N_27851,N_24263,N_25086);
and U27852 (N_27852,N_24775,N_25580);
and U27853 (N_27853,N_25073,N_24144);
nand U27854 (N_27854,N_25726,N_24577);
nand U27855 (N_27855,N_25885,N_25269);
nor U27856 (N_27856,N_25738,N_24943);
or U27857 (N_27857,N_24615,N_24972);
and U27858 (N_27858,N_24737,N_25404);
xor U27859 (N_27859,N_25139,N_24885);
xnor U27860 (N_27860,N_24012,N_24165);
nand U27861 (N_27861,N_24303,N_25543);
or U27862 (N_27862,N_25200,N_24478);
xnor U27863 (N_27863,N_24727,N_24821);
nor U27864 (N_27864,N_25255,N_25903);
nand U27865 (N_27865,N_24312,N_25876);
xor U27866 (N_27866,N_24106,N_24986);
xnor U27867 (N_27867,N_25246,N_25903);
nor U27868 (N_27868,N_24443,N_24012);
nand U27869 (N_27869,N_25351,N_25285);
nand U27870 (N_27870,N_25175,N_25270);
and U27871 (N_27871,N_24016,N_24270);
xnor U27872 (N_27872,N_24223,N_25849);
nor U27873 (N_27873,N_25882,N_25815);
or U27874 (N_27874,N_25844,N_24870);
xor U27875 (N_27875,N_25499,N_25800);
nand U27876 (N_27876,N_24164,N_25709);
nor U27877 (N_27877,N_24796,N_25314);
xnor U27878 (N_27878,N_24794,N_24719);
nor U27879 (N_27879,N_24465,N_25904);
or U27880 (N_27880,N_25823,N_25155);
nand U27881 (N_27881,N_25879,N_25887);
xnor U27882 (N_27882,N_24041,N_25146);
nand U27883 (N_27883,N_24953,N_24373);
nand U27884 (N_27884,N_24966,N_25236);
nor U27885 (N_27885,N_24490,N_25749);
nand U27886 (N_27886,N_24094,N_24005);
nor U27887 (N_27887,N_24841,N_25710);
nand U27888 (N_27888,N_25422,N_24792);
nand U27889 (N_27889,N_24948,N_25196);
nand U27890 (N_27890,N_24610,N_25826);
nor U27891 (N_27891,N_25345,N_24462);
and U27892 (N_27892,N_25190,N_25710);
nand U27893 (N_27893,N_24211,N_25170);
xor U27894 (N_27894,N_24962,N_24328);
nand U27895 (N_27895,N_25020,N_25228);
and U27896 (N_27896,N_24432,N_25666);
and U27897 (N_27897,N_25952,N_25971);
xnor U27898 (N_27898,N_24008,N_25840);
xor U27899 (N_27899,N_25352,N_24384);
and U27900 (N_27900,N_25794,N_24464);
nand U27901 (N_27901,N_24015,N_25825);
nor U27902 (N_27902,N_25589,N_25733);
nor U27903 (N_27903,N_25554,N_24907);
nand U27904 (N_27904,N_24945,N_24250);
nor U27905 (N_27905,N_24111,N_24528);
nand U27906 (N_27906,N_24875,N_24735);
or U27907 (N_27907,N_24468,N_25083);
or U27908 (N_27908,N_25100,N_25442);
nand U27909 (N_27909,N_24542,N_25558);
and U27910 (N_27910,N_24731,N_24726);
or U27911 (N_27911,N_24704,N_25940);
nand U27912 (N_27912,N_25622,N_25104);
and U27913 (N_27913,N_25603,N_25875);
nor U27914 (N_27914,N_25405,N_24859);
nor U27915 (N_27915,N_24648,N_25960);
nand U27916 (N_27916,N_25466,N_24107);
or U27917 (N_27917,N_25546,N_25669);
or U27918 (N_27918,N_24556,N_24386);
xnor U27919 (N_27919,N_24591,N_24920);
xnor U27920 (N_27920,N_25582,N_25971);
and U27921 (N_27921,N_25124,N_24521);
nand U27922 (N_27922,N_24097,N_25476);
and U27923 (N_27923,N_25826,N_25540);
nor U27924 (N_27924,N_24319,N_25923);
nand U27925 (N_27925,N_25653,N_25555);
nor U27926 (N_27926,N_25058,N_25525);
nand U27927 (N_27927,N_24152,N_24886);
and U27928 (N_27928,N_24396,N_24406);
nand U27929 (N_27929,N_24658,N_25797);
and U27930 (N_27930,N_25328,N_25312);
and U27931 (N_27931,N_24283,N_24372);
nor U27932 (N_27932,N_24216,N_25508);
or U27933 (N_27933,N_25453,N_24412);
nor U27934 (N_27934,N_24779,N_24868);
nor U27935 (N_27935,N_25413,N_24556);
and U27936 (N_27936,N_25139,N_25448);
and U27937 (N_27937,N_24401,N_25999);
xor U27938 (N_27938,N_25877,N_25083);
nand U27939 (N_27939,N_25233,N_25617);
nor U27940 (N_27940,N_24897,N_25890);
or U27941 (N_27941,N_24198,N_24658);
nand U27942 (N_27942,N_24130,N_24420);
and U27943 (N_27943,N_24075,N_24972);
xor U27944 (N_27944,N_24529,N_25376);
nor U27945 (N_27945,N_25607,N_24732);
or U27946 (N_27946,N_25350,N_25857);
and U27947 (N_27947,N_25445,N_24314);
and U27948 (N_27948,N_25879,N_25462);
or U27949 (N_27949,N_24513,N_25600);
xnor U27950 (N_27950,N_25962,N_25730);
or U27951 (N_27951,N_24763,N_24569);
and U27952 (N_27952,N_25426,N_24140);
xnor U27953 (N_27953,N_24589,N_24751);
nor U27954 (N_27954,N_24091,N_24671);
and U27955 (N_27955,N_24652,N_24150);
nor U27956 (N_27956,N_25655,N_25780);
nand U27957 (N_27957,N_24911,N_25772);
nor U27958 (N_27958,N_25039,N_25206);
nor U27959 (N_27959,N_24003,N_24799);
and U27960 (N_27960,N_25997,N_25024);
nand U27961 (N_27961,N_25115,N_25140);
nor U27962 (N_27962,N_25794,N_25313);
or U27963 (N_27963,N_25266,N_24314);
nand U27964 (N_27964,N_25905,N_24578);
nand U27965 (N_27965,N_25308,N_24108);
nor U27966 (N_27966,N_25280,N_24189);
or U27967 (N_27967,N_24551,N_24370);
or U27968 (N_27968,N_25462,N_25442);
and U27969 (N_27969,N_24169,N_24323);
and U27970 (N_27970,N_24013,N_24318);
nor U27971 (N_27971,N_25034,N_24695);
and U27972 (N_27972,N_25259,N_25935);
or U27973 (N_27973,N_24442,N_24681);
nand U27974 (N_27974,N_25936,N_25721);
and U27975 (N_27975,N_25008,N_25068);
and U27976 (N_27976,N_24898,N_24610);
and U27977 (N_27977,N_25220,N_25925);
and U27978 (N_27978,N_25984,N_24214);
or U27979 (N_27979,N_25834,N_24446);
and U27980 (N_27980,N_24952,N_24238);
nor U27981 (N_27981,N_25110,N_25276);
xor U27982 (N_27982,N_25349,N_25596);
nand U27983 (N_27983,N_25429,N_25597);
nor U27984 (N_27984,N_25956,N_25953);
or U27985 (N_27985,N_24804,N_25390);
or U27986 (N_27986,N_25264,N_25232);
nor U27987 (N_27987,N_24160,N_25278);
or U27988 (N_27988,N_25171,N_25845);
and U27989 (N_27989,N_24478,N_25504);
xor U27990 (N_27990,N_25722,N_25400);
or U27991 (N_27991,N_25619,N_24999);
nand U27992 (N_27992,N_24191,N_24055);
or U27993 (N_27993,N_25923,N_24839);
nand U27994 (N_27994,N_25846,N_24726);
xnor U27995 (N_27995,N_24365,N_24809);
nand U27996 (N_27996,N_25157,N_25326);
or U27997 (N_27997,N_24101,N_25233);
nand U27998 (N_27998,N_24724,N_24897);
and U27999 (N_27999,N_25634,N_25339);
or U28000 (N_28000,N_26153,N_26446);
nor U28001 (N_28001,N_27847,N_27287);
xor U28002 (N_28002,N_27357,N_27265);
or U28003 (N_28003,N_26002,N_26457);
and U28004 (N_28004,N_26104,N_26490);
nor U28005 (N_28005,N_26932,N_27743);
nor U28006 (N_28006,N_26098,N_26456);
or U28007 (N_28007,N_27311,N_26889);
and U28008 (N_28008,N_26813,N_27748);
xnor U28009 (N_28009,N_26840,N_26601);
nor U28010 (N_28010,N_26673,N_27304);
xnor U28011 (N_28011,N_27728,N_26450);
and U28012 (N_28012,N_26691,N_26690);
xnor U28013 (N_28013,N_27073,N_27064);
nor U28014 (N_28014,N_26864,N_26349);
and U28015 (N_28015,N_26692,N_27333);
xor U28016 (N_28016,N_26614,N_27288);
xor U28017 (N_28017,N_26848,N_27985);
nor U28018 (N_28018,N_27734,N_27250);
nor U28019 (N_28019,N_26133,N_26972);
xor U28020 (N_28020,N_26677,N_27114);
xor U28021 (N_28021,N_27701,N_26005);
and U28022 (N_28022,N_26508,N_27087);
or U28023 (N_28023,N_27075,N_26917);
nor U28024 (N_28024,N_26925,N_26953);
or U28025 (N_28025,N_27101,N_26333);
nor U28026 (N_28026,N_26383,N_27371);
or U28027 (N_28027,N_27082,N_27295);
or U28028 (N_28028,N_27200,N_26150);
nand U28029 (N_28029,N_27724,N_27320);
xor U28030 (N_28030,N_27566,N_27406);
or U28031 (N_28031,N_27279,N_26777);
nand U28032 (N_28032,N_27548,N_27430);
and U28033 (N_28033,N_26334,N_26482);
or U28034 (N_28034,N_27874,N_27573);
nor U28035 (N_28035,N_27219,N_27414);
nand U28036 (N_28036,N_26294,N_27811);
xor U28037 (N_28037,N_26548,N_27793);
nor U28038 (N_28038,N_27998,N_27307);
nand U28039 (N_28039,N_27987,N_27753);
nor U28040 (N_28040,N_27834,N_27084);
and U28041 (N_28041,N_27280,N_26979);
and U28042 (N_28042,N_26912,N_27079);
and U28043 (N_28043,N_26125,N_26453);
or U28044 (N_28044,N_26113,N_27722);
and U28045 (N_28045,N_27435,N_26035);
nand U28046 (N_28046,N_26866,N_27096);
xor U28047 (N_28047,N_26720,N_26189);
and U28048 (N_28048,N_26049,N_27169);
or U28049 (N_28049,N_26998,N_27737);
xnor U28050 (N_28050,N_27469,N_26760);
nor U28051 (N_28051,N_26629,N_27606);
or U28052 (N_28052,N_26513,N_26080);
nand U28053 (N_28053,N_27090,N_27652);
nor U28054 (N_28054,N_26209,N_26352);
and U28055 (N_28055,N_26694,N_26213);
nand U28056 (N_28056,N_27958,N_27116);
and U28057 (N_28057,N_26770,N_27954);
nor U28058 (N_28058,N_27057,N_26410);
nand U28059 (N_28059,N_27345,N_27343);
or U28060 (N_28060,N_26372,N_27608);
or U28061 (N_28061,N_27058,N_27459);
xor U28062 (N_28062,N_27645,N_26245);
and U28063 (N_28063,N_26085,N_26552);
or U28064 (N_28064,N_26031,N_26585);
and U28065 (N_28065,N_27381,N_26847);
xor U28066 (N_28066,N_27156,N_27892);
or U28067 (N_28067,N_26368,N_26818);
and U28068 (N_28068,N_27106,N_27177);
xnor U28069 (N_28069,N_27820,N_27434);
nor U28070 (N_28070,N_27241,N_26976);
and U28071 (N_28071,N_27878,N_27155);
xnor U28072 (N_28072,N_27591,N_27425);
nand U28073 (N_28073,N_27725,N_26221);
or U28074 (N_28074,N_27884,N_26498);
nor U28075 (N_28075,N_27401,N_27593);
nor U28076 (N_28076,N_27668,N_27137);
or U28077 (N_28077,N_26656,N_26906);
xnor U28078 (N_28078,N_26949,N_26657);
nor U28079 (N_28079,N_27331,N_26991);
xnor U28080 (N_28080,N_27220,N_26149);
and U28081 (N_28081,N_27682,N_26225);
nor U28082 (N_28082,N_26533,N_26921);
nand U28083 (N_28083,N_27324,N_26215);
nand U28084 (N_28084,N_26117,N_27512);
nand U28085 (N_28085,N_26184,N_26556);
xor U28086 (N_28086,N_26995,N_27902);
nor U28087 (N_28087,N_27749,N_26536);
or U28088 (N_28088,N_27797,N_26028);
and U28089 (N_28089,N_27654,N_26766);
and U28090 (N_28090,N_27831,N_27936);
or U28091 (N_28091,N_27230,N_27862);
nand U28092 (N_28092,N_27491,N_27024);
xnor U28093 (N_28093,N_27258,N_26255);
nor U28094 (N_28094,N_26808,N_26404);
nor U28095 (N_28095,N_27589,N_26195);
xor U28096 (N_28096,N_27395,N_26735);
xor U28097 (N_28097,N_26233,N_26376);
or U28098 (N_28098,N_26897,N_26929);
xnor U28099 (N_28099,N_26017,N_26935);
nor U28100 (N_28100,N_27359,N_26780);
xor U28101 (N_28101,N_27118,N_27933);
or U28102 (N_28102,N_27123,N_27947);
nor U28103 (N_28103,N_26711,N_27899);
nor U28104 (N_28104,N_27868,N_26105);
or U28105 (N_28105,N_27502,N_27590);
nor U28106 (N_28106,N_26712,N_27182);
nor U28107 (N_28107,N_26197,N_27270);
nand U28108 (N_28108,N_27126,N_26721);
nor U28109 (N_28109,N_26648,N_26415);
xor U28110 (N_28110,N_27976,N_27050);
or U28111 (N_28111,N_27035,N_26623);
xor U28112 (N_28112,N_27442,N_27227);
nand U28113 (N_28113,N_27198,N_27691);
xor U28114 (N_28114,N_26768,N_26190);
nor U28115 (N_28115,N_27363,N_26553);
nand U28116 (N_28116,N_26874,N_27329);
or U28117 (N_28117,N_26667,N_27763);
nor U28118 (N_28118,N_26761,N_27323);
nand U28119 (N_28119,N_27239,N_26163);
nor U28120 (N_28120,N_27208,N_26488);
and U28121 (N_28121,N_26962,N_27009);
nor U28122 (N_28122,N_27635,N_27089);
and U28123 (N_28123,N_27322,N_26134);
or U28124 (N_28124,N_26638,N_26480);
or U28125 (N_28125,N_27263,N_27594);
nand U28126 (N_28126,N_26382,N_26241);
nor U28127 (N_28127,N_27253,N_26625);
nor U28128 (N_28128,N_27383,N_26007);
or U28129 (N_28129,N_27676,N_26619);
and U28130 (N_28130,N_27928,N_27575);
or U28131 (N_28131,N_27729,N_26425);
or U28132 (N_28132,N_26173,N_26913);
xnor U28133 (N_28133,N_27153,N_26434);
xor U28134 (N_28134,N_26403,N_26736);
nor U28135 (N_28135,N_27223,N_26545);
xnor U28136 (N_28136,N_26716,N_27833);
or U28137 (N_28137,N_26154,N_26414);
nand U28138 (N_28138,N_27949,N_27555);
nand U28139 (N_28139,N_26162,N_26527);
xnor U28140 (N_28140,N_27648,N_27229);
and U28141 (N_28141,N_27694,N_27337);
nand U28142 (N_28142,N_27054,N_27489);
and U28143 (N_28143,N_26988,N_27146);
nand U28144 (N_28144,N_27744,N_26634);
nor U28145 (N_28145,N_26033,N_26621);
nand U28146 (N_28146,N_27471,N_26965);
and U28147 (N_28147,N_26474,N_26320);
nor U28148 (N_28148,N_27008,N_26140);
nand U28149 (N_28149,N_27276,N_26170);
or U28150 (N_28150,N_27463,N_26534);
or U28151 (N_28151,N_27755,N_26120);
xor U28152 (N_28152,N_27309,N_27112);
or U28153 (N_28153,N_26001,N_26159);
nand U28154 (N_28154,N_27745,N_26811);
and U28155 (N_28155,N_26771,N_26332);
nor U28156 (N_28156,N_26336,N_26769);
and U28157 (N_28157,N_26027,N_26681);
xor U28158 (N_28158,N_26158,N_27045);
nor U28159 (N_28159,N_27992,N_26139);
xor U28160 (N_28160,N_27599,N_26697);
nand U28161 (N_28161,N_27438,N_26265);
or U28162 (N_28162,N_27474,N_26807);
or U28163 (N_28163,N_26119,N_26858);
nor U28164 (N_28164,N_26798,N_27607);
nand U28165 (N_28165,N_26964,N_26520);
nand U28166 (N_28166,N_26014,N_27747);
nor U28167 (N_28167,N_27201,N_27792);
and U28168 (N_28168,N_26362,N_26039);
and U28169 (N_28169,N_27521,N_26460);
or U28170 (N_28170,N_26042,N_27735);
and U28171 (N_28171,N_27873,N_26514);
nand U28172 (N_28172,N_27937,N_26495);
and U28173 (N_28173,N_26633,N_27557);
and U28174 (N_28174,N_27213,N_27879);
nor U28175 (N_28175,N_26369,N_26090);
xor U28176 (N_28176,N_27056,N_27245);
and U28177 (N_28177,N_27060,N_26008);
xnor U28178 (N_28178,N_26538,N_27254);
nor U28179 (N_28179,N_27558,N_26996);
or U28180 (N_28180,N_26575,N_27780);
xor U28181 (N_28181,N_27188,N_27571);
nor U28182 (N_28182,N_27273,N_26955);
or U28183 (N_28183,N_27040,N_26584);
xor U28184 (N_28184,N_27789,N_27779);
nor U28185 (N_28185,N_27742,N_27181);
or U28186 (N_28186,N_26114,N_26523);
nand U28187 (N_28187,N_27563,N_26224);
and U28188 (N_28188,N_26386,N_27974);
and U28189 (N_28189,N_26805,N_26212);
nand U28190 (N_28190,N_26872,N_27605);
and U28191 (N_28191,N_26728,N_26249);
and U28192 (N_28192,N_26849,N_27487);
xnor U28193 (N_28193,N_27470,N_26370);
nor U28194 (N_28194,N_26725,N_26083);
xor U28195 (N_28195,N_26941,N_27460);
nor U28196 (N_28196,N_26572,N_26343);
nand U28197 (N_28197,N_27016,N_26016);
xor U28198 (N_28198,N_26791,N_26714);
or U28199 (N_28199,N_26522,N_27720);
nand U28200 (N_28200,N_27167,N_27003);
and U28201 (N_28201,N_27825,N_26810);
nor U28202 (N_28202,N_27516,N_26229);
nor U28203 (N_28203,N_27214,N_27835);
xnor U28204 (N_28204,N_26846,N_26885);
xor U28205 (N_28205,N_27236,N_27826);
or U28206 (N_28206,N_26240,N_26898);
or U28207 (N_28207,N_26351,N_27653);
nor U28208 (N_28208,N_26501,N_26610);
nor U28209 (N_28209,N_27247,N_27740);
nand U28210 (N_28210,N_27961,N_27634);
nor U28211 (N_28211,N_27917,N_27598);
or U28212 (N_28212,N_26424,N_26263);
and U28213 (N_28213,N_26377,N_26177);
nor U28214 (N_28214,N_26160,N_27864);
and U28215 (N_28215,N_26959,N_27702);
nor U28216 (N_28216,N_26081,N_27712);
xor U28217 (N_28217,N_27316,N_27759);
or U28218 (N_28218,N_26228,N_26686);
nor U28219 (N_28219,N_27643,N_27205);
nor U28220 (N_28220,N_26561,N_27492);
or U28221 (N_28221,N_27889,N_26128);
xnor U28222 (N_28222,N_27404,N_27582);
nor U28223 (N_28223,N_26797,N_26844);
nand U28224 (N_28224,N_26298,N_26069);
nor U28225 (N_28225,N_27681,N_26837);
and U28226 (N_28226,N_26850,N_27901);
xnor U28227 (N_28227,N_26266,N_27308);
nand U28228 (N_28228,N_26015,N_27658);
or U28229 (N_28229,N_26067,N_27911);
and U28230 (N_28230,N_26792,N_27586);
xor U28231 (N_28231,N_26824,N_26470);
and U28232 (N_28232,N_27001,N_27128);
nor U28233 (N_28233,N_27986,N_27750);
or U28234 (N_28234,N_26075,N_27120);
xor U28235 (N_28235,N_26822,N_26429);
nand U28236 (N_28236,N_27536,N_27072);
nor U28237 (N_28237,N_27785,N_26662);
and U28238 (N_28238,N_27687,N_27437);
nor U28239 (N_28239,N_27765,N_27529);
and U28240 (N_28240,N_27511,N_27385);
nand U28241 (N_28241,N_26291,N_26367);
and U28242 (N_28242,N_27962,N_27685);
nand U28243 (N_28243,N_27147,N_27637);
nor U28244 (N_28244,N_26900,N_27477);
nor U28245 (N_28245,N_27168,N_27409);
nand U28246 (N_28246,N_26518,N_26471);
xor U28247 (N_28247,N_27275,N_26682);
and U28248 (N_28248,N_27508,N_27127);
nand U28249 (N_28249,N_26688,N_27569);
xor U28250 (N_28250,N_27875,N_26264);
and U28251 (N_28251,N_27538,N_27303);
xnor U28252 (N_28252,N_27154,N_27669);
and U28253 (N_28253,N_26658,N_27306);
nor U28254 (N_28254,N_27335,N_27380);
xor U28255 (N_28255,N_27392,N_27775);
xnor U28256 (N_28256,N_27352,N_26702);
and U28257 (N_28257,N_27327,N_27952);
or U28258 (N_28258,N_27194,N_27618);
nor U28259 (N_28259,N_26216,N_27751);
xor U28260 (N_28260,N_27549,N_26786);
and U28261 (N_28261,N_27390,N_27458);
or U28262 (N_28262,N_26193,N_26003);
xnor U28263 (N_28263,N_27195,N_26011);
nor U28264 (N_28264,N_26056,N_27207);
nor U28265 (N_28265,N_26500,N_26079);
and U28266 (N_28266,N_26919,N_26109);
or U28267 (N_28267,N_26137,N_26743);
and U28268 (N_28268,N_27115,N_27131);
nand U28269 (N_28269,N_26757,N_27523);
nor U28270 (N_28270,N_26420,N_26468);
nand U28271 (N_28271,N_27543,N_26793);
xnor U28272 (N_28272,N_26254,N_27703);
and U28273 (N_28273,N_26051,N_27932);
nand U28274 (N_28274,N_26430,N_26586);
xor U28275 (N_28275,N_27157,N_27382);
nor U28276 (N_28276,N_27240,N_27465);
nand U28277 (N_28277,N_26293,N_26401);
and U28278 (N_28278,N_26999,N_26116);
xnor U28279 (N_28279,N_26274,N_27570);
nor U28280 (N_28280,N_27863,N_27774);
nor U28281 (N_28281,N_26304,N_26306);
or U28282 (N_28282,N_26243,N_27579);
xor U28283 (N_28283,N_26645,N_27778);
and U28284 (N_28284,N_27766,N_27503);
nand U28285 (N_28285,N_27528,N_26724);
and U28286 (N_28286,N_26580,N_27821);
xnor U28287 (N_28287,N_27286,N_27143);
nand U28288 (N_28288,N_27039,N_26799);
xnor U28289 (N_28289,N_27592,N_26717);
nor U28290 (N_28290,N_27705,N_26175);
xnor U28291 (N_28291,N_26022,N_26344);
xor U28292 (N_28292,N_27302,N_26251);
or U28293 (N_28293,N_26458,N_26188);
nand U28294 (N_28294,N_26568,N_26151);
or U28295 (N_28295,N_26271,N_27867);
nor U28296 (N_28296,N_27413,N_26834);
xor U28297 (N_28297,N_27232,N_27321);
nand U28298 (N_28298,N_26540,N_26603);
nor U28299 (N_28299,N_26841,N_26705);
or U28300 (N_28300,N_26882,N_27522);
and U28301 (N_28301,N_26400,N_26816);
nand U28302 (N_28302,N_27365,N_26559);
xor U28303 (N_28303,N_26359,N_26338);
xor U28304 (N_28304,N_26587,N_26931);
nor U28305 (N_28305,N_27913,N_27228);
xnor U28306 (N_28306,N_27042,N_27514);
nand U28307 (N_28307,N_27272,N_26958);
xor U28308 (N_28308,N_27074,N_26064);
and U28309 (N_28309,N_27994,N_27104);
or U28310 (N_28310,N_27204,N_26499);
and U28311 (N_28311,N_27581,N_27451);
and U28312 (N_28312,N_26172,N_26695);
or U28313 (N_28313,N_26968,N_27912);
nor U28314 (N_28314,N_27944,N_26655);
nor U28315 (N_28315,N_26024,N_27004);
and U28316 (N_28316,N_26709,N_26497);
and U28317 (N_28317,N_26218,N_27449);
xor U28318 (N_28318,N_27597,N_27047);
or U28319 (N_28319,N_27909,N_27827);
nor U28320 (N_28320,N_27876,N_27113);
and U28321 (N_28321,N_26803,N_26779);
nor U28322 (N_28322,N_26704,N_27025);
and U28323 (N_28323,N_27368,N_27010);
and U28324 (N_28324,N_26018,N_27726);
or U28325 (N_28325,N_26182,N_27824);
and U28326 (N_28326,N_27289,N_27979);
and U28327 (N_28327,N_27386,N_27028);
nor U28328 (N_28328,N_26186,N_27739);
nand U28329 (N_28329,N_27017,N_26853);
or U28330 (N_28330,N_26896,N_26099);
and U28331 (N_28331,N_27362,N_27387);
and U28332 (N_28332,N_26867,N_27354);
nor U28333 (N_28333,N_27699,N_26647);
and U28334 (N_28334,N_27325,N_27071);
nand U28335 (N_28335,N_27452,N_26396);
xor U28336 (N_28336,N_27539,N_27193);
nor U28337 (N_28337,N_26804,N_27577);
nor U28338 (N_28338,N_27540,N_27659);
and U28339 (N_28339,N_26719,N_27138);
nor U28340 (N_28340,N_27542,N_27092);
xnor U28341 (N_28341,N_26544,N_26305);
and U28342 (N_28342,N_27723,N_27269);
or U28343 (N_28343,N_26687,N_27145);
xor U28344 (N_28344,N_27799,N_26438);
nand U28345 (N_28345,N_27866,N_27209);
nand U28346 (N_28346,N_27527,N_26418);
nor U28347 (N_28347,N_26675,N_27180);
nand U28348 (N_28348,N_27215,N_26985);
or U28349 (N_28349,N_27218,N_27099);
nor U28350 (N_28350,N_26387,N_27412);
and U28351 (N_28351,N_26993,N_27211);
nand U28352 (N_28352,N_26578,N_26181);
xnor U28353 (N_28353,N_27537,N_27358);
nand U28354 (N_28354,N_26169,N_26699);
or U28355 (N_28355,N_27282,N_26258);
nor U28356 (N_28356,N_26337,N_26341);
nor U28357 (N_28357,N_27500,N_26239);
or U28358 (N_28358,N_26776,N_27688);
xnor U28359 (N_28359,N_26307,N_26318);
and U28360 (N_28360,N_26141,N_26605);
and U28361 (N_28361,N_27077,N_26023);
or U28362 (N_28362,N_26969,N_27963);
nand U28363 (N_28363,N_27741,N_26136);
xor U28364 (N_28364,N_26406,N_26875);
and U28365 (N_28365,N_27464,N_26787);
and U28366 (N_28366,N_27709,N_27633);
and U28367 (N_28367,N_26364,N_27915);
and U28368 (N_28368,N_26427,N_27495);
and U28369 (N_28369,N_27271,N_27185);
nor U28370 (N_28370,N_27107,N_27367);
xnor U28371 (N_28371,N_26895,N_26781);
xor U28372 (N_28372,N_26554,N_26296);
and U28373 (N_28373,N_27559,N_26244);
and U28374 (N_28374,N_26983,N_26506);
nor U28375 (N_28375,N_27670,N_26835);
nand U28376 (N_28376,N_26641,N_27429);
or U28377 (N_28377,N_27388,N_27910);
or U28378 (N_28378,N_26636,N_26130);
or U28379 (N_28379,N_26502,N_27697);
nor U28380 (N_28380,N_26507,N_27501);
and U28381 (N_28381,N_27475,N_26004);
nand U28382 (N_28382,N_27150,N_27338);
and U28383 (N_28383,N_26600,N_27574);
nor U28384 (N_28384,N_26063,N_27266);
and U28385 (N_28385,N_27069,N_26103);
or U28386 (N_28386,N_27890,N_27224);
nor U28387 (N_28387,N_26135,N_27922);
and U28388 (N_28388,N_26746,N_26970);
xor U28389 (N_28389,N_26801,N_26576);
nand U28390 (N_28390,N_26166,N_27334);
or U28391 (N_28391,N_26185,N_27373);
and U28392 (N_28392,N_27795,N_26562);
nor U28393 (N_28393,N_26577,N_27353);
and U28394 (N_28394,N_26558,N_27408);
xnor U28395 (N_28395,N_27485,N_27070);
xnor U28396 (N_28396,N_27830,N_27715);
nor U28397 (N_28397,N_27718,N_26280);
xor U28398 (N_28398,N_26363,N_26171);
nor U28399 (N_28399,N_26459,N_27533);
or U28400 (N_28400,N_27545,N_27350);
and U28401 (N_28401,N_26237,N_27706);
xnor U28402 (N_28402,N_27342,N_26309);
xnor U28403 (N_28403,N_27950,N_26591);
and U28404 (N_28404,N_26532,N_26530);
and U28405 (N_28405,N_27340,N_27535);
nand U28406 (N_28406,N_27339,N_27907);
xnor U28407 (N_28407,N_26358,N_27033);
nand U28408 (N_28408,N_26944,N_26744);
nor U28409 (N_28409,N_26951,N_26029);
nand U28410 (N_28410,N_26250,N_26062);
nor U28411 (N_28411,N_26903,N_26515);
nor U28412 (N_28412,N_27488,N_27777);
nand U28413 (N_28413,N_27203,N_27552);
nand U28414 (N_28414,N_27020,N_26025);
xnor U28415 (N_28415,N_27030,N_27479);
xor U28416 (N_28416,N_27317,N_26191);
xor U28417 (N_28417,N_27291,N_26628);
nor U28418 (N_28418,N_27807,N_27233);
or U28419 (N_28419,N_26392,N_27615);
nor U28420 (N_28420,N_26129,N_26829);
nand U28421 (N_28421,N_26065,N_26060);
nand U28422 (N_28422,N_26618,N_26013);
xor U28423 (N_28423,N_27490,N_26248);
nor U28424 (N_28424,N_27657,N_26200);
or U28425 (N_28425,N_26557,N_26879);
xnor U28426 (N_28426,N_27956,N_26464);
nand U28427 (N_28427,N_26087,N_27315);
nand U28428 (N_28428,N_26748,N_27776);
or U28429 (N_28429,N_26624,N_27731);
and U28430 (N_28430,N_27088,N_27173);
and U28431 (N_28431,N_27292,N_26143);
or U28432 (N_28432,N_26930,N_27190);
and U28433 (N_28433,N_27256,N_26583);
nor U28434 (N_28434,N_27832,N_27556);
nand U28435 (N_28435,N_27666,N_27930);
xnor U28436 (N_28436,N_26204,N_26282);
or U28437 (N_28437,N_27617,N_26521);
and U28438 (N_28438,N_26142,N_27671);
or U28439 (N_28439,N_27945,N_27225);
or U28440 (N_28440,N_26990,N_27631);
nand U28441 (N_28441,N_27441,N_27237);
or U28442 (N_28442,N_26977,N_27132);
and U28443 (N_28443,N_27360,N_27692);
nand U28444 (N_28444,N_26432,N_26071);
nand U28445 (N_28445,N_27984,N_26205);
nand U28446 (N_28446,N_26000,N_26830);
nor U28447 (N_28447,N_27496,N_26426);
nand U28448 (N_28448,N_26974,N_27453);
or U28449 (N_28449,N_26541,N_27328);
xor U28450 (N_28450,N_27419,N_27898);
nand U28451 (N_28451,N_27758,N_26617);
or U28452 (N_28452,N_26108,N_26884);
or U28453 (N_28453,N_27544,N_27134);
xnor U28454 (N_28454,N_26503,N_27038);
xnor U28455 (N_28455,N_26772,N_26978);
or U28456 (N_28456,N_27431,N_27921);
nand U28457 (N_28457,N_26402,N_27843);
xor U28458 (N_28458,N_26942,N_27858);
and U28459 (N_28459,N_26321,N_26272);
xnor U28460 (N_28460,N_27052,N_27663);
or U28461 (N_28461,N_26411,N_27923);
or U28462 (N_28462,N_27274,N_26510);
and U28463 (N_28463,N_26353,N_26226);
and U28464 (N_28464,N_27293,N_26484);
nand U28465 (N_28465,N_26894,N_27816);
or U28466 (N_28466,N_27013,N_26784);
nor U28467 (N_28467,N_26433,N_26052);
nor U28468 (N_28468,N_27175,N_26325);
nand U28469 (N_28469,N_27100,N_27497);
and U28470 (N_28470,N_27919,N_27160);
and U28471 (N_28471,N_26389,N_27897);
nor U28472 (N_28472,N_27130,N_27103);
xor U28473 (N_28473,N_26152,N_26689);
or U28474 (N_28474,N_26660,N_26214);
nand U28475 (N_28475,N_26219,N_26046);
and U28476 (N_28476,N_26997,N_27526);
nand U28477 (N_28477,N_27877,N_26236);
xnor U28478 (N_28478,N_27708,N_27370);
and U28479 (N_28479,N_27852,N_27716);
or U28480 (N_28480,N_27619,N_26581);
nor U28481 (N_28481,N_26230,N_26276);
xnor U28482 (N_28482,N_27732,N_27026);
xor U28483 (N_28483,N_27319,N_27184);
or U28484 (N_28484,N_27920,N_26910);
or U28485 (N_28485,N_26680,N_26040);
xnor U28486 (N_28486,N_26696,N_26448);
xnor U28487 (N_28487,N_27908,N_27448);
nor U28488 (N_28488,N_26542,N_26398);
or U28489 (N_28489,N_27761,N_26729);
and U28490 (N_28490,N_26615,N_26412);
nor U28491 (N_28491,N_26920,N_27332);
and U28492 (N_28492,N_26227,N_27818);
or U28493 (N_28493,N_26089,N_27969);
and U28494 (N_28494,N_26038,N_27202);
and U28495 (N_28495,N_26179,N_26371);
nor U28496 (N_28496,N_27454,N_26279);
and U28497 (N_28497,N_27841,N_27651);
nand U28498 (N_28498,N_26823,N_27046);
nand U28499 (N_28499,N_27476,N_26180);
nand U28500 (N_28500,N_27356,N_27674);
nand U28501 (N_28501,N_26435,N_27813);
xor U28502 (N_28502,N_27461,N_26281);
nor U28503 (N_28503,N_26517,N_26700);
nand U28504 (N_28504,N_26685,N_26519);
or U28505 (N_28505,N_27769,N_27672);
nor U28506 (N_28506,N_27296,N_27817);
nand U28507 (N_28507,N_27860,N_26911);
nand U28508 (N_28508,N_27609,N_27836);
and U28509 (N_28509,N_27613,N_26317);
nor U28510 (N_28510,N_27081,N_26854);
or U28511 (N_28511,N_27252,N_26222);
and U28512 (N_28512,N_26762,N_26118);
and U28513 (N_28513,N_26408,N_27136);
and U28514 (N_28514,N_27399,N_26311);
xnor U28515 (N_28515,N_27098,N_27277);
xor U28516 (N_28516,N_26683,N_26340);
or U28517 (N_28517,N_26549,N_27596);
xnor U28518 (N_28518,N_27894,N_26322);
nor U28519 (N_28519,N_27007,N_27517);
nor U28520 (N_28520,N_27513,N_27000);
and U28521 (N_28521,N_26940,N_26441);
xor U28522 (N_28522,N_27346,N_27267);
or U28523 (N_28523,N_26860,N_27690);
xnor U28524 (N_28524,N_26528,N_26981);
and U28525 (N_28525,N_27133,N_27762);
xor U28526 (N_28526,N_27600,N_26066);
nand U28527 (N_28527,N_27372,N_27713);
and U28528 (N_28528,N_27796,N_27585);
xor U28529 (N_28529,N_27554,N_26314);
xnor U28530 (N_28530,N_27059,N_27015);
and U28531 (N_28531,N_26388,N_27400);
xor U28532 (N_28532,N_27886,N_26308);
nand U28533 (N_28533,N_26883,N_27604);
or U28534 (N_28534,N_26379,N_26312);
and U28535 (N_28535,N_27805,N_27804);
nor U28536 (N_28536,N_27384,N_27394);
nand U28537 (N_28537,N_27621,N_27649);
nor U28538 (N_28538,N_27347,N_26943);
and U28539 (N_28539,N_26345,N_26828);
and U28540 (N_28540,N_27149,N_27192);
xnor U28541 (N_28541,N_26659,N_26324);
xnor U28542 (N_28542,N_26492,N_26933);
and U28543 (N_28543,N_26234,N_26631);
nor U28544 (N_28544,N_26339,N_26201);
nand U28545 (N_28545,N_26019,N_27620);
nor U28546 (N_28546,N_26095,N_26892);
or U28547 (N_28547,N_26948,N_27756);
xor U28548 (N_28548,N_27719,N_26147);
nor U28549 (N_28549,N_27298,N_27547);
nor U28550 (N_28550,N_26257,N_27595);
xnor U28551 (N_28551,N_26084,N_26782);
nor U28552 (N_28552,N_27809,N_26788);
xor U28553 (N_28553,N_27611,N_26354);
and U28554 (N_28554,N_27973,N_26082);
or U28555 (N_28555,N_27022,N_26284);
xnor U28556 (N_28556,N_27140,N_26622);
nor U28557 (N_28557,N_27065,N_26509);
xor U28558 (N_28558,N_27080,N_26394);
and U28559 (N_28559,N_26901,N_26543);
xor U28560 (N_28560,N_26865,N_27124);
xnor U28561 (N_28561,N_27393,N_26292);
nor U28562 (N_28562,N_26937,N_27632);
xnor U28563 (N_28563,N_27176,N_27473);
nor U28564 (N_28564,N_26127,N_27760);
xor U28565 (N_28565,N_27294,N_26329);
or U28566 (N_28566,N_27838,N_27283);
xor U28567 (N_28567,N_27447,N_27861);
or U28568 (N_28568,N_27565,N_27736);
nand U28569 (N_28569,N_27376,N_26939);
nor U28570 (N_28570,N_26923,N_27191);
and U28571 (N_28571,N_26323,N_27960);
xnor U28572 (N_28572,N_27925,N_27330);
xnor U28573 (N_28573,N_27561,N_27967);
nor U28574 (N_28574,N_27183,N_26419);
nand U28575 (N_28575,N_26670,N_26909);
xnor U28576 (N_28576,N_26767,N_27405);
xnor U28577 (N_28577,N_27810,N_27091);
nor U28578 (N_28578,N_26607,N_26242);
nand U28579 (N_28579,N_26365,N_26698);
or U28580 (N_28580,N_27187,N_26870);
and U28581 (N_28581,N_27752,N_26789);
or U28582 (N_28582,N_27403,N_27630);
xor U28583 (N_28583,N_27377,N_27942);
nor U28584 (N_28584,N_27534,N_26146);
xnor U28585 (N_28585,N_26131,N_26378);
nand U28586 (N_28586,N_26836,N_27951);
and U28587 (N_28587,N_27679,N_26535);
nand U28588 (N_28588,N_26632,N_26693);
nor U28589 (N_28589,N_27800,N_27642);
and U28590 (N_28590,N_26775,N_26058);
xor U28591 (N_28591,N_27002,N_26211);
xnor U28592 (N_28592,N_26061,N_26703);
and U28593 (N_28593,N_26992,N_26812);
and U28594 (N_28594,N_26021,N_26863);
nor U28595 (N_28595,N_27102,N_26102);
nor U28596 (N_28596,N_27484,N_27626);
or U28597 (N_28597,N_27842,N_26451);
nor U28598 (N_28598,N_26132,N_27163);
nand U28599 (N_28599,N_27667,N_26391);
nand U28600 (N_28600,N_26444,N_26256);
nand U28601 (N_28601,N_27206,N_27174);
xnor U28602 (N_28602,N_26348,N_27815);
or U28603 (N_28603,N_26934,N_27231);
nor U28604 (N_28604,N_26774,N_26302);
nor U28605 (N_28605,N_27446,N_27019);
xnor U28606 (N_28606,N_26072,N_26455);
or U28607 (N_28607,N_26861,N_26914);
and U28608 (N_28608,N_27704,N_26547);
nor U28609 (N_28609,N_26194,N_27186);
nor U28610 (N_28610,N_26253,N_26316);
or U28611 (N_28611,N_27782,N_26395);
xnor U28612 (N_28612,N_27865,N_27122);
nand U28613 (N_28613,N_26740,N_26413);
nor U28614 (N_28614,N_27062,N_26165);
nor U28615 (N_28615,N_26054,N_27420);
nor U28616 (N_28616,N_27341,N_26765);
xor U28617 (N_28617,N_27374,N_26034);
nor U28618 (N_28618,N_26091,N_26174);
and U28619 (N_28619,N_26890,N_27264);
and U28620 (N_28620,N_27402,N_27216);
or U28621 (N_28621,N_27480,N_26873);
and U28622 (N_28622,N_27764,N_26286);
nor U28623 (N_28623,N_26278,N_27217);
nand U28624 (N_28624,N_27803,N_27439);
xnor U28625 (N_28625,N_26739,N_27410);
or U28626 (N_28626,N_27794,N_26439);
xnor U28627 (N_28627,N_26504,N_27110);
and U28628 (N_28628,N_26888,N_27941);
xor U28629 (N_28629,N_26374,N_27221);
or U28630 (N_28630,N_26707,N_27853);
or U28631 (N_28631,N_27444,N_26199);
nand U28632 (N_28632,N_27646,N_26952);
nand U28633 (N_28633,N_27562,N_27111);
nand U28634 (N_28634,N_27550,N_27313);
nor U28635 (N_28635,N_26891,N_26327);
nand U28636 (N_28636,N_27520,N_27105);
nor U28637 (N_28637,N_26833,N_26796);
or U28638 (N_28638,N_27900,N_26806);
nand U28639 (N_28639,N_27602,N_27851);
and U28640 (N_28640,N_27970,N_27870);
and U28641 (N_28641,N_27733,N_27006);
and U28642 (N_28642,N_26407,N_26626);
and U28643 (N_28643,N_26288,N_27248);
xnor U28644 (N_28644,N_26537,N_26176);
and U28645 (N_28645,N_27965,N_26431);
nor U28646 (N_28646,N_27018,N_26068);
xnor U28647 (N_28647,N_26144,N_26232);
and U28648 (N_28648,N_27415,N_27462);
nor U28649 (N_28649,N_27977,N_26220);
xnor U28650 (N_28650,N_27916,N_26857);
xor U28651 (N_28651,N_27771,N_26546);
xor U28652 (N_28652,N_26594,N_27164);
or U28653 (N_28653,N_27773,N_26155);
xnor U28654 (N_28654,N_26202,N_27159);
nand U28655 (N_28655,N_26512,N_27975);
nand U28656 (N_28656,N_26723,N_27802);
nor U28657 (N_28657,N_27011,N_26946);
nor U28658 (N_28658,N_27391,N_27855);
xnor U28659 (N_28659,N_27152,N_26773);
xor U28660 (N_28660,N_27044,N_26764);
xor U28661 (N_28661,N_26259,N_26566);
or U28662 (N_28662,N_27336,N_26469);
nor U28663 (N_28663,N_26347,N_27989);
or U28664 (N_28664,N_27037,N_26393);
nor U28665 (N_28665,N_27883,N_27675);
nor U28666 (N_28666,N_27781,N_26361);
nor U28667 (N_28667,N_27560,N_27746);
xnor U28668 (N_28668,N_27603,N_27814);
xor U28669 (N_28669,N_26531,N_26701);
xnor U28670 (N_28670,N_27957,N_27727);
nand U28671 (N_28671,N_26252,N_27524);
nand U28672 (N_28672,N_27839,N_27189);
or U28673 (N_28673,N_26669,N_26663);
or U28674 (N_28674,N_26472,N_26217);
nand U28675 (N_28675,N_26262,N_27297);
nand U28676 (N_28676,N_27455,N_26635);
nand U28677 (N_28677,N_26355,N_26582);
nor U28678 (N_28678,N_27999,N_26859);
nand U28679 (N_28679,N_27828,N_26945);
or U28680 (N_28680,N_26496,N_26713);
nand U28681 (N_28681,N_27398,N_27310);
nor U28682 (N_28682,N_26465,N_26094);
nand U28683 (N_28683,N_27695,N_27641);
nor U28684 (N_28684,N_26167,N_26477);
and U28685 (N_28685,N_27083,N_27859);
and U28686 (N_28686,N_27129,N_27940);
and U28687 (N_28687,N_26475,N_27212);
and U28688 (N_28688,N_27314,N_27572);
or U28689 (N_28689,N_27678,N_27553);
or U28690 (N_28690,N_27023,N_26516);
nand U28691 (N_28691,N_27178,N_26421);
nand U28692 (N_28692,N_27005,N_27515);
and U28693 (N_28693,N_27721,N_27445);
or U28694 (N_28694,N_26907,N_27119);
or U28695 (N_28695,N_27109,N_26124);
nor U28696 (N_28696,N_26295,N_26975);
nor U28697 (N_28697,N_27436,N_27197);
and U28698 (N_28698,N_27993,N_27684);
and U28699 (N_28699,N_26550,N_26260);
nor U28700 (N_28700,N_27063,N_27696);
or U28701 (N_28701,N_27361,N_26356);
nor U28702 (N_28702,N_26449,N_26954);
or U28703 (N_28703,N_27968,N_27788);
nand U28704 (N_28704,N_26041,N_27036);
nor U28705 (N_28705,N_27397,N_26984);
nand U28706 (N_28706,N_26986,N_26678);
nand U28707 (N_28707,N_26203,N_26032);
or U28708 (N_28708,N_27141,N_26752);
nand U28709 (N_28709,N_27067,N_26126);
xnor U28710 (N_28710,N_27872,N_27882);
xnor U28711 (N_28711,N_26009,N_26454);
and U28712 (N_28712,N_27300,N_26926);
xnor U28713 (N_28713,N_26715,N_27840);
nor U28714 (N_28714,N_26246,N_27507);
nor U28715 (N_28715,N_26827,N_26285);
xnor U28716 (N_28716,N_27066,N_26101);
xnor U28717 (N_28717,N_27483,N_26437);
or U28718 (N_28718,N_27355,N_26639);
and U28719 (N_28719,N_26462,N_26722);
xor U28720 (N_28720,N_27996,N_26574);
or U28721 (N_28721,N_26967,N_26881);
or U28722 (N_28722,N_26405,N_26445);
xnor U28723 (N_28723,N_27541,N_26110);
nand U28724 (N_28724,N_26661,N_27158);
xnor U28725 (N_28725,N_27144,N_26564);
xor U28726 (N_28726,N_27914,N_27095);
and U28727 (N_28727,N_26093,N_27693);
or U28728 (N_28728,N_26971,N_26684);
xor U28729 (N_28729,N_27837,N_27519);
or U28730 (N_28730,N_26758,N_26595);
nand U28731 (N_28731,N_27093,N_26487);
and U28732 (N_28732,N_26428,N_26273);
nor U28733 (N_28733,N_26800,N_26442);
xor U28734 (N_28734,N_26856,N_27854);
xor U28735 (N_28735,N_26904,N_27432);
nand U28736 (N_28736,N_26121,N_26915);
xor U28737 (N_28737,N_27964,N_27664);
nand U28738 (N_28738,N_27172,N_26640);
or U28739 (N_28739,N_26599,N_27650);
nand U28740 (N_28740,N_27481,N_27982);
nand U28741 (N_28741,N_27790,N_26461);
nand U28742 (N_28742,N_26111,N_27567);
nand U28743 (N_28743,N_27784,N_26741);
and U28744 (N_28744,N_27179,N_26037);
or U28745 (N_28745,N_26328,N_26357);
nor U28746 (N_28746,N_27349,N_27578);
and U28747 (N_28747,N_27783,N_26055);
xnor U28748 (N_28748,N_27959,N_27587);
nand U28749 (N_28749,N_26073,N_27426);
and U28750 (N_28750,N_26613,N_27656);
nor U28751 (N_28751,N_27369,N_26763);
or U28752 (N_28752,N_26529,N_27148);
xnor U28753 (N_28753,N_27757,N_26668);
and U28754 (N_28754,N_26012,N_27972);
or U28755 (N_28755,N_27418,N_27121);
and U28756 (N_28756,N_27953,N_26596);
or U28757 (N_28757,N_26718,N_26731);
xnor U28758 (N_28758,N_27640,N_26196);
and U28759 (N_28759,N_27012,N_26331);
nor U28760 (N_28760,N_27351,N_27423);
or U28761 (N_28761,N_26936,N_26646);
xor U28762 (N_28762,N_26973,N_26077);
and U28763 (N_28763,N_26597,N_26479);
nor U28764 (N_28764,N_26183,N_27786);
or U28765 (N_28765,N_27770,N_26778);
xnor U28766 (N_28766,N_27829,N_26570);
and U28767 (N_28767,N_26563,N_27893);
xor U28768 (N_28768,N_27717,N_26106);
nand U28769 (N_28769,N_26360,N_26839);
nand U28770 (N_28770,N_27710,N_27326);
nand U28771 (N_28771,N_26593,N_26652);
and U28772 (N_28772,N_26381,N_27904);
nand U28773 (N_28773,N_26006,N_27767);
nor U28774 (N_28774,N_27857,N_27210);
xor U28775 (N_28775,N_27407,N_27238);
nor U28776 (N_28776,N_26604,N_26313);
nand U28777 (N_28777,N_27628,N_27457);
nand U28778 (N_28778,N_27966,N_27629);
xnor U28779 (N_28779,N_27978,N_27139);
nand U28780 (N_28780,N_26423,N_26145);
or U28781 (N_28781,N_26096,N_26611);
xnor U28782 (N_28782,N_26238,N_27924);
nor U28783 (N_28783,N_26602,N_26838);
xnor U28784 (N_28784,N_27808,N_27416);
xor U28785 (N_28785,N_27662,N_26494);
and U28786 (N_28786,N_27499,N_27268);
nand U28787 (N_28787,N_26452,N_26380);
nand U28788 (N_28788,N_27094,N_27299);
nor U28789 (N_28789,N_27312,N_27568);
or U28790 (N_28790,N_27887,N_27806);
or U28791 (N_28791,N_26122,N_27823);
and U28792 (N_28792,N_26053,N_27261);
xnor U28793 (N_28793,N_26598,N_26825);
nor U28794 (N_28794,N_27616,N_27260);
nor U28795 (N_28795,N_27869,N_26961);
nor U28796 (N_28796,N_26070,N_27896);
nand U28797 (N_28797,N_26869,N_27085);
xor U28798 (N_28798,N_26738,N_26730);
nand U28799 (N_28799,N_26397,N_26960);
or U28800 (N_28800,N_26270,N_26505);
xnor U28801 (N_28801,N_26283,N_26855);
nand U28802 (N_28802,N_27700,N_26539);
nor U28803 (N_28803,N_27378,N_26436);
or U28804 (N_28804,N_26737,N_26588);
xnor U28805 (N_28805,N_26036,N_26569);
or U28806 (N_28806,N_27711,N_26966);
and U28807 (N_28807,N_27162,N_26187);
nor U28808 (N_28808,N_26198,N_26287);
xor U28809 (N_28809,N_27934,N_26235);
and U28810 (N_28810,N_27918,N_27639);
nor U28811 (N_28811,N_26493,N_26315);
xor U28812 (N_28812,N_27305,N_26277);
and U28813 (N_28813,N_27622,N_27812);
xnor U28814 (N_28814,N_27125,N_27844);
or U28815 (N_28815,N_26342,N_27510);
or U28816 (N_28816,N_26524,N_26989);
or U28817 (N_28817,N_27798,N_26612);
nor U28818 (N_28818,N_26010,N_27680);
or U28819 (N_28819,N_26086,N_27504);
xnor U28820 (N_28820,N_27588,N_27677);
nor U28821 (N_28821,N_26326,N_27906);
or U28822 (N_28822,N_27166,N_26573);
xnor U28823 (N_28823,N_26845,N_26821);
xor U28824 (N_28824,N_26672,N_26299);
and U28825 (N_28825,N_26790,N_26609);
and U28826 (N_28826,N_26168,N_27730);
or U28827 (N_28827,N_27644,N_26463);
xnor U28828 (N_28828,N_26123,N_27466);
and U28829 (N_28829,N_26366,N_27366);
or U28830 (N_28830,N_26275,N_26044);
and U28831 (N_28831,N_26592,N_27885);
xnor U28832 (N_28832,N_27021,N_26310);
xor U28833 (N_28833,N_26048,N_27281);
xor U28834 (N_28834,N_26476,N_26950);
nor U28835 (N_28835,N_27053,N_27888);
and U28836 (N_28836,N_26207,N_27031);
nor U28837 (N_28837,N_26795,N_26745);
xnor U28838 (N_28838,N_27506,N_26409);
and U28839 (N_28839,N_26491,N_26100);
nand U28840 (N_28840,N_26871,N_27518);
xor U28841 (N_28841,N_27135,N_26115);
and U28842 (N_28842,N_26350,N_27856);
xnor U28843 (N_28843,N_26733,N_27981);
nand U28844 (N_28844,N_27086,N_27049);
and U28845 (N_28845,N_26247,N_27482);
and U28846 (N_28846,N_27428,N_27108);
xnor U28847 (N_28847,N_27284,N_26928);
nor U28848 (N_28848,N_26802,N_27478);
or U28849 (N_28849,N_26440,N_26868);
nand U28850 (N_28850,N_27683,N_27255);
nand U28851 (N_28851,N_27850,N_26589);
xor U28852 (N_28852,N_27754,N_26385);
and U28853 (N_28853,N_26076,N_27905);
or U28854 (N_28854,N_26817,N_27427);
nor U28855 (N_28855,N_27625,N_27249);
or U28856 (N_28856,N_27498,N_26783);
nor U28857 (N_28857,N_26815,N_27525);
nor U28858 (N_28858,N_26759,N_26478);
xor U28859 (N_28859,N_27655,N_26050);
xnor U28860 (N_28860,N_27881,N_26297);
nand U28861 (N_28861,N_26303,N_27244);
and U28862 (N_28862,N_26525,N_26300);
and U28863 (N_28863,N_27097,N_27801);
nor U28864 (N_28864,N_27623,N_27903);
or U28865 (N_28865,N_27259,N_27530);
nand U28866 (N_28866,N_26417,N_27440);
or U28867 (N_28867,N_27714,N_26608);
and U28868 (N_28868,N_27421,N_27845);
and U28869 (N_28869,N_26876,N_26727);
nand U28870 (N_28870,N_26208,N_26862);
nor U28871 (N_28871,N_27532,N_27318);
and U28872 (N_28872,N_27068,N_26092);
nor U28873 (N_28873,N_27278,N_26742);
or U28874 (N_28874,N_26905,N_27980);
nor U28875 (N_28875,N_27014,N_27971);
xnor U28876 (N_28876,N_26330,N_26571);
or U28877 (N_28877,N_27027,N_26319);
nand U28878 (N_28878,N_26653,N_27467);
and U28879 (N_28879,N_27389,N_26918);
and U28880 (N_28880,N_27624,N_26138);
xor U28881 (N_28881,N_27364,N_26223);
or U28882 (N_28882,N_27055,N_27226);
nand U28883 (N_28883,N_26710,N_26706);
nor U28884 (N_28884,N_26708,N_27531);
or U28885 (N_28885,N_26749,N_26980);
xor U28886 (N_28886,N_26074,N_26422);
xor U28887 (N_28887,N_26664,N_26616);
nor U28888 (N_28888,N_27032,N_26726);
nand U28889 (N_28889,N_26447,N_27988);
and U28890 (N_28890,N_27636,N_26902);
or U28891 (N_28891,N_26644,N_26097);
or U28892 (N_28892,N_26261,N_26290);
and U28893 (N_28893,N_27871,N_27290);
xor U28894 (N_28894,N_27375,N_27142);
and U28895 (N_28895,N_26047,N_26908);
xnor U28896 (N_28896,N_26030,N_27926);
or U28897 (N_28897,N_27707,N_26606);
and U28898 (N_28898,N_27161,N_26642);
nor U28899 (N_28899,N_26590,N_26399);
and U28900 (N_28900,N_27041,N_26753);
or U28901 (N_28901,N_27564,N_26637);
nor U28902 (N_28902,N_27583,N_26852);
xor U28903 (N_28903,N_26057,N_26269);
and U28904 (N_28904,N_27846,N_26877);
and U28905 (N_28905,N_26289,N_26043);
nand U28906 (N_28906,N_26107,N_27242);
and U28907 (N_28907,N_26164,N_27849);
nor U28908 (N_28908,N_27061,N_26734);
nor U28909 (N_28909,N_27234,N_27472);
nor U28910 (N_28910,N_26676,N_26947);
or U28911 (N_28911,N_26088,N_27078);
nor U28912 (N_28912,N_27051,N_27151);
xnor U28913 (N_28913,N_27660,N_27938);
and U28914 (N_28914,N_26045,N_26210);
nand U28915 (N_28915,N_26148,N_27199);
or U28916 (N_28916,N_26679,N_27997);
or U28917 (N_28917,N_26567,N_27584);
nand U28918 (N_28918,N_27698,N_26473);
or U28919 (N_28919,N_26809,N_26511);
nor U28920 (N_28920,N_27580,N_26630);
and U28921 (N_28921,N_26732,N_27379);
nand U28922 (N_28922,N_27243,N_26938);
nor U28923 (N_28923,N_27983,N_26794);
and U28924 (N_28924,N_26814,N_26551);
or U28925 (N_28925,N_27257,N_26579);
and U28926 (N_28926,N_27955,N_26922);
xor U28927 (N_28927,N_27927,N_27943);
or U28928 (N_28928,N_26443,N_27251);
or U28929 (N_28929,N_26526,N_26671);
nor U28930 (N_28930,N_27546,N_26489);
or U28931 (N_28931,N_27450,N_26982);
or U28932 (N_28932,N_26390,N_27895);
and U28933 (N_28933,N_27689,N_27246);
nand U28934 (N_28934,N_26157,N_26842);
xor U28935 (N_28935,N_26643,N_27995);
nand U28936 (N_28936,N_27948,N_27034);
nand U28937 (N_28937,N_26192,N_27787);
nor U28938 (N_28938,N_26924,N_26956);
and U28939 (N_28939,N_27468,N_26156);
or U28940 (N_28940,N_27411,N_26267);
or U28941 (N_28941,N_26674,N_26346);
nor U28942 (N_28942,N_26651,N_26820);
nand U28943 (N_28943,N_26994,N_27262);
nand U28944 (N_28944,N_27117,N_26916);
and U28945 (N_28945,N_26886,N_27772);
nand U28946 (N_28946,N_26755,N_26384);
or U28947 (N_28947,N_26756,N_26927);
xnor U28948 (N_28948,N_27505,N_27551);
xnor U28949 (N_28949,N_26754,N_26178);
xnor U28950 (N_28950,N_27396,N_27043);
nand U28951 (N_28951,N_26466,N_27768);
or U28952 (N_28952,N_26231,N_27647);
nand U28953 (N_28953,N_27929,N_26785);
nand U28954 (N_28954,N_26851,N_27738);
xnor U28955 (N_28955,N_27171,N_26649);
or U28956 (N_28956,N_26650,N_26747);
nor U28957 (N_28957,N_27456,N_27301);
xnor U28958 (N_28958,N_26832,N_27935);
nand U28959 (N_28959,N_26751,N_26826);
nand U28960 (N_28960,N_26750,N_26899);
xnor U28961 (N_28961,N_26020,N_27348);
xor U28962 (N_28962,N_26831,N_26627);
and U28963 (N_28963,N_26560,N_26620);
nand U28964 (N_28964,N_27222,N_26887);
xor U28965 (N_28965,N_27686,N_26963);
or U28966 (N_28966,N_26878,N_27880);
nor U28967 (N_28967,N_27285,N_27601);
nor U28968 (N_28968,N_26665,N_26373);
nand U28969 (N_28969,N_27443,N_26893);
nor U28970 (N_28970,N_26206,N_26819);
nor U28971 (N_28971,N_27931,N_26161);
and U28972 (N_28972,N_26375,N_27822);
or U28973 (N_28973,N_26026,N_27486);
xnor U28974 (N_28974,N_27433,N_27673);
nand U28975 (N_28975,N_26481,N_26666);
and U28976 (N_28976,N_27891,N_26486);
nor U28977 (N_28977,N_27819,N_26957);
or U28978 (N_28978,N_27417,N_27990);
or U28979 (N_28979,N_27939,N_27422);
and U28980 (N_28980,N_27627,N_26416);
xnor U28981 (N_28981,N_26301,N_26654);
or U28982 (N_28982,N_27076,N_26485);
nor U28983 (N_28983,N_27665,N_27165);
xnor U28984 (N_28984,N_27791,N_26483);
xor U28985 (N_28985,N_26555,N_26843);
and U28986 (N_28986,N_27661,N_27610);
or U28987 (N_28987,N_26565,N_27029);
nor U28988 (N_28988,N_27991,N_27196);
and U28989 (N_28989,N_27614,N_27638);
and U28990 (N_28990,N_27946,N_27344);
nand U28991 (N_28991,N_26467,N_27048);
xor U28992 (N_28992,N_27509,N_26268);
or U28993 (N_28993,N_26112,N_26335);
nor U28994 (N_28994,N_26880,N_26078);
and U28995 (N_28995,N_27576,N_27424);
or U28996 (N_28996,N_26987,N_27612);
and U28997 (N_28997,N_27170,N_27235);
nor U28998 (N_28998,N_26059,N_27493);
xor U28999 (N_28999,N_27848,N_27494);
xor U29000 (N_29000,N_26801,N_26480);
xor U29001 (N_29001,N_27275,N_27775);
xor U29002 (N_29002,N_27117,N_27725);
and U29003 (N_29003,N_26552,N_27887);
xnor U29004 (N_29004,N_26708,N_26363);
and U29005 (N_29005,N_26015,N_27131);
and U29006 (N_29006,N_27222,N_26041);
nand U29007 (N_29007,N_27431,N_27107);
and U29008 (N_29008,N_26485,N_27154);
nand U29009 (N_29009,N_27836,N_27146);
nor U29010 (N_29010,N_26191,N_27257);
or U29011 (N_29011,N_26033,N_27356);
nor U29012 (N_29012,N_27971,N_27351);
nand U29013 (N_29013,N_27784,N_26135);
and U29014 (N_29014,N_27838,N_26824);
and U29015 (N_29015,N_27750,N_27025);
nand U29016 (N_29016,N_26927,N_26975);
and U29017 (N_29017,N_27330,N_26269);
nor U29018 (N_29018,N_26751,N_26582);
and U29019 (N_29019,N_26026,N_26952);
or U29020 (N_29020,N_27462,N_27673);
nand U29021 (N_29021,N_26919,N_26144);
and U29022 (N_29022,N_26011,N_26255);
or U29023 (N_29023,N_27686,N_27084);
nand U29024 (N_29024,N_26667,N_27560);
nand U29025 (N_29025,N_26342,N_26899);
and U29026 (N_29026,N_27255,N_26644);
or U29027 (N_29027,N_26495,N_26617);
and U29028 (N_29028,N_27510,N_27281);
nand U29029 (N_29029,N_27961,N_27178);
and U29030 (N_29030,N_27362,N_27916);
nand U29031 (N_29031,N_27146,N_27243);
xor U29032 (N_29032,N_26487,N_27467);
or U29033 (N_29033,N_26153,N_27150);
and U29034 (N_29034,N_27251,N_27802);
nor U29035 (N_29035,N_26164,N_27754);
and U29036 (N_29036,N_26015,N_26483);
xnor U29037 (N_29037,N_26575,N_27336);
nand U29038 (N_29038,N_26009,N_26610);
nor U29039 (N_29039,N_27199,N_27406);
and U29040 (N_29040,N_27340,N_26822);
nand U29041 (N_29041,N_26890,N_26033);
nand U29042 (N_29042,N_27872,N_27414);
and U29043 (N_29043,N_27718,N_27055);
or U29044 (N_29044,N_27494,N_26548);
nand U29045 (N_29045,N_27290,N_26689);
nand U29046 (N_29046,N_26778,N_26176);
nand U29047 (N_29047,N_26851,N_26575);
nand U29048 (N_29048,N_26502,N_27988);
and U29049 (N_29049,N_26872,N_26600);
xor U29050 (N_29050,N_27760,N_27012);
or U29051 (N_29051,N_26265,N_27916);
and U29052 (N_29052,N_27723,N_26897);
xor U29053 (N_29053,N_26805,N_27648);
nand U29054 (N_29054,N_26539,N_26818);
or U29055 (N_29055,N_26970,N_27580);
or U29056 (N_29056,N_26933,N_27190);
or U29057 (N_29057,N_27944,N_26670);
or U29058 (N_29058,N_26789,N_27875);
xnor U29059 (N_29059,N_26570,N_27858);
nand U29060 (N_29060,N_27993,N_27562);
nor U29061 (N_29061,N_27510,N_26979);
and U29062 (N_29062,N_27291,N_26498);
xor U29063 (N_29063,N_26553,N_26525);
xor U29064 (N_29064,N_26276,N_27653);
nand U29065 (N_29065,N_26297,N_27806);
xnor U29066 (N_29066,N_27943,N_26860);
or U29067 (N_29067,N_27095,N_27088);
nor U29068 (N_29068,N_27126,N_27122);
or U29069 (N_29069,N_26645,N_26785);
nand U29070 (N_29070,N_27299,N_26278);
and U29071 (N_29071,N_26697,N_26033);
and U29072 (N_29072,N_26580,N_26196);
xnor U29073 (N_29073,N_26321,N_26864);
nand U29074 (N_29074,N_27864,N_27382);
nor U29075 (N_29075,N_27914,N_26500);
and U29076 (N_29076,N_27554,N_27727);
xor U29077 (N_29077,N_26672,N_26800);
and U29078 (N_29078,N_27238,N_26900);
nand U29079 (N_29079,N_26399,N_26640);
nor U29080 (N_29080,N_26376,N_26713);
xnor U29081 (N_29081,N_27244,N_26813);
or U29082 (N_29082,N_27416,N_27199);
and U29083 (N_29083,N_26048,N_27644);
xnor U29084 (N_29084,N_26085,N_26691);
or U29085 (N_29085,N_26861,N_27565);
nor U29086 (N_29086,N_26573,N_27227);
or U29087 (N_29087,N_26620,N_26009);
nand U29088 (N_29088,N_26785,N_27902);
xnor U29089 (N_29089,N_26802,N_27337);
nand U29090 (N_29090,N_27633,N_27318);
nor U29091 (N_29091,N_27797,N_26572);
or U29092 (N_29092,N_26912,N_27272);
nand U29093 (N_29093,N_27379,N_27565);
nand U29094 (N_29094,N_26520,N_27189);
nor U29095 (N_29095,N_26094,N_26916);
or U29096 (N_29096,N_27935,N_27617);
or U29097 (N_29097,N_27886,N_27525);
nand U29098 (N_29098,N_26912,N_26835);
nor U29099 (N_29099,N_26504,N_26310);
or U29100 (N_29100,N_27662,N_26649);
and U29101 (N_29101,N_27287,N_26465);
or U29102 (N_29102,N_27641,N_27877);
xnor U29103 (N_29103,N_26884,N_26268);
nand U29104 (N_29104,N_26509,N_27662);
nor U29105 (N_29105,N_27169,N_26696);
xor U29106 (N_29106,N_27135,N_26582);
or U29107 (N_29107,N_27740,N_27103);
or U29108 (N_29108,N_26600,N_26725);
xnor U29109 (N_29109,N_27999,N_26189);
or U29110 (N_29110,N_26545,N_26090);
nor U29111 (N_29111,N_26023,N_27075);
xnor U29112 (N_29112,N_27777,N_27374);
nand U29113 (N_29113,N_27098,N_26825);
nor U29114 (N_29114,N_27488,N_27216);
or U29115 (N_29115,N_26263,N_27456);
xnor U29116 (N_29116,N_26378,N_27610);
and U29117 (N_29117,N_27089,N_27837);
nor U29118 (N_29118,N_27203,N_26568);
or U29119 (N_29119,N_27526,N_27033);
nand U29120 (N_29120,N_27837,N_27090);
nand U29121 (N_29121,N_26824,N_26862);
or U29122 (N_29122,N_26443,N_26775);
nand U29123 (N_29123,N_27013,N_26161);
xor U29124 (N_29124,N_27382,N_27419);
or U29125 (N_29125,N_27477,N_27128);
nand U29126 (N_29126,N_27484,N_26304);
nand U29127 (N_29127,N_26858,N_26397);
xor U29128 (N_29128,N_27667,N_26897);
and U29129 (N_29129,N_27457,N_26718);
nor U29130 (N_29130,N_26670,N_26224);
nor U29131 (N_29131,N_27271,N_27710);
xnor U29132 (N_29132,N_26788,N_26770);
and U29133 (N_29133,N_27723,N_26952);
and U29134 (N_29134,N_27861,N_26952);
and U29135 (N_29135,N_27893,N_27292);
xnor U29136 (N_29136,N_27531,N_27955);
nand U29137 (N_29137,N_27888,N_26060);
xnor U29138 (N_29138,N_27713,N_27174);
xnor U29139 (N_29139,N_27694,N_26129);
xor U29140 (N_29140,N_26190,N_26314);
nand U29141 (N_29141,N_26738,N_26013);
nand U29142 (N_29142,N_27704,N_27410);
nand U29143 (N_29143,N_26975,N_27737);
xnor U29144 (N_29144,N_27254,N_27193);
nor U29145 (N_29145,N_27955,N_26748);
or U29146 (N_29146,N_27083,N_26905);
and U29147 (N_29147,N_26519,N_26788);
and U29148 (N_29148,N_26222,N_26120);
xor U29149 (N_29149,N_26871,N_26508);
xor U29150 (N_29150,N_27487,N_27700);
nand U29151 (N_29151,N_27792,N_26475);
xnor U29152 (N_29152,N_26563,N_26931);
or U29153 (N_29153,N_26077,N_27942);
or U29154 (N_29154,N_26065,N_26186);
nand U29155 (N_29155,N_27460,N_26024);
xor U29156 (N_29156,N_27208,N_26685);
xnor U29157 (N_29157,N_27003,N_27504);
and U29158 (N_29158,N_27343,N_27238);
xnor U29159 (N_29159,N_27363,N_27786);
nor U29160 (N_29160,N_26549,N_27507);
xor U29161 (N_29161,N_27414,N_27867);
nand U29162 (N_29162,N_26637,N_26519);
nand U29163 (N_29163,N_26201,N_26696);
or U29164 (N_29164,N_27737,N_27367);
nand U29165 (N_29165,N_27204,N_26564);
or U29166 (N_29166,N_27425,N_26779);
xor U29167 (N_29167,N_26263,N_26369);
nand U29168 (N_29168,N_27943,N_27860);
and U29169 (N_29169,N_26462,N_27165);
xor U29170 (N_29170,N_27091,N_26495);
nor U29171 (N_29171,N_26438,N_27964);
nor U29172 (N_29172,N_26083,N_26155);
or U29173 (N_29173,N_27683,N_26047);
xor U29174 (N_29174,N_27879,N_27324);
nor U29175 (N_29175,N_27009,N_27270);
nand U29176 (N_29176,N_26538,N_27192);
nor U29177 (N_29177,N_26312,N_27459);
and U29178 (N_29178,N_27763,N_26901);
nand U29179 (N_29179,N_27788,N_27158);
and U29180 (N_29180,N_27239,N_26630);
or U29181 (N_29181,N_26862,N_26910);
or U29182 (N_29182,N_26259,N_27395);
or U29183 (N_29183,N_27217,N_27820);
nand U29184 (N_29184,N_26534,N_27239);
xnor U29185 (N_29185,N_26848,N_27585);
nand U29186 (N_29186,N_27775,N_26204);
nand U29187 (N_29187,N_26119,N_26155);
nor U29188 (N_29188,N_27592,N_27588);
nand U29189 (N_29189,N_26417,N_27564);
or U29190 (N_29190,N_27079,N_27509);
nor U29191 (N_29191,N_27272,N_27309);
nor U29192 (N_29192,N_27252,N_27339);
xnor U29193 (N_29193,N_26071,N_27438);
nor U29194 (N_29194,N_27265,N_27348);
or U29195 (N_29195,N_27667,N_27934);
nor U29196 (N_29196,N_26500,N_27507);
xor U29197 (N_29197,N_26104,N_27382);
or U29198 (N_29198,N_26229,N_27069);
and U29199 (N_29199,N_27900,N_27806);
nand U29200 (N_29200,N_26363,N_27611);
xnor U29201 (N_29201,N_27486,N_26040);
nand U29202 (N_29202,N_27037,N_27346);
xor U29203 (N_29203,N_26900,N_26089);
nor U29204 (N_29204,N_26221,N_26644);
or U29205 (N_29205,N_27263,N_27240);
xnor U29206 (N_29206,N_27631,N_27572);
nand U29207 (N_29207,N_26597,N_26971);
nor U29208 (N_29208,N_26530,N_27611);
nor U29209 (N_29209,N_26416,N_27437);
and U29210 (N_29210,N_27299,N_27895);
and U29211 (N_29211,N_27467,N_26591);
nor U29212 (N_29212,N_26639,N_26928);
nand U29213 (N_29213,N_26633,N_27857);
xor U29214 (N_29214,N_27492,N_26278);
and U29215 (N_29215,N_27229,N_27451);
or U29216 (N_29216,N_27337,N_27272);
nor U29217 (N_29217,N_27541,N_27766);
or U29218 (N_29218,N_26009,N_26471);
or U29219 (N_29219,N_26577,N_26105);
and U29220 (N_29220,N_26367,N_27843);
and U29221 (N_29221,N_26140,N_27438);
or U29222 (N_29222,N_27960,N_27210);
nor U29223 (N_29223,N_26410,N_26054);
xnor U29224 (N_29224,N_27360,N_27884);
and U29225 (N_29225,N_27380,N_26879);
nor U29226 (N_29226,N_27821,N_26561);
nor U29227 (N_29227,N_27947,N_27839);
xnor U29228 (N_29228,N_26021,N_26529);
nor U29229 (N_29229,N_27507,N_26755);
and U29230 (N_29230,N_26169,N_26045);
or U29231 (N_29231,N_27241,N_26051);
nor U29232 (N_29232,N_26777,N_26371);
xnor U29233 (N_29233,N_27566,N_27241);
xor U29234 (N_29234,N_26281,N_26203);
xor U29235 (N_29235,N_27328,N_27194);
and U29236 (N_29236,N_27035,N_26171);
nor U29237 (N_29237,N_26200,N_26906);
nand U29238 (N_29238,N_27226,N_26431);
xor U29239 (N_29239,N_26335,N_27544);
nand U29240 (N_29240,N_27402,N_27417);
or U29241 (N_29241,N_27075,N_27303);
xnor U29242 (N_29242,N_27181,N_27258);
nand U29243 (N_29243,N_26762,N_26176);
xor U29244 (N_29244,N_26773,N_26215);
or U29245 (N_29245,N_27717,N_26243);
or U29246 (N_29246,N_27642,N_26029);
xor U29247 (N_29247,N_27229,N_26333);
xnor U29248 (N_29248,N_27051,N_26156);
nor U29249 (N_29249,N_26893,N_27876);
nand U29250 (N_29250,N_27422,N_26307);
xor U29251 (N_29251,N_27035,N_26100);
xor U29252 (N_29252,N_26917,N_27898);
nor U29253 (N_29253,N_27649,N_27193);
and U29254 (N_29254,N_27416,N_27674);
xor U29255 (N_29255,N_26971,N_27943);
or U29256 (N_29256,N_26293,N_27027);
nand U29257 (N_29257,N_26732,N_26714);
xor U29258 (N_29258,N_27492,N_26820);
nand U29259 (N_29259,N_26695,N_26983);
or U29260 (N_29260,N_26676,N_27096);
nand U29261 (N_29261,N_26141,N_27048);
xnor U29262 (N_29262,N_26997,N_27880);
xor U29263 (N_29263,N_26250,N_26365);
nor U29264 (N_29264,N_27693,N_27416);
or U29265 (N_29265,N_27935,N_27091);
or U29266 (N_29266,N_27985,N_26894);
nand U29267 (N_29267,N_27021,N_26041);
and U29268 (N_29268,N_26272,N_27631);
or U29269 (N_29269,N_27559,N_27740);
and U29270 (N_29270,N_26083,N_26792);
and U29271 (N_29271,N_27529,N_26052);
and U29272 (N_29272,N_27146,N_27478);
xor U29273 (N_29273,N_26644,N_26560);
xor U29274 (N_29274,N_27776,N_26192);
nand U29275 (N_29275,N_27897,N_26256);
nor U29276 (N_29276,N_27611,N_27661);
and U29277 (N_29277,N_26663,N_26226);
or U29278 (N_29278,N_27215,N_26355);
and U29279 (N_29279,N_26272,N_27197);
nor U29280 (N_29280,N_26109,N_27592);
and U29281 (N_29281,N_26399,N_26414);
xnor U29282 (N_29282,N_26024,N_27951);
xor U29283 (N_29283,N_27764,N_26287);
and U29284 (N_29284,N_26609,N_27559);
nor U29285 (N_29285,N_27310,N_27788);
or U29286 (N_29286,N_26800,N_26474);
xor U29287 (N_29287,N_26004,N_27880);
and U29288 (N_29288,N_26369,N_26761);
and U29289 (N_29289,N_26283,N_27280);
nor U29290 (N_29290,N_26674,N_26266);
or U29291 (N_29291,N_26846,N_26908);
nor U29292 (N_29292,N_27450,N_26430);
or U29293 (N_29293,N_26775,N_26835);
nand U29294 (N_29294,N_27347,N_27415);
xnor U29295 (N_29295,N_26725,N_26801);
nand U29296 (N_29296,N_27179,N_26763);
nor U29297 (N_29297,N_27618,N_26142);
nand U29298 (N_29298,N_26092,N_27543);
and U29299 (N_29299,N_27235,N_26316);
xnor U29300 (N_29300,N_26016,N_26731);
nand U29301 (N_29301,N_26476,N_27531);
nor U29302 (N_29302,N_26773,N_27460);
nand U29303 (N_29303,N_27311,N_26949);
xor U29304 (N_29304,N_27153,N_26800);
nor U29305 (N_29305,N_27097,N_26823);
or U29306 (N_29306,N_26107,N_26845);
and U29307 (N_29307,N_26662,N_27731);
and U29308 (N_29308,N_27255,N_26715);
nor U29309 (N_29309,N_26393,N_27205);
nor U29310 (N_29310,N_27135,N_26621);
xor U29311 (N_29311,N_26165,N_27038);
or U29312 (N_29312,N_26923,N_27417);
xor U29313 (N_29313,N_26980,N_26423);
xor U29314 (N_29314,N_27310,N_27326);
and U29315 (N_29315,N_26048,N_27881);
xor U29316 (N_29316,N_27318,N_26373);
and U29317 (N_29317,N_26754,N_27061);
xor U29318 (N_29318,N_27820,N_26011);
nor U29319 (N_29319,N_27470,N_26211);
or U29320 (N_29320,N_26574,N_27181);
nand U29321 (N_29321,N_26696,N_27209);
or U29322 (N_29322,N_26627,N_26743);
or U29323 (N_29323,N_26309,N_26154);
nand U29324 (N_29324,N_27306,N_26831);
nor U29325 (N_29325,N_26946,N_27847);
and U29326 (N_29326,N_26121,N_27348);
xnor U29327 (N_29327,N_27354,N_26803);
nand U29328 (N_29328,N_27753,N_27649);
or U29329 (N_29329,N_27748,N_26509);
or U29330 (N_29330,N_26929,N_26998);
nor U29331 (N_29331,N_27030,N_27421);
or U29332 (N_29332,N_26317,N_26942);
nand U29333 (N_29333,N_27151,N_26824);
nand U29334 (N_29334,N_27416,N_26213);
and U29335 (N_29335,N_27700,N_27401);
and U29336 (N_29336,N_26444,N_27520);
xor U29337 (N_29337,N_27545,N_26274);
nand U29338 (N_29338,N_27293,N_27200);
or U29339 (N_29339,N_27350,N_26683);
nand U29340 (N_29340,N_27205,N_26864);
nor U29341 (N_29341,N_27911,N_26372);
nor U29342 (N_29342,N_26867,N_26389);
nor U29343 (N_29343,N_26221,N_26692);
nor U29344 (N_29344,N_26258,N_27559);
and U29345 (N_29345,N_27639,N_27039);
xor U29346 (N_29346,N_26727,N_27278);
and U29347 (N_29347,N_26210,N_27215);
xor U29348 (N_29348,N_26838,N_26025);
nand U29349 (N_29349,N_26169,N_27767);
nor U29350 (N_29350,N_27874,N_26235);
or U29351 (N_29351,N_26488,N_27832);
nor U29352 (N_29352,N_27708,N_26588);
and U29353 (N_29353,N_27960,N_26170);
xor U29354 (N_29354,N_26798,N_27125);
nand U29355 (N_29355,N_27785,N_27872);
xor U29356 (N_29356,N_27416,N_27646);
or U29357 (N_29357,N_27449,N_27210);
or U29358 (N_29358,N_26894,N_27801);
and U29359 (N_29359,N_26250,N_27819);
nor U29360 (N_29360,N_26103,N_27197);
or U29361 (N_29361,N_27611,N_26024);
xor U29362 (N_29362,N_27127,N_27118);
and U29363 (N_29363,N_27100,N_26841);
nand U29364 (N_29364,N_26714,N_26954);
nand U29365 (N_29365,N_27101,N_26101);
nor U29366 (N_29366,N_26882,N_27948);
xor U29367 (N_29367,N_26733,N_26978);
nor U29368 (N_29368,N_26799,N_26579);
nor U29369 (N_29369,N_26383,N_27900);
nand U29370 (N_29370,N_27418,N_26576);
nor U29371 (N_29371,N_27082,N_27946);
nor U29372 (N_29372,N_27660,N_26997);
xor U29373 (N_29373,N_27978,N_26102);
xor U29374 (N_29374,N_26289,N_27945);
nand U29375 (N_29375,N_27426,N_27012);
nand U29376 (N_29376,N_27110,N_26790);
nor U29377 (N_29377,N_26642,N_27143);
xor U29378 (N_29378,N_26531,N_26792);
nand U29379 (N_29379,N_26699,N_27278);
or U29380 (N_29380,N_27282,N_26597);
nand U29381 (N_29381,N_26489,N_27570);
or U29382 (N_29382,N_27280,N_27131);
or U29383 (N_29383,N_27548,N_27682);
nand U29384 (N_29384,N_26740,N_27111);
nand U29385 (N_29385,N_27528,N_26572);
and U29386 (N_29386,N_27857,N_27861);
nand U29387 (N_29387,N_26357,N_26347);
or U29388 (N_29388,N_27384,N_27835);
and U29389 (N_29389,N_26060,N_27842);
or U29390 (N_29390,N_27834,N_26665);
xnor U29391 (N_29391,N_27522,N_26542);
nor U29392 (N_29392,N_26580,N_26797);
nor U29393 (N_29393,N_26557,N_26342);
nor U29394 (N_29394,N_27391,N_26584);
nand U29395 (N_29395,N_27422,N_26343);
nand U29396 (N_29396,N_27824,N_26585);
xor U29397 (N_29397,N_26841,N_27411);
or U29398 (N_29398,N_26966,N_27305);
or U29399 (N_29399,N_27034,N_26017);
nand U29400 (N_29400,N_27722,N_26757);
or U29401 (N_29401,N_27004,N_27016);
nand U29402 (N_29402,N_26136,N_27654);
nand U29403 (N_29403,N_26804,N_26645);
and U29404 (N_29404,N_27692,N_27958);
xnor U29405 (N_29405,N_26788,N_26634);
nand U29406 (N_29406,N_26859,N_26915);
or U29407 (N_29407,N_27579,N_27453);
and U29408 (N_29408,N_27883,N_26840);
nor U29409 (N_29409,N_27223,N_27000);
nand U29410 (N_29410,N_27704,N_27375);
xor U29411 (N_29411,N_26505,N_26481);
nand U29412 (N_29412,N_27961,N_27472);
nand U29413 (N_29413,N_26794,N_27114);
xnor U29414 (N_29414,N_26725,N_26249);
xor U29415 (N_29415,N_26619,N_27416);
and U29416 (N_29416,N_27788,N_26881);
and U29417 (N_29417,N_26111,N_27118);
nor U29418 (N_29418,N_27233,N_26170);
or U29419 (N_29419,N_27040,N_26553);
xnor U29420 (N_29420,N_27814,N_27601);
or U29421 (N_29421,N_27053,N_26662);
nor U29422 (N_29422,N_27652,N_26854);
nor U29423 (N_29423,N_27217,N_27763);
or U29424 (N_29424,N_27656,N_26382);
or U29425 (N_29425,N_26325,N_26642);
xnor U29426 (N_29426,N_26937,N_27296);
and U29427 (N_29427,N_26500,N_26431);
and U29428 (N_29428,N_26019,N_27538);
nor U29429 (N_29429,N_26221,N_27370);
nand U29430 (N_29430,N_26326,N_26840);
nor U29431 (N_29431,N_27039,N_27362);
xnor U29432 (N_29432,N_26371,N_27379);
and U29433 (N_29433,N_26234,N_26642);
xnor U29434 (N_29434,N_26726,N_26605);
nor U29435 (N_29435,N_27382,N_26565);
xnor U29436 (N_29436,N_26413,N_27321);
nor U29437 (N_29437,N_27673,N_26327);
or U29438 (N_29438,N_27622,N_27217);
nand U29439 (N_29439,N_27620,N_27670);
xor U29440 (N_29440,N_27918,N_27186);
nand U29441 (N_29441,N_26825,N_26354);
nor U29442 (N_29442,N_27858,N_27207);
nand U29443 (N_29443,N_26348,N_26538);
nor U29444 (N_29444,N_27097,N_26593);
or U29445 (N_29445,N_26290,N_26674);
xnor U29446 (N_29446,N_26152,N_27514);
nand U29447 (N_29447,N_27130,N_26443);
and U29448 (N_29448,N_26107,N_26803);
xnor U29449 (N_29449,N_27491,N_26743);
nor U29450 (N_29450,N_27269,N_26021);
nand U29451 (N_29451,N_27698,N_27435);
xor U29452 (N_29452,N_27720,N_27332);
xor U29453 (N_29453,N_27476,N_27222);
nand U29454 (N_29454,N_26583,N_27688);
or U29455 (N_29455,N_27686,N_26409);
or U29456 (N_29456,N_26300,N_26882);
nor U29457 (N_29457,N_26082,N_27710);
xnor U29458 (N_29458,N_26307,N_26194);
xor U29459 (N_29459,N_26604,N_26102);
nor U29460 (N_29460,N_26636,N_27871);
and U29461 (N_29461,N_26714,N_26979);
or U29462 (N_29462,N_27805,N_27213);
nor U29463 (N_29463,N_27931,N_26801);
or U29464 (N_29464,N_26590,N_27047);
xnor U29465 (N_29465,N_26080,N_26944);
or U29466 (N_29466,N_27771,N_26187);
or U29467 (N_29467,N_26276,N_27231);
nand U29468 (N_29468,N_26262,N_27861);
xnor U29469 (N_29469,N_26136,N_27540);
nor U29470 (N_29470,N_26908,N_26038);
xor U29471 (N_29471,N_27123,N_26248);
or U29472 (N_29472,N_26098,N_26564);
xor U29473 (N_29473,N_26919,N_27647);
xnor U29474 (N_29474,N_27785,N_26340);
xor U29475 (N_29475,N_26231,N_26639);
nand U29476 (N_29476,N_26871,N_27527);
and U29477 (N_29477,N_26916,N_26938);
xnor U29478 (N_29478,N_27126,N_27294);
xor U29479 (N_29479,N_26198,N_27998);
nor U29480 (N_29480,N_26557,N_27176);
nor U29481 (N_29481,N_26315,N_26921);
xor U29482 (N_29482,N_26945,N_27367);
nand U29483 (N_29483,N_26942,N_26614);
and U29484 (N_29484,N_26135,N_26469);
or U29485 (N_29485,N_27601,N_26991);
nand U29486 (N_29486,N_26878,N_26026);
or U29487 (N_29487,N_26319,N_26621);
xnor U29488 (N_29488,N_26632,N_26297);
nor U29489 (N_29489,N_26875,N_27929);
xor U29490 (N_29490,N_27809,N_27308);
nand U29491 (N_29491,N_26818,N_26082);
nand U29492 (N_29492,N_26114,N_27496);
nand U29493 (N_29493,N_27674,N_27690);
and U29494 (N_29494,N_26281,N_27091);
xnor U29495 (N_29495,N_27540,N_27244);
nor U29496 (N_29496,N_26500,N_26471);
nor U29497 (N_29497,N_27112,N_27657);
and U29498 (N_29498,N_27818,N_26977);
or U29499 (N_29499,N_26925,N_26161);
xor U29500 (N_29500,N_26592,N_27486);
and U29501 (N_29501,N_27244,N_26098);
nand U29502 (N_29502,N_26314,N_27212);
nor U29503 (N_29503,N_27172,N_26616);
xnor U29504 (N_29504,N_27273,N_26601);
nor U29505 (N_29505,N_26307,N_27282);
nand U29506 (N_29506,N_26583,N_27308);
nor U29507 (N_29507,N_26428,N_27541);
or U29508 (N_29508,N_27999,N_26432);
nand U29509 (N_29509,N_27261,N_26057);
or U29510 (N_29510,N_27245,N_27190);
and U29511 (N_29511,N_26713,N_27861);
or U29512 (N_29512,N_26849,N_26883);
and U29513 (N_29513,N_27982,N_27333);
and U29514 (N_29514,N_27789,N_27944);
nor U29515 (N_29515,N_26986,N_26968);
xor U29516 (N_29516,N_27433,N_27509);
xor U29517 (N_29517,N_26122,N_27527);
or U29518 (N_29518,N_27183,N_27492);
nor U29519 (N_29519,N_27560,N_26097);
or U29520 (N_29520,N_27969,N_26223);
nor U29521 (N_29521,N_27624,N_27618);
or U29522 (N_29522,N_26547,N_27465);
nand U29523 (N_29523,N_27724,N_26393);
or U29524 (N_29524,N_26675,N_27391);
xor U29525 (N_29525,N_27624,N_27589);
xor U29526 (N_29526,N_27970,N_27357);
xnor U29527 (N_29527,N_26073,N_27262);
nor U29528 (N_29528,N_27894,N_26003);
and U29529 (N_29529,N_27982,N_27950);
or U29530 (N_29530,N_27009,N_26139);
nand U29531 (N_29531,N_26881,N_27862);
nor U29532 (N_29532,N_26109,N_26122);
nor U29533 (N_29533,N_27600,N_27612);
xor U29534 (N_29534,N_26009,N_27199);
nand U29535 (N_29535,N_27972,N_26906);
and U29536 (N_29536,N_27126,N_26867);
and U29537 (N_29537,N_27269,N_27985);
or U29538 (N_29538,N_26648,N_27751);
nor U29539 (N_29539,N_26809,N_27446);
and U29540 (N_29540,N_27009,N_27302);
or U29541 (N_29541,N_26935,N_26467);
nor U29542 (N_29542,N_26847,N_27441);
nor U29543 (N_29543,N_26765,N_27182);
or U29544 (N_29544,N_27308,N_26093);
nand U29545 (N_29545,N_27675,N_27248);
xor U29546 (N_29546,N_27452,N_27377);
nand U29547 (N_29547,N_27146,N_26079);
nand U29548 (N_29548,N_27009,N_26521);
xnor U29549 (N_29549,N_26675,N_26144);
and U29550 (N_29550,N_26178,N_26976);
nand U29551 (N_29551,N_27450,N_27762);
or U29552 (N_29552,N_26917,N_26531);
and U29553 (N_29553,N_27061,N_27145);
and U29554 (N_29554,N_26384,N_26448);
nor U29555 (N_29555,N_27518,N_27370);
xnor U29556 (N_29556,N_26248,N_26190);
nand U29557 (N_29557,N_27269,N_26070);
xor U29558 (N_29558,N_26869,N_26122);
or U29559 (N_29559,N_27231,N_27316);
and U29560 (N_29560,N_26603,N_27902);
nor U29561 (N_29561,N_27170,N_26912);
or U29562 (N_29562,N_26124,N_26592);
or U29563 (N_29563,N_26120,N_26530);
nand U29564 (N_29564,N_27776,N_26045);
or U29565 (N_29565,N_26394,N_27333);
and U29566 (N_29566,N_27176,N_27279);
nor U29567 (N_29567,N_26277,N_27999);
nor U29568 (N_29568,N_27349,N_26503);
xnor U29569 (N_29569,N_26324,N_26829);
or U29570 (N_29570,N_27540,N_27384);
nand U29571 (N_29571,N_26227,N_26341);
nor U29572 (N_29572,N_27745,N_27767);
nor U29573 (N_29573,N_26356,N_27234);
nand U29574 (N_29574,N_26764,N_27841);
nor U29575 (N_29575,N_26813,N_26664);
nand U29576 (N_29576,N_27740,N_27768);
nand U29577 (N_29577,N_26769,N_27559);
nand U29578 (N_29578,N_27879,N_27233);
nand U29579 (N_29579,N_27689,N_27025);
nor U29580 (N_29580,N_26912,N_26304);
nand U29581 (N_29581,N_27744,N_27091);
and U29582 (N_29582,N_26853,N_26531);
nand U29583 (N_29583,N_27131,N_27587);
xnor U29584 (N_29584,N_26078,N_26864);
or U29585 (N_29585,N_26841,N_27710);
or U29586 (N_29586,N_26488,N_26373);
nand U29587 (N_29587,N_27228,N_26117);
and U29588 (N_29588,N_26066,N_27923);
or U29589 (N_29589,N_26517,N_27535);
or U29590 (N_29590,N_26101,N_27311);
nor U29591 (N_29591,N_26508,N_27399);
and U29592 (N_29592,N_27898,N_27089);
nand U29593 (N_29593,N_27312,N_26104);
nand U29594 (N_29594,N_27877,N_26539);
nor U29595 (N_29595,N_27029,N_26765);
xnor U29596 (N_29596,N_27187,N_27846);
xor U29597 (N_29597,N_27204,N_27983);
nor U29598 (N_29598,N_26752,N_26009);
nor U29599 (N_29599,N_27931,N_26431);
xor U29600 (N_29600,N_26497,N_26292);
nor U29601 (N_29601,N_26330,N_26924);
nor U29602 (N_29602,N_26878,N_27504);
xnor U29603 (N_29603,N_26637,N_26483);
xor U29604 (N_29604,N_26124,N_27496);
nand U29605 (N_29605,N_27652,N_26890);
nand U29606 (N_29606,N_26479,N_26638);
nor U29607 (N_29607,N_26895,N_27377);
xor U29608 (N_29608,N_26426,N_26677);
or U29609 (N_29609,N_27229,N_26102);
and U29610 (N_29610,N_26394,N_27168);
nor U29611 (N_29611,N_27488,N_27702);
xor U29612 (N_29612,N_26112,N_27588);
or U29613 (N_29613,N_27926,N_26070);
and U29614 (N_29614,N_26007,N_27147);
or U29615 (N_29615,N_27161,N_26476);
xor U29616 (N_29616,N_27731,N_27650);
or U29617 (N_29617,N_27193,N_27918);
xnor U29618 (N_29618,N_26077,N_27636);
nor U29619 (N_29619,N_27060,N_26402);
nor U29620 (N_29620,N_26067,N_26798);
and U29621 (N_29621,N_26661,N_26419);
nor U29622 (N_29622,N_26659,N_27389);
xor U29623 (N_29623,N_27285,N_27468);
or U29624 (N_29624,N_27978,N_27700);
nand U29625 (N_29625,N_26668,N_27877);
and U29626 (N_29626,N_26913,N_27819);
xor U29627 (N_29627,N_27469,N_26571);
nor U29628 (N_29628,N_27519,N_26131);
xor U29629 (N_29629,N_26268,N_26081);
nand U29630 (N_29630,N_26372,N_27188);
xnor U29631 (N_29631,N_27980,N_27514);
and U29632 (N_29632,N_27900,N_27238);
nor U29633 (N_29633,N_27352,N_26122);
and U29634 (N_29634,N_27115,N_27334);
xor U29635 (N_29635,N_27990,N_26595);
or U29636 (N_29636,N_27537,N_26387);
nand U29637 (N_29637,N_27773,N_26024);
or U29638 (N_29638,N_26461,N_27132);
and U29639 (N_29639,N_27222,N_26006);
nor U29640 (N_29640,N_27197,N_26385);
xor U29641 (N_29641,N_27927,N_27597);
nand U29642 (N_29642,N_26132,N_27032);
xor U29643 (N_29643,N_27611,N_27877);
and U29644 (N_29644,N_26739,N_27174);
nor U29645 (N_29645,N_27498,N_27372);
or U29646 (N_29646,N_26883,N_27308);
and U29647 (N_29647,N_27242,N_26550);
or U29648 (N_29648,N_27630,N_27327);
and U29649 (N_29649,N_27697,N_27035);
or U29650 (N_29650,N_26288,N_27696);
nor U29651 (N_29651,N_26152,N_26743);
nor U29652 (N_29652,N_27689,N_26817);
and U29653 (N_29653,N_27533,N_26060);
nand U29654 (N_29654,N_26670,N_26364);
or U29655 (N_29655,N_27745,N_26437);
nand U29656 (N_29656,N_27127,N_27601);
or U29657 (N_29657,N_26970,N_27590);
xor U29658 (N_29658,N_26990,N_26107);
and U29659 (N_29659,N_26396,N_26564);
nand U29660 (N_29660,N_27578,N_27553);
and U29661 (N_29661,N_26579,N_27692);
nor U29662 (N_29662,N_26240,N_27075);
xnor U29663 (N_29663,N_27058,N_26165);
xnor U29664 (N_29664,N_27020,N_27555);
xor U29665 (N_29665,N_26023,N_27199);
xor U29666 (N_29666,N_27669,N_26568);
nor U29667 (N_29667,N_26460,N_26787);
and U29668 (N_29668,N_27360,N_27897);
or U29669 (N_29669,N_26741,N_27305);
or U29670 (N_29670,N_26234,N_27539);
nor U29671 (N_29671,N_27219,N_27167);
and U29672 (N_29672,N_27652,N_27954);
nand U29673 (N_29673,N_26163,N_27478);
and U29674 (N_29674,N_26757,N_27455);
nor U29675 (N_29675,N_27324,N_26183);
xor U29676 (N_29676,N_26980,N_27331);
and U29677 (N_29677,N_26028,N_27098);
or U29678 (N_29678,N_27815,N_27339);
nor U29679 (N_29679,N_27674,N_26345);
xnor U29680 (N_29680,N_26270,N_27817);
xor U29681 (N_29681,N_27714,N_26588);
xor U29682 (N_29682,N_26474,N_26263);
nand U29683 (N_29683,N_27152,N_27226);
nor U29684 (N_29684,N_26041,N_27450);
xor U29685 (N_29685,N_27631,N_26563);
or U29686 (N_29686,N_27506,N_26530);
or U29687 (N_29687,N_27792,N_27381);
nor U29688 (N_29688,N_27725,N_26248);
xnor U29689 (N_29689,N_27653,N_27110);
nand U29690 (N_29690,N_26866,N_27425);
or U29691 (N_29691,N_26167,N_27581);
xnor U29692 (N_29692,N_27092,N_27334);
and U29693 (N_29693,N_26435,N_26250);
and U29694 (N_29694,N_27364,N_26421);
nand U29695 (N_29695,N_26388,N_26489);
and U29696 (N_29696,N_26856,N_27784);
or U29697 (N_29697,N_26169,N_26711);
or U29698 (N_29698,N_26599,N_27516);
xor U29699 (N_29699,N_27710,N_26088);
xnor U29700 (N_29700,N_26825,N_27860);
and U29701 (N_29701,N_26948,N_27785);
nor U29702 (N_29702,N_26599,N_27346);
nand U29703 (N_29703,N_26356,N_26375);
and U29704 (N_29704,N_27039,N_26562);
and U29705 (N_29705,N_27880,N_26522);
nand U29706 (N_29706,N_27739,N_26644);
nor U29707 (N_29707,N_26441,N_27607);
nor U29708 (N_29708,N_26029,N_27433);
nand U29709 (N_29709,N_27338,N_26595);
nand U29710 (N_29710,N_27838,N_26841);
xnor U29711 (N_29711,N_26233,N_27522);
nand U29712 (N_29712,N_26956,N_27740);
or U29713 (N_29713,N_27530,N_26562);
or U29714 (N_29714,N_26306,N_27504);
xnor U29715 (N_29715,N_26787,N_26648);
nand U29716 (N_29716,N_27817,N_26974);
nor U29717 (N_29717,N_26137,N_27976);
and U29718 (N_29718,N_27463,N_27128);
and U29719 (N_29719,N_26764,N_27291);
xor U29720 (N_29720,N_26913,N_26872);
or U29721 (N_29721,N_26030,N_26431);
xor U29722 (N_29722,N_26269,N_26720);
or U29723 (N_29723,N_27745,N_26030);
or U29724 (N_29724,N_26206,N_26570);
or U29725 (N_29725,N_27801,N_26228);
or U29726 (N_29726,N_26629,N_26193);
or U29727 (N_29727,N_27733,N_27213);
nand U29728 (N_29728,N_27467,N_27879);
or U29729 (N_29729,N_26961,N_26861);
or U29730 (N_29730,N_26311,N_27606);
nand U29731 (N_29731,N_27532,N_27421);
xnor U29732 (N_29732,N_26281,N_26850);
nor U29733 (N_29733,N_26112,N_26415);
nor U29734 (N_29734,N_27590,N_26691);
or U29735 (N_29735,N_26288,N_27493);
or U29736 (N_29736,N_27434,N_27200);
or U29737 (N_29737,N_26641,N_26530);
nand U29738 (N_29738,N_27975,N_27180);
nor U29739 (N_29739,N_26853,N_27603);
nor U29740 (N_29740,N_26237,N_26820);
nor U29741 (N_29741,N_26563,N_26479);
nand U29742 (N_29742,N_26883,N_26662);
nor U29743 (N_29743,N_27598,N_26455);
nand U29744 (N_29744,N_26306,N_27031);
or U29745 (N_29745,N_27591,N_26647);
xnor U29746 (N_29746,N_26990,N_27020);
nor U29747 (N_29747,N_26373,N_26009);
xnor U29748 (N_29748,N_27392,N_26661);
xor U29749 (N_29749,N_26553,N_26761);
or U29750 (N_29750,N_27926,N_27540);
nor U29751 (N_29751,N_27776,N_27771);
or U29752 (N_29752,N_27713,N_26309);
nand U29753 (N_29753,N_27564,N_26432);
and U29754 (N_29754,N_26773,N_27673);
xnor U29755 (N_29755,N_26230,N_26940);
nor U29756 (N_29756,N_27669,N_27110);
and U29757 (N_29757,N_26807,N_26193);
and U29758 (N_29758,N_27724,N_26745);
nand U29759 (N_29759,N_27722,N_26686);
xor U29760 (N_29760,N_26648,N_27967);
and U29761 (N_29761,N_27460,N_27970);
xnor U29762 (N_29762,N_27020,N_26666);
nand U29763 (N_29763,N_26039,N_27729);
or U29764 (N_29764,N_26398,N_26252);
nand U29765 (N_29765,N_26563,N_26654);
xor U29766 (N_29766,N_26329,N_27709);
xor U29767 (N_29767,N_26720,N_27478);
xnor U29768 (N_29768,N_27035,N_27125);
or U29769 (N_29769,N_26948,N_27175);
or U29770 (N_29770,N_26803,N_27509);
nand U29771 (N_29771,N_26887,N_27671);
nand U29772 (N_29772,N_26762,N_27502);
and U29773 (N_29773,N_26701,N_26628);
nand U29774 (N_29774,N_26864,N_27789);
or U29775 (N_29775,N_27517,N_27429);
nor U29776 (N_29776,N_27085,N_27248);
and U29777 (N_29777,N_26315,N_26719);
nor U29778 (N_29778,N_26452,N_27408);
nand U29779 (N_29779,N_26416,N_26664);
nand U29780 (N_29780,N_26018,N_27019);
xor U29781 (N_29781,N_27067,N_27951);
xnor U29782 (N_29782,N_26054,N_27434);
and U29783 (N_29783,N_27928,N_26764);
nor U29784 (N_29784,N_27000,N_26598);
nand U29785 (N_29785,N_27295,N_27997);
nand U29786 (N_29786,N_26968,N_26682);
nor U29787 (N_29787,N_26880,N_26680);
and U29788 (N_29788,N_26795,N_27157);
or U29789 (N_29789,N_26782,N_26555);
nand U29790 (N_29790,N_26256,N_27223);
nand U29791 (N_29791,N_27832,N_27497);
or U29792 (N_29792,N_26428,N_27474);
nand U29793 (N_29793,N_26511,N_26712);
nor U29794 (N_29794,N_26885,N_26156);
or U29795 (N_29795,N_26090,N_26629);
and U29796 (N_29796,N_27152,N_26231);
and U29797 (N_29797,N_27568,N_26726);
or U29798 (N_29798,N_26532,N_26599);
and U29799 (N_29799,N_27997,N_26632);
xnor U29800 (N_29800,N_27559,N_26581);
nor U29801 (N_29801,N_26773,N_26798);
xor U29802 (N_29802,N_26429,N_26767);
xor U29803 (N_29803,N_26342,N_26868);
or U29804 (N_29804,N_27339,N_27865);
nor U29805 (N_29805,N_27740,N_26021);
or U29806 (N_29806,N_26900,N_26710);
nor U29807 (N_29807,N_26551,N_27256);
or U29808 (N_29808,N_26382,N_27173);
xor U29809 (N_29809,N_26172,N_27633);
xor U29810 (N_29810,N_27807,N_26587);
and U29811 (N_29811,N_27351,N_27520);
xnor U29812 (N_29812,N_27095,N_26050);
and U29813 (N_29813,N_27762,N_27521);
nor U29814 (N_29814,N_26267,N_27486);
or U29815 (N_29815,N_26580,N_27308);
nor U29816 (N_29816,N_27134,N_26196);
nor U29817 (N_29817,N_26053,N_27694);
and U29818 (N_29818,N_26849,N_26856);
xor U29819 (N_29819,N_27653,N_26656);
or U29820 (N_29820,N_27632,N_27156);
xor U29821 (N_29821,N_26347,N_27792);
or U29822 (N_29822,N_26940,N_27066);
nor U29823 (N_29823,N_27507,N_26361);
or U29824 (N_29824,N_27608,N_26031);
nor U29825 (N_29825,N_26116,N_27282);
and U29826 (N_29826,N_26249,N_27353);
or U29827 (N_29827,N_27326,N_27251);
nand U29828 (N_29828,N_27888,N_26417);
or U29829 (N_29829,N_27457,N_26196);
or U29830 (N_29830,N_26017,N_27699);
nor U29831 (N_29831,N_26314,N_27329);
xnor U29832 (N_29832,N_27364,N_27161);
nand U29833 (N_29833,N_26515,N_26833);
or U29834 (N_29834,N_26511,N_27745);
and U29835 (N_29835,N_27359,N_27884);
or U29836 (N_29836,N_27223,N_26702);
or U29837 (N_29837,N_27003,N_27397);
and U29838 (N_29838,N_26394,N_27535);
nand U29839 (N_29839,N_27233,N_26429);
and U29840 (N_29840,N_27900,N_27928);
nor U29841 (N_29841,N_26929,N_27289);
and U29842 (N_29842,N_26884,N_27424);
nor U29843 (N_29843,N_26331,N_26045);
xor U29844 (N_29844,N_26975,N_27990);
nor U29845 (N_29845,N_26302,N_27248);
nand U29846 (N_29846,N_26555,N_26203);
or U29847 (N_29847,N_26110,N_27385);
nand U29848 (N_29848,N_27769,N_27633);
nand U29849 (N_29849,N_27078,N_27314);
nand U29850 (N_29850,N_26108,N_27518);
nand U29851 (N_29851,N_27217,N_26763);
nor U29852 (N_29852,N_27999,N_26801);
nand U29853 (N_29853,N_26278,N_27081);
nand U29854 (N_29854,N_26511,N_27136);
nand U29855 (N_29855,N_27017,N_27394);
and U29856 (N_29856,N_26307,N_26106);
xnor U29857 (N_29857,N_27622,N_27791);
nor U29858 (N_29858,N_27286,N_27068);
or U29859 (N_29859,N_27658,N_26938);
or U29860 (N_29860,N_26483,N_26052);
nor U29861 (N_29861,N_26547,N_26233);
and U29862 (N_29862,N_26830,N_27212);
xor U29863 (N_29863,N_26230,N_26687);
or U29864 (N_29864,N_27244,N_27374);
nand U29865 (N_29865,N_27500,N_26154);
nor U29866 (N_29866,N_26177,N_27327);
or U29867 (N_29867,N_26162,N_26962);
nand U29868 (N_29868,N_27306,N_26007);
nand U29869 (N_29869,N_26865,N_27320);
nor U29870 (N_29870,N_27697,N_27146);
or U29871 (N_29871,N_27876,N_27002);
and U29872 (N_29872,N_26918,N_26616);
and U29873 (N_29873,N_27672,N_26624);
or U29874 (N_29874,N_27320,N_27736);
and U29875 (N_29875,N_26034,N_26027);
and U29876 (N_29876,N_27505,N_27391);
and U29877 (N_29877,N_26087,N_27127);
and U29878 (N_29878,N_27328,N_26828);
xor U29879 (N_29879,N_26564,N_27109);
nand U29880 (N_29880,N_27402,N_27228);
xor U29881 (N_29881,N_27438,N_26219);
nand U29882 (N_29882,N_26688,N_26146);
or U29883 (N_29883,N_26107,N_26862);
or U29884 (N_29884,N_27151,N_27288);
nand U29885 (N_29885,N_26072,N_27540);
nor U29886 (N_29886,N_26189,N_26632);
nand U29887 (N_29887,N_27142,N_26108);
nor U29888 (N_29888,N_26000,N_26510);
or U29889 (N_29889,N_26525,N_27817);
nor U29890 (N_29890,N_27508,N_27333);
xor U29891 (N_29891,N_27178,N_27421);
nand U29892 (N_29892,N_26018,N_26040);
nor U29893 (N_29893,N_27315,N_27156);
nand U29894 (N_29894,N_26915,N_27880);
nor U29895 (N_29895,N_27351,N_26895);
nand U29896 (N_29896,N_27729,N_27845);
or U29897 (N_29897,N_27213,N_26193);
or U29898 (N_29898,N_26750,N_26465);
nand U29899 (N_29899,N_26275,N_27554);
nand U29900 (N_29900,N_27330,N_27991);
nor U29901 (N_29901,N_27030,N_26720);
nand U29902 (N_29902,N_27934,N_26883);
or U29903 (N_29903,N_27646,N_26454);
and U29904 (N_29904,N_27045,N_27985);
nor U29905 (N_29905,N_27842,N_27602);
nor U29906 (N_29906,N_27163,N_26015);
and U29907 (N_29907,N_27031,N_26361);
nor U29908 (N_29908,N_26151,N_26028);
and U29909 (N_29909,N_27893,N_27497);
nor U29910 (N_29910,N_26800,N_27438);
and U29911 (N_29911,N_26918,N_26271);
nand U29912 (N_29912,N_27135,N_26863);
or U29913 (N_29913,N_27834,N_27375);
nand U29914 (N_29914,N_27733,N_27172);
nor U29915 (N_29915,N_26529,N_26562);
and U29916 (N_29916,N_26122,N_27241);
nor U29917 (N_29917,N_27865,N_27474);
and U29918 (N_29918,N_27893,N_27258);
nor U29919 (N_29919,N_27610,N_27843);
xnor U29920 (N_29920,N_27464,N_27129);
nand U29921 (N_29921,N_26671,N_27515);
nor U29922 (N_29922,N_27271,N_26622);
or U29923 (N_29923,N_27958,N_27531);
nand U29924 (N_29924,N_27710,N_27527);
and U29925 (N_29925,N_26927,N_26404);
nand U29926 (N_29926,N_26890,N_26401);
nand U29927 (N_29927,N_26707,N_26909);
and U29928 (N_29928,N_26031,N_26559);
or U29929 (N_29929,N_27032,N_26040);
and U29930 (N_29930,N_26101,N_26067);
nand U29931 (N_29931,N_26792,N_27110);
or U29932 (N_29932,N_27381,N_27447);
and U29933 (N_29933,N_27190,N_27341);
or U29934 (N_29934,N_27666,N_27357);
or U29935 (N_29935,N_27079,N_27931);
or U29936 (N_29936,N_26867,N_27731);
xnor U29937 (N_29937,N_26071,N_26114);
nand U29938 (N_29938,N_27607,N_26326);
and U29939 (N_29939,N_27085,N_26144);
nand U29940 (N_29940,N_27804,N_27344);
or U29941 (N_29941,N_26124,N_27355);
nand U29942 (N_29942,N_26602,N_26459);
or U29943 (N_29943,N_26819,N_26036);
or U29944 (N_29944,N_26293,N_26272);
nand U29945 (N_29945,N_26016,N_27978);
xnor U29946 (N_29946,N_27372,N_27370);
xor U29947 (N_29947,N_27214,N_26629);
nor U29948 (N_29948,N_27905,N_27580);
nand U29949 (N_29949,N_27094,N_26734);
and U29950 (N_29950,N_27123,N_27810);
and U29951 (N_29951,N_26554,N_26593);
nand U29952 (N_29952,N_27579,N_27571);
xnor U29953 (N_29953,N_26305,N_27370);
or U29954 (N_29954,N_27316,N_27530);
or U29955 (N_29955,N_27321,N_26488);
nor U29956 (N_29956,N_26566,N_27839);
nand U29957 (N_29957,N_26070,N_26816);
nor U29958 (N_29958,N_27271,N_26665);
and U29959 (N_29959,N_26830,N_27809);
nand U29960 (N_29960,N_27417,N_26961);
nor U29961 (N_29961,N_26457,N_26804);
nand U29962 (N_29962,N_26376,N_27498);
xor U29963 (N_29963,N_26315,N_26557);
nand U29964 (N_29964,N_26403,N_26973);
nor U29965 (N_29965,N_26061,N_26974);
nor U29966 (N_29966,N_26651,N_26089);
xor U29967 (N_29967,N_26338,N_27887);
and U29968 (N_29968,N_26190,N_27054);
xnor U29969 (N_29969,N_27667,N_27524);
or U29970 (N_29970,N_27308,N_26821);
and U29971 (N_29971,N_26083,N_27451);
nand U29972 (N_29972,N_27021,N_26693);
xor U29973 (N_29973,N_26351,N_26628);
xor U29974 (N_29974,N_27859,N_27330);
or U29975 (N_29975,N_27961,N_27113);
nand U29976 (N_29976,N_26896,N_26671);
nand U29977 (N_29977,N_27670,N_27514);
nand U29978 (N_29978,N_26690,N_27058);
or U29979 (N_29979,N_26670,N_27134);
xnor U29980 (N_29980,N_26327,N_27864);
and U29981 (N_29981,N_27233,N_27824);
or U29982 (N_29982,N_27054,N_26921);
or U29983 (N_29983,N_27873,N_26201);
or U29984 (N_29984,N_26750,N_26605);
or U29985 (N_29985,N_27999,N_27854);
nor U29986 (N_29986,N_26994,N_26349);
xnor U29987 (N_29987,N_26365,N_26169);
or U29988 (N_29988,N_27782,N_26133);
nor U29989 (N_29989,N_27106,N_26288);
and U29990 (N_29990,N_27978,N_26921);
nand U29991 (N_29991,N_27006,N_26862);
and U29992 (N_29992,N_27312,N_26300);
xor U29993 (N_29993,N_26855,N_27579);
xor U29994 (N_29994,N_27675,N_27366);
nand U29995 (N_29995,N_26263,N_26993);
nand U29996 (N_29996,N_26731,N_26542);
nor U29997 (N_29997,N_27594,N_26304);
nand U29998 (N_29998,N_26112,N_26866);
xor U29999 (N_29999,N_26878,N_27385);
nor UO_0 (O_0,N_29868,N_28474);
or UO_1 (O_1,N_28892,N_28303);
nor UO_2 (O_2,N_28513,N_28129);
nor UO_3 (O_3,N_29306,N_29672);
nor UO_4 (O_4,N_29141,N_28629);
and UO_5 (O_5,N_28985,N_29162);
nand UO_6 (O_6,N_28295,N_28644);
or UO_7 (O_7,N_29484,N_29611);
and UO_8 (O_8,N_29147,N_28789);
nor UO_9 (O_9,N_29858,N_28328);
xor UO_10 (O_10,N_28000,N_29145);
and UO_11 (O_11,N_28854,N_29377);
xnor UO_12 (O_12,N_28778,N_29144);
and UO_13 (O_13,N_29985,N_29091);
and UO_14 (O_14,N_28201,N_28735);
nor UO_15 (O_15,N_28554,N_28332);
and UO_16 (O_16,N_28533,N_29287);
or UO_17 (O_17,N_28902,N_28917);
or UO_18 (O_18,N_28458,N_29729);
and UO_19 (O_19,N_29875,N_28802);
nor UO_20 (O_20,N_29195,N_29876);
or UO_21 (O_21,N_28991,N_28769);
or UO_22 (O_22,N_29515,N_28733);
and UO_23 (O_23,N_28023,N_28349);
xnor UO_24 (O_24,N_29624,N_28298);
nand UO_25 (O_25,N_29790,N_28687);
or UO_26 (O_26,N_28326,N_29295);
and UO_27 (O_27,N_29165,N_28026);
nand UO_28 (O_28,N_29955,N_29978);
xnor UO_29 (O_29,N_28098,N_28357);
or UO_30 (O_30,N_28764,N_29601);
and UO_31 (O_31,N_29084,N_28128);
xor UO_32 (O_32,N_29528,N_28369);
or UO_33 (O_33,N_29372,N_28439);
nand UO_34 (O_34,N_28220,N_28099);
xor UO_35 (O_35,N_28924,N_29704);
nor UO_36 (O_36,N_28397,N_29213);
and UO_37 (O_37,N_29090,N_28017);
xnor UO_38 (O_38,N_28324,N_28910);
nor UO_39 (O_39,N_28176,N_29284);
and UO_40 (O_40,N_28333,N_29166);
or UO_41 (O_41,N_28530,N_29417);
xnor UO_42 (O_42,N_29553,N_29524);
and UO_43 (O_43,N_28879,N_29029);
nor UO_44 (O_44,N_29664,N_29730);
nand UO_45 (O_45,N_29842,N_28024);
or UO_46 (O_46,N_28509,N_28813);
and UO_47 (O_47,N_29971,N_29440);
nand UO_48 (O_48,N_28732,N_28634);
nor UO_49 (O_49,N_28962,N_29873);
nor UO_50 (O_50,N_28981,N_28928);
and UO_51 (O_51,N_28388,N_28245);
nand UO_52 (O_52,N_29131,N_28231);
xnor UO_53 (O_53,N_28641,N_28174);
xnor UO_54 (O_54,N_28102,N_29623);
nand UO_55 (O_55,N_29050,N_29206);
xnor UO_56 (O_56,N_28539,N_29738);
nor UO_57 (O_57,N_28811,N_29191);
or UO_58 (O_58,N_28689,N_29374);
and UO_59 (O_59,N_29902,N_29411);
nor UO_60 (O_60,N_29519,N_28932);
and UO_61 (O_61,N_29156,N_28125);
nor UO_62 (O_62,N_29444,N_29547);
or UO_63 (O_63,N_28771,N_28524);
or UO_64 (O_64,N_28786,N_29916);
nand UO_65 (O_65,N_28422,N_28006);
xor UO_66 (O_66,N_28100,N_28543);
or UO_67 (O_67,N_28287,N_29840);
nor UO_68 (O_68,N_28294,N_29402);
or UO_69 (O_69,N_28885,N_29341);
xnor UO_70 (O_70,N_28268,N_29757);
xnor UO_71 (O_71,N_29817,N_28829);
or UO_72 (O_72,N_28720,N_28659);
xnor UO_73 (O_73,N_28149,N_29111);
or UO_74 (O_74,N_28471,N_29115);
xor UO_75 (O_75,N_29708,N_28886);
xnor UO_76 (O_76,N_29752,N_29210);
or UO_77 (O_77,N_28156,N_28107);
nor UO_78 (O_78,N_29001,N_28219);
and UO_79 (O_79,N_29671,N_29311);
nor UO_80 (O_80,N_28404,N_28865);
or UO_81 (O_81,N_29563,N_29371);
nand UO_82 (O_82,N_29514,N_29074);
nor UO_83 (O_83,N_28187,N_29520);
nand UO_84 (O_84,N_28817,N_29655);
nand UO_85 (O_85,N_29953,N_29567);
and UO_86 (O_86,N_28657,N_29215);
nor UO_87 (O_87,N_29745,N_28348);
nor UO_88 (O_88,N_28613,N_29496);
or UO_89 (O_89,N_29022,N_29260);
nor UO_90 (O_90,N_28822,N_28588);
xor UO_91 (O_91,N_28140,N_29312);
nand UO_92 (O_92,N_29245,N_29118);
or UO_93 (O_93,N_28647,N_29964);
nor UO_94 (O_94,N_28618,N_28267);
and UO_95 (O_95,N_28546,N_28265);
nand UO_96 (O_96,N_28807,N_29353);
nand UO_97 (O_97,N_28331,N_29650);
nand UO_98 (O_98,N_28581,N_28446);
nand UO_99 (O_99,N_29635,N_29716);
or UO_100 (O_100,N_29951,N_28449);
nor UO_101 (O_101,N_29913,N_29238);
or UO_102 (O_102,N_29645,N_28645);
nand UO_103 (O_103,N_28352,N_28234);
nor UO_104 (O_104,N_28034,N_29930);
xnor UO_105 (O_105,N_29552,N_29854);
nor UO_106 (O_106,N_29651,N_28749);
and UO_107 (O_107,N_28361,N_28240);
nand UO_108 (O_108,N_28428,N_28461);
xnor UO_109 (O_109,N_28013,N_28435);
nor UO_110 (O_110,N_28716,N_28721);
or UO_111 (O_111,N_28041,N_29430);
xor UO_112 (O_112,N_29850,N_29468);
xnor UO_113 (O_113,N_29797,N_28269);
nor UO_114 (O_114,N_28358,N_28289);
xnor UO_115 (O_115,N_29862,N_28061);
or UO_116 (O_116,N_28230,N_29682);
nor UO_117 (O_117,N_29820,N_29420);
or UO_118 (O_118,N_28650,N_29719);
xnor UO_119 (O_119,N_28929,N_28171);
nand UO_120 (O_120,N_28906,N_28150);
nand UO_121 (O_121,N_29944,N_28598);
and UO_122 (O_122,N_29934,N_28405);
nor UO_123 (O_123,N_29229,N_28677);
xnor UO_124 (O_124,N_29660,N_29346);
xor UO_125 (O_125,N_29825,N_28915);
and UO_126 (O_126,N_28092,N_29431);
xor UO_127 (O_127,N_29523,N_28907);
and UO_128 (O_128,N_28393,N_29779);
nor UO_129 (O_129,N_29300,N_28266);
nand UO_130 (O_130,N_29591,N_28763);
nor UO_131 (O_131,N_29365,N_28978);
nand UO_132 (O_132,N_29816,N_28052);
and UO_133 (O_133,N_29448,N_29460);
xnor UO_134 (O_134,N_29441,N_29390);
xor UO_135 (O_135,N_28712,N_29721);
xor UO_136 (O_136,N_28561,N_29235);
xor UO_137 (O_137,N_28237,N_28473);
nand UO_138 (O_138,N_29775,N_28105);
and UO_139 (O_139,N_28726,N_28481);
nor UO_140 (O_140,N_28842,N_28195);
or UO_141 (O_141,N_29322,N_29389);
nand UO_142 (O_142,N_29539,N_28384);
or UO_143 (O_143,N_28632,N_28517);
nand UO_144 (O_144,N_28489,N_29271);
nand UO_145 (O_145,N_29694,N_29011);
and UO_146 (O_146,N_29218,N_29697);
nor UO_147 (O_147,N_28126,N_28706);
xnor UO_148 (O_148,N_29072,N_29356);
or UO_149 (O_149,N_29408,N_28457);
or UO_150 (O_150,N_29297,N_28680);
xnor UO_151 (O_151,N_28299,N_28567);
nor UO_152 (O_152,N_29424,N_29965);
nand UO_153 (O_153,N_29616,N_28708);
nor UO_154 (O_154,N_29178,N_28002);
nor UO_155 (O_155,N_29387,N_29332);
xor UO_156 (O_156,N_29681,N_29193);
or UO_157 (O_157,N_29990,N_29239);
or UO_158 (O_158,N_29846,N_29288);
and UO_159 (O_159,N_28636,N_29693);
and UO_160 (O_160,N_28127,N_28313);
xor UO_161 (O_161,N_28531,N_28623);
nor UO_162 (O_162,N_28470,N_28551);
nor UO_163 (O_163,N_28182,N_28057);
xnor UO_164 (O_164,N_29807,N_29626);
and UO_165 (O_165,N_29548,N_29622);
and UO_166 (O_166,N_28091,N_29740);
nand UO_167 (O_167,N_28516,N_29199);
nand UO_168 (O_168,N_29502,N_29543);
nor UO_169 (O_169,N_28027,N_28916);
nor UO_170 (O_170,N_28258,N_29061);
and UO_171 (O_171,N_28438,N_29168);
xor UO_172 (O_172,N_29109,N_29443);
or UO_173 (O_173,N_29247,N_29362);
and UO_174 (O_174,N_29002,N_28994);
xor UO_175 (O_175,N_28407,N_28445);
xnor UO_176 (O_176,N_28600,N_28047);
nor UO_177 (O_177,N_29452,N_29824);
xor UO_178 (O_178,N_28083,N_29856);
and UO_179 (O_179,N_29851,N_28007);
nand UO_180 (O_180,N_29703,N_29637);
nor UO_181 (O_181,N_28003,N_28610);
and UO_182 (O_182,N_29941,N_29568);
and UO_183 (O_183,N_29897,N_28717);
nand UO_184 (O_184,N_28164,N_29052);
xor UO_185 (O_185,N_28897,N_29410);
and UO_186 (O_186,N_29019,N_28323);
and UO_187 (O_187,N_28893,N_29056);
xnor UO_188 (O_188,N_29059,N_28968);
and UO_189 (O_189,N_28946,N_28825);
xnor UO_190 (O_190,N_29844,N_28077);
and UO_191 (O_191,N_29989,N_29778);
nor UO_192 (O_192,N_28711,N_28232);
or UO_193 (O_193,N_28396,N_28049);
or UO_194 (O_194,N_29764,N_29878);
xor UO_195 (O_195,N_29426,N_28983);
and UO_196 (O_196,N_29170,N_28227);
nor UO_197 (O_197,N_28365,N_29025);
xnor UO_198 (O_198,N_28690,N_28974);
xor UO_199 (O_199,N_29291,N_28197);
xor UO_200 (O_200,N_28812,N_29077);
xnor UO_201 (O_201,N_29344,N_28300);
and UO_202 (O_202,N_28198,N_29422);
xor UO_203 (O_203,N_28819,N_28982);
and UO_204 (O_204,N_28661,N_28109);
xor UO_205 (O_205,N_29244,N_29483);
and UO_206 (O_206,N_29108,N_29017);
or UO_207 (O_207,N_28165,N_28288);
nand UO_208 (O_208,N_29838,N_29273);
nor UO_209 (O_209,N_28071,N_28669);
nor UO_210 (O_210,N_29892,N_29434);
nand UO_211 (O_211,N_29909,N_29834);
or UO_212 (O_212,N_28599,N_28878);
xnor UO_213 (O_213,N_28980,N_29835);
and UO_214 (O_214,N_28167,N_29119);
nand UO_215 (O_215,N_28591,N_29429);
nand UO_216 (O_216,N_29639,N_29340);
or UO_217 (O_217,N_28360,N_28311);
nor UO_218 (O_218,N_28961,N_29146);
xor UO_219 (O_219,N_28005,N_28930);
xor UO_220 (O_220,N_28483,N_29004);
or UO_221 (O_221,N_29038,N_28903);
nand UO_222 (O_222,N_29678,N_29554);
xnor UO_223 (O_223,N_29604,N_28593);
nor UO_224 (O_224,N_28501,N_28821);
or UO_225 (O_225,N_29805,N_29958);
or UO_226 (O_226,N_29026,N_28949);
and UO_227 (O_227,N_28325,N_29970);
or UO_228 (O_228,N_28199,N_29647);
xor UO_229 (O_229,N_29728,N_28922);
or UO_230 (O_230,N_28875,N_29290);
or UO_231 (O_231,N_29453,N_29125);
and UO_232 (O_232,N_29500,N_29915);
nand UO_233 (O_233,N_28018,N_28620);
or UO_234 (O_234,N_28188,N_29919);
nor UO_235 (O_235,N_28568,N_28111);
and UO_236 (O_236,N_28606,N_28364);
nor UO_237 (O_237,N_29883,N_28996);
or UO_238 (O_238,N_29319,N_28837);
nand UO_239 (O_239,N_28465,N_28609);
and UO_240 (O_240,N_29602,N_29078);
nor UO_241 (O_241,N_29559,N_29925);
and UO_242 (O_242,N_29298,N_28538);
nand UO_243 (O_243,N_28162,N_28448);
and UO_244 (O_244,N_28355,N_28894);
and UO_245 (O_245,N_29605,N_28212);
and UO_246 (O_246,N_29041,N_29134);
nor UO_247 (O_247,N_29761,N_29644);
or UO_248 (O_248,N_28029,N_28054);
nand UO_249 (O_249,N_28498,N_29252);
nor UO_250 (O_250,N_29413,N_29636);
nor UO_251 (O_251,N_29427,N_29907);
or UO_252 (O_252,N_29870,N_28208);
or UO_253 (O_253,N_29254,N_28969);
xor UO_254 (O_254,N_29133,N_28801);
xor UO_255 (O_255,N_29766,N_29330);
nand UO_256 (O_256,N_29081,N_28663);
nand UO_257 (O_257,N_29898,N_29815);
nor UO_258 (O_258,N_28056,N_28139);
nand UO_259 (O_259,N_29760,N_29580);
nor UO_260 (O_260,N_28014,N_28860);
xnor UO_261 (O_261,N_28800,N_29348);
and UO_262 (O_262,N_29927,N_28876);
and UO_263 (O_263,N_29201,N_28975);
xor UO_264 (O_264,N_29836,N_29711);
and UO_265 (O_265,N_29795,N_29618);
nor UO_266 (O_266,N_29584,N_29446);
and UO_267 (O_267,N_28437,N_28114);
nor UO_268 (O_268,N_29378,N_29498);
and UO_269 (O_269,N_29590,N_28226);
and UO_270 (O_270,N_29649,N_29606);
and UO_271 (O_271,N_28345,N_29739);
nand UO_272 (O_272,N_28228,N_29905);
nand UO_273 (O_273,N_29734,N_29037);
xor UO_274 (O_274,N_29046,N_29407);
or UO_275 (O_275,N_28637,N_28851);
or UO_276 (O_276,N_28069,N_29717);
xnor UO_277 (O_277,N_29171,N_28296);
or UO_278 (O_278,N_28466,N_28891);
nor UO_279 (O_279,N_28713,N_28389);
xor UO_280 (O_280,N_29024,N_28490);
nor UO_281 (O_281,N_29073,N_29327);
xor UO_282 (O_282,N_29819,N_28161);
nand UO_283 (O_283,N_29105,N_29759);
and UO_284 (O_284,N_29124,N_29656);
xnor UO_285 (O_285,N_28134,N_29304);
or UO_286 (O_286,N_29230,N_28584);
xnor UO_287 (O_287,N_29360,N_28253);
nor UO_288 (O_288,N_28214,N_28774);
xor UO_289 (O_289,N_28883,N_29347);
nor UO_290 (O_290,N_28122,N_29653);
nor UO_291 (O_291,N_29954,N_29801);
nand UO_292 (O_292,N_29474,N_28725);
and UO_293 (O_293,N_29541,N_28196);
nor UO_294 (O_294,N_28064,N_28904);
or UO_295 (O_295,N_29555,N_29397);
xnor UO_296 (O_296,N_28523,N_29732);
nand UO_297 (O_297,N_28642,N_29275);
or UO_298 (O_298,N_29343,N_29943);
or UO_299 (O_299,N_29363,N_28455);
xor UO_300 (O_300,N_28674,N_29532);
or UO_301 (O_301,N_28247,N_28502);
nor UO_302 (O_302,N_28412,N_28339);
nand UO_303 (O_303,N_28039,N_29487);
and UO_304 (O_304,N_29456,N_29279);
xnor UO_305 (O_305,N_28900,N_28803);
xnor UO_306 (O_306,N_29083,N_28491);
or UO_307 (O_307,N_28415,N_29464);
nor UO_308 (O_308,N_28011,N_28032);
nand UO_309 (O_309,N_28486,N_28304);
and UO_310 (O_310,N_29465,N_28124);
or UO_311 (O_311,N_29065,N_29710);
or UO_312 (O_312,N_28571,N_28381);
and UO_313 (O_313,N_28291,N_28565);
nand UO_314 (O_314,N_28849,N_28096);
nand UO_315 (O_315,N_28037,N_28989);
xor UO_316 (O_316,N_29035,N_28792);
and UO_317 (O_317,N_29910,N_29324);
xnor UO_318 (O_318,N_29629,N_29673);
nor UO_319 (O_319,N_29993,N_29966);
nand UO_320 (O_320,N_28675,N_28948);
xor UO_321 (O_321,N_29471,N_28261);
nor UO_322 (O_322,N_28464,N_28478);
and UO_323 (O_323,N_29110,N_28863);
xnor UO_324 (O_324,N_29712,N_29659);
nand UO_325 (O_325,N_29047,N_28432);
nor UO_326 (O_326,N_29299,N_29936);
and UO_327 (O_327,N_28714,N_28979);
nor UO_328 (O_328,N_28635,N_29163);
or UO_329 (O_329,N_29490,N_29478);
and UO_330 (O_330,N_28617,N_28068);
nand UO_331 (O_331,N_29981,N_29294);
and UO_332 (O_332,N_29316,N_28757);
xor UO_333 (O_333,N_29048,N_28649);
nand UO_334 (O_334,N_28814,N_28236);
nand UO_335 (O_335,N_29744,N_28806);
nand UO_336 (O_336,N_29224,N_28387);
nor UO_337 (O_337,N_29253,N_28877);
xor UO_338 (O_338,N_29725,N_28235);
or UO_339 (O_339,N_28104,N_29718);
xnor UO_340 (O_340,N_29153,N_28500);
nor UO_341 (O_341,N_29830,N_28282);
and UO_342 (O_342,N_28604,N_29724);
xor UO_343 (O_343,N_28505,N_29207);
or UO_344 (O_344,N_28153,N_28520);
and UO_345 (O_345,N_29695,N_29173);
and UO_346 (O_346,N_29013,N_28777);
xor UO_347 (O_347,N_28089,N_29665);
and UO_348 (O_348,N_29385,N_28694);
or UO_349 (O_349,N_28559,N_29136);
or UO_350 (O_350,N_28737,N_29317);
and UO_351 (O_351,N_29544,N_28085);
or UO_352 (O_352,N_28507,N_29589);
xnor UO_353 (O_353,N_28537,N_28354);
or UO_354 (O_354,N_28882,N_29242);
nand UO_355 (O_355,N_28960,N_28366);
or UO_356 (O_356,N_29039,N_29803);
nor UO_357 (O_357,N_29194,N_28662);
xnor UO_358 (O_358,N_28577,N_29351);
and UO_359 (O_359,N_29986,N_28004);
and UO_360 (O_360,N_29786,N_29578);
and UO_361 (O_361,N_28009,N_29612);
or UO_362 (O_362,N_28857,N_28351);
nand UO_363 (O_363,N_28884,N_29747);
or UO_364 (O_364,N_28084,N_29848);
and UO_365 (O_365,N_29009,N_28276);
nor UO_366 (O_366,N_28654,N_29505);
xnor UO_367 (O_367,N_29438,N_28142);
or UO_368 (O_368,N_29669,N_28673);
nor UO_369 (O_369,N_29379,N_28444);
or UO_370 (O_370,N_29450,N_29433);
nand UO_371 (O_371,N_28353,N_28705);
or UO_372 (O_372,N_29564,N_29551);
xor UO_373 (O_373,N_28416,N_28211);
nor UO_374 (O_374,N_29234,N_28036);
nand UO_375 (O_375,N_28492,N_28738);
nand UO_376 (O_376,N_29727,N_28552);
or UO_377 (O_377,N_28545,N_28377);
xor UO_378 (O_378,N_28828,N_29506);
or UO_379 (O_379,N_29219,N_29049);
and UO_380 (O_380,N_29000,N_28012);
xor UO_381 (O_381,N_28881,N_28867);
xor UO_382 (O_382,N_28751,N_29281);
nand UO_383 (O_383,N_29619,N_29722);
xnor UO_384 (O_384,N_28776,N_28651);
xor UO_385 (O_385,N_29228,N_29236);
nor UO_386 (O_386,N_28586,N_29685);
or UO_387 (O_387,N_28221,N_29699);
or UO_388 (O_388,N_29227,N_28193);
nor UO_389 (O_389,N_29391,N_29055);
and UO_390 (O_390,N_29741,N_28958);
nor UO_391 (O_391,N_29042,N_29068);
nor UO_392 (O_392,N_29791,N_29398);
nor UO_393 (O_393,N_29837,N_28146);
nand UO_394 (O_394,N_28191,N_29154);
or UO_395 (O_395,N_29096,N_28999);
nand UO_396 (O_396,N_29093,N_29977);
or UO_397 (O_397,N_28159,N_29648);
or UO_398 (O_398,N_28033,N_29597);
xor UO_399 (O_399,N_29044,N_28990);
nor UO_400 (O_400,N_28755,N_29302);
nor UO_401 (O_401,N_28409,N_28818);
or UO_402 (O_402,N_29674,N_29089);
or UO_403 (O_403,N_29489,N_29203);
nand UO_404 (O_404,N_28678,N_28823);
xnor UO_405 (O_405,N_29501,N_29871);
xor UO_406 (O_406,N_29032,N_28976);
nor UO_407 (O_407,N_28556,N_28587);
and UO_408 (O_408,N_28805,N_28627);
nand UO_409 (O_409,N_28986,N_28206);
or UO_410 (O_410,N_28336,N_29008);
nor UO_411 (O_411,N_28558,N_29799);
xnor UO_412 (O_412,N_29904,N_29890);
nand UO_413 (O_413,N_29337,N_29662);
xor UO_414 (O_414,N_28223,N_29384);
nand UO_415 (O_415,N_29097,N_28855);
nand UO_416 (O_416,N_28992,N_28392);
nand UO_417 (O_417,N_28548,N_28430);
nor UO_418 (O_418,N_28178,N_29646);
xnor UO_419 (O_419,N_28482,N_28233);
nor UO_420 (O_420,N_28053,N_28493);
xor UO_421 (O_421,N_28270,N_28209);
nor UO_422 (O_422,N_29928,N_29114);
or UO_423 (O_423,N_29040,N_28512);
nand UO_424 (O_424,N_28506,N_29517);
and UO_425 (O_425,N_28145,N_28936);
nand UO_426 (O_426,N_28756,N_28147);
or UO_427 (O_427,N_28967,N_29885);
nand UO_428 (O_428,N_29908,N_28427);
nand UO_429 (O_429,N_29172,N_29075);
xnor UO_430 (O_430,N_28569,N_29933);
nand UO_431 (O_431,N_28843,N_28399);
and UO_432 (O_432,N_29696,N_28487);
xor UO_433 (O_433,N_29027,N_29720);
and UO_434 (O_434,N_28977,N_29668);
or UO_435 (O_435,N_29099,N_29071);
nand UO_436 (O_436,N_28656,N_29030);
nand UO_437 (O_437,N_28484,N_29866);
xor UO_438 (O_438,N_28433,N_29959);
nor UO_439 (O_439,N_29789,N_28648);
or UO_440 (O_440,N_29676,N_28031);
and UO_441 (O_441,N_29395,N_28964);
or UO_442 (O_442,N_28938,N_29600);
and UO_443 (O_443,N_29473,N_28138);
or UO_444 (O_444,N_29293,N_29888);
or UO_445 (O_445,N_28108,N_28872);
or UO_446 (O_446,N_28421,N_29918);
or UO_447 (O_447,N_28462,N_28779);
or UO_448 (O_448,N_29182,N_28852);
or UO_449 (O_449,N_29007,N_29526);
nor UO_450 (O_450,N_29882,N_28601);
xnor UO_451 (O_451,N_29571,N_29968);
or UO_452 (O_452,N_28622,N_28784);
nand UO_453 (O_453,N_28927,N_29045);
nor UO_454 (O_454,N_29536,N_29416);
nor UO_455 (O_455,N_28692,N_29537);
and UO_456 (O_456,N_29823,N_28218);
nand UO_457 (O_457,N_28639,N_29157);
or UO_458 (O_458,N_28959,N_28862);
and UO_459 (O_459,N_28781,N_28783);
or UO_460 (O_460,N_28861,N_29307);
or UO_461 (O_461,N_29204,N_29021);
xor UO_462 (O_462,N_29034,N_28955);
nor UO_463 (O_463,N_28186,N_29183);
xor UO_464 (O_464,N_29631,N_28790);
nor UO_465 (O_465,N_29216,N_29036);
xor UO_466 (O_466,N_29043,N_29995);
and UO_467 (O_467,N_29872,N_29278);
xnor UO_468 (O_468,N_28170,N_29280);
xor UO_469 (O_469,N_29628,N_28244);
nor UO_470 (O_470,N_28497,N_28788);
nor UO_471 (O_471,N_29126,N_28425);
or UO_472 (O_472,N_29509,N_29533);
nor UO_473 (O_473,N_28603,N_28463);
or UO_474 (O_474,N_29463,N_28723);
nand UO_475 (O_475,N_28136,N_29177);
or UO_476 (O_476,N_29342,N_28321);
nor UO_477 (O_477,N_28204,N_28504);
nand UO_478 (O_478,N_29894,N_29282);
and UO_479 (O_479,N_29583,N_28155);
and UO_480 (O_480,N_29076,N_29485);
or UO_481 (O_481,N_28592,N_28665);
nand UO_482 (O_482,N_28271,N_28625);
nor UO_483 (O_483,N_28225,N_29736);
or UO_484 (O_484,N_29421,N_28844);
xor UO_485 (O_485,N_29367,N_29792);
and UO_486 (O_486,N_29237,N_29366);
and UO_487 (O_487,N_29094,N_29960);
and UO_488 (O_488,N_28275,N_28540);
and UO_489 (O_489,N_28408,N_29504);
and UO_490 (O_490,N_28762,N_28008);
or UO_491 (O_491,N_28615,N_28450);
xnor UO_492 (O_492,N_28447,N_29845);
or UO_493 (O_493,N_29376,N_28988);
or UO_494 (O_494,N_28987,N_29494);
nand UO_495 (O_495,N_28241,N_28736);
nor UO_496 (O_496,N_29814,N_28536);
or UO_497 (O_497,N_28185,N_29777);
nand UO_498 (O_498,N_29809,N_29063);
and UO_499 (O_499,N_28330,N_29394);
and UO_500 (O_500,N_28488,N_28515);
and UO_501 (O_501,N_29661,N_29570);
nor UO_502 (O_502,N_29373,N_29217);
and UO_503 (O_503,N_29289,N_28183);
xor UO_504 (O_504,N_29436,N_29999);
and UO_505 (O_505,N_28496,N_29497);
or UO_506 (O_506,N_29499,N_28312);
xor UO_507 (O_507,N_28525,N_29976);
xnor UO_508 (O_508,N_28579,N_28472);
nor UO_509 (O_509,N_28320,N_28526);
xor UO_510 (O_510,N_28110,N_28745);
nand UO_511 (O_511,N_29012,N_28257);
or UO_512 (O_512,N_28341,N_29608);
nor UO_513 (O_513,N_28356,N_29263);
and UO_514 (O_514,N_28179,N_28835);
and UO_515 (O_515,N_28688,N_29707);
xnor UO_516 (O_516,N_28190,N_28379);
nand UO_517 (O_517,N_29102,N_28597);
and UO_518 (O_518,N_29270,N_29577);
and UO_519 (O_519,N_28385,N_29788);
xnor UO_520 (O_520,N_29804,N_29205);
and UO_521 (O_521,N_29272,N_29381);
or UO_522 (O_522,N_29774,N_28638);
xor UO_523 (O_523,N_28741,N_28547);
nand UO_524 (O_524,N_28021,N_28826);
nor UO_525 (O_525,N_29161,N_28905);
xor UO_526 (O_526,N_29470,N_28562);
and UO_527 (O_527,N_29190,N_29683);
xor UO_528 (O_528,N_29117,N_29869);
nor UO_529 (O_529,N_29603,N_28797);
or UO_530 (O_530,N_28914,N_28532);
nand UO_531 (O_531,N_29652,N_29266);
xor UO_532 (O_532,N_29691,N_29392);
nand UO_533 (O_533,N_29654,N_28703);
and UO_534 (O_534,N_29558,N_29208);
nand UO_535 (O_535,N_28203,N_29518);
and UO_536 (O_536,N_28112,N_28660);
nor UO_537 (O_537,N_29911,N_29246);
nand UO_538 (O_538,N_28947,N_29286);
xor UO_539 (O_539,N_29810,N_29947);
or UO_540 (O_540,N_29967,N_29403);
nand UO_541 (O_541,N_29946,N_28350);
xnor UO_542 (O_542,N_29053,N_28582);
and UO_543 (O_543,N_29891,N_28939);
xor UO_544 (O_544,N_28742,N_29511);
and UO_545 (O_545,N_29961,N_29594);
and UO_546 (O_546,N_29129,N_29188);
or UO_547 (O_547,N_28724,N_29014);
nand UO_548 (O_548,N_28963,N_29301);
and UO_549 (O_549,N_29896,N_28535);
nor UO_550 (O_550,N_28279,N_29458);
nand UO_551 (O_551,N_28414,N_28436);
xor UO_552 (O_552,N_28693,N_28163);
xnor UO_553 (O_553,N_28238,N_29406);
and UO_554 (O_554,N_28135,N_29714);
and UO_555 (O_555,N_29285,N_28951);
nor UO_556 (O_556,N_28941,N_28334);
and UO_557 (O_557,N_28619,N_29480);
and UO_558 (O_558,N_28046,N_29220);
xnor UO_559 (O_559,N_29447,N_28696);
nor UO_560 (O_560,N_29914,N_28133);
nand UO_561 (O_561,N_28094,N_29625);
xor UO_562 (O_562,N_28215,N_29773);
nand UO_563 (O_563,N_29614,N_28684);
or UO_564 (O_564,N_28666,N_28752);
and UO_565 (O_565,N_28728,N_28698);
and UO_566 (O_566,N_29122,N_29546);
nand UO_567 (O_567,N_29132,N_29527);
xor UO_568 (O_568,N_29582,N_28451);
and UO_569 (O_569,N_29956,N_29399);
xor UO_570 (O_570,N_28454,N_28957);
nand UO_571 (O_571,N_28050,N_28971);
xor UO_572 (O_572,N_29051,N_28670);
xnor UO_573 (O_573,N_29482,N_29962);
nor UO_574 (O_574,N_28671,N_28317);
nand UO_575 (O_575,N_29249,N_28177);
and UO_576 (O_576,N_28263,N_29715);
xor UO_577 (O_577,N_29200,N_29860);
nand UO_578 (O_578,N_29586,N_28925);
xor UO_579 (O_579,N_29550,N_28503);
or UO_580 (O_580,N_28920,N_28459);
xor UO_581 (O_581,N_28534,N_29475);
xor UO_582 (O_582,N_28059,N_29225);
nand UO_583 (O_583,N_29139,N_29187);
nand UO_584 (O_584,N_28997,N_29833);
xor UO_585 (O_585,N_28722,N_28700);
or UO_586 (O_586,N_29643,N_29657);
nand UO_587 (O_587,N_29549,N_29261);
or UO_588 (O_588,N_29018,N_28719);
nor UO_589 (O_589,N_28283,N_28923);
and UO_590 (O_590,N_28252,N_29886);
xnor UO_591 (O_591,N_29857,N_28250);
xnor UO_592 (O_592,N_29679,N_28580);
and UO_593 (O_593,N_29388,N_28995);
nor UO_594 (O_594,N_28544,N_28895);
xor UO_595 (O_595,N_28376,N_28016);
nand UO_596 (O_596,N_29748,N_28097);
nand UO_597 (O_597,N_29321,N_28704);
nor UO_598 (O_598,N_29015,N_28431);
xnor UO_599 (O_599,N_28701,N_29214);
or UO_600 (O_600,N_29737,N_29926);
nor UO_601 (O_601,N_29924,N_28585);
xor UO_602 (O_602,N_29853,N_29743);
xor UO_603 (O_603,N_28429,N_29749);
nor UO_604 (O_604,N_28519,N_28194);
or UO_605 (O_605,N_29581,N_28888);
nand UO_606 (O_606,N_28390,N_29808);
nand UO_607 (O_607,N_28750,N_28643);
or UO_608 (O_608,N_29409,N_28499);
xor UO_609 (O_609,N_29355,N_28840);
xnor UO_610 (O_610,N_29684,N_28772);
and UO_611 (O_611,N_29753,N_28322);
nor UO_612 (O_612,N_29400,N_28522);
and UO_613 (O_613,N_29973,N_29561);
nor UO_614 (O_614,N_28766,N_29491);
and UO_615 (O_615,N_28469,N_28166);
or UO_616 (O_616,N_28251,N_29486);
nor UO_617 (O_617,N_29326,N_28281);
or UO_618 (O_618,N_29345,N_28911);
nand UO_619 (O_619,N_29135,N_28799);
xnor UO_620 (O_620,N_29663,N_29405);
xnor UO_621 (O_621,N_29798,N_28087);
nor UO_622 (O_622,N_28456,N_29787);
nor UO_623 (O_623,N_29359,N_28933);
xor UO_624 (O_624,N_28073,N_28419);
and UO_625 (O_625,N_28744,N_29095);
and UO_626 (O_626,N_28676,N_28020);
nor UO_627 (O_627,N_29950,N_28395);
nand UO_628 (O_628,N_29451,N_29839);
or UO_629 (O_629,N_28943,N_28555);
nor UO_630 (O_630,N_28563,N_28273);
or UO_631 (O_631,N_29107,N_29852);
and UO_632 (O_632,N_29781,N_29516);
or UO_633 (O_633,N_29726,N_28148);
nand UO_634 (O_634,N_29880,N_29477);
nor UO_635 (O_635,N_28919,N_29325);
xnor UO_636 (O_636,N_29466,N_29917);
nor UO_637 (O_637,N_29865,N_29492);
nand UO_638 (O_638,N_28834,N_28151);
nand UO_639 (O_639,N_29016,N_28595);
nor UO_640 (O_640,N_28113,N_28727);
nor UO_641 (O_641,N_29338,N_28378);
and UO_642 (O_642,N_29627,N_28782);
or UO_643 (O_643,N_29525,N_29112);
or UO_644 (O_644,N_29507,N_29262);
nor UO_645 (O_645,N_29189,N_29929);
nand UO_646 (O_646,N_29151,N_28815);
or UO_647 (O_647,N_28424,N_29086);
xor UO_648 (O_648,N_29698,N_28402);
and UO_649 (O_649,N_29361,N_28137);
or UO_650 (O_650,N_29881,N_29423);
or UO_651 (O_651,N_29920,N_29358);
xnor UO_652 (O_652,N_29185,N_29945);
xnor UO_653 (O_653,N_29314,N_28301);
xor UO_654 (O_654,N_28278,N_28434);
xnor UO_655 (O_655,N_28106,N_29687);
nand UO_656 (O_656,N_28743,N_28890);
xnor UO_657 (O_657,N_29957,N_28868);
and UO_658 (O_658,N_28841,N_28363);
and UO_659 (O_659,N_28767,N_29454);
or UO_660 (O_660,N_29879,N_28318);
nand UO_661 (O_661,N_29887,N_28590);
xnor UO_662 (O_662,N_29476,N_29149);
nor UO_663 (O_663,N_28874,N_28901);
and UO_664 (O_664,N_29308,N_28566);
nand UO_665 (O_665,N_29522,N_28889);
xor UO_666 (O_666,N_28088,N_28753);
nand UO_667 (O_667,N_29248,N_28045);
nand UO_668 (O_668,N_29771,N_29069);
and UO_669 (O_669,N_28418,N_28658);
and UO_670 (O_670,N_29949,N_28864);
and UO_671 (O_671,N_29972,N_28410);
nor UO_672 (O_672,N_28607,N_28255);
xor UO_673 (O_673,N_28172,N_29983);
nor UO_674 (O_674,N_28667,N_28787);
and UO_675 (O_675,N_28168,N_28411);
xor UO_676 (O_676,N_29283,N_28626);
nand UO_677 (O_677,N_28343,N_29383);
and UO_678 (O_678,N_29596,N_29257);
and UO_679 (O_679,N_28899,N_29763);
and UO_680 (O_680,N_28131,N_28605);
and UO_681 (O_681,N_28965,N_29512);
nand UO_682 (O_682,N_29884,N_29585);
xnor UO_683 (O_683,N_28594,N_29607);
or UO_684 (O_684,N_29142,N_29092);
nor UO_685 (O_685,N_28372,N_28804);
xnor UO_686 (O_686,N_28847,N_29412);
and UO_687 (O_687,N_29418,N_28391);
nand UO_688 (O_688,N_29310,N_29938);
nand UO_689 (O_689,N_29889,N_28293);
or UO_690 (O_690,N_28773,N_29855);
xor UO_691 (O_691,N_29057,N_29899);
or UO_692 (O_692,N_29562,N_28624);
xnor UO_693 (O_693,N_28476,N_28426);
or UO_694 (O_694,N_28896,N_29784);
nand UO_695 (O_695,N_28770,N_29331);
nand UO_696 (O_696,N_29713,N_29859);
or UO_697 (O_697,N_29680,N_29382);
nor UO_698 (O_698,N_28075,N_28557);
nor UO_699 (O_699,N_29082,N_28175);
or UO_700 (O_700,N_28329,N_29640);
xor UO_701 (O_701,N_28368,N_28010);
xor UO_702 (O_702,N_28836,N_28827);
xnor UO_703 (O_703,N_28508,N_29935);
nor UO_704 (O_704,N_29202,N_28335);
and UO_705 (O_705,N_28090,N_28453);
xor UO_706 (O_706,N_28918,N_29617);
nand UO_707 (O_707,N_28935,N_29137);
or UO_708 (O_708,N_29370,N_28810);
xor UO_709 (O_709,N_28710,N_28970);
and UO_710 (O_710,N_29277,N_29828);
or UO_711 (O_711,N_28141,N_29979);
and UO_712 (O_712,N_29576,N_28413);
nor UO_713 (O_713,N_28400,N_29264);
and UO_714 (O_714,N_28859,N_29241);
nand UO_715 (O_715,N_29731,N_28467);
and UO_716 (O_716,N_29123,N_29221);
or UO_717 (O_717,N_29103,N_28856);
nand UO_718 (O_718,N_29542,N_29148);
and UO_719 (O_719,N_28846,N_28602);
nand UO_720 (O_720,N_29256,N_28830);
nand UO_721 (O_721,N_28785,N_28180);
or UO_722 (O_722,N_29020,N_28060);
or UO_723 (O_723,N_29259,N_28748);
or UO_724 (O_724,N_28216,N_28292);
nor UO_725 (O_725,N_29783,N_28833);
xnor UO_726 (O_726,N_29991,N_28316);
nand UO_727 (O_727,N_28460,N_28078);
xor UO_728 (O_728,N_29980,N_29592);
nor UO_729 (O_729,N_28475,N_29579);
or UO_730 (O_730,N_29425,N_29572);
nor UO_731 (O_731,N_28154,N_29735);
xor UO_732 (O_732,N_29158,N_29634);
nand UO_733 (O_733,N_29831,N_29992);
xor UO_734 (O_734,N_28937,N_28117);
nor UO_735 (O_735,N_28873,N_28553);
or UO_736 (O_736,N_28699,N_29702);
or UO_737 (O_737,N_28406,N_29811);
nand UO_738 (O_738,N_28596,N_28375);
nand UO_739 (O_739,N_29912,N_28734);
xor UO_740 (O_740,N_28729,N_28808);
or UO_741 (O_741,N_28373,N_29667);
xnor UO_742 (O_742,N_29328,N_29066);
nand UO_743 (O_743,N_28646,N_28342);
and UO_744 (O_744,N_28319,N_28306);
xnor UO_745 (O_745,N_29415,N_29159);
nand UO_746 (O_746,N_29333,N_29642);
or UO_747 (O_747,N_28119,N_29952);
or UO_748 (O_748,N_28367,N_28015);
xnor UO_749 (O_749,N_29140,N_28079);
and UO_750 (O_750,N_28760,N_29006);
and UO_751 (O_751,N_29437,N_29755);
and UO_752 (O_752,N_29067,N_29354);
nand UO_753 (O_753,N_28796,N_28972);
nand UO_754 (O_754,N_28051,N_29160);
nand UO_755 (O_755,N_28277,N_28200);
xor UO_756 (O_756,N_28246,N_29419);
and UO_757 (O_757,N_28583,N_28984);
nor UO_758 (O_758,N_29569,N_29688);
and UO_759 (O_759,N_29469,N_28956);
or UO_760 (O_760,N_28668,N_29033);
xor UO_761 (O_761,N_28839,N_28993);
xnor UO_762 (O_762,N_29513,N_29849);
and UO_763 (O_763,N_28274,N_29847);
nand UO_764 (O_764,N_29127,N_28260);
nand UO_765 (O_765,N_29723,N_29832);
nor UO_766 (O_766,N_28417,N_29404);
and UO_767 (O_767,N_29121,N_29556);
and UO_768 (O_768,N_29670,N_28793);
and UO_769 (O_769,N_29689,N_29770);
and UO_770 (O_770,N_28305,N_29375);
xnor UO_771 (O_771,N_28853,N_28249);
nand UO_772 (O_772,N_29794,N_28944);
or UO_773 (O_773,N_29843,N_28442);
nand UO_774 (O_774,N_29198,N_29292);
xor UO_775 (O_775,N_29329,N_29174);
xnor UO_776 (O_776,N_29369,N_29462);
or UO_777 (O_777,N_29255,N_28739);
xnor UO_778 (O_778,N_29467,N_29922);
nor UO_779 (O_779,N_28327,N_28758);
xnor UO_780 (O_780,N_28731,N_29232);
and UO_781 (O_781,N_28043,N_28572);
xnor UO_782 (O_782,N_29138,N_29776);
or UO_783 (O_783,N_28820,N_29258);
and UO_784 (O_784,N_29900,N_29495);
xor UO_785 (O_785,N_28653,N_28908);
or UO_786 (O_786,N_28374,N_28510);
or UO_787 (O_787,N_28380,N_28101);
or UO_788 (O_788,N_29530,N_29901);
nand UO_789 (O_789,N_28308,N_28284);
and UO_790 (O_790,N_29574,N_29762);
xnor UO_791 (O_791,N_29079,N_29357);
xor UO_792 (O_792,N_29481,N_29867);
nor UO_793 (O_793,N_29593,N_29472);
and UO_794 (O_794,N_29461,N_29352);
xnor UO_795 (O_795,N_29772,N_28794);
nand UO_796 (O_796,N_28576,N_28256);
nor UO_797 (O_797,N_29128,N_29829);
xnor UO_798 (O_798,N_28495,N_29315);
and UO_799 (O_799,N_29005,N_28309);
nor UO_800 (O_800,N_28887,N_29806);
xor UO_801 (O_801,N_28074,N_28691);
xor UO_802 (O_802,N_28062,N_29610);
nand UO_803 (O_803,N_29414,N_28816);
xor UO_804 (O_804,N_29010,N_29802);
or UO_805 (O_805,N_28798,N_28272);
xnor UO_806 (O_806,N_28616,N_28589);
and UO_807 (O_807,N_29746,N_28118);
nor UO_808 (O_808,N_28440,N_28479);
xor UO_809 (O_809,N_29062,N_29742);
nand UO_810 (O_810,N_28264,N_29250);
or UO_811 (O_811,N_29538,N_28210);
or UO_812 (O_812,N_28359,N_28514);
nor UO_813 (O_813,N_28880,N_29164);
or UO_814 (O_814,N_29540,N_29998);
nor UO_815 (O_815,N_28560,N_28423);
and UO_816 (O_816,N_29143,N_28130);
nand UO_817 (O_817,N_28574,N_28001);
xnor UO_818 (O_818,N_29969,N_28123);
nand UO_819 (O_819,N_29557,N_29152);
and UO_820 (O_820,N_28103,N_29488);
nand UO_821 (O_821,N_28192,N_28362);
nor UO_822 (O_822,N_29296,N_29609);
or UO_823 (O_823,N_29796,N_29903);
and UO_824 (O_824,N_29459,N_28952);
nor UO_825 (O_825,N_28382,N_28254);
nor UO_826 (O_826,N_29003,N_28152);
or UO_827 (O_827,N_29632,N_29800);
nor UO_828 (O_828,N_29931,N_29641);
or UO_829 (O_829,N_29895,N_29982);
xnor UO_830 (O_830,N_29101,N_29176);
or UO_831 (O_831,N_29812,N_29274);
xnor UO_832 (O_832,N_28550,N_28921);
xor UO_833 (O_833,N_28337,N_28630);
or UO_834 (O_834,N_28695,N_28239);
or UO_835 (O_835,N_28371,N_29087);
nor UO_836 (O_836,N_28028,N_29180);
xor UO_837 (O_837,N_29169,N_28310);
and UO_838 (O_838,N_28898,N_28954);
nand UO_839 (O_839,N_29701,N_28575);
xnor UO_840 (O_840,N_29751,N_29630);
nor UO_841 (O_841,N_28093,N_28869);
nand UO_842 (O_842,N_28664,N_29621);
nand UO_843 (O_843,N_29080,N_29212);
xor UO_844 (O_844,N_28682,N_28913);
nor UO_845 (O_845,N_29060,N_28121);
nand UO_846 (O_846,N_29994,N_29184);
and UO_847 (O_847,N_28628,N_29428);
xnor UO_848 (O_848,N_28871,N_29181);
or UO_849 (O_849,N_29226,N_28370);
nor UO_850 (O_850,N_29826,N_29276);
and UO_851 (O_851,N_28683,N_28768);
or UO_852 (O_852,N_29615,N_29613);
nor UO_853 (O_853,N_28386,N_28866);
nand UO_854 (O_854,N_28243,N_29573);
nand UO_855 (O_855,N_28631,N_28791);
nor UO_856 (O_856,N_29932,N_29334);
nor UO_857 (O_857,N_28222,N_28759);
or UO_858 (O_858,N_29937,N_28953);
nor UO_859 (O_859,N_29455,N_29064);
or UO_860 (O_860,N_29785,N_28035);
nor UO_861 (O_861,N_28702,N_28132);
nand UO_862 (O_862,N_28614,N_29268);
nor UO_863 (O_863,N_29058,N_29975);
or UO_864 (O_864,N_29449,N_29827);
nor UO_865 (O_865,N_29700,N_28115);
xnor UO_866 (O_866,N_28205,N_29690);
and UO_867 (O_867,N_29666,N_28931);
xor UO_868 (O_868,N_28485,N_29309);
xor UO_869 (O_869,N_29211,N_28848);
or UO_870 (O_870,N_28116,N_28080);
xnor UO_871 (O_871,N_28314,N_28912);
and UO_872 (O_872,N_28019,N_29209);
xor UO_873 (O_873,N_29186,N_29893);
or UO_874 (O_874,N_28754,N_28795);
xnor UO_875 (O_875,N_28612,N_28740);
nor UO_876 (O_876,N_29923,N_28809);
xnor UO_877 (O_877,N_28030,N_28573);
or UO_878 (O_878,N_29758,N_28926);
or UO_879 (O_879,N_28248,N_28765);
nor UO_880 (O_880,N_28242,N_28055);
and UO_881 (O_881,N_28082,N_28213);
nor UO_882 (O_882,N_28297,N_29588);
or UO_883 (O_883,N_29821,N_29435);
nand UO_884 (O_884,N_29756,N_28184);
or UO_885 (O_885,N_28824,N_29243);
xnor UO_886 (O_886,N_29769,N_28143);
nor UO_887 (O_887,N_28518,N_28640);
or UO_888 (O_888,N_28686,N_28679);
nand UO_889 (O_889,N_28063,N_29088);
xnor UO_890 (O_890,N_28542,N_29638);
nand UO_891 (O_891,N_28038,N_29997);
xor UO_892 (O_892,N_29028,N_28058);
nor UO_893 (O_893,N_29813,N_28511);
xor UO_894 (O_894,N_29442,N_28850);
and UO_895 (O_895,N_29534,N_28067);
or UO_896 (O_896,N_29948,N_29675);
and UO_897 (O_897,N_29987,N_28966);
and UO_898 (O_898,N_28302,N_29921);
xnor UO_899 (O_899,N_28202,N_28549);
and UO_900 (O_900,N_29323,N_29305);
nand UO_901 (O_901,N_29054,N_28909);
or UO_902 (O_902,N_29861,N_29106);
xor UO_903 (O_903,N_29531,N_28076);
nor UO_904 (O_904,N_29070,N_28746);
or UO_905 (O_905,N_29368,N_28025);
nor UO_906 (O_906,N_28672,N_29598);
nand UO_907 (O_907,N_28570,N_29222);
and UO_908 (O_908,N_29963,N_28998);
and UO_909 (O_909,N_28401,N_28715);
and UO_910 (O_910,N_28040,N_29877);
nand UO_911 (O_911,N_28173,N_29233);
nand UO_912 (O_912,N_29692,N_28564);
and UO_913 (O_913,N_28307,N_29432);
nor UO_914 (O_914,N_28441,N_28621);
xnor UO_915 (O_915,N_29535,N_29767);
or UO_916 (O_916,N_29479,N_29822);
or UO_917 (O_917,N_29940,N_29620);
or UO_918 (O_918,N_29709,N_29508);
nor UO_919 (O_919,N_28945,N_29633);
nor UO_920 (O_920,N_28290,N_29231);
nor UO_921 (O_921,N_29313,N_28383);
nand UO_922 (O_922,N_28081,N_28528);
nand UO_923 (O_923,N_29336,N_29782);
nor UO_924 (O_924,N_29023,N_28611);
and UO_925 (O_925,N_29396,N_29706);
or UO_926 (O_926,N_28285,N_28633);
nor UO_927 (O_927,N_29350,N_28229);
and UO_928 (O_928,N_28347,N_29793);
or UO_929 (O_929,N_29364,N_29393);
xnor UO_930 (O_930,N_28494,N_28346);
xor UO_931 (O_931,N_29104,N_28120);
xnor UO_932 (O_932,N_28286,N_29939);
or UO_933 (O_933,N_29658,N_29733);
and UO_934 (O_934,N_29818,N_29196);
and UO_935 (O_935,N_28022,N_28315);
xnor UO_936 (O_936,N_28042,N_29545);
xnor UO_937 (O_937,N_29349,N_29335);
nand UO_938 (O_938,N_29560,N_29874);
nand UO_939 (O_939,N_29705,N_29267);
nor UO_940 (O_940,N_29130,N_29113);
nor UO_941 (O_941,N_28169,N_28217);
or UO_942 (O_942,N_28942,N_29677);
nand UO_943 (O_943,N_29599,N_29167);
and UO_944 (O_944,N_29116,N_28709);
xnor UO_945 (O_945,N_28344,N_29754);
nand UO_946 (O_946,N_29339,N_29031);
nand UO_947 (O_947,N_28870,N_28160);
nand UO_948 (O_948,N_29445,N_29386);
nand UO_949 (O_949,N_28452,N_28707);
xnor UO_950 (O_950,N_28207,N_28398);
xor UO_951 (O_951,N_29269,N_28832);
nand UO_952 (O_952,N_28338,N_29566);
and UO_953 (O_953,N_28477,N_29988);
and UO_954 (O_954,N_29529,N_29251);
nor UO_955 (O_955,N_28652,N_28845);
xnor UO_956 (O_956,N_28403,N_28761);
xor UO_957 (O_957,N_29942,N_28443);
nor UO_958 (O_958,N_29380,N_28681);
xor UO_959 (O_959,N_28086,N_29863);
nand UO_960 (O_960,N_28858,N_29303);
xor UO_961 (O_961,N_29318,N_28950);
or UO_962 (O_962,N_28070,N_29503);
and UO_963 (O_963,N_29197,N_29192);
or UO_964 (O_964,N_28095,N_28655);
or UO_965 (O_965,N_28468,N_28973);
xnor UO_966 (O_966,N_28718,N_29265);
or UO_967 (O_967,N_29179,N_28838);
or UO_968 (O_968,N_28420,N_29401);
nand UO_969 (O_969,N_29085,N_28224);
xnor UO_970 (O_970,N_28259,N_29595);
nand UO_971 (O_971,N_28775,N_29120);
nor UO_972 (O_972,N_28044,N_28747);
nand UO_973 (O_973,N_28780,N_28144);
xor UO_974 (O_974,N_28340,N_29565);
or UO_975 (O_975,N_29098,N_29223);
and UO_976 (O_976,N_28048,N_28578);
and UO_977 (O_977,N_28940,N_29906);
or UO_978 (O_978,N_29686,N_28157);
and UO_979 (O_979,N_29984,N_29575);
xor UO_980 (O_980,N_29864,N_28697);
xnor UO_981 (O_981,N_28262,N_28529);
nor UO_982 (O_982,N_28066,N_29320);
and UO_983 (O_983,N_29457,N_29510);
and UO_984 (O_984,N_29155,N_28685);
nand UO_985 (O_985,N_29439,N_29996);
xnor UO_986 (O_986,N_28934,N_28608);
xor UO_987 (O_987,N_28065,N_29521);
nor UO_988 (O_988,N_29240,N_28158);
or UO_989 (O_989,N_29841,N_28831);
and UO_990 (O_990,N_28521,N_28072);
nor UO_991 (O_991,N_28730,N_28394);
nor UO_992 (O_992,N_29587,N_28541);
and UO_993 (O_993,N_29175,N_29768);
nand UO_994 (O_994,N_29100,N_28181);
and UO_995 (O_995,N_28280,N_29780);
and UO_996 (O_996,N_29765,N_29150);
and UO_997 (O_997,N_28189,N_29493);
nand UO_998 (O_998,N_28480,N_28527);
nand UO_999 (O_999,N_29750,N_29974);
nor UO_1000 (O_1000,N_28112,N_28781);
and UO_1001 (O_1001,N_29756,N_29504);
or UO_1002 (O_1002,N_29554,N_29529);
nor UO_1003 (O_1003,N_28084,N_28076);
or UO_1004 (O_1004,N_28861,N_28639);
xnor UO_1005 (O_1005,N_28024,N_29061);
xor UO_1006 (O_1006,N_29512,N_28049);
and UO_1007 (O_1007,N_29634,N_29022);
nand UO_1008 (O_1008,N_28814,N_28010);
nor UO_1009 (O_1009,N_29315,N_29945);
nor UO_1010 (O_1010,N_28412,N_29390);
nor UO_1011 (O_1011,N_28179,N_29765);
nand UO_1012 (O_1012,N_28479,N_28147);
nand UO_1013 (O_1013,N_29421,N_28152);
nor UO_1014 (O_1014,N_29175,N_28952);
nand UO_1015 (O_1015,N_28539,N_28675);
xor UO_1016 (O_1016,N_29103,N_29515);
and UO_1017 (O_1017,N_29531,N_28619);
nand UO_1018 (O_1018,N_29745,N_28130);
and UO_1019 (O_1019,N_29553,N_28360);
nand UO_1020 (O_1020,N_29093,N_29126);
nand UO_1021 (O_1021,N_28899,N_28499);
and UO_1022 (O_1022,N_28466,N_29817);
nand UO_1023 (O_1023,N_28311,N_28754);
nor UO_1024 (O_1024,N_28382,N_28856);
and UO_1025 (O_1025,N_29380,N_29109);
or UO_1026 (O_1026,N_28112,N_29310);
nand UO_1027 (O_1027,N_29900,N_28536);
nand UO_1028 (O_1028,N_29541,N_28320);
nand UO_1029 (O_1029,N_29197,N_28048);
and UO_1030 (O_1030,N_29714,N_29108);
and UO_1031 (O_1031,N_28145,N_28750);
nand UO_1032 (O_1032,N_28655,N_28784);
or UO_1033 (O_1033,N_28635,N_28038);
and UO_1034 (O_1034,N_29418,N_28654);
and UO_1035 (O_1035,N_28663,N_29464);
xnor UO_1036 (O_1036,N_29539,N_29958);
nor UO_1037 (O_1037,N_28489,N_29579);
nor UO_1038 (O_1038,N_29263,N_29618);
or UO_1039 (O_1039,N_29436,N_29167);
nor UO_1040 (O_1040,N_29813,N_29555);
xor UO_1041 (O_1041,N_28812,N_29617);
xor UO_1042 (O_1042,N_28638,N_28983);
nor UO_1043 (O_1043,N_28728,N_28929);
nand UO_1044 (O_1044,N_29645,N_29591);
or UO_1045 (O_1045,N_29961,N_28606);
nor UO_1046 (O_1046,N_28098,N_28981);
or UO_1047 (O_1047,N_29299,N_28611);
xor UO_1048 (O_1048,N_29733,N_28466);
xor UO_1049 (O_1049,N_28498,N_29509);
or UO_1050 (O_1050,N_29061,N_29893);
or UO_1051 (O_1051,N_29869,N_29413);
nor UO_1052 (O_1052,N_28503,N_29334);
nor UO_1053 (O_1053,N_29871,N_29212);
or UO_1054 (O_1054,N_28431,N_29006);
xnor UO_1055 (O_1055,N_29782,N_29686);
or UO_1056 (O_1056,N_28396,N_28709);
nor UO_1057 (O_1057,N_29536,N_29731);
or UO_1058 (O_1058,N_28410,N_28156);
and UO_1059 (O_1059,N_28380,N_28108);
or UO_1060 (O_1060,N_29234,N_29038);
and UO_1061 (O_1061,N_28265,N_29328);
nand UO_1062 (O_1062,N_28234,N_29907);
xnor UO_1063 (O_1063,N_29161,N_29090);
or UO_1064 (O_1064,N_28554,N_29095);
nand UO_1065 (O_1065,N_28239,N_29693);
xor UO_1066 (O_1066,N_29355,N_29765);
nand UO_1067 (O_1067,N_29759,N_28541);
xnor UO_1068 (O_1068,N_29469,N_29232);
xor UO_1069 (O_1069,N_29227,N_28577);
xnor UO_1070 (O_1070,N_29128,N_29238);
or UO_1071 (O_1071,N_29023,N_28019);
or UO_1072 (O_1072,N_28495,N_29693);
or UO_1073 (O_1073,N_28394,N_29148);
nand UO_1074 (O_1074,N_29355,N_28285);
nor UO_1075 (O_1075,N_29806,N_29210);
nand UO_1076 (O_1076,N_28562,N_28805);
nor UO_1077 (O_1077,N_29690,N_28737);
or UO_1078 (O_1078,N_28104,N_29404);
nor UO_1079 (O_1079,N_28551,N_29208);
xnor UO_1080 (O_1080,N_28734,N_29174);
xor UO_1081 (O_1081,N_29179,N_28721);
nand UO_1082 (O_1082,N_28071,N_29126);
nor UO_1083 (O_1083,N_29887,N_28410);
xnor UO_1084 (O_1084,N_29212,N_29991);
and UO_1085 (O_1085,N_28963,N_29904);
nor UO_1086 (O_1086,N_28164,N_28038);
nor UO_1087 (O_1087,N_28481,N_29269);
nand UO_1088 (O_1088,N_29424,N_29520);
nand UO_1089 (O_1089,N_29192,N_29944);
nand UO_1090 (O_1090,N_29903,N_29657);
xor UO_1091 (O_1091,N_28379,N_29802);
nand UO_1092 (O_1092,N_28982,N_29326);
xnor UO_1093 (O_1093,N_28502,N_28516);
nand UO_1094 (O_1094,N_29766,N_29350);
nor UO_1095 (O_1095,N_28634,N_29964);
nand UO_1096 (O_1096,N_29593,N_28545);
xor UO_1097 (O_1097,N_28936,N_28297);
and UO_1098 (O_1098,N_29466,N_28469);
nor UO_1099 (O_1099,N_29111,N_29899);
xnor UO_1100 (O_1100,N_29613,N_28740);
nor UO_1101 (O_1101,N_28491,N_29761);
or UO_1102 (O_1102,N_28185,N_28335);
nand UO_1103 (O_1103,N_28641,N_28106);
nand UO_1104 (O_1104,N_29180,N_29610);
xor UO_1105 (O_1105,N_28325,N_28079);
and UO_1106 (O_1106,N_28293,N_29978);
nand UO_1107 (O_1107,N_28129,N_28787);
nand UO_1108 (O_1108,N_28902,N_29533);
or UO_1109 (O_1109,N_29339,N_28695);
and UO_1110 (O_1110,N_29843,N_29056);
nor UO_1111 (O_1111,N_28017,N_29840);
and UO_1112 (O_1112,N_29962,N_29150);
nor UO_1113 (O_1113,N_28798,N_28218);
nand UO_1114 (O_1114,N_28138,N_29866);
nand UO_1115 (O_1115,N_29985,N_28820);
nor UO_1116 (O_1116,N_28081,N_29604);
or UO_1117 (O_1117,N_29204,N_28860);
xnor UO_1118 (O_1118,N_28095,N_28282);
nor UO_1119 (O_1119,N_29705,N_28226);
and UO_1120 (O_1120,N_28037,N_28697);
nor UO_1121 (O_1121,N_28967,N_29880);
nand UO_1122 (O_1122,N_29865,N_29545);
nand UO_1123 (O_1123,N_28844,N_29096);
nor UO_1124 (O_1124,N_28306,N_28295);
or UO_1125 (O_1125,N_29174,N_28106);
nor UO_1126 (O_1126,N_28903,N_28111);
nand UO_1127 (O_1127,N_29911,N_29794);
nand UO_1128 (O_1128,N_28602,N_29515);
xor UO_1129 (O_1129,N_28861,N_29025);
xnor UO_1130 (O_1130,N_28130,N_29036);
or UO_1131 (O_1131,N_28142,N_29732);
nor UO_1132 (O_1132,N_28416,N_29171);
and UO_1133 (O_1133,N_29363,N_29504);
nand UO_1134 (O_1134,N_29800,N_29892);
xor UO_1135 (O_1135,N_29921,N_28320);
xnor UO_1136 (O_1136,N_29300,N_29706);
or UO_1137 (O_1137,N_29758,N_29441);
xnor UO_1138 (O_1138,N_28334,N_29525);
and UO_1139 (O_1139,N_28658,N_29875);
and UO_1140 (O_1140,N_29132,N_29457);
and UO_1141 (O_1141,N_29851,N_29364);
xor UO_1142 (O_1142,N_29913,N_28328);
or UO_1143 (O_1143,N_28575,N_29543);
nand UO_1144 (O_1144,N_28295,N_28757);
xnor UO_1145 (O_1145,N_28148,N_29966);
or UO_1146 (O_1146,N_28609,N_28107);
xnor UO_1147 (O_1147,N_29193,N_28742);
nand UO_1148 (O_1148,N_29332,N_29893);
or UO_1149 (O_1149,N_29362,N_28985);
nand UO_1150 (O_1150,N_29273,N_29853);
and UO_1151 (O_1151,N_29441,N_29242);
and UO_1152 (O_1152,N_28538,N_29304);
nor UO_1153 (O_1153,N_28801,N_28818);
and UO_1154 (O_1154,N_29337,N_29474);
nand UO_1155 (O_1155,N_28839,N_28983);
xor UO_1156 (O_1156,N_29700,N_28605);
or UO_1157 (O_1157,N_28160,N_28190);
and UO_1158 (O_1158,N_29670,N_28864);
nand UO_1159 (O_1159,N_28304,N_28057);
or UO_1160 (O_1160,N_28746,N_29851);
or UO_1161 (O_1161,N_29757,N_29574);
or UO_1162 (O_1162,N_29725,N_29492);
nor UO_1163 (O_1163,N_29521,N_28579);
and UO_1164 (O_1164,N_28502,N_28386);
xnor UO_1165 (O_1165,N_28920,N_28405);
nor UO_1166 (O_1166,N_29565,N_28585);
or UO_1167 (O_1167,N_29447,N_29288);
nand UO_1168 (O_1168,N_28915,N_28509);
nor UO_1169 (O_1169,N_29592,N_28993);
nand UO_1170 (O_1170,N_28428,N_28320);
nor UO_1171 (O_1171,N_28186,N_28975);
nand UO_1172 (O_1172,N_28082,N_28904);
nor UO_1173 (O_1173,N_28492,N_28935);
or UO_1174 (O_1174,N_29630,N_28860);
xor UO_1175 (O_1175,N_28588,N_28212);
xnor UO_1176 (O_1176,N_29169,N_29376);
or UO_1177 (O_1177,N_28440,N_28605);
nand UO_1178 (O_1178,N_28830,N_29999);
xnor UO_1179 (O_1179,N_28461,N_28334);
nand UO_1180 (O_1180,N_29438,N_29050);
and UO_1181 (O_1181,N_28812,N_29870);
xor UO_1182 (O_1182,N_28484,N_28933);
and UO_1183 (O_1183,N_29223,N_28127);
nor UO_1184 (O_1184,N_28628,N_29590);
nand UO_1185 (O_1185,N_29946,N_28818);
xor UO_1186 (O_1186,N_29097,N_28293);
or UO_1187 (O_1187,N_28892,N_28466);
nand UO_1188 (O_1188,N_28127,N_29005);
nand UO_1189 (O_1189,N_29836,N_29363);
or UO_1190 (O_1190,N_28518,N_29469);
nor UO_1191 (O_1191,N_29213,N_28160);
and UO_1192 (O_1192,N_29701,N_28651);
or UO_1193 (O_1193,N_29532,N_28524);
or UO_1194 (O_1194,N_28133,N_29503);
or UO_1195 (O_1195,N_28382,N_29997);
xnor UO_1196 (O_1196,N_28564,N_29826);
or UO_1197 (O_1197,N_28010,N_28435);
nand UO_1198 (O_1198,N_29557,N_29374);
and UO_1199 (O_1199,N_28059,N_29352);
xor UO_1200 (O_1200,N_28973,N_29089);
xnor UO_1201 (O_1201,N_29292,N_28925);
nand UO_1202 (O_1202,N_29030,N_28294);
nor UO_1203 (O_1203,N_28927,N_29403);
xor UO_1204 (O_1204,N_29737,N_29837);
or UO_1205 (O_1205,N_28040,N_28950);
nor UO_1206 (O_1206,N_29276,N_29131);
nand UO_1207 (O_1207,N_28690,N_29423);
nor UO_1208 (O_1208,N_29941,N_29070);
or UO_1209 (O_1209,N_29996,N_29763);
and UO_1210 (O_1210,N_29978,N_29851);
nor UO_1211 (O_1211,N_28601,N_29492);
or UO_1212 (O_1212,N_29274,N_29314);
nand UO_1213 (O_1213,N_28313,N_29275);
nor UO_1214 (O_1214,N_29800,N_28751);
or UO_1215 (O_1215,N_29815,N_29476);
or UO_1216 (O_1216,N_28248,N_28651);
or UO_1217 (O_1217,N_29979,N_28665);
and UO_1218 (O_1218,N_28280,N_28063);
nand UO_1219 (O_1219,N_28065,N_29507);
and UO_1220 (O_1220,N_29900,N_29959);
or UO_1221 (O_1221,N_28235,N_28281);
or UO_1222 (O_1222,N_28128,N_29992);
nand UO_1223 (O_1223,N_28374,N_28620);
nand UO_1224 (O_1224,N_28377,N_29010);
nand UO_1225 (O_1225,N_28621,N_28687);
xnor UO_1226 (O_1226,N_29499,N_29565);
or UO_1227 (O_1227,N_28137,N_28485);
nor UO_1228 (O_1228,N_28601,N_28357);
and UO_1229 (O_1229,N_28135,N_28965);
and UO_1230 (O_1230,N_29706,N_29346);
xor UO_1231 (O_1231,N_29031,N_29296);
nor UO_1232 (O_1232,N_28729,N_29791);
or UO_1233 (O_1233,N_28262,N_29982);
or UO_1234 (O_1234,N_29715,N_29806);
nand UO_1235 (O_1235,N_29060,N_29135);
or UO_1236 (O_1236,N_28277,N_28648);
nand UO_1237 (O_1237,N_28234,N_29554);
nand UO_1238 (O_1238,N_29999,N_28096);
nor UO_1239 (O_1239,N_29352,N_28187);
nand UO_1240 (O_1240,N_28650,N_29549);
and UO_1241 (O_1241,N_29579,N_28329);
or UO_1242 (O_1242,N_29502,N_28070);
or UO_1243 (O_1243,N_29683,N_28314);
xor UO_1244 (O_1244,N_28002,N_29788);
or UO_1245 (O_1245,N_29708,N_29980);
and UO_1246 (O_1246,N_28951,N_28576);
or UO_1247 (O_1247,N_29644,N_28205);
or UO_1248 (O_1248,N_28725,N_29420);
and UO_1249 (O_1249,N_29883,N_29057);
nor UO_1250 (O_1250,N_28301,N_28564);
xor UO_1251 (O_1251,N_28447,N_28866);
xor UO_1252 (O_1252,N_28557,N_28731);
and UO_1253 (O_1253,N_29891,N_28618);
xnor UO_1254 (O_1254,N_28133,N_28631);
xnor UO_1255 (O_1255,N_29818,N_28195);
nand UO_1256 (O_1256,N_29060,N_29468);
or UO_1257 (O_1257,N_29707,N_29076);
nand UO_1258 (O_1258,N_29934,N_29248);
nand UO_1259 (O_1259,N_28811,N_28110);
or UO_1260 (O_1260,N_29151,N_28126);
xor UO_1261 (O_1261,N_29949,N_28632);
nor UO_1262 (O_1262,N_28716,N_29158);
nand UO_1263 (O_1263,N_29777,N_29752);
xor UO_1264 (O_1264,N_28408,N_29587);
and UO_1265 (O_1265,N_29586,N_28090);
or UO_1266 (O_1266,N_29996,N_28203);
or UO_1267 (O_1267,N_29668,N_29152);
xor UO_1268 (O_1268,N_28466,N_29317);
xnor UO_1269 (O_1269,N_29241,N_29939);
and UO_1270 (O_1270,N_29204,N_29502);
xor UO_1271 (O_1271,N_28140,N_29586);
and UO_1272 (O_1272,N_28366,N_29185);
nand UO_1273 (O_1273,N_29371,N_29637);
and UO_1274 (O_1274,N_28458,N_28371);
xnor UO_1275 (O_1275,N_29946,N_28146);
and UO_1276 (O_1276,N_29514,N_29997);
xor UO_1277 (O_1277,N_28265,N_28623);
and UO_1278 (O_1278,N_29955,N_29167);
and UO_1279 (O_1279,N_29477,N_29328);
or UO_1280 (O_1280,N_28034,N_29682);
nand UO_1281 (O_1281,N_28484,N_28162);
or UO_1282 (O_1282,N_28424,N_29434);
nand UO_1283 (O_1283,N_29356,N_28130);
xor UO_1284 (O_1284,N_29181,N_29621);
xnor UO_1285 (O_1285,N_28116,N_28937);
and UO_1286 (O_1286,N_28359,N_28336);
nand UO_1287 (O_1287,N_29159,N_28250);
or UO_1288 (O_1288,N_29830,N_29967);
nor UO_1289 (O_1289,N_29498,N_29047);
and UO_1290 (O_1290,N_28202,N_28884);
nand UO_1291 (O_1291,N_28091,N_28797);
nor UO_1292 (O_1292,N_29613,N_28894);
nor UO_1293 (O_1293,N_29131,N_29871);
nor UO_1294 (O_1294,N_28155,N_29550);
and UO_1295 (O_1295,N_28128,N_28357);
and UO_1296 (O_1296,N_29378,N_28976);
xor UO_1297 (O_1297,N_28506,N_29141);
xnor UO_1298 (O_1298,N_29668,N_28389);
nor UO_1299 (O_1299,N_29089,N_29873);
or UO_1300 (O_1300,N_29186,N_29347);
xor UO_1301 (O_1301,N_29916,N_29969);
xnor UO_1302 (O_1302,N_28525,N_28199);
or UO_1303 (O_1303,N_29276,N_29891);
nor UO_1304 (O_1304,N_29323,N_29230);
nand UO_1305 (O_1305,N_28328,N_28899);
nor UO_1306 (O_1306,N_28285,N_29882);
nand UO_1307 (O_1307,N_28724,N_29794);
nand UO_1308 (O_1308,N_28189,N_28062);
nor UO_1309 (O_1309,N_28751,N_29395);
nand UO_1310 (O_1310,N_28851,N_28497);
nand UO_1311 (O_1311,N_28136,N_28695);
nor UO_1312 (O_1312,N_29555,N_28876);
and UO_1313 (O_1313,N_28115,N_29232);
or UO_1314 (O_1314,N_28908,N_28348);
nor UO_1315 (O_1315,N_29999,N_29373);
xor UO_1316 (O_1316,N_29092,N_28657);
nor UO_1317 (O_1317,N_29172,N_28035);
and UO_1318 (O_1318,N_28998,N_29824);
nor UO_1319 (O_1319,N_28447,N_29913);
nand UO_1320 (O_1320,N_29806,N_29370);
nand UO_1321 (O_1321,N_29188,N_28768);
nor UO_1322 (O_1322,N_28002,N_28464);
and UO_1323 (O_1323,N_28111,N_29330);
and UO_1324 (O_1324,N_29313,N_28992);
nor UO_1325 (O_1325,N_29844,N_29491);
nor UO_1326 (O_1326,N_28841,N_29349);
nand UO_1327 (O_1327,N_29899,N_29220);
nand UO_1328 (O_1328,N_28760,N_29621);
xnor UO_1329 (O_1329,N_28174,N_29109);
xnor UO_1330 (O_1330,N_29539,N_28136);
xor UO_1331 (O_1331,N_28220,N_29435);
nor UO_1332 (O_1332,N_28592,N_28204);
nand UO_1333 (O_1333,N_29908,N_29927);
xnor UO_1334 (O_1334,N_29469,N_29159);
xnor UO_1335 (O_1335,N_29103,N_28772);
nand UO_1336 (O_1336,N_29142,N_28833);
nor UO_1337 (O_1337,N_29505,N_29956);
and UO_1338 (O_1338,N_29173,N_29098);
xor UO_1339 (O_1339,N_28099,N_29271);
and UO_1340 (O_1340,N_29407,N_28028);
or UO_1341 (O_1341,N_29408,N_28606);
xor UO_1342 (O_1342,N_28255,N_29292);
and UO_1343 (O_1343,N_29046,N_29197);
xor UO_1344 (O_1344,N_29760,N_28976);
nand UO_1345 (O_1345,N_28695,N_29532);
nand UO_1346 (O_1346,N_28075,N_28408);
xor UO_1347 (O_1347,N_28885,N_28355);
xor UO_1348 (O_1348,N_28492,N_28554);
xor UO_1349 (O_1349,N_29098,N_28303);
and UO_1350 (O_1350,N_28478,N_29352);
nor UO_1351 (O_1351,N_28590,N_28658);
or UO_1352 (O_1352,N_28107,N_29723);
nor UO_1353 (O_1353,N_29344,N_29921);
and UO_1354 (O_1354,N_29895,N_28496);
xnor UO_1355 (O_1355,N_28673,N_28529);
xnor UO_1356 (O_1356,N_28521,N_28446);
nor UO_1357 (O_1357,N_29349,N_29294);
or UO_1358 (O_1358,N_29746,N_28811);
nor UO_1359 (O_1359,N_28540,N_28743);
nand UO_1360 (O_1360,N_29340,N_29013);
nor UO_1361 (O_1361,N_28512,N_28243);
and UO_1362 (O_1362,N_28162,N_28759);
or UO_1363 (O_1363,N_28608,N_28376);
nand UO_1364 (O_1364,N_28700,N_29095);
nor UO_1365 (O_1365,N_28606,N_28797);
or UO_1366 (O_1366,N_28184,N_29406);
nor UO_1367 (O_1367,N_29403,N_29135);
or UO_1368 (O_1368,N_29931,N_29988);
nand UO_1369 (O_1369,N_29206,N_29424);
nand UO_1370 (O_1370,N_28374,N_29679);
xnor UO_1371 (O_1371,N_28568,N_29615);
nand UO_1372 (O_1372,N_28640,N_28224);
nand UO_1373 (O_1373,N_28587,N_28663);
xor UO_1374 (O_1374,N_29039,N_29834);
and UO_1375 (O_1375,N_28450,N_29413);
xnor UO_1376 (O_1376,N_29903,N_29139);
nor UO_1377 (O_1377,N_28696,N_28990);
or UO_1378 (O_1378,N_29319,N_28944);
nand UO_1379 (O_1379,N_29202,N_28115);
nor UO_1380 (O_1380,N_29828,N_28292);
nand UO_1381 (O_1381,N_29511,N_28680);
nor UO_1382 (O_1382,N_29169,N_29730);
xor UO_1383 (O_1383,N_29437,N_29824);
nor UO_1384 (O_1384,N_29962,N_28945);
nand UO_1385 (O_1385,N_28378,N_29284);
or UO_1386 (O_1386,N_28373,N_29770);
and UO_1387 (O_1387,N_29659,N_29823);
or UO_1388 (O_1388,N_29207,N_29577);
nand UO_1389 (O_1389,N_28987,N_28158);
nand UO_1390 (O_1390,N_28969,N_29377);
nand UO_1391 (O_1391,N_28976,N_29686);
nand UO_1392 (O_1392,N_28797,N_28727);
and UO_1393 (O_1393,N_28809,N_28039);
and UO_1394 (O_1394,N_28111,N_29913);
xor UO_1395 (O_1395,N_29421,N_28946);
nor UO_1396 (O_1396,N_29846,N_28709);
or UO_1397 (O_1397,N_29784,N_29202);
nor UO_1398 (O_1398,N_29852,N_28431);
or UO_1399 (O_1399,N_29758,N_29583);
and UO_1400 (O_1400,N_29063,N_29717);
nand UO_1401 (O_1401,N_29678,N_28527);
nand UO_1402 (O_1402,N_29218,N_29696);
nor UO_1403 (O_1403,N_29080,N_29564);
or UO_1404 (O_1404,N_29691,N_29862);
nor UO_1405 (O_1405,N_28041,N_28116);
or UO_1406 (O_1406,N_28802,N_29935);
nand UO_1407 (O_1407,N_28392,N_29457);
nand UO_1408 (O_1408,N_29397,N_29063);
and UO_1409 (O_1409,N_28921,N_29615);
nand UO_1410 (O_1410,N_29647,N_29356);
and UO_1411 (O_1411,N_28126,N_29058);
or UO_1412 (O_1412,N_29080,N_28797);
or UO_1413 (O_1413,N_29739,N_29442);
and UO_1414 (O_1414,N_28052,N_28819);
or UO_1415 (O_1415,N_29224,N_28462);
and UO_1416 (O_1416,N_28562,N_28048);
xnor UO_1417 (O_1417,N_29716,N_29523);
nor UO_1418 (O_1418,N_28366,N_29779);
and UO_1419 (O_1419,N_29271,N_29290);
nor UO_1420 (O_1420,N_29502,N_28542);
or UO_1421 (O_1421,N_28133,N_28600);
nor UO_1422 (O_1422,N_29186,N_29659);
or UO_1423 (O_1423,N_28839,N_29286);
and UO_1424 (O_1424,N_28347,N_28123);
or UO_1425 (O_1425,N_29041,N_29219);
nor UO_1426 (O_1426,N_28735,N_29505);
and UO_1427 (O_1427,N_28158,N_29906);
nand UO_1428 (O_1428,N_28783,N_28657);
and UO_1429 (O_1429,N_29561,N_28555);
nor UO_1430 (O_1430,N_28166,N_28602);
and UO_1431 (O_1431,N_29245,N_28731);
nand UO_1432 (O_1432,N_28214,N_29273);
or UO_1433 (O_1433,N_29344,N_28003);
nor UO_1434 (O_1434,N_28002,N_28649);
nor UO_1435 (O_1435,N_29045,N_28561);
or UO_1436 (O_1436,N_29976,N_29013);
nand UO_1437 (O_1437,N_28754,N_29245);
or UO_1438 (O_1438,N_28091,N_29187);
nor UO_1439 (O_1439,N_28737,N_29064);
and UO_1440 (O_1440,N_29776,N_29878);
nand UO_1441 (O_1441,N_29248,N_29855);
xnor UO_1442 (O_1442,N_28317,N_29295);
xor UO_1443 (O_1443,N_28834,N_28735);
or UO_1444 (O_1444,N_28509,N_28578);
xnor UO_1445 (O_1445,N_28617,N_29267);
nand UO_1446 (O_1446,N_28477,N_28214);
xor UO_1447 (O_1447,N_29685,N_28852);
and UO_1448 (O_1448,N_29485,N_29138);
and UO_1449 (O_1449,N_28498,N_28339);
nor UO_1450 (O_1450,N_29141,N_29070);
and UO_1451 (O_1451,N_29389,N_28668);
xnor UO_1452 (O_1452,N_29274,N_29459);
nand UO_1453 (O_1453,N_28806,N_29358);
nand UO_1454 (O_1454,N_29908,N_29696);
nand UO_1455 (O_1455,N_28953,N_28244);
or UO_1456 (O_1456,N_29932,N_29830);
or UO_1457 (O_1457,N_29475,N_29451);
and UO_1458 (O_1458,N_28285,N_28820);
nor UO_1459 (O_1459,N_29300,N_28600);
or UO_1460 (O_1460,N_28663,N_29402);
or UO_1461 (O_1461,N_29704,N_29753);
xor UO_1462 (O_1462,N_28506,N_28628);
or UO_1463 (O_1463,N_28886,N_28606);
xor UO_1464 (O_1464,N_29952,N_28468);
xor UO_1465 (O_1465,N_29390,N_29230);
xnor UO_1466 (O_1466,N_29252,N_28267);
xor UO_1467 (O_1467,N_29480,N_29348);
and UO_1468 (O_1468,N_28098,N_29914);
nor UO_1469 (O_1469,N_29320,N_29433);
nand UO_1470 (O_1470,N_28434,N_28719);
and UO_1471 (O_1471,N_28031,N_29069);
or UO_1472 (O_1472,N_28805,N_28998);
xnor UO_1473 (O_1473,N_28524,N_28145);
xnor UO_1474 (O_1474,N_29443,N_29757);
and UO_1475 (O_1475,N_29996,N_28870);
nor UO_1476 (O_1476,N_28280,N_28560);
or UO_1477 (O_1477,N_29700,N_28364);
nor UO_1478 (O_1478,N_28122,N_28743);
nor UO_1479 (O_1479,N_29944,N_28222);
xor UO_1480 (O_1480,N_29204,N_29123);
nand UO_1481 (O_1481,N_29087,N_29723);
nor UO_1482 (O_1482,N_29878,N_28759);
nor UO_1483 (O_1483,N_28587,N_28354);
xor UO_1484 (O_1484,N_29032,N_29357);
or UO_1485 (O_1485,N_29299,N_29196);
and UO_1486 (O_1486,N_29694,N_28444);
nor UO_1487 (O_1487,N_28881,N_28440);
xor UO_1488 (O_1488,N_29225,N_29672);
xor UO_1489 (O_1489,N_28338,N_29037);
nand UO_1490 (O_1490,N_28741,N_29550);
nand UO_1491 (O_1491,N_28858,N_28038);
xnor UO_1492 (O_1492,N_28340,N_29172);
nand UO_1493 (O_1493,N_28852,N_28218);
and UO_1494 (O_1494,N_28369,N_28921);
xor UO_1495 (O_1495,N_28993,N_29444);
or UO_1496 (O_1496,N_29682,N_28075);
or UO_1497 (O_1497,N_29389,N_28050);
nand UO_1498 (O_1498,N_29079,N_28125);
nand UO_1499 (O_1499,N_29477,N_28951);
and UO_1500 (O_1500,N_28044,N_28921);
and UO_1501 (O_1501,N_29820,N_29917);
and UO_1502 (O_1502,N_29058,N_29772);
and UO_1503 (O_1503,N_28951,N_28386);
and UO_1504 (O_1504,N_28843,N_28591);
nand UO_1505 (O_1505,N_29044,N_29583);
xnor UO_1506 (O_1506,N_28204,N_29173);
nand UO_1507 (O_1507,N_28245,N_28844);
or UO_1508 (O_1508,N_28613,N_29722);
xnor UO_1509 (O_1509,N_29204,N_29881);
or UO_1510 (O_1510,N_28323,N_29363);
xnor UO_1511 (O_1511,N_28283,N_29594);
and UO_1512 (O_1512,N_29365,N_28705);
nor UO_1513 (O_1513,N_28634,N_29161);
nor UO_1514 (O_1514,N_29719,N_29279);
nand UO_1515 (O_1515,N_29370,N_28111);
nand UO_1516 (O_1516,N_28910,N_28311);
or UO_1517 (O_1517,N_29745,N_28881);
and UO_1518 (O_1518,N_29618,N_29935);
nand UO_1519 (O_1519,N_29141,N_28163);
and UO_1520 (O_1520,N_29028,N_29346);
nand UO_1521 (O_1521,N_28439,N_28096);
xor UO_1522 (O_1522,N_28223,N_28665);
nand UO_1523 (O_1523,N_28342,N_29194);
xnor UO_1524 (O_1524,N_29187,N_29424);
xor UO_1525 (O_1525,N_29620,N_28330);
xnor UO_1526 (O_1526,N_28162,N_29818);
nor UO_1527 (O_1527,N_29238,N_29105);
and UO_1528 (O_1528,N_29116,N_28176);
nor UO_1529 (O_1529,N_29517,N_29560);
xor UO_1530 (O_1530,N_28603,N_29753);
and UO_1531 (O_1531,N_28143,N_28712);
xnor UO_1532 (O_1532,N_28662,N_28328);
nor UO_1533 (O_1533,N_29850,N_28340);
or UO_1534 (O_1534,N_28140,N_28710);
or UO_1535 (O_1535,N_29119,N_28610);
or UO_1536 (O_1536,N_29700,N_29361);
xor UO_1537 (O_1537,N_29382,N_28641);
nor UO_1538 (O_1538,N_28784,N_28828);
nor UO_1539 (O_1539,N_28525,N_29128);
nand UO_1540 (O_1540,N_28293,N_28071);
nor UO_1541 (O_1541,N_28115,N_29146);
nor UO_1542 (O_1542,N_29790,N_29504);
or UO_1543 (O_1543,N_28582,N_29108);
and UO_1544 (O_1544,N_29645,N_29716);
xor UO_1545 (O_1545,N_29646,N_28245);
nor UO_1546 (O_1546,N_29735,N_29927);
or UO_1547 (O_1547,N_29820,N_28421);
nor UO_1548 (O_1548,N_29280,N_29134);
nor UO_1549 (O_1549,N_29663,N_29368);
xor UO_1550 (O_1550,N_29627,N_28468);
nor UO_1551 (O_1551,N_28054,N_29050);
or UO_1552 (O_1552,N_28588,N_29036);
and UO_1553 (O_1553,N_28449,N_29191);
or UO_1554 (O_1554,N_29891,N_28087);
nor UO_1555 (O_1555,N_29532,N_28102);
xor UO_1556 (O_1556,N_29539,N_29637);
xnor UO_1557 (O_1557,N_28247,N_29484);
xor UO_1558 (O_1558,N_28589,N_28622);
or UO_1559 (O_1559,N_28343,N_29280);
xnor UO_1560 (O_1560,N_28939,N_28930);
nand UO_1561 (O_1561,N_29563,N_28608);
nand UO_1562 (O_1562,N_28521,N_29146);
nor UO_1563 (O_1563,N_29633,N_28361);
nand UO_1564 (O_1564,N_28082,N_29211);
nand UO_1565 (O_1565,N_29182,N_28854);
and UO_1566 (O_1566,N_29046,N_28553);
or UO_1567 (O_1567,N_29570,N_28715);
and UO_1568 (O_1568,N_29759,N_29264);
nor UO_1569 (O_1569,N_29825,N_29675);
or UO_1570 (O_1570,N_29382,N_29481);
xor UO_1571 (O_1571,N_28757,N_29167);
and UO_1572 (O_1572,N_28847,N_29149);
or UO_1573 (O_1573,N_29594,N_28332);
xnor UO_1574 (O_1574,N_28967,N_29841);
nand UO_1575 (O_1575,N_28418,N_28645);
nand UO_1576 (O_1576,N_29484,N_28387);
nand UO_1577 (O_1577,N_29843,N_28969);
or UO_1578 (O_1578,N_28437,N_29260);
nand UO_1579 (O_1579,N_29340,N_29785);
xnor UO_1580 (O_1580,N_28390,N_29398);
nand UO_1581 (O_1581,N_28718,N_28227);
or UO_1582 (O_1582,N_29949,N_28950);
nand UO_1583 (O_1583,N_29158,N_28656);
nor UO_1584 (O_1584,N_29861,N_29993);
nor UO_1585 (O_1585,N_28857,N_29853);
nand UO_1586 (O_1586,N_29240,N_29763);
and UO_1587 (O_1587,N_29528,N_29980);
nand UO_1588 (O_1588,N_28845,N_29446);
and UO_1589 (O_1589,N_28698,N_28110);
xnor UO_1590 (O_1590,N_29212,N_29537);
nor UO_1591 (O_1591,N_29981,N_29520);
and UO_1592 (O_1592,N_29422,N_28764);
xnor UO_1593 (O_1593,N_28335,N_28742);
nor UO_1594 (O_1594,N_29756,N_28903);
nor UO_1595 (O_1595,N_29839,N_28087);
nand UO_1596 (O_1596,N_28821,N_29804);
or UO_1597 (O_1597,N_28405,N_28912);
and UO_1598 (O_1598,N_28707,N_28948);
xnor UO_1599 (O_1599,N_28959,N_29656);
nand UO_1600 (O_1600,N_29833,N_28559);
and UO_1601 (O_1601,N_29971,N_28790);
nand UO_1602 (O_1602,N_29926,N_28178);
nand UO_1603 (O_1603,N_29172,N_29145);
and UO_1604 (O_1604,N_29937,N_28884);
or UO_1605 (O_1605,N_28231,N_28712);
and UO_1606 (O_1606,N_29819,N_29768);
and UO_1607 (O_1607,N_29637,N_29207);
or UO_1608 (O_1608,N_28292,N_28911);
nand UO_1609 (O_1609,N_29473,N_29958);
xor UO_1610 (O_1610,N_28750,N_28673);
and UO_1611 (O_1611,N_28316,N_29427);
and UO_1612 (O_1612,N_29885,N_28238);
xnor UO_1613 (O_1613,N_29684,N_29737);
or UO_1614 (O_1614,N_29141,N_29847);
and UO_1615 (O_1615,N_29716,N_28525);
and UO_1616 (O_1616,N_28003,N_29286);
or UO_1617 (O_1617,N_28198,N_28180);
or UO_1618 (O_1618,N_29491,N_28241);
nor UO_1619 (O_1619,N_28252,N_29087);
nor UO_1620 (O_1620,N_28599,N_28800);
nor UO_1621 (O_1621,N_28373,N_28826);
xor UO_1622 (O_1622,N_29257,N_29922);
or UO_1623 (O_1623,N_28369,N_28789);
or UO_1624 (O_1624,N_29851,N_28199);
or UO_1625 (O_1625,N_29199,N_28953);
nand UO_1626 (O_1626,N_29730,N_28188);
or UO_1627 (O_1627,N_29535,N_29967);
and UO_1628 (O_1628,N_28660,N_28434);
and UO_1629 (O_1629,N_29950,N_29260);
nand UO_1630 (O_1630,N_29382,N_28904);
or UO_1631 (O_1631,N_29724,N_28830);
xnor UO_1632 (O_1632,N_28869,N_29842);
or UO_1633 (O_1633,N_28958,N_28414);
xor UO_1634 (O_1634,N_29753,N_29207);
nand UO_1635 (O_1635,N_28037,N_28352);
and UO_1636 (O_1636,N_28795,N_29011);
nand UO_1637 (O_1637,N_29668,N_29124);
nand UO_1638 (O_1638,N_29737,N_29422);
nand UO_1639 (O_1639,N_29006,N_29647);
or UO_1640 (O_1640,N_29426,N_28527);
nor UO_1641 (O_1641,N_29669,N_29290);
xor UO_1642 (O_1642,N_29558,N_29347);
nand UO_1643 (O_1643,N_28340,N_28353);
nor UO_1644 (O_1644,N_29455,N_28681);
and UO_1645 (O_1645,N_29339,N_29697);
xor UO_1646 (O_1646,N_29758,N_28091);
nand UO_1647 (O_1647,N_28232,N_29147);
nand UO_1648 (O_1648,N_28071,N_28182);
nor UO_1649 (O_1649,N_28054,N_28939);
nor UO_1650 (O_1650,N_28844,N_29302);
nand UO_1651 (O_1651,N_29654,N_28332);
and UO_1652 (O_1652,N_28526,N_29820);
or UO_1653 (O_1653,N_28814,N_29735);
xor UO_1654 (O_1654,N_28285,N_29050);
and UO_1655 (O_1655,N_29518,N_28271);
nand UO_1656 (O_1656,N_28394,N_28488);
or UO_1657 (O_1657,N_29991,N_28791);
nor UO_1658 (O_1658,N_28728,N_28484);
or UO_1659 (O_1659,N_29756,N_29918);
or UO_1660 (O_1660,N_28877,N_29000);
nor UO_1661 (O_1661,N_29119,N_28644);
and UO_1662 (O_1662,N_28482,N_28187);
nor UO_1663 (O_1663,N_28888,N_29684);
xor UO_1664 (O_1664,N_29545,N_29888);
and UO_1665 (O_1665,N_29841,N_28306);
nand UO_1666 (O_1666,N_29498,N_29858);
and UO_1667 (O_1667,N_28081,N_29386);
xnor UO_1668 (O_1668,N_28130,N_29308);
and UO_1669 (O_1669,N_29619,N_28837);
nor UO_1670 (O_1670,N_29619,N_29209);
or UO_1671 (O_1671,N_29322,N_28653);
xnor UO_1672 (O_1672,N_28780,N_28310);
nand UO_1673 (O_1673,N_28266,N_29722);
and UO_1674 (O_1674,N_29306,N_28429);
nand UO_1675 (O_1675,N_28503,N_29466);
nor UO_1676 (O_1676,N_29930,N_29924);
xor UO_1677 (O_1677,N_28054,N_29318);
xor UO_1678 (O_1678,N_29523,N_28570);
nor UO_1679 (O_1679,N_28516,N_29366);
and UO_1680 (O_1680,N_28780,N_28831);
xor UO_1681 (O_1681,N_29193,N_28177);
or UO_1682 (O_1682,N_28666,N_29161);
nor UO_1683 (O_1683,N_29544,N_29284);
and UO_1684 (O_1684,N_29006,N_28280);
nor UO_1685 (O_1685,N_29704,N_28245);
nand UO_1686 (O_1686,N_29216,N_28241);
nor UO_1687 (O_1687,N_28005,N_28366);
nor UO_1688 (O_1688,N_29756,N_29953);
nor UO_1689 (O_1689,N_28454,N_28013);
xor UO_1690 (O_1690,N_28248,N_29292);
and UO_1691 (O_1691,N_29070,N_29740);
nor UO_1692 (O_1692,N_28953,N_28983);
and UO_1693 (O_1693,N_28542,N_28712);
or UO_1694 (O_1694,N_28033,N_29605);
and UO_1695 (O_1695,N_29451,N_29974);
nor UO_1696 (O_1696,N_28002,N_28657);
xor UO_1697 (O_1697,N_28679,N_29373);
nor UO_1698 (O_1698,N_29753,N_28344);
xnor UO_1699 (O_1699,N_28290,N_28965);
xnor UO_1700 (O_1700,N_29304,N_29394);
or UO_1701 (O_1701,N_29981,N_29420);
nand UO_1702 (O_1702,N_28930,N_28897);
xnor UO_1703 (O_1703,N_29668,N_29951);
and UO_1704 (O_1704,N_28944,N_29476);
or UO_1705 (O_1705,N_29975,N_29019);
and UO_1706 (O_1706,N_29767,N_29566);
and UO_1707 (O_1707,N_29976,N_29208);
nor UO_1708 (O_1708,N_28681,N_29740);
nand UO_1709 (O_1709,N_29684,N_29084);
nand UO_1710 (O_1710,N_29051,N_29501);
nand UO_1711 (O_1711,N_28816,N_28187);
xnor UO_1712 (O_1712,N_29757,N_29328);
and UO_1713 (O_1713,N_29971,N_29394);
nor UO_1714 (O_1714,N_29093,N_29942);
nor UO_1715 (O_1715,N_28536,N_29816);
and UO_1716 (O_1716,N_29127,N_28817);
xor UO_1717 (O_1717,N_29119,N_28230);
and UO_1718 (O_1718,N_28271,N_29521);
xnor UO_1719 (O_1719,N_28378,N_29832);
nand UO_1720 (O_1720,N_29900,N_29629);
or UO_1721 (O_1721,N_28983,N_28547);
or UO_1722 (O_1722,N_28706,N_29651);
or UO_1723 (O_1723,N_28758,N_29392);
nand UO_1724 (O_1724,N_28212,N_28811);
and UO_1725 (O_1725,N_29976,N_28755);
or UO_1726 (O_1726,N_29490,N_29151);
and UO_1727 (O_1727,N_29549,N_29193);
xnor UO_1728 (O_1728,N_29569,N_29645);
nor UO_1729 (O_1729,N_29335,N_29184);
and UO_1730 (O_1730,N_29537,N_29127);
or UO_1731 (O_1731,N_29526,N_28208);
nand UO_1732 (O_1732,N_28384,N_28543);
xor UO_1733 (O_1733,N_28334,N_28506);
and UO_1734 (O_1734,N_28583,N_28265);
or UO_1735 (O_1735,N_28805,N_29257);
nand UO_1736 (O_1736,N_29051,N_28236);
nand UO_1737 (O_1737,N_28408,N_29342);
and UO_1738 (O_1738,N_29523,N_28648);
xor UO_1739 (O_1739,N_29991,N_28398);
nand UO_1740 (O_1740,N_28034,N_28127);
or UO_1741 (O_1741,N_28561,N_28710);
and UO_1742 (O_1742,N_28871,N_29212);
and UO_1743 (O_1743,N_29637,N_28585);
nand UO_1744 (O_1744,N_28034,N_29285);
nor UO_1745 (O_1745,N_29682,N_28170);
or UO_1746 (O_1746,N_28599,N_28920);
nand UO_1747 (O_1747,N_29084,N_28026);
nor UO_1748 (O_1748,N_29913,N_29829);
nand UO_1749 (O_1749,N_29658,N_29490);
nor UO_1750 (O_1750,N_28725,N_29509);
or UO_1751 (O_1751,N_28146,N_29620);
and UO_1752 (O_1752,N_28210,N_29171);
nor UO_1753 (O_1753,N_29556,N_28715);
nand UO_1754 (O_1754,N_29109,N_29792);
and UO_1755 (O_1755,N_29871,N_28956);
nand UO_1756 (O_1756,N_29648,N_28895);
or UO_1757 (O_1757,N_29195,N_28261);
nor UO_1758 (O_1758,N_29096,N_29952);
and UO_1759 (O_1759,N_28123,N_29702);
or UO_1760 (O_1760,N_28949,N_28182);
xor UO_1761 (O_1761,N_28006,N_29177);
or UO_1762 (O_1762,N_29130,N_29723);
or UO_1763 (O_1763,N_29053,N_29588);
nor UO_1764 (O_1764,N_29105,N_28441);
xnor UO_1765 (O_1765,N_29914,N_28921);
xor UO_1766 (O_1766,N_29097,N_28851);
or UO_1767 (O_1767,N_29366,N_29849);
or UO_1768 (O_1768,N_28040,N_29405);
or UO_1769 (O_1769,N_29832,N_28350);
and UO_1770 (O_1770,N_28856,N_29609);
or UO_1771 (O_1771,N_29272,N_29324);
nor UO_1772 (O_1772,N_29510,N_28895);
nand UO_1773 (O_1773,N_29957,N_29973);
nand UO_1774 (O_1774,N_29894,N_29125);
nor UO_1775 (O_1775,N_28447,N_29265);
nand UO_1776 (O_1776,N_28502,N_28143);
xnor UO_1777 (O_1777,N_28888,N_28883);
or UO_1778 (O_1778,N_28296,N_29477);
nor UO_1779 (O_1779,N_28179,N_29368);
or UO_1780 (O_1780,N_29400,N_29254);
and UO_1781 (O_1781,N_28566,N_29661);
nand UO_1782 (O_1782,N_28849,N_29871);
nor UO_1783 (O_1783,N_28421,N_28945);
nand UO_1784 (O_1784,N_28193,N_28934);
xor UO_1785 (O_1785,N_29455,N_29631);
xor UO_1786 (O_1786,N_28237,N_29423);
or UO_1787 (O_1787,N_28541,N_28012);
xnor UO_1788 (O_1788,N_29607,N_29139);
and UO_1789 (O_1789,N_29251,N_29680);
nand UO_1790 (O_1790,N_29508,N_29906);
nand UO_1791 (O_1791,N_29362,N_29095);
or UO_1792 (O_1792,N_28813,N_29885);
or UO_1793 (O_1793,N_29359,N_29258);
and UO_1794 (O_1794,N_28855,N_28478);
nor UO_1795 (O_1795,N_28690,N_29575);
nor UO_1796 (O_1796,N_28034,N_29205);
and UO_1797 (O_1797,N_28589,N_28967);
xor UO_1798 (O_1798,N_29432,N_28897);
or UO_1799 (O_1799,N_28328,N_29903);
or UO_1800 (O_1800,N_28075,N_29135);
xnor UO_1801 (O_1801,N_29081,N_28047);
nand UO_1802 (O_1802,N_28262,N_29438);
or UO_1803 (O_1803,N_28185,N_29313);
xnor UO_1804 (O_1804,N_29219,N_28274);
nand UO_1805 (O_1805,N_29397,N_28373);
or UO_1806 (O_1806,N_29023,N_28968);
xnor UO_1807 (O_1807,N_28204,N_29495);
xor UO_1808 (O_1808,N_29839,N_28958);
and UO_1809 (O_1809,N_28112,N_28782);
and UO_1810 (O_1810,N_29068,N_28808);
or UO_1811 (O_1811,N_29558,N_29518);
xor UO_1812 (O_1812,N_28661,N_29543);
nor UO_1813 (O_1813,N_28391,N_29824);
or UO_1814 (O_1814,N_29215,N_29716);
nor UO_1815 (O_1815,N_29585,N_28806);
and UO_1816 (O_1816,N_29961,N_28454);
or UO_1817 (O_1817,N_28885,N_29851);
or UO_1818 (O_1818,N_29181,N_29246);
or UO_1819 (O_1819,N_28500,N_29732);
or UO_1820 (O_1820,N_28819,N_29010);
or UO_1821 (O_1821,N_28717,N_28049);
xor UO_1822 (O_1822,N_28409,N_28121);
nand UO_1823 (O_1823,N_29758,N_29123);
or UO_1824 (O_1824,N_29103,N_29369);
and UO_1825 (O_1825,N_28164,N_29678);
nand UO_1826 (O_1826,N_29357,N_28617);
or UO_1827 (O_1827,N_29903,N_28014);
nor UO_1828 (O_1828,N_28928,N_29101);
and UO_1829 (O_1829,N_29239,N_29105);
nand UO_1830 (O_1830,N_28737,N_28920);
xor UO_1831 (O_1831,N_28576,N_29000);
nand UO_1832 (O_1832,N_28366,N_29306);
xor UO_1833 (O_1833,N_29861,N_28599);
and UO_1834 (O_1834,N_28718,N_28927);
nor UO_1835 (O_1835,N_29014,N_28976);
or UO_1836 (O_1836,N_28153,N_29981);
or UO_1837 (O_1837,N_29124,N_28945);
xor UO_1838 (O_1838,N_29941,N_29643);
and UO_1839 (O_1839,N_28719,N_28681);
xnor UO_1840 (O_1840,N_29377,N_29011);
nor UO_1841 (O_1841,N_28521,N_28260);
nor UO_1842 (O_1842,N_29041,N_29060);
nand UO_1843 (O_1843,N_29629,N_28274);
and UO_1844 (O_1844,N_28284,N_28910);
or UO_1845 (O_1845,N_28891,N_28367);
xnor UO_1846 (O_1846,N_28650,N_28552);
xnor UO_1847 (O_1847,N_28083,N_28591);
nand UO_1848 (O_1848,N_28344,N_29037);
nand UO_1849 (O_1849,N_29973,N_28041);
and UO_1850 (O_1850,N_28936,N_29828);
and UO_1851 (O_1851,N_29455,N_29377);
and UO_1852 (O_1852,N_28593,N_28123);
nand UO_1853 (O_1853,N_28378,N_28152);
and UO_1854 (O_1854,N_28731,N_28492);
nor UO_1855 (O_1855,N_28938,N_28959);
nor UO_1856 (O_1856,N_28501,N_28512);
nand UO_1857 (O_1857,N_29565,N_28156);
nand UO_1858 (O_1858,N_29911,N_29279);
xor UO_1859 (O_1859,N_29912,N_28432);
nor UO_1860 (O_1860,N_29057,N_29941);
or UO_1861 (O_1861,N_28515,N_29490);
and UO_1862 (O_1862,N_28535,N_29935);
or UO_1863 (O_1863,N_29564,N_29732);
nand UO_1864 (O_1864,N_29631,N_29367);
nor UO_1865 (O_1865,N_29980,N_28212);
and UO_1866 (O_1866,N_28929,N_29168);
nor UO_1867 (O_1867,N_28104,N_29532);
nor UO_1868 (O_1868,N_28349,N_28804);
and UO_1869 (O_1869,N_28816,N_28810);
or UO_1870 (O_1870,N_29856,N_29500);
xnor UO_1871 (O_1871,N_28582,N_29209);
nand UO_1872 (O_1872,N_28160,N_28210);
nor UO_1873 (O_1873,N_28719,N_29770);
xor UO_1874 (O_1874,N_28085,N_29066);
xor UO_1875 (O_1875,N_29763,N_28330);
and UO_1876 (O_1876,N_29258,N_29991);
nand UO_1877 (O_1877,N_29673,N_29822);
or UO_1878 (O_1878,N_28347,N_29115);
xnor UO_1879 (O_1879,N_28113,N_29833);
xnor UO_1880 (O_1880,N_29324,N_29689);
nor UO_1881 (O_1881,N_28147,N_29211);
or UO_1882 (O_1882,N_28417,N_28389);
nand UO_1883 (O_1883,N_29409,N_29278);
and UO_1884 (O_1884,N_29134,N_28124);
xnor UO_1885 (O_1885,N_28352,N_29679);
nand UO_1886 (O_1886,N_29614,N_29966);
nand UO_1887 (O_1887,N_29218,N_28533);
nand UO_1888 (O_1888,N_28925,N_29729);
nor UO_1889 (O_1889,N_29159,N_29100);
xor UO_1890 (O_1890,N_29050,N_29252);
or UO_1891 (O_1891,N_28202,N_28976);
xnor UO_1892 (O_1892,N_28400,N_29773);
or UO_1893 (O_1893,N_29272,N_28827);
nand UO_1894 (O_1894,N_28014,N_28317);
and UO_1895 (O_1895,N_28396,N_28417);
or UO_1896 (O_1896,N_28239,N_28779);
nand UO_1897 (O_1897,N_29123,N_29206);
nor UO_1898 (O_1898,N_28862,N_29035);
nor UO_1899 (O_1899,N_29041,N_29170);
nand UO_1900 (O_1900,N_28608,N_28949);
nor UO_1901 (O_1901,N_29799,N_28112);
xnor UO_1902 (O_1902,N_28031,N_29956);
or UO_1903 (O_1903,N_28718,N_28058);
and UO_1904 (O_1904,N_29726,N_29271);
nor UO_1905 (O_1905,N_29724,N_29757);
and UO_1906 (O_1906,N_29767,N_29466);
xnor UO_1907 (O_1907,N_29285,N_29066);
nor UO_1908 (O_1908,N_28754,N_28603);
or UO_1909 (O_1909,N_29099,N_28930);
nand UO_1910 (O_1910,N_29971,N_28910);
or UO_1911 (O_1911,N_29813,N_28262);
and UO_1912 (O_1912,N_28307,N_28334);
nor UO_1913 (O_1913,N_29317,N_28370);
and UO_1914 (O_1914,N_29016,N_28944);
or UO_1915 (O_1915,N_28601,N_29816);
xor UO_1916 (O_1916,N_28420,N_28202);
nand UO_1917 (O_1917,N_28707,N_29930);
and UO_1918 (O_1918,N_29137,N_29340);
and UO_1919 (O_1919,N_28141,N_28136);
xor UO_1920 (O_1920,N_28557,N_29603);
nand UO_1921 (O_1921,N_29529,N_29588);
nand UO_1922 (O_1922,N_28315,N_28892);
and UO_1923 (O_1923,N_29201,N_29013);
and UO_1924 (O_1924,N_29425,N_28640);
and UO_1925 (O_1925,N_28876,N_29972);
xor UO_1926 (O_1926,N_29611,N_28753);
or UO_1927 (O_1927,N_29195,N_29873);
and UO_1928 (O_1928,N_28355,N_29799);
and UO_1929 (O_1929,N_29121,N_29661);
nand UO_1930 (O_1930,N_29843,N_29611);
and UO_1931 (O_1931,N_28626,N_28908);
nor UO_1932 (O_1932,N_28589,N_29049);
xor UO_1933 (O_1933,N_28580,N_29127);
nor UO_1934 (O_1934,N_29910,N_28171);
or UO_1935 (O_1935,N_28479,N_29702);
nand UO_1936 (O_1936,N_29038,N_28762);
and UO_1937 (O_1937,N_29672,N_28932);
or UO_1938 (O_1938,N_28019,N_28306);
or UO_1939 (O_1939,N_28558,N_28040);
nand UO_1940 (O_1940,N_29405,N_29200);
nor UO_1941 (O_1941,N_29051,N_29893);
or UO_1942 (O_1942,N_29634,N_28084);
and UO_1943 (O_1943,N_28878,N_28514);
nand UO_1944 (O_1944,N_28868,N_28860);
xnor UO_1945 (O_1945,N_29637,N_28466);
nor UO_1946 (O_1946,N_28722,N_29619);
and UO_1947 (O_1947,N_29313,N_28825);
xor UO_1948 (O_1948,N_29472,N_29293);
xnor UO_1949 (O_1949,N_29110,N_28229);
xnor UO_1950 (O_1950,N_28737,N_29791);
and UO_1951 (O_1951,N_28076,N_29647);
and UO_1952 (O_1952,N_28410,N_29825);
xor UO_1953 (O_1953,N_28550,N_28367);
xor UO_1954 (O_1954,N_29704,N_29280);
xor UO_1955 (O_1955,N_28227,N_28110);
xor UO_1956 (O_1956,N_28979,N_28943);
nand UO_1957 (O_1957,N_29494,N_29460);
and UO_1958 (O_1958,N_29001,N_29236);
xnor UO_1959 (O_1959,N_29406,N_28086);
or UO_1960 (O_1960,N_28635,N_29252);
nor UO_1961 (O_1961,N_28482,N_28303);
and UO_1962 (O_1962,N_29596,N_29486);
and UO_1963 (O_1963,N_28223,N_28097);
and UO_1964 (O_1964,N_28883,N_28331);
or UO_1965 (O_1965,N_29765,N_29528);
nand UO_1966 (O_1966,N_29997,N_29063);
or UO_1967 (O_1967,N_29796,N_29241);
or UO_1968 (O_1968,N_29085,N_29495);
or UO_1969 (O_1969,N_29869,N_28636);
nand UO_1970 (O_1970,N_29820,N_28051);
nand UO_1971 (O_1971,N_28904,N_29095);
or UO_1972 (O_1972,N_28541,N_29917);
nor UO_1973 (O_1973,N_29165,N_28703);
nor UO_1974 (O_1974,N_29424,N_28627);
xnor UO_1975 (O_1975,N_29256,N_28709);
nand UO_1976 (O_1976,N_29934,N_29606);
nor UO_1977 (O_1977,N_28981,N_28460);
nor UO_1978 (O_1978,N_29275,N_28298);
or UO_1979 (O_1979,N_29248,N_29308);
nor UO_1980 (O_1980,N_28033,N_28661);
and UO_1981 (O_1981,N_28787,N_29520);
and UO_1982 (O_1982,N_28682,N_29255);
nand UO_1983 (O_1983,N_28525,N_29789);
nand UO_1984 (O_1984,N_28797,N_28145);
nand UO_1985 (O_1985,N_28656,N_28946);
and UO_1986 (O_1986,N_29995,N_29713);
xor UO_1987 (O_1987,N_29774,N_29266);
nor UO_1988 (O_1988,N_28434,N_28800);
nand UO_1989 (O_1989,N_29269,N_29187);
and UO_1990 (O_1990,N_29311,N_28006);
nand UO_1991 (O_1991,N_29402,N_29442);
or UO_1992 (O_1992,N_28411,N_29400);
or UO_1993 (O_1993,N_29522,N_28306);
nand UO_1994 (O_1994,N_29710,N_29814);
xor UO_1995 (O_1995,N_29511,N_29334);
nand UO_1996 (O_1996,N_29694,N_29594);
nor UO_1997 (O_1997,N_28209,N_28005);
or UO_1998 (O_1998,N_28849,N_28726);
xnor UO_1999 (O_1999,N_29520,N_28706);
or UO_2000 (O_2000,N_29927,N_29459);
and UO_2001 (O_2001,N_28870,N_28476);
nor UO_2002 (O_2002,N_29129,N_28563);
nand UO_2003 (O_2003,N_28415,N_28155);
nor UO_2004 (O_2004,N_28418,N_29632);
or UO_2005 (O_2005,N_29895,N_29843);
xor UO_2006 (O_2006,N_29816,N_28884);
xnor UO_2007 (O_2007,N_28697,N_28484);
xor UO_2008 (O_2008,N_28081,N_29884);
xor UO_2009 (O_2009,N_29071,N_28010);
or UO_2010 (O_2010,N_28628,N_28502);
nand UO_2011 (O_2011,N_29907,N_29393);
or UO_2012 (O_2012,N_28822,N_28701);
or UO_2013 (O_2013,N_29896,N_29192);
and UO_2014 (O_2014,N_28043,N_28632);
nand UO_2015 (O_2015,N_28190,N_28407);
xor UO_2016 (O_2016,N_28903,N_28190);
nor UO_2017 (O_2017,N_29256,N_28239);
xor UO_2018 (O_2018,N_28232,N_28347);
or UO_2019 (O_2019,N_29521,N_29543);
and UO_2020 (O_2020,N_28638,N_29090);
and UO_2021 (O_2021,N_29264,N_28945);
nand UO_2022 (O_2022,N_29910,N_28351);
xor UO_2023 (O_2023,N_28634,N_28714);
or UO_2024 (O_2024,N_29243,N_28901);
and UO_2025 (O_2025,N_28424,N_29039);
xnor UO_2026 (O_2026,N_29690,N_28302);
nand UO_2027 (O_2027,N_28213,N_29653);
nand UO_2028 (O_2028,N_29383,N_28785);
nor UO_2029 (O_2029,N_28167,N_29314);
or UO_2030 (O_2030,N_28956,N_28175);
xnor UO_2031 (O_2031,N_29508,N_28862);
nand UO_2032 (O_2032,N_29434,N_28159);
or UO_2033 (O_2033,N_29138,N_28505);
xor UO_2034 (O_2034,N_28136,N_28381);
xnor UO_2035 (O_2035,N_29964,N_29018);
nor UO_2036 (O_2036,N_28088,N_28256);
xnor UO_2037 (O_2037,N_28411,N_28215);
and UO_2038 (O_2038,N_28297,N_29651);
xnor UO_2039 (O_2039,N_29149,N_28323);
nor UO_2040 (O_2040,N_28693,N_29608);
xnor UO_2041 (O_2041,N_29555,N_28351);
xnor UO_2042 (O_2042,N_28872,N_28231);
and UO_2043 (O_2043,N_29033,N_29256);
nand UO_2044 (O_2044,N_29265,N_29163);
xor UO_2045 (O_2045,N_29321,N_29708);
xor UO_2046 (O_2046,N_29856,N_29088);
nand UO_2047 (O_2047,N_29198,N_29116);
and UO_2048 (O_2048,N_29956,N_29504);
nand UO_2049 (O_2049,N_28798,N_28735);
xnor UO_2050 (O_2050,N_29136,N_28870);
nand UO_2051 (O_2051,N_28252,N_28535);
nand UO_2052 (O_2052,N_29048,N_28665);
nand UO_2053 (O_2053,N_28868,N_28728);
nand UO_2054 (O_2054,N_29751,N_29302);
nand UO_2055 (O_2055,N_28125,N_29737);
and UO_2056 (O_2056,N_28118,N_28522);
nor UO_2057 (O_2057,N_29993,N_28199);
xor UO_2058 (O_2058,N_29161,N_29107);
xor UO_2059 (O_2059,N_28157,N_29649);
xor UO_2060 (O_2060,N_29595,N_29370);
nor UO_2061 (O_2061,N_29836,N_28332);
xor UO_2062 (O_2062,N_29712,N_29647);
nand UO_2063 (O_2063,N_29326,N_28652);
xnor UO_2064 (O_2064,N_29940,N_29709);
and UO_2065 (O_2065,N_28213,N_28174);
xor UO_2066 (O_2066,N_29588,N_28756);
nor UO_2067 (O_2067,N_28595,N_28174);
xnor UO_2068 (O_2068,N_29272,N_28366);
and UO_2069 (O_2069,N_29350,N_29824);
xor UO_2070 (O_2070,N_28728,N_29691);
nor UO_2071 (O_2071,N_28572,N_29915);
nor UO_2072 (O_2072,N_28376,N_28913);
and UO_2073 (O_2073,N_29983,N_29158);
nor UO_2074 (O_2074,N_29922,N_29233);
nor UO_2075 (O_2075,N_29161,N_28495);
and UO_2076 (O_2076,N_28976,N_29541);
nand UO_2077 (O_2077,N_28942,N_29058);
nand UO_2078 (O_2078,N_28739,N_29032);
nor UO_2079 (O_2079,N_28454,N_29844);
or UO_2080 (O_2080,N_28102,N_29497);
nor UO_2081 (O_2081,N_28414,N_28881);
or UO_2082 (O_2082,N_28186,N_29453);
or UO_2083 (O_2083,N_28818,N_28349);
or UO_2084 (O_2084,N_29550,N_29619);
or UO_2085 (O_2085,N_29899,N_28785);
xor UO_2086 (O_2086,N_28906,N_28090);
nand UO_2087 (O_2087,N_29040,N_28713);
xor UO_2088 (O_2088,N_29610,N_28303);
or UO_2089 (O_2089,N_29283,N_29689);
nand UO_2090 (O_2090,N_29394,N_29043);
xnor UO_2091 (O_2091,N_29261,N_29760);
nor UO_2092 (O_2092,N_29485,N_28364);
or UO_2093 (O_2093,N_28321,N_28249);
and UO_2094 (O_2094,N_29074,N_29680);
xor UO_2095 (O_2095,N_28326,N_28977);
xor UO_2096 (O_2096,N_29415,N_28756);
nor UO_2097 (O_2097,N_29967,N_29521);
nor UO_2098 (O_2098,N_29835,N_29853);
xnor UO_2099 (O_2099,N_29897,N_28521);
nand UO_2100 (O_2100,N_29226,N_28375);
and UO_2101 (O_2101,N_28948,N_29895);
xor UO_2102 (O_2102,N_29359,N_29370);
nor UO_2103 (O_2103,N_28037,N_28085);
nand UO_2104 (O_2104,N_29482,N_29361);
nor UO_2105 (O_2105,N_29805,N_28088);
or UO_2106 (O_2106,N_28036,N_29594);
and UO_2107 (O_2107,N_29987,N_29707);
xor UO_2108 (O_2108,N_28876,N_29824);
or UO_2109 (O_2109,N_29738,N_28294);
nand UO_2110 (O_2110,N_29155,N_29035);
nand UO_2111 (O_2111,N_28828,N_29115);
nand UO_2112 (O_2112,N_28352,N_28140);
or UO_2113 (O_2113,N_29867,N_29161);
nand UO_2114 (O_2114,N_29886,N_28357);
nand UO_2115 (O_2115,N_28692,N_28436);
nand UO_2116 (O_2116,N_28986,N_29030);
and UO_2117 (O_2117,N_28295,N_28227);
and UO_2118 (O_2118,N_29398,N_28271);
xnor UO_2119 (O_2119,N_29215,N_28620);
and UO_2120 (O_2120,N_29528,N_29820);
nor UO_2121 (O_2121,N_29092,N_28395);
or UO_2122 (O_2122,N_28713,N_29452);
or UO_2123 (O_2123,N_29356,N_28437);
nor UO_2124 (O_2124,N_29091,N_28255);
nand UO_2125 (O_2125,N_29962,N_28609);
nand UO_2126 (O_2126,N_29573,N_28801);
and UO_2127 (O_2127,N_28992,N_29633);
or UO_2128 (O_2128,N_29764,N_29644);
and UO_2129 (O_2129,N_29354,N_29257);
and UO_2130 (O_2130,N_29819,N_28118);
xnor UO_2131 (O_2131,N_29946,N_29412);
xnor UO_2132 (O_2132,N_28465,N_29548);
and UO_2133 (O_2133,N_28514,N_28557);
nor UO_2134 (O_2134,N_29039,N_29186);
nor UO_2135 (O_2135,N_28371,N_29006);
xnor UO_2136 (O_2136,N_28899,N_28160);
nor UO_2137 (O_2137,N_28929,N_29467);
or UO_2138 (O_2138,N_29943,N_29371);
nand UO_2139 (O_2139,N_29570,N_28620);
xor UO_2140 (O_2140,N_29249,N_29355);
xor UO_2141 (O_2141,N_28879,N_29060);
nor UO_2142 (O_2142,N_29147,N_29063);
xor UO_2143 (O_2143,N_29502,N_28811);
or UO_2144 (O_2144,N_29230,N_29301);
xor UO_2145 (O_2145,N_28170,N_28439);
or UO_2146 (O_2146,N_28519,N_29756);
xor UO_2147 (O_2147,N_29386,N_28191);
nor UO_2148 (O_2148,N_28666,N_29463);
nand UO_2149 (O_2149,N_28351,N_29169);
and UO_2150 (O_2150,N_29755,N_29261);
xor UO_2151 (O_2151,N_28190,N_29014);
xor UO_2152 (O_2152,N_28236,N_28036);
and UO_2153 (O_2153,N_29074,N_29033);
or UO_2154 (O_2154,N_29103,N_28118);
nor UO_2155 (O_2155,N_28836,N_29325);
and UO_2156 (O_2156,N_29663,N_28115);
nand UO_2157 (O_2157,N_28928,N_29574);
and UO_2158 (O_2158,N_28157,N_28255);
or UO_2159 (O_2159,N_28220,N_28394);
nand UO_2160 (O_2160,N_29538,N_28099);
nor UO_2161 (O_2161,N_29946,N_28203);
nor UO_2162 (O_2162,N_29369,N_29835);
nand UO_2163 (O_2163,N_29979,N_29347);
nand UO_2164 (O_2164,N_28733,N_29843);
or UO_2165 (O_2165,N_29668,N_28982);
nor UO_2166 (O_2166,N_29852,N_29381);
nand UO_2167 (O_2167,N_28264,N_29293);
xor UO_2168 (O_2168,N_28908,N_28065);
or UO_2169 (O_2169,N_29483,N_28342);
or UO_2170 (O_2170,N_29028,N_28646);
nand UO_2171 (O_2171,N_29098,N_29740);
nand UO_2172 (O_2172,N_29106,N_29153);
nor UO_2173 (O_2173,N_29862,N_29944);
and UO_2174 (O_2174,N_28723,N_29565);
nand UO_2175 (O_2175,N_29247,N_29394);
and UO_2176 (O_2176,N_28815,N_29778);
or UO_2177 (O_2177,N_28754,N_29489);
and UO_2178 (O_2178,N_28915,N_29135);
nand UO_2179 (O_2179,N_28647,N_29054);
nor UO_2180 (O_2180,N_28791,N_29699);
nand UO_2181 (O_2181,N_29491,N_28248);
nand UO_2182 (O_2182,N_28457,N_28007);
and UO_2183 (O_2183,N_29032,N_29095);
or UO_2184 (O_2184,N_28685,N_28771);
and UO_2185 (O_2185,N_28588,N_29875);
nand UO_2186 (O_2186,N_28192,N_28916);
nand UO_2187 (O_2187,N_28398,N_28826);
or UO_2188 (O_2188,N_28171,N_29308);
xnor UO_2189 (O_2189,N_29043,N_29685);
xnor UO_2190 (O_2190,N_29245,N_29191);
xnor UO_2191 (O_2191,N_28054,N_29491);
or UO_2192 (O_2192,N_28292,N_28144);
and UO_2193 (O_2193,N_29317,N_28029);
or UO_2194 (O_2194,N_28986,N_28260);
and UO_2195 (O_2195,N_28011,N_28065);
xor UO_2196 (O_2196,N_29409,N_29914);
and UO_2197 (O_2197,N_28478,N_28036);
or UO_2198 (O_2198,N_29754,N_29899);
nor UO_2199 (O_2199,N_29430,N_29833);
or UO_2200 (O_2200,N_29615,N_28626);
nand UO_2201 (O_2201,N_29357,N_29084);
xnor UO_2202 (O_2202,N_29300,N_28096);
and UO_2203 (O_2203,N_29278,N_29573);
or UO_2204 (O_2204,N_28050,N_29763);
and UO_2205 (O_2205,N_28346,N_29498);
or UO_2206 (O_2206,N_28055,N_28942);
and UO_2207 (O_2207,N_29877,N_28459);
and UO_2208 (O_2208,N_28567,N_28839);
and UO_2209 (O_2209,N_29518,N_28879);
nand UO_2210 (O_2210,N_29843,N_29709);
nor UO_2211 (O_2211,N_29941,N_28248);
or UO_2212 (O_2212,N_29462,N_29770);
and UO_2213 (O_2213,N_28535,N_29979);
nand UO_2214 (O_2214,N_29927,N_29119);
and UO_2215 (O_2215,N_29062,N_28634);
and UO_2216 (O_2216,N_29401,N_28626);
xor UO_2217 (O_2217,N_29087,N_28372);
and UO_2218 (O_2218,N_28386,N_29818);
nor UO_2219 (O_2219,N_28275,N_28508);
and UO_2220 (O_2220,N_29967,N_28598);
nor UO_2221 (O_2221,N_29502,N_28742);
nor UO_2222 (O_2222,N_29228,N_29143);
nand UO_2223 (O_2223,N_29886,N_29902);
or UO_2224 (O_2224,N_28072,N_29096);
or UO_2225 (O_2225,N_28470,N_29415);
or UO_2226 (O_2226,N_28019,N_29024);
or UO_2227 (O_2227,N_28573,N_29701);
nand UO_2228 (O_2228,N_28702,N_29805);
nand UO_2229 (O_2229,N_28747,N_28902);
and UO_2230 (O_2230,N_29787,N_29395);
xor UO_2231 (O_2231,N_28000,N_28154);
nand UO_2232 (O_2232,N_29163,N_28721);
or UO_2233 (O_2233,N_28262,N_28844);
xnor UO_2234 (O_2234,N_28489,N_28071);
xor UO_2235 (O_2235,N_28638,N_29610);
or UO_2236 (O_2236,N_29205,N_29695);
xor UO_2237 (O_2237,N_29903,N_29789);
and UO_2238 (O_2238,N_28710,N_28897);
and UO_2239 (O_2239,N_29586,N_29980);
nor UO_2240 (O_2240,N_28010,N_28316);
xnor UO_2241 (O_2241,N_29831,N_28911);
nor UO_2242 (O_2242,N_29816,N_29280);
or UO_2243 (O_2243,N_28670,N_28928);
nor UO_2244 (O_2244,N_28949,N_28037);
nor UO_2245 (O_2245,N_29823,N_29705);
nand UO_2246 (O_2246,N_28056,N_28748);
nor UO_2247 (O_2247,N_29369,N_28737);
and UO_2248 (O_2248,N_29765,N_29093);
nand UO_2249 (O_2249,N_28874,N_28036);
nor UO_2250 (O_2250,N_29695,N_28304);
and UO_2251 (O_2251,N_29707,N_29877);
nand UO_2252 (O_2252,N_28338,N_29886);
and UO_2253 (O_2253,N_29825,N_28647);
or UO_2254 (O_2254,N_29658,N_28294);
or UO_2255 (O_2255,N_29773,N_29822);
and UO_2256 (O_2256,N_28970,N_28993);
nor UO_2257 (O_2257,N_29452,N_29790);
nor UO_2258 (O_2258,N_29878,N_28112);
nor UO_2259 (O_2259,N_29601,N_28223);
nand UO_2260 (O_2260,N_28786,N_28140);
xor UO_2261 (O_2261,N_28684,N_29710);
or UO_2262 (O_2262,N_29282,N_29687);
nor UO_2263 (O_2263,N_29576,N_29932);
nand UO_2264 (O_2264,N_29272,N_29725);
nand UO_2265 (O_2265,N_28563,N_29203);
and UO_2266 (O_2266,N_29808,N_29464);
nand UO_2267 (O_2267,N_28204,N_29294);
and UO_2268 (O_2268,N_28394,N_28640);
or UO_2269 (O_2269,N_29531,N_29841);
nand UO_2270 (O_2270,N_28194,N_28607);
nor UO_2271 (O_2271,N_29586,N_29081);
xnor UO_2272 (O_2272,N_29888,N_29912);
or UO_2273 (O_2273,N_29868,N_28043);
xnor UO_2274 (O_2274,N_28589,N_29044);
or UO_2275 (O_2275,N_28421,N_28834);
xnor UO_2276 (O_2276,N_28618,N_28443);
nand UO_2277 (O_2277,N_28606,N_28642);
nand UO_2278 (O_2278,N_28517,N_28262);
xnor UO_2279 (O_2279,N_29345,N_29053);
and UO_2280 (O_2280,N_29037,N_28009);
or UO_2281 (O_2281,N_29576,N_29551);
or UO_2282 (O_2282,N_28267,N_29894);
or UO_2283 (O_2283,N_29280,N_28575);
nand UO_2284 (O_2284,N_29169,N_29958);
nor UO_2285 (O_2285,N_28542,N_29553);
nand UO_2286 (O_2286,N_29389,N_29315);
or UO_2287 (O_2287,N_28661,N_29254);
nand UO_2288 (O_2288,N_28335,N_29778);
and UO_2289 (O_2289,N_29779,N_29103);
nand UO_2290 (O_2290,N_29503,N_29717);
nor UO_2291 (O_2291,N_29218,N_29472);
or UO_2292 (O_2292,N_28372,N_29366);
or UO_2293 (O_2293,N_29377,N_28607);
and UO_2294 (O_2294,N_29477,N_29455);
or UO_2295 (O_2295,N_29487,N_28683);
nand UO_2296 (O_2296,N_29856,N_29049);
nor UO_2297 (O_2297,N_28671,N_29430);
and UO_2298 (O_2298,N_28251,N_29968);
nand UO_2299 (O_2299,N_29867,N_28229);
or UO_2300 (O_2300,N_28987,N_29133);
xnor UO_2301 (O_2301,N_29880,N_29141);
xnor UO_2302 (O_2302,N_29333,N_29300);
or UO_2303 (O_2303,N_28921,N_28771);
nand UO_2304 (O_2304,N_29774,N_28371);
or UO_2305 (O_2305,N_29325,N_29374);
or UO_2306 (O_2306,N_29462,N_28783);
xor UO_2307 (O_2307,N_28482,N_29946);
nor UO_2308 (O_2308,N_28600,N_28717);
xnor UO_2309 (O_2309,N_28905,N_29503);
xor UO_2310 (O_2310,N_29736,N_28414);
nand UO_2311 (O_2311,N_29940,N_28847);
nor UO_2312 (O_2312,N_29752,N_29765);
nand UO_2313 (O_2313,N_28053,N_28417);
or UO_2314 (O_2314,N_28243,N_28170);
xnor UO_2315 (O_2315,N_28900,N_28215);
or UO_2316 (O_2316,N_29945,N_28469);
or UO_2317 (O_2317,N_29437,N_29308);
and UO_2318 (O_2318,N_29799,N_28195);
and UO_2319 (O_2319,N_29201,N_29507);
and UO_2320 (O_2320,N_29602,N_28825);
nand UO_2321 (O_2321,N_29546,N_28067);
nor UO_2322 (O_2322,N_29271,N_28895);
nand UO_2323 (O_2323,N_28943,N_28659);
or UO_2324 (O_2324,N_29466,N_29262);
nand UO_2325 (O_2325,N_28320,N_28160);
nand UO_2326 (O_2326,N_29384,N_28225);
or UO_2327 (O_2327,N_29131,N_28658);
xnor UO_2328 (O_2328,N_29908,N_29399);
nor UO_2329 (O_2329,N_29045,N_28728);
nor UO_2330 (O_2330,N_28541,N_29911);
or UO_2331 (O_2331,N_28012,N_29123);
xnor UO_2332 (O_2332,N_29208,N_28833);
nand UO_2333 (O_2333,N_28534,N_28796);
or UO_2334 (O_2334,N_28213,N_29012);
nand UO_2335 (O_2335,N_29775,N_29448);
xnor UO_2336 (O_2336,N_28465,N_29417);
nor UO_2337 (O_2337,N_28164,N_28716);
and UO_2338 (O_2338,N_28319,N_29047);
xor UO_2339 (O_2339,N_29653,N_29666);
nor UO_2340 (O_2340,N_29962,N_29704);
xnor UO_2341 (O_2341,N_28586,N_29987);
or UO_2342 (O_2342,N_29289,N_28804);
xor UO_2343 (O_2343,N_29151,N_28829);
nor UO_2344 (O_2344,N_28266,N_29342);
and UO_2345 (O_2345,N_28112,N_28051);
nand UO_2346 (O_2346,N_28228,N_28396);
nand UO_2347 (O_2347,N_29453,N_29446);
or UO_2348 (O_2348,N_29260,N_28492);
nand UO_2349 (O_2349,N_29808,N_29638);
nor UO_2350 (O_2350,N_28473,N_28802);
xnor UO_2351 (O_2351,N_28413,N_28720);
nand UO_2352 (O_2352,N_28400,N_29665);
xor UO_2353 (O_2353,N_28333,N_29037);
nor UO_2354 (O_2354,N_29640,N_28876);
nand UO_2355 (O_2355,N_29691,N_28029);
nor UO_2356 (O_2356,N_29369,N_29675);
or UO_2357 (O_2357,N_28626,N_29383);
and UO_2358 (O_2358,N_28816,N_29082);
xor UO_2359 (O_2359,N_29537,N_29866);
nand UO_2360 (O_2360,N_28737,N_29812);
xnor UO_2361 (O_2361,N_28424,N_28979);
nor UO_2362 (O_2362,N_28936,N_29547);
xor UO_2363 (O_2363,N_29168,N_28014);
xor UO_2364 (O_2364,N_29834,N_29135);
or UO_2365 (O_2365,N_28573,N_29975);
nand UO_2366 (O_2366,N_28563,N_28595);
nor UO_2367 (O_2367,N_29302,N_29715);
nand UO_2368 (O_2368,N_28731,N_28927);
nand UO_2369 (O_2369,N_29662,N_28603);
and UO_2370 (O_2370,N_29502,N_28129);
or UO_2371 (O_2371,N_29054,N_29403);
xnor UO_2372 (O_2372,N_28320,N_29753);
xnor UO_2373 (O_2373,N_28716,N_28125);
and UO_2374 (O_2374,N_29702,N_29200);
nand UO_2375 (O_2375,N_29251,N_28566);
or UO_2376 (O_2376,N_29736,N_29546);
and UO_2377 (O_2377,N_29810,N_28944);
xnor UO_2378 (O_2378,N_29142,N_29150);
nor UO_2379 (O_2379,N_28551,N_28715);
xor UO_2380 (O_2380,N_29651,N_28963);
xor UO_2381 (O_2381,N_28126,N_28429);
nand UO_2382 (O_2382,N_29474,N_28448);
nor UO_2383 (O_2383,N_29803,N_28119);
and UO_2384 (O_2384,N_28080,N_29296);
or UO_2385 (O_2385,N_29214,N_29972);
nand UO_2386 (O_2386,N_28157,N_28921);
nor UO_2387 (O_2387,N_29586,N_29862);
or UO_2388 (O_2388,N_29802,N_28253);
nand UO_2389 (O_2389,N_28724,N_29453);
and UO_2390 (O_2390,N_29719,N_28293);
and UO_2391 (O_2391,N_28192,N_29308);
nand UO_2392 (O_2392,N_28014,N_28646);
or UO_2393 (O_2393,N_29370,N_29133);
nor UO_2394 (O_2394,N_28761,N_28339);
xnor UO_2395 (O_2395,N_28396,N_29092);
nand UO_2396 (O_2396,N_29369,N_29770);
nor UO_2397 (O_2397,N_29997,N_28244);
nand UO_2398 (O_2398,N_28298,N_28733);
nor UO_2399 (O_2399,N_28068,N_28353);
or UO_2400 (O_2400,N_29465,N_29521);
xnor UO_2401 (O_2401,N_28895,N_29867);
nor UO_2402 (O_2402,N_29392,N_29927);
or UO_2403 (O_2403,N_29788,N_29918);
nor UO_2404 (O_2404,N_29513,N_29026);
nand UO_2405 (O_2405,N_29395,N_29589);
and UO_2406 (O_2406,N_28887,N_29365);
nand UO_2407 (O_2407,N_29730,N_28081);
nand UO_2408 (O_2408,N_29953,N_28126);
xnor UO_2409 (O_2409,N_29063,N_29072);
or UO_2410 (O_2410,N_29675,N_28808);
nor UO_2411 (O_2411,N_29328,N_29933);
and UO_2412 (O_2412,N_29815,N_28779);
or UO_2413 (O_2413,N_28020,N_28997);
or UO_2414 (O_2414,N_29008,N_29595);
nor UO_2415 (O_2415,N_29863,N_28034);
and UO_2416 (O_2416,N_29811,N_28930);
or UO_2417 (O_2417,N_28866,N_28366);
and UO_2418 (O_2418,N_28778,N_29002);
or UO_2419 (O_2419,N_28776,N_28658);
xor UO_2420 (O_2420,N_29760,N_29240);
or UO_2421 (O_2421,N_28908,N_28474);
nand UO_2422 (O_2422,N_29661,N_28775);
xor UO_2423 (O_2423,N_29882,N_29271);
xnor UO_2424 (O_2424,N_29889,N_28981);
nand UO_2425 (O_2425,N_29015,N_29646);
nor UO_2426 (O_2426,N_28446,N_28306);
or UO_2427 (O_2427,N_29510,N_29524);
nand UO_2428 (O_2428,N_28296,N_28541);
xor UO_2429 (O_2429,N_29775,N_28406);
or UO_2430 (O_2430,N_28396,N_28628);
or UO_2431 (O_2431,N_29318,N_29577);
nor UO_2432 (O_2432,N_29719,N_28741);
nand UO_2433 (O_2433,N_29351,N_29687);
nand UO_2434 (O_2434,N_28131,N_29936);
nand UO_2435 (O_2435,N_28434,N_29157);
and UO_2436 (O_2436,N_28808,N_28327);
nor UO_2437 (O_2437,N_28458,N_29644);
and UO_2438 (O_2438,N_28270,N_29722);
xor UO_2439 (O_2439,N_29014,N_29303);
xor UO_2440 (O_2440,N_28046,N_29124);
and UO_2441 (O_2441,N_29919,N_29140);
nor UO_2442 (O_2442,N_28462,N_29333);
nand UO_2443 (O_2443,N_28679,N_28200);
nor UO_2444 (O_2444,N_29798,N_29954);
nand UO_2445 (O_2445,N_28517,N_28806);
xnor UO_2446 (O_2446,N_29089,N_28092);
nand UO_2447 (O_2447,N_28978,N_28909);
xnor UO_2448 (O_2448,N_28198,N_29469);
xor UO_2449 (O_2449,N_29807,N_28961);
nand UO_2450 (O_2450,N_28135,N_28779);
and UO_2451 (O_2451,N_29674,N_28155);
and UO_2452 (O_2452,N_28218,N_28007);
and UO_2453 (O_2453,N_28434,N_28350);
nand UO_2454 (O_2454,N_28741,N_28690);
or UO_2455 (O_2455,N_28603,N_29417);
or UO_2456 (O_2456,N_28762,N_28639);
nand UO_2457 (O_2457,N_29541,N_29085);
or UO_2458 (O_2458,N_29278,N_28245);
nor UO_2459 (O_2459,N_29319,N_28070);
nor UO_2460 (O_2460,N_28095,N_28716);
xnor UO_2461 (O_2461,N_29450,N_29308);
xor UO_2462 (O_2462,N_28902,N_28665);
nand UO_2463 (O_2463,N_28025,N_29287);
xnor UO_2464 (O_2464,N_28072,N_29266);
nand UO_2465 (O_2465,N_29359,N_29952);
nand UO_2466 (O_2466,N_29871,N_28440);
nor UO_2467 (O_2467,N_29975,N_28553);
and UO_2468 (O_2468,N_29283,N_28600);
xor UO_2469 (O_2469,N_29385,N_28027);
nand UO_2470 (O_2470,N_29582,N_28889);
or UO_2471 (O_2471,N_28164,N_29135);
nor UO_2472 (O_2472,N_29847,N_28101);
xor UO_2473 (O_2473,N_29547,N_28242);
nand UO_2474 (O_2474,N_28430,N_29018);
xor UO_2475 (O_2475,N_28794,N_28319);
nand UO_2476 (O_2476,N_29098,N_29997);
and UO_2477 (O_2477,N_28015,N_29097);
nand UO_2478 (O_2478,N_28165,N_28313);
xor UO_2479 (O_2479,N_28699,N_28226);
nand UO_2480 (O_2480,N_28226,N_29418);
or UO_2481 (O_2481,N_29914,N_29461);
nor UO_2482 (O_2482,N_28957,N_28675);
and UO_2483 (O_2483,N_28429,N_29353);
or UO_2484 (O_2484,N_28522,N_29542);
or UO_2485 (O_2485,N_28108,N_29219);
xor UO_2486 (O_2486,N_28517,N_29429);
and UO_2487 (O_2487,N_28376,N_28042);
and UO_2488 (O_2488,N_28102,N_29056);
and UO_2489 (O_2489,N_29558,N_28781);
nor UO_2490 (O_2490,N_28057,N_29118);
nand UO_2491 (O_2491,N_28497,N_28992);
nand UO_2492 (O_2492,N_28743,N_29765);
nor UO_2493 (O_2493,N_29252,N_28474);
nor UO_2494 (O_2494,N_29999,N_29722);
and UO_2495 (O_2495,N_28483,N_29252);
and UO_2496 (O_2496,N_28912,N_29856);
or UO_2497 (O_2497,N_29395,N_29763);
nor UO_2498 (O_2498,N_28364,N_28947);
nor UO_2499 (O_2499,N_29011,N_29133);
nand UO_2500 (O_2500,N_28906,N_28577);
xor UO_2501 (O_2501,N_29171,N_28323);
and UO_2502 (O_2502,N_29210,N_28477);
xnor UO_2503 (O_2503,N_28479,N_29159);
xor UO_2504 (O_2504,N_28447,N_28760);
nor UO_2505 (O_2505,N_28713,N_29236);
nor UO_2506 (O_2506,N_28686,N_29693);
nand UO_2507 (O_2507,N_29187,N_28270);
xor UO_2508 (O_2508,N_28235,N_28894);
xor UO_2509 (O_2509,N_29915,N_28063);
or UO_2510 (O_2510,N_28414,N_29505);
nand UO_2511 (O_2511,N_29627,N_29301);
or UO_2512 (O_2512,N_29917,N_29415);
nand UO_2513 (O_2513,N_28693,N_28438);
and UO_2514 (O_2514,N_28657,N_28075);
nor UO_2515 (O_2515,N_29296,N_28284);
nand UO_2516 (O_2516,N_28555,N_28568);
nor UO_2517 (O_2517,N_28549,N_29014);
or UO_2518 (O_2518,N_29769,N_29105);
or UO_2519 (O_2519,N_29092,N_29231);
or UO_2520 (O_2520,N_28871,N_29951);
or UO_2521 (O_2521,N_29271,N_29769);
xnor UO_2522 (O_2522,N_28445,N_29209);
xor UO_2523 (O_2523,N_28291,N_28101);
and UO_2524 (O_2524,N_28506,N_29294);
xor UO_2525 (O_2525,N_28098,N_28396);
nor UO_2526 (O_2526,N_28039,N_28941);
nand UO_2527 (O_2527,N_28587,N_29060);
and UO_2528 (O_2528,N_28372,N_29878);
xor UO_2529 (O_2529,N_28380,N_29193);
nor UO_2530 (O_2530,N_28861,N_28780);
xor UO_2531 (O_2531,N_28784,N_28448);
and UO_2532 (O_2532,N_29352,N_29659);
and UO_2533 (O_2533,N_29945,N_29604);
or UO_2534 (O_2534,N_29986,N_29633);
or UO_2535 (O_2535,N_29041,N_29944);
or UO_2536 (O_2536,N_29700,N_29761);
nor UO_2537 (O_2537,N_28322,N_28408);
xnor UO_2538 (O_2538,N_28330,N_28288);
xnor UO_2539 (O_2539,N_29813,N_29620);
xnor UO_2540 (O_2540,N_29902,N_29906);
nand UO_2541 (O_2541,N_28367,N_29582);
or UO_2542 (O_2542,N_29963,N_28491);
nand UO_2543 (O_2543,N_28484,N_28865);
nand UO_2544 (O_2544,N_29141,N_28695);
nor UO_2545 (O_2545,N_29905,N_28405);
or UO_2546 (O_2546,N_29144,N_28335);
and UO_2547 (O_2547,N_29329,N_29308);
and UO_2548 (O_2548,N_28694,N_28792);
and UO_2549 (O_2549,N_28775,N_29395);
nand UO_2550 (O_2550,N_28422,N_28530);
and UO_2551 (O_2551,N_29690,N_28272);
and UO_2552 (O_2552,N_29923,N_28085);
and UO_2553 (O_2553,N_28621,N_29541);
or UO_2554 (O_2554,N_29043,N_29477);
xor UO_2555 (O_2555,N_29689,N_29355);
or UO_2556 (O_2556,N_29146,N_29712);
and UO_2557 (O_2557,N_29919,N_28357);
xnor UO_2558 (O_2558,N_28647,N_29254);
or UO_2559 (O_2559,N_28143,N_29508);
and UO_2560 (O_2560,N_29527,N_28208);
nand UO_2561 (O_2561,N_29703,N_28171);
nand UO_2562 (O_2562,N_29893,N_29523);
nand UO_2563 (O_2563,N_28407,N_28966);
nand UO_2564 (O_2564,N_28134,N_29523);
or UO_2565 (O_2565,N_29057,N_28385);
and UO_2566 (O_2566,N_29363,N_29394);
nand UO_2567 (O_2567,N_28740,N_29465);
and UO_2568 (O_2568,N_29070,N_29165);
nor UO_2569 (O_2569,N_29036,N_28767);
nand UO_2570 (O_2570,N_28062,N_29563);
and UO_2571 (O_2571,N_29501,N_28721);
xor UO_2572 (O_2572,N_28350,N_29013);
nand UO_2573 (O_2573,N_28998,N_28873);
nor UO_2574 (O_2574,N_28552,N_29055);
xor UO_2575 (O_2575,N_28725,N_28580);
or UO_2576 (O_2576,N_29359,N_28199);
and UO_2577 (O_2577,N_29202,N_29379);
nand UO_2578 (O_2578,N_28371,N_28028);
or UO_2579 (O_2579,N_28288,N_28692);
nor UO_2580 (O_2580,N_29595,N_29131);
or UO_2581 (O_2581,N_29025,N_29034);
or UO_2582 (O_2582,N_29662,N_28417);
or UO_2583 (O_2583,N_29420,N_29932);
xnor UO_2584 (O_2584,N_28073,N_28071);
and UO_2585 (O_2585,N_29688,N_28505);
and UO_2586 (O_2586,N_29173,N_29677);
or UO_2587 (O_2587,N_29216,N_28609);
xnor UO_2588 (O_2588,N_29431,N_28308);
nand UO_2589 (O_2589,N_28728,N_29675);
nand UO_2590 (O_2590,N_29899,N_28230);
or UO_2591 (O_2591,N_29373,N_28816);
nand UO_2592 (O_2592,N_28861,N_28516);
xnor UO_2593 (O_2593,N_29356,N_28707);
and UO_2594 (O_2594,N_28692,N_29592);
xnor UO_2595 (O_2595,N_29691,N_28267);
nor UO_2596 (O_2596,N_28572,N_29183);
nand UO_2597 (O_2597,N_29221,N_29424);
nor UO_2598 (O_2598,N_29394,N_28975);
and UO_2599 (O_2599,N_29053,N_28445);
and UO_2600 (O_2600,N_29365,N_28461);
xor UO_2601 (O_2601,N_29680,N_28878);
nor UO_2602 (O_2602,N_28564,N_29242);
or UO_2603 (O_2603,N_28403,N_29579);
and UO_2604 (O_2604,N_29913,N_28398);
nor UO_2605 (O_2605,N_29111,N_28967);
nand UO_2606 (O_2606,N_29765,N_29277);
xor UO_2607 (O_2607,N_28995,N_28749);
nor UO_2608 (O_2608,N_28392,N_28100);
and UO_2609 (O_2609,N_28095,N_28785);
nand UO_2610 (O_2610,N_29791,N_28400);
xor UO_2611 (O_2611,N_28499,N_28434);
and UO_2612 (O_2612,N_28342,N_29979);
and UO_2613 (O_2613,N_29325,N_28650);
nor UO_2614 (O_2614,N_28655,N_28141);
xor UO_2615 (O_2615,N_29206,N_29986);
and UO_2616 (O_2616,N_28293,N_28272);
and UO_2617 (O_2617,N_28413,N_29464);
nor UO_2618 (O_2618,N_29016,N_29195);
nand UO_2619 (O_2619,N_29857,N_29945);
nor UO_2620 (O_2620,N_29622,N_28985);
and UO_2621 (O_2621,N_28706,N_29983);
or UO_2622 (O_2622,N_29186,N_29300);
nor UO_2623 (O_2623,N_29480,N_29618);
nand UO_2624 (O_2624,N_28158,N_28047);
and UO_2625 (O_2625,N_29649,N_28819);
nor UO_2626 (O_2626,N_29846,N_29824);
and UO_2627 (O_2627,N_29043,N_28564);
or UO_2628 (O_2628,N_28998,N_28225);
nand UO_2629 (O_2629,N_28987,N_28123);
nor UO_2630 (O_2630,N_28411,N_28095);
nand UO_2631 (O_2631,N_28350,N_28426);
xor UO_2632 (O_2632,N_29027,N_28559);
and UO_2633 (O_2633,N_28876,N_28753);
nand UO_2634 (O_2634,N_28914,N_28491);
or UO_2635 (O_2635,N_28394,N_28100);
or UO_2636 (O_2636,N_28184,N_29035);
xor UO_2637 (O_2637,N_29931,N_28367);
or UO_2638 (O_2638,N_29340,N_28105);
nor UO_2639 (O_2639,N_28198,N_28254);
nand UO_2640 (O_2640,N_28835,N_29889);
nand UO_2641 (O_2641,N_28828,N_29566);
nand UO_2642 (O_2642,N_29408,N_28187);
nand UO_2643 (O_2643,N_28668,N_28888);
nand UO_2644 (O_2644,N_28487,N_28821);
nand UO_2645 (O_2645,N_29946,N_28443);
and UO_2646 (O_2646,N_29783,N_28759);
xor UO_2647 (O_2647,N_28543,N_28386);
and UO_2648 (O_2648,N_29829,N_29865);
nand UO_2649 (O_2649,N_29876,N_28157);
xnor UO_2650 (O_2650,N_29064,N_29267);
or UO_2651 (O_2651,N_29622,N_29757);
and UO_2652 (O_2652,N_28828,N_29716);
nand UO_2653 (O_2653,N_29057,N_29255);
xor UO_2654 (O_2654,N_28664,N_28015);
and UO_2655 (O_2655,N_29532,N_29974);
or UO_2656 (O_2656,N_29564,N_29710);
nand UO_2657 (O_2657,N_28067,N_29883);
and UO_2658 (O_2658,N_29683,N_29836);
nand UO_2659 (O_2659,N_28897,N_28362);
and UO_2660 (O_2660,N_29416,N_29993);
nand UO_2661 (O_2661,N_28960,N_29390);
nor UO_2662 (O_2662,N_29193,N_29239);
nand UO_2663 (O_2663,N_29359,N_29698);
nor UO_2664 (O_2664,N_29921,N_28467);
nor UO_2665 (O_2665,N_28721,N_29283);
xor UO_2666 (O_2666,N_28206,N_29076);
nand UO_2667 (O_2667,N_28418,N_29220);
and UO_2668 (O_2668,N_29337,N_28852);
xor UO_2669 (O_2669,N_29069,N_28580);
nand UO_2670 (O_2670,N_28100,N_28233);
or UO_2671 (O_2671,N_29445,N_28441);
or UO_2672 (O_2672,N_28860,N_28098);
xnor UO_2673 (O_2673,N_29247,N_28720);
nand UO_2674 (O_2674,N_28707,N_29712);
nor UO_2675 (O_2675,N_28972,N_29584);
nand UO_2676 (O_2676,N_28882,N_28162);
xnor UO_2677 (O_2677,N_28423,N_28276);
nand UO_2678 (O_2678,N_29566,N_28358);
xnor UO_2679 (O_2679,N_29484,N_28225);
or UO_2680 (O_2680,N_28072,N_28975);
nand UO_2681 (O_2681,N_29668,N_28362);
nor UO_2682 (O_2682,N_28260,N_29824);
or UO_2683 (O_2683,N_28591,N_29885);
xnor UO_2684 (O_2684,N_28287,N_29035);
xor UO_2685 (O_2685,N_29319,N_29811);
nand UO_2686 (O_2686,N_28902,N_28304);
nor UO_2687 (O_2687,N_28143,N_29452);
or UO_2688 (O_2688,N_29457,N_29565);
and UO_2689 (O_2689,N_29382,N_28298);
or UO_2690 (O_2690,N_28592,N_29598);
or UO_2691 (O_2691,N_28270,N_28672);
nor UO_2692 (O_2692,N_29461,N_29759);
nand UO_2693 (O_2693,N_29170,N_29159);
nor UO_2694 (O_2694,N_28782,N_28126);
nand UO_2695 (O_2695,N_29734,N_28386);
nor UO_2696 (O_2696,N_29139,N_29721);
nand UO_2697 (O_2697,N_28126,N_29744);
nor UO_2698 (O_2698,N_28560,N_28898);
and UO_2699 (O_2699,N_28545,N_29031);
xnor UO_2700 (O_2700,N_29171,N_28194);
or UO_2701 (O_2701,N_29675,N_29122);
or UO_2702 (O_2702,N_29909,N_29640);
or UO_2703 (O_2703,N_28312,N_28308);
nor UO_2704 (O_2704,N_29713,N_28452);
nand UO_2705 (O_2705,N_29821,N_28922);
xnor UO_2706 (O_2706,N_28727,N_28504);
xor UO_2707 (O_2707,N_28492,N_28763);
or UO_2708 (O_2708,N_29032,N_29356);
nand UO_2709 (O_2709,N_29282,N_28340);
xor UO_2710 (O_2710,N_29881,N_28462);
nor UO_2711 (O_2711,N_28618,N_29873);
xor UO_2712 (O_2712,N_29770,N_29329);
nand UO_2713 (O_2713,N_29784,N_28019);
or UO_2714 (O_2714,N_28767,N_29476);
nor UO_2715 (O_2715,N_28647,N_29844);
xor UO_2716 (O_2716,N_28693,N_28900);
xnor UO_2717 (O_2717,N_28965,N_28861);
or UO_2718 (O_2718,N_29104,N_29772);
xor UO_2719 (O_2719,N_29472,N_29254);
nand UO_2720 (O_2720,N_29264,N_28057);
or UO_2721 (O_2721,N_29158,N_28793);
or UO_2722 (O_2722,N_29316,N_28670);
xor UO_2723 (O_2723,N_29001,N_29461);
nand UO_2724 (O_2724,N_29061,N_28456);
nor UO_2725 (O_2725,N_29730,N_29414);
and UO_2726 (O_2726,N_29518,N_28195);
nand UO_2727 (O_2727,N_29882,N_29926);
and UO_2728 (O_2728,N_28967,N_29145);
xnor UO_2729 (O_2729,N_28464,N_29552);
or UO_2730 (O_2730,N_28327,N_28446);
xnor UO_2731 (O_2731,N_29389,N_28659);
nand UO_2732 (O_2732,N_28372,N_28896);
nor UO_2733 (O_2733,N_28594,N_28784);
xnor UO_2734 (O_2734,N_29796,N_28145);
xor UO_2735 (O_2735,N_28247,N_29047);
xnor UO_2736 (O_2736,N_28514,N_29988);
nor UO_2737 (O_2737,N_29245,N_29163);
xnor UO_2738 (O_2738,N_28936,N_29158);
nand UO_2739 (O_2739,N_29194,N_28193);
or UO_2740 (O_2740,N_28088,N_28010);
nor UO_2741 (O_2741,N_29451,N_28761);
nand UO_2742 (O_2742,N_29272,N_28114);
nand UO_2743 (O_2743,N_28682,N_28309);
xor UO_2744 (O_2744,N_29887,N_29671);
or UO_2745 (O_2745,N_29489,N_29947);
nand UO_2746 (O_2746,N_29756,N_29912);
nor UO_2747 (O_2747,N_28721,N_28545);
nand UO_2748 (O_2748,N_29175,N_29142);
xnor UO_2749 (O_2749,N_29333,N_28000);
xor UO_2750 (O_2750,N_28456,N_29923);
xor UO_2751 (O_2751,N_28668,N_29563);
and UO_2752 (O_2752,N_29354,N_28528);
nor UO_2753 (O_2753,N_29136,N_28920);
or UO_2754 (O_2754,N_29909,N_29262);
or UO_2755 (O_2755,N_28053,N_29425);
xnor UO_2756 (O_2756,N_28903,N_29853);
and UO_2757 (O_2757,N_29938,N_28544);
and UO_2758 (O_2758,N_29000,N_29028);
xnor UO_2759 (O_2759,N_29736,N_28228);
and UO_2760 (O_2760,N_28669,N_28312);
nor UO_2761 (O_2761,N_29586,N_28003);
nand UO_2762 (O_2762,N_28113,N_28120);
xor UO_2763 (O_2763,N_28978,N_28533);
or UO_2764 (O_2764,N_28765,N_29402);
and UO_2765 (O_2765,N_29913,N_29314);
and UO_2766 (O_2766,N_29519,N_29984);
and UO_2767 (O_2767,N_28956,N_29480);
nor UO_2768 (O_2768,N_29318,N_28096);
or UO_2769 (O_2769,N_28664,N_29789);
nor UO_2770 (O_2770,N_28497,N_28176);
and UO_2771 (O_2771,N_29417,N_28268);
xnor UO_2772 (O_2772,N_28593,N_29301);
nor UO_2773 (O_2773,N_28495,N_29890);
nor UO_2774 (O_2774,N_29600,N_28382);
and UO_2775 (O_2775,N_29390,N_28643);
xor UO_2776 (O_2776,N_28729,N_29365);
nand UO_2777 (O_2777,N_28634,N_29747);
or UO_2778 (O_2778,N_29496,N_28968);
nand UO_2779 (O_2779,N_28090,N_28958);
or UO_2780 (O_2780,N_29775,N_28753);
and UO_2781 (O_2781,N_29972,N_29344);
nor UO_2782 (O_2782,N_28474,N_28911);
and UO_2783 (O_2783,N_29839,N_28037);
and UO_2784 (O_2784,N_28717,N_29801);
nor UO_2785 (O_2785,N_29690,N_29408);
or UO_2786 (O_2786,N_29082,N_29923);
or UO_2787 (O_2787,N_28165,N_29674);
nand UO_2788 (O_2788,N_29208,N_28331);
or UO_2789 (O_2789,N_28561,N_29001);
and UO_2790 (O_2790,N_29747,N_28580);
or UO_2791 (O_2791,N_29652,N_29477);
and UO_2792 (O_2792,N_28161,N_28636);
nor UO_2793 (O_2793,N_29277,N_28905);
xor UO_2794 (O_2794,N_29017,N_29388);
or UO_2795 (O_2795,N_28444,N_29456);
xnor UO_2796 (O_2796,N_29038,N_29120);
and UO_2797 (O_2797,N_28146,N_29854);
nor UO_2798 (O_2798,N_28512,N_28665);
xnor UO_2799 (O_2799,N_28278,N_29469);
nor UO_2800 (O_2800,N_28186,N_29880);
nand UO_2801 (O_2801,N_28686,N_28886);
nor UO_2802 (O_2802,N_28287,N_28878);
xor UO_2803 (O_2803,N_28673,N_28369);
or UO_2804 (O_2804,N_29708,N_28899);
nand UO_2805 (O_2805,N_29520,N_28463);
nor UO_2806 (O_2806,N_29163,N_29125);
and UO_2807 (O_2807,N_29362,N_28681);
xor UO_2808 (O_2808,N_29900,N_29098);
nor UO_2809 (O_2809,N_29883,N_29800);
xor UO_2810 (O_2810,N_28425,N_29089);
and UO_2811 (O_2811,N_29701,N_28726);
nand UO_2812 (O_2812,N_28468,N_29182);
nor UO_2813 (O_2813,N_28946,N_28048);
nand UO_2814 (O_2814,N_29664,N_29621);
or UO_2815 (O_2815,N_28028,N_28421);
xnor UO_2816 (O_2816,N_28408,N_29647);
or UO_2817 (O_2817,N_29128,N_28506);
and UO_2818 (O_2818,N_28250,N_29190);
or UO_2819 (O_2819,N_28619,N_29490);
and UO_2820 (O_2820,N_28930,N_29707);
or UO_2821 (O_2821,N_28438,N_28478);
or UO_2822 (O_2822,N_29076,N_29294);
nor UO_2823 (O_2823,N_29006,N_28052);
or UO_2824 (O_2824,N_28312,N_29596);
nand UO_2825 (O_2825,N_28767,N_29532);
nor UO_2826 (O_2826,N_28589,N_28236);
or UO_2827 (O_2827,N_29560,N_29734);
and UO_2828 (O_2828,N_29887,N_29103);
or UO_2829 (O_2829,N_28031,N_28814);
nand UO_2830 (O_2830,N_29429,N_28694);
nor UO_2831 (O_2831,N_28626,N_29203);
nor UO_2832 (O_2832,N_29060,N_29600);
and UO_2833 (O_2833,N_28520,N_28586);
xor UO_2834 (O_2834,N_28265,N_29173);
or UO_2835 (O_2835,N_28346,N_28843);
nand UO_2836 (O_2836,N_29614,N_29738);
or UO_2837 (O_2837,N_28294,N_28324);
xnor UO_2838 (O_2838,N_29877,N_28482);
and UO_2839 (O_2839,N_28574,N_28196);
xnor UO_2840 (O_2840,N_29764,N_28329);
nand UO_2841 (O_2841,N_29113,N_28296);
and UO_2842 (O_2842,N_28433,N_28243);
nor UO_2843 (O_2843,N_29455,N_28215);
nor UO_2844 (O_2844,N_28280,N_29636);
xor UO_2845 (O_2845,N_29321,N_28395);
nor UO_2846 (O_2846,N_29481,N_29881);
nand UO_2847 (O_2847,N_28876,N_29427);
nor UO_2848 (O_2848,N_29572,N_29638);
and UO_2849 (O_2849,N_28882,N_28442);
nor UO_2850 (O_2850,N_29820,N_28401);
and UO_2851 (O_2851,N_28851,N_29122);
or UO_2852 (O_2852,N_29086,N_28042);
or UO_2853 (O_2853,N_28229,N_28899);
and UO_2854 (O_2854,N_28686,N_28248);
nand UO_2855 (O_2855,N_28904,N_29048);
nor UO_2856 (O_2856,N_29584,N_28463);
or UO_2857 (O_2857,N_28995,N_28999);
nand UO_2858 (O_2858,N_29755,N_29655);
or UO_2859 (O_2859,N_29888,N_28791);
xnor UO_2860 (O_2860,N_29350,N_28222);
and UO_2861 (O_2861,N_28580,N_29039);
xor UO_2862 (O_2862,N_28235,N_29225);
and UO_2863 (O_2863,N_28973,N_29846);
xor UO_2864 (O_2864,N_28444,N_28535);
xnor UO_2865 (O_2865,N_29008,N_29647);
or UO_2866 (O_2866,N_29415,N_29584);
xnor UO_2867 (O_2867,N_29070,N_29167);
nand UO_2868 (O_2868,N_29017,N_29649);
and UO_2869 (O_2869,N_28722,N_28259);
or UO_2870 (O_2870,N_28318,N_28003);
or UO_2871 (O_2871,N_29787,N_28731);
and UO_2872 (O_2872,N_29895,N_28754);
or UO_2873 (O_2873,N_29182,N_29210);
or UO_2874 (O_2874,N_29236,N_28082);
or UO_2875 (O_2875,N_28773,N_29267);
nand UO_2876 (O_2876,N_28495,N_28889);
xor UO_2877 (O_2877,N_28801,N_28072);
or UO_2878 (O_2878,N_28003,N_29679);
and UO_2879 (O_2879,N_29094,N_28166);
nand UO_2880 (O_2880,N_29883,N_28717);
nand UO_2881 (O_2881,N_28802,N_28521);
nand UO_2882 (O_2882,N_29204,N_28570);
or UO_2883 (O_2883,N_28951,N_29907);
or UO_2884 (O_2884,N_28574,N_28594);
xor UO_2885 (O_2885,N_29286,N_29025);
nand UO_2886 (O_2886,N_29840,N_28805);
or UO_2887 (O_2887,N_29519,N_28780);
xor UO_2888 (O_2888,N_29927,N_29520);
xnor UO_2889 (O_2889,N_28283,N_28975);
and UO_2890 (O_2890,N_28393,N_29939);
or UO_2891 (O_2891,N_29089,N_28493);
xnor UO_2892 (O_2892,N_28159,N_28978);
nand UO_2893 (O_2893,N_29594,N_29887);
and UO_2894 (O_2894,N_28379,N_29599);
or UO_2895 (O_2895,N_29381,N_28174);
or UO_2896 (O_2896,N_29175,N_29505);
or UO_2897 (O_2897,N_28325,N_28309);
xnor UO_2898 (O_2898,N_29364,N_29191);
or UO_2899 (O_2899,N_28775,N_28647);
and UO_2900 (O_2900,N_28600,N_29545);
and UO_2901 (O_2901,N_29560,N_28442);
nor UO_2902 (O_2902,N_29618,N_29140);
or UO_2903 (O_2903,N_28505,N_29069);
xnor UO_2904 (O_2904,N_29036,N_29767);
nand UO_2905 (O_2905,N_28324,N_28834);
and UO_2906 (O_2906,N_29420,N_28068);
nand UO_2907 (O_2907,N_28153,N_28154);
nand UO_2908 (O_2908,N_28867,N_29144);
and UO_2909 (O_2909,N_29016,N_29013);
and UO_2910 (O_2910,N_29523,N_29421);
nand UO_2911 (O_2911,N_29363,N_28899);
nand UO_2912 (O_2912,N_29452,N_29035);
nor UO_2913 (O_2913,N_28902,N_28997);
xnor UO_2914 (O_2914,N_29607,N_29389);
nor UO_2915 (O_2915,N_28773,N_29880);
and UO_2916 (O_2916,N_29704,N_28297);
or UO_2917 (O_2917,N_28561,N_29798);
nor UO_2918 (O_2918,N_28562,N_29541);
or UO_2919 (O_2919,N_29920,N_29984);
and UO_2920 (O_2920,N_28978,N_28657);
and UO_2921 (O_2921,N_29223,N_28244);
or UO_2922 (O_2922,N_29289,N_28304);
nor UO_2923 (O_2923,N_28976,N_29737);
nor UO_2924 (O_2924,N_28997,N_28386);
nor UO_2925 (O_2925,N_28029,N_28111);
nor UO_2926 (O_2926,N_29031,N_29640);
or UO_2927 (O_2927,N_28319,N_28492);
xnor UO_2928 (O_2928,N_29211,N_28469);
or UO_2929 (O_2929,N_28946,N_29837);
or UO_2930 (O_2930,N_29697,N_29461);
and UO_2931 (O_2931,N_29869,N_29547);
and UO_2932 (O_2932,N_29238,N_29453);
or UO_2933 (O_2933,N_29390,N_28047);
and UO_2934 (O_2934,N_28394,N_29562);
nor UO_2935 (O_2935,N_29792,N_29651);
or UO_2936 (O_2936,N_28191,N_28651);
and UO_2937 (O_2937,N_29809,N_29933);
nor UO_2938 (O_2938,N_28679,N_29614);
nor UO_2939 (O_2939,N_28954,N_29348);
xor UO_2940 (O_2940,N_29171,N_29608);
and UO_2941 (O_2941,N_29507,N_29699);
nor UO_2942 (O_2942,N_29921,N_28837);
or UO_2943 (O_2943,N_28944,N_28273);
nand UO_2944 (O_2944,N_28817,N_28952);
and UO_2945 (O_2945,N_29794,N_28465);
nor UO_2946 (O_2946,N_28209,N_29248);
and UO_2947 (O_2947,N_29178,N_28395);
nand UO_2948 (O_2948,N_29917,N_28863);
xnor UO_2949 (O_2949,N_28881,N_28723);
xnor UO_2950 (O_2950,N_28203,N_28788);
or UO_2951 (O_2951,N_29882,N_28887);
and UO_2952 (O_2952,N_28479,N_28953);
xor UO_2953 (O_2953,N_28871,N_29524);
and UO_2954 (O_2954,N_29860,N_28571);
nand UO_2955 (O_2955,N_29026,N_29639);
or UO_2956 (O_2956,N_29938,N_29103);
nor UO_2957 (O_2957,N_28880,N_29603);
nor UO_2958 (O_2958,N_28773,N_29809);
nand UO_2959 (O_2959,N_28356,N_29594);
xnor UO_2960 (O_2960,N_29055,N_29615);
and UO_2961 (O_2961,N_29699,N_29109);
nand UO_2962 (O_2962,N_28512,N_29058);
xnor UO_2963 (O_2963,N_28369,N_28202);
or UO_2964 (O_2964,N_28152,N_29676);
nor UO_2965 (O_2965,N_29615,N_28472);
and UO_2966 (O_2966,N_29593,N_28896);
nor UO_2967 (O_2967,N_28191,N_29608);
and UO_2968 (O_2968,N_28370,N_29584);
or UO_2969 (O_2969,N_29360,N_29985);
xor UO_2970 (O_2970,N_29064,N_29859);
xnor UO_2971 (O_2971,N_29346,N_29629);
xor UO_2972 (O_2972,N_28310,N_29945);
nand UO_2973 (O_2973,N_29619,N_28043);
nand UO_2974 (O_2974,N_28958,N_29198);
or UO_2975 (O_2975,N_29094,N_28495);
or UO_2976 (O_2976,N_29050,N_28223);
or UO_2977 (O_2977,N_29421,N_28706);
or UO_2978 (O_2978,N_29246,N_28276);
or UO_2979 (O_2979,N_29315,N_29773);
nor UO_2980 (O_2980,N_29853,N_29198);
xor UO_2981 (O_2981,N_28069,N_29442);
and UO_2982 (O_2982,N_28659,N_28103);
nor UO_2983 (O_2983,N_28356,N_29933);
nand UO_2984 (O_2984,N_29260,N_29721);
or UO_2985 (O_2985,N_29740,N_28239);
nor UO_2986 (O_2986,N_29721,N_29435);
nand UO_2987 (O_2987,N_29397,N_29033);
or UO_2988 (O_2988,N_28235,N_28412);
and UO_2989 (O_2989,N_29750,N_29213);
or UO_2990 (O_2990,N_28003,N_28460);
or UO_2991 (O_2991,N_28027,N_29701);
nor UO_2992 (O_2992,N_29120,N_28241);
nor UO_2993 (O_2993,N_28152,N_29625);
and UO_2994 (O_2994,N_28538,N_28167);
and UO_2995 (O_2995,N_28839,N_29016);
and UO_2996 (O_2996,N_28762,N_28910);
xnor UO_2997 (O_2997,N_29195,N_28464);
nand UO_2998 (O_2998,N_28107,N_28932);
and UO_2999 (O_2999,N_28810,N_29256);
nor UO_3000 (O_3000,N_28719,N_28734);
or UO_3001 (O_3001,N_28983,N_29675);
and UO_3002 (O_3002,N_28388,N_28265);
xor UO_3003 (O_3003,N_28071,N_28219);
and UO_3004 (O_3004,N_29516,N_28470);
or UO_3005 (O_3005,N_28422,N_29238);
and UO_3006 (O_3006,N_28210,N_29497);
nor UO_3007 (O_3007,N_28242,N_28187);
or UO_3008 (O_3008,N_28342,N_28110);
and UO_3009 (O_3009,N_29225,N_28307);
nand UO_3010 (O_3010,N_29398,N_28651);
and UO_3011 (O_3011,N_29274,N_29565);
or UO_3012 (O_3012,N_29766,N_28943);
or UO_3013 (O_3013,N_29103,N_29313);
xor UO_3014 (O_3014,N_28958,N_28317);
and UO_3015 (O_3015,N_28415,N_28729);
nor UO_3016 (O_3016,N_28836,N_29203);
xnor UO_3017 (O_3017,N_28032,N_28511);
or UO_3018 (O_3018,N_28043,N_28215);
nor UO_3019 (O_3019,N_28577,N_28045);
and UO_3020 (O_3020,N_28633,N_29130);
or UO_3021 (O_3021,N_29605,N_29540);
nor UO_3022 (O_3022,N_28780,N_29508);
or UO_3023 (O_3023,N_29241,N_29089);
nor UO_3024 (O_3024,N_29335,N_29176);
nor UO_3025 (O_3025,N_29647,N_29780);
nor UO_3026 (O_3026,N_29237,N_29460);
and UO_3027 (O_3027,N_28029,N_28556);
or UO_3028 (O_3028,N_28974,N_29365);
and UO_3029 (O_3029,N_28542,N_28465);
nand UO_3030 (O_3030,N_29738,N_28602);
nand UO_3031 (O_3031,N_28082,N_29403);
and UO_3032 (O_3032,N_28238,N_28387);
nand UO_3033 (O_3033,N_28776,N_28536);
nor UO_3034 (O_3034,N_28402,N_29540);
and UO_3035 (O_3035,N_29016,N_29846);
nand UO_3036 (O_3036,N_28451,N_29380);
xor UO_3037 (O_3037,N_28960,N_29793);
nand UO_3038 (O_3038,N_28360,N_29738);
nor UO_3039 (O_3039,N_29980,N_28326);
and UO_3040 (O_3040,N_29539,N_28251);
nor UO_3041 (O_3041,N_28310,N_29804);
xor UO_3042 (O_3042,N_28282,N_29127);
or UO_3043 (O_3043,N_29468,N_29181);
and UO_3044 (O_3044,N_29308,N_29589);
or UO_3045 (O_3045,N_28196,N_28599);
and UO_3046 (O_3046,N_29884,N_28694);
nand UO_3047 (O_3047,N_28132,N_28589);
xor UO_3048 (O_3048,N_28005,N_28204);
xnor UO_3049 (O_3049,N_28683,N_28188);
or UO_3050 (O_3050,N_28425,N_28368);
or UO_3051 (O_3051,N_29747,N_28109);
or UO_3052 (O_3052,N_29596,N_29964);
xor UO_3053 (O_3053,N_28908,N_28757);
and UO_3054 (O_3054,N_29143,N_28281);
and UO_3055 (O_3055,N_28661,N_28582);
and UO_3056 (O_3056,N_28965,N_29016);
and UO_3057 (O_3057,N_29155,N_28518);
nor UO_3058 (O_3058,N_29008,N_29452);
or UO_3059 (O_3059,N_28598,N_28451);
nor UO_3060 (O_3060,N_29104,N_28522);
xnor UO_3061 (O_3061,N_28736,N_28985);
nor UO_3062 (O_3062,N_28482,N_29637);
nand UO_3063 (O_3063,N_29501,N_29235);
xnor UO_3064 (O_3064,N_29282,N_28622);
and UO_3065 (O_3065,N_29326,N_29920);
or UO_3066 (O_3066,N_28996,N_28437);
xnor UO_3067 (O_3067,N_29747,N_29082);
xor UO_3068 (O_3068,N_28097,N_28808);
nor UO_3069 (O_3069,N_28186,N_28760);
and UO_3070 (O_3070,N_29459,N_29698);
and UO_3071 (O_3071,N_29885,N_28614);
nand UO_3072 (O_3072,N_29971,N_28957);
nor UO_3073 (O_3073,N_28599,N_28377);
nor UO_3074 (O_3074,N_28680,N_28381);
or UO_3075 (O_3075,N_29530,N_28731);
or UO_3076 (O_3076,N_29772,N_29022);
xor UO_3077 (O_3077,N_29774,N_29177);
xor UO_3078 (O_3078,N_29558,N_29070);
and UO_3079 (O_3079,N_28347,N_28006);
xor UO_3080 (O_3080,N_28271,N_29689);
nand UO_3081 (O_3081,N_28541,N_28109);
xnor UO_3082 (O_3082,N_29389,N_28545);
nand UO_3083 (O_3083,N_29311,N_29484);
nand UO_3084 (O_3084,N_28497,N_28545);
or UO_3085 (O_3085,N_28257,N_28306);
xnor UO_3086 (O_3086,N_29219,N_29848);
xor UO_3087 (O_3087,N_29498,N_29197);
nand UO_3088 (O_3088,N_29664,N_29232);
xor UO_3089 (O_3089,N_28635,N_28553);
and UO_3090 (O_3090,N_28073,N_28870);
and UO_3091 (O_3091,N_29798,N_29296);
or UO_3092 (O_3092,N_29834,N_28795);
or UO_3093 (O_3093,N_29128,N_29823);
xor UO_3094 (O_3094,N_29721,N_29295);
nor UO_3095 (O_3095,N_28667,N_28476);
nor UO_3096 (O_3096,N_29462,N_29608);
nor UO_3097 (O_3097,N_28871,N_28462);
and UO_3098 (O_3098,N_28419,N_28121);
xnor UO_3099 (O_3099,N_29820,N_28963);
nor UO_3100 (O_3100,N_29806,N_29683);
nand UO_3101 (O_3101,N_28286,N_28148);
or UO_3102 (O_3102,N_29778,N_29290);
and UO_3103 (O_3103,N_28926,N_29676);
xnor UO_3104 (O_3104,N_28914,N_29489);
or UO_3105 (O_3105,N_28858,N_29309);
xnor UO_3106 (O_3106,N_29736,N_28494);
nand UO_3107 (O_3107,N_29224,N_29805);
nand UO_3108 (O_3108,N_29822,N_28546);
xnor UO_3109 (O_3109,N_28946,N_28282);
or UO_3110 (O_3110,N_28155,N_28512);
or UO_3111 (O_3111,N_29601,N_29047);
xor UO_3112 (O_3112,N_29057,N_28891);
or UO_3113 (O_3113,N_29875,N_28473);
nand UO_3114 (O_3114,N_28827,N_29576);
and UO_3115 (O_3115,N_28147,N_28900);
nor UO_3116 (O_3116,N_28566,N_29024);
nand UO_3117 (O_3117,N_29065,N_29972);
xnor UO_3118 (O_3118,N_28071,N_28311);
or UO_3119 (O_3119,N_29687,N_28824);
nor UO_3120 (O_3120,N_29314,N_28587);
xnor UO_3121 (O_3121,N_29712,N_29277);
and UO_3122 (O_3122,N_28089,N_28485);
xor UO_3123 (O_3123,N_28418,N_29991);
nor UO_3124 (O_3124,N_29146,N_29578);
or UO_3125 (O_3125,N_28734,N_29934);
xor UO_3126 (O_3126,N_28661,N_29887);
or UO_3127 (O_3127,N_29770,N_29454);
or UO_3128 (O_3128,N_29330,N_28487);
nor UO_3129 (O_3129,N_28019,N_29223);
xnor UO_3130 (O_3130,N_28436,N_28787);
nor UO_3131 (O_3131,N_29741,N_29755);
nand UO_3132 (O_3132,N_29823,N_29877);
nand UO_3133 (O_3133,N_28417,N_29624);
or UO_3134 (O_3134,N_29897,N_29906);
xor UO_3135 (O_3135,N_29364,N_28702);
xor UO_3136 (O_3136,N_29116,N_28160);
nand UO_3137 (O_3137,N_28485,N_29901);
nor UO_3138 (O_3138,N_29929,N_28673);
nand UO_3139 (O_3139,N_29113,N_28611);
and UO_3140 (O_3140,N_29495,N_28762);
or UO_3141 (O_3141,N_29877,N_29844);
xor UO_3142 (O_3142,N_28849,N_29132);
and UO_3143 (O_3143,N_28888,N_29368);
nor UO_3144 (O_3144,N_29521,N_28577);
nor UO_3145 (O_3145,N_29836,N_28673);
and UO_3146 (O_3146,N_28611,N_28868);
or UO_3147 (O_3147,N_29190,N_29375);
or UO_3148 (O_3148,N_28289,N_28105);
and UO_3149 (O_3149,N_28198,N_29480);
xor UO_3150 (O_3150,N_29203,N_28153);
and UO_3151 (O_3151,N_28112,N_28462);
and UO_3152 (O_3152,N_29542,N_29249);
and UO_3153 (O_3153,N_28031,N_28515);
and UO_3154 (O_3154,N_29684,N_29414);
xnor UO_3155 (O_3155,N_29912,N_28501);
and UO_3156 (O_3156,N_29204,N_28266);
xnor UO_3157 (O_3157,N_29792,N_28627);
and UO_3158 (O_3158,N_29244,N_29329);
nand UO_3159 (O_3159,N_29605,N_29262);
or UO_3160 (O_3160,N_29208,N_29425);
nand UO_3161 (O_3161,N_29820,N_28611);
and UO_3162 (O_3162,N_28808,N_28648);
nor UO_3163 (O_3163,N_29908,N_29031);
nor UO_3164 (O_3164,N_28483,N_28061);
and UO_3165 (O_3165,N_28718,N_28517);
xnor UO_3166 (O_3166,N_28038,N_28901);
or UO_3167 (O_3167,N_28749,N_29986);
nand UO_3168 (O_3168,N_28244,N_29149);
or UO_3169 (O_3169,N_29409,N_29035);
nor UO_3170 (O_3170,N_28140,N_29541);
nand UO_3171 (O_3171,N_29407,N_28789);
xnor UO_3172 (O_3172,N_28753,N_29397);
and UO_3173 (O_3173,N_28742,N_28496);
nand UO_3174 (O_3174,N_28816,N_28855);
or UO_3175 (O_3175,N_28859,N_29127);
nor UO_3176 (O_3176,N_28103,N_28410);
and UO_3177 (O_3177,N_28910,N_28968);
nand UO_3178 (O_3178,N_29137,N_28458);
nand UO_3179 (O_3179,N_28177,N_29168);
nor UO_3180 (O_3180,N_28966,N_28714);
or UO_3181 (O_3181,N_28375,N_28245);
xnor UO_3182 (O_3182,N_29997,N_29503);
nand UO_3183 (O_3183,N_29302,N_28138);
nor UO_3184 (O_3184,N_28583,N_29001);
and UO_3185 (O_3185,N_28212,N_29840);
xnor UO_3186 (O_3186,N_28376,N_29430);
nor UO_3187 (O_3187,N_29165,N_28639);
nand UO_3188 (O_3188,N_28046,N_28675);
nand UO_3189 (O_3189,N_28358,N_28882);
nand UO_3190 (O_3190,N_28332,N_28411);
nand UO_3191 (O_3191,N_29960,N_29577);
or UO_3192 (O_3192,N_28766,N_29813);
and UO_3193 (O_3193,N_28522,N_28550);
nand UO_3194 (O_3194,N_29202,N_29443);
and UO_3195 (O_3195,N_28183,N_29620);
nand UO_3196 (O_3196,N_28364,N_29775);
xor UO_3197 (O_3197,N_28515,N_29605);
xnor UO_3198 (O_3198,N_29271,N_29321);
or UO_3199 (O_3199,N_28474,N_29308);
or UO_3200 (O_3200,N_29077,N_28343);
or UO_3201 (O_3201,N_29159,N_29902);
xnor UO_3202 (O_3202,N_29157,N_28521);
or UO_3203 (O_3203,N_29499,N_28562);
and UO_3204 (O_3204,N_29656,N_29341);
and UO_3205 (O_3205,N_28082,N_28820);
xnor UO_3206 (O_3206,N_28902,N_29437);
and UO_3207 (O_3207,N_29697,N_29621);
nor UO_3208 (O_3208,N_29252,N_29792);
nand UO_3209 (O_3209,N_28896,N_29264);
nand UO_3210 (O_3210,N_29237,N_28845);
nor UO_3211 (O_3211,N_28569,N_29251);
nand UO_3212 (O_3212,N_28748,N_28339);
and UO_3213 (O_3213,N_29794,N_28060);
nor UO_3214 (O_3214,N_28118,N_28238);
nor UO_3215 (O_3215,N_29713,N_29521);
nor UO_3216 (O_3216,N_29228,N_29767);
or UO_3217 (O_3217,N_28057,N_29774);
or UO_3218 (O_3218,N_28005,N_29028);
or UO_3219 (O_3219,N_29169,N_29108);
nand UO_3220 (O_3220,N_29967,N_29088);
nand UO_3221 (O_3221,N_29190,N_28121);
and UO_3222 (O_3222,N_29346,N_29147);
xnor UO_3223 (O_3223,N_29450,N_29694);
nand UO_3224 (O_3224,N_29251,N_28105);
nor UO_3225 (O_3225,N_29561,N_28708);
or UO_3226 (O_3226,N_29090,N_29134);
and UO_3227 (O_3227,N_28523,N_28145);
xnor UO_3228 (O_3228,N_29106,N_29353);
xor UO_3229 (O_3229,N_29000,N_29596);
nand UO_3230 (O_3230,N_29270,N_28051);
nand UO_3231 (O_3231,N_28186,N_28930);
and UO_3232 (O_3232,N_28895,N_28498);
or UO_3233 (O_3233,N_29346,N_28476);
nand UO_3234 (O_3234,N_28651,N_29432);
nand UO_3235 (O_3235,N_29927,N_28896);
xor UO_3236 (O_3236,N_28476,N_28351);
nor UO_3237 (O_3237,N_28110,N_28884);
and UO_3238 (O_3238,N_28338,N_28768);
or UO_3239 (O_3239,N_29244,N_28548);
or UO_3240 (O_3240,N_28474,N_28266);
nand UO_3241 (O_3241,N_29296,N_29386);
and UO_3242 (O_3242,N_28730,N_28339);
xnor UO_3243 (O_3243,N_28450,N_29974);
nor UO_3244 (O_3244,N_29846,N_28555);
nor UO_3245 (O_3245,N_29582,N_28796);
nor UO_3246 (O_3246,N_28785,N_29441);
nor UO_3247 (O_3247,N_28048,N_29054);
or UO_3248 (O_3248,N_29590,N_28223);
nor UO_3249 (O_3249,N_29400,N_29471);
nand UO_3250 (O_3250,N_28759,N_28853);
xor UO_3251 (O_3251,N_29940,N_29615);
nand UO_3252 (O_3252,N_28950,N_28982);
nor UO_3253 (O_3253,N_28991,N_29080);
xor UO_3254 (O_3254,N_28729,N_29249);
nand UO_3255 (O_3255,N_28921,N_28211);
nand UO_3256 (O_3256,N_28142,N_29403);
and UO_3257 (O_3257,N_29654,N_29101);
or UO_3258 (O_3258,N_28172,N_28264);
or UO_3259 (O_3259,N_28134,N_28232);
nor UO_3260 (O_3260,N_29407,N_28038);
nand UO_3261 (O_3261,N_28615,N_29290);
and UO_3262 (O_3262,N_28959,N_28019);
nor UO_3263 (O_3263,N_28623,N_29801);
and UO_3264 (O_3264,N_29509,N_29474);
or UO_3265 (O_3265,N_28635,N_29887);
xor UO_3266 (O_3266,N_29589,N_28911);
nor UO_3267 (O_3267,N_29075,N_28768);
nor UO_3268 (O_3268,N_29589,N_29389);
nand UO_3269 (O_3269,N_29874,N_29568);
and UO_3270 (O_3270,N_28927,N_28903);
nand UO_3271 (O_3271,N_29307,N_29948);
nor UO_3272 (O_3272,N_28013,N_28661);
nand UO_3273 (O_3273,N_29520,N_28216);
xor UO_3274 (O_3274,N_29134,N_28023);
nand UO_3275 (O_3275,N_28509,N_29699);
and UO_3276 (O_3276,N_29981,N_29485);
xor UO_3277 (O_3277,N_29355,N_28289);
or UO_3278 (O_3278,N_28781,N_28177);
and UO_3279 (O_3279,N_29604,N_29714);
or UO_3280 (O_3280,N_29432,N_28217);
nor UO_3281 (O_3281,N_29304,N_29632);
xor UO_3282 (O_3282,N_28365,N_28063);
nand UO_3283 (O_3283,N_28429,N_28663);
nand UO_3284 (O_3284,N_28876,N_28204);
and UO_3285 (O_3285,N_28901,N_28615);
or UO_3286 (O_3286,N_28277,N_29986);
nand UO_3287 (O_3287,N_29966,N_29373);
xor UO_3288 (O_3288,N_29325,N_29350);
or UO_3289 (O_3289,N_28630,N_29743);
and UO_3290 (O_3290,N_28276,N_29605);
xor UO_3291 (O_3291,N_28984,N_28374);
xor UO_3292 (O_3292,N_28750,N_29599);
or UO_3293 (O_3293,N_28062,N_28800);
nor UO_3294 (O_3294,N_29952,N_28234);
nand UO_3295 (O_3295,N_29346,N_29561);
nand UO_3296 (O_3296,N_29808,N_28595);
xnor UO_3297 (O_3297,N_29272,N_29675);
or UO_3298 (O_3298,N_28519,N_29380);
nand UO_3299 (O_3299,N_28572,N_29716);
nor UO_3300 (O_3300,N_29068,N_29086);
and UO_3301 (O_3301,N_29245,N_28267);
xor UO_3302 (O_3302,N_29260,N_28569);
xor UO_3303 (O_3303,N_28666,N_29335);
and UO_3304 (O_3304,N_28614,N_29320);
xor UO_3305 (O_3305,N_29520,N_29558);
nor UO_3306 (O_3306,N_29780,N_29600);
xor UO_3307 (O_3307,N_29020,N_28268);
xnor UO_3308 (O_3308,N_28792,N_29000);
and UO_3309 (O_3309,N_28328,N_28602);
or UO_3310 (O_3310,N_29074,N_29088);
or UO_3311 (O_3311,N_29543,N_29643);
or UO_3312 (O_3312,N_29696,N_29687);
xnor UO_3313 (O_3313,N_29929,N_29140);
nand UO_3314 (O_3314,N_28899,N_29119);
nand UO_3315 (O_3315,N_28431,N_29212);
and UO_3316 (O_3316,N_29675,N_29657);
and UO_3317 (O_3317,N_29979,N_28464);
nor UO_3318 (O_3318,N_29091,N_28850);
nand UO_3319 (O_3319,N_29070,N_29014);
and UO_3320 (O_3320,N_29563,N_29137);
nor UO_3321 (O_3321,N_28575,N_29834);
nand UO_3322 (O_3322,N_29153,N_29378);
and UO_3323 (O_3323,N_29565,N_29330);
and UO_3324 (O_3324,N_28509,N_29207);
nor UO_3325 (O_3325,N_29946,N_29668);
nor UO_3326 (O_3326,N_29731,N_29533);
and UO_3327 (O_3327,N_28678,N_28226);
xnor UO_3328 (O_3328,N_29903,N_28819);
and UO_3329 (O_3329,N_28477,N_28674);
xnor UO_3330 (O_3330,N_28374,N_28500);
xnor UO_3331 (O_3331,N_28584,N_28416);
xnor UO_3332 (O_3332,N_29649,N_28869);
nand UO_3333 (O_3333,N_29266,N_29150);
nand UO_3334 (O_3334,N_29795,N_29660);
xor UO_3335 (O_3335,N_28640,N_28425);
nor UO_3336 (O_3336,N_29494,N_29680);
nor UO_3337 (O_3337,N_28894,N_28484);
nand UO_3338 (O_3338,N_29894,N_29150);
or UO_3339 (O_3339,N_28560,N_28789);
nor UO_3340 (O_3340,N_29098,N_28002);
xor UO_3341 (O_3341,N_29387,N_29626);
nor UO_3342 (O_3342,N_29873,N_28089);
and UO_3343 (O_3343,N_28596,N_28304);
xor UO_3344 (O_3344,N_29762,N_28943);
nand UO_3345 (O_3345,N_29123,N_28559);
or UO_3346 (O_3346,N_29283,N_28048);
nor UO_3347 (O_3347,N_28661,N_29220);
xnor UO_3348 (O_3348,N_29944,N_29710);
xor UO_3349 (O_3349,N_28971,N_28275);
xnor UO_3350 (O_3350,N_28161,N_28083);
or UO_3351 (O_3351,N_29061,N_28051);
and UO_3352 (O_3352,N_28458,N_29887);
xnor UO_3353 (O_3353,N_28627,N_29895);
nor UO_3354 (O_3354,N_29982,N_28267);
or UO_3355 (O_3355,N_28428,N_29191);
nor UO_3356 (O_3356,N_28174,N_29287);
nand UO_3357 (O_3357,N_28133,N_29049);
xor UO_3358 (O_3358,N_29139,N_29059);
xor UO_3359 (O_3359,N_28206,N_29273);
xor UO_3360 (O_3360,N_28806,N_29913);
and UO_3361 (O_3361,N_28604,N_29188);
xor UO_3362 (O_3362,N_29424,N_28329);
xnor UO_3363 (O_3363,N_28902,N_28800);
nor UO_3364 (O_3364,N_29416,N_29128);
or UO_3365 (O_3365,N_28872,N_29550);
nand UO_3366 (O_3366,N_28705,N_28714);
xor UO_3367 (O_3367,N_29616,N_29229);
and UO_3368 (O_3368,N_29629,N_28007);
nor UO_3369 (O_3369,N_29826,N_29005);
and UO_3370 (O_3370,N_29915,N_29391);
or UO_3371 (O_3371,N_28526,N_29708);
nand UO_3372 (O_3372,N_29901,N_29706);
or UO_3373 (O_3373,N_29657,N_29241);
or UO_3374 (O_3374,N_29694,N_28136);
or UO_3375 (O_3375,N_28796,N_28996);
xor UO_3376 (O_3376,N_29652,N_28704);
nand UO_3377 (O_3377,N_29048,N_29225);
nand UO_3378 (O_3378,N_28352,N_28339);
or UO_3379 (O_3379,N_28201,N_28922);
xnor UO_3380 (O_3380,N_28058,N_29984);
or UO_3381 (O_3381,N_29305,N_28795);
or UO_3382 (O_3382,N_28056,N_29931);
nor UO_3383 (O_3383,N_28164,N_28667);
or UO_3384 (O_3384,N_28025,N_29810);
xor UO_3385 (O_3385,N_28527,N_28970);
nor UO_3386 (O_3386,N_29431,N_28797);
nand UO_3387 (O_3387,N_29615,N_28110);
nor UO_3388 (O_3388,N_28683,N_29912);
and UO_3389 (O_3389,N_29654,N_29881);
nand UO_3390 (O_3390,N_28160,N_28235);
and UO_3391 (O_3391,N_29298,N_28033);
xnor UO_3392 (O_3392,N_29181,N_29053);
xnor UO_3393 (O_3393,N_28780,N_28631);
nor UO_3394 (O_3394,N_28112,N_28894);
xor UO_3395 (O_3395,N_29154,N_29502);
or UO_3396 (O_3396,N_29388,N_28011);
xor UO_3397 (O_3397,N_28101,N_28357);
and UO_3398 (O_3398,N_28410,N_29562);
and UO_3399 (O_3399,N_29281,N_29608);
nor UO_3400 (O_3400,N_28247,N_28711);
xnor UO_3401 (O_3401,N_29008,N_28615);
or UO_3402 (O_3402,N_28441,N_29123);
and UO_3403 (O_3403,N_28399,N_29070);
and UO_3404 (O_3404,N_29453,N_29374);
nor UO_3405 (O_3405,N_28266,N_29636);
or UO_3406 (O_3406,N_29265,N_29714);
or UO_3407 (O_3407,N_29944,N_29157);
nor UO_3408 (O_3408,N_28180,N_28700);
or UO_3409 (O_3409,N_28662,N_29611);
nand UO_3410 (O_3410,N_28475,N_28662);
nor UO_3411 (O_3411,N_29742,N_29941);
or UO_3412 (O_3412,N_28969,N_28932);
nor UO_3413 (O_3413,N_28599,N_29750);
nand UO_3414 (O_3414,N_28990,N_29810);
and UO_3415 (O_3415,N_28439,N_28477);
nand UO_3416 (O_3416,N_28564,N_29188);
nand UO_3417 (O_3417,N_28302,N_28879);
and UO_3418 (O_3418,N_29988,N_29869);
nand UO_3419 (O_3419,N_29893,N_29765);
and UO_3420 (O_3420,N_28704,N_28502);
xnor UO_3421 (O_3421,N_28111,N_28304);
xnor UO_3422 (O_3422,N_29410,N_29709);
and UO_3423 (O_3423,N_28947,N_28512);
or UO_3424 (O_3424,N_28941,N_29247);
nand UO_3425 (O_3425,N_28378,N_29973);
and UO_3426 (O_3426,N_29363,N_28747);
and UO_3427 (O_3427,N_28418,N_28424);
or UO_3428 (O_3428,N_29378,N_29705);
and UO_3429 (O_3429,N_28975,N_29289);
or UO_3430 (O_3430,N_29570,N_28151);
and UO_3431 (O_3431,N_28656,N_29091);
nand UO_3432 (O_3432,N_28286,N_28192);
xor UO_3433 (O_3433,N_28490,N_28798);
nand UO_3434 (O_3434,N_28873,N_29816);
nor UO_3435 (O_3435,N_28909,N_28087);
xor UO_3436 (O_3436,N_28580,N_29199);
nand UO_3437 (O_3437,N_29259,N_28293);
or UO_3438 (O_3438,N_29786,N_29089);
xnor UO_3439 (O_3439,N_28576,N_29701);
nand UO_3440 (O_3440,N_28942,N_28264);
nor UO_3441 (O_3441,N_28827,N_28624);
or UO_3442 (O_3442,N_28730,N_29537);
nand UO_3443 (O_3443,N_28315,N_28528);
nor UO_3444 (O_3444,N_29571,N_28490);
nand UO_3445 (O_3445,N_29133,N_28804);
xnor UO_3446 (O_3446,N_28179,N_28669);
and UO_3447 (O_3447,N_29374,N_28711);
and UO_3448 (O_3448,N_29558,N_29289);
xnor UO_3449 (O_3449,N_28105,N_29077);
xor UO_3450 (O_3450,N_29141,N_29340);
xor UO_3451 (O_3451,N_28330,N_29155);
or UO_3452 (O_3452,N_29323,N_29366);
nor UO_3453 (O_3453,N_28699,N_28693);
xnor UO_3454 (O_3454,N_29033,N_28970);
xnor UO_3455 (O_3455,N_29778,N_28090);
and UO_3456 (O_3456,N_28503,N_28426);
xor UO_3457 (O_3457,N_29847,N_29364);
nor UO_3458 (O_3458,N_29166,N_29485);
or UO_3459 (O_3459,N_29949,N_28010);
and UO_3460 (O_3460,N_28394,N_28676);
or UO_3461 (O_3461,N_28231,N_29178);
nand UO_3462 (O_3462,N_28285,N_28471);
nor UO_3463 (O_3463,N_29561,N_29652);
nand UO_3464 (O_3464,N_29605,N_29051);
nor UO_3465 (O_3465,N_28316,N_28491);
or UO_3466 (O_3466,N_29399,N_28788);
nand UO_3467 (O_3467,N_28364,N_28325);
nor UO_3468 (O_3468,N_28944,N_28730);
nor UO_3469 (O_3469,N_28680,N_29781);
nor UO_3470 (O_3470,N_29734,N_29775);
nor UO_3471 (O_3471,N_29533,N_28932);
nor UO_3472 (O_3472,N_29837,N_28162);
or UO_3473 (O_3473,N_29966,N_29547);
nand UO_3474 (O_3474,N_28467,N_28562);
or UO_3475 (O_3475,N_29412,N_28133);
nand UO_3476 (O_3476,N_29056,N_28469);
or UO_3477 (O_3477,N_28398,N_29046);
or UO_3478 (O_3478,N_28534,N_29324);
nor UO_3479 (O_3479,N_28076,N_29329);
nor UO_3480 (O_3480,N_29881,N_28246);
xnor UO_3481 (O_3481,N_28292,N_28636);
xor UO_3482 (O_3482,N_29504,N_28039);
nand UO_3483 (O_3483,N_29050,N_29581);
nand UO_3484 (O_3484,N_29605,N_29800);
nand UO_3485 (O_3485,N_29978,N_29793);
nor UO_3486 (O_3486,N_29470,N_29489);
nand UO_3487 (O_3487,N_28277,N_28482);
or UO_3488 (O_3488,N_28019,N_29864);
xnor UO_3489 (O_3489,N_29189,N_29532);
and UO_3490 (O_3490,N_28228,N_29079);
or UO_3491 (O_3491,N_28988,N_29208);
and UO_3492 (O_3492,N_29551,N_28961);
nand UO_3493 (O_3493,N_28335,N_28098);
or UO_3494 (O_3494,N_29787,N_29289);
and UO_3495 (O_3495,N_29699,N_28573);
or UO_3496 (O_3496,N_29088,N_28912);
nor UO_3497 (O_3497,N_29873,N_29746);
nor UO_3498 (O_3498,N_28410,N_29165);
nor UO_3499 (O_3499,N_28412,N_29371);
endmodule