module basic_500_3000_500_40_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_127,In_207);
nand U1 (N_1,In_372,In_111);
or U2 (N_2,In_223,In_276);
nand U3 (N_3,In_295,In_343);
nor U4 (N_4,In_355,In_216);
or U5 (N_5,In_282,In_492);
and U6 (N_6,In_48,In_51);
and U7 (N_7,In_378,In_381);
or U8 (N_8,In_102,In_28);
nor U9 (N_9,In_497,In_93);
nor U10 (N_10,In_362,In_14);
nand U11 (N_11,In_297,In_442);
and U12 (N_12,In_142,In_323);
xor U13 (N_13,In_20,In_112);
xor U14 (N_14,In_346,In_166);
or U15 (N_15,In_59,In_107);
xor U16 (N_16,In_251,In_270);
xor U17 (N_17,In_13,In_244);
or U18 (N_18,In_65,In_337);
nor U19 (N_19,In_45,In_475);
nor U20 (N_20,In_214,In_481);
xor U21 (N_21,In_80,In_453);
xnor U22 (N_22,In_185,In_449);
nor U23 (N_23,In_479,In_370);
xor U24 (N_24,In_236,In_240);
or U25 (N_25,In_228,In_376);
and U26 (N_26,In_265,In_252);
nor U27 (N_27,In_458,In_472);
and U28 (N_28,In_73,In_291);
or U29 (N_29,In_336,In_243);
xnor U30 (N_30,In_206,In_181);
and U31 (N_31,In_180,In_115);
and U32 (N_32,In_198,In_79);
nand U33 (N_33,In_315,In_134);
and U34 (N_34,In_101,In_221);
and U35 (N_35,In_394,In_220);
nor U36 (N_36,In_173,In_229);
nor U37 (N_37,In_385,In_188);
nor U38 (N_38,In_470,In_304);
or U39 (N_39,In_130,In_390);
and U40 (N_40,In_190,In_247);
and U41 (N_41,In_170,In_47);
and U42 (N_42,In_483,In_361);
and U43 (N_43,In_363,In_420);
nor U44 (N_44,In_8,In_338);
or U45 (N_45,In_283,In_113);
and U46 (N_46,In_482,In_91);
xor U47 (N_47,In_488,In_473);
xnor U48 (N_48,In_409,In_259);
nor U49 (N_49,In_135,In_201);
or U50 (N_50,In_10,In_341);
and U51 (N_51,In_143,In_37);
or U52 (N_52,In_396,In_395);
xor U53 (N_53,In_455,In_391);
nor U54 (N_54,In_212,In_52);
nor U55 (N_55,In_490,In_493);
nand U56 (N_56,In_7,In_242);
or U57 (N_57,In_208,In_99);
nor U58 (N_58,In_429,In_196);
xnor U59 (N_59,In_366,In_157);
nand U60 (N_60,In_219,In_86);
xor U61 (N_61,In_178,In_64);
xor U62 (N_62,In_21,In_271);
or U63 (N_63,In_422,In_72);
nor U64 (N_64,In_284,In_414);
xor U65 (N_65,In_81,In_119);
or U66 (N_66,In_9,In_68);
xor U67 (N_67,In_485,In_36);
xnor U68 (N_68,In_451,In_76);
and U69 (N_69,In_1,In_330);
and U70 (N_70,In_75,In_0);
and U71 (N_71,In_344,In_371);
and U72 (N_72,In_167,In_11);
xnor U73 (N_73,In_327,In_224);
nand U74 (N_74,In_313,In_419);
xnor U75 (N_75,In_233,In_268);
and U76 (N_76,In_487,In_289);
or U77 (N_77,In_95,In_345);
or U78 (N_78,In_300,In_12);
nor U79 (N_79,N_51,In_164);
xor U80 (N_80,In_88,In_132);
and U81 (N_81,In_110,In_24);
and U82 (N_82,In_447,In_23);
and U83 (N_83,In_392,N_52);
nor U84 (N_84,In_154,In_77);
nor U85 (N_85,In_286,In_160);
and U86 (N_86,In_287,In_58);
nor U87 (N_87,N_31,In_427);
or U88 (N_88,N_73,In_365);
nand U89 (N_89,In_298,In_386);
xor U90 (N_90,In_41,In_440);
nand U91 (N_91,In_263,In_17);
nor U92 (N_92,In_393,N_41);
or U93 (N_93,In_328,N_64);
nor U94 (N_94,In_177,In_147);
or U95 (N_95,N_32,In_83);
nor U96 (N_96,N_10,In_406);
and U97 (N_97,In_424,In_197);
nor U98 (N_98,In_126,In_29);
xor U99 (N_99,In_98,N_55);
or U100 (N_100,In_278,In_184);
or U101 (N_101,In_261,In_159);
or U102 (N_102,In_31,In_257);
or U103 (N_103,In_152,In_137);
and U104 (N_104,In_74,In_27);
or U105 (N_105,In_90,In_163);
xor U106 (N_106,In_39,In_433);
or U107 (N_107,In_303,In_443);
xor U108 (N_108,N_57,N_24);
nor U109 (N_109,In_441,In_404);
nand U110 (N_110,In_250,In_253);
and U111 (N_111,In_174,In_122);
nor U112 (N_112,N_56,N_33);
nor U113 (N_113,N_30,In_105);
and U114 (N_114,In_260,N_36);
xnor U115 (N_115,In_462,In_4);
nand U116 (N_116,N_12,In_437);
xnor U117 (N_117,N_43,In_375);
nor U118 (N_118,N_8,In_281);
nor U119 (N_119,In_418,In_210);
and U120 (N_120,In_168,In_117);
xnor U121 (N_121,In_156,In_353);
or U122 (N_122,In_349,In_499);
nand U123 (N_123,In_494,In_162);
nand U124 (N_124,In_288,In_231);
nor U125 (N_125,In_428,In_3);
nor U126 (N_126,In_426,In_311);
nand U127 (N_127,In_457,N_44);
and U128 (N_128,In_348,In_292);
xnor U129 (N_129,In_33,In_465);
or U130 (N_130,In_118,In_123);
nand U131 (N_131,In_466,In_397);
nor U132 (N_132,N_38,In_193);
and U133 (N_133,In_6,In_96);
xnor U134 (N_134,In_321,In_32);
and U135 (N_135,In_171,In_301);
or U136 (N_136,In_408,In_498);
nor U137 (N_137,In_120,In_71);
or U138 (N_138,N_14,In_367);
nand U139 (N_139,N_40,N_67);
or U140 (N_140,In_484,In_149);
nand U141 (N_141,In_213,In_275);
or U142 (N_142,N_23,In_104);
or U143 (N_143,In_238,In_186);
nor U144 (N_144,In_266,In_432);
nor U145 (N_145,In_460,In_279);
and U146 (N_146,In_205,In_165);
nor U147 (N_147,N_34,In_489);
xor U148 (N_148,N_15,In_176);
and U149 (N_149,In_44,N_37);
nor U150 (N_150,N_112,In_255);
nand U151 (N_151,In_30,N_110);
and U152 (N_152,In_187,N_115);
nand U153 (N_153,N_16,N_58);
xnor U154 (N_154,In_351,N_146);
nand U155 (N_155,In_431,N_91);
nand U156 (N_156,In_438,N_26);
nand U157 (N_157,In_241,In_446);
nand U158 (N_158,In_218,In_182);
nand U159 (N_159,In_459,In_425);
nor U160 (N_160,N_116,N_61);
xnor U161 (N_161,In_245,In_89);
nand U162 (N_162,In_309,In_379);
or U163 (N_163,N_28,In_435);
nor U164 (N_164,In_129,In_399);
xnor U165 (N_165,In_85,In_2);
nand U166 (N_166,N_6,N_128);
nor U167 (N_167,In_380,In_121);
nand U168 (N_168,In_153,In_342);
or U169 (N_169,In_320,In_161);
and U170 (N_170,In_421,In_50);
xor U171 (N_171,N_66,In_139);
nand U172 (N_172,In_388,In_100);
xor U173 (N_173,N_22,In_230);
and U174 (N_174,In_329,In_175);
nor U175 (N_175,In_352,In_25);
nand U176 (N_176,In_310,In_467);
nand U177 (N_177,In_317,N_69);
nand U178 (N_178,In_179,In_172);
nand U179 (N_179,N_42,N_96);
xnor U180 (N_180,In_114,In_62);
nand U181 (N_181,N_21,In_412);
nand U182 (N_182,In_146,In_215);
nor U183 (N_183,N_90,In_128);
and U184 (N_184,N_45,In_34);
or U185 (N_185,N_106,In_359);
nor U186 (N_186,N_80,N_11);
or U187 (N_187,N_105,In_464);
and U188 (N_188,In_290,N_50);
nor U189 (N_189,In_326,In_456);
or U190 (N_190,In_67,In_273);
or U191 (N_191,N_139,In_200);
and U192 (N_192,In_314,In_192);
or U193 (N_193,In_293,In_203);
or U194 (N_194,N_7,In_299);
xnor U195 (N_195,In_97,In_264);
xor U196 (N_196,N_93,N_63);
and U197 (N_197,In_254,In_439);
or U198 (N_198,In_61,N_123);
or U199 (N_199,In_140,N_77);
xor U200 (N_200,In_148,In_354);
nor U201 (N_201,N_48,N_39);
or U202 (N_202,In_384,N_72);
xnor U203 (N_203,In_225,N_95);
or U204 (N_204,In_491,In_331);
xor U205 (N_205,In_5,In_237);
nand U206 (N_206,N_13,N_46);
or U207 (N_207,N_136,N_125);
xnor U208 (N_208,In_249,In_461);
and U209 (N_209,In_138,In_26);
nor U210 (N_210,N_133,In_46);
nor U211 (N_211,N_74,N_19);
and U212 (N_212,N_111,N_86);
nor U213 (N_213,In_158,In_169);
nor U214 (N_214,N_101,In_125);
xnor U215 (N_215,In_16,In_478);
and U216 (N_216,In_410,In_191);
xor U217 (N_217,N_147,In_407);
and U218 (N_218,In_53,N_49);
nor U219 (N_219,N_92,In_217);
and U220 (N_220,N_5,In_108);
xor U221 (N_221,In_22,N_113);
nand U222 (N_222,N_138,In_54);
xor U223 (N_223,N_75,In_66);
nor U224 (N_224,In_222,N_29);
nor U225 (N_225,N_177,N_65);
or U226 (N_226,N_179,N_201);
or U227 (N_227,In_350,N_195);
or U228 (N_228,N_224,N_126);
or U229 (N_229,In_377,N_193);
nor U230 (N_230,N_202,N_59);
or U231 (N_231,N_71,N_214);
xor U232 (N_232,In_280,In_486);
xnor U233 (N_233,In_382,In_204);
nor U234 (N_234,In_209,N_185);
nor U235 (N_235,In_103,N_194);
nand U236 (N_236,In_106,N_180);
nor U237 (N_237,In_468,In_415);
xnor U238 (N_238,N_166,N_109);
or U239 (N_239,In_63,In_199);
or U240 (N_240,In_450,N_78);
and U241 (N_241,N_25,In_306);
nor U242 (N_242,N_187,In_189);
nor U243 (N_243,In_194,In_340);
and U244 (N_244,N_221,N_134);
nand U245 (N_245,N_216,In_302);
xnor U246 (N_246,In_133,N_4);
or U247 (N_247,N_114,In_389);
xor U248 (N_248,N_169,In_423);
and U249 (N_249,In_471,N_18);
xnor U250 (N_250,In_307,In_92);
and U251 (N_251,N_100,In_38);
nand U252 (N_252,N_144,In_496);
nor U253 (N_253,N_127,In_454);
nor U254 (N_254,N_160,In_402);
nor U255 (N_255,In_144,N_121);
nand U256 (N_256,N_152,In_347);
nor U257 (N_257,N_17,N_182);
nand U258 (N_258,N_9,In_335);
nor U259 (N_259,N_119,In_87);
xnor U260 (N_260,In_124,N_184);
xnor U261 (N_261,In_416,In_294);
and U262 (N_262,N_186,N_178);
or U263 (N_263,N_130,In_19);
xor U264 (N_264,N_210,In_403);
and U265 (N_265,N_108,N_165);
xor U266 (N_266,N_197,In_43);
nand U267 (N_267,N_217,N_35);
and U268 (N_268,In_369,In_84);
nand U269 (N_269,N_137,In_131);
nor U270 (N_270,N_120,In_463);
xnor U271 (N_271,N_82,N_163);
xnor U272 (N_272,N_79,In_35);
and U273 (N_273,N_175,N_156);
nor U274 (N_274,N_173,N_200);
and U275 (N_275,N_206,N_209);
nand U276 (N_276,In_413,N_199);
or U277 (N_277,N_203,N_47);
nor U278 (N_278,In_151,In_82);
and U279 (N_279,In_411,N_222);
nor U280 (N_280,In_274,In_322);
and U281 (N_281,N_87,In_364);
and U282 (N_282,In_436,In_339);
and U283 (N_283,In_232,In_248);
xnor U284 (N_284,N_154,N_97);
xnor U285 (N_285,In_495,N_161);
nand U286 (N_286,N_159,In_296);
xor U287 (N_287,In_383,N_89);
and U288 (N_288,N_212,N_102);
nor U289 (N_289,N_129,N_70);
nand U290 (N_290,In_305,In_15);
or U291 (N_291,N_99,In_116);
and U292 (N_292,In_357,N_149);
or U293 (N_293,N_213,N_142);
xnor U294 (N_294,In_69,In_202);
xor U295 (N_295,In_476,In_49);
xnor U296 (N_296,In_183,In_42);
nand U297 (N_297,In_318,N_54);
and U298 (N_298,In_387,In_398);
nor U299 (N_299,In_258,In_57);
xor U300 (N_300,In_312,In_400);
nand U301 (N_301,N_191,N_60);
xor U302 (N_302,N_172,N_238);
or U303 (N_303,In_272,N_170);
nor U304 (N_304,N_265,N_183);
or U305 (N_305,N_150,N_245);
nor U306 (N_306,N_76,N_241);
and U307 (N_307,N_246,N_207);
xor U308 (N_308,N_223,N_215);
or U309 (N_309,N_225,N_274);
or U310 (N_310,N_263,In_325);
nand U311 (N_311,N_1,N_299);
or U312 (N_312,In_267,N_249);
nand U313 (N_313,N_252,N_275);
nor U314 (N_314,In_474,N_268);
xor U315 (N_315,N_198,N_255);
or U316 (N_316,N_167,In_401);
nor U317 (N_317,In_334,In_94);
and U318 (N_318,N_267,N_230);
nand U319 (N_319,N_155,N_288);
xor U320 (N_320,N_290,In_227);
xnor U321 (N_321,N_164,In_356);
nor U322 (N_322,N_242,N_151);
and U323 (N_323,In_316,In_60);
nor U324 (N_324,N_118,In_469);
xor U325 (N_325,N_84,N_2);
and U326 (N_326,N_143,N_189);
or U327 (N_327,In_246,N_219);
and U328 (N_328,N_282,N_253);
nor U329 (N_329,In_374,N_248);
or U330 (N_330,N_62,N_107);
xor U331 (N_331,N_289,N_281);
xor U332 (N_332,In_150,N_237);
or U333 (N_333,N_243,In_332);
or U334 (N_334,In_234,N_244);
nor U335 (N_335,N_266,N_81);
or U336 (N_336,N_284,N_251);
nand U337 (N_337,N_204,N_280);
nor U338 (N_338,N_285,N_291);
and U339 (N_339,In_235,N_20);
or U340 (N_340,N_132,In_333);
and U341 (N_341,N_258,N_273);
or U342 (N_342,N_188,N_27);
xnor U343 (N_343,N_234,N_98);
and U344 (N_344,N_3,In_211);
nand U345 (N_345,In_358,N_153);
or U346 (N_346,In_373,N_278);
xor U347 (N_347,N_103,N_171);
nand U348 (N_348,In_480,N_260);
xnor U349 (N_349,N_148,N_88);
xor U350 (N_350,N_233,In_195);
and U351 (N_351,N_272,N_218);
or U352 (N_352,In_285,N_83);
xor U353 (N_353,In_452,In_324);
nor U354 (N_354,N_264,N_279);
nand U355 (N_355,N_259,In_444);
nor U356 (N_356,N_262,In_262);
and U357 (N_357,N_158,In_136);
nand U358 (N_358,N_190,N_141);
nand U359 (N_359,In_445,N_122);
xor U360 (N_360,N_256,In_417);
nand U361 (N_361,N_261,N_117);
xor U362 (N_362,N_297,In_308);
nor U363 (N_363,N_276,N_140);
or U364 (N_364,N_226,N_168);
and U365 (N_365,In_448,N_298);
xor U366 (N_366,N_257,N_250);
nor U367 (N_367,N_247,N_270);
nor U368 (N_368,In_70,N_294);
or U369 (N_369,N_239,N_85);
and U370 (N_370,N_157,N_211);
xor U371 (N_371,In_18,In_319);
nor U372 (N_372,In_269,N_231);
and U373 (N_373,N_162,N_235);
and U374 (N_374,N_205,N_196);
nand U375 (N_375,N_332,N_271);
and U376 (N_376,N_232,N_372);
nand U377 (N_377,N_325,N_295);
and U378 (N_378,N_287,N_293);
nor U379 (N_379,N_316,N_339);
and U380 (N_380,N_94,N_220);
nor U381 (N_381,N_351,N_240);
nor U382 (N_382,N_307,N_334);
nand U383 (N_383,N_208,N_336);
xnor U384 (N_384,In_277,N_353);
and U385 (N_385,N_371,In_226);
nand U386 (N_386,N_365,N_292);
xor U387 (N_387,N_254,N_174);
xnor U388 (N_388,N_341,N_312);
or U389 (N_389,N_350,N_314);
nor U390 (N_390,N_361,N_370);
or U391 (N_391,N_313,N_344);
or U392 (N_392,N_296,N_328);
and U393 (N_393,N_304,N_342);
nand U394 (N_394,N_367,N_277);
or U395 (N_395,N_228,N_311);
and U396 (N_396,In_430,N_318);
nor U397 (N_397,N_355,N_352);
or U398 (N_398,N_340,In_56);
or U399 (N_399,N_323,N_368);
xor U400 (N_400,N_335,N_300);
and U401 (N_401,N_301,N_181);
nand U402 (N_402,N_236,N_331);
or U403 (N_403,In_40,N_135);
or U404 (N_404,N_283,N_326);
or U405 (N_405,N_104,N_357);
nor U406 (N_406,In_368,N_333);
and U407 (N_407,In_141,N_374);
nor U408 (N_408,N_349,In_256);
and U409 (N_409,N_322,N_68);
xnor U410 (N_410,N_324,N_303);
xor U411 (N_411,N_309,N_345);
nand U412 (N_412,N_362,N_346);
xor U413 (N_413,N_356,N_305);
and U414 (N_414,N_229,N_373);
or U415 (N_415,N_306,N_329);
nand U416 (N_416,In_55,N_369);
or U417 (N_417,N_319,N_269);
and U418 (N_418,In_78,N_321);
and U419 (N_419,In_239,N_359);
nor U420 (N_420,In_109,N_0);
and U421 (N_421,In_155,N_364);
nand U422 (N_422,N_363,N_343);
and U423 (N_423,In_405,N_337);
nor U424 (N_424,N_338,In_360);
nor U425 (N_425,N_366,N_192);
nor U426 (N_426,N_347,N_317);
nor U427 (N_427,N_320,In_477);
nand U428 (N_428,N_227,N_176);
nor U429 (N_429,N_327,N_348);
nand U430 (N_430,N_53,N_358);
or U431 (N_431,N_302,In_434);
or U432 (N_432,N_310,N_360);
nor U433 (N_433,N_308,N_286);
nor U434 (N_434,N_315,N_354);
nor U435 (N_435,N_124,N_131);
nand U436 (N_436,In_145,N_330);
and U437 (N_437,N_145,N_350);
xor U438 (N_438,N_283,N_295);
xor U439 (N_439,N_327,N_104);
and U440 (N_440,N_355,N_308);
and U441 (N_441,N_343,N_366);
nand U442 (N_442,N_240,In_78);
and U443 (N_443,N_344,In_256);
and U444 (N_444,N_332,N_313);
xnor U445 (N_445,N_349,N_327);
xnor U446 (N_446,N_311,N_337);
or U447 (N_447,N_332,N_316);
nand U448 (N_448,N_364,N_366);
or U449 (N_449,N_307,N_320);
xor U450 (N_450,N_430,N_382);
nor U451 (N_451,N_394,N_447);
nor U452 (N_452,N_378,N_409);
or U453 (N_453,N_403,N_421);
xor U454 (N_454,N_385,N_396);
nand U455 (N_455,N_386,N_445);
xor U456 (N_456,N_392,N_397);
and U457 (N_457,N_381,N_434);
and U458 (N_458,N_398,N_376);
xnor U459 (N_459,N_418,N_429);
nor U460 (N_460,N_390,N_395);
or U461 (N_461,N_414,N_415);
or U462 (N_462,N_375,N_432);
xor U463 (N_463,N_438,N_399);
or U464 (N_464,N_448,N_419);
nor U465 (N_465,N_393,N_391);
nand U466 (N_466,N_424,N_413);
nand U467 (N_467,N_431,N_389);
xnor U468 (N_468,N_443,N_405);
nand U469 (N_469,N_411,N_406);
or U470 (N_470,N_422,N_433);
nand U471 (N_471,N_423,N_449);
nand U472 (N_472,N_426,N_439);
xor U473 (N_473,N_420,N_402);
nand U474 (N_474,N_444,N_440);
and U475 (N_475,N_435,N_401);
xor U476 (N_476,N_427,N_383);
and U477 (N_477,N_412,N_446);
nor U478 (N_478,N_417,N_380);
nand U479 (N_479,N_425,N_379);
and U480 (N_480,N_442,N_410);
xor U481 (N_481,N_408,N_437);
nor U482 (N_482,N_384,N_404);
and U483 (N_483,N_377,N_400);
or U484 (N_484,N_407,N_441);
nor U485 (N_485,N_436,N_428);
xnor U486 (N_486,N_388,N_387);
or U487 (N_487,N_416,N_388);
or U488 (N_488,N_444,N_382);
xnor U489 (N_489,N_409,N_439);
xnor U490 (N_490,N_384,N_424);
nand U491 (N_491,N_448,N_430);
xnor U492 (N_492,N_414,N_434);
nor U493 (N_493,N_385,N_404);
nand U494 (N_494,N_395,N_446);
xor U495 (N_495,N_399,N_421);
nand U496 (N_496,N_447,N_414);
xnor U497 (N_497,N_420,N_424);
or U498 (N_498,N_442,N_424);
nand U499 (N_499,N_402,N_426);
xnor U500 (N_500,N_436,N_412);
xnor U501 (N_501,N_391,N_411);
nor U502 (N_502,N_441,N_424);
or U503 (N_503,N_448,N_433);
or U504 (N_504,N_399,N_393);
and U505 (N_505,N_447,N_422);
nor U506 (N_506,N_404,N_425);
xnor U507 (N_507,N_433,N_382);
and U508 (N_508,N_385,N_426);
or U509 (N_509,N_414,N_440);
and U510 (N_510,N_412,N_431);
and U511 (N_511,N_432,N_416);
xor U512 (N_512,N_383,N_439);
nand U513 (N_513,N_432,N_384);
and U514 (N_514,N_408,N_398);
or U515 (N_515,N_417,N_386);
nand U516 (N_516,N_442,N_377);
nand U517 (N_517,N_406,N_431);
nor U518 (N_518,N_443,N_433);
xor U519 (N_519,N_392,N_448);
nor U520 (N_520,N_404,N_392);
or U521 (N_521,N_437,N_432);
nor U522 (N_522,N_438,N_396);
nor U523 (N_523,N_382,N_415);
nand U524 (N_524,N_384,N_410);
xor U525 (N_525,N_458,N_474);
and U526 (N_526,N_475,N_473);
nor U527 (N_527,N_495,N_461);
xnor U528 (N_528,N_491,N_468);
or U529 (N_529,N_483,N_499);
xor U530 (N_530,N_524,N_459);
or U531 (N_531,N_500,N_471);
and U532 (N_532,N_479,N_456);
xor U533 (N_533,N_450,N_514);
nor U534 (N_534,N_511,N_487);
or U535 (N_535,N_455,N_463);
nor U536 (N_536,N_466,N_454);
nor U537 (N_537,N_465,N_451);
nor U538 (N_538,N_470,N_518);
nor U539 (N_539,N_453,N_472);
and U540 (N_540,N_507,N_478);
and U541 (N_541,N_515,N_488);
nor U542 (N_542,N_521,N_484);
nor U543 (N_543,N_496,N_481);
nor U544 (N_544,N_502,N_508);
nand U545 (N_545,N_510,N_489);
nor U546 (N_546,N_477,N_452);
and U547 (N_547,N_501,N_517);
or U548 (N_548,N_505,N_509);
and U549 (N_549,N_513,N_490);
xnor U550 (N_550,N_503,N_516);
nand U551 (N_551,N_467,N_482);
nor U552 (N_552,N_486,N_457);
xor U553 (N_553,N_523,N_485);
nand U554 (N_554,N_504,N_519);
nor U555 (N_555,N_464,N_469);
nand U556 (N_556,N_480,N_462);
nand U557 (N_557,N_497,N_493);
and U558 (N_558,N_460,N_522);
nand U559 (N_559,N_512,N_520);
xor U560 (N_560,N_506,N_498);
and U561 (N_561,N_476,N_492);
nand U562 (N_562,N_494,N_466);
or U563 (N_563,N_524,N_456);
or U564 (N_564,N_510,N_471);
nor U565 (N_565,N_485,N_499);
and U566 (N_566,N_482,N_509);
nand U567 (N_567,N_466,N_490);
xor U568 (N_568,N_483,N_498);
nand U569 (N_569,N_458,N_502);
xor U570 (N_570,N_495,N_498);
xnor U571 (N_571,N_454,N_492);
or U572 (N_572,N_516,N_487);
nand U573 (N_573,N_459,N_495);
or U574 (N_574,N_498,N_512);
and U575 (N_575,N_486,N_472);
xnor U576 (N_576,N_517,N_502);
or U577 (N_577,N_500,N_515);
xor U578 (N_578,N_479,N_523);
and U579 (N_579,N_484,N_462);
nand U580 (N_580,N_483,N_497);
nand U581 (N_581,N_464,N_478);
and U582 (N_582,N_473,N_485);
and U583 (N_583,N_455,N_483);
nor U584 (N_584,N_486,N_458);
and U585 (N_585,N_500,N_460);
nor U586 (N_586,N_468,N_504);
xnor U587 (N_587,N_487,N_450);
nor U588 (N_588,N_452,N_469);
and U589 (N_589,N_508,N_478);
and U590 (N_590,N_491,N_510);
xor U591 (N_591,N_490,N_524);
xor U592 (N_592,N_499,N_500);
xor U593 (N_593,N_489,N_478);
nand U594 (N_594,N_509,N_457);
or U595 (N_595,N_450,N_462);
and U596 (N_596,N_472,N_519);
or U597 (N_597,N_499,N_481);
nand U598 (N_598,N_472,N_479);
nand U599 (N_599,N_463,N_479);
nor U600 (N_600,N_578,N_573);
nand U601 (N_601,N_543,N_561);
or U602 (N_602,N_591,N_534);
nor U603 (N_603,N_586,N_549);
nand U604 (N_604,N_540,N_583);
nand U605 (N_605,N_544,N_564);
xor U606 (N_606,N_597,N_587);
nor U607 (N_607,N_565,N_547);
nor U608 (N_608,N_568,N_556);
or U609 (N_609,N_593,N_570);
nor U610 (N_610,N_563,N_557);
or U611 (N_611,N_538,N_580);
nand U612 (N_612,N_577,N_589);
nor U613 (N_613,N_584,N_574);
or U614 (N_614,N_541,N_537);
or U615 (N_615,N_588,N_559);
nand U616 (N_616,N_536,N_548);
and U617 (N_617,N_542,N_530);
or U618 (N_618,N_558,N_582);
xor U619 (N_619,N_529,N_553);
nor U620 (N_620,N_579,N_528);
and U621 (N_621,N_572,N_569);
xnor U622 (N_622,N_525,N_535);
or U623 (N_623,N_527,N_566);
and U624 (N_624,N_545,N_571);
nand U625 (N_625,N_594,N_560);
or U626 (N_626,N_552,N_555);
nor U627 (N_627,N_595,N_567);
and U628 (N_628,N_581,N_576);
xor U629 (N_629,N_575,N_551);
nor U630 (N_630,N_533,N_554);
xor U631 (N_631,N_596,N_590);
xor U632 (N_632,N_562,N_598);
and U633 (N_633,N_550,N_546);
and U634 (N_634,N_539,N_526);
nor U635 (N_635,N_531,N_592);
xnor U636 (N_636,N_532,N_599);
and U637 (N_637,N_585,N_563);
or U638 (N_638,N_534,N_599);
nand U639 (N_639,N_549,N_553);
or U640 (N_640,N_558,N_548);
or U641 (N_641,N_535,N_590);
and U642 (N_642,N_573,N_535);
and U643 (N_643,N_533,N_566);
and U644 (N_644,N_548,N_572);
xor U645 (N_645,N_563,N_583);
nand U646 (N_646,N_564,N_557);
nor U647 (N_647,N_531,N_565);
or U648 (N_648,N_541,N_549);
nor U649 (N_649,N_569,N_568);
nand U650 (N_650,N_529,N_568);
or U651 (N_651,N_588,N_529);
or U652 (N_652,N_531,N_552);
nor U653 (N_653,N_538,N_594);
and U654 (N_654,N_537,N_566);
and U655 (N_655,N_577,N_586);
nor U656 (N_656,N_562,N_534);
xor U657 (N_657,N_534,N_598);
nand U658 (N_658,N_532,N_556);
and U659 (N_659,N_555,N_533);
nor U660 (N_660,N_534,N_577);
nand U661 (N_661,N_555,N_586);
nand U662 (N_662,N_569,N_533);
xnor U663 (N_663,N_598,N_560);
nand U664 (N_664,N_561,N_568);
xnor U665 (N_665,N_577,N_549);
nor U666 (N_666,N_576,N_554);
nor U667 (N_667,N_536,N_555);
or U668 (N_668,N_548,N_564);
xnor U669 (N_669,N_573,N_591);
and U670 (N_670,N_557,N_560);
nor U671 (N_671,N_553,N_595);
xor U672 (N_672,N_589,N_568);
or U673 (N_673,N_539,N_562);
nand U674 (N_674,N_540,N_537);
xnor U675 (N_675,N_644,N_658);
nand U676 (N_676,N_619,N_612);
nand U677 (N_677,N_645,N_626);
and U678 (N_678,N_672,N_636);
nand U679 (N_679,N_641,N_615);
nor U680 (N_680,N_625,N_665);
nor U681 (N_681,N_621,N_662);
nand U682 (N_682,N_666,N_611);
xnor U683 (N_683,N_671,N_655);
nor U684 (N_684,N_617,N_667);
or U685 (N_685,N_670,N_635);
or U686 (N_686,N_620,N_642);
and U687 (N_687,N_648,N_606);
and U688 (N_688,N_634,N_650);
nor U689 (N_689,N_649,N_622);
nor U690 (N_690,N_654,N_628);
nor U691 (N_691,N_630,N_601);
nand U692 (N_692,N_613,N_652);
or U693 (N_693,N_656,N_614);
and U694 (N_694,N_623,N_638);
xnor U695 (N_695,N_661,N_674);
xor U696 (N_696,N_624,N_647);
xnor U697 (N_697,N_609,N_663);
and U698 (N_698,N_633,N_637);
xnor U699 (N_699,N_664,N_603);
xnor U700 (N_700,N_643,N_627);
or U701 (N_701,N_639,N_631);
xnor U702 (N_702,N_657,N_646);
and U703 (N_703,N_629,N_604);
nor U704 (N_704,N_659,N_653);
nor U705 (N_705,N_673,N_668);
or U706 (N_706,N_632,N_618);
or U707 (N_707,N_600,N_605);
nand U708 (N_708,N_660,N_669);
or U709 (N_709,N_651,N_607);
nand U710 (N_710,N_640,N_616);
xnor U711 (N_711,N_602,N_610);
and U712 (N_712,N_608,N_609);
nor U713 (N_713,N_624,N_618);
and U714 (N_714,N_640,N_659);
nand U715 (N_715,N_649,N_672);
nand U716 (N_716,N_655,N_605);
xor U717 (N_717,N_603,N_607);
or U718 (N_718,N_648,N_673);
nand U719 (N_719,N_657,N_618);
xnor U720 (N_720,N_600,N_632);
and U721 (N_721,N_652,N_671);
nor U722 (N_722,N_601,N_650);
and U723 (N_723,N_627,N_622);
or U724 (N_724,N_610,N_656);
and U725 (N_725,N_647,N_626);
nor U726 (N_726,N_655,N_649);
nand U727 (N_727,N_653,N_649);
and U728 (N_728,N_641,N_645);
nand U729 (N_729,N_624,N_607);
and U730 (N_730,N_672,N_609);
and U731 (N_731,N_631,N_625);
or U732 (N_732,N_660,N_659);
xnor U733 (N_733,N_608,N_670);
xor U734 (N_734,N_602,N_622);
and U735 (N_735,N_619,N_663);
xor U736 (N_736,N_653,N_612);
xnor U737 (N_737,N_648,N_653);
and U738 (N_738,N_608,N_618);
and U739 (N_739,N_621,N_633);
nor U740 (N_740,N_657,N_627);
xor U741 (N_741,N_625,N_658);
nand U742 (N_742,N_646,N_626);
nand U743 (N_743,N_631,N_642);
nor U744 (N_744,N_625,N_657);
xor U745 (N_745,N_655,N_654);
xor U746 (N_746,N_626,N_654);
xnor U747 (N_747,N_635,N_647);
nand U748 (N_748,N_614,N_637);
nor U749 (N_749,N_616,N_647);
nor U750 (N_750,N_685,N_689);
and U751 (N_751,N_683,N_749);
nor U752 (N_752,N_719,N_733);
or U753 (N_753,N_738,N_735);
xnor U754 (N_754,N_744,N_710);
or U755 (N_755,N_705,N_713);
and U756 (N_756,N_675,N_740);
or U757 (N_757,N_741,N_697);
and U758 (N_758,N_731,N_682);
xnor U759 (N_759,N_717,N_684);
and U760 (N_760,N_727,N_709);
nor U761 (N_761,N_721,N_677);
and U762 (N_762,N_678,N_732);
nand U763 (N_763,N_723,N_726);
or U764 (N_764,N_686,N_700);
nand U765 (N_765,N_688,N_745);
and U766 (N_766,N_747,N_711);
nor U767 (N_767,N_725,N_681);
and U768 (N_768,N_728,N_702);
nor U769 (N_769,N_720,N_692);
or U770 (N_770,N_724,N_715);
nand U771 (N_771,N_714,N_742);
or U772 (N_772,N_696,N_698);
or U773 (N_773,N_708,N_739);
and U774 (N_774,N_695,N_748);
or U775 (N_775,N_707,N_716);
or U776 (N_776,N_680,N_687);
or U777 (N_777,N_712,N_736);
xor U778 (N_778,N_703,N_679);
and U779 (N_779,N_734,N_690);
xor U780 (N_780,N_737,N_701);
nor U781 (N_781,N_676,N_722);
and U782 (N_782,N_743,N_704);
or U783 (N_783,N_729,N_694);
xnor U784 (N_784,N_699,N_746);
and U785 (N_785,N_691,N_706);
nor U786 (N_786,N_730,N_718);
or U787 (N_787,N_693,N_686);
xnor U788 (N_788,N_703,N_738);
nand U789 (N_789,N_688,N_679);
or U790 (N_790,N_718,N_678);
xnor U791 (N_791,N_725,N_687);
nor U792 (N_792,N_690,N_695);
nand U793 (N_793,N_715,N_701);
and U794 (N_794,N_725,N_728);
xor U795 (N_795,N_736,N_702);
and U796 (N_796,N_696,N_714);
nor U797 (N_797,N_740,N_677);
or U798 (N_798,N_687,N_706);
nor U799 (N_799,N_717,N_679);
and U800 (N_800,N_748,N_744);
nand U801 (N_801,N_738,N_709);
xor U802 (N_802,N_678,N_685);
and U803 (N_803,N_746,N_742);
nand U804 (N_804,N_713,N_709);
xor U805 (N_805,N_722,N_693);
nand U806 (N_806,N_749,N_737);
xnor U807 (N_807,N_711,N_745);
nor U808 (N_808,N_715,N_705);
nor U809 (N_809,N_741,N_747);
or U810 (N_810,N_693,N_719);
nor U811 (N_811,N_704,N_721);
and U812 (N_812,N_715,N_696);
nor U813 (N_813,N_714,N_738);
and U814 (N_814,N_707,N_738);
or U815 (N_815,N_737,N_675);
nand U816 (N_816,N_687,N_717);
xnor U817 (N_817,N_731,N_718);
or U818 (N_818,N_678,N_734);
and U819 (N_819,N_704,N_716);
nor U820 (N_820,N_721,N_720);
nand U821 (N_821,N_702,N_705);
nor U822 (N_822,N_748,N_749);
nor U823 (N_823,N_738,N_733);
nor U824 (N_824,N_705,N_723);
or U825 (N_825,N_760,N_761);
or U826 (N_826,N_822,N_792);
and U827 (N_827,N_755,N_811);
and U828 (N_828,N_753,N_776);
xor U829 (N_829,N_784,N_812);
or U830 (N_830,N_762,N_751);
and U831 (N_831,N_789,N_764);
nor U832 (N_832,N_782,N_759);
xnor U833 (N_833,N_806,N_758);
or U834 (N_834,N_799,N_818);
xnor U835 (N_835,N_791,N_815);
nor U836 (N_836,N_805,N_769);
xnor U837 (N_837,N_777,N_785);
and U838 (N_838,N_816,N_775);
nor U839 (N_839,N_824,N_795);
nand U840 (N_840,N_780,N_800);
nor U841 (N_841,N_754,N_798);
nor U842 (N_842,N_809,N_796);
and U843 (N_843,N_787,N_810);
or U844 (N_844,N_814,N_783);
nor U845 (N_845,N_803,N_763);
and U846 (N_846,N_765,N_821);
or U847 (N_847,N_808,N_804);
nor U848 (N_848,N_773,N_807);
nand U849 (N_849,N_786,N_823);
or U850 (N_850,N_757,N_768);
nor U851 (N_851,N_801,N_819);
xor U852 (N_852,N_756,N_790);
or U853 (N_853,N_770,N_817);
nand U854 (N_854,N_788,N_752);
or U855 (N_855,N_779,N_797);
and U856 (N_856,N_750,N_802);
or U857 (N_857,N_771,N_794);
xor U858 (N_858,N_772,N_778);
or U859 (N_859,N_774,N_820);
or U860 (N_860,N_766,N_813);
and U861 (N_861,N_781,N_793);
and U862 (N_862,N_767,N_818);
and U863 (N_863,N_777,N_779);
nand U864 (N_864,N_795,N_787);
nand U865 (N_865,N_790,N_755);
and U866 (N_866,N_822,N_802);
and U867 (N_867,N_763,N_755);
nor U868 (N_868,N_792,N_795);
and U869 (N_869,N_754,N_781);
xnor U870 (N_870,N_806,N_753);
or U871 (N_871,N_810,N_786);
and U872 (N_872,N_786,N_791);
or U873 (N_873,N_815,N_819);
or U874 (N_874,N_764,N_802);
nor U875 (N_875,N_779,N_773);
nand U876 (N_876,N_766,N_759);
and U877 (N_877,N_795,N_823);
or U878 (N_878,N_782,N_751);
nor U879 (N_879,N_803,N_774);
nand U880 (N_880,N_812,N_757);
nor U881 (N_881,N_800,N_763);
or U882 (N_882,N_755,N_791);
xnor U883 (N_883,N_821,N_782);
nor U884 (N_884,N_823,N_798);
nor U885 (N_885,N_785,N_751);
nand U886 (N_886,N_796,N_781);
xnor U887 (N_887,N_774,N_770);
nor U888 (N_888,N_820,N_754);
nor U889 (N_889,N_772,N_756);
nand U890 (N_890,N_770,N_810);
nor U891 (N_891,N_785,N_771);
and U892 (N_892,N_801,N_817);
nand U893 (N_893,N_789,N_819);
xor U894 (N_894,N_806,N_821);
and U895 (N_895,N_809,N_784);
nor U896 (N_896,N_811,N_760);
xnor U897 (N_897,N_820,N_805);
and U898 (N_898,N_768,N_758);
or U899 (N_899,N_772,N_786);
and U900 (N_900,N_830,N_856);
and U901 (N_901,N_867,N_832);
nor U902 (N_902,N_860,N_852);
nand U903 (N_903,N_836,N_854);
and U904 (N_904,N_898,N_894);
xor U905 (N_905,N_829,N_825);
or U906 (N_906,N_897,N_850);
nand U907 (N_907,N_877,N_881);
xnor U908 (N_908,N_853,N_861);
or U909 (N_909,N_866,N_875);
nand U910 (N_910,N_889,N_845);
nor U911 (N_911,N_882,N_833);
nand U912 (N_912,N_858,N_879);
or U913 (N_913,N_855,N_847);
nand U914 (N_914,N_884,N_887);
and U915 (N_915,N_828,N_865);
or U916 (N_916,N_834,N_859);
nor U917 (N_917,N_873,N_841);
nand U918 (N_918,N_840,N_844);
and U919 (N_919,N_863,N_885);
nand U920 (N_920,N_868,N_891);
or U921 (N_921,N_886,N_848);
xnor U922 (N_922,N_831,N_872);
nand U923 (N_923,N_862,N_837);
xor U924 (N_924,N_838,N_892);
xor U925 (N_925,N_899,N_827);
nand U926 (N_926,N_896,N_874);
or U927 (N_927,N_893,N_839);
or U928 (N_928,N_870,N_888);
or U929 (N_929,N_876,N_843);
and U930 (N_930,N_871,N_826);
and U931 (N_931,N_842,N_869);
xor U932 (N_932,N_895,N_883);
or U933 (N_933,N_878,N_880);
or U934 (N_934,N_857,N_851);
nor U935 (N_935,N_835,N_864);
or U936 (N_936,N_846,N_849);
xnor U937 (N_937,N_890,N_891);
xor U938 (N_938,N_849,N_896);
nand U939 (N_939,N_898,N_872);
or U940 (N_940,N_860,N_899);
nor U941 (N_941,N_866,N_872);
nor U942 (N_942,N_839,N_881);
or U943 (N_943,N_853,N_879);
nor U944 (N_944,N_849,N_873);
nor U945 (N_945,N_876,N_842);
or U946 (N_946,N_855,N_874);
and U947 (N_947,N_839,N_859);
nand U948 (N_948,N_885,N_856);
xnor U949 (N_949,N_854,N_884);
xnor U950 (N_950,N_838,N_857);
or U951 (N_951,N_885,N_887);
nand U952 (N_952,N_867,N_862);
and U953 (N_953,N_866,N_878);
nor U954 (N_954,N_875,N_874);
nand U955 (N_955,N_890,N_856);
xor U956 (N_956,N_830,N_828);
and U957 (N_957,N_887,N_865);
xnor U958 (N_958,N_831,N_867);
xnor U959 (N_959,N_836,N_844);
and U960 (N_960,N_852,N_829);
nor U961 (N_961,N_836,N_879);
xnor U962 (N_962,N_882,N_870);
nor U963 (N_963,N_885,N_849);
nor U964 (N_964,N_850,N_838);
xor U965 (N_965,N_859,N_844);
xor U966 (N_966,N_842,N_859);
nor U967 (N_967,N_858,N_895);
xor U968 (N_968,N_887,N_896);
xor U969 (N_969,N_889,N_850);
or U970 (N_970,N_891,N_888);
xor U971 (N_971,N_860,N_859);
nand U972 (N_972,N_878,N_890);
or U973 (N_973,N_870,N_853);
and U974 (N_974,N_833,N_855);
xor U975 (N_975,N_914,N_953);
xor U976 (N_976,N_928,N_945);
xnor U977 (N_977,N_970,N_921);
nor U978 (N_978,N_918,N_920);
and U979 (N_979,N_917,N_939);
or U980 (N_980,N_947,N_927);
xor U981 (N_981,N_956,N_904);
nand U982 (N_982,N_941,N_968);
xor U983 (N_983,N_926,N_930);
or U984 (N_984,N_922,N_929);
and U985 (N_985,N_907,N_958);
nand U986 (N_986,N_906,N_903);
or U987 (N_987,N_938,N_905);
nand U988 (N_988,N_960,N_901);
and U989 (N_989,N_965,N_932);
or U990 (N_990,N_944,N_915);
or U991 (N_991,N_925,N_940);
nand U992 (N_992,N_910,N_974);
or U993 (N_993,N_924,N_950);
nor U994 (N_994,N_942,N_959);
nand U995 (N_995,N_909,N_967);
xor U996 (N_996,N_951,N_972);
xor U997 (N_997,N_916,N_943);
nor U998 (N_998,N_955,N_946);
nor U999 (N_999,N_933,N_911);
or U1000 (N_1000,N_971,N_966);
nor U1001 (N_1001,N_919,N_935);
xor U1002 (N_1002,N_957,N_952);
xnor U1003 (N_1003,N_931,N_948);
nor U1004 (N_1004,N_961,N_937);
or U1005 (N_1005,N_954,N_936);
and U1006 (N_1006,N_923,N_962);
or U1007 (N_1007,N_969,N_913);
xor U1008 (N_1008,N_934,N_963);
xnor U1009 (N_1009,N_912,N_900);
nand U1010 (N_1010,N_964,N_902);
nand U1011 (N_1011,N_908,N_973);
xnor U1012 (N_1012,N_949,N_930);
nor U1013 (N_1013,N_955,N_945);
and U1014 (N_1014,N_970,N_936);
and U1015 (N_1015,N_950,N_939);
or U1016 (N_1016,N_909,N_950);
nand U1017 (N_1017,N_922,N_940);
nor U1018 (N_1018,N_972,N_921);
nor U1019 (N_1019,N_918,N_919);
nand U1020 (N_1020,N_974,N_912);
or U1021 (N_1021,N_957,N_954);
xnor U1022 (N_1022,N_921,N_957);
or U1023 (N_1023,N_919,N_927);
xor U1024 (N_1024,N_939,N_945);
and U1025 (N_1025,N_917,N_913);
and U1026 (N_1026,N_965,N_940);
nand U1027 (N_1027,N_902,N_939);
nand U1028 (N_1028,N_909,N_940);
and U1029 (N_1029,N_944,N_971);
or U1030 (N_1030,N_958,N_905);
or U1031 (N_1031,N_958,N_941);
nor U1032 (N_1032,N_972,N_932);
nand U1033 (N_1033,N_972,N_958);
or U1034 (N_1034,N_911,N_909);
xnor U1035 (N_1035,N_905,N_945);
nor U1036 (N_1036,N_924,N_947);
or U1037 (N_1037,N_924,N_945);
or U1038 (N_1038,N_904,N_963);
or U1039 (N_1039,N_944,N_917);
nand U1040 (N_1040,N_929,N_909);
or U1041 (N_1041,N_974,N_948);
nor U1042 (N_1042,N_960,N_957);
nand U1043 (N_1043,N_954,N_934);
and U1044 (N_1044,N_920,N_909);
nor U1045 (N_1045,N_968,N_918);
and U1046 (N_1046,N_948,N_967);
or U1047 (N_1047,N_964,N_916);
nor U1048 (N_1048,N_928,N_974);
or U1049 (N_1049,N_916,N_946);
xnor U1050 (N_1050,N_1021,N_1039);
or U1051 (N_1051,N_1018,N_1010);
nand U1052 (N_1052,N_981,N_1030);
nor U1053 (N_1053,N_1045,N_1008);
and U1054 (N_1054,N_1009,N_1014);
nor U1055 (N_1055,N_1028,N_1044);
and U1056 (N_1056,N_1013,N_992);
nand U1057 (N_1057,N_1016,N_994);
xnor U1058 (N_1058,N_1001,N_1042);
xor U1059 (N_1059,N_1049,N_978);
nor U1060 (N_1060,N_979,N_1047);
and U1061 (N_1061,N_1002,N_997);
xnor U1062 (N_1062,N_1015,N_1048);
xor U1063 (N_1063,N_986,N_1037);
nor U1064 (N_1064,N_1007,N_1012);
nor U1065 (N_1065,N_1036,N_1000);
xnor U1066 (N_1066,N_1040,N_1027);
xor U1067 (N_1067,N_1038,N_1019);
nand U1068 (N_1068,N_982,N_1017);
or U1069 (N_1069,N_1025,N_1024);
xor U1070 (N_1070,N_1005,N_993);
and U1071 (N_1071,N_995,N_989);
and U1072 (N_1072,N_991,N_980);
nor U1073 (N_1073,N_1004,N_1033);
nand U1074 (N_1074,N_1006,N_990);
or U1075 (N_1075,N_1035,N_1022);
nor U1076 (N_1076,N_984,N_1020);
or U1077 (N_1077,N_1026,N_988);
nor U1078 (N_1078,N_985,N_1032);
or U1079 (N_1079,N_996,N_1023);
and U1080 (N_1080,N_977,N_1041);
or U1081 (N_1081,N_983,N_1011);
xnor U1082 (N_1082,N_1043,N_1046);
and U1083 (N_1083,N_1029,N_1034);
nor U1084 (N_1084,N_975,N_1031);
or U1085 (N_1085,N_987,N_1003);
nor U1086 (N_1086,N_976,N_999);
nor U1087 (N_1087,N_998,N_979);
or U1088 (N_1088,N_1015,N_978);
nand U1089 (N_1089,N_1004,N_989);
nor U1090 (N_1090,N_993,N_1038);
xor U1091 (N_1091,N_998,N_980);
or U1092 (N_1092,N_985,N_986);
or U1093 (N_1093,N_1044,N_984);
and U1094 (N_1094,N_979,N_987);
and U1095 (N_1095,N_1022,N_1047);
nor U1096 (N_1096,N_978,N_983);
nand U1097 (N_1097,N_1009,N_975);
and U1098 (N_1098,N_1019,N_979);
or U1099 (N_1099,N_1048,N_1005);
nand U1100 (N_1100,N_1034,N_1009);
xor U1101 (N_1101,N_1015,N_1040);
nor U1102 (N_1102,N_1041,N_1031);
nand U1103 (N_1103,N_1018,N_997);
nor U1104 (N_1104,N_1023,N_1005);
or U1105 (N_1105,N_978,N_976);
or U1106 (N_1106,N_1035,N_1049);
nor U1107 (N_1107,N_1028,N_1018);
and U1108 (N_1108,N_1040,N_983);
nor U1109 (N_1109,N_1008,N_1041);
and U1110 (N_1110,N_1015,N_981);
nand U1111 (N_1111,N_1008,N_1007);
xor U1112 (N_1112,N_1026,N_1003);
or U1113 (N_1113,N_1018,N_999);
xor U1114 (N_1114,N_990,N_1029);
nor U1115 (N_1115,N_1021,N_1014);
or U1116 (N_1116,N_1006,N_1021);
nand U1117 (N_1117,N_1006,N_1027);
and U1118 (N_1118,N_1032,N_1036);
nor U1119 (N_1119,N_1018,N_1015);
nand U1120 (N_1120,N_989,N_1010);
or U1121 (N_1121,N_1019,N_1043);
or U1122 (N_1122,N_975,N_1000);
and U1123 (N_1123,N_1011,N_985);
nor U1124 (N_1124,N_1003,N_1046);
or U1125 (N_1125,N_1074,N_1088);
or U1126 (N_1126,N_1096,N_1122);
and U1127 (N_1127,N_1118,N_1110);
or U1128 (N_1128,N_1058,N_1090);
or U1129 (N_1129,N_1121,N_1123);
or U1130 (N_1130,N_1078,N_1069);
nand U1131 (N_1131,N_1097,N_1051);
or U1132 (N_1132,N_1102,N_1113);
xnor U1133 (N_1133,N_1063,N_1066);
or U1134 (N_1134,N_1100,N_1111);
and U1135 (N_1135,N_1072,N_1079);
and U1136 (N_1136,N_1085,N_1115);
or U1137 (N_1137,N_1095,N_1077);
or U1138 (N_1138,N_1089,N_1119);
nand U1139 (N_1139,N_1117,N_1065);
xor U1140 (N_1140,N_1124,N_1059);
or U1141 (N_1141,N_1086,N_1106);
xnor U1142 (N_1142,N_1101,N_1092);
nand U1143 (N_1143,N_1112,N_1104);
or U1144 (N_1144,N_1105,N_1091);
nand U1145 (N_1145,N_1070,N_1050);
nand U1146 (N_1146,N_1099,N_1055);
nor U1147 (N_1147,N_1068,N_1108);
xor U1148 (N_1148,N_1083,N_1109);
nand U1149 (N_1149,N_1080,N_1120);
xnor U1150 (N_1150,N_1084,N_1116);
xor U1151 (N_1151,N_1081,N_1053);
and U1152 (N_1152,N_1114,N_1103);
or U1153 (N_1153,N_1082,N_1057);
and U1154 (N_1154,N_1061,N_1052);
nor U1155 (N_1155,N_1087,N_1076);
nand U1156 (N_1156,N_1067,N_1075);
nand U1157 (N_1157,N_1062,N_1098);
and U1158 (N_1158,N_1060,N_1093);
and U1159 (N_1159,N_1056,N_1064);
and U1160 (N_1160,N_1071,N_1073);
xnor U1161 (N_1161,N_1094,N_1107);
nand U1162 (N_1162,N_1054,N_1085);
nor U1163 (N_1163,N_1115,N_1084);
xor U1164 (N_1164,N_1063,N_1091);
nand U1165 (N_1165,N_1075,N_1051);
nand U1166 (N_1166,N_1058,N_1098);
xor U1167 (N_1167,N_1117,N_1089);
xnor U1168 (N_1168,N_1087,N_1062);
and U1169 (N_1169,N_1097,N_1087);
nor U1170 (N_1170,N_1109,N_1077);
or U1171 (N_1171,N_1115,N_1056);
nand U1172 (N_1172,N_1054,N_1111);
nor U1173 (N_1173,N_1099,N_1074);
nor U1174 (N_1174,N_1067,N_1058);
or U1175 (N_1175,N_1090,N_1071);
and U1176 (N_1176,N_1106,N_1076);
xor U1177 (N_1177,N_1058,N_1077);
nand U1178 (N_1178,N_1058,N_1076);
nor U1179 (N_1179,N_1093,N_1112);
or U1180 (N_1180,N_1086,N_1097);
nor U1181 (N_1181,N_1080,N_1063);
nand U1182 (N_1182,N_1112,N_1120);
or U1183 (N_1183,N_1105,N_1123);
nand U1184 (N_1184,N_1065,N_1091);
and U1185 (N_1185,N_1074,N_1054);
nor U1186 (N_1186,N_1123,N_1069);
nand U1187 (N_1187,N_1124,N_1073);
xor U1188 (N_1188,N_1124,N_1063);
nand U1189 (N_1189,N_1050,N_1056);
xor U1190 (N_1190,N_1120,N_1078);
nand U1191 (N_1191,N_1093,N_1076);
nand U1192 (N_1192,N_1114,N_1098);
and U1193 (N_1193,N_1081,N_1075);
and U1194 (N_1194,N_1103,N_1073);
nor U1195 (N_1195,N_1089,N_1120);
xnor U1196 (N_1196,N_1109,N_1118);
and U1197 (N_1197,N_1085,N_1072);
xnor U1198 (N_1198,N_1054,N_1055);
xnor U1199 (N_1199,N_1115,N_1107);
nand U1200 (N_1200,N_1175,N_1155);
or U1201 (N_1201,N_1187,N_1190);
nand U1202 (N_1202,N_1189,N_1182);
and U1203 (N_1203,N_1154,N_1146);
xor U1204 (N_1204,N_1188,N_1173);
and U1205 (N_1205,N_1156,N_1153);
nand U1206 (N_1206,N_1135,N_1178);
or U1207 (N_1207,N_1134,N_1139);
xor U1208 (N_1208,N_1129,N_1198);
and U1209 (N_1209,N_1150,N_1165);
or U1210 (N_1210,N_1192,N_1147);
nand U1211 (N_1211,N_1195,N_1183);
or U1212 (N_1212,N_1161,N_1169);
or U1213 (N_1213,N_1136,N_1138);
nand U1214 (N_1214,N_1177,N_1171);
and U1215 (N_1215,N_1185,N_1149);
or U1216 (N_1216,N_1167,N_1151);
and U1217 (N_1217,N_1186,N_1143);
nor U1218 (N_1218,N_1191,N_1128);
nor U1219 (N_1219,N_1170,N_1125);
nor U1220 (N_1220,N_1132,N_1141);
nand U1221 (N_1221,N_1174,N_1162);
nand U1222 (N_1222,N_1157,N_1159);
nor U1223 (N_1223,N_1148,N_1194);
and U1224 (N_1224,N_1152,N_1180);
xor U1225 (N_1225,N_1179,N_1184);
and U1226 (N_1226,N_1140,N_1193);
nor U1227 (N_1227,N_1196,N_1199);
nor U1228 (N_1228,N_1145,N_1144);
nor U1229 (N_1229,N_1158,N_1164);
or U1230 (N_1230,N_1168,N_1197);
and U1231 (N_1231,N_1137,N_1166);
nor U1232 (N_1232,N_1130,N_1133);
or U1233 (N_1233,N_1126,N_1160);
nor U1234 (N_1234,N_1176,N_1172);
or U1235 (N_1235,N_1181,N_1163);
or U1236 (N_1236,N_1142,N_1131);
and U1237 (N_1237,N_1127,N_1163);
nor U1238 (N_1238,N_1185,N_1190);
nor U1239 (N_1239,N_1164,N_1125);
nor U1240 (N_1240,N_1175,N_1139);
nand U1241 (N_1241,N_1147,N_1129);
and U1242 (N_1242,N_1153,N_1157);
nor U1243 (N_1243,N_1170,N_1162);
and U1244 (N_1244,N_1160,N_1159);
nand U1245 (N_1245,N_1164,N_1193);
and U1246 (N_1246,N_1184,N_1164);
nor U1247 (N_1247,N_1145,N_1130);
nor U1248 (N_1248,N_1156,N_1151);
nor U1249 (N_1249,N_1129,N_1192);
nand U1250 (N_1250,N_1148,N_1151);
xnor U1251 (N_1251,N_1196,N_1127);
nand U1252 (N_1252,N_1162,N_1139);
nor U1253 (N_1253,N_1162,N_1129);
or U1254 (N_1254,N_1144,N_1152);
nor U1255 (N_1255,N_1181,N_1178);
nand U1256 (N_1256,N_1138,N_1132);
and U1257 (N_1257,N_1163,N_1189);
nor U1258 (N_1258,N_1180,N_1183);
and U1259 (N_1259,N_1167,N_1173);
xor U1260 (N_1260,N_1177,N_1145);
xor U1261 (N_1261,N_1190,N_1154);
nand U1262 (N_1262,N_1182,N_1143);
nand U1263 (N_1263,N_1126,N_1145);
nor U1264 (N_1264,N_1187,N_1146);
xor U1265 (N_1265,N_1186,N_1149);
xor U1266 (N_1266,N_1182,N_1186);
or U1267 (N_1267,N_1199,N_1190);
and U1268 (N_1268,N_1199,N_1163);
and U1269 (N_1269,N_1195,N_1160);
and U1270 (N_1270,N_1139,N_1199);
xnor U1271 (N_1271,N_1165,N_1192);
nand U1272 (N_1272,N_1170,N_1134);
nand U1273 (N_1273,N_1137,N_1146);
xnor U1274 (N_1274,N_1131,N_1129);
xnor U1275 (N_1275,N_1258,N_1248);
xnor U1276 (N_1276,N_1236,N_1219);
and U1277 (N_1277,N_1255,N_1237);
nor U1278 (N_1278,N_1214,N_1239);
nand U1279 (N_1279,N_1228,N_1229);
nand U1280 (N_1280,N_1262,N_1270);
xor U1281 (N_1281,N_1227,N_1225);
or U1282 (N_1282,N_1268,N_1200);
nand U1283 (N_1283,N_1218,N_1230);
xnor U1284 (N_1284,N_1211,N_1204);
nand U1285 (N_1285,N_1254,N_1234);
xnor U1286 (N_1286,N_1203,N_1201);
xor U1287 (N_1287,N_1244,N_1264);
nor U1288 (N_1288,N_1210,N_1231);
or U1289 (N_1289,N_1208,N_1261);
and U1290 (N_1290,N_1265,N_1246);
nand U1291 (N_1291,N_1256,N_1250);
nor U1292 (N_1292,N_1274,N_1216);
xor U1293 (N_1293,N_1252,N_1217);
or U1294 (N_1294,N_1226,N_1220);
or U1295 (N_1295,N_1207,N_1260);
or U1296 (N_1296,N_1202,N_1266);
or U1297 (N_1297,N_1232,N_1247);
nor U1298 (N_1298,N_1253,N_1263);
or U1299 (N_1299,N_1235,N_1249);
xnor U1300 (N_1300,N_1257,N_1213);
and U1301 (N_1301,N_1221,N_1272);
xor U1302 (N_1302,N_1233,N_1271);
nor U1303 (N_1303,N_1267,N_1243);
xnor U1304 (N_1304,N_1241,N_1212);
and U1305 (N_1305,N_1259,N_1269);
or U1306 (N_1306,N_1238,N_1223);
xnor U1307 (N_1307,N_1206,N_1222);
and U1308 (N_1308,N_1240,N_1251);
or U1309 (N_1309,N_1209,N_1215);
or U1310 (N_1310,N_1273,N_1205);
nor U1311 (N_1311,N_1224,N_1242);
or U1312 (N_1312,N_1245,N_1217);
xnor U1313 (N_1313,N_1244,N_1218);
nor U1314 (N_1314,N_1206,N_1233);
nand U1315 (N_1315,N_1201,N_1217);
nor U1316 (N_1316,N_1209,N_1244);
and U1317 (N_1317,N_1252,N_1268);
and U1318 (N_1318,N_1253,N_1234);
or U1319 (N_1319,N_1254,N_1264);
or U1320 (N_1320,N_1235,N_1236);
and U1321 (N_1321,N_1227,N_1258);
nor U1322 (N_1322,N_1265,N_1207);
or U1323 (N_1323,N_1265,N_1248);
nor U1324 (N_1324,N_1233,N_1227);
xor U1325 (N_1325,N_1233,N_1268);
and U1326 (N_1326,N_1229,N_1267);
xor U1327 (N_1327,N_1246,N_1241);
and U1328 (N_1328,N_1210,N_1214);
or U1329 (N_1329,N_1200,N_1212);
and U1330 (N_1330,N_1267,N_1261);
and U1331 (N_1331,N_1271,N_1260);
or U1332 (N_1332,N_1244,N_1205);
and U1333 (N_1333,N_1263,N_1247);
or U1334 (N_1334,N_1263,N_1272);
or U1335 (N_1335,N_1218,N_1270);
nand U1336 (N_1336,N_1227,N_1232);
nand U1337 (N_1337,N_1212,N_1267);
nand U1338 (N_1338,N_1247,N_1213);
and U1339 (N_1339,N_1201,N_1251);
nand U1340 (N_1340,N_1220,N_1210);
xor U1341 (N_1341,N_1266,N_1252);
xor U1342 (N_1342,N_1270,N_1255);
and U1343 (N_1343,N_1256,N_1243);
nand U1344 (N_1344,N_1264,N_1255);
nor U1345 (N_1345,N_1259,N_1218);
nor U1346 (N_1346,N_1272,N_1206);
nor U1347 (N_1347,N_1233,N_1226);
or U1348 (N_1348,N_1233,N_1232);
nor U1349 (N_1349,N_1248,N_1274);
xnor U1350 (N_1350,N_1326,N_1275);
xor U1351 (N_1351,N_1338,N_1343);
and U1352 (N_1352,N_1283,N_1325);
and U1353 (N_1353,N_1311,N_1292);
and U1354 (N_1354,N_1304,N_1286);
nand U1355 (N_1355,N_1293,N_1305);
or U1356 (N_1356,N_1333,N_1330);
or U1357 (N_1357,N_1277,N_1298);
xnor U1358 (N_1358,N_1300,N_1335);
and U1359 (N_1359,N_1297,N_1288);
nand U1360 (N_1360,N_1310,N_1282);
nor U1361 (N_1361,N_1322,N_1328);
nand U1362 (N_1362,N_1341,N_1306);
or U1363 (N_1363,N_1342,N_1315);
nand U1364 (N_1364,N_1294,N_1295);
and U1365 (N_1365,N_1321,N_1284);
or U1366 (N_1366,N_1278,N_1337);
nand U1367 (N_1367,N_1329,N_1279);
xnor U1368 (N_1368,N_1280,N_1302);
or U1369 (N_1369,N_1303,N_1345);
nor U1370 (N_1370,N_1301,N_1340);
nand U1371 (N_1371,N_1291,N_1320);
or U1372 (N_1372,N_1307,N_1289);
xnor U1373 (N_1373,N_1276,N_1332);
and U1374 (N_1374,N_1324,N_1313);
and U1375 (N_1375,N_1319,N_1334);
nor U1376 (N_1376,N_1348,N_1309);
nor U1377 (N_1377,N_1339,N_1327);
or U1378 (N_1378,N_1331,N_1349);
nand U1379 (N_1379,N_1312,N_1314);
and U1380 (N_1380,N_1323,N_1299);
or U1381 (N_1381,N_1346,N_1317);
nand U1382 (N_1382,N_1336,N_1308);
and U1383 (N_1383,N_1316,N_1281);
and U1384 (N_1384,N_1285,N_1287);
nand U1385 (N_1385,N_1347,N_1290);
and U1386 (N_1386,N_1296,N_1344);
nand U1387 (N_1387,N_1318,N_1296);
xor U1388 (N_1388,N_1313,N_1347);
and U1389 (N_1389,N_1319,N_1322);
or U1390 (N_1390,N_1285,N_1349);
nand U1391 (N_1391,N_1288,N_1287);
and U1392 (N_1392,N_1331,N_1347);
and U1393 (N_1393,N_1326,N_1342);
nand U1394 (N_1394,N_1321,N_1288);
and U1395 (N_1395,N_1300,N_1279);
nand U1396 (N_1396,N_1277,N_1328);
or U1397 (N_1397,N_1316,N_1341);
and U1398 (N_1398,N_1297,N_1275);
nor U1399 (N_1399,N_1303,N_1315);
nand U1400 (N_1400,N_1321,N_1319);
nand U1401 (N_1401,N_1316,N_1320);
xnor U1402 (N_1402,N_1324,N_1301);
nor U1403 (N_1403,N_1277,N_1339);
and U1404 (N_1404,N_1325,N_1299);
xnor U1405 (N_1405,N_1332,N_1279);
and U1406 (N_1406,N_1280,N_1331);
nand U1407 (N_1407,N_1331,N_1277);
and U1408 (N_1408,N_1344,N_1331);
nand U1409 (N_1409,N_1286,N_1311);
xnor U1410 (N_1410,N_1349,N_1290);
xnor U1411 (N_1411,N_1326,N_1286);
and U1412 (N_1412,N_1336,N_1292);
nand U1413 (N_1413,N_1326,N_1298);
and U1414 (N_1414,N_1346,N_1339);
nor U1415 (N_1415,N_1308,N_1330);
xor U1416 (N_1416,N_1319,N_1326);
nor U1417 (N_1417,N_1304,N_1324);
nor U1418 (N_1418,N_1345,N_1286);
or U1419 (N_1419,N_1336,N_1344);
and U1420 (N_1420,N_1320,N_1298);
or U1421 (N_1421,N_1339,N_1283);
xnor U1422 (N_1422,N_1322,N_1280);
nor U1423 (N_1423,N_1292,N_1317);
and U1424 (N_1424,N_1332,N_1286);
xnor U1425 (N_1425,N_1414,N_1357);
nor U1426 (N_1426,N_1420,N_1376);
nor U1427 (N_1427,N_1375,N_1393);
xor U1428 (N_1428,N_1421,N_1402);
nor U1429 (N_1429,N_1359,N_1404);
nand U1430 (N_1430,N_1391,N_1352);
nor U1431 (N_1431,N_1382,N_1356);
nand U1432 (N_1432,N_1423,N_1364);
or U1433 (N_1433,N_1384,N_1388);
xor U1434 (N_1434,N_1387,N_1371);
nor U1435 (N_1435,N_1383,N_1409);
xnor U1436 (N_1436,N_1385,N_1373);
xnor U1437 (N_1437,N_1401,N_1370);
nand U1438 (N_1438,N_1374,N_1407);
nor U1439 (N_1439,N_1406,N_1412);
and U1440 (N_1440,N_1367,N_1411);
xnor U1441 (N_1441,N_1405,N_1377);
xnor U1442 (N_1442,N_1397,N_1419);
and U1443 (N_1443,N_1368,N_1355);
nand U1444 (N_1444,N_1395,N_1369);
nor U1445 (N_1445,N_1410,N_1362);
and U1446 (N_1446,N_1390,N_1415);
and U1447 (N_1447,N_1408,N_1378);
xnor U1448 (N_1448,N_1379,N_1417);
xor U1449 (N_1449,N_1396,N_1389);
nor U1450 (N_1450,N_1351,N_1350);
or U1451 (N_1451,N_1424,N_1403);
xor U1452 (N_1452,N_1372,N_1358);
and U1453 (N_1453,N_1354,N_1386);
xnor U1454 (N_1454,N_1399,N_1363);
or U1455 (N_1455,N_1392,N_1400);
or U1456 (N_1456,N_1366,N_1418);
nor U1457 (N_1457,N_1381,N_1380);
nand U1458 (N_1458,N_1398,N_1413);
and U1459 (N_1459,N_1360,N_1422);
xnor U1460 (N_1460,N_1365,N_1394);
or U1461 (N_1461,N_1416,N_1353);
and U1462 (N_1462,N_1361,N_1420);
nor U1463 (N_1463,N_1372,N_1405);
xnor U1464 (N_1464,N_1369,N_1358);
or U1465 (N_1465,N_1418,N_1378);
or U1466 (N_1466,N_1382,N_1384);
nor U1467 (N_1467,N_1381,N_1370);
nand U1468 (N_1468,N_1370,N_1392);
xnor U1469 (N_1469,N_1354,N_1387);
or U1470 (N_1470,N_1358,N_1386);
xnor U1471 (N_1471,N_1375,N_1417);
or U1472 (N_1472,N_1382,N_1403);
nand U1473 (N_1473,N_1410,N_1370);
or U1474 (N_1474,N_1378,N_1401);
or U1475 (N_1475,N_1373,N_1353);
xnor U1476 (N_1476,N_1394,N_1375);
xnor U1477 (N_1477,N_1373,N_1406);
nand U1478 (N_1478,N_1374,N_1359);
xor U1479 (N_1479,N_1363,N_1365);
nor U1480 (N_1480,N_1413,N_1391);
nand U1481 (N_1481,N_1416,N_1422);
nand U1482 (N_1482,N_1354,N_1398);
and U1483 (N_1483,N_1379,N_1380);
nor U1484 (N_1484,N_1417,N_1364);
or U1485 (N_1485,N_1375,N_1411);
and U1486 (N_1486,N_1350,N_1382);
or U1487 (N_1487,N_1402,N_1419);
and U1488 (N_1488,N_1382,N_1360);
xnor U1489 (N_1489,N_1360,N_1418);
nand U1490 (N_1490,N_1419,N_1369);
and U1491 (N_1491,N_1407,N_1371);
nor U1492 (N_1492,N_1397,N_1363);
nor U1493 (N_1493,N_1424,N_1369);
xnor U1494 (N_1494,N_1417,N_1416);
xnor U1495 (N_1495,N_1356,N_1408);
nand U1496 (N_1496,N_1380,N_1421);
and U1497 (N_1497,N_1408,N_1350);
xor U1498 (N_1498,N_1382,N_1399);
nor U1499 (N_1499,N_1373,N_1354);
xor U1500 (N_1500,N_1429,N_1465);
or U1501 (N_1501,N_1438,N_1468);
and U1502 (N_1502,N_1442,N_1449);
or U1503 (N_1503,N_1466,N_1448);
nor U1504 (N_1504,N_1475,N_1499);
nand U1505 (N_1505,N_1444,N_1474);
nand U1506 (N_1506,N_1464,N_1472);
or U1507 (N_1507,N_1480,N_1446);
nor U1508 (N_1508,N_1498,N_1487);
or U1509 (N_1509,N_1436,N_1494);
nor U1510 (N_1510,N_1484,N_1452);
or U1511 (N_1511,N_1492,N_1447);
and U1512 (N_1512,N_1485,N_1454);
xnor U1513 (N_1513,N_1469,N_1431);
nand U1514 (N_1514,N_1482,N_1427);
and U1515 (N_1515,N_1489,N_1440);
nand U1516 (N_1516,N_1432,N_1483);
nand U1517 (N_1517,N_1434,N_1453);
xnor U1518 (N_1518,N_1425,N_1467);
nor U1519 (N_1519,N_1470,N_1481);
nor U1520 (N_1520,N_1456,N_1450);
xnor U1521 (N_1521,N_1497,N_1443);
or U1522 (N_1522,N_1439,N_1476);
or U1523 (N_1523,N_1441,N_1491);
nor U1524 (N_1524,N_1437,N_1457);
and U1525 (N_1525,N_1496,N_1435);
nor U1526 (N_1526,N_1477,N_1428);
or U1527 (N_1527,N_1479,N_1462);
nand U1528 (N_1528,N_1486,N_1430);
nor U1529 (N_1529,N_1460,N_1493);
nand U1530 (N_1530,N_1461,N_1426);
and U1531 (N_1531,N_1463,N_1433);
xnor U1532 (N_1532,N_1459,N_1458);
or U1533 (N_1533,N_1451,N_1455);
xnor U1534 (N_1534,N_1478,N_1471);
xnor U1535 (N_1535,N_1445,N_1495);
nor U1536 (N_1536,N_1490,N_1488);
and U1537 (N_1537,N_1473,N_1440);
nand U1538 (N_1538,N_1466,N_1434);
nand U1539 (N_1539,N_1463,N_1434);
or U1540 (N_1540,N_1481,N_1429);
and U1541 (N_1541,N_1473,N_1429);
nand U1542 (N_1542,N_1439,N_1478);
nand U1543 (N_1543,N_1465,N_1471);
nand U1544 (N_1544,N_1481,N_1425);
or U1545 (N_1545,N_1455,N_1487);
xor U1546 (N_1546,N_1498,N_1483);
xor U1547 (N_1547,N_1456,N_1493);
xnor U1548 (N_1548,N_1458,N_1470);
xnor U1549 (N_1549,N_1472,N_1490);
xnor U1550 (N_1550,N_1445,N_1448);
nand U1551 (N_1551,N_1454,N_1495);
or U1552 (N_1552,N_1473,N_1483);
and U1553 (N_1553,N_1481,N_1462);
and U1554 (N_1554,N_1450,N_1471);
xor U1555 (N_1555,N_1455,N_1498);
nor U1556 (N_1556,N_1435,N_1465);
xnor U1557 (N_1557,N_1475,N_1486);
and U1558 (N_1558,N_1463,N_1472);
nand U1559 (N_1559,N_1471,N_1499);
xnor U1560 (N_1560,N_1453,N_1450);
and U1561 (N_1561,N_1472,N_1452);
xor U1562 (N_1562,N_1441,N_1460);
nor U1563 (N_1563,N_1441,N_1446);
nor U1564 (N_1564,N_1475,N_1440);
xor U1565 (N_1565,N_1461,N_1462);
nor U1566 (N_1566,N_1462,N_1488);
nor U1567 (N_1567,N_1459,N_1444);
nor U1568 (N_1568,N_1426,N_1493);
xnor U1569 (N_1569,N_1459,N_1462);
xnor U1570 (N_1570,N_1477,N_1453);
xor U1571 (N_1571,N_1494,N_1493);
xor U1572 (N_1572,N_1485,N_1440);
or U1573 (N_1573,N_1442,N_1464);
nand U1574 (N_1574,N_1431,N_1476);
or U1575 (N_1575,N_1548,N_1533);
nor U1576 (N_1576,N_1563,N_1549);
xor U1577 (N_1577,N_1558,N_1532);
nor U1578 (N_1578,N_1570,N_1517);
nand U1579 (N_1579,N_1574,N_1528);
or U1580 (N_1580,N_1514,N_1553);
xnor U1581 (N_1581,N_1531,N_1510);
xor U1582 (N_1582,N_1568,N_1545);
or U1583 (N_1583,N_1527,N_1509);
xor U1584 (N_1584,N_1519,N_1542);
or U1585 (N_1585,N_1511,N_1551);
nor U1586 (N_1586,N_1518,N_1508);
nor U1587 (N_1587,N_1536,N_1515);
nor U1588 (N_1588,N_1572,N_1506);
and U1589 (N_1589,N_1559,N_1550);
nand U1590 (N_1590,N_1562,N_1513);
and U1591 (N_1591,N_1530,N_1525);
xor U1592 (N_1592,N_1537,N_1507);
xor U1593 (N_1593,N_1544,N_1500);
nor U1594 (N_1594,N_1566,N_1573);
nand U1595 (N_1595,N_1535,N_1556);
nor U1596 (N_1596,N_1529,N_1541);
and U1597 (N_1597,N_1539,N_1521);
xor U1598 (N_1598,N_1540,N_1526);
or U1599 (N_1599,N_1522,N_1557);
or U1600 (N_1600,N_1524,N_1552);
nor U1601 (N_1601,N_1546,N_1571);
xor U1602 (N_1602,N_1504,N_1520);
nor U1603 (N_1603,N_1569,N_1502);
nor U1604 (N_1604,N_1555,N_1543);
and U1605 (N_1605,N_1538,N_1565);
and U1606 (N_1606,N_1501,N_1547);
xnor U1607 (N_1607,N_1561,N_1512);
nor U1608 (N_1608,N_1560,N_1534);
and U1609 (N_1609,N_1564,N_1567);
xnor U1610 (N_1610,N_1554,N_1505);
or U1611 (N_1611,N_1516,N_1523);
xnor U1612 (N_1612,N_1503,N_1536);
xor U1613 (N_1613,N_1546,N_1547);
nor U1614 (N_1614,N_1548,N_1532);
nand U1615 (N_1615,N_1538,N_1563);
or U1616 (N_1616,N_1503,N_1510);
or U1617 (N_1617,N_1561,N_1546);
xor U1618 (N_1618,N_1557,N_1548);
or U1619 (N_1619,N_1521,N_1527);
and U1620 (N_1620,N_1562,N_1517);
nor U1621 (N_1621,N_1501,N_1518);
nor U1622 (N_1622,N_1543,N_1501);
nand U1623 (N_1623,N_1559,N_1545);
nand U1624 (N_1624,N_1547,N_1529);
nor U1625 (N_1625,N_1546,N_1573);
nor U1626 (N_1626,N_1525,N_1509);
xor U1627 (N_1627,N_1570,N_1573);
and U1628 (N_1628,N_1525,N_1519);
xor U1629 (N_1629,N_1554,N_1541);
and U1630 (N_1630,N_1505,N_1543);
or U1631 (N_1631,N_1508,N_1506);
and U1632 (N_1632,N_1562,N_1544);
nor U1633 (N_1633,N_1560,N_1566);
nand U1634 (N_1634,N_1523,N_1545);
nand U1635 (N_1635,N_1573,N_1515);
or U1636 (N_1636,N_1562,N_1520);
nand U1637 (N_1637,N_1561,N_1543);
xnor U1638 (N_1638,N_1544,N_1540);
or U1639 (N_1639,N_1537,N_1516);
or U1640 (N_1640,N_1502,N_1547);
xnor U1641 (N_1641,N_1534,N_1557);
nand U1642 (N_1642,N_1508,N_1503);
or U1643 (N_1643,N_1545,N_1525);
or U1644 (N_1644,N_1520,N_1555);
or U1645 (N_1645,N_1557,N_1502);
nor U1646 (N_1646,N_1512,N_1549);
nand U1647 (N_1647,N_1529,N_1566);
or U1648 (N_1648,N_1532,N_1513);
or U1649 (N_1649,N_1539,N_1518);
and U1650 (N_1650,N_1635,N_1631);
or U1651 (N_1651,N_1598,N_1614);
nor U1652 (N_1652,N_1584,N_1643);
xnor U1653 (N_1653,N_1596,N_1600);
nand U1654 (N_1654,N_1627,N_1576);
nand U1655 (N_1655,N_1593,N_1634);
xnor U1656 (N_1656,N_1620,N_1621);
or U1657 (N_1657,N_1647,N_1626);
or U1658 (N_1658,N_1586,N_1649);
nor U1659 (N_1659,N_1644,N_1613);
nand U1660 (N_1660,N_1630,N_1646);
nor U1661 (N_1661,N_1594,N_1622);
nand U1662 (N_1662,N_1633,N_1578);
nor U1663 (N_1663,N_1628,N_1616);
nand U1664 (N_1664,N_1624,N_1583);
nor U1665 (N_1665,N_1588,N_1629);
nand U1666 (N_1666,N_1605,N_1619);
nand U1667 (N_1667,N_1601,N_1625);
nand U1668 (N_1668,N_1607,N_1597);
nand U1669 (N_1669,N_1582,N_1580);
nand U1670 (N_1670,N_1589,N_1592);
and U1671 (N_1671,N_1608,N_1617);
nand U1672 (N_1672,N_1577,N_1637);
and U1673 (N_1673,N_1642,N_1590);
and U1674 (N_1674,N_1587,N_1606);
or U1675 (N_1675,N_1611,N_1615);
nor U1676 (N_1676,N_1640,N_1603);
nor U1677 (N_1677,N_1623,N_1610);
and U1678 (N_1678,N_1599,N_1595);
or U1679 (N_1679,N_1602,N_1632);
xnor U1680 (N_1680,N_1612,N_1579);
nor U1681 (N_1681,N_1604,N_1585);
xnor U1682 (N_1682,N_1641,N_1609);
nand U1683 (N_1683,N_1638,N_1618);
or U1684 (N_1684,N_1591,N_1636);
or U1685 (N_1685,N_1575,N_1645);
nor U1686 (N_1686,N_1648,N_1639);
xnor U1687 (N_1687,N_1581,N_1605);
nor U1688 (N_1688,N_1626,N_1640);
nor U1689 (N_1689,N_1623,N_1627);
and U1690 (N_1690,N_1627,N_1596);
nor U1691 (N_1691,N_1625,N_1623);
or U1692 (N_1692,N_1610,N_1577);
xor U1693 (N_1693,N_1622,N_1618);
nand U1694 (N_1694,N_1597,N_1625);
xnor U1695 (N_1695,N_1599,N_1597);
nor U1696 (N_1696,N_1584,N_1577);
nand U1697 (N_1697,N_1601,N_1622);
nor U1698 (N_1698,N_1645,N_1647);
nor U1699 (N_1699,N_1619,N_1648);
xor U1700 (N_1700,N_1638,N_1598);
xnor U1701 (N_1701,N_1589,N_1641);
or U1702 (N_1702,N_1629,N_1610);
nor U1703 (N_1703,N_1615,N_1635);
xnor U1704 (N_1704,N_1601,N_1594);
nand U1705 (N_1705,N_1603,N_1586);
and U1706 (N_1706,N_1646,N_1641);
nand U1707 (N_1707,N_1647,N_1633);
xnor U1708 (N_1708,N_1593,N_1622);
or U1709 (N_1709,N_1626,N_1646);
xnor U1710 (N_1710,N_1578,N_1597);
or U1711 (N_1711,N_1591,N_1647);
or U1712 (N_1712,N_1579,N_1609);
nor U1713 (N_1713,N_1577,N_1586);
nand U1714 (N_1714,N_1613,N_1641);
nor U1715 (N_1715,N_1640,N_1576);
or U1716 (N_1716,N_1598,N_1628);
xor U1717 (N_1717,N_1606,N_1634);
and U1718 (N_1718,N_1644,N_1588);
or U1719 (N_1719,N_1579,N_1582);
and U1720 (N_1720,N_1584,N_1616);
nor U1721 (N_1721,N_1644,N_1609);
or U1722 (N_1722,N_1649,N_1646);
nor U1723 (N_1723,N_1645,N_1632);
nand U1724 (N_1724,N_1612,N_1609);
xor U1725 (N_1725,N_1657,N_1695);
nand U1726 (N_1726,N_1680,N_1686);
and U1727 (N_1727,N_1684,N_1698);
xnor U1728 (N_1728,N_1663,N_1714);
xnor U1729 (N_1729,N_1717,N_1670);
nand U1730 (N_1730,N_1713,N_1671);
xor U1731 (N_1731,N_1652,N_1719);
nor U1732 (N_1732,N_1666,N_1668);
or U1733 (N_1733,N_1669,N_1706);
or U1734 (N_1734,N_1677,N_1707);
and U1735 (N_1735,N_1682,N_1672);
and U1736 (N_1736,N_1693,N_1712);
xor U1737 (N_1737,N_1715,N_1673);
nand U1738 (N_1738,N_1690,N_1667);
xnor U1739 (N_1739,N_1718,N_1724);
or U1740 (N_1740,N_1700,N_1709);
or U1741 (N_1741,N_1716,N_1662);
nand U1742 (N_1742,N_1651,N_1687);
and U1743 (N_1743,N_1650,N_1702);
or U1744 (N_1744,N_1692,N_1661);
nor U1745 (N_1745,N_1688,N_1659);
or U1746 (N_1746,N_1665,N_1655);
xnor U1747 (N_1747,N_1676,N_1678);
xor U1748 (N_1748,N_1683,N_1703);
or U1749 (N_1749,N_1691,N_1656);
nand U1750 (N_1750,N_1664,N_1704);
nand U1751 (N_1751,N_1694,N_1701);
and U1752 (N_1752,N_1658,N_1721);
nor U1753 (N_1753,N_1689,N_1711);
xnor U1754 (N_1754,N_1697,N_1720);
and U1755 (N_1755,N_1674,N_1679);
nand U1756 (N_1756,N_1722,N_1653);
and U1757 (N_1757,N_1710,N_1681);
nor U1758 (N_1758,N_1723,N_1699);
or U1759 (N_1759,N_1654,N_1708);
or U1760 (N_1760,N_1660,N_1675);
and U1761 (N_1761,N_1696,N_1705);
or U1762 (N_1762,N_1685,N_1709);
nand U1763 (N_1763,N_1665,N_1682);
and U1764 (N_1764,N_1659,N_1714);
and U1765 (N_1765,N_1706,N_1673);
xor U1766 (N_1766,N_1671,N_1710);
or U1767 (N_1767,N_1711,N_1690);
nor U1768 (N_1768,N_1654,N_1721);
or U1769 (N_1769,N_1654,N_1685);
or U1770 (N_1770,N_1699,N_1656);
xor U1771 (N_1771,N_1652,N_1701);
nand U1772 (N_1772,N_1695,N_1717);
or U1773 (N_1773,N_1723,N_1708);
or U1774 (N_1774,N_1708,N_1657);
xnor U1775 (N_1775,N_1662,N_1659);
nor U1776 (N_1776,N_1652,N_1718);
xor U1777 (N_1777,N_1702,N_1709);
or U1778 (N_1778,N_1707,N_1678);
nand U1779 (N_1779,N_1669,N_1690);
nand U1780 (N_1780,N_1689,N_1697);
or U1781 (N_1781,N_1718,N_1719);
xnor U1782 (N_1782,N_1686,N_1694);
nand U1783 (N_1783,N_1660,N_1724);
or U1784 (N_1784,N_1718,N_1654);
nand U1785 (N_1785,N_1677,N_1669);
xor U1786 (N_1786,N_1671,N_1662);
nor U1787 (N_1787,N_1653,N_1712);
or U1788 (N_1788,N_1652,N_1662);
nor U1789 (N_1789,N_1657,N_1655);
or U1790 (N_1790,N_1704,N_1650);
nand U1791 (N_1791,N_1697,N_1690);
xor U1792 (N_1792,N_1658,N_1689);
nor U1793 (N_1793,N_1702,N_1654);
and U1794 (N_1794,N_1707,N_1710);
nand U1795 (N_1795,N_1693,N_1671);
or U1796 (N_1796,N_1699,N_1696);
and U1797 (N_1797,N_1661,N_1703);
nand U1798 (N_1798,N_1683,N_1702);
and U1799 (N_1799,N_1724,N_1694);
nand U1800 (N_1800,N_1787,N_1751);
nor U1801 (N_1801,N_1789,N_1763);
or U1802 (N_1802,N_1798,N_1778);
or U1803 (N_1803,N_1737,N_1792);
xnor U1804 (N_1804,N_1777,N_1757);
nor U1805 (N_1805,N_1727,N_1775);
nor U1806 (N_1806,N_1740,N_1790);
and U1807 (N_1807,N_1748,N_1743);
and U1808 (N_1808,N_1794,N_1750);
nand U1809 (N_1809,N_1761,N_1739);
nand U1810 (N_1810,N_1797,N_1734);
nor U1811 (N_1811,N_1753,N_1744);
nand U1812 (N_1812,N_1793,N_1758);
or U1813 (N_1813,N_1731,N_1745);
nand U1814 (N_1814,N_1738,N_1772);
nand U1815 (N_1815,N_1741,N_1735);
nor U1816 (N_1816,N_1783,N_1780);
or U1817 (N_1817,N_1725,N_1776);
nand U1818 (N_1818,N_1733,N_1770);
nor U1819 (N_1819,N_1785,N_1768);
nor U1820 (N_1820,N_1764,N_1786);
nor U1821 (N_1821,N_1742,N_1781);
nor U1822 (N_1822,N_1728,N_1766);
xnor U1823 (N_1823,N_1730,N_1732);
nor U1824 (N_1824,N_1726,N_1749);
or U1825 (N_1825,N_1784,N_1769);
xnor U1826 (N_1826,N_1779,N_1796);
nand U1827 (N_1827,N_1754,N_1759);
nor U1828 (N_1828,N_1774,N_1795);
or U1829 (N_1829,N_1755,N_1736);
nand U1830 (N_1830,N_1799,N_1791);
xor U1831 (N_1831,N_1765,N_1729);
xor U1832 (N_1832,N_1773,N_1760);
nand U1833 (N_1833,N_1767,N_1746);
and U1834 (N_1834,N_1756,N_1752);
xor U1835 (N_1835,N_1762,N_1788);
xnor U1836 (N_1836,N_1771,N_1782);
and U1837 (N_1837,N_1747,N_1727);
and U1838 (N_1838,N_1731,N_1790);
nand U1839 (N_1839,N_1727,N_1766);
xnor U1840 (N_1840,N_1754,N_1789);
xnor U1841 (N_1841,N_1766,N_1798);
nand U1842 (N_1842,N_1745,N_1733);
nand U1843 (N_1843,N_1792,N_1777);
nand U1844 (N_1844,N_1791,N_1753);
nand U1845 (N_1845,N_1750,N_1725);
and U1846 (N_1846,N_1755,N_1738);
and U1847 (N_1847,N_1748,N_1793);
xor U1848 (N_1848,N_1733,N_1749);
xor U1849 (N_1849,N_1726,N_1759);
and U1850 (N_1850,N_1767,N_1749);
xor U1851 (N_1851,N_1761,N_1743);
xor U1852 (N_1852,N_1797,N_1759);
and U1853 (N_1853,N_1757,N_1734);
and U1854 (N_1854,N_1795,N_1744);
nor U1855 (N_1855,N_1786,N_1768);
or U1856 (N_1856,N_1793,N_1726);
nor U1857 (N_1857,N_1738,N_1771);
and U1858 (N_1858,N_1754,N_1795);
and U1859 (N_1859,N_1744,N_1764);
nor U1860 (N_1860,N_1788,N_1725);
or U1861 (N_1861,N_1764,N_1748);
nand U1862 (N_1862,N_1744,N_1789);
nor U1863 (N_1863,N_1768,N_1787);
nor U1864 (N_1864,N_1758,N_1784);
xor U1865 (N_1865,N_1764,N_1795);
xnor U1866 (N_1866,N_1785,N_1772);
and U1867 (N_1867,N_1773,N_1729);
and U1868 (N_1868,N_1743,N_1792);
nand U1869 (N_1869,N_1735,N_1796);
nand U1870 (N_1870,N_1736,N_1774);
nand U1871 (N_1871,N_1767,N_1762);
or U1872 (N_1872,N_1733,N_1776);
xor U1873 (N_1873,N_1791,N_1792);
xnor U1874 (N_1874,N_1759,N_1785);
and U1875 (N_1875,N_1858,N_1829);
xnor U1876 (N_1876,N_1860,N_1850);
xnor U1877 (N_1877,N_1833,N_1871);
nand U1878 (N_1878,N_1801,N_1810);
or U1879 (N_1879,N_1846,N_1865);
nand U1880 (N_1880,N_1814,N_1836);
and U1881 (N_1881,N_1843,N_1855);
and U1882 (N_1882,N_1842,N_1808);
xnor U1883 (N_1883,N_1873,N_1831);
or U1884 (N_1884,N_1867,N_1838);
xor U1885 (N_1885,N_1821,N_1849);
nand U1886 (N_1886,N_1813,N_1805);
and U1887 (N_1887,N_1863,N_1844);
xor U1888 (N_1888,N_1857,N_1806);
and U1889 (N_1889,N_1822,N_1807);
nand U1890 (N_1890,N_1839,N_1804);
nand U1891 (N_1891,N_1841,N_1866);
and U1892 (N_1892,N_1809,N_1802);
or U1893 (N_1893,N_1853,N_1874);
nand U1894 (N_1894,N_1816,N_1832);
xor U1895 (N_1895,N_1823,N_1826);
nand U1896 (N_1896,N_1869,N_1854);
or U1897 (N_1897,N_1872,N_1848);
xnor U1898 (N_1898,N_1800,N_1812);
xnor U1899 (N_1899,N_1862,N_1856);
nand U1900 (N_1900,N_1824,N_1837);
nor U1901 (N_1901,N_1861,N_1864);
xnor U1902 (N_1902,N_1859,N_1840);
or U1903 (N_1903,N_1825,N_1830);
or U1904 (N_1904,N_1851,N_1847);
and U1905 (N_1905,N_1815,N_1834);
or U1906 (N_1906,N_1827,N_1818);
xor U1907 (N_1907,N_1820,N_1819);
xnor U1908 (N_1908,N_1868,N_1811);
and U1909 (N_1909,N_1828,N_1803);
nand U1910 (N_1910,N_1845,N_1852);
or U1911 (N_1911,N_1817,N_1835);
and U1912 (N_1912,N_1870,N_1854);
nor U1913 (N_1913,N_1812,N_1835);
nand U1914 (N_1914,N_1847,N_1856);
and U1915 (N_1915,N_1863,N_1805);
and U1916 (N_1916,N_1844,N_1828);
and U1917 (N_1917,N_1808,N_1855);
or U1918 (N_1918,N_1861,N_1852);
and U1919 (N_1919,N_1809,N_1830);
and U1920 (N_1920,N_1816,N_1821);
nand U1921 (N_1921,N_1868,N_1832);
and U1922 (N_1922,N_1838,N_1868);
nor U1923 (N_1923,N_1845,N_1807);
nor U1924 (N_1924,N_1808,N_1844);
xnor U1925 (N_1925,N_1831,N_1861);
nand U1926 (N_1926,N_1850,N_1844);
and U1927 (N_1927,N_1865,N_1842);
or U1928 (N_1928,N_1833,N_1831);
and U1929 (N_1929,N_1845,N_1853);
nand U1930 (N_1930,N_1828,N_1864);
xor U1931 (N_1931,N_1853,N_1847);
nor U1932 (N_1932,N_1844,N_1820);
and U1933 (N_1933,N_1866,N_1873);
nor U1934 (N_1934,N_1812,N_1851);
nor U1935 (N_1935,N_1858,N_1802);
nand U1936 (N_1936,N_1831,N_1835);
xor U1937 (N_1937,N_1839,N_1802);
nor U1938 (N_1938,N_1858,N_1868);
or U1939 (N_1939,N_1856,N_1846);
or U1940 (N_1940,N_1824,N_1810);
and U1941 (N_1941,N_1800,N_1814);
nor U1942 (N_1942,N_1842,N_1812);
nor U1943 (N_1943,N_1832,N_1863);
and U1944 (N_1944,N_1832,N_1866);
xnor U1945 (N_1945,N_1816,N_1848);
and U1946 (N_1946,N_1811,N_1824);
xor U1947 (N_1947,N_1804,N_1850);
nand U1948 (N_1948,N_1873,N_1804);
nor U1949 (N_1949,N_1871,N_1824);
nor U1950 (N_1950,N_1899,N_1889);
xor U1951 (N_1951,N_1944,N_1922);
xor U1952 (N_1952,N_1923,N_1878);
nor U1953 (N_1953,N_1928,N_1925);
nor U1954 (N_1954,N_1941,N_1909);
or U1955 (N_1955,N_1883,N_1879);
or U1956 (N_1956,N_1919,N_1902);
and U1957 (N_1957,N_1932,N_1916);
and U1958 (N_1958,N_1890,N_1900);
and U1959 (N_1959,N_1891,N_1897);
nand U1960 (N_1960,N_1904,N_1882);
nand U1961 (N_1961,N_1888,N_1937);
nor U1962 (N_1962,N_1906,N_1905);
xor U1963 (N_1963,N_1915,N_1930);
xnor U1964 (N_1964,N_1877,N_1920);
xnor U1965 (N_1965,N_1896,N_1885);
or U1966 (N_1966,N_1945,N_1875);
and U1967 (N_1967,N_1907,N_1929);
and U1968 (N_1968,N_1876,N_1943);
nor U1969 (N_1969,N_1949,N_1946);
nor U1970 (N_1970,N_1917,N_1947);
and U1971 (N_1971,N_1939,N_1908);
nand U1972 (N_1972,N_1942,N_1881);
nor U1973 (N_1973,N_1936,N_1893);
nand U1974 (N_1974,N_1895,N_1912);
nand U1975 (N_1975,N_1910,N_1924);
and U1976 (N_1976,N_1886,N_1901);
xor U1977 (N_1977,N_1948,N_1918);
nand U1978 (N_1978,N_1940,N_1880);
nor U1979 (N_1979,N_1892,N_1921);
and U1980 (N_1980,N_1914,N_1903);
nand U1981 (N_1981,N_1913,N_1935);
xnor U1982 (N_1982,N_1926,N_1884);
nor U1983 (N_1983,N_1927,N_1934);
or U1984 (N_1984,N_1931,N_1933);
nand U1985 (N_1985,N_1938,N_1898);
and U1986 (N_1986,N_1894,N_1911);
or U1987 (N_1987,N_1887,N_1900);
and U1988 (N_1988,N_1899,N_1881);
nand U1989 (N_1989,N_1896,N_1914);
nor U1990 (N_1990,N_1949,N_1916);
and U1991 (N_1991,N_1929,N_1911);
nor U1992 (N_1992,N_1911,N_1884);
and U1993 (N_1993,N_1875,N_1878);
nor U1994 (N_1994,N_1940,N_1932);
nand U1995 (N_1995,N_1906,N_1926);
xnor U1996 (N_1996,N_1893,N_1894);
and U1997 (N_1997,N_1906,N_1943);
xor U1998 (N_1998,N_1914,N_1930);
nor U1999 (N_1999,N_1883,N_1940);
nand U2000 (N_2000,N_1901,N_1936);
nand U2001 (N_2001,N_1927,N_1888);
xor U2002 (N_2002,N_1916,N_1912);
and U2003 (N_2003,N_1889,N_1898);
nand U2004 (N_2004,N_1885,N_1942);
nand U2005 (N_2005,N_1944,N_1920);
xnor U2006 (N_2006,N_1947,N_1898);
or U2007 (N_2007,N_1940,N_1903);
xnor U2008 (N_2008,N_1887,N_1898);
nand U2009 (N_2009,N_1918,N_1906);
or U2010 (N_2010,N_1949,N_1889);
and U2011 (N_2011,N_1934,N_1936);
nand U2012 (N_2012,N_1905,N_1902);
and U2013 (N_2013,N_1908,N_1945);
nand U2014 (N_2014,N_1876,N_1933);
nand U2015 (N_2015,N_1878,N_1882);
xnor U2016 (N_2016,N_1941,N_1940);
or U2017 (N_2017,N_1924,N_1949);
nand U2018 (N_2018,N_1927,N_1947);
xor U2019 (N_2019,N_1894,N_1907);
or U2020 (N_2020,N_1918,N_1923);
nor U2021 (N_2021,N_1886,N_1883);
xnor U2022 (N_2022,N_1897,N_1942);
xor U2023 (N_2023,N_1907,N_1932);
nand U2024 (N_2024,N_1897,N_1945);
or U2025 (N_2025,N_2014,N_2023);
and U2026 (N_2026,N_1993,N_1990);
nand U2027 (N_2027,N_1962,N_1996);
xnor U2028 (N_2028,N_1986,N_2022);
or U2029 (N_2029,N_1952,N_1994);
nor U2030 (N_2030,N_1981,N_1964);
nand U2031 (N_2031,N_1997,N_1992);
and U2032 (N_2032,N_1960,N_1979);
nor U2033 (N_2033,N_2008,N_1951);
nand U2034 (N_2034,N_2020,N_2007);
and U2035 (N_2035,N_1984,N_2001);
xnor U2036 (N_2036,N_1968,N_2013);
xor U2037 (N_2037,N_1976,N_2019);
xnor U2038 (N_2038,N_1963,N_1989);
nand U2039 (N_2039,N_2024,N_2010);
xnor U2040 (N_2040,N_1957,N_2018);
xnor U2041 (N_2041,N_1959,N_1958);
xor U2042 (N_2042,N_2005,N_2009);
nor U2043 (N_2043,N_1980,N_2012);
xor U2044 (N_2044,N_1998,N_1985);
or U2045 (N_2045,N_1973,N_2003);
or U2046 (N_2046,N_2006,N_1961);
nor U2047 (N_2047,N_2017,N_1982);
nand U2048 (N_2048,N_2015,N_1965);
nand U2049 (N_2049,N_1988,N_1956);
nor U2050 (N_2050,N_1977,N_1971);
xnor U2051 (N_2051,N_1991,N_1978);
nand U2052 (N_2052,N_1983,N_1967);
or U2053 (N_2053,N_2000,N_2002);
or U2054 (N_2054,N_1970,N_1999);
xor U2055 (N_2055,N_1955,N_2021);
nand U2056 (N_2056,N_1950,N_2004);
and U2057 (N_2057,N_1969,N_1974);
nand U2058 (N_2058,N_2016,N_1966);
or U2059 (N_2059,N_1972,N_1975);
nor U2060 (N_2060,N_2011,N_1954);
or U2061 (N_2061,N_1987,N_1953);
nor U2062 (N_2062,N_1995,N_1969);
nand U2063 (N_2063,N_1962,N_1993);
or U2064 (N_2064,N_1983,N_1957);
or U2065 (N_2065,N_1999,N_2003);
or U2066 (N_2066,N_2012,N_1968);
nand U2067 (N_2067,N_2004,N_1966);
nor U2068 (N_2068,N_2020,N_1974);
or U2069 (N_2069,N_1981,N_2018);
xnor U2070 (N_2070,N_2022,N_1979);
nand U2071 (N_2071,N_1960,N_2020);
nand U2072 (N_2072,N_1974,N_1970);
xnor U2073 (N_2073,N_2007,N_1963);
xor U2074 (N_2074,N_1997,N_2019);
nand U2075 (N_2075,N_1986,N_1974);
nand U2076 (N_2076,N_1976,N_2004);
nand U2077 (N_2077,N_1979,N_1972);
xor U2078 (N_2078,N_2000,N_1962);
and U2079 (N_2079,N_1998,N_1959);
and U2080 (N_2080,N_1996,N_1986);
and U2081 (N_2081,N_1977,N_1975);
nor U2082 (N_2082,N_1980,N_1978);
xor U2083 (N_2083,N_1950,N_1984);
or U2084 (N_2084,N_1977,N_1965);
nor U2085 (N_2085,N_1959,N_1986);
or U2086 (N_2086,N_1989,N_2024);
nor U2087 (N_2087,N_1978,N_1957);
nor U2088 (N_2088,N_1985,N_2002);
nand U2089 (N_2089,N_1960,N_1982);
and U2090 (N_2090,N_1965,N_1976);
nor U2091 (N_2091,N_2019,N_1978);
xnor U2092 (N_2092,N_2024,N_1962);
or U2093 (N_2093,N_1994,N_1963);
nand U2094 (N_2094,N_1957,N_1952);
and U2095 (N_2095,N_1969,N_2002);
xor U2096 (N_2096,N_2019,N_1952);
and U2097 (N_2097,N_2008,N_2011);
and U2098 (N_2098,N_2009,N_1971);
or U2099 (N_2099,N_1981,N_1983);
nor U2100 (N_2100,N_2071,N_2030);
nand U2101 (N_2101,N_2051,N_2096);
or U2102 (N_2102,N_2099,N_2053);
xnor U2103 (N_2103,N_2081,N_2095);
and U2104 (N_2104,N_2078,N_2029);
nand U2105 (N_2105,N_2097,N_2027);
and U2106 (N_2106,N_2069,N_2025);
or U2107 (N_2107,N_2037,N_2082);
nand U2108 (N_2108,N_2085,N_2087);
and U2109 (N_2109,N_2094,N_2047);
nor U2110 (N_2110,N_2038,N_2072);
nor U2111 (N_2111,N_2068,N_2028);
nor U2112 (N_2112,N_2031,N_2083);
xor U2113 (N_2113,N_2035,N_2086);
and U2114 (N_2114,N_2057,N_2052);
and U2115 (N_2115,N_2064,N_2055);
nand U2116 (N_2116,N_2040,N_2026);
nand U2117 (N_2117,N_2032,N_2080);
nand U2118 (N_2118,N_2044,N_2059);
xor U2119 (N_2119,N_2084,N_2060);
and U2120 (N_2120,N_2089,N_2073);
and U2121 (N_2121,N_2043,N_2063);
nor U2122 (N_2122,N_2049,N_2046);
or U2123 (N_2123,N_2056,N_2061);
nand U2124 (N_2124,N_2054,N_2033);
nor U2125 (N_2125,N_2067,N_2045);
xnor U2126 (N_2126,N_2042,N_2077);
and U2127 (N_2127,N_2041,N_2065);
and U2128 (N_2128,N_2062,N_2074);
xor U2129 (N_2129,N_2088,N_2050);
nand U2130 (N_2130,N_2090,N_2034);
xnor U2131 (N_2131,N_2076,N_2092);
and U2132 (N_2132,N_2048,N_2091);
xor U2133 (N_2133,N_2070,N_2036);
nand U2134 (N_2134,N_2079,N_2098);
xnor U2135 (N_2135,N_2093,N_2058);
xnor U2136 (N_2136,N_2066,N_2075);
nor U2137 (N_2137,N_2039,N_2069);
nand U2138 (N_2138,N_2052,N_2038);
or U2139 (N_2139,N_2080,N_2062);
nor U2140 (N_2140,N_2057,N_2094);
nor U2141 (N_2141,N_2064,N_2088);
xnor U2142 (N_2142,N_2064,N_2092);
and U2143 (N_2143,N_2084,N_2092);
xnor U2144 (N_2144,N_2071,N_2046);
nand U2145 (N_2145,N_2084,N_2094);
xnor U2146 (N_2146,N_2090,N_2046);
nand U2147 (N_2147,N_2041,N_2051);
nor U2148 (N_2148,N_2060,N_2049);
or U2149 (N_2149,N_2060,N_2037);
xor U2150 (N_2150,N_2048,N_2096);
or U2151 (N_2151,N_2063,N_2091);
nor U2152 (N_2152,N_2058,N_2033);
nor U2153 (N_2153,N_2042,N_2039);
nand U2154 (N_2154,N_2089,N_2075);
and U2155 (N_2155,N_2050,N_2098);
and U2156 (N_2156,N_2090,N_2037);
or U2157 (N_2157,N_2043,N_2054);
nor U2158 (N_2158,N_2073,N_2067);
or U2159 (N_2159,N_2071,N_2039);
or U2160 (N_2160,N_2061,N_2034);
or U2161 (N_2161,N_2032,N_2057);
nor U2162 (N_2162,N_2062,N_2043);
or U2163 (N_2163,N_2053,N_2030);
nor U2164 (N_2164,N_2066,N_2041);
and U2165 (N_2165,N_2090,N_2026);
nor U2166 (N_2166,N_2040,N_2044);
nor U2167 (N_2167,N_2034,N_2048);
or U2168 (N_2168,N_2073,N_2079);
nor U2169 (N_2169,N_2091,N_2067);
nor U2170 (N_2170,N_2031,N_2036);
xnor U2171 (N_2171,N_2089,N_2093);
and U2172 (N_2172,N_2089,N_2085);
and U2173 (N_2173,N_2050,N_2047);
and U2174 (N_2174,N_2048,N_2049);
or U2175 (N_2175,N_2149,N_2143);
xor U2176 (N_2176,N_2162,N_2104);
or U2177 (N_2177,N_2113,N_2107);
nand U2178 (N_2178,N_2170,N_2125);
or U2179 (N_2179,N_2174,N_2127);
or U2180 (N_2180,N_2139,N_2126);
or U2181 (N_2181,N_2160,N_2101);
and U2182 (N_2182,N_2136,N_2103);
xor U2183 (N_2183,N_2150,N_2166);
xor U2184 (N_2184,N_2155,N_2128);
and U2185 (N_2185,N_2120,N_2114);
nor U2186 (N_2186,N_2124,N_2137);
nor U2187 (N_2187,N_2112,N_2133);
or U2188 (N_2188,N_2167,N_2157);
and U2189 (N_2189,N_2116,N_2152);
and U2190 (N_2190,N_2154,N_2148);
nand U2191 (N_2191,N_2161,N_2151);
nor U2192 (N_2192,N_2119,N_2122);
nand U2193 (N_2193,N_2158,N_2140);
xor U2194 (N_2194,N_2138,N_2169);
nand U2195 (N_2195,N_2134,N_2121);
nand U2196 (N_2196,N_2145,N_2135);
nor U2197 (N_2197,N_2168,N_2171);
nor U2198 (N_2198,N_2118,N_2159);
nand U2199 (N_2199,N_2111,N_2144);
xnor U2200 (N_2200,N_2117,N_2156);
xnor U2201 (N_2201,N_2129,N_2163);
or U2202 (N_2202,N_2108,N_2146);
nand U2203 (N_2203,N_2173,N_2109);
nand U2204 (N_2204,N_2110,N_2164);
and U2205 (N_2205,N_2141,N_2172);
xor U2206 (N_2206,N_2115,N_2131);
and U2207 (N_2207,N_2142,N_2130);
nor U2208 (N_2208,N_2102,N_2165);
or U2209 (N_2209,N_2106,N_2123);
nand U2210 (N_2210,N_2147,N_2132);
and U2211 (N_2211,N_2153,N_2100);
xnor U2212 (N_2212,N_2105,N_2174);
nand U2213 (N_2213,N_2117,N_2110);
nand U2214 (N_2214,N_2153,N_2131);
or U2215 (N_2215,N_2141,N_2164);
nand U2216 (N_2216,N_2164,N_2107);
xor U2217 (N_2217,N_2151,N_2165);
and U2218 (N_2218,N_2156,N_2148);
nor U2219 (N_2219,N_2100,N_2164);
nor U2220 (N_2220,N_2122,N_2105);
nor U2221 (N_2221,N_2103,N_2114);
and U2222 (N_2222,N_2108,N_2163);
and U2223 (N_2223,N_2137,N_2126);
nor U2224 (N_2224,N_2143,N_2121);
xnor U2225 (N_2225,N_2127,N_2113);
nand U2226 (N_2226,N_2151,N_2172);
nor U2227 (N_2227,N_2171,N_2137);
nand U2228 (N_2228,N_2109,N_2122);
and U2229 (N_2229,N_2121,N_2147);
or U2230 (N_2230,N_2167,N_2165);
nor U2231 (N_2231,N_2122,N_2150);
or U2232 (N_2232,N_2139,N_2127);
nor U2233 (N_2233,N_2127,N_2152);
xnor U2234 (N_2234,N_2155,N_2125);
and U2235 (N_2235,N_2148,N_2166);
xor U2236 (N_2236,N_2138,N_2112);
and U2237 (N_2237,N_2103,N_2165);
xor U2238 (N_2238,N_2156,N_2147);
nor U2239 (N_2239,N_2154,N_2126);
or U2240 (N_2240,N_2107,N_2152);
xnor U2241 (N_2241,N_2168,N_2147);
and U2242 (N_2242,N_2144,N_2123);
nor U2243 (N_2243,N_2130,N_2134);
and U2244 (N_2244,N_2173,N_2165);
nand U2245 (N_2245,N_2147,N_2113);
nor U2246 (N_2246,N_2109,N_2169);
nor U2247 (N_2247,N_2105,N_2141);
nand U2248 (N_2248,N_2114,N_2122);
and U2249 (N_2249,N_2108,N_2119);
nor U2250 (N_2250,N_2176,N_2227);
nor U2251 (N_2251,N_2241,N_2232);
xor U2252 (N_2252,N_2202,N_2247);
nor U2253 (N_2253,N_2183,N_2182);
nand U2254 (N_2254,N_2235,N_2203);
nor U2255 (N_2255,N_2223,N_2192);
or U2256 (N_2256,N_2220,N_2237);
nand U2257 (N_2257,N_2199,N_2204);
nor U2258 (N_2258,N_2217,N_2189);
xnor U2259 (N_2259,N_2224,N_2218);
nand U2260 (N_2260,N_2248,N_2181);
or U2261 (N_2261,N_2210,N_2234);
xor U2262 (N_2262,N_2242,N_2231);
or U2263 (N_2263,N_2221,N_2195);
xor U2264 (N_2264,N_2185,N_2191);
and U2265 (N_2265,N_2187,N_2238);
or U2266 (N_2266,N_2193,N_2215);
nor U2267 (N_2267,N_2179,N_2206);
nor U2268 (N_2268,N_2212,N_2236);
and U2269 (N_2269,N_2209,N_2226);
xor U2270 (N_2270,N_2225,N_2178);
and U2271 (N_2271,N_2239,N_2188);
and U2272 (N_2272,N_2208,N_2249);
or U2273 (N_2273,N_2184,N_2197);
nand U2274 (N_2274,N_2177,N_2200);
or U2275 (N_2275,N_2196,N_2245);
and U2276 (N_2276,N_2230,N_2211);
nor U2277 (N_2277,N_2180,N_2233);
or U2278 (N_2278,N_2243,N_2228);
nor U2279 (N_2279,N_2240,N_2194);
nor U2280 (N_2280,N_2216,N_2246);
and U2281 (N_2281,N_2201,N_2205);
or U2282 (N_2282,N_2214,N_2207);
nor U2283 (N_2283,N_2175,N_2186);
nor U2284 (N_2284,N_2190,N_2229);
xor U2285 (N_2285,N_2198,N_2219);
and U2286 (N_2286,N_2222,N_2244);
nand U2287 (N_2287,N_2213,N_2202);
and U2288 (N_2288,N_2235,N_2196);
nand U2289 (N_2289,N_2196,N_2190);
and U2290 (N_2290,N_2184,N_2244);
and U2291 (N_2291,N_2178,N_2245);
and U2292 (N_2292,N_2183,N_2207);
and U2293 (N_2293,N_2239,N_2225);
nand U2294 (N_2294,N_2181,N_2237);
nor U2295 (N_2295,N_2217,N_2233);
nor U2296 (N_2296,N_2194,N_2175);
nand U2297 (N_2297,N_2226,N_2199);
xor U2298 (N_2298,N_2178,N_2243);
nand U2299 (N_2299,N_2190,N_2185);
nand U2300 (N_2300,N_2198,N_2249);
nand U2301 (N_2301,N_2198,N_2234);
nand U2302 (N_2302,N_2231,N_2240);
or U2303 (N_2303,N_2244,N_2198);
nand U2304 (N_2304,N_2180,N_2177);
and U2305 (N_2305,N_2222,N_2185);
and U2306 (N_2306,N_2222,N_2217);
and U2307 (N_2307,N_2178,N_2199);
xnor U2308 (N_2308,N_2245,N_2205);
or U2309 (N_2309,N_2215,N_2208);
or U2310 (N_2310,N_2177,N_2212);
nand U2311 (N_2311,N_2226,N_2203);
or U2312 (N_2312,N_2185,N_2196);
xor U2313 (N_2313,N_2218,N_2206);
or U2314 (N_2314,N_2215,N_2198);
or U2315 (N_2315,N_2236,N_2182);
and U2316 (N_2316,N_2203,N_2225);
nor U2317 (N_2317,N_2195,N_2177);
or U2318 (N_2318,N_2183,N_2208);
nor U2319 (N_2319,N_2247,N_2175);
or U2320 (N_2320,N_2244,N_2179);
nor U2321 (N_2321,N_2202,N_2212);
xor U2322 (N_2322,N_2241,N_2231);
nor U2323 (N_2323,N_2235,N_2238);
nand U2324 (N_2324,N_2196,N_2188);
and U2325 (N_2325,N_2253,N_2261);
xnor U2326 (N_2326,N_2271,N_2267);
and U2327 (N_2327,N_2305,N_2318);
nand U2328 (N_2328,N_2292,N_2311);
nor U2329 (N_2329,N_2295,N_2279);
or U2330 (N_2330,N_2301,N_2255);
and U2331 (N_2331,N_2262,N_2323);
nor U2332 (N_2332,N_2317,N_2257);
and U2333 (N_2333,N_2312,N_2288);
xor U2334 (N_2334,N_2324,N_2307);
nand U2335 (N_2335,N_2313,N_2314);
xnor U2336 (N_2336,N_2287,N_2276);
or U2337 (N_2337,N_2254,N_2274);
xnor U2338 (N_2338,N_2315,N_2250);
or U2339 (N_2339,N_2283,N_2316);
or U2340 (N_2340,N_2281,N_2264);
and U2341 (N_2341,N_2258,N_2273);
and U2342 (N_2342,N_2310,N_2259);
nand U2343 (N_2343,N_2319,N_2263);
xnor U2344 (N_2344,N_2270,N_2282);
nand U2345 (N_2345,N_2252,N_2256);
xnor U2346 (N_2346,N_2251,N_2293);
and U2347 (N_2347,N_2304,N_2278);
or U2348 (N_2348,N_2309,N_2320);
or U2349 (N_2349,N_2306,N_2322);
nor U2350 (N_2350,N_2280,N_2266);
and U2351 (N_2351,N_2321,N_2289);
xor U2352 (N_2352,N_2290,N_2284);
or U2353 (N_2353,N_2286,N_2303);
or U2354 (N_2354,N_2298,N_2260);
or U2355 (N_2355,N_2308,N_2299);
xnor U2356 (N_2356,N_2285,N_2296);
or U2357 (N_2357,N_2269,N_2302);
nor U2358 (N_2358,N_2275,N_2277);
and U2359 (N_2359,N_2294,N_2291);
or U2360 (N_2360,N_2265,N_2268);
or U2361 (N_2361,N_2297,N_2300);
xor U2362 (N_2362,N_2272,N_2293);
nor U2363 (N_2363,N_2320,N_2257);
nand U2364 (N_2364,N_2281,N_2310);
and U2365 (N_2365,N_2314,N_2316);
and U2366 (N_2366,N_2262,N_2283);
nor U2367 (N_2367,N_2298,N_2294);
and U2368 (N_2368,N_2311,N_2262);
xnor U2369 (N_2369,N_2258,N_2306);
nand U2370 (N_2370,N_2266,N_2303);
nand U2371 (N_2371,N_2250,N_2300);
xor U2372 (N_2372,N_2273,N_2295);
nand U2373 (N_2373,N_2319,N_2253);
nand U2374 (N_2374,N_2260,N_2259);
nand U2375 (N_2375,N_2317,N_2260);
nor U2376 (N_2376,N_2256,N_2300);
nand U2377 (N_2377,N_2322,N_2268);
or U2378 (N_2378,N_2252,N_2281);
and U2379 (N_2379,N_2271,N_2283);
nand U2380 (N_2380,N_2319,N_2272);
nand U2381 (N_2381,N_2301,N_2298);
and U2382 (N_2382,N_2303,N_2301);
and U2383 (N_2383,N_2300,N_2265);
or U2384 (N_2384,N_2252,N_2270);
or U2385 (N_2385,N_2321,N_2315);
xor U2386 (N_2386,N_2324,N_2303);
or U2387 (N_2387,N_2284,N_2256);
xor U2388 (N_2388,N_2312,N_2285);
nor U2389 (N_2389,N_2284,N_2302);
nand U2390 (N_2390,N_2265,N_2324);
nand U2391 (N_2391,N_2304,N_2316);
or U2392 (N_2392,N_2322,N_2262);
and U2393 (N_2393,N_2299,N_2315);
nand U2394 (N_2394,N_2250,N_2307);
xor U2395 (N_2395,N_2250,N_2298);
or U2396 (N_2396,N_2253,N_2321);
and U2397 (N_2397,N_2256,N_2304);
nand U2398 (N_2398,N_2265,N_2292);
and U2399 (N_2399,N_2289,N_2261);
and U2400 (N_2400,N_2355,N_2365);
nor U2401 (N_2401,N_2335,N_2369);
xnor U2402 (N_2402,N_2397,N_2344);
xnor U2403 (N_2403,N_2342,N_2395);
xnor U2404 (N_2404,N_2398,N_2372);
nor U2405 (N_2405,N_2377,N_2332);
nor U2406 (N_2406,N_2384,N_2378);
nor U2407 (N_2407,N_2383,N_2396);
and U2408 (N_2408,N_2327,N_2340);
nand U2409 (N_2409,N_2390,N_2333);
nor U2410 (N_2410,N_2362,N_2366);
or U2411 (N_2411,N_2367,N_2371);
nand U2412 (N_2412,N_2331,N_2364);
and U2413 (N_2413,N_2393,N_2379);
xnor U2414 (N_2414,N_2357,N_2353);
or U2415 (N_2415,N_2345,N_2354);
nor U2416 (N_2416,N_2339,N_2389);
and U2417 (N_2417,N_2368,N_2386);
nand U2418 (N_2418,N_2326,N_2352);
and U2419 (N_2419,N_2328,N_2338);
or U2420 (N_2420,N_2336,N_2376);
xnor U2421 (N_2421,N_2346,N_2381);
nand U2422 (N_2422,N_2399,N_2382);
and U2423 (N_2423,N_2387,N_2348);
nor U2424 (N_2424,N_2388,N_2350);
or U2425 (N_2425,N_2374,N_2337);
and U2426 (N_2426,N_2341,N_2361);
and U2427 (N_2427,N_2370,N_2347);
or U2428 (N_2428,N_2385,N_2363);
and U2429 (N_2429,N_2392,N_2356);
xnor U2430 (N_2430,N_2330,N_2360);
and U2431 (N_2431,N_2329,N_2394);
or U2432 (N_2432,N_2359,N_2334);
and U2433 (N_2433,N_2391,N_2375);
nor U2434 (N_2434,N_2349,N_2351);
or U2435 (N_2435,N_2358,N_2343);
xor U2436 (N_2436,N_2380,N_2373);
and U2437 (N_2437,N_2325,N_2371);
xor U2438 (N_2438,N_2398,N_2378);
nand U2439 (N_2439,N_2395,N_2367);
xnor U2440 (N_2440,N_2349,N_2382);
xnor U2441 (N_2441,N_2390,N_2362);
nor U2442 (N_2442,N_2346,N_2340);
and U2443 (N_2443,N_2335,N_2355);
or U2444 (N_2444,N_2389,N_2349);
and U2445 (N_2445,N_2351,N_2390);
nand U2446 (N_2446,N_2378,N_2347);
or U2447 (N_2447,N_2365,N_2357);
nand U2448 (N_2448,N_2342,N_2327);
xnor U2449 (N_2449,N_2377,N_2329);
nor U2450 (N_2450,N_2380,N_2372);
xnor U2451 (N_2451,N_2326,N_2376);
and U2452 (N_2452,N_2374,N_2353);
and U2453 (N_2453,N_2346,N_2397);
nand U2454 (N_2454,N_2388,N_2383);
nand U2455 (N_2455,N_2360,N_2346);
or U2456 (N_2456,N_2357,N_2393);
xnor U2457 (N_2457,N_2369,N_2395);
nor U2458 (N_2458,N_2372,N_2341);
nand U2459 (N_2459,N_2331,N_2339);
nand U2460 (N_2460,N_2394,N_2352);
nor U2461 (N_2461,N_2352,N_2332);
or U2462 (N_2462,N_2398,N_2371);
or U2463 (N_2463,N_2399,N_2354);
nand U2464 (N_2464,N_2379,N_2345);
xor U2465 (N_2465,N_2377,N_2339);
xnor U2466 (N_2466,N_2398,N_2394);
nor U2467 (N_2467,N_2359,N_2368);
nand U2468 (N_2468,N_2338,N_2359);
or U2469 (N_2469,N_2343,N_2368);
nand U2470 (N_2470,N_2342,N_2382);
nand U2471 (N_2471,N_2328,N_2372);
nor U2472 (N_2472,N_2348,N_2358);
nand U2473 (N_2473,N_2357,N_2351);
or U2474 (N_2474,N_2365,N_2343);
and U2475 (N_2475,N_2440,N_2415);
xor U2476 (N_2476,N_2428,N_2469);
nand U2477 (N_2477,N_2412,N_2403);
nor U2478 (N_2478,N_2462,N_2472);
nand U2479 (N_2479,N_2427,N_2402);
nand U2480 (N_2480,N_2406,N_2441);
nor U2481 (N_2481,N_2445,N_2407);
xor U2482 (N_2482,N_2401,N_2444);
xnor U2483 (N_2483,N_2409,N_2465);
nor U2484 (N_2484,N_2416,N_2466);
and U2485 (N_2485,N_2405,N_2429);
or U2486 (N_2486,N_2458,N_2468);
nand U2487 (N_2487,N_2404,N_2437);
nand U2488 (N_2488,N_2408,N_2417);
nor U2489 (N_2489,N_2449,N_2450);
nand U2490 (N_2490,N_2433,N_2448);
and U2491 (N_2491,N_2459,N_2470);
nor U2492 (N_2492,N_2432,N_2424);
and U2493 (N_2493,N_2426,N_2463);
nor U2494 (N_2494,N_2410,N_2461);
nor U2495 (N_2495,N_2423,N_2414);
nor U2496 (N_2496,N_2454,N_2455);
nand U2497 (N_2497,N_2452,N_2447);
xor U2498 (N_2498,N_2439,N_2413);
or U2499 (N_2499,N_2436,N_2467);
nor U2500 (N_2500,N_2464,N_2421);
nor U2501 (N_2501,N_2418,N_2456);
or U2502 (N_2502,N_2434,N_2460);
nor U2503 (N_2503,N_2435,N_2451);
nor U2504 (N_2504,N_2431,N_2473);
xnor U2505 (N_2505,N_2425,N_2446);
nor U2506 (N_2506,N_2422,N_2430);
or U2507 (N_2507,N_2453,N_2443);
and U2508 (N_2508,N_2442,N_2419);
nand U2509 (N_2509,N_2457,N_2420);
nor U2510 (N_2510,N_2474,N_2471);
xnor U2511 (N_2511,N_2400,N_2438);
or U2512 (N_2512,N_2411,N_2410);
xnor U2513 (N_2513,N_2442,N_2421);
or U2514 (N_2514,N_2450,N_2438);
and U2515 (N_2515,N_2419,N_2412);
and U2516 (N_2516,N_2457,N_2439);
xor U2517 (N_2517,N_2424,N_2464);
or U2518 (N_2518,N_2465,N_2433);
nor U2519 (N_2519,N_2412,N_2418);
nor U2520 (N_2520,N_2415,N_2411);
or U2521 (N_2521,N_2436,N_2449);
nor U2522 (N_2522,N_2419,N_2409);
nor U2523 (N_2523,N_2414,N_2458);
or U2524 (N_2524,N_2444,N_2448);
nand U2525 (N_2525,N_2474,N_2437);
or U2526 (N_2526,N_2411,N_2463);
and U2527 (N_2527,N_2415,N_2417);
or U2528 (N_2528,N_2460,N_2468);
nor U2529 (N_2529,N_2447,N_2450);
nand U2530 (N_2530,N_2434,N_2436);
xor U2531 (N_2531,N_2464,N_2428);
nand U2532 (N_2532,N_2468,N_2403);
xnor U2533 (N_2533,N_2449,N_2460);
and U2534 (N_2534,N_2404,N_2416);
or U2535 (N_2535,N_2402,N_2434);
and U2536 (N_2536,N_2413,N_2436);
and U2537 (N_2537,N_2412,N_2442);
xnor U2538 (N_2538,N_2410,N_2455);
or U2539 (N_2539,N_2426,N_2410);
xnor U2540 (N_2540,N_2419,N_2469);
and U2541 (N_2541,N_2400,N_2435);
nand U2542 (N_2542,N_2459,N_2462);
nand U2543 (N_2543,N_2411,N_2447);
nor U2544 (N_2544,N_2460,N_2472);
and U2545 (N_2545,N_2426,N_2418);
xor U2546 (N_2546,N_2406,N_2438);
or U2547 (N_2547,N_2413,N_2442);
and U2548 (N_2548,N_2462,N_2425);
and U2549 (N_2549,N_2464,N_2439);
or U2550 (N_2550,N_2528,N_2527);
nor U2551 (N_2551,N_2513,N_2493);
nor U2552 (N_2552,N_2518,N_2495);
xnor U2553 (N_2553,N_2536,N_2492);
nor U2554 (N_2554,N_2515,N_2525);
nand U2555 (N_2555,N_2545,N_2486);
and U2556 (N_2556,N_2510,N_2544);
nand U2557 (N_2557,N_2478,N_2514);
nor U2558 (N_2558,N_2549,N_2508);
or U2559 (N_2559,N_2509,N_2479);
nor U2560 (N_2560,N_2497,N_2532);
nand U2561 (N_2561,N_2506,N_2489);
nor U2562 (N_2562,N_2543,N_2476);
or U2563 (N_2563,N_2477,N_2530);
xor U2564 (N_2564,N_2524,N_2542);
and U2565 (N_2565,N_2523,N_2526);
and U2566 (N_2566,N_2534,N_2539);
or U2567 (N_2567,N_2485,N_2487);
and U2568 (N_2568,N_2482,N_2507);
and U2569 (N_2569,N_2517,N_2546);
and U2570 (N_2570,N_2496,N_2538);
xnor U2571 (N_2571,N_2535,N_2522);
and U2572 (N_2572,N_2502,N_2537);
nor U2573 (N_2573,N_2480,N_2500);
and U2574 (N_2574,N_2520,N_2511);
xnor U2575 (N_2575,N_2505,N_2503);
and U2576 (N_2576,N_2491,N_2494);
nor U2577 (N_2577,N_2501,N_2481);
nand U2578 (N_2578,N_2531,N_2490);
or U2579 (N_2579,N_2512,N_2529);
nor U2580 (N_2580,N_2540,N_2488);
or U2581 (N_2581,N_2547,N_2504);
nand U2582 (N_2582,N_2541,N_2533);
xnor U2583 (N_2583,N_2498,N_2521);
and U2584 (N_2584,N_2483,N_2499);
xnor U2585 (N_2585,N_2519,N_2516);
nand U2586 (N_2586,N_2475,N_2548);
or U2587 (N_2587,N_2484,N_2534);
and U2588 (N_2588,N_2531,N_2536);
nor U2589 (N_2589,N_2492,N_2546);
and U2590 (N_2590,N_2523,N_2481);
or U2591 (N_2591,N_2531,N_2519);
nand U2592 (N_2592,N_2544,N_2518);
xor U2593 (N_2593,N_2527,N_2476);
nor U2594 (N_2594,N_2543,N_2477);
xnor U2595 (N_2595,N_2513,N_2516);
nand U2596 (N_2596,N_2527,N_2490);
or U2597 (N_2597,N_2527,N_2487);
or U2598 (N_2598,N_2521,N_2530);
and U2599 (N_2599,N_2544,N_2535);
nand U2600 (N_2600,N_2478,N_2512);
xor U2601 (N_2601,N_2482,N_2480);
xor U2602 (N_2602,N_2516,N_2545);
and U2603 (N_2603,N_2490,N_2521);
xnor U2604 (N_2604,N_2528,N_2549);
xor U2605 (N_2605,N_2520,N_2483);
nor U2606 (N_2606,N_2538,N_2548);
or U2607 (N_2607,N_2489,N_2528);
or U2608 (N_2608,N_2535,N_2537);
nor U2609 (N_2609,N_2480,N_2541);
xnor U2610 (N_2610,N_2500,N_2495);
nor U2611 (N_2611,N_2547,N_2535);
and U2612 (N_2612,N_2509,N_2529);
and U2613 (N_2613,N_2494,N_2539);
xor U2614 (N_2614,N_2503,N_2481);
or U2615 (N_2615,N_2546,N_2542);
xnor U2616 (N_2616,N_2475,N_2533);
or U2617 (N_2617,N_2527,N_2502);
xnor U2618 (N_2618,N_2543,N_2479);
nand U2619 (N_2619,N_2521,N_2549);
and U2620 (N_2620,N_2536,N_2475);
xor U2621 (N_2621,N_2511,N_2499);
or U2622 (N_2622,N_2483,N_2503);
and U2623 (N_2623,N_2489,N_2536);
xor U2624 (N_2624,N_2528,N_2536);
xnor U2625 (N_2625,N_2568,N_2583);
or U2626 (N_2626,N_2557,N_2552);
nor U2627 (N_2627,N_2598,N_2614);
and U2628 (N_2628,N_2564,N_2559);
xor U2629 (N_2629,N_2572,N_2602);
or U2630 (N_2630,N_2571,N_2594);
nand U2631 (N_2631,N_2605,N_2619);
and U2632 (N_2632,N_2609,N_2582);
xnor U2633 (N_2633,N_2587,N_2613);
nand U2634 (N_2634,N_2595,N_2560);
xnor U2635 (N_2635,N_2610,N_2577);
and U2636 (N_2636,N_2580,N_2578);
and U2637 (N_2637,N_2551,N_2563);
and U2638 (N_2638,N_2593,N_2561);
nor U2639 (N_2639,N_2620,N_2597);
or U2640 (N_2640,N_2622,N_2573);
nor U2641 (N_2641,N_2588,N_2608);
xnor U2642 (N_2642,N_2624,N_2565);
xor U2643 (N_2643,N_2621,N_2604);
nand U2644 (N_2644,N_2612,N_2584);
and U2645 (N_2645,N_2611,N_2556);
xnor U2646 (N_2646,N_2574,N_2615);
nand U2647 (N_2647,N_2569,N_2555);
nand U2648 (N_2648,N_2562,N_2567);
or U2649 (N_2649,N_2600,N_2599);
nor U2650 (N_2650,N_2566,N_2581);
nand U2651 (N_2651,N_2606,N_2601);
xor U2652 (N_2652,N_2586,N_2575);
nor U2653 (N_2653,N_2616,N_2607);
nor U2654 (N_2654,N_2590,N_2592);
and U2655 (N_2655,N_2579,N_2554);
nor U2656 (N_2656,N_2623,N_2576);
or U2657 (N_2657,N_2553,N_2589);
nand U2658 (N_2658,N_2550,N_2596);
xnor U2659 (N_2659,N_2558,N_2570);
or U2660 (N_2660,N_2618,N_2617);
nor U2661 (N_2661,N_2585,N_2591);
xor U2662 (N_2662,N_2603,N_2583);
nand U2663 (N_2663,N_2564,N_2572);
nand U2664 (N_2664,N_2607,N_2623);
xor U2665 (N_2665,N_2557,N_2619);
nand U2666 (N_2666,N_2579,N_2597);
and U2667 (N_2667,N_2579,N_2576);
xnor U2668 (N_2668,N_2613,N_2611);
nand U2669 (N_2669,N_2563,N_2624);
nand U2670 (N_2670,N_2612,N_2551);
nor U2671 (N_2671,N_2553,N_2602);
and U2672 (N_2672,N_2621,N_2554);
and U2673 (N_2673,N_2589,N_2563);
nand U2674 (N_2674,N_2593,N_2553);
and U2675 (N_2675,N_2573,N_2556);
xnor U2676 (N_2676,N_2554,N_2595);
or U2677 (N_2677,N_2576,N_2566);
or U2678 (N_2678,N_2551,N_2622);
nor U2679 (N_2679,N_2553,N_2597);
nor U2680 (N_2680,N_2590,N_2559);
xor U2681 (N_2681,N_2619,N_2592);
nor U2682 (N_2682,N_2607,N_2590);
nand U2683 (N_2683,N_2552,N_2612);
nor U2684 (N_2684,N_2580,N_2592);
and U2685 (N_2685,N_2620,N_2592);
xnor U2686 (N_2686,N_2553,N_2598);
nand U2687 (N_2687,N_2578,N_2551);
nor U2688 (N_2688,N_2619,N_2613);
xor U2689 (N_2689,N_2594,N_2579);
or U2690 (N_2690,N_2580,N_2576);
xnor U2691 (N_2691,N_2590,N_2620);
nand U2692 (N_2692,N_2586,N_2566);
xnor U2693 (N_2693,N_2584,N_2622);
xor U2694 (N_2694,N_2565,N_2597);
and U2695 (N_2695,N_2601,N_2571);
nand U2696 (N_2696,N_2623,N_2556);
and U2697 (N_2697,N_2571,N_2579);
or U2698 (N_2698,N_2563,N_2562);
nor U2699 (N_2699,N_2619,N_2622);
or U2700 (N_2700,N_2674,N_2649);
nor U2701 (N_2701,N_2656,N_2664);
and U2702 (N_2702,N_2690,N_2638);
nand U2703 (N_2703,N_2695,N_2644);
and U2704 (N_2704,N_2641,N_2680);
nor U2705 (N_2705,N_2698,N_2645);
and U2706 (N_2706,N_2679,N_2682);
or U2707 (N_2707,N_2689,N_2697);
or U2708 (N_2708,N_2667,N_2658);
or U2709 (N_2709,N_2655,N_2654);
or U2710 (N_2710,N_2643,N_2665);
or U2711 (N_2711,N_2684,N_2663);
xnor U2712 (N_2712,N_2669,N_2692);
xnor U2713 (N_2713,N_2632,N_2677);
xor U2714 (N_2714,N_2651,N_2659);
or U2715 (N_2715,N_2635,N_2666);
and U2716 (N_2716,N_2696,N_2660);
nor U2717 (N_2717,N_2691,N_2630);
xnor U2718 (N_2718,N_2676,N_2685);
or U2719 (N_2719,N_2650,N_2661);
xor U2720 (N_2720,N_2647,N_2683);
xnor U2721 (N_2721,N_2694,N_2672);
nor U2722 (N_2722,N_2626,N_2699);
or U2723 (N_2723,N_2688,N_2625);
or U2724 (N_2724,N_2671,N_2637);
or U2725 (N_2725,N_2662,N_2652);
or U2726 (N_2726,N_2687,N_2627);
and U2727 (N_2727,N_2675,N_2668);
nor U2728 (N_2728,N_2642,N_2686);
xor U2729 (N_2729,N_2633,N_2628);
xnor U2730 (N_2730,N_2629,N_2673);
nand U2731 (N_2731,N_2640,N_2636);
xor U2732 (N_2732,N_2648,N_2681);
or U2733 (N_2733,N_2653,N_2693);
xnor U2734 (N_2734,N_2634,N_2639);
xor U2735 (N_2735,N_2678,N_2646);
or U2736 (N_2736,N_2631,N_2670);
nand U2737 (N_2737,N_2657,N_2670);
nand U2738 (N_2738,N_2670,N_2688);
xor U2739 (N_2739,N_2662,N_2645);
nor U2740 (N_2740,N_2651,N_2647);
xnor U2741 (N_2741,N_2648,N_2626);
nor U2742 (N_2742,N_2652,N_2668);
and U2743 (N_2743,N_2633,N_2690);
or U2744 (N_2744,N_2641,N_2646);
xor U2745 (N_2745,N_2668,N_2634);
and U2746 (N_2746,N_2682,N_2634);
nor U2747 (N_2747,N_2678,N_2682);
nand U2748 (N_2748,N_2660,N_2651);
xnor U2749 (N_2749,N_2671,N_2698);
nor U2750 (N_2750,N_2660,N_2675);
or U2751 (N_2751,N_2647,N_2663);
and U2752 (N_2752,N_2633,N_2627);
nor U2753 (N_2753,N_2642,N_2631);
nor U2754 (N_2754,N_2692,N_2690);
nand U2755 (N_2755,N_2686,N_2629);
xor U2756 (N_2756,N_2676,N_2662);
and U2757 (N_2757,N_2659,N_2642);
nor U2758 (N_2758,N_2685,N_2686);
nand U2759 (N_2759,N_2665,N_2639);
nor U2760 (N_2760,N_2626,N_2625);
or U2761 (N_2761,N_2647,N_2684);
and U2762 (N_2762,N_2631,N_2626);
and U2763 (N_2763,N_2630,N_2670);
nor U2764 (N_2764,N_2654,N_2684);
xor U2765 (N_2765,N_2672,N_2679);
nor U2766 (N_2766,N_2649,N_2640);
or U2767 (N_2767,N_2693,N_2684);
and U2768 (N_2768,N_2652,N_2686);
or U2769 (N_2769,N_2645,N_2657);
and U2770 (N_2770,N_2675,N_2654);
nand U2771 (N_2771,N_2654,N_2669);
nand U2772 (N_2772,N_2686,N_2656);
nor U2773 (N_2773,N_2697,N_2666);
or U2774 (N_2774,N_2661,N_2665);
and U2775 (N_2775,N_2742,N_2712);
nand U2776 (N_2776,N_2714,N_2773);
or U2777 (N_2777,N_2727,N_2730);
and U2778 (N_2778,N_2719,N_2752);
nor U2779 (N_2779,N_2713,N_2743);
and U2780 (N_2780,N_2709,N_2729);
nor U2781 (N_2781,N_2753,N_2736);
or U2782 (N_2782,N_2750,N_2728);
or U2783 (N_2783,N_2759,N_2756);
or U2784 (N_2784,N_2744,N_2731);
or U2785 (N_2785,N_2774,N_2717);
or U2786 (N_2786,N_2772,N_2751);
nor U2787 (N_2787,N_2757,N_2765);
and U2788 (N_2788,N_2723,N_2741);
or U2789 (N_2789,N_2761,N_2734);
xor U2790 (N_2790,N_2739,N_2748);
or U2791 (N_2791,N_2725,N_2770);
xnor U2792 (N_2792,N_2746,N_2771);
nand U2793 (N_2793,N_2706,N_2705);
nor U2794 (N_2794,N_2720,N_2747);
nor U2795 (N_2795,N_2733,N_2763);
and U2796 (N_2796,N_2767,N_2754);
or U2797 (N_2797,N_2721,N_2769);
and U2798 (N_2798,N_2716,N_2708);
nor U2799 (N_2799,N_2738,N_2764);
xor U2800 (N_2800,N_2768,N_2718);
xor U2801 (N_2801,N_2737,N_2762);
nor U2802 (N_2802,N_2703,N_2711);
xnor U2803 (N_2803,N_2755,N_2726);
nand U2804 (N_2804,N_2704,N_2760);
or U2805 (N_2805,N_2710,N_2735);
nor U2806 (N_2806,N_2740,N_2701);
and U2807 (N_2807,N_2724,N_2715);
xnor U2808 (N_2808,N_2766,N_2732);
xor U2809 (N_2809,N_2707,N_2749);
and U2810 (N_2810,N_2758,N_2722);
or U2811 (N_2811,N_2702,N_2700);
and U2812 (N_2812,N_2745,N_2731);
and U2813 (N_2813,N_2718,N_2727);
nor U2814 (N_2814,N_2724,N_2764);
nor U2815 (N_2815,N_2762,N_2750);
nand U2816 (N_2816,N_2701,N_2738);
xnor U2817 (N_2817,N_2735,N_2738);
nor U2818 (N_2818,N_2754,N_2748);
and U2819 (N_2819,N_2766,N_2739);
xor U2820 (N_2820,N_2737,N_2723);
xnor U2821 (N_2821,N_2726,N_2700);
nand U2822 (N_2822,N_2741,N_2729);
xnor U2823 (N_2823,N_2750,N_2770);
nor U2824 (N_2824,N_2762,N_2758);
and U2825 (N_2825,N_2731,N_2729);
xnor U2826 (N_2826,N_2709,N_2730);
and U2827 (N_2827,N_2747,N_2763);
nand U2828 (N_2828,N_2768,N_2755);
xnor U2829 (N_2829,N_2734,N_2758);
and U2830 (N_2830,N_2735,N_2704);
or U2831 (N_2831,N_2711,N_2713);
and U2832 (N_2832,N_2732,N_2751);
xor U2833 (N_2833,N_2704,N_2734);
and U2834 (N_2834,N_2745,N_2761);
nand U2835 (N_2835,N_2705,N_2733);
nor U2836 (N_2836,N_2732,N_2721);
and U2837 (N_2837,N_2762,N_2735);
or U2838 (N_2838,N_2755,N_2731);
or U2839 (N_2839,N_2750,N_2712);
or U2840 (N_2840,N_2706,N_2774);
nand U2841 (N_2841,N_2739,N_2722);
xnor U2842 (N_2842,N_2770,N_2751);
xor U2843 (N_2843,N_2711,N_2735);
and U2844 (N_2844,N_2763,N_2719);
nor U2845 (N_2845,N_2751,N_2762);
nor U2846 (N_2846,N_2709,N_2763);
and U2847 (N_2847,N_2711,N_2756);
nor U2848 (N_2848,N_2736,N_2738);
nand U2849 (N_2849,N_2743,N_2761);
and U2850 (N_2850,N_2848,N_2844);
xnor U2851 (N_2851,N_2819,N_2800);
nand U2852 (N_2852,N_2789,N_2793);
and U2853 (N_2853,N_2808,N_2825);
nand U2854 (N_2854,N_2802,N_2834);
xor U2855 (N_2855,N_2784,N_2846);
nand U2856 (N_2856,N_2780,N_2847);
or U2857 (N_2857,N_2810,N_2826);
nand U2858 (N_2858,N_2842,N_2790);
or U2859 (N_2859,N_2816,N_2836);
nor U2860 (N_2860,N_2783,N_2849);
nor U2861 (N_2861,N_2817,N_2794);
nor U2862 (N_2862,N_2832,N_2839);
nor U2863 (N_2863,N_2797,N_2776);
and U2864 (N_2864,N_2812,N_2779);
and U2865 (N_2865,N_2804,N_2803);
or U2866 (N_2866,N_2830,N_2796);
and U2867 (N_2867,N_2811,N_2809);
nor U2868 (N_2868,N_2824,N_2791);
and U2869 (N_2869,N_2795,N_2781);
xnor U2870 (N_2870,N_2840,N_2823);
xor U2871 (N_2871,N_2843,N_2805);
and U2872 (N_2872,N_2806,N_2833);
or U2873 (N_2873,N_2828,N_2807);
nand U2874 (N_2874,N_2831,N_2821);
or U2875 (N_2875,N_2814,N_2788);
xor U2876 (N_2876,N_2815,N_2782);
nor U2877 (N_2877,N_2775,N_2829);
or U2878 (N_2878,N_2822,N_2799);
nor U2879 (N_2879,N_2798,N_2792);
nor U2880 (N_2880,N_2818,N_2786);
xor U2881 (N_2881,N_2820,N_2837);
or U2882 (N_2882,N_2838,N_2785);
xor U2883 (N_2883,N_2778,N_2827);
or U2884 (N_2884,N_2841,N_2787);
nand U2885 (N_2885,N_2835,N_2801);
or U2886 (N_2886,N_2845,N_2813);
xnor U2887 (N_2887,N_2777,N_2808);
nor U2888 (N_2888,N_2807,N_2810);
or U2889 (N_2889,N_2813,N_2775);
nor U2890 (N_2890,N_2836,N_2832);
and U2891 (N_2891,N_2782,N_2836);
nand U2892 (N_2892,N_2801,N_2782);
or U2893 (N_2893,N_2781,N_2837);
nand U2894 (N_2894,N_2835,N_2800);
xnor U2895 (N_2895,N_2807,N_2808);
or U2896 (N_2896,N_2845,N_2795);
nor U2897 (N_2897,N_2820,N_2827);
or U2898 (N_2898,N_2833,N_2837);
xnor U2899 (N_2899,N_2830,N_2831);
and U2900 (N_2900,N_2806,N_2779);
or U2901 (N_2901,N_2807,N_2846);
xnor U2902 (N_2902,N_2810,N_2832);
and U2903 (N_2903,N_2837,N_2818);
nor U2904 (N_2904,N_2849,N_2820);
nor U2905 (N_2905,N_2802,N_2821);
and U2906 (N_2906,N_2783,N_2845);
nand U2907 (N_2907,N_2826,N_2780);
xor U2908 (N_2908,N_2831,N_2790);
nor U2909 (N_2909,N_2818,N_2844);
nor U2910 (N_2910,N_2794,N_2815);
xnor U2911 (N_2911,N_2846,N_2840);
nand U2912 (N_2912,N_2797,N_2793);
or U2913 (N_2913,N_2838,N_2815);
or U2914 (N_2914,N_2792,N_2781);
xnor U2915 (N_2915,N_2823,N_2780);
nor U2916 (N_2916,N_2788,N_2784);
nand U2917 (N_2917,N_2811,N_2795);
nor U2918 (N_2918,N_2779,N_2832);
or U2919 (N_2919,N_2828,N_2803);
xor U2920 (N_2920,N_2828,N_2849);
xnor U2921 (N_2921,N_2814,N_2849);
nand U2922 (N_2922,N_2775,N_2796);
or U2923 (N_2923,N_2801,N_2824);
nor U2924 (N_2924,N_2776,N_2820);
nand U2925 (N_2925,N_2900,N_2881);
xnor U2926 (N_2926,N_2909,N_2910);
and U2927 (N_2927,N_2878,N_2911);
and U2928 (N_2928,N_2860,N_2863);
xnor U2929 (N_2929,N_2893,N_2866);
xnor U2930 (N_2930,N_2886,N_2869);
nor U2931 (N_2931,N_2907,N_2915);
nor U2932 (N_2932,N_2875,N_2885);
or U2933 (N_2933,N_2872,N_2922);
and U2934 (N_2934,N_2865,N_2917);
xor U2935 (N_2935,N_2914,N_2884);
and U2936 (N_2936,N_2851,N_2924);
nand U2937 (N_2937,N_2853,N_2916);
or U2938 (N_2938,N_2888,N_2880);
nand U2939 (N_2939,N_2904,N_2858);
nand U2940 (N_2940,N_2918,N_2857);
or U2941 (N_2941,N_2891,N_2852);
nor U2942 (N_2942,N_2890,N_2864);
xor U2943 (N_2943,N_2855,N_2882);
nor U2944 (N_2944,N_2873,N_2870);
and U2945 (N_2945,N_2902,N_2901);
nor U2946 (N_2946,N_2896,N_2897);
or U2947 (N_2947,N_2894,N_2854);
and U2948 (N_2948,N_2887,N_2895);
nor U2949 (N_2949,N_2913,N_2859);
nor U2950 (N_2950,N_2921,N_2908);
xor U2951 (N_2951,N_2850,N_2903);
or U2952 (N_2952,N_2899,N_2867);
nand U2953 (N_2953,N_2862,N_2898);
nand U2954 (N_2954,N_2877,N_2892);
and U2955 (N_2955,N_2920,N_2905);
nor U2956 (N_2956,N_2919,N_2856);
or U2957 (N_2957,N_2889,N_2879);
nor U2958 (N_2958,N_2861,N_2868);
xnor U2959 (N_2959,N_2906,N_2871);
nor U2960 (N_2960,N_2923,N_2876);
and U2961 (N_2961,N_2874,N_2912);
and U2962 (N_2962,N_2883,N_2913);
and U2963 (N_2963,N_2905,N_2862);
xor U2964 (N_2964,N_2894,N_2866);
or U2965 (N_2965,N_2867,N_2892);
xnor U2966 (N_2966,N_2901,N_2858);
xnor U2967 (N_2967,N_2920,N_2855);
or U2968 (N_2968,N_2852,N_2897);
nand U2969 (N_2969,N_2859,N_2914);
xnor U2970 (N_2970,N_2890,N_2900);
xor U2971 (N_2971,N_2863,N_2924);
or U2972 (N_2972,N_2904,N_2852);
and U2973 (N_2973,N_2890,N_2873);
and U2974 (N_2974,N_2898,N_2872);
nor U2975 (N_2975,N_2889,N_2861);
nor U2976 (N_2976,N_2909,N_2864);
nor U2977 (N_2977,N_2920,N_2878);
nand U2978 (N_2978,N_2890,N_2868);
and U2979 (N_2979,N_2912,N_2894);
nand U2980 (N_2980,N_2855,N_2923);
nor U2981 (N_2981,N_2921,N_2889);
and U2982 (N_2982,N_2872,N_2879);
and U2983 (N_2983,N_2860,N_2855);
or U2984 (N_2984,N_2893,N_2916);
or U2985 (N_2985,N_2873,N_2911);
and U2986 (N_2986,N_2864,N_2873);
xor U2987 (N_2987,N_2884,N_2923);
and U2988 (N_2988,N_2887,N_2866);
or U2989 (N_2989,N_2916,N_2896);
and U2990 (N_2990,N_2883,N_2879);
or U2991 (N_2991,N_2852,N_2869);
and U2992 (N_2992,N_2895,N_2911);
nor U2993 (N_2993,N_2879,N_2914);
nor U2994 (N_2994,N_2881,N_2897);
and U2995 (N_2995,N_2871,N_2872);
nor U2996 (N_2996,N_2904,N_2868);
and U2997 (N_2997,N_2896,N_2909);
nor U2998 (N_2998,N_2921,N_2858);
xor U2999 (N_2999,N_2919,N_2898);
xor UO_0 (O_0,N_2961,N_2999);
nand UO_1 (O_1,N_2990,N_2975);
and UO_2 (O_2,N_2988,N_2942);
xor UO_3 (O_3,N_2976,N_2943);
and UO_4 (O_4,N_2957,N_2955);
nand UO_5 (O_5,N_2974,N_2964);
nand UO_6 (O_6,N_2987,N_2989);
or UO_7 (O_7,N_2926,N_2968);
nor UO_8 (O_8,N_2962,N_2929);
nand UO_9 (O_9,N_2956,N_2945);
nor UO_10 (O_10,N_2972,N_2951);
nand UO_11 (O_11,N_2946,N_2969);
nand UO_12 (O_12,N_2941,N_2973);
nor UO_13 (O_13,N_2934,N_2939);
nor UO_14 (O_14,N_2992,N_2959);
and UO_15 (O_15,N_2938,N_2935);
nor UO_16 (O_16,N_2940,N_2978);
and UO_17 (O_17,N_2984,N_2965);
xor UO_18 (O_18,N_2958,N_2947);
nand UO_19 (O_19,N_2971,N_2928);
nand UO_20 (O_20,N_2994,N_2970);
nor UO_21 (O_21,N_2931,N_2967);
nor UO_22 (O_22,N_2949,N_2979);
or UO_23 (O_23,N_2930,N_2966);
xnor UO_24 (O_24,N_2991,N_2977);
xnor UO_25 (O_25,N_2986,N_2980);
xnor UO_26 (O_26,N_2960,N_2937);
xor UO_27 (O_27,N_2997,N_2954);
nor UO_28 (O_28,N_2944,N_2932);
and UO_29 (O_29,N_2950,N_2995);
nor UO_30 (O_30,N_2952,N_2996);
nand UO_31 (O_31,N_2953,N_2998);
nand UO_32 (O_32,N_2925,N_2933);
nor UO_33 (O_33,N_2985,N_2927);
or UO_34 (O_34,N_2993,N_2983);
nand UO_35 (O_35,N_2981,N_2948);
nor UO_36 (O_36,N_2963,N_2936);
or UO_37 (O_37,N_2982,N_2998);
or UO_38 (O_38,N_2928,N_2935);
nand UO_39 (O_39,N_2981,N_2991);
and UO_40 (O_40,N_2939,N_2973);
and UO_41 (O_41,N_2989,N_2931);
xor UO_42 (O_42,N_2981,N_2990);
or UO_43 (O_43,N_2940,N_2936);
xor UO_44 (O_44,N_2956,N_2987);
and UO_45 (O_45,N_2937,N_2949);
or UO_46 (O_46,N_2956,N_2928);
and UO_47 (O_47,N_2929,N_2957);
nand UO_48 (O_48,N_2963,N_2937);
and UO_49 (O_49,N_2971,N_2934);
and UO_50 (O_50,N_2992,N_2940);
and UO_51 (O_51,N_2926,N_2960);
and UO_52 (O_52,N_2950,N_2985);
and UO_53 (O_53,N_2973,N_2931);
nor UO_54 (O_54,N_2950,N_2963);
or UO_55 (O_55,N_2949,N_2984);
or UO_56 (O_56,N_2998,N_2958);
and UO_57 (O_57,N_2954,N_2976);
nor UO_58 (O_58,N_2999,N_2953);
nor UO_59 (O_59,N_2929,N_2954);
nor UO_60 (O_60,N_2956,N_2939);
nor UO_61 (O_61,N_2968,N_2981);
or UO_62 (O_62,N_2983,N_2986);
xor UO_63 (O_63,N_2956,N_2947);
nor UO_64 (O_64,N_2979,N_2984);
nand UO_65 (O_65,N_2944,N_2950);
xnor UO_66 (O_66,N_2950,N_2958);
nor UO_67 (O_67,N_2940,N_2943);
or UO_68 (O_68,N_2978,N_2992);
nor UO_69 (O_69,N_2949,N_2941);
nand UO_70 (O_70,N_2961,N_2950);
and UO_71 (O_71,N_2927,N_2932);
and UO_72 (O_72,N_2974,N_2961);
or UO_73 (O_73,N_2994,N_2992);
nor UO_74 (O_74,N_2963,N_2971);
nand UO_75 (O_75,N_2940,N_2968);
nor UO_76 (O_76,N_2985,N_2977);
nand UO_77 (O_77,N_2965,N_2938);
nand UO_78 (O_78,N_2971,N_2981);
nor UO_79 (O_79,N_2985,N_2928);
xnor UO_80 (O_80,N_2990,N_2949);
or UO_81 (O_81,N_2978,N_2951);
xor UO_82 (O_82,N_2993,N_2936);
or UO_83 (O_83,N_2980,N_2988);
xnor UO_84 (O_84,N_2944,N_2937);
nand UO_85 (O_85,N_2965,N_2964);
and UO_86 (O_86,N_2976,N_2969);
nand UO_87 (O_87,N_2925,N_2953);
nand UO_88 (O_88,N_2941,N_2925);
nor UO_89 (O_89,N_2929,N_2941);
nand UO_90 (O_90,N_2930,N_2985);
xor UO_91 (O_91,N_2968,N_2962);
nor UO_92 (O_92,N_2994,N_2971);
nor UO_93 (O_93,N_2975,N_2944);
nand UO_94 (O_94,N_2974,N_2978);
xnor UO_95 (O_95,N_2990,N_2986);
nor UO_96 (O_96,N_2925,N_2955);
nand UO_97 (O_97,N_2939,N_2980);
xor UO_98 (O_98,N_2968,N_2995);
and UO_99 (O_99,N_2942,N_2969);
nand UO_100 (O_100,N_2962,N_2963);
nand UO_101 (O_101,N_2973,N_2932);
nor UO_102 (O_102,N_2942,N_2931);
nand UO_103 (O_103,N_2948,N_2958);
nor UO_104 (O_104,N_2936,N_2943);
and UO_105 (O_105,N_2997,N_2960);
and UO_106 (O_106,N_2963,N_2927);
xnor UO_107 (O_107,N_2937,N_2927);
xor UO_108 (O_108,N_2945,N_2950);
xnor UO_109 (O_109,N_2946,N_2930);
and UO_110 (O_110,N_2950,N_2939);
or UO_111 (O_111,N_2964,N_2949);
or UO_112 (O_112,N_2997,N_2948);
nor UO_113 (O_113,N_2999,N_2984);
or UO_114 (O_114,N_2942,N_2959);
nor UO_115 (O_115,N_2974,N_2953);
nor UO_116 (O_116,N_2970,N_2946);
nand UO_117 (O_117,N_2986,N_2997);
nor UO_118 (O_118,N_2932,N_2962);
and UO_119 (O_119,N_2939,N_2991);
nor UO_120 (O_120,N_2929,N_2950);
and UO_121 (O_121,N_2932,N_2940);
xnor UO_122 (O_122,N_2949,N_2931);
xnor UO_123 (O_123,N_2955,N_2933);
or UO_124 (O_124,N_2968,N_2991);
nor UO_125 (O_125,N_2960,N_2963);
or UO_126 (O_126,N_2925,N_2993);
nand UO_127 (O_127,N_2977,N_2976);
and UO_128 (O_128,N_2980,N_2977);
and UO_129 (O_129,N_2949,N_2987);
nand UO_130 (O_130,N_2932,N_2929);
nand UO_131 (O_131,N_2977,N_2967);
or UO_132 (O_132,N_2964,N_2954);
nand UO_133 (O_133,N_2966,N_2981);
nand UO_134 (O_134,N_2964,N_2933);
or UO_135 (O_135,N_2995,N_2943);
xnor UO_136 (O_136,N_2965,N_2935);
xor UO_137 (O_137,N_2935,N_2926);
xor UO_138 (O_138,N_2963,N_2979);
and UO_139 (O_139,N_2930,N_2975);
and UO_140 (O_140,N_2936,N_2985);
and UO_141 (O_141,N_2964,N_2987);
and UO_142 (O_142,N_2999,N_2996);
and UO_143 (O_143,N_2937,N_2987);
and UO_144 (O_144,N_2986,N_2973);
nand UO_145 (O_145,N_2993,N_2966);
nor UO_146 (O_146,N_2936,N_2989);
nor UO_147 (O_147,N_2987,N_2946);
or UO_148 (O_148,N_2978,N_2928);
xnor UO_149 (O_149,N_2992,N_2939);
nor UO_150 (O_150,N_2946,N_2964);
nand UO_151 (O_151,N_2984,N_2967);
and UO_152 (O_152,N_2961,N_2981);
xor UO_153 (O_153,N_2927,N_2935);
or UO_154 (O_154,N_2958,N_2937);
or UO_155 (O_155,N_2960,N_2989);
nor UO_156 (O_156,N_2946,N_2984);
nand UO_157 (O_157,N_2952,N_2944);
xnor UO_158 (O_158,N_2972,N_2967);
nand UO_159 (O_159,N_2997,N_2977);
or UO_160 (O_160,N_2959,N_2979);
xnor UO_161 (O_161,N_2925,N_2961);
nor UO_162 (O_162,N_2950,N_2993);
nand UO_163 (O_163,N_2987,N_2971);
nor UO_164 (O_164,N_2944,N_2979);
nor UO_165 (O_165,N_2985,N_2988);
or UO_166 (O_166,N_2961,N_2964);
nand UO_167 (O_167,N_2952,N_2933);
xnor UO_168 (O_168,N_2987,N_2982);
nor UO_169 (O_169,N_2947,N_2965);
and UO_170 (O_170,N_2972,N_2931);
nor UO_171 (O_171,N_2992,N_2968);
and UO_172 (O_172,N_2988,N_2976);
xor UO_173 (O_173,N_2928,N_2927);
or UO_174 (O_174,N_2925,N_2982);
xor UO_175 (O_175,N_2982,N_2991);
nand UO_176 (O_176,N_2957,N_2941);
and UO_177 (O_177,N_2982,N_2972);
nor UO_178 (O_178,N_2940,N_2948);
xor UO_179 (O_179,N_2991,N_2945);
and UO_180 (O_180,N_2953,N_2985);
and UO_181 (O_181,N_2977,N_2960);
and UO_182 (O_182,N_2939,N_2977);
nand UO_183 (O_183,N_2987,N_2928);
and UO_184 (O_184,N_2943,N_2999);
or UO_185 (O_185,N_2994,N_2998);
nand UO_186 (O_186,N_2934,N_2994);
nor UO_187 (O_187,N_2965,N_2983);
and UO_188 (O_188,N_2947,N_2960);
nor UO_189 (O_189,N_2971,N_2943);
nor UO_190 (O_190,N_2951,N_2963);
nor UO_191 (O_191,N_2959,N_2963);
and UO_192 (O_192,N_2990,N_2979);
nand UO_193 (O_193,N_2982,N_2941);
nor UO_194 (O_194,N_2975,N_2996);
nand UO_195 (O_195,N_2953,N_2964);
and UO_196 (O_196,N_2946,N_2949);
or UO_197 (O_197,N_2938,N_2971);
nor UO_198 (O_198,N_2930,N_2947);
nor UO_199 (O_199,N_2994,N_2982);
or UO_200 (O_200,N_2997,N_2941);
xnor UO_201 (O_201,N_2935,N_2954);
or UO_202 (O_202,N_2931,N_2994);
xor UO_203 (O_203,N_2985,N_2938);
and UO_204 (O_204,N_2928,N_2973);
and UO_205 (O_205,N_2953,N_2933);
nor UO_206 (O_206,N_2925,N_2945);
and UO_207 (O_207,N_2984,N_2959);
and UO_208 (O_208,N_2958,N_2951);
nand UO_209 (O_209,N_2964,N_2960);
nor UO_210 (O_210,N_2934,N_2950);
or UO_211 (O_211,N_2997,N_2926);
and UO_212 (O_212,N_2967,N_2926);
and UO_213 (O_213,N_2926,N_2982);
nor UO_214 (O_214,N_2963,N_2945);
or UO_215 (O_215,N_2951,N_2974);
or UO_216 (O_216,N_2989,N_2994);
and UO_217 (O_217,N_2982,N_2997);
and UO_218 (O_218,N_2944,N_2955);
and UO_219 (O_219,N_2983,N_2947);
nor UO_220 (O_220,N_2985,N_2980);
xor UO_221 (O_221,N_2974,N_2930);
nand UO_222 (O_222,N_2983,N_2926);
nor UO_223 (O_223,N_2991,N_2930);
nor UO_224 (O_224,N_2927,N_2973);
nor UO_225 (O_225,N_2946,N_2982);
nand UO_226 (O_226,N_2981,N_2955);
xor UO_227 (O_227,N_2936,N_2976);
or UO_228 (O_228,N_2979,N_2975);
nand UO_229 (O_229,N_2940,N_2977);
or UO_230 (O_230,N_2934,N_2933);
nor UO_231 (O_231,N_2947,N_2942);
nor UO_232 (O_232,N_2933,N_2979);
or UO_233 (O_233,N_2937,N_2999);
xnor UO_234 (O_234,N_2954,N_2949);
and UO_235 (O_235,N_2955,N_2985);
xor UO_236 (O_236,N_2964,N_2984);
nand UO_237 (O_237,N_2952,N_2960);
nor UO_238 (O_238,N_2953,N_2967);
and UO_239 (O_239,N_2926,N_2995);
or UO_240 (O_240,N_2936,N_2980);
or UO_241 (O_241,N_2998,N_2967);
or UO_242 (O_242,N_2947,N_2999);
xnor UO_243 (O_243,N_2940,N_2980);
and UO_244 (O_244,N_2932,N_2992);
xor UO_245 (O_245,N_2937,N_2946);
nand UO_246 (O_246,N_2957,N_2950);
or UO_247 (O_247,N_2979,N_2928);
nand UO_248 (O_248,N_2944,N_2987);
nor UO_249 (O_249,N_2956,N_2986);
or UO_250 (O_250,N_2929,N_2964);
nand UO_251 (O_251,N_2978,N_2963);
and UO_252 (O_252,N_2955,N_2969);
and UO_253 (O_253,N_2945,N_2992);
nand UO_254 (O_254,N_2998,N_2986);
nor UO_255 (O_255,N_2979,N_2942);
or UO_256 (O_256,N_2976,N_2956);
nand UO_257 (O_257,N_2965,N_2957);
nand UO_258 (O_258,N_2996,N_2963);
or UO_259 (O_259,N_2977,N_2995);
nand UO_260 (O_260,N_2960,N_2984);
nand UO_261 (O_261,N_2976,N_2992);
and UO_262 (O_262,N_2927,N_2942);
or UO_263 (O_263,N_2958,N_2968);
nor UO_264 (O_264,N_2928,N_2977);
and UO_265 (O_265,N_2989,N_2944);
or UO_266 (O_266,N_2976,N_2984);
and UO_267 (O_267,N_2998,N_2974);
nand UO_268 (O_268,N_2952,N_2972);
and UO_269 (O_269,N_2944,N_2956);
nor UO_270 (O_270,N_2954,N_2944);
nand UO_271 (O_271,N_2987,N_2993);
nor UO_272 (O_272,N_2995,N_2949);
and UO_273 (O_273,N_2973,N_2996);
xor UO_274 (O_274,N_2955,N_2984);
nand UO_275 (O_275,N_2977,N_2932);
xor UO_276 (O_276,N_2934,N_2942);
xnor UO_277 (O_277,N_2929,N_2928);
and UO_278 (O_278,N_2967,N_2973);
nand UO_279 (O_279,N_2955,N_2931);
nor UO_280 (O_280,N_2946,N_2972);
or UO_281 (O_281,N_2950,N_2974);
nand UO_282 (O_282,N_2930,N_2952);
or UO_283 (O_283,N_2939,N_2969);
nor UO_284 (O_284,N_2925,N_2969);
nor UO_285 (O_285,N_2951,N_2992);
nor UO_286 (O_286,N_2943,N_2953);
nand UO_287 (O_287,N_2981,N_2999);
nor UO_288 (O_288,N_2931,N_2927);
and UO_289 (O_289,N_2992,N_2972);
nand UO_290 (O_290,N_2989,N_2949);
xor UO_291 (O_291,N_2978,N_2958);
nand UO_292 (O_292,N_2942,N_2996);
nor UO_293 (O_293,N_2983,N_2956);
and UO_294 (O_294,N_2956,N_2950);
or UO_295 (O_295,N_2936,N_2992);
xor UO_296 (O_296,N_2968,N_2949);
xor UO_297 (O_297,N_2977,N_2966);
and UO_298 (O_298,N_2961,N_2976);
or UO_299 (O_299,N_2929,N_2955);
nor UO_300 (O_300,N_2932,N_2976);
xnor UO_301 (O_301,N_2935,N_2973);
nand UO_302 (O_302,N_2979,N_2962);
nand UO_303 (O_303,N_2995,N_2930);
xnor UO_304 (O_304,N_2985,N_2982);
nand UO_305 (O_305,N_2977,N_2951);
or UO_306 (O_306,N_2964,N_2995);
and UO_307 (O_307,N_2992,N_2950);
xnor UO_308 (O_308,N_2942,N_2946);
nand UO_309 (O_309,N_2935,N_2967);
xor UO_310 (O_310,N_2944,N_2960);
nor UO_311 (O_311,N_2983,N_2996);
nor UO_312 (O_312,N_2946,N_2935);
xnor UO_313 (O_313,N_2978,N_2930);
nor UO_314 (O_314,N_2973,N_2974);
or UO_315 (O_315,N_2931,N_2957);
nor UO_316 (O_316,N_2966,N_2948);
nor UO_317 (O_317,N_2991,N_2975);
and UO_318 (O_318,N_2997,N_2971);
and UO_319 (O_319,N_2955,N_2928);
nor UO_320 (O_320,N_2990,N_2944);
or UO_321 (O_321,N_2973,N_2951);
nor UO_322 (O_322,N_2938,N_2997);
xor UO_323 (O_323,N_2957,N_2937);
nand UO_324 (O_324,N_2987,N_2959);
or UO_325 (O_325,N_2997,N_2946);
and UO_326 (O_326,N_2994,N_2933);
nor UO_327 (O_327,N_2959,N_2928);
nor UO_328 (O_328,N_2957,N_2995);
nor UO_329 (O_329,N_2978,N_2969);
and UO_330 (O_330,N_2977,N_2988);
and UO_331 (O_331,N_2976,N_2986);
or UO_332 (O_332,N_2960,N_2957);
nor UO_333 (O_333,N_2968,N_2978);
nor UO_334 (O_334,N_2944,N_2978);
nor UO_335 (O_335,N_2977,N_2999);
xnor UO_336 (O_336,N_2999,N_2992);
and UO_337 (O_337,N_2948,N_2935);
nand UO_338 (O_338,N_2933,N_2937);
and UO_339 (O_339,N_2955,N_2980);
nand UO_340 (O_340,N_2938,N_2934);
or UO_341 (O_341,N_2936,N_2949);
and UO_342 (O_342,N_2972,N_2976);
and UO_343 (O_343,N_2986,N_2930);
xor UO_344 (O_344,N_2980,N_2992);
nand UO_345 (O_345,N_2947,N_2987);
nand UO_346 (O_346,N_2935,N_2959);
or UO_347 (O_347,N_2993,N_2938);
or UO_348 (O_348,N_2960,N_2950);
xor UO_349 (O_349,N_2928,N_2947);
nand UO_350 (O_350,N_2979,N_2983);
or UO_351 (O_351,N_2939,N_2990);
or UO_352 (O_352,N_2959,N_2943);
nand UO_353 (O_353,N_2959,N_2951);
xor UO_354 (O_354,N_2994,N_2987);
nor UO_355 (O_355,N_2978,N_2939);
nand UO_356 (O_356,N_2958,N_2940);
and UO_357 (O_357,N_2953,N_2962);
nand UO_358 (O_358,N_2984,N_2936);
or UO_359 (O_359,N_2972,N_2995);
and UO_360 (O_360,N_2972,N_2998);
nand UO_361 (O_361,N_2959,N_2955);
nand UO_362 (O_362,N_2984,N_2986);
nor UO_363 (O_363,N_2959,N_2939);
and UO_364 (O_364,N_2985,N_2942);
nand UO_365 (O_365,N_2930,N_2970);
nand UO_366 (O_366,N_2986,N_2996);
or UO_367 (O_367,N_2978,N_2950);
and UO_368 (O_368,N_2986,N_2972);
nor UO_369 (O_369,N_2964,N_2975);
or UO_370 (O_370,N_2985,N_2981);
or UO_371 (O_371,N_2985,N_2956);
and UO_372 (O_372,N_2986,N_2948);
nor UO_373 (O_373,N_2989,N_2942);
and UO_374 (O_374,N_2941,N_2989);
nor UO_375 (O_375,N_2931,N_2954);
nand UO_376 (O_376,N_2998,N_2995);
or UO_377 (O_377,N_2973,N_2938);
nand UO_378 (O_378,N_2939,N_2942);
nor UO_379 (O_379,N_2943,N_2950);
or UO_380 (O_380,N_2980,N_2996);
and UO_381 (O_381,N_2997,N_2966);
or UO_382 (O_382,N_2985,N_2944);
and UO_383 (O_383,N_2938,N_2989);
or UO_384 (O_384,N_2965,N_2946);
nor UO_385 (O_385,N_2972,N_2938);
xor UO_386 (O_386,N_2958,N_2938);
and UO_387 (O_387,N_2963,N_2939);
or UO_388 (O_388,N_2975,N_2963);
nor UO_389 (O_389,N_2990,N_2951);
nor UO_390 (O_390,N_2931,N_2950);
nor UO_391 (O_391,N_2965,N_2961);
xnor UO_392 (O_392,N_2960,N_2955);
nand UO_393 (O_393,N_2941,N_2947);
nand UO_394 (O_394,N_2973,N_2956);
nand UO_395 (O_395,N_2968,N_2935);
and UO_396 (O_396,N_2954,N_2946);
xor UO_397 (O_397,N_2955,N_2936);
and UO_398 (O_398,N_2981,N_2946);
nand UO_399 (O_399,N_2951,N_2926);
nor UO_400 (O_400,N_2982,N_2954);
or UO_401 (O_401,N_2936,N_2932);
nand UO_402 (O_402,N_2977,N_2947);
xor UO_403 (O_403,N_2936,N_2958);
nand UO_404 (O_404,N_2950,N_2936);
and UO_405 (O_405,N_2968,N_2985);
nor UO_406 (O_406,N_2970,N_2972);
nand UO_407 (O_407,N_2971,N_2925);
xor UO_408 (O_408,N_2942,N_2956);
or UO_409 (O_409,N_2951,N_2979);
nor UO_410 (O_410,N_2945,N_2989);
nor UO_411 (O_411,N_2974,N_2965);
xnor UO_412 (O_412,N_2928,N_2953);
nor UO_413 (O_413,N_2933,N_2970);
xor UO_414 (O_414,N_2963,N_2955);
and UO_415 (O_415,N_2944,N_2936);
nor UO_416 (O_416,N_2929,N_2986);
xnor UO_417 (O_417,N_2982,N_2989);
nor UO_418 (O_418,N_2957,N_2982);
and UO_419 (O_419,N_2969,N_2968);
and UO_420 (O_420,N_2999,N_2979);
xor UO_421 (O_421,N_2950,N_2940);
nor UO_422 (O_422,N_2952,N_2997);
or UO_423 (O_423,N_2974,N_2983);
and UO_424 (O_424,N_2979,N_2961);
nand UO_425 (O_425,N_2984,N_2966);
nor UO_426 (O_426,N_2995,N_2947);
xnor UO_427 (O_427,N_2943,N_2927);
nand UO_428 (O_428,N_2976,N_2951);
nand UO_429 (O_429,N_2964,N_2948);
and UO_430 (O_430,N_2954,N_2938);
or UO_431 (O_431,N_2979,N_2925);
nor UO_432 (O_432,N_2928,N_2991);
or UO_433 (O_433,N_2992,N_2946);
xor UO_434 (O_434,N_2986,N_2966);
xnor UO_435 (O_435,N_2957,N_2940);
xnor UO_436 (O_436,N_2972,N_2954);
and UO_437 (O_437,N_2997,N_2939);
nor UO_438 (O_438,N_2988,N_2996);
and UO_439 (O_439,N_2953,N_2945);
or UO_440 (O_440,N_2935,N_2951);
or UO_441 (O_441,N_2993,N_2972);
and UO_442 (O_442,N_2989,N_2990);
nor UO_443 (O_443,N_2946,N_2963);
xnor UO_444 (O_444,N_2969,N_2965);
or UO_445 (O_445,N_2941,N_2963);
nor UO_446 (O_446,N_2996,N_2965);
or UO_447 (O_447,N_2976,N_2940);
xor UO_448 (O_448,N_2942,N_2940);
nand UO_449 (O_449,N_2990,N_2995);
xnor UO_450 (O_450,N_2933,N_2983);
nand UO_451 (O_451,N_2971,N_2984);
nand UO_452 (O_452,N_2953,N_2996);
nor UO_453 (O_453,N_2973,N_2949);
or UO_454 (O_454,N_2993,N_2995);
and UO_455 (O_455,N_2973,N_2972);
or UO_456 (O_456,N_2935,N_2976);
and UO_457 (O_457,N_2996,N_2970);
nand UO_458 (O_458,N_2961,N_2987);
nor UO_459 (O_459,N_2978,N_2995);
nor UO_460 (O_460,N_2974,N_2934);
xor UO_461 (O_461,N_2945,N_2986);
or UO_462 (O_462,N_2979,N_2966);
or UO_463 (O_463,N_2977,N_2931);
or UO_464 (O_464,N_2986,N_2934);
xor UO_465 (O_465,N_2989,N_2961);
nand UO_466 (O_466,N_2955,N_2937);
or UO_467 (O_467,N_2997,N_2950);
xor UO_468 (O_468,N_2979,N_2994);
xor UO_469 (O_469,N_2977,N_2930);
or UO_470 (O_470,N_2996,N_2984);
xor UO_471 (O_471,N_2975,N_2926);
xnor UO_472 (O_472,N_2989,N_2986);
and UO_473 (O_473,N_2981,N_2953);
nand UO_474 (O_474,N_2999,N_2929);
or UO_475 (O_475,N_2963,N_2933);
nand UO_476 (O_476,N_2969,N_2980);
nand UO_477 (O_477,N_2995,N_2937);
nand UO_478 (O_478,N_2952,N_2954);
nor UO_479 (O_479,N_2928,N_2995);
xnor UO_480 (O_480,N_2976,N_2996);
nor UO_481 (O_481,N_2926,N_2934);
or UO_482 (O_482,N_2990,N_2938);
nor UO_483 (O_483,N_2971,N_2982);
and UO_484 (O_484,N_2963,N_2982);
nand UO_485 (O_485,N_2978,N_2925);
nor UO_486 (O_486,N_2962,N_2985);
nand UO_487 (O_487,N_2985,N_2947);
nand UO_488 (O_488,N_2942,N_2975);
nand UO_489 (O_489,N_2957,N_2971);
nor UO_490 (O_490,N_2965,N_2967);
nand UO_491 (O_491,N_2965,N_2966);
nand UO_492 (O_492,N_2943,N_2987);
or UO_493 (O_493,N_2999,N_2942);
or UO_494 (O_494,N_2964,N_2968);
or UO_495 (O_495,N_2953,N_2978);
or UO_496 (O_496,N_2987,N_2992);
xnor UO_497 (O_497,N_2956,N_2996);
nor UO_498 (O_498,N_2932,N_2934);
nand UO_499 (O_499,N_2939,N_2951);
endmodule