module basic_1000_10000_1500_10_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_38,In_879);
or U1 (N_1,In_399,In_331);
nand U2 (N_2,In_592,In_178);
nand U3 (N_3,In_71,In_885);
and U4 (N_4,In_395,In_924);
nand U5 (N_5,In_710,In_638);
or U6 (N_6,In_257,In_859);
nand U7 (N_7,In_367,In_597);
nor U8 (N_8,In_905,In_610);
or U9 (N_9,In_670,In_931);
and U10 (N_10,In_543,In_474);
xnor U11 (N_11,In_700,In_66);
nor U12 (N_12,In_968,In_351);
or U13 (N_13,In_504,In_138);
and U14 (N_14,In_45,In_645);
nand U15 (N_15,In_761,In_42);
nor U16 (N_16,In_908,In_196);
or U17 (N_17,In_759,In_280);
and U18 (N_18,In_371,In_807);
nand U19 (N_19,In_104,In_920);
nor U20 (N_20,In_277,In_758);
nor U21 (N_21,In_602,In_70);
nand U22 (N_22,In_169,In_40);
xor U23 (N_23,In_37,In_381);
xor U24 (N_24,In_890,In_157);
or U25 (N_25,In_883,In_869);
nand U26 (N_26,In_339,In_994);
and U27 (N_27,In_526,In_158);
or U28 (N_28,In_407,In_631);
nor U29 (N_29,In_240,In_820);
xor U30 (N_30,In_334,In_507);
and U31 (N_31,In_545,In_460);
nand U32 (N_32,In_141,In_11);
nor U33 (N_33,In_753,In_176);
nand U34 (N_34,In_58,In_706);
and U35 (N_35,In_798,In_957);
nor U36 (N_36,In_802,In_296);
or U37 (N_37,In_168,In_637);
xor U38 (N_38,In_396,In_958);
or U39 (N_39,In_223,In_677);
xnor U40 (N_40,In_711,In_363);
or U41 (N_41,In_875,In_906);
xor U42 (N_42,In_995,In_94);
or U43 (N_43,In_854,In_934);
and U44 (N_44,In_531,In_208);
nor U45 (N_45,In_326,In_946);
nand U46 (N_46,In_659,In_85);
and U47 (N_47,In_726,In_27);
xor U48 (N_48,In_292,In_671);
and U49 (N_49,In_375,In_118);
nor U50 (N_50,In_213,In_693);
nand U51 (N_51,In_812,In_254);
nor U52 (N_52,In_311,In_727);
nand U53 (N_53,In_201,In_180);
or U54 (N_54,In_166,In_751);
or U55 (N_55,In_252,In_356);
nand U56 (N_56,In_835,In_943);
and U57 (N_57,In_225,In_792);
or U58 (N_58,In_830,In_956);
and U59 (N_59,In_839,In_676);
or U60 (N_60,In_762,In_817);
nand U61 (N_61,In_337,In_805);
or U62 (N_62,In_725,In_86);
and U63 (N_63,In_886,In_480);
nor U64 (N_64,In_465,In_33);
or U65 (N_65,In_198,In_188);
nor U66 (N_66,In_861,In_980);
nand U67 (N_67,In_224,In_183);
xnor U68 (N_68,In_205,In_982);
or U69 (N_69,In_662,In_343);
and U70 (N_70,In_773,In_728);
and U71 (N_71,In_453,In_193);
nor U72 (N_72,In_954,In_495);
xnor U73 (N_73,In_437,In_10);
or U74 (N_74,In_642,In_698);
xor U75 (N_75,In_16,In_630);
nor U76 (N_76,In_272,In_22);
or U77 (N_77,In_528,In_264);
nor U78 (N_78,In_215,In_1);
nor U79 (N_79,In_632,In_900);
nand U80 (N_80,In_942,In_179);
nor U81 (N_81,In_44,In_595);
or U82 (N_82,In_527,In_394);
or U83 (N_83,In_837,In_133);
and U84 (N_84,In_865,In_56);
or U85 (N_85,In_189,In_987);
or U86 (N_86,In_406,In_628);
and U87 (N_87,In_578,In_534);
and U88 (N_88,In_82,In_867);
nand U89 (N_89,In_226,In_944);
nand U90 (N_90,In_986,In_23);
xor U91 (N_91,In_540,In_397);
nand U92 (N_92,In_61,In_350);
nor U93 (N_93,In_888,In_919);
nand U94 (N_94,In_7,In_409);
nor U95 (N_95,In_818,In_473);
and U96 (N_96,In_788,In_64);
nor U97 (N_97,In_449,In_521);
and U98 (N_98,In_243,In_652);
or U99 (N_99,In_90,In_742);
or U100 (N_100,In_911,In_53);
or U101 (N_101,In_787,In_947);
nand U102 (N_102,In_562,In_868);
xor U103 (N_103,In_232,In_748);
and U104 (N_104,In_194,In_450);
and U105 (N_105,In_953,In_997);
nand U106 (N_106,In_466,In_236);
and U107 (N_107,In_616,In_784);
and U108 (N_108,In_413,In_569);
nor U109 (N_109,In_889,In_320);
or U110 (N_110,In_800,In_490);
and U111 (N_111,In_846,In_596);
nor U112 (N_112,In_649,In_845);
nor U113 (N_113,In_467,In_96);
nor U114 (N_114,In_503,In_945);
or U115 (N_115,In_195,In_657);
xnor U116 (N_116,In_511,In_689);
or U117 (N_117,In_357,In_36);
nor U118 (N_118,In_952,In_472);
nor U119 (N_119,In_881,In_667);
xor U120 (N_120,In_855,In_216);
nand U121 (N_121,In_77,In_147);
and U122 (N_122,In_778,In_414);
xnor U123 (N_123,In_156,In_585);
nor U124 (N_124,In_59,In_162);
nand U125 (N_125,In_563,In_163);
nor U126 (N_126,In_813,In_523);
nand U127 (N_127,In_288,In_591);
nor U128 (N_128,In_419,In_28);
nor U129 (N_129,In_332,In_404);
nor U130 (N_130,In_456,In_873);
nand U131 (N_131,In_127,In_750);
nand U132 (N_132,In_43,In_432);
nor U133 (N_133,In_244,In_341);
and U134 (N_134,In_468,In_191);
nor U135 (N_135,In_546,In_768);
nor U136 (N_136,In_791,In_478);
or U137 (N_137,In_650,In_744);
xnor U138 (N_138,In_145,In_427);
and U139 (N_139,In_826,In_187);
and U140 (N_140,In_423,In_458);
or U141 (N_141,In_993,In_114);
and U142 (N_142,In_228,In_740);
nand U143 (N_143,In_72,In_69);
xnor U144 (N_144,In_418,In_832);
nand U145 (N_145,In_874,In_68);
nand U146 (N_146,In_603,In_15);
and U147 (N_147,In_655,In_428);
xnor U148 (N_148,In_779,In_471);
nor U149 (N_149,In_629,In_705);
nor U150 (N_150,In_2,In_197);
nor U151 (N_151,In_338,In_488);
or U152 (N_152,In_828,In_661);
nor U153 (N_153,In_360,In_261);
nand U154 (N_154,In_576,In_314);
or U155 (N_155,In_653,In_789);
or U156 (N_156,In_310,In_312);
and U157 (N_157,In_513,In_416);
nor U158 (N_158,In_134,In_441);
nand U159 (N_159,In_482,In_305);
nor U160 (N_160,In_489,In_870);
or U161 (N_161,In_524,In_673);
and U162 (N_162,In_303,In_249);
or U163 (N_163,In_590,In_581);
nand U164 (N_164,In_206,In_119);
nor U165 (N_165,In_278,In_716);
xor U166 (N_166,In_799,In_864);
and U167 (N_167,In_283,In_568);
or U168 (N_168,In_965,In_763);
nand U169 (N_169,In_810,In_365);
and U170 (N_170,In_608,In_439);
or U171 (N_171,In_695,In_424);
nor U172 (N_172,In_109,In_959);
or U173 (N_173,In_8,In_697);
nor U174 (N_174,In_398,In_914);
and U175 (N_175,In_151,In_101);
or U176 (N_176,In_464,In_829);
nor U177 (N_177,In_937,In_186);
nand U178 (N_178,In_739,In_366);
nand U179 (N_179,In_455,In_79);
nor U180 (N_180,In_627,In_301);
and U181 (N_181,In_75,In_654);
nor U182 (N_182,In_690,In_493);
and U183 (N_183,In_843,In_315);
and U184 (N_184,In_410,In_512);
nor U185 (N_185,In_614,In_125);
nand U186 (N_186,In_160,In_408);
nand U187 (N_187,In_459,In_483);
nor U188 (N_188,In_260,In_626);
and U189 (N_189,In_594,In_856);
nor U190 (N_190,In_391,In_892);
and U191 (N_191,In_926,In_227);
and U192 (N_192,In_267,In_620);
nand U193 (N_193,In_538,In_373);
and U194 (N_194,In_378,In_979);
nor U195 (N_195,In_938,In_295);
nand U196 (N_196,In_918,In_76);
and U197 (N_197,In_734,In_34);
or U198 (N_198,In_775,In_374);
nand U199 (N_199,In_539,In_477);
or U200 (N_200,In_47,In_348);
nand U201 (N_201,In_731,In_701);
nand U202 (N_202,In_207,In_896);
nand U203 (N_203,In_411,In_962);
nor U204 (N_204,In_730,In_929);
or U205 (N_205,In_971,In_492);
and U206 (N_206,In_74,In_939);
and U207 (N_207,In_440,In_549);
and U208 (N_208,In_951,In_785);
and U209 (N_209,In_840,In_403);
or U210 (N_210,In_200,In_684);
and U211 (N_211,In_850,In_89);
and U212 (N_212,In_308,In_48);
and U213 (N_213,In_299,In_152);
and U214 (N_214,In_816,In_841);
xnor U215 (N_215,In_290,In_497);
or U216 (N_216,In_173,In_412);
nand U217 (N_217,In_170,In_532);
nor U218 (N_218,In_164,In_382);
or U219 (N_219,In_553,In_558);
or U220 (N_220,In_346,In_322);
or U221 (N_221,In_755,In_990);
and U222 (N_222,In_379,In_364);
or U223 (N_223,In_651,In_714);
or U224 (N_224,In_964,In_340);
nand U225 (N_225,In_81,In_948);
and U226 (N_226,In_849,In_910);
and U227 (N_227,In_229,In_936);
nor U228 (N_228,In_390,In_804);
nand U229 (N_229,In_421,In_289);
nor U230 (N_230,In_344,In_30);
and U231 (N_231,In_978,In_913);
xnor U232 (N_232,In_143,In_589);
nor U233 (N_233,In_606,In_611);
xor U234 (N_234,In_88,In_370);
nor U235 (N_235,In_192,In_362);
nand U236 (N_236,In_24,In_872);
nand U237 (N_237,In_447,In_239);
nor U238 (N_238,In_126,In_430);
or U239 (N_239,In_970,In_902);
or U240 (N_240,In_559,In_199);
nor U241 (N_241,In_479,In_781);
nor U242 (N_242,In_831,In_794);
nand U243 (N_243,In_185,In_230);
nand U244 (N_244,In_112,In_570);
nor U245 (N_245,In_517,In_612);
nor U246 (N_246,In_117,In_67);
or U247 (N_247,In_674,In_694);
nor U248 (N_248,In_102,In_454);
nand U249 (N_249,In_369,In_756);
or U250 (N_250,In_878,In_498);
nand U251 (N_251,In_722,In_83);
or U252 (N_252,In_636,In_641);
and U253 (N_253,In_501,In_715);
or U254 (N_254,In_552,In_52);
nor U255 (N_255,In_3,In_294);
xnor U256 (N_256,In_274,In_159);
or U257 (N_257,In_675,In_564);
xor U258 (N_258,In_644,In_177);
nor U259 (N_259,In_767,In_898);
nand U260 (N_260,In_721,In_827);
nor U261 (N_261,In_123,In_231);
nor U262 (N_262,In_385,In_702);
xor U263 (N_263,In_359,In_237);
nor U264 (N_264,In_848,In_933);
and U265 (N_265,In_941,In_907);
and U266 (N_266,In_729,In_451);
and U267 (N_267,In_98,In_745);
and U268 (N_268,In_733,In_664);
and U269 (N_269,In_882,In_271);
nand U270 (N_270,In_887,In_613);
nor U271 (N_271,In_108,In_577);
xor U272 (N_272,In_723,In_258);
nor U273 (N_273,In_685,In_646);
nor U274 (N_274,In_121,In_448);
xor U275 (N_275,In_130,In_536);
nand U276 (N_276,In_836,In_949);
nand U277 (N_277,In_361,In_372);
nand U278 (N_278,In_273,In_678);
nand U279 (N_279,In_304,In_647);
nand U280 (N_280,In_897,In_87);
and U281 (N_281,In_438,In_182);
or U282 (N_282,In_55,In_317);
nor U283 (N_283,In_318,In_420);
nor U284 (N_284,In_91,In_822);
nor U285 (N_285,In_253,In_853);
and U286 (N_286,In_509,In_604);
nor U287 (N_287,In_680,In_431);
nor U288 (N_288,In_144,In_737);
xnor U289 (N_289,In_648,In_99);
and U290 (N_290,In_62,In_541);
xnor U291 (N_291,In_858,In_245);
nor U292 (N_292,In_203,In_550);
or U293 (N_293,In_525,In_901);
nand U294 (N_294,In_5,In_452);
nand U295 (N_295,In_210,In_209);
nor U296 (N_296,In_247,In_150);
xnor U297 (N_297,In_422,In_508);
nand U298 (N_298,In_530,In_623);
nand U299 (N_299,In_19,In_884);
nor U300 (N_300,In_921,In_974);
and U301 (N_301,In_443,In_586);
and U302 (N_302,In_703,In_633);
nand U303 (N_303,In_686,In_746);
and U304 (N_304,In_4,In_214);
nand U305 (N_305,In_860,In_222);
or U306 (N_306,In_769,In_73);
nand U307 (N_307,In_640,In_969);
and U308 (N_308,In_960,In_707);
nor U309 (N_309,In_916,In_621);
nor U310 (N_310,In_146,In_302);
and U311 (N_311,In_579,In_485);
and U312 (N_312,In_772,In_107);
nor U313 (N_313,In_405,In_457);
nand U314 (N_314,In_863,In_128);
and U315 (N_315,In_866,In_354);
and U316 (N_316,In_29,In_12);
nand U317 (N_317,In_851,In_298);
and U318 (N_318,In_174,In_599);
nor U319 (N_319,In_246,In_821);
nand U320 (N_320,In_148,In_35);
or U321 (N_321,In_401,In_266);
nor U322 (N_322,In_708,In_461);
xnor U323 (N_323,In_129,In_393);
and U324 (N_324,In_270,In_241);
nor U325 (N_325,In_415,In_609);
nor U326 (N_326,In_462,In_446);
or U327 (N_327,In_801,In_732);
and U328 (N_328,In_32,In_560);
and U329 (N_329,In_475,In_780);
nor U330 (N_330,In_487,In_442);
nor U331 (N_331,In_388,In_622);
nand U332 (N_332,In_469,In_593);
nand U333 (N_333,In_814,In_218);
nand U334 (N_334,In_704,In_14);
and U335 (N_335,In_400,In_566);
nand U336 (N_336,In_793,In_97);
xor U337 (N_337,In_329,In_54);
nand U338 (N_338,In_65,In_238);
nor U339 (N_339,In_899,In_165);
or U340 (N_340,In_699,In_383);
nor U341 (N_341,In_154,In_551);
nor U342 (N_342,In_389,In_279);
and U343 (N_343,In_668,In_204);
and U344 (N_344,In_63,In_476);
xnor U345 (N_345,In_547,In_132);
and U346 (N_346,In_893,In_309);
or U347 (N_347,In_724,In_743);
nor U348 (N_348,In_41,In_998);
nand U349 (N_349,In_248,In_556);
nor U350 (N_350,In_571,In_605);
or U351 (N_351,In_757,In_752);
and U352 (N_352,In_561,In_0);
and U353 (N_353,In_542,In_306);
or U354 (N_354,In_287,In_696);
nand U355 (N_355,In_580,In_808);
nand U356 (N_356,In_93,In_712);
or U357 (N_357,In_766,In_21);
nand U358 (N_358,In_219,In_328);
xor U359 (N_359,In_983,In_297);
or U360 (N_360,In_774,In_516);
nand U361 (N_361,In_754,In_679);
nor U362 (N_362,In_358,In_131);
and U363 (N_363,In_481,In_909);
and U364 (N_364,In_17,In_928);
or U365 (N_365,In_352,In_984);
xnor U366 (N_366,In_484,In_996);
xnor U367 (N_367,In_323,In_796);
xnor U368 (N_368,In_220,In_790);
and U369 (N_369,In_417,In_286);
and U370 (N_370,In_377,In_262);
or U371 (N_371,In_683,In_293);
and U372 (N_372,In_307,In_575);
or U373 (N_373,In_51,In_124);
or U374 (N_374,In_717,In_316);
or U375 (N_375,In_242,In_565);
and U376 (N_376,In_925,In_520);
xnor U377 (N_377,In_738,In_190);
and U378 (N_378,In_434,In_6);
nor U379 (N_379,In_834,In_895);
and U380 (N_380,In_663,In_300);
nand U381 (N_381,In_506,In_284);
and U382 (N_382,In_991,In_115);
or U383 (N_383,In_588,In_172);
and U384 (N_384,In_666,In_347);
nand U385 (N_385,In_184,In_838);
and U386 (N_386,In_782,In_573);
nand U387 (N_387,In_555,In_135);
nor U388 (N_388,In_31,In_342);
nand U389 (N_389,In_665,In_202);
nand U390 (N_390,In_847,In_345);
nor U391 (N_391,In_463,In_321);
or U392 (N_392,In_276,In_607);
and U393 (N_393,In_291,In_966);
and U394 (N_394,In_786,In_880);
and U395 (N_395,In_435,In_100);
xor U396 (N_396,In_672,In_494);
and U397 (N_397,In_598,In_852);
xor U398 (N_398,In_999,In_537);
or U399 (N_399,In_429,In_353);
and U400 (N_400,In_9,In_903);
nand U401 (N_401,In_325,In_384);
nor U402 (N_402,In_368,In_735);
nand U403 (N_403,In_122,In_445);
or U404 (N_404,In_39,In_268);
and U405 (N_405,In_795,In_349);
or U406 (N_406,In_49,In_574);
or U407 (N_407,In_857,In_502);
nand U408 (N_408,In_444,In_103);
nand U409 (N_409,In_634,In_330);
or U410 (N_410,In_660,In_922);
and U411 (N_411,In_234,In_217);
and U412 (N_412,In_977,In_747);
and U413 (N_413,In_624,In_263);
nor U414 (N_414,In_819,In_572);
nor U415 (N_415,In_80,In_324);
nand U416 (N_416,In_967,In_486);
xnor U417 (N_417,In_60,In_691);
nor U418 (N_418,In_681,In_741);
and U419 (N_419,In_961,In_989);
and U420 (N_420,In_142,In_877);
and U421 (N_421,In_256,In_335);
nor U422 (N_422,In_842,In_776);
nor U423 (N_423,In_113,In_518);
and U424 (N_424,In_376,In_615);
nand U425 (N_425,In_402,In_777);
nand U426 (N_426,In_387,In_535);
nor U427 (N_427,In_930,In_149);
or U428 (N_428,In_171,In_643);
or U429 (N_429,In_491,In_770);
and U430 (N_430,In_932,In_600);
xor U431 (N_431,In_140,In_713);
and U432 (N_432,In_554,In_20);
xnor U433 (N_433,In_567,In_106);
nand U434 (N_434,In_582,In_815);
nand U435 (N_435,In_265,In_601);
or U436 (N_436,In_269,In_797);
and U437 (N_437,In_18,In_282);
and U438 (N_438,In_25,In_904);
xnor U439 (N_439,In_136,In_927);
xor U440 (N_440,In_514,In_78);
nor U441 (N_441,In_221,In_692);
and U442 (N_442,In_250,In_894);
or U443 (N_443,In_57,In_718);
or U444 (N_444,In_105,In_26);
or U445 (N_445,In_765,In_235);
nor U446 (N_446,In_688,In_811);
nor U447 (N_447,In_935,In_529);
nand U448 (N_448,In_720,In_809);
nand U449 (N_449,In_940,In_386);
nand U450 (N_450,In_824,In_496);
xor U451 (N_451,In_285,In_656);
nor U452 (N_452,In_233,In_46);
xnor U453 (N_453,In_181,In_275);
nor U454 (N_454,In_625,In_871);
or U455 (N_455,In_619,In_505);
nor U456 (N_456,In_584,In_380);
or U457 (N_457,In_319,In_963);
nor U458 (N_458,In_139,In_587);
nor U459 (N_459,In_736,In_862);
or U460 (N_460,In_955,In_500);
nand U461 (N_461,In_771,In_392);
nand U462 (N_462,In_618,In_973);
or U463 (N_463,In_803,In_825);
nand U464 (N_464,In_433,In_917);
nand U465 (N_465,In_639,In_992);
and U466 (N_466,In_544,In_912);
nand U467 (N_467,In_635,In_583);
nor U468 (N_468,In_120,In_155);
nor U469 (N_469,In_425,In_617);
xnor U470 (N_470,In_50,In_972);
or U471 (N_471,In_709,In_211);
and U472 (N_472,In_658,In_985);
or U473 (N_473,In_84,In_167);
nand U474 (N_474,In_259,In_281);
and U475 (N_475,In_764,In_981);
and U476 (N_476,In_175,In_950);
and U477 (N_477,In_212,In_153);
and U478 (N_478,In_876,In_111);
or U479 (N_479,In_251,In_333);
nand U480 (N_480,In_533,In_687);
xnor U481 (N_481,In_510,In_975);
nand U482 (N_482,In_336,In_823);
nor U483 (N_483,In_749,In_499);
nand U484 (N_484,In_95,In_313);
nor U485 (N_485,In_844,In_783);
nor U486 (N_486,In_161,In_116);
or U487 (N_487,In_436,In_682);
and U488 (N_488,In_519,In_806);
and U489 (N_489,In_669,In_355);
nor U490 (N_490,In_137,In_515);
nor U491 (N_491,In_833,In_426);
nand U492 (N_492,In_988,In_470);
xor U493 (N_493,In_760,In_891);
nor U494 (N_494,In_522,In_719);
or U495 (N_495,In_923,In_557);
and U496 (N_496,In_110,In_327);
and U497 (N_497,In_976,In_255);
nor U498 (N_498,In_13,In_92);
nand U499 (N_499,In_548,In_915);
nor U500 (N_500,In_598,In_579);
or U501 (N_501,In_627,In_824);
or U502 (N_502,In_837,In_581);
nor U503 (N_503,In_278,In_230);
nor U504 (N_504,In_681,In_587);
nor U505 (N_505,In_436,In_689);
xor U506 (N_506,In_942,In_645);
nand U507 (N_507,In_571,In_980);
nand U508 (N_508,In_127,In_170);
nor U509 (N_509,In_289,In_324);
and U510 (N_510,In_543,In_414);
and U511 (N_511,In_714,In_316);
or U512 (N_512,In_398,In_35);
xor U513 (N_513,In_24,In_388);
or U514 (N_514,In_666,In_572);
nor U515 (N_515,In_723,In_710);
nand U516 (N_516,In_113,In_240);
xnor U517 (N_517,In_624,In_750);
or U518 (N_518,In_6,In_47);
nor U519 (N_519,In_321,In_772);
or U520 (N_520,In_891,In_925);
or U521 (N_521,In_851,In_227);
and U522 (N_522,In_299,In_955);
or U523 (N_523,In_945,In_344);
and U524 (N_524,In_145,In_957);
and U525 (N_525,In_100,In_770);
nand U526 (N_526,In_867,In_612);
and U527 (N_527,In_347,In_844);
nor U528 (N_528,In_326,In_985);
nand U529 (N_529,In_216,In_903);
or U530 (N_530,In_643,In_554);
nor U531 (N_531,In_169,In_846);
or U532 (N_532,In_349,In_144);
or U533 (N_533,In_933,In_294);
nand U534 (N_534,In_567,In_976);
nor U535 (N_535,In_80,In_110);
and U536 (N_536,In_749,In_695);
or U537 (N_537,In_127,In_955);
nand U538 (N_538,In_387,In_658);
or U539 (N_539,In_487,In_962);
nor U540 (N_540,In_411,In_324);
and U541 (N_541,In_108,In_344);
or U542 (N_542,In_137,In_961);
nand U543 (N_543,In_775,In_369);
nand U544 (N_544,In_805,In_909);
nor U545 (N_545,In_519,In_489);
and U546 (N_546,In_12,In_46);
nand U547 (N_547,In_180,In_438);
or U548 (N_548,In_819,In_615);
nand U549 (N_549,In_785,In_935);
or U550 (N_550,In_797,In_703);
nor U551 (N_551,In_794,In_65);
nor U552 (N_552,In_560,In_591);
and U553 (N_553,In_239,In_138);
nand U554 (N_554,In_184,In_583);
or U555 (N_555,In_791,In_514);
nand U556 (N_556,In_465,In_151);
and U557 (N_557,In_177,In_561);
or U558 (N_558,In_844,In_260);
or U559 (N_559,In_695,In_318);
nand U560 (N_560,In_290,In_543);
or U561 (N_561,In_474,In_183);
nand U562 (N_562,In_854,In_203);
and U563 (N_563,In_127,In_900);
nor U564 (N_564,In_477,In_530);
or U565 (N_565,In_965,In_769);
nand U566 (N_566,In_90,In_146);
or U567 (N_567,In_483,In_678);
or U568 (N_568,In_212,In_620);
and U569 (N_569,In_653,In_694);
and U570 (N_570,In_591,In_305);
xor U571 (N_571,In_369,In_444);
xnor U572 (N_572,In_869,In_957);
or U573 (N_573,In_371,In_112);
nand U574 (N_574,In_317,In_163);
nor U575 (N_575,In_160,In_667);
nand U576 (N_576,In_9,In_376);
or U577 (N_577,In_963,In_546);
xnor U578 (N_578,In_484,In_306);
and U579 (N_579,In_795,In_720);
and U580 (N_580,In_126,In_832);
and U581 (N_581,In_83,In_867);
or U582 (N_582,In_452,In_883);
and U583 (N_583,In_163,In_840);
or U584 (N_584,In_894,In_853);
nor U585 (N_585,In_24,In_858);
or U586 (N_586,In_56,In_247);
nand U587 (N_587,In_355,In_551);
nand U588 (N_588,In_381,In_482);
nor U589 (N_589,In_865,In_690);
nor U590 (N_590,In_817,In_788);
nor U591 (N_591,In_626,In_737);
nor U592 (N_592,In_447,In_798);
nor U593 (N_593,In_967,In_371);
nand U594 (N_594,In_91,In_34);
or U595 (N_595,In_115,In_222);
nor U596 (N_596,In_835,In_358);
xnor U597 (N_597,In_356,In_919);
or U598 (N_598,In_221,In_178);
nand U599 (N_599,In_763,In_764);
nand U600 (N_600,In_41,In_646);
xor U601 (N_601,In_202,In_360);
or U602 (N_602,In_873,In_648);
or U603 (N_603,In_854,In_295);
and U604 (N_604,In_530,In_266);
nor U605 (N_605,In_483,In_255);
or U606 (N_606,In_278,In_126);
xnor U607 (N_607,In_711,In_563);
or U608 (N_608,In_308,In_402);
or U609 (N_609,In_228,In_331);
and U610 (N_610,In_740,In_80);
or U611 (N_611,In_105,In_998);
xnor U612 (N_612,In_63,In_135);
nand U613 (N_613,In_428,In_433);
and U614 (N_614,In_832,In_203);
xnor U615 (N_615,In_100,In_975);
and U616 (N_616,In_964,In_991);
or U617 (N_617,In_380,In_825);
nor U618 (N_618,In_371,In_760);
nor U619 (N_619,In_965,In_999);
or U620 (N_620,In_59,In_305);
or U621 (N_621,In_824,In_932);
or U622 (N_622,In_558,In_192);
nor U623 (N_623,In_781,In_431);
nand U624 (N_624,In_775,In_215);
or U625 (N_625,In_754,In_44);
xnor U626 (N_626,In_898,In_62);
xor U627 (N_627,In_554,In_930);
or U628 (N_628,In_951,In_402);
nor U629 (N_629,In_777,In_875);
xnor U630 (N_630,In_306,In_143);
or U631 (N_631,In_862,In_424);
or U632 (N_632,In_452,In_644);
and U633 (N_633,In_526,In_926);
or U634 (N_634,In_188,In_499);
or U635 (N_635,In_770,In_909);
nor U636 (N_636,In_664,In_242);
nand U637 (N_637,In_386,In_518);
or U638 (N_638,In_66,In_555);
nor U639 (N_639,In_336,In_381);
and U640 (N_640,In_904,In_390);
or U641 (N_641,In_19,In_563);
xor U642 (N_642,In_164,In_139);
or U643 (N_643,In_202,In_359);
or U644 (N_644,In_287,In_633);
and U645 (N_645,In_877,In_50);
and U646 (N_646,In_463,In_740);
nor U647 (N_647,In_699,In_365);
nand U648 (N_648,In_505,In_787);
and U649 (N_649,In_145,In_393);
or U650 (N_650,In_382,In_431);
and U651 (N_651,In_906,In_434);
and U652 (N_652,In_143,In_137);
and U653 (N_653,In_912,In_518);
or U654 (N_654,In_310,In_815);
nand U655 (N_655,In_933,In_729);
and U656 (N_656,In_31,In_688);
or U657 (N_657,In_779,In_340);
nand U658 (N_658,In_340,In_898);
or U659 (N_659,In_79,In_891);
and U660 (N_660,In_677,In_804);
or U661 (N_661,In_321,In_141);
nor U662 (N_662,In_734,In_595);
and U663 (N_663,In_610,In_186);
and U664 (N_664,In_895,In_587);
and U665 (N_665,In_34,In_27);
nor U666 (N_666,In_274,In_225);
nor U667 (N_667,In_394,In_766);
or U668 (N_668,In_617,In_860);
and U669 (N_669,In_55,In_496);
nor U670 (N_670,In_662,In_30);
or U671 (N_671,In_848,In_657);
xor U672 (N_672,In_486,In_152);
nand U673 (N_673,In_779,In_438);
nand U674 (N_674,In_493,In_22);
xor U675 (N_675,In_78,In_182);
and U676 (N_676,In_858,In_345);
nand U677 (N_677,In_536,In_899);
nand U678 (N_678,In_750,In_338);
nand U679 (N_679,In_561,In_65);
and U680 (N_680,In_648,In_779);
and U681 (N_681,In_521,In_45);
or U682 (N_682,In_447,In_649);
or U683 (N_683,In_15,In_708);
nand U684 (N_684,In_218,In_456);
or U685 (N_685,In_591,In_446);
nand U686 (N_686,In_132,In_300);
and U687 (N_687,In_679,In_884);
and U688 (N_688,In_270,In_207);
and U689 (N_689,In_238,In_919);
nor U690 (N_690,In_637,In_249);
nor U691 (N_691,In_783,In_833);
or U692 (N_692,In_400,In_7);
nor U693 (N_693,In_252,In_328);
nand U694 (N_694,In_989,In_224);
xor U695 (N_695,In_314,In_647);
nor U696 (N_696,In_173,In_268);
or U697 (N_697,In_490,In_617);
or U698 (N_698,In_939,In_964);
or U699 (N_699,In_407,In_490);
nor U700 (N_700,In_802,In_645);
nand U701 (N_701,In_766,In_987);
and U702 (N_702,In_26,In_869);
nor U703 (N_703,In_279,In_183);
or U704 (N_704,In_861,In_708);
nand U705 (N_705,In_985,In_267);
nand U706 (N_706,In_107,In_908);
nor U707 (N_707,In_608,In_993);
xor U708 (N_708,In_866,In_406);
or U709 (N_709,In_392,In_870);
nor U710 (N_710,In_381,In_764);
and U711 (N_711,In_879,In_71);
or U712 (N_712,In_79,In_842);
or U713 (N_713,In_926,In_546);
nand U714 (N_714,In_338,In_729);
nor U715 (N_715,In_902,In_541);
nand U716 (N_716,In_772,In_454);
xnor U717 (N_717,In_231,In_999);
nand U718 (N_718,In_174,In_887);
or U719 (N_719,In_684,In_650);
nor U720 (N_720,In_230,In_948);
nand U721 (N_721,In_904,In_972);
and U722 (N_722,In_363,In_744);
and U723 (N_723,In_898,In_289);
and U724 (N_724,In_64,In_461);
nand U725 (N_725,In_220,In_965);
nand U726 (N_726,In_901,In_750);
nand U727 (N_727,In_640,In_384);
or U728 (N_728,In_413,In_552);
xor U729 (N_729,In_423,In_564);
or U730 (N_730,In_339,In_960);
and U731 (N_731,In_589,In_465);
nor U732 (N_732,In_688,In_517);
or U733 (N_733,In_660,In_801);
or U734 (N_734,In_681,In_651);
xor U735 (N_735,In_724,In_284);
and U736 (N_736,In_932,In_14);
nand U737 (N_737,In_867,In_798);
nor U738 (N_738,In_449,In_487);
nand U739 (N_739,In_972,In_376);
and U740 (N_740,In_542,In_822);
xnor U741 (N_741,In_367,In_812);
nor U742 (N_742,In_810,In_620);
nor U743 (N_743,In_952,In_167);
or U744 (N_744,In_296,In_433);
and U745 (N_745,In_75,In_82);
and U746 (N_746,In_831,In_423);
or U747 (N_747,In_71,In_630);
nor U748 (N_748,In_481,In_703);
and U749 (N_749,In_324,In_958);
xnor U750 (N_750,In_454,In_836);
nor U751 (N_751,In_566,In_103);
and U752 (N_752,In_509,In_158);
nand U753 (N_753,In_898,In_214);
and U754 (N_754,In_389,In_84);
nor U755 (N_755,In_177,In_276);
nand U756 (N_756,In_272,In_751);
nor U757 (N_757,In_811,In_703);
nor U758 (N_758,In_854,In_642);
or U759 (N_759,In_533,In_950);
or U760 (N_760,In_862,In_791);
or U761 (N_761,In_209,In_295);
or U762 (N_762,In_441,In_905);
or U763 (N_763,In_594,In_821);
nor U764 (N_764,In_464,In_858);
nor U765 (N_765,In_521,In_784);
nand U766 (N_766,In_303,In_879);
and U767 (N_767,In_675,In_431);
nand U768 (N_768,In_611,In_673);
and U769 (N_769,In_62,In_699);
or U770 (N_770,In_596,In_427);
and U771 (N_771,In_866,In_312);
or U772 (N_772,In_897,In_286);
nor U773 (N_773,In_446,In_946);
or U774 (N_774,In_560,In_476);
nor U775 (N_775,In_392,In_666);
and U776 (N_776,In_25,In_906);
nor U777 (N_777,In_22,In_291);
and U778 (N_778,In_928,In_418);
or U779 (N_779,In_915,In_490);
nor U780 (N_780,In_863,In_821);
nor U781 (N_781,In_524,In_135);
and U782 (N_782,In_743,In_136);
or U783 (N_783,In_922,In_866);
and U784 (N_784,In_107,In_264);
or U785 (N_785,In_389,In_302);
nor U786 (N_786,In_927,In_797);
and U787 (N_787,In_21,In_90);
and U788 (N_788,In_5,In_415);
and U789 (N_789,In_373,In_860);
or U790 (N_790,In_62,In_737);
nor U791 (N_791,In_495,In_701);
nor U792 (N_792,In_310,In_5);
nand U793 (N_793,In_979,In_230);
nor U794 (N_794,In_88,In_655);
nor U795 (N_795,In_611,In_566);
nand U796 (N_796,In_284,In_823);
nand U797 (N_797,In_54,In_225);
xnor U798 (N_798,In_513,In_382);
and U799 (N_799,In_187,In_393);
or U800 (N_800,In_451,In_134);
and U801 (N_801,In_854,In_159);
nor U802 (N_802,In_576,In_73);
or U803 (N_803,In_926,In_885);
and U804 (N_804,In_798,In_550);
and U805 (N_805,In_94,In_267);
xnor U806 (N_806,In_334,In_29);
nand U807 (N_807,In_242,In_539);
nand U808 (N_808,In_196,In_708);
or U809 (N_809,In_322,In_384);
nor U810 (N_810,In_486,In_329);
nand U811 (N_811,In_201,In_421);
nor U812 (N_812,In_713,In_687);
and U813 (N_813,In_446,In_827);
nor U814 (N_814,In_646,In_155);
nand U815 (N_815,In_640,In_52);
nand U816 (N_816,In_258,In_985);
nand U817 (N_817,In_322,In_57);
and U818 (N_818,In_50,In_230);
and U819 (N_819,In_93,In_976);
and U820 (N_820,In_281,In_15);
nand U821 (N_821,In_757,In_365);
nor U822 (N_822,In_930,In_771);
nand U823 (N_823,In_944,In_480);
xor U824 (N_824,In_743,In_952);
or U825 (N_825,In_577,In_507);
or U826 (N_826,In_840,In_676);
xnor U827 (N_827,In_2,In_745);
and U828 (N_828,In_132,In_67);
and U829 (N_829,In_642,In_460);
nand U830 (N_830,In_732,In_164);
xnor U831 (N_831,In_527,In_321);
nand U832 (N_832,In_174,In_886);
nor U833 (N_833,In_985,In_857);
nor U834 (N_834,In_542,In_890);
nor U835 (N_835,In_442,In_499);
nand U836 (N_836,In_667,In_32);
or U837 (N_837,In_140,In_604);
nor U838 (N_838,In_548,In_97);
nand U839 (N_839,In_304,In_122);
or U840 (N_840,In_249,In_909);
or U841 (N_841,In_749,In_81);
or U842 (N_842,In_808,In_117);
or U843 (N_843,In_646,In_327);
nand U844 (N_844,In_570,In_648);
or U845 (N_845,In_554,In_851);
or U846 (N_846,In_774,In_698);
nand U847 (N_847,In_645,In_392);
nor U848 (N_848,In_695,In_134);
nor U849 (N_849,In_11,In_876);
nand U850 (N_850,In_201,In_362);
or U851 (N_851,In_744,In_409);
xor U852 (N_852,In_205,In_789);
nor U853 (N_853,In_587,In_594);
nand U854 (N_854,In_608,In_760);
nor U855 (N_855,In_18,In_564);
or U856 (N_856,In_631,In_348);
and U857 (N_857,In_123,In_533);
and U858 (N_858,In_743,In_951);
and U859 (N_859,In_657,In_489);
or U860 (N_860,In_913,In_537);
nor U861 (N_861,In_335,In_367);
xor U862 (N_862,In_123,In_199);
and U863 (N_863,In_777,In_472);
or U864 (N_864,In_704,In_396);
nand U865 (N_865,In_470,In_30);
nand U866 (N_866,In_207,In_526);
and U867 (N_867,In_211,In_479);
nor U868 (N_868,In_47,In_340);
nand U869 (N_869,In_412,In_704);
or U870 (N_870,In_495,In_113);
nand U871 (N_871,In_393,In_571);
nor U872 (N_872,In_768,In_38);
and U873 (N_873,In_964,In_526);
nor U874 (N_874,In_775,In_263);
or U875 (N_875,In_904,In_712);
or U876 (N_876,In_857,In_897);
or U877 (N_877,In_917,In_887);
xor U878 (N_878,In_595,In_857);
nand U879 (N_879,In_311,In_144);
or U880 (N_880,In_534,In_388);
nand U881 (N_881,In_337,In_113);
nor U882 (N_882,In_987,In_601);
and U883 (N_883,In_289,In_594);
nor U884 (N_884,In_38,In_431);
nor U885 (N_885,In_627,In_358);
and U886 (N_886,In_677,In_486);
nor U887 (N_887,In_459,In_116);
nor U888 (N_888,In_519,In_425);
nor U889 (N_889,In_506,In_249);
nand U890 (N_890,In_241,In_27);
nand U891 (N_891,In_459,In_690);
and U892 (N_892,In_833,In_612);
or U893 (N_893,In_514,In_669);
nor U894 (N_894,In_857,In_922);
and U895 (N_895,In_221,In_617);
nor U896 (N_896,In_302,In_727);
nand U897 (N_897,In_274,In_848);
nand U898 (N_898,In_792,In_991);
or U899 (N_899,In_496,In_243);
or U900 (N_900,In_332,In_534);
or U901 (N_901,In_151,In_121);
nor U902 (N_902,In_242,In_347);
or U903 (N_903,In_388,In_479);
or U904 (N_904,In_695,In_869);
nor U905 (N_905,In_747,In_494);
nand U906 (N_906,In_620,In_545);
nand U907 (N_907,In_438,In_285);
or U908 (N_908,In_949,In_874);
xnor U909 (N_909,In_63,In_731);
or U910 (N_910,In_852,In_72);
or U911 (N_911,In_528,In_224);
or U912 (N_912,In_372,In_386);
or U913 (N_913,In_833,In_670);
nand U914 (N_914,In_980,In_703);
and U915 (N_915,In_589,In_686);
nand U916 (N_916,In_484,In_575);
nand U917 (N_917,In_700,In_786);
and U918 (N_918,In_594,In_239);
nand U919 (N_919,In_72,In_531);
or U920 (N_920,In_857,In_746);
nor U921 (N_921,In_937,In_197);
and U922 (N_922,In_465,In_140);
nand U923 (N_923,In_832,In_409);
or U924 (N_924,In_397,In_472);
nor U925 (N_925,In_836,In_494);
xnor U926 (N_926,In_554,In_532);
and U927 (N_927,In_74,In_610);
nor U928 (N_928,In_866,In_855);
nor U929 (N_929,In_936,In_539);
xor U930 (N_930,In_78,In_812);
or U931 (N_931,In_662,In_836);
nor U932 (N_932,In_882,In_94);
nor U933 (N_933,In_118,In_428);
nor U934 (N_934,In_791,In_824);
nor U935 (N_935,In_796,In_1);
and U936 (N_936,In_380,In_942);
and U937 (N_937,In_304,In_58);
or U938 (N_938,In_249,In_109);
nand U939 (N_939,In_172,In_761);
or U940 (N_940,In_369,In_429);
or U941 (N_941,In_345,In_881);
nor U942 (N_942,In_768,In_886);
or U943 (N_943,In_282,In_980);
nand U944 (N_944,In_239,In_784);
or U945 (N_945,In_876,In_289);
xnor U946 (N_946,In_515,In_120);
or U947 (N_947,In_637,In_820);
or U948 (N_948,In_127,In_604);
xnor U949 (N_949,In_9,In_261);
nor U950 (N_950,In_443,In_580);
nor U951 (N_951,In_748,In_107);
nor U952 (N_952,In_312,In_889);
xor U953 (N_953,In_881,In_665);
and U954 (N_954,In_434,In_430);
nand U955 (N_955,In_13,In_79);
or U956 (N_956,In_804,In_421);
and U957 (N_957,In_948,In_503);
or U958 (N_958,In_244,In_125);
nor U959 (N_959,In_779,In_806);
or U960 (N_960,In_797,In_65);
xor U961 (N_961,In_310,In_180);
nor U962 (N_962,In_327,In_301);
nor U963 (N_963,In_854,In_959);
and U964 (N_964,In_426,In_958);
nand U965 (N_965,In_217,In_737);
and U966 (N_966,In_451,In_398);
and U967 (N_967,In_624,In_683);
nand U968 (N_968,In_459,In_789);
or U969 (N_969,In_686,In_660);
and U970 (N_970,In_957,In_269);
nand U971 (N_971,In_56,In_330);
or U972 (N_972,In_532,In_327);
nand U973 (N_973,In_131,In_315);
nand U974 (N_974,In_943,In_508);
nor U975 (N_975,In_352,In_149);
nand U976 (N_976,In_663,In_783);
xnor U977 (N_977,In_827,In_247);
xor U978 (N_978,In_646,In_773);
nand U979 (N_979,In_14,In_542);
nand U980 (N_980,In_367,In_283);
and U981 (N_981,In_439,In_430);
and U982 (N_982,In_287,In_947);
nor U983 (N_983,In_463,In_212);
and U984 (N_984,In_725,In_500);
or U985 (N_985,In_451,In_971);
nand U986 (N_986,In_116,In_691);
nand U987 (N_987,In_390,In_221);
and U988 (N_988,In_687,In_670);
and U989 (N_989,In_249,In_924);
xor U990 (N_990,In_157,In_80);
nand U991 (N_991,In_713,In_545);
nand U992 (N_992,In_532,In_273);
or U993 (N_993,In_609,In_24);
and U994 (N_994,In_532,In_51);
and U995 (N_995,In_524,In_610);
nor U996 (N_996,In_825,In_788);
nor U997 (N_997,In_340,In_531);
or U998 (N_998,In_925,In_170);
and U999 (N_999,In_23,In_520);
xor U1000 (N_1000,N_847,N_132);
and U1001 (N_1001,N_771,N_598);
nor U1002 (N_1002,N_407,N_921);
or U1003 (N_1003,N_295,N_7);
and U1004 (N_1004,N_900,N_973);
nand U1005 (N_1005,N_650,N_588);
nand U1006 (N_1006,N_501,N_106);
nor U1007 (N_1007,N_35,N_675);
nand U1008 (N_1008,N_478,N_517);
nor U1009 (N_1009,N_961,N_547);
nand U1010 (N_1010,N_601,N_279);
nand U1011 (N_1011,N_493,N_509);
nand U1012 (N_1012,N_191,N_740);
nor U1013 (N_1013,N_991,N_82);
or U1014 (N_1014,N_880,N_281);
and U1015 (N_1015,N_352,N_895);
nor U1016 (N_1016,N_987,N_248);
nand U1017 (N_1017,N_477,N_275);
and U1018 (N_1018,N_386,N_757);
nand U1019 (N_1019,N_508,N_178);
and U1020 (N_1020,N_765,N_129);
or U1021 (N_1021,N_858,N_676);
and U1022 (N_1022,N_181,N_343);
and U1023 (N_1023,N_773,N_241);
and U1024 (N_1024,N_428,N_375);
or U1025 (N_1025,N_339,N_879);
or U1026 (N_1026,N_750,N_350);
and U1027 (N_1027,N_513,N_671);
and U1028 (N_1028,N_538,N_171);
nand U1029 (N_1029,N_26,N_760);
or U1030 (N_1030,N_716,N_310);
nand U1031 (N_1031,N_977,N_292);
and U1032 (N_1032,N_767,N_460);
or U1033 (N_1033,N_330,N_652);
nand U1034 (N_1034,N_646,N_523);
nand U1035 (N_1035,N_144,N_23);
xnor U1036 (N_1036,N_86,N_368);
or U1037 (N_1037,N_678,N_423);
nand U1038 (N_1038,N_440,N_358);
and U1039 (N_1039,N_79,N_585);
nand U1040 (N_1040,N_974,N_496);
and U1041 (N_1041,N_525,N_134);
and U1042 (N_1042,N_314,N_192);
nor U1043 (N_1043,N_663,N_438);
nor U1044 (N_1044,N_491,N_862);
nand U1045 (N_1045,N_246,N_211);
and U1046 (N_1046,N_833,N_944);
nand U1047 (N_1047,N_50,N_487);
xor U1048 (N_1048,N_69,N_831);
or U1049 (N_1049,N_537,N_532);
xor U1050 (N_1050,N_391,N_571);
or U1051 (N_1051,N_317,N_2);
and U1052 (N_1052,N_115,N_484);
xnor U1053 (N_1053,N_968,N_320);
and U1054 (N_1054,N_872,N_963);
nor U1055 (N_1055,N_693,N_159);
nand U1056 (N_1056,N_296,N_869);
and U1057 (N_1057,N_15,N_27);
nand U1058 (N_1058,N_369,N_175);
xnor U1059 (N_1059,N_566,N_709);
or U1060 (N_1060,N_474,N_836);
or U1061 (N_1061,N_975,N_970);
nand U1062 (N_1062,N_940,N_202);
and U1063 (N_1063,N_575,N_190);
nand U1064 (N_1064,N_146,N_516);
nor U1065 (N_1065,N_626,N_586);
nand U1066 (N_1066,N_432,N_639);
nor U1067 (N_1067,N_848,N_988);
or U1068 (N_1068,N_274,N_955);
or U1069 (N_1069,N_59,N_521);
xnor U1070 (N_1070,N_835,N_867);
nor U1071 (N_1071,N_700,N_12);
nor U1072 (N_1072,N_463,N_374);
nor U1073 (N_1073,N_483,N_128);
or U1074 (N_1074,N_109,N_36);
xor U1075 (N_1075,N_793,N_347);
or U1076 (N_1076,N_567,N_498);
or U1077 (N_1077,N_398,N_897);
and U1078 (N_1078,N_24,N_265);
nand U1079 (N_1079,N_489,N_759);
and U1080 (N_1080,N_683,N_734);
and U1081 (N_1081,N_738,N_906);
xor U1082 (N_1082,N_307,N_136);
and U1083 (N_1083,N_408,N_455);
xor U1084 (N_1084,N_332,N_469);
xor U1085 (N_1085,N_229,N_593);
and U1086 (N_1086,N_643,N_545);
and U1087 (N_1087,N_298,N_31);
nor U1088 (N_1088,N_362,N_666);
nor U1089 (N_1089,N_338,N_905);
nand U1090 (N_1090,N_511,N_9);
nand U1091 (N_1091,N_885,N_889);
or U1092 (N_1092,N_551,N_719);
nand U1093 (N_1093,N_605,N_449);
and U1094 (N_1094,N_637,N_365);
nor U1095 (N_1095,N_874,N_742);
and U1096 (N_1096,N_990,N_454);
or U1097 (N_1097,N_948,N_475);
nand U1098 (N_1098,N_63,N_470);
or U1099 (N_1099,N_183,N_635);
nand U1100 (N_1100,N_66,N_758);
nor U1101 (N_1101,N_770,N_749);
nand U1102 (N_1102,N_435,N_766);
nand U1103 (N_1103,N_62,N_213);
nand U1104 (N_1104,N_964,N_776);
and U1105 (N_1105,N_844,N_592);
nor U1106 (N_1106,N_723,N_558);
xor U1107 (N_1107,N_752,N_792);
nor U1108 (N_1108,N_807,N_284);
or U1109 (N_1109,N_80,N_762);
and U1110 (N_1110,N_779,N_239);
or U1111 (N_1111,N_283,N_473);
nand U1112 (N_1112,N_222,N_941);
nand U1113 (N_1113,N_170,N_708);
nand U1114 (N_1114,N_176,N_240);
or U1115 (N_1115,N_92,N_249);
and U1116 (N_1116,N_777,N_808);
nor U1117 (N_1117,N_390,N_866);
nor U1118 (N_1118,N_913,N_231);
nand U1119 (N_1119,N_813,N_658);
or U1120 (N_1120,N_138,N_821);
nand U1121 (N_1121,N_632,N_465);
and U1122 (N_1122,N_452,N_290);
nand U1123 (N_1123,N_72,N_110);
and U1124 (N_1124,N_647,N_286);
nand U1125 (N_1125,N_490,N_945);
and U1126 (N_1126,N_252,N_361);
and U1127 (N_1127,N_322,N_818);
and U1128 (N_1128,N_817,N_809);
nor U1129 (N_1129,N_805,N_285);
and U1130 (N_1130,N_340,N_837);
nor U1131 (N_1131,N_3,N_662);
xor U1132 (N_1132,N_70,N_495);
nand U1133 (N_1133,N_754,N_325);
or U1134 (N_1134,N_270,N_166);
nand U1135 (N_1135,N_417,N_731);
and U1136 (N_1136,N_989,N_316);
nand U1137 (N_1137,N_367,N_297);
or U1138 (N_1138,N_439,N_238);
nand U1139 (N_1139,N_38,N_868);
nand U1140 (N_1140,N_71,N_604);
nand U1141 (N_1141,N_137,N_370);
and U1142 (N_1142,N_691,N_419);
nor U1143 (N_1143,N_565,N_55);
or U1144 (N_1144,N_4,N_346);
nand U1145 (N_1145,N_729,N_717);
nor U1146 (N_1146,N_242,N_94);
nor U1147 (N_1147,N_881,N_573);
xnor U1148 (N_1148,N_788,N_140);
nor U1149 (N_1149,N_783,N_43);
or U1150 (N_1150,N_780,N_235);
xor U1151 (N_1151,N_851,N_116);
nand U1152 (N_1152,N_834,N_562);
nor U1153 (N_1153,N_706,N_822);
or U1154 (N_1154,N_450,N_642);
nand U1155 (N_1155,N_257,N_896);
or U1156 (N_1156,N_713,N_11);
and U1157 (N_1157,N_486,N_447);
nor U1158 (N_1158,N_617,N_823);
nand U1159 (N_1159,N_506,N_512);
xor U1160 (N_1160,N_707,N_841);
or U1161 (N_1161,N_670,N_621);
nor U1162 (N_1162,N_10,N_445);
nand U1163 (N_1163,N_654,N_425);
nand U1164 (N_1164,N_267,N_595);
nand U1165 (N_1165,N_406,N_113);
nand U1166 (N_1166,N_207,N_306);
or U1167 (N_1167,N_392,N_173);
and U1168 (N_1168,N_378,N_220);
nand U1169 (N_1169,N_324,N_157);
xnor U1170 (N_1170,N_158,N_300);
nor U1171 (N_1171,N_319,N_811);
or U1172 (N_1172,N_411,N_177);
or U1173 (N_1173,N_920,N_388);
nor U1174 (N_1174,N_25,N_755);
xor U1175 (N_1175,N_39,N_19);
xnor U1176 (N_1176,N_978,N_403);
and U1177 (N_1177,N_204,N_364);
and U1178 (N_1178,N_255,N_48);
nor U1179 (N_1179,N_289,N_769);
and U1180 (N_1180,N_58,N_927);
and U1181 (N_1181,N_57,N_739);
xor U1182 (N_1182,N_942,N_276);
nor U1183 (N_1183,N_433,N_100);
and U1184 (N_1184,N_414,N_225);
xor U1185 (N_1185,N_812,N_520);
nor U1186 (N_1186,N_221,N_680);
or U1187 (N_1187,N_745,N_627);
or U1188 (N_1188,N_893,N_429);
or U1189 (N_1189,N_382,N_857);
or U1190 (N_1190,N_278,N_502);
or U1191 (N_1191,N_967,N_29);
nor U1192 (N_1192,N_591,N_568);
or U1193 (N_1193,N_44,N_499);
nor U1194 (N_1194,N_826,N_854);
nand U1195 (N_1195,N_917,N_715);
nor U1196 (N_1196,N_803,N_219);
or U1197 (N_1197,N_665,N_187);
and U1198 (N_1198,N_802,N_272);
nand U1199 (N_1199,N_355,N_957);
nor U1200 (N_1200,N_200,N_54);
or U1201 (N_1201,N_623,N_476);
nand U1202 (N_1202,N_301,N_18);
nand U1203 (N_1203,N_774,N_611);
nand U1204 (N_1204,N_622,N_827);
or U1205 (N_1205,N_795,N_661);
nand U1206 (N_1206,N_539,N_315);
and U1207 (N_1207,N_172,N_702);
nor U1208 (N_1208,N_956,N_97);
nor U1209 (N_1209,N_462,N_609);
nor U1210 (N_1210,N_580,N_442);
nor U1211 (N_1211,N_842,N_32);
nor U1212 (N_1212,N_832,N_481);
and U1213 (N_1213,N_838,N_543);
nor U1214 (N_1214,N_494,N_720);
or U1215 (N_1215,N_799,N_381);
or U1216 (N_1216,N_198,N_466);
and U1217 (N_1217,N_16,N_308);
and U1218 (N_1218,N_559,N_883);
and U1219 (N_1219,N_689,N_946);
nand U1220 (N_1220,N_224,N_724);
or U1221 (N_1221,N_934,N_553);
and U1222 (N_1222,N_633,N_130);
nand U1223 (N_1223,N_856,N_966);
xor U1224 (N_1224,N_142,N_437);
nor U1225 (N_1225,N_886,N_93);
and U1226 (N_1226,N_725,N_864);
nor U1227 (N_1227,N_596,N_215);
or U1228 (N_1228,N_395,N_933);
and U1229 (N_1229,N_163,N_205);
nor U1230 (N_1230,N_563,N_356);
nor U1231 (N_1231,N_925,N_959);
nor U1232 (N_1232,N_540,N_287);
nor U1233 (N_1233,N_935,N_840);
nand U1234 (N_1234,N_684,N_529);
and U1235 (N_1235,N_243,N_519);
xnor U1236 (N_1236,N_131,N_542);
xnor U1237 (N_1237,N_262,N_87);
nor U1238 (N_1238,N_612,N_907);
nand U1239 (N_1239,N_816,N_409);
nand U1240 (N_1240,N_114,N_351);
nand U1241 (N_1241,N_572,N_227);
xnor U1242 (N_1242,N_357,N_51);
or U1243 (N_1243,N_589,N_651);
or U1244 (N_1244,N_263,N_986);
xnor U1245 (N_1245,N_943,N_126);
and U1246 (N_1246,N_534,N_712);
or U1247 (N_1247,N_412,N_504);
and U1248 (N_1248,N_471,N_251);
nand U1249 (N_1249,N_122,N_953);
nor U1250 (N_1250,N_574,N_971);
and U1251 (N_1251,N_149,N_174);
nor U1252 (N_1252,N_960,N_794);
and U1253 (N_1253,N_860,N_898);
nor U1254 (N_1254,N_8,N_620);
or U1255 (N_1255,N_461,N_859);
nor U1256 (N_1256,N_160,N_148);
and U1257 (N_1257,N_640,N_326);
nor U1258 (N_1258,N_522,N_981);
nand U1259 (N_1259,N_839,N_424);
xor U1260 (N_1260,N_787,N_217);
and U1261 (N_1261,N_485,N_74);
nand U1262 (N_1262,N_653,N_746);
or U1263 (N_1263,N_914,N_228);
xnor U1264 (N_1264,N_333,N_107);
nor U1265 (N_1265,N_915,N_656);
or U1266 (N_1266,N_22,N_550);
xnor U1267 (N_1267,N_448,N_353);
nand U1268 (N_1268,N_376,N_150);
nor U1269 (N_1269,N_904,N_902);
xnor U1270 (N_1270,N_711,N_815);
nand U1271 (N_1271,N_825,N_396);
nand U1272 (N_1272,N_732,N_560);
or U1273 (N_1273,N_687,N_954);
nand U1274 (N_1274,N_488,N_664);
or U1275 (N_1275,N_965,N_630);
or U1276 (N_1276,N_806,N_33);
nand U1277 (N_1277,N_120,N_668);
nor U1278 (N_1278,N_726,N_245);
nor U1279 (N_1279,N_727,N_830);
or U1280 (N_1280,N_884,N_692);
nor U1281 (N_1281,N_579,N_518);
and U1282 (N_1282,N_101,N_625);
and U1283 (N_1283,N_983,N_436);
nor U1284 (N_1284,N_309,N_528);
nand U1285 (N_1285,N_819,N_185);
nor U1286 (N_1286,N_446,N_359);
nor U1287 (N_1287,N_548,N_103);
or U1288 (N_1288,N_90,N_434);
and U1289 (N_1289,N_912,N_195);
and U1290 (N_1290,N_697,N_189);
and U1291 (N_1291,N_261,N_634);
nand U1292 (N_1292,N_61,N_682);
and U1293 (N_1293,N_141,N_778);
or U1294 (N_1294,N_418,N_282);
or U1295 (N_1295,N_169,N_401);
nor U1296 (N_1296,N_863,N_570);
nor U1297 (N_1297,N_404,N_569);
nor U1298 (N_1298,N_871,N_196);
nor U1299 (N_1299,N_124,N_852);
and U1300 (N_1300,N_603,N_329);
nand U1301 (N_1301,N_824,N_302);
or U1302 (N_1302,N_464,N_784);
or U1303 (N_1303,N_164,N_952);
or U1304 (N_1304,N_197,N_894);
or U1305 (N_1305,N_413,N_613);
nand U1306 (N_1306,N_344,N_781);
nand U1307 (N_1307,N_610,N_405);
nor U1308 (N_1308,N_53,N_936);
nor U1309 (N_1309,N_797,N_703);
and U1310 (N_1310,N_667,N_919);
or U1311 (N_1311,N_76,N_162);
nor U1312 (N_1312,N_645,N_372);
nor U1313 (N_1313,N_363,N_422);
xor U1314 (N_1314,N_695,N_236);
or U1315 (N_1315,N_273,N_736);
or U1316 (N_1316,N_145,N_212);
nor U1317 (N_1317,N_600,N_996);
nor U1318 (N_1318,N_312,N_800);
or U1319 (N_1319,N_785,N_599);
or U1320 (N_1320,N_584,N_354);
and U1321 (N_1321,N_334,N_379);
nand U1322 (N_1322,N_139,N_976);
and U1323 (N_1323,N_349,N_648);
nand U1324 (N_1324,N_741,N_546);
xor U1325 (N_1325,N_660,N_688);
nor U1326 (N_1326,N_744,N_323);
nor U1327 (N_1327,N_533,N_108);
or U1328 (N_1328,N_577,N_421);
nand U1329 (N_1329,N_397,N_638);
nand U1330 (N_1330,N_237,N_81);
or U1331 (N_1331,N_135,N_524);
and U1332 (N_1332,N_47,N_56);
and U1333 (N_1333,N_756,N_250);
and U1334 (N_1334,N_582,N_234);
and U1335 (N_1335,N_728,N_321);
nor U1336 (N_1336,N_557,N_467);
nor U1337 (N_1337,N_28,N_345);
nand U1338 (N_1338,N_256,N_194);
and U1339 (N_1339,N_468,N_718);
or U1340 (N_1340,N_394,N_336);
xor U1341 (N_1341,N_444,N_969);
nor U1342 (N_1342,N_208,N_606);
nand U1343 (N_1343,N_510,N_430);
nor U1344 (N_1344,N_628,N_427);
nor U1345 (N_1345,N_861,N_210);
nor U1346 (N_1346,N_400,N_125);
and U1347 (N_1347,N_153,N_655);
xnor U1348 (N_1348,N_52,N_167);
nand U1349 (N_1349,N_143,N_313);
or U1350 (N_1350,N_916,N_73);
nor U1351 (N_1351,N_698,N_541);
and U1352 (N_1352,N_791,N_188);
and U1353 (N_1353,N_747,N_458);
or U1354 (N_1354,N_865,N_119);
and U1355 (N_1355,N_492,N_615);
nand U1356 (N_1356,N_253,N_796);
nor U1357 (N_1357,N_266,N_83);
and U1358 (N_1358,N_931,N_891);
nor U1359 (N_1359,N_223,N_121);
xor U1360 (N_1360,N_393,N_932);
nand U1361 (N_1361,N_133,N_385);
nor U1362 (N_1362,N_280,N_994);
and U1363 (N_1363,N_980,N_152);
or U1364 (N_1364,N_514,N_288);
and U1365 (N_1365,N_89,N_118);
or U1366 (N_1366,N_14,N_992);
or U1367 (N_1367,N_939,N_46);
nand U1368 (N_1368,N_503,N_68);
nor U1369 (N_1369,N_201,N_705);
or U1370 (N_1370,N_426,N_922);
and U1371 (N_1371,N_318,N_993);
nand U1372 (N_1372,N_649,N_305);
or U1373 (N_1373,N_6,N_673);
and U1374 (N_1374,N_371,N_843);
and U1375 (N_1375,N_764,N_686);
nand U1376 (N_1376,N_619,N_576);
nand U1377 (N_1377,N_497,N_938);
nor U1378 (N_1378,N_387,N_772);
nor U1379 (N_1379,N_979,N_402);
and U1380 (N_1380,N_578,N_416);
nand U1381 (N_1381,N_636,N_342);
nand U1382 (N_1382,N_214,N_230);
xor U1383 (N_1383,N_768,N_327);
and U1384 (N_1384,N_685,N_694);
nand U1385 (N_1385,N_184,N_679);
nand U1386 (N_1386,N_453,N_311);
nand U1387 (N_1387,N_155,N_882);
nand U1388 (N_1388,N_722,N_681);
and U1389 (N_1389,N_65,N_982);
nand U1390 (N_1390,N_929,N_875);
and U1391 (N_1391,N_677,N_264);
and U1392 (N_1392,N_853,N_701);
nand U1393 (N_1393,N_730,N_45);
and U1394 (N_1394,N_899,N_618);
or U1395 (N_1395,N_151,N_218);
xnor U1396 (N_1396,N_870,N_226);
nand U1397 (N_1397,N_180,N_104);
or U1398 (N_1398,N_696,N_49);
nand U1399 (N_1399,N_587,N_5);
and U1400 (N_1400,N_377,N_482);
nand U1401 (N_1401,N_798,N_761);
or U1402 (N_1402,N_549,N_737);
nor U1403 (N_1403,N_810,N_99);
nor U1404 (N_1404,N_244,N_735);
and U1405 (N_1405,N_34,N_674);
and U1406 (N_1406,N_583,N_530);
nor U1407 (N_1407,N_556,N_304);
xor U1408 (N_1408,N_850,N_294);
nor U1409 (N_1409,N_457,N_105);
nand U1410 (N_1410,N_233,N_947);
nand U1411 (N_1411,N_958,N_303);
or U1412 (N_1412,N_456,N_254);
nor U1413 (N_1413,N_877,N_67);
nand U1414 (N_1414,N_98,N_814);
or U1415 (N_1415,N_64,N_182);
or U1416 (N_1416,N_951,N_607);
nor U1417 (N_1417,N_179,N_552);
nor U1418 (N_1418,N_930,N_928);
xor U1419 (N_1419,N_804,N_908);
and U1420 (N_1420,N_876,N_845);
or U1421 (N_1421,N_828,N_112);
and U1422 (N_1422,N_641,N_561);
nor U1423 (N_1423,N_892,N_1);
xor U1424 (N_1424,N_209,N_995);
or U1425 (N_1425,N_88,N_581);
nand U1426 (N_1426,N_614,N_366);
and U1427 (N_1427,N_984,N_926);
and U1428 (N_1428,N_998,N_111);
and U1429 (N_1429,N_84,N_710);
or U1430 (N_1430,N_335,N_507);
or U1431 (N_1431,N_269,N_629);
and U1432 (N_1432,N_78,N_41);
or U1433 (N_1433,N_594,N_399);
nand U1434 (N_1434,N_75,N_554);
nor U1435 (N_1435,N_505,N_901);
or U1436 (N_1436,N_360,N_997);
xor U1437 (N_1437,N_268,N_602);
or U1438 (N_1438,N_743,N_555);
nor U1439 (N_1439,N_431,N_690);
and U1440 (N_1440,N_659,N_515);
nand U1441 (N_1441,N_751,N_985);
nor U1442 (N_1442,N_888,N_937);
and U1443 (N_1443,N_704,N_373);
nand U1444 (N_1444,N_293,N_216);
or U1445 (N_1445,N_500,N_672);
nor U1446 (N_1446,N_443,N_910);
or U1447 (N_1447,N_42,N_631);
nor U1448 (N_1448,N_855,N_829);
nor U1449 (N_1449,N_535,N_60);
xor U1450 (N_1450,N_247,N_161);
nand U1451 (N_1451,N_203,N_410);
nand U1452 (N_1452,N_102,N_873);
xnor U1453 (N_1453,N_564,N_260);
or U1454 (N_1454,N_123,N_790);
xor U1455 (N_1455,N_962,N_590);
and U1456 (N_1456,N_232,N_949);
or U1457 (N_1457,N_472,N_801);
xor U1458 (N_1458,N_348,N_903);
and U1459 (N_1459,N_753,N_384);
xor U1460 (N_1460,N_331,N_782);
nor U1461 (N_1461,N_480,N_459);
or U1462 (N_1462,N_616,N_117);
or U1463 (N_1463,N_714,N_156);
nor U1464 (N_1464,N_91,N_299);
nand U1465 (N_1465,N_40,N_748);
or U1466 (N_1466,N_918,N_337);
and U1467 (N_1467,N_789,N_544);
nor U1468 (N_1468,N_20,N_96);
or U1469 (N_1469,N_291,N_186);
nand U1470 (N_1470,N_657,N_154);
and U1471 (N_1471,N_820,N_950);
nand U1472 (N_1472,N_441,N_341);
nand U1473 (N_1473,N_624,N_999);
nor U1474 (N_1474,N_206,N_911);
or U1475 (N_1475,N_597,N_644);
nand U1476 (N_1476,N_531,N_127);
and U1477 (N_1477,N_147,N_380);
nor U1478 (N_1478,N_890,N_699);
nand U1479 (N_1479,N_85,N_849);
or U1480 (N_1480,N_30,N_193);
and U1481 (N_1481,N_763,N_17);
and U1482 (N_1482,N_95,N_271);
nor U1483 (N_1483,N_526,N_878);
xor U1484 (N_1484,N_258,N_13);
and U1485 (N_1485,N_479,N_923);
nor U1486 (N_1486,N_37,N_846);
and U1487 (N_1487,N_415,N_972);
or U1488 (N_1488,N_608,N_199);
and U1489 (N_1489,N_786,N_527);
and U1490 (N_1490,N_328,N_21);
and U1491 (N_1491,N_536,N_669);
nor U1492 (N_1492,N_0,N_451);
or U1493 (N_1493,N_277,N_721);
nand U1494 (N_1494,N_389,N_887);
and U1495 (N_1495,N_775,N_259);
xor U1496 (N_1496,N_77,N_924);
nand U1497 (N_1497,N_733,N_165);
or U1498 (N_1498,N_420,N_909);
or U1499 (N_1499,N_168,N_383);
nand U1500 (N_1500,N_601,N_319);
or U1501 (N_1501,N_362,N_35);
and U1502 (N_1502,N_464,N_831);
and U1503 (N_1503,N_482,N_263);
or U1504 (N_1504,N_251,N_838);
and U1505 (N_1505,N_393,N_97);
nand U1506 (N_1506,N_163,N_723);
and U1507 (N_1507,N_941,N_946);
nand U1508 (N_1508,N_749,N_136);
nand U1509 (N_1509,N_388,N_831);
nand U1510 (N_1510,N_519,N_23);
nand U1511 (N_1511,N_295,N_138);
or U1512 (N_1512,N_967,N_794);
or U1513 (N_1513,N_114,N_111);
nand U1514 (N_1514,N_204,N_932);
or U1515 (N_1515,N_968,N_12);
xor U1516 (N_1516,N_329,N_190);
nand U1517 (N_1517,N_481,N_45);
and U1518 (N_1518,N_139,N_670);
nor U1519 (N_1519,N_680,N_984);
and U1520 (N_1520,N_607,N_771);
nand U1521 (N_1521,N_823,N_57);
nand U1522 (N_1522,N_876,N_175);
nor U1523 (N_1523,N_542,N_501);
nor U1524 (N_1524,N_309,N_13);
nor U1525 (N_1525,N_184,N_812);
nor U1526 (N_1526,N_658,N_517);
and U1527 (N_1527,N_297,N_959);
and U1528 (N_1528,N_494,N_958);
or U1529 (N_1529,N_693,N_664);
nor U1530 (N_1530,N_938,N_848);
nand U1531 (N_1531,N_705,N_260);
or U1532 (N_1532,N_927,N_192);
nand U1533 (N_1533,N_202,N_449);
nand U1534 (N_1534,N_71,N_241);
or U1535 (N_1535,N_559,N_343);
or U1536 (N_1536,N_212,N_835);
nor U1537 (N_1537,N_998,N_513);
nor U1538 (N_1538,N_610,N_501);
and U1539 (N_1539,N_543,N_653);
nor U1540 (N_1540,N_296,N_365);
and U1541 (N_1541,N_377,N_955);
nand U1542 (N_1542,N_440,N_139);
nand U1543 (N_1543,N_319,N_181);
xor U1544 (N_1544,N_915,N_590);
nand U1545 (N_1545,N_951,N_80);
nor U1546 (N_1546,N_821,N_481);
and U1547 (N_1547,N_104,N_677);
xnor U1548 (N_1548,N_859,N_823);
nand U1549 (N_1549,N_271,N_997);
or U1550 (N_1550,N_188,N_117);
and U1551 (N_1551,N_920,N_206);
nand U1552 (N_1552,N_190,N_394);
or U1553 (N_1553,N_23,N_857);
nor U1554 (N_1554,N_326,N_452);
nor U1555 (N_1555,N_717,N_778);
nor U1556 (N_1556,N_804,N_912);
and U1557 (N_1557,N_615,N_858);
xnor U1558 (N_1558,N_42,N_803);
and U1559 (N_1559,N_366,N_34);
nor U1560 (N_1560,N_51,N_467);
or U1561 (N_1561,N_210,N_965);
and U1562 (N_1562,N_936,N_266);
and U1563 (N_1563,N_167,N_825);
nor U1564 (N_1564,N_762,N_274);
nor U1565 (N_1565,N_515,N_549);
or U1566 (N_1566,N_18,N_705);
xnor U1567 (N_1567,N_938,N_121);
and U1568 (N_1568,N_198,N_962);
nor U1569 (N_1569,N_782,N_399);
and U1570 (N_1570,N_919,N_202);
or U1571 (N_1571,N_157,N_46);
xnor U1572 (N_1572,N_792,N_465);
nor U1573 (N_1573,N_466,N_495);
nand U1574 (N_1574,N_540,N_519);
or U1575 (N_1575,N_885,N_816);
nor U1576 (N_1576,N_528,N_108);
and U1577 (N_1577,N_170,N_522);
and U1578 (N_1578,N_286,N_797);
or U1579 (N_1579,N_162,N_35);
nand U1580 (N_1580,N_159,N_859);
or U1581 (N_1581,N_14,N_311);
nor U1582 (N_1582,N_360,N_49);
xnor U1583 (N_1583,N_888,N_799);
and U1584 (N_1584,N_168,N_15);
nand U1585 (N_1585,N_477,N_622);
or U1586 (N_1586,N_492,N_393);
and U1587 (N_1587,N_313,N_196);
or U1588 (N_1588,N_187,N_218);
nor U1589 (N_1589,N_178,N_531);
or U1590 (N_1590,N_147,N_95);
xor U1591 (N_1591,N_357,N_110);
and U1592 (N_1592,N_205,N_553);
xnor U1593 (N_1593,N_339,N_407);
xnor U1594 (N_1594,N_568,N_442);
nand U1595 (N_1595,N_576,N_243);
and U1596 (N_1596,N_28,N_108);
nand U1597 (N_1597,N_380,N_839);
and U1598 (N_1598,N_724,N_321);
and U1599 (N_1599,N_273,N_944);
and U1600 (N_1600,N_489,N_182);
or U1601 (N_1601,N_396,N_690);
xnor U1602 (N_1602,N_524,N_774);
and U1603 (N_1603,N_216,N_16);
or U1604 (N_1604,N_538,N_774);
nand U1605 (N_1605,N_991,N_322);
nand U1606 (N_1606,N_587,N_367);
xnor U1607 (N_1607,N_177,N_812);
nand U1608 (N_1608,N_764,N_309);
nand U1609 (N_1609,N_74,N_315);
nor U1610 (N_1610,N_544,N_444);
or U1611 (N_1611,N_580,N_69);
nor U1612 (N_1612,N_72,N_334);
or U1613 (N_1613,N_454,N_2);
nand U1614 (N_1614,N_41,N_569);
or U1615 (N_1615,N_962,N_949);
and U1616 (N_1616,N_684,N_106);
or U1617 (N_1617,N_424,N_259);
or U1618 (N_1618,N_12,N_476);
nand U1619 (N_1619,N_729,N_967);
xor U1620 (N_1620,N_662,N_638);
nand U1621 (N_1621,N_881,N_541);
or U1622 (N_1622,N_514,N_437);
or U1623 (N_1623,N_755,N_220);
nor U1624 (N_1624,N_836,N_697);
and U1625 (N_1625,N_420,N_79);
or U1626 (N_1626,N_520,N_811);
or U1627 (N_1627,N_129,N_157);
nor U1628 (N_1628,N_737,N_692);
nand U1629 (N_1629,N_705,N_757);
and U1630 (N_1630,N_282,N_722);
xor U1631 (N_1631,N_156,N_12);
nor U1632 (N_1632,N_296,N_379);
xor U1633 (N_1633,N_459,N_386);
xor U1634 (N_1634,N_295,N_808);
and U1635 (N_1635,N_738,N_24);
and U1636 (N_1636,N_206,N_416);
nand U1637 (N_1637,N_851,N_533);
and U1638 (N_1638,N_953,N_124);
nand U1639 (N_1639,N_875,N_498);
xor U1640 (N_1640,N_721,N_994);
or U1641 (N_1641,N_874,N_461);
or U1642 (N_1642,N_572,N_243);
nand U1643 (N_1643,N_752,N_398);
and U1644 (N_1644,N_604,N_721);
nand U1645 (N_1645,N_794,N_205);
nand U1646 (N_1646,N_756,N_418);
and U1647 (N_1647,N_644,N_73);
and U1648 (N_1648,N_768,N_526);
nor U1649 (N_1649,N_650,N_348);
or U1650 (N_1650,N_919,N_613);
nor U1651 (N_1651,N_793,N_521);
and U1652 (N_1652,N_892,N_49);
and U1653 (N_1653,N_545,N_682);
nand U1654 (N_1654,N_665,N_206);
xnor U1655 (N_1655,N_38,N_828);
nand U1656 (N_1656,N_829,N_562);
nor U1657 (N_1657,N_592,N_197);
nand U1658 (N_1658,N_674,N_442);
xor U1659 (N_1659,N_550,N_706);
nor U1660 (N_1660,N_34,N_877);
nand U1661 (N_1661,N_836,N_517);
nor U1662 (N_1662,N_958,N_968);
nor U1663 (N_1663,N_312,N_872);
nand U1664 (N_1664,N_641,N_858);
or U1665 (N_1665,N_691,N_953);
xor U1666 (N_1666,N_664,N_57);
nand U1667 (N_1667,N_160,N_343);
nor U1668 (N_1668,N_521,N_547);
or U1669 (N_1669,N_827,N_419);
nor U1670 (N_1670,N_497,N_770);
or U1671 (N_1671,N_7,N_802);
nand U1672 (N_1672,N_568,N_893);
nand U1673 (N_1673,N_867,N_154);
and U1674 (N_1674,N_762,N_118);
or U1675 (N_1675,N_281,N_977);
and U1676 (N_1676,N_768,N_810);
or U1677 (N_1677,N_70,N_822);
nor U1678 (N_1678,N_114,N_246);
and U1679 (N_1679,N_282,N_155);
and U1680 (N_1680,N_432,N_655);
nand U1681 (N_1681,N_576,N_85);
nand U1682 (N_1682,N_71,N_772);
or U1683 (N_1683,N_610,N_561);
or U1684 (N_1684,N_954,N_525);
nand U1685 (N_1685,N_584,N_263);
nor U1686 (N_1686,N_690,N_267);
nor U1687 (N_1687,N_641,N_703);
nor U1688 (N_1688,N_121,N_769);
nor U1689 (N_1689,N_195,N_979);
or U1690 (N_1690,N_185,N_167);
and U1691 (N_1691,N_123,N_926);
and U1692 (N_1692,N_212,N_467);
nor U1693 (N_1693,N_677,N_444);
or U1694 (N_1694,N_828,N_631);
xor U1695 (N_1695,N_887,N_259);
and U1696 (N_1696,N_243,N_127);
nor U1697 (N_1697,N_82,N_928);
nor U1698 (N_1698,N_5,N_265);
and U1699 (N_1699,N_338,N_5);
or U1700 (N_1700,N_73,N_231);
or U1701 (N_1701,N_550,N_501);
nand U1702 (N_1702,N_382,N_186);
and U1703 (N_1703,N_864,N_699);
or U1704 (N_1704,N_561,N_482);
and U1705 (N_1705,N_780,N_510);
and U1706 (N_1706,N_953,N_734);
nand U1707 (N_1707,N_743,N_277);
and U1708 (N_1708,N_429,N_505);
nand U1709 (N_1709,N_241,N_996);
xnor U1710 (N_1710,N_685,N_64);
and U1711 (N_1711,N_80,N_932);
or U1712 (N_1712,N_643,N_689);
or U1713 (N_1713,N_245,N_8);
and U1714 (N_1714,N_778,N_900);
nand U1715 (N_1715,N_636,N_338);
nor U1716 (N_1716,N_178,N_417);
and U1717 (N_1717,N_477,N_493);
nor U1718 (N_1718,N_13,N_954);
and U1719 (N_1719,N_728,N_328);
and U1720 (N_1720,N_230,N_323);
xor U1721 (N_1721,N_539,N_908);
nor U1722 (N_1722,N_32,N_632);
and U1723 (N_1723,N_655,N_781);
xnor U1724 (N_1724,N_102,N_999);
or U1725 (N_1725,N_516,N_544);
and U1726 (N_1726,N_305,N_578);
nand U1727 (N_1727,N_678,N_758);
xnor U1728 (N_1728,N_328,N_552);
and U1729 (N_1729,N_200,N_384);
xor U1730 (N_1730,N_395,N_403);
nand U1731 (N_1731,N_733,N_710);
nor U1732 (N_1732,N_28,N_609);
or U1733 (N_1733,N_577,N_429);
and U1734 (N_1734,N_834,N_501);
and U1735 (N_1735,N_67,N_693);
and U1736 (N_1736,N_58,N_906);
and U1737 (N_1737,N_690,N_337);
and U1738 (N_1738,N_458,N_4);
or U1739 (N_1739,N_265,N_842);
nor U1740 (N_1740,N_541,N_394);
nor U1741 (N_1741,N_410,N_403);
nor U1742 (N_1742,N_388,N_123);
nor U1743 (N_1743,N_697,N_528);
nand U1744 (N_1744,N_606,N_73);
nor U1745 (N_1745,N_275,N_995);
and U1746 (N_1746,N_210,N_148);
nor U1747 (N_1747,N_910,N_112);
nor U1748 (N_1748,N_997,N_267);
or U1749 (N_1749,N_540,N_642);
nor U1750 (N_1750,N_395,N_851);
and U1751 (N_1751,N_34,N_839);
nor U1752 (N_1752,N_157,N_921);
nand U1753 (N_1753,N_926,N_702);
nor U1754 (N_1754,N_722,N_303);
nor U1755 (N_1755,N_239,N_894);
nand U1756 (N_1756,N_840,N_918);
nor U1757 (N_1757,N_812,N_59);
nor U1758 (N_1758,N_470,N_862);
and U1759 (N_1759,N_654,N_749);
or U1760 (N_1760,N_118,N_178);
nor U1761 (N_1761,N_238,N_295);
or U1762 (N_1762,N_997,N_928);
or U1763 (N_1763,N_387,N_613);
nor U1764 (N_1764,N_960,N_396);
and U1765 (N_1765,N_658,N_170);
or U1766 (N_1766,N_241,N_613);
xor U1767 (N_1767,N_98,N_726);
nor U1768 (N_1768,N_199,N_650);
nor U1769 (N_1769,N_110,N_522);
and U1770 (N_1770,N_929,N_589);
or U1771 (N_1771,N_822,N_68);
or U1772 (N_1772,N_293,N_367);
nand U1773 (N_1773,N_978,N_188);
nor U1774 (N_1774,N_514,N_799);
or U1775 (N_1775,N_622,N_931);
nand U1776 (N_1776,N_202,N_330);
or U1777 (N_1777,N_11,N_449);
nor U1778 (N_1778,N_492,N_767);
or U1779 (N_1779,N_275,N_156);
or U1780 (N_1780,N_778,N_689);
or U1781 (N_1781,N_868,N_779);
nor U1782 (N_1782,N_306,N_5);
and U1783 (N_1783,N_509,N_31);
nand U1784 (N_1784,N_970,N_855);
nand U1785 (N_1785,N_907,N_147);
and U1786 (N_1786,N_590,N_874);
nor U1787 (N_1787,N_958,N_376);
nor U1788 (N_1788,N_575,N_268);
nor U1789 (N_1789,N_662,N_288);
nor U1790 (N_1790,N_921,N_728);
nand U1791 (N_1791,N_747,N_530);
or U1792 (N_1792,N_376,N_887);
nand U1793 (N_1793,N_847,N_240);
and U1794 (N_1794,N_75,N_653);
and U1795 (N_1795,N_575,N_208);
nand U1796 (N_1796,N_680,N_295);
nand U1797 (N_1797,N_451,N_710);
nor U1798 (N_1798,N_154,N_386);
nand U1799 (N_1799,N_231,N_527);
and U1800 (N_1800,N_478,N_922);
or U1801 (N_1801,N_564,N_159);
or U1802 (N_1802,N_116,N_258);
nand U1803 (N_1803,N_848,N_980);
nor U1804 (N_1804,N_80,N_56);
or U1805 (N_1805,N_888,N_406);
or U1806 (N_1806,N_800,N_713);
or U1807 (N_1807,N_821,N_547);
or U1808 (N_1808,N_304,N_843);
and U1809 (N_1809,N_507,N_731);
nand U1810 (N_1810,N_849,N_362);
and U1811 (N_1811,N_145,N_771);
nand U1812 (N_1812,N_404,N_522);
nand U1813 (N_1813,N_196,N_934);
xnor U1814 (N_1814,N_40,N_636);
nor U1815 (N_1815,N_251,N_358);
and U1816 (N_1816,N_784,N_124);
xor U1817 (N_1817,N_19,N_121);
and U1818 (N_1818,N_28,N_142);
xnor U1819 (N_1819,N_648,N_860);
or U1820 (N_1820,N_668,N_866);
nand U1821 (N_1821,N_487,N_427);
and U1822 (N_1822,N_18,N_834);
or U1823 (N_1823,N_232,N_716);
nand U1824 (N_1824,N_386,N_742);
or U1825 (N_1825,N_67,N_946);
or U1826 (N_1826,N_539,N_996);
nor U1827 (N_1827,N_652,N_16);
and U1828 (N_1828,N_645,N_711);
and U1829 (N_1829,N_581,N_870);
nand U1830 (N_1830,N_29,N_355);
or U1831 (N_1831,N_251,N_918);
xor U1832 (N_1832,N_829,N_512);
xnor U1833 (N_1833,N_326,N_592);
or U1834 (N_1834,N_173,N_753);
nand U1835 (N_1835,N_706,N_650);
nor U1836 (N_1836,N_604,N_276);
or U1837 (N_1837,N_556,N_77);
nor U1838 (N_1838,N_229,N_143);
nand U1839 (N_1839,N_218,N_657);
and U1840 (N_1840,N_438,N_570);
and U1841 (N_1841,N_691,N_391);
xnor U1842 (N_1842,N_609,N_965);
nand U1843 (N_1843,N_313,N_147);
or U1844 (N_1844,N_230,N_365);
nand U1845 (N_1845,N_378,N_151);
and U1846 (N_1846,N_638,N_619);
and U1847 (N_1847,N_490,N_102);
or U1848 (N_1848,N_766,N_380);
and U1849 (N_1849,N_787,N_775);
nand U1850 (N_1850,N_531,N_618);
and U1851 (N_1851,N_95,N_495);
or U1852 (N_1852,N_539,N_339);
nor U1853 (N_1853,N_742,N_215);
or U1854 (N_1854,N_330,N_725);
and U1855 (N_1855,N_12,N_685);
nor U1856 (N_1856,N_282,N_947);
nand U1857 (N_1857,N_834,N_973);
or U1858 (N_1858,N_292,N_664);
or U1859 (N_1859,N_663,N_220);
nand U1860 (N_1860,N_253,N_826);
and U1861 (N_1861,N_208,N_632);
nand U1862 (N_1862,N_290,N_876);
xor U1863 (N_1863,N_758,N_789);
nor U1864 (N_1864,N_819,N_209);
and U1865 (N_1865,N_387,N_299);
nor U1866 (N_1866,N_733,N_573);
xor U1867 (N_1867,N_514,N_440);
nor U1868 (N_1868,N_111,N_7);
and U1869 (N_1869,N_145,N_493);
or U1870 (N_1870,N_842,N_529);
xnor U1871 (N_1871,N_936,N_140);
nor U1872 (N_1872,N_411,N_412);
and U1873 (N_1873,N_416,N_767);
or U1874 (N_1874,N_782,N_846);
and U1875 (N_1875,N_833,N_410);
nand U1876 (N_1876,N_943,N_119);
nor U1877 (N_1877,N_27,N_601);
nor U1878 (N_1878,N_782,N_838);
or U1879 (N_1879,N_402,N_120);
nand U1880 (N_1880,N_606,N_739);
xnor U1881 (N_1881,N_557,N_155);
and U1882 (N_1882,N_27,N_315);
xor U1883 (N_1883,N_44,N_921);
and U1884 (N_1884,N_568,N_260);
nor U1885 (N_1885,N_689,N_427);
and U1886 (N_1886,N_987,N_107);
and U1887 (N_1887,N_764,N_317);
nand U1888 (N_1888,N_280,N_875);
nand U1889 (N_1889,N_352,N_854);
nand U1890 (N_1890,N_512,N_501);
and U1891 (N_1891,N_3,N_688);
and U1892 (N_1892,N_485,N_953);
nand U1893 (N_1893,N_75,N_882);
xor U1894 (N_1894,N_805,N_929);
or U1895 (N_1895,N_382,N_19);
nor U1896 (N_1896,N_332,N_732);
nand U1897 (N_1897,N_407,N_90);
nand U1898 (N_1898,N_78,N_659);
and U1899 (N_1899,N_767,N_750);
or U1900 (N_1900,N_45,N_378);
xnor U1901 (N_1901,N_647,N_549);
nor U1902 (N_1902,N_114,N_504);
nand U1903 (N_1903,N_781,N_580);
nor U1904 (N_1904,N_173,N_608);
nor U1905 (N_1905,N_185,N_511);
or U1906 (N_1906,N_739,N_292);
and U1907 (N_1907,N_382,N_457);
xor U1908 (N_1908,N_283,N_310);
and U1909 (N_1909,N_922,N_975);
nor U1910 (N_1910,N_492,N_713);
nand U1911 (N_1911,N_191,N_492);
or U1912 (N_1912,N_92,N_379);
or U1913 (N_1913,N_957,N_484);
nand U1914 (N_1914,N_528,N_541);
xnor U1915 (N_1915,N_753,N_286);
nand U1916 (N_1916,N_514,N_712);
and U1917 (N_1917,N_709,N_25);
and U1918 (N_1918,N_668,N_355);
nand U1919 (N_1919,N_65,N_252);
or U1920 (N_1920,N_510,N_805);
nor U1921 (N_1921,N_357,N_703);
and U1922 (N_1922,N_764,N_419);
and U1923 (N_1923,N_643,N_594);
or U1924 (N_1924,N_828,N_676);
and U1925 (N_1925,N_674,N_301);
or U1926 (N_1926,N_657,N_446);
xnor U1927 (N_1927,N_237,N_819);
or U1928 (N_1928,N_78,N_746);
nand U1929 (N_1929,N_989,N_209);
nor U1930 (N_1930,N_722,N_737);
nor U1931 (N_1931,N_142,N_654);
and U1932 (N_1932,N_297,N_456);
nand U1933 (N_1933,N_455,N_451);
and U1934 (N_1934,N_762,N_212);
xnor U1935 (N_1935,N_194,N_191);
and U1936 (N_1936,N_63,N_475);
nor U1937 (N_1937,N_322,N_797);
or U1938 (N_1938,N_991,N_856);
and U1939 (N_1939,N_468,N_682);
nor U1940 (N_1940,N_439,N_200);
and U1941 (N_1941,N_167,N_10);
or U1942 (N_1942,N_267,N_557);
nor U1943 (N_1943,N_567,N_527);
and U1944 (N_1944,N_295,N_512);
and U1945 (N_1945,N_683,N_377);
nor U1946 (N_1946,N_266,N_972);
nand U1947 (N_1947,N_804,N_91);
and U1948 (N_1948,N_751,N_512);
xor U1949 (N_1949,N_612,N_798);
nand U1950 (N_1950,N_889,N_48);
nand U1951 (N_1951,N_63,N_992);
and U1952 (N_1952,N_383,N_286);
nand U1953 (N_1953,N_743,N_585);
and U1954 (N_1954,N_758,N_204);
or U1955 (N_1955,N_628,N_491);
nand U1956 (N_1956,N_529,N_16);
xnor U1957 (N_1957,N_38,N_692);
or U1958 (N_1958,N_410,N_606);
nand U1959 (N_1959,N_809,N_517);
nand U1960 (N_1960,N_615,N_547);
nor U1961 (N_1961,N_111,N_688);
nor U1962 (N_1962,N_914,N_34);
or U1963 (N_1963,N_627,N_597);
nand U1964 (N_1964,N_161,N_578);
and U1965 (N_1965,N_682,N_139);
nand U1966 (N_1966,N_746,N_9);
and U1967 (N_1967,N_100,N_806);
nor U1968 (N_1968,N_149,N_689);
and U1969 (N_1969,N_614,N_914);
or U1970 (N_1970,N_919,N_906);
nand U1971 (N_1971,N_524,N_852);
or U1972 (N_1972,N_452,N_87);
and U1973 (N_1973,N_919,N_501);
or U1974 (N_1974,N_15,N_643);
nand U1975 (N_1975,N_121,N_271);
nor U1976 (N_1976,N_304,N_788);
nand U1977 (N_1977,N_657,N_462);
or U1978 (N_1978,N_81,N_882);
xnor U1979 (N_1979,N_242,N_98);
xnor U1980 (N_1980,N_940,N_412);
xnor U1981 (N_1981,N_271,N_177);
and U1982 (N_1982,N_198,N_802);
nor U1983 (N_1983,N_374,N_755);
nand U1984 (N_1984,N_713,N_533);
nor U1985 (N_1985,N_392,N_907);
nor U1986 (N_1986,N_51,N_828);
and U1987 (N_1987,N_561,N_901);
nand U1988 (N_1988,N_220,N_870);
nand U1989 (N_1989,N_817,N_265);
or U1990 (N_1990,N_102,N_97);
nand U1991 (N_1991,N_202,N_525);
and U1992 (N_1992,N_624,N_36);
xor U1993 (N_1993,N_372,N_171);
or U1994 (N_1994,N_117,N_955);
nor U1995 (N_1995,N_40,N_92);
and U1996 (N_1996,N_989,N_324);
or U1997 (N_1997,N_187,N_940);
and U1998 (N_1998,N_976,N_974);
or U1999 (N_1999,N_242,N_497);
nor U2000 (N_2000,N_1726,N_1751);
or U2001 (N_2001,N_1570,N_1446);
nand U2002 (N_2002,N_1492,N_1970);
nor U2003 (N_2003,N_1364,N_1824);
nor U2004 (N_2004,N_1049,N_1300);
and U2005 (N_2005,N_1964,N_1999);
nand U2006 (N_2006,N_1563,N_1417);
nand U2007 (N_2007,N_1222,N_1474);
nand U2008 (N_2008,N_1822,N_1249);
and U2009 (N_2009,N_1915,N_1293);
nand U2010 (N_2010,N_1643,N_1745);
or U2011 (N_2011,N_1242,N_1285);
nor U2012 (N_2012,N_1121,N_1012);
and U2013 (N_2013,N_1157,N_1835);
nand U2014 (N_2014,N_1821,N_1163);
xnor U2015 (N_2015,N_1944,N_1609);
or U2016 (N_2016,N_1206,N_1568);
and U2017 (N_2017,N_1036,N_1830);
and U2018 (N_2018,N_1599,N_1968);
nand U2019 (N_2019,N_1502,N_1829);
or U2020 (N_2020,N_1008,N_1045);
and U2021 (N_2021,N_1062,N_1001);
and U2022 (N_2022,N_1865,N_1733);
nor U2023 (N_2023,N_1578,N_1017);
or U2024 (N_2024,N_1527,N_1781);
nand U2025 (N_2025,N_1436,N_1391);
and U2026 (N_2026,N_1434,N_1201);
and U2027 (N_2027,N_1357,N_1681);
and U2028 (N_2028,N_1621,N_1481);
nand U2029 (N_2029,N_1234,N_1287);
nand U2030 (N_2030,N_1272,N_1267);
or U2031 (N_2031,N_1322,N_1808);
and U2032 (N_2032,N_1345,N_1675);
and U2033 (N_2033,N_1542,N_1101);
nand U2034 (N_2034,N_1102,N_1535);
and U2035 (N_2035,N_1512,N_1583);
and U2036 (N_2036,N_1940,N_1370);
or U2037 (N_2037,N_1847,N_1320);
nor U2038 (N_2038,N_1288,N_1277);
nor U2039 (N_2039,N_1591,N_1715);
xnor U2040 (N_2040,N_1831,N_1221);
or U2041 (N_2041,N_1392,N_1368);
nor U2042 (N_2042,N_1039,N_1683);
nor U2043 (N_2043,N_1034,N_1554);
or U2044 (N_2044,N_1615,N_1185);
and U2045 (N_2045,N_1735,N_1150);
nand U2046 (N_2046,N_1212,N_1190);
or U2047 (N_2047,N_1099,N_1213);
nand U2048 (N_2048,N_1027,N_1893);
or U2049 (N_2049,N_1953,N_1306);
nor U2050 (N_2050,N_1038,N_1962);
xor U2051 (N_2051,N_1172,N_1812);
nor U2052 (N_2052,N_1601,N_1861);
or U2053 (N_2053,N_1878,N_1916);
nand U2054 (N_2054,N_1333,N_1700);
nand U2055 (N_2055,N_1404,N_1985);
nor U2056 (N_2056,N_1389,N_1562);
xor U2057 (N_2057,N_1005,N_1476);
nor U2058 (N_2058,N_1956,N_1314);
xnor U2059 (N_2059,N_1097,N_1973);
and U2060 (N_2060,N_1498,N_1536);
xor U2061 (N_2061,N_1044,N_1667);
nand U2062 (N_2062,N_1807,N_1084);
xnor U2063 (N_2063,N_1367,N_1676);
nor U2064 (N_2064,N_1655,N_1886);
nor U2065 (N_2065,N_1432,N_1445);
or U2066 (N_2066,N_1025,N_1278);
nand U2067 (N_2067,N_1620,N_1647);
or U2068 (N_2068,N_1522,N_1879);
and U2069 (N_2069,N_1447,N_1261);
and U2070 (N_2070,N_1604,N_1187);
nor U2071 (N_2071,N_1672,N_1792);
and U2072 (N_2072,N_1454,N_1144);
and U2073 (N_2073,N_1086,N_1900);
and U2074 (N_2074,N_1855,N_1938);
and U2075 (N_2075,N_1632,N_1466);
nor U2076 (N_2076,N_1580,N_1074);
or U2077 (N_2077,N_1301,N_1550);
xor U2078 (N_2078,N_1603,N_1828);
nand U2079 (N_2079,N_1087,N_1024);
nor U2080 (N_2080,N_1903,N_1375);
xnor U2081 (N_2081,N_1585,N_1203);
or U2082 (N_2082,N_1959,N_1505);
nand U2083 (N_2083,N_1553,N_1456);
nand U2084 (N_2084,N_1720,N_1266);
xnor U2085 (N_2085,N_1529,N_1537);
nand U2086 (N_2086,N_1011,N_1707);
or U2087 (N_2087,N_1761,N_1794);
and U2088 (N_2088,N_1588,N_1227);
xnor U2089 (N_2089,N_1495,N_1079);
nand U2090 (N_2090,N_1414,N_1351);
nor U2091 (N_2091,N_1166,N_1022);
nand U2092 (N_2092,N_1584,N_1216);
nor U2093 (N_2093,N_1067,N_1625);
or U2094 (N_2094,N_1590,N_1437);
and U2095 (N_2095,N_1941,N_1549);
or U2096 (N_2096,N_1159,N_1983);
nor U2097 (N_2097,N_1654,N_1613);
nand U2098 (N_2098,N_1050,N_1698);
nand U2099 (N_2099,N_1308,N_1862);
or U2100 (N_2100,N_1165,N_1282);
or U2101 (N_2101,N_1708,N_1352);
or U2102 (N_2102,N_1449,N_1104);
or U2103 (N_2103,N_1534,N_1988);
or U2104 (N_2104,N_1366,N_1825);
nor U2105 (N_2105,N_1302,N_1774);
nand U2106 (N_2106,N_1094,N_1678);
xnor U2107 (N_2107,N_1523,N_1219);
or U2108 (N_2108,N_1612,N_1026);
nor U2109 (N_2109,N_1056,N_1530);
and U2110 (N_2110,N_1813,N_1650);
or U2111 (N_2111,N_1853,N_1054);
or U2112 (N_2112,N_1021,N_1003);
nor U2113 (N_2113,N_1051,N_1348);
or U2114 (N_2114,N_1371,N_1421);
nand U2115 (N_2115,N_1838,N_1564);
or U2116 (N_2116,N_1799,N_1856);
nor U2117 (N_2117,N_1491,N_1233);
and U2118 (N_2118,N_1737,N_1410);
or U2119 (N_2119,N_1326,N_1633);
nand U2120 (N_2120,N_1706,N_1118);
and U2121 (N_2121,N_1451,N_1089);
and U2122 (N_2122,N_1137,N_1639);
or U2123 (N_2123,N_1228,N_1197);
and U2124 (N_2124,N_1384,N_1096);
and U2125 (N_2125,N_1532,N_1070);
nor U2126 (N_2126,N_1264,N_1624);
nand U2127 (N_2127,N_1939,N_1839);
xor U2128 (N_2128,N_1385,N_1194);
or U2129 (N_2129,N_1377,N_1161);
and U2130 (N_2130,N_1395,N_1778);
nor U2131 (N_2131,N_1468,N_1969);
xnor U2132 (N_2132,N_1577,N_1690);
nor U2133 (N_2133,N_1411,N_1037);
nand U2134 (N_2134,N_1184,N_1902);
nor U2135 (N_2135,N_1611,N_1763);
nor U2136 (N_2136,N_1283,N_1866);
xnor U2137 (N_2137,N_1006,N_1112);
or U2138 (N_2138,N_1975,N_1355);
or U2139 (N_2139,N_1732,N_1400);
or U2140 (N_2140,N_1494,N_1134);
and U2141 (N_2141,N_1873,N_1842);
or U2142 (N_2142,N_1606,N_1775);
or U2143 (N_2143,N_1519,N_1111);
xnor U2144 (N_2144,N_1235,N_1817);
or U2145 (N_2145,N_1214,N_1365);
or U2146 (N_2146,N_1889,N_1891);
nor U2147 (N_2147,N_1296,N_1605);
nand U2148 (N_2148,N_1061,N_1338);
or U2149 (N_2149,N_1191,N_1107);
xnor U2150 (N_2150,N_1046,N_1120);
nand U2151 (N_2151,N_1617,N_1630);
and U2152 (N_2152,N_1488,N_1115);
or U2153 (N_2153,N_1731,N_1147);
and U2154 (N_2154,N_1057,N_1415);
nand U2155 (N_2155,N_1782,N_1608);
nor U2156 (N_2156,N_1279,N_1823);
and U2157 (N_2157,N_1618,N_1472);
nand U2158 (N_2158,N_1518,N_1709);
nor U2159 (N_2159,N_1321,N_1933);
nand U2160 (N_2160,N_1907,N_1133);
nand U2161 (N_2161,N_1635,N_1232);
nor U2162 (N_2162,N_1188,N_1131);
nor U2163 (N_2163,N_1425,N_1149);
nor U2164 (N_2164,N_1546,N_1381);
nor U2165 (N_2165,N_1260,N_1575);
and U2166 (N_2166,N_1085,N_1090);
nand U2167 (N_2167,N_1356,N_1660);
nor U2168 (N_2168,N_1652,N_1153);
nand U2169 (N_2169,N_1487,N_1480);
nand U2170 (N_2170,N_1042,N_1141);
xor U2171 (N_2171,N_1286,N_1353);
nand U2172 (N_2172,N_1990,N_1937);
nor U2173 (N_2173,N_1503,N_1091);
or U2174 (N_2174,N_1884,N_1475);
nand U2175 (N_2175,N_1610,N_1092);
nand U2176 (N_2176,N_1435,N_1229);
nand U2177 (N_2177,N_1173,N_1904);
or U2178 (N_2178,N_1028,N_1573);
and U2179 (N_2179,N_1734,N_1772);
or U2180 (N_2180,N_1559,N_1909);
nand U2181 (N_2181,N_1183,N_1545);
nand U2182 (N_2182,N_1509,N_1656);
nor U2183 (N_2183,N_1696,N_1803);
and U2184 (N_2184,N_1402,N_1066);
xor U2185 (N_2185,N_1463,N_1294);
nand U2186 (N_2186,N_1342,N_1752);
xnor U2187 (N_2187,N_1925,N_1511);
nor U2188 (N_2188,N_1258,N_1832);
or U2189 (N_2189,N_1030,N_1015);
nand U2190 (N_2190,N_1507,N_1297);
and U2191 (N_2191,N_1299,N_1238);
nor U2192 (N_2192,N_1957,N_1344);
and U2193 (N_2193,N_1117,N_1255);
or U2194 (N_2194,N_1789,N_1156);
nand U2195 (N_2195,N_1477,N_1019);
nor U2196 (N_2196,N_1952,N_1547);
nand U2197 (N_2197,N_1848,N_1020);
and U2198 (N_2198,N_1883,N_1629);
and U2199 (N_2199,N_1424,N_1976);
or U2200 (N_2200,N_1557,N_1148);
xor U2201 (N_2201,N_1685,N_1926);
and U2202 (N_2202,N_1478,N_1710);
nand U2203 (N_2203,N_1671,N_1533);
and U2204 (N_2204,N_1440,N_1482);
or U2205 (N_2205,N_1922,N_1651);
nor U2206 (N_2206,N_1524,N_1493);
nand U2207 (N_2207,N_1958,N_1325);
or U2208 (N_2208,N_1467,N_1510);
nor U2209 (N_2209,N_1363,N_1140);
nor U2210 (N_2210,N_1064,N_1243);
nand U2211 (N_2211,N_1899,N_1721);
or U2212 (N_2212,N_1490,N_1935);
nand U2213 (N_2213,N_1628,N_1182);
and U2214 (N_2214,N_1949,N_1598);
nand U2215 (N_2215,N_1428,N_1442);
and U2216 (N_2216,N_1984,N_1174);
nor U2217 (N_2217,N_1426,N_1041);
nor U2218 (N_2218,N_1677,N_1138);
or U2219 (N_2219,N_1589,N_1974);
or U2220 (N_2220,N_1892,N_1747);
nand U2221 (N_2221,N_1016,N_1077);
nor U2222 (N_2222,N_1836,N_1506);
or U2223 (N_2223,N_1465,N_1906);
nor U2224 (N_2224,N_1749,N_1776);
nor U2225 (N_2225,N_1179,N_1080);
nor U2226 (N_2226,N_1035,N_1566);
nand U2227 (N_2227,N_1796,N_1429);
nand U2228 (N_2228,N_1380,N_1082);
and U2229 (N_2229,N_1431,N_1693);
and U2230 (N_2230,N_1418,N_1397);
nand U2231 (N_2231,N_1544,N_1723);
or U2232 (N_2232,N_1311,N_1770);
and U2233 (N_2233,N_1127,N_1768);
and U2234 (N_2234,N_1180,N_1000);
or U2235 (N_2235,N_1398,N_1664);
nor U2236 (N_2236,N_1572,N_1728);
nor U2237 (N_2237,N_1211,N_1586);
or U2238 (N_2238,N_1315,N_1558);
xnor U2239 (N_2239,N_1863,N_1614);
and U2240 (N_2240,N_1644,N_1849);
and U2241 (N_2241,N_1078,N_1059);
and U2242 (N_2242,N_1323,N_1433);
and U2243 (N_2243,N_1200,N_1661);
xor U2244 (N_2244,N_1162,N_1210);
and U2245 (N_2245,N_1245,N_1483);
and U2246 (N_2246,N_1827,N_1053);
and U2247 (N_2247,N_1724,N_1125);
nor U2248 (N_2248,N_1443,N_1539);
nand U2249 (N_2249,N_1921,N_1122);
nand U2250 (N_2250,N_1631,N_1170);
xor U2251 (N_2251,N_1390,N_1779);
or U2252 (N_2252,N_1209,N_1762);
and U2253 (N_2253,N_1936,N_1199);
or U2254 (N_2254,N_1928,N_1945);
or U2255 (N_2255,N_1666,N_1874);
and U2256 (N_2256,N_1627,N_1977);
or U2257 (N_2257,N_1877,N_1388);
nand U2258 (N_2258,N_1815,N_1753);
or U2259 (N_2259,N_1638,N_1119);
nor U2260 (N_2260,N_1335,N_1453);
nor U2261 (N_2261,N_1459,N_1237);
and U2262 (N_2262,N_1581,N_1961);
nor U2263 (N_2263,N_1670,N_1126);
nor U2264 (N_2264,N_1576,N_1504);
xor U2265 (N_2265,N_1354,N_1450);
and U2266 (N_2266,N_1387,N_1919);
nand U2267 (N_2267,N_1766,N_1247);
or U2268 (N_2268,N_1596,N_1382);
nand U2269 (N_2269,N_1095,N_1595);
nor U2270 (N_2270,N_1181,N_1955);
and U2271 (N_2271,N_1309,N_1997);
xnor U2272 (N_2272,N_1489,N_1154);
or U2273 (N_2273,N_1637,N_1273);
nand U2274 (N_2274,N_1204,N_1018);
and U2275 (N_2275,N_1526,N_1754);
nor U2276 (N_2276,N_1236,N_1259);
or U2277 (N_2277,N_1420,N_1727);
and U2278 (N_2278,N_1816,N_1826);
and U2279 (N_2279,N_1202,N_1324);
or U2280 (N_2280,N_1850,N_1641);
or U2281 (N_2281,N_1508,N_1729);
or U2282 (N_2282,N_1640,N_1911);
and U2283 (N_2283,N_1248,N_1275);
nor U2284 (N_2284,N_1994,N_1905);
xor U2285 (N_2285,N_1464,N_1818);
nor U2286 (N_2286,N_1555,N_1561);
nor U2287 (N_2287,N_1602,N_1291);
or U2288 (N_2288,N_1452,N_1784);
nand U2289 (N_2289,N_1594,N_1177);
nand U2290 (N_2290,N_1801,N_1719);
or U2291 (N_2291,N_1755,N_1864);
nor U2292 (N_2292,N_1810,N_1393);
or U2293 (N_2293,N_1995,N_1551);
xor U2294 (N_2294,N_1350,N_1256);
nand U2295 (N_2295,N_1205,N_1341);
nand U2296 (N_2296,N_1725,N_1673);
nor U2297 (N_2297,N_1569,N_1110);
or U2298 (N_2298,N_1337,N_1951);
xor U2299 (N_2299,N_1556,N_1742);
nand U2300 (N_2300,N_1088,N_1800);
nor U2301 (N_2301,N_1113,N_1739);
nand U2302 (N_2302,N_1979,N_1010);
nor U2303 (N_2303,N_1416,N_1422);
nand U2304 (N_2304,N_1132,N_1047);
xor U2305 (N_2305,N_1890,N_1600);
nor U2306 (N_2306,N_1339,N_1298);
xnor U2307 (N_2307,N_1695,N_1499);
nand U2308 (N_2308,N_1697,N_1448);
and U2309 (N_2309,N_1854,N_1330);
and U2310 (N_2310,N_1517,N_1901);
or U2311 (N_2311,N_1623,N_1531);
and U2312 (N_2312,N_1691,N_1744);
and U2313 (N_2313,N_1767,N_1152);
nor U2314 (N_2314,N_1845,N_1423);
or U2315 (N_2315,N_1250,N_1662);
or U2316 (N_2316,N_1646,N_1819);
or U2317 (N_2317,N_1269,N_1978);
nand U2318 (N_2318,N_1262,N_1934);
or U2319 (N_2319,N_1791,N_1307);
or U2320 (N_2320,N_1765,N_1332);
or U2321 (N_2321,N_1738,N_1318);
and U2322 (N_2322,N_1931,N_1178);
nand U2323 (N_2323,N_1193,N_1023);
nor U2324 (N_2324,N_1303,N_1083);
nand U2325 (N_2325,N_1783,N_1328);
and U2326 (N_2326,N_1396,N_1100);
or U2327 (N_2327,N_1841,N_1859);
and U2328 (N_2328,N_1648,N_1574);
nor U2329 (N_2329,N_1963,N_1760);
or U2330 (N_2330,N_1276,N_1642);
and U2331 (N_2331,N_1349,N_1362);
or U2332 (N_2332,N_1746,N_1567);
nor U2333 (N_2333,N_1918,N_1653);
nand U2334 (N_2334,N_1058,N_1109);
nand U2335 (N_2335,N_1773,N_1699);
nor U2336 (N_2336,N_1674,N_1972);
nand U2337 (N_2337,N_1541,N_1868);
nor U2338 (N_2338,N_1917,N_1319);
nand U2339 (N_2339,N_1930,N_1469);
and U2340 (N_2340,N_1966,N_1920);
nor U2341 (N_2341,N_1254,N_1947);
nor U2342 (N_2342,N_1441,N_1871);
nor U2343 (N_2343,N_1718,N_1063);
nand U2344 (N_2344,N_1274,N_1663);
nand U2345 (N_2345,N_1497,N_1155);
nand U2346 (N_2346,N_1960,N_1002);
or U2347 (N_2347,N_1657,N_1270);
and U2348 (N_2348,N_1457,N_1128);
nand U2349 (N_2349,N_1607,N_1484);
nor U2350 (N_2350,N_1649,N_1797);
nor U2351 (N_2351,N_1694,N_1548);
nor U2352 (N_2352,N_1251,N_1785);
and U2353 (N_2353,N_1769,N_1597);
and U2354 (N_2354,N_1386,N_1013);
or U2355 (N_2355,N_1130,N_1914);
or U2356 (N_2356,N_1712,N_1171);
and U2357 (N_2357,N_1971,N_1679);
nor U2358 (N_2358,N_1814,N_1908);
and U2359 (N_2359,N_1076,N_1593);
and U2360 (N_2360,N_1032,N_1327);
nand U2361 (N_2361,N_1924,N_1081);
nor U2362 (N_2362,N_1129,N_1403);
or U2363 (N_2363,N_1515,N_1912);
nor U2364 (N_2364,N_1406,N_1145);
nor U2365 (N_2365,N_1896,N_1317);
and U2366 (N_2366,N_1462,N_1427);
and U2367 (N_2367,N_1834,N_1516);
xor U2368 (N_2368,N_1031,N_1965);
nand U2369 (N_2369,N_1992,N_1383);
and U2370 (N_2370,N_1682,N_1833);
nor U2371 (N_2371,N_1169,N_1659);
or U2372 (N_2372,N_1852,N_1790);
nor U2373 (N_2373,N_1098,N_1486);
or U2374 (N_2374,N_1993,N_1991);
or U2375 (N_2375,N_1175,N_1713);
or U2376 (N_2376,N_1135,N_1316);
xor U2377 (N_2377,N_1980,N_1336);
xor U2378 (N_2378,N_1281,N_1804);
or U2379 (N_2379,N_1347,N_1029);
xor U2380 (N_2380,N_1579,N_1343);
xor U2381 (N_2381,N_1750,N_1413);
and U2382 (N_2382,N_1870,N_1186);
or U2383 (N_2383,N_1705,N_1052);
and U2384 (N_2384,N_1802,N_1704);
and U2385 (N_2385,N_1701,N_1379);
and U2386 (N_2386,N_1927,N_1571);
and U2387 (N_2387,N_1060,N_1711);
nor U2388 (N_2388,N_1195,N_1263);
nand U2389 (N_2389,N_1882,N_1473);
xor U2390 (N_2390,N_1369,N_1894);
xor U2391 (N_2391,N_1479,N_1124);
nor U2392 (N_2392,N_1872,N_1736);
and U2393 (N_2393,N_1312,N_1888);
or U2394 (N_2394,N_1207,N_1334);
nor U2395 (N_2395,N_1844,N_1795);
nor U2396 (N_2396,N_1461,N_1717);
nor U2397 (N_2397,N_1998,N_1858);
nand U2398 (N_2398,N_1780,N_1224);
nand U2399 (N_2399,N_1239,N_1876);
nor U2400 (N_2400,N_1756,N_1636);
and U2401 (N_2401,N_1684,N_1967);
or U2402 (N_2402,N_1048,N_1881);
nor U2403 (N_2403,N_1217,N_1072);
and U2404 (N_2404,N_1552,N_1714);
nand U2405 (N_2405,N_1996,N_1645);
nor U2406 (N_2406,N_1412,N_1942);
or U2407 (N_2407,N_1716,N_1009);
or U2408 (N_2408,N_1284,N_1764);
nor U2409 (N_2409,N_1361,N_1004);
and U2410 (N_2410,N_1840,N_1843);
xnor U2411 (N_2411,N_1358,N_1798);
nand U2412 (N_2412,N_1869,N_1225);
nor U2413 (N_2413,N_1168,N_1669);
nor U2414 (N_2414,N_1688,N_1218);
nand U2415 (N_2415,N_1405,N_1265);
xor U2416 (N_2416,N_1913,N_1068);
nand U2417 (N_2417,N_1582,N_1455);
and U2418 (N_2418,N_1528,N_1268);
or U2419 (N_2419,N_1658,N_1360);
nor U2420 (N_2420,N_1758,N_1820);
and U2421 (N_2421,N_1065,N_1932);
nor U2422 (N_2422,N_1143,N_1394);
nand U2423 (N_2423,N_1313,N_1167);
and U2424 (N_2424,N_1787,N_1208);
nand U2425 (N_2425,N_1292,N_1857);
and U2426 (N_2426,N_1895,N_1252);
xor U2427 (N_2427,N_1176,N_1231);
xnor U2428 (N_2428,N_1687,N_1771);
and U2429 (N_2429,N_1875,N_1565);
and U2430 (N_2430,N_1189,N_1142);
nor U2431 (N_2431,N_1592,N_1409);
or U2432 (N_2432,N_1289,N_1280);
nor U2433 (N_2433,N_1069,N_1376);
nor U2434 (N_2434,N_1340,N_1192);
nand U2435 (N_2435,N_1634,N_1106);
xor U2436 (N_2436,N_1033,N_1525);
and U2437 (N_2437,N_1740,N_1867);
nand U2438 (N_2438,N_1226,N_1923);
nor U2439 (N_2439,N_1788,N_1310);
or U2440 (N_2440,N_1806,N_1253);
nor U2441 (N_2441,N_1943,N_1543);
nand U2442 (N_2442,N_1444,N_1014);
or U2443 (N_2443,N_1910,N_1230);
or U2444 (N_2444,N_1500,N_1271);
nand U2445 (N_2445,N_1103,N_1329);
nand U2446 (N_2446,N_1793,N_1692);
nand U2447 (N_2447,N_1501,N_1407);
or U2448 (N_2448,N_1485,N_1240);
nor U2449 (N_2449,N_1374,N_1946);
nand U2450 (N_2450,N_1898,N_1075);
or U2451 (N_2451,N_1430,N_1860);
nand U2452 (N_2452,N_1439,N_1160);
or U2453 (N_2453,N_1887,N_1587);
or U2454 (N_2454,N_1880,N_1851);
nand U2455 (N_2455,N_1616,N_1471);
or U2456 (N_2456,N_1989,N_1460);
nor U2457 (N_2457,N_1811,N_1702);
nand U2458 (N_2458,N_1123,N_1139);
nor U2459 (N_2459,N_1986,N_1540);
nor U2460 (N_2460,N_1007,N_1680);
nand U2461 (N_2461,N_1304,N_1223);
nor U2462 (N_2462,N_1105,N_1560);
or U2463 (N_2463,N_1241,N_1722);
nand U2464 (N_2464,N_1055,N_1257);
nand U2465 (N_2465,N_1689,N_1196);
and U2466 (N_2466,N_1215,N_1626);
nand U2467 (N_2467,N_1748,N_1198);
and U2468 (N_2468,N_1786,N_1136);
or U2469 (N_2469,N_1146,N_1981);
or U2470 (N_2470,N_1846,N_1521);
nor U2471 (N_2471,N_1114,N_1743);
and U2472 (N_2472,N_1346,N_1513);
nand U2473 (N_2473,N_1244,N_1458);
or U2474 (N_2474,N_1837,N_1885);
or U2475 (N_2475,N_1246,N_1419);
and U2476 (N_2476,N_1151,N_1220);
nand U2477 (N_2477,N_1897,N_1950);
or U2478 (N_2478,N_1158,N_1757);
nand U2479 (N_2479,N_1686,N_1703);
nor U2480 (N_2480,N_1496,N_1378);
nor U2481 (N_2481,N_1359,N_1665);
nand U2482 (N_2482,N_1401,N_1777);
nor U2483 (N_2483,N_1073,N_1305);
nand U2484 (N_2484,N_1948,N_1093);
nor U2485 (N_2485,N_1619,N_1438);
xnor U2486 (N_2486,N_1805,N_1987);
and U2487 (N_2487,N_1373,N_1372);
or U2488 (N_2488,N_1043,N_1116);
nand U2489 (N_2489,N_1295,N_1954);
or U2490 (N_2490,N_1290,N_1759);
nand U2491 (N_2491,N_1071,N_1040);
nor U2492 (N_2492,N_1399,N_1809);
xor U2493 (N_2493,N_1164,N_1331);
nor U2494 (N_2494,N_1408,N_1982);
nor U2495 (N_2495,N_1622,N_1470);
xor U2496 (N_2496,N_1520,N_1538);
xor U2497 (N_2497,N_1108,N_1741);
and U2498 (N_2498,N_1730,N_1929);
nand U2499 (N_2499,N_1514,N_1668);
and U2500 (N_2500,N_1591,N_1194);
nor U2501 (N_2501,N_1280,N_1585);
or U2502 (N_2502,N_1909,N_1346);
and U2503 (N_2503,N_1112,N_1517);
xor U2504 (N_2504,N_1912,N_1531);
and U2505 (N_2505,N_1108,N_1425);
or U2506 (N_2506,N_1199,N_1060);
nor U2507 (N_2507,N_1164,N_1320);
or U2508 (N_2508,N_1122,N_1272);
and U2509 (N_2509,N_1411,N_1659);
and U2510 (N_2510,N_1178,N_1008);
nand U2511 (N_2511,N_1027,N_1094);
or U2512 (N_2512,N_1476,N_1913);
nor U2513 (N_2513,N_1610,N_1634);
or U2514 (N_2514,N_1271,N_1486);
or U2515 (N_2515,N_1139,N_1161);
or U2516 (N_2516,N_1532,N_1976);
nand U2517 (N_2517,N_1282,N_1791);
and U2518 (N_2518,N_1097,N_1413);
nor U2519 (N_2519,N_1459,N_1434);
and U2520 (N_2520,N_1127,N_1572);
nor U2521 (N_2521,N_1867,N_1154);
or U2522 (N_2522,N_1089,N_1943);
xor U2523 (N_2523,N_1821,N_1933);
nand U2524 (N_2524,N_1188,N_1013);
or U2525 (N_2525,N_1067,N_1201);
nor U2526 (N_2526,N_1044,N_1712);
nand U2527 (N_2527,N_1392,N_1493);
nor U2528 (N_2528,N_1922,N_1917);
or U2529 (N_2529,N_1822,N_1166);
or U2530 (N_2530,N_1808,N_1934);
nor U2531 (N_2531,N_1395,N_1835);
xor U2532 (N_2532,N_1350,N_1473);
nor U2533 (N_2533,N_1755,N_1924);
and U2534 (N_2534,N_1712,N_1012);
or U2535 (N_2535,N_1459,N_1392);
xor U2536 (N_2536,N_1217,N_1629);
nand U2537 (N_2537,N_1432,N_1459);
nand U2538 (N_2538,N_1624,N_1458);
nor U2539 (N_2539,N_1945,N_1380);
and U2540 (N_2540,N_1846,N_1464);
or U2541 (N_2541,N_1238,N_1187);
or U2542 (N_2542,N_1452,N_1460);
or U2543 (N_2543,N_1904,N_1337);
nor U2544 (N_2544,N_1981,N_1950);
or U2545 (N_2545,N_1044,N_1901);
nand U2546 (N_2546,N_1686,N_1393);
nand U2547 (N_2547,N_1651,N_1539);
or U2548 (N_2548,N_1199,N_1387);
nand U2549 (N_2549,N_1982,N_1858);
nor U2550 (N_2550,N_1481,N_1040);
and U2551 (N_2551,N_1228,N_1329);
or U2552 (N_2552,N_1623,N_1809);
or U2553 (N_2553,N_1335,N_1677);
and U2554 (N_2554,N_1014,N_1309);
nand U2555 (N_2555,N_1319,N_1336);
nand U2556 (N_2556,N_1077,N_1944);
or U2557 (N_2557,N_1655,N_1016);
or U2558 (N_2558,N_1747,N_1656);
and U2559 (N_2559,N_1273,N_1878);
nor U2560 (N_2560,N_1338,N_1330);
nor U2561 (N_2561,N_1750,N_1244);
nand U2562 (N_2562,N_1248,N_1930);
nand U2563 (N_2563,N_1242,N_1088);
nand U2564 (N_2564,N_1309,N_1960);
and U2565 (N_2565,N_1938,N_1522);
or U2566 (N_2566,N_1397,N_1394);
nor U2567 (N_2567,N_1236,N_1245);
nor U2568 (N_2568,N_1917,N_1581);
or U2569 (N_2569,N_1903,N_1449);
and U2570 (N_2570,N_1858,N_1802);
and U2571 (N_2571,N_1676,N_1582);
and U2572 (N_2572,N_1355,N_1661);
and U2573 (N_2573,N_1472,N_1065);
xnor U2574 (N_2574,N_1273,N_1613);
and U2575 (N_2575,N_1355,N_1923);
nor U2576 (N_2576,N_1382,N_1591);
nand U2577 (N_2577,N_1695,N_1379);
or U2578 (N_2578,N_1659,N_1962);
or U2579 (N_2579,N_1177,N_1428);
or U2580 (N_2580,N_1797,N_1890);
nand U2581 (N_2581,N_1004,N_1374);
and U2582 (N_2582,N_1773,N_1129);
nand U2583 (N_2583,N_1526,N_1759);
nand U2584 (N_2584,N_1608,N_1248);
and U2585 (N_2585,N_1355,N_1166);
and U2586 (N_2586,N_1980,N_1076);
or U2587 (N_2587,N_1661,N_1016);
or U2588 (N_2588,N_1785,N_1499);
nand U2589 (N_2589,N_1481,N_1352);
or U2590 (N_2590,N_1787,N_1011);
or U2591 (N_2591,N_1156,N_1073);
and U2592 (N_2592,N_1104,N_1695);
or U2593 (N_2593,N_1161,N_1678);
nor U2594 (N_2594,N_1989,N_1352);
or U2595 (N_2595,N_1137,N_1812);
or U2596 (N_2596,N_1184,N_1948);
and U2597 (N_2597,N_1196,N_1416);
nor U2598 (N_2598,N_1282,N_1158);
or U2599 (N_2599,N_1372,N_1344);
and U2600 (N_2600,N_1222,N_1205);
nor U2601 (N_2601,N_1359,N_1097);
or U2602 (N_2602,N_1215,N_1039);
nor U2603 (N_2603,N_1693,N_1320);
xor U2604 (N_2604,N_1774,N_1527);
or U2605 (N_2605,N_1615,N_1370);
and U2606 (N_2606,N_1049,N_1424);
nand U2607 (N_2607,N_1443,N_1896);
or U2608 (N_2608,N_1337,N_1667);
or U2609 (N_2609,N_1939,N_1646);
nor U2610 (N_2610,N_1456,N_1463);
or U2611 (N_2611,N_1541,N_1342);
or U2612 (N_2612,N_1854,N_1649);
and U2613 (N_2613,N_1935,N_1325);
or U2614 (N_2614,N_1579,N_1847);
and U2615 (N_2615,N_1205,N_1054);
xnor U2616 (N_2616,N_1384,N_1463);
nor U2617 (N_2617,N_1154,N_1610);
and U2618 (N_2618,N_1694,N_1153);
and U2619 (N_2619,N_1541,N_1272);
and U2620 (N_2620,N_1385,N_1269);
nor U2621 (N_2621,N_1941,N_1552);
nand U2622 (N_2622,N_1455,N_1076);
nor U2623 (N_2623,N_1643,N_1068);
xnor U2624 (N_2624,N_1890,N_1535);
nor U2625 (N_2625,N_1630,N_1169);
and U2626 (N_2626,N_1719,N_1643);
nand U2627 (N_2627,N_1313,N_1562);
nor U2628 (N_2628,N_1312,N_1320);
or U2629 (N_2629,N_1121,N_1031);
and U2630 (N_2630,N_1868,N_1632);
and U2631 (N_2631,N_1843,N_1895);
xor U2632 (N_2632,N_1990,N_1169);
nor U2633 (N_2633,N_1122,N_1400);
nor U2634 (N_2634,N_1714,N_1750);
and U2635 (N_2635,N_1947,N_1966);
nor U2636 (N_2636,N_1030,N_1035);
or U2637 (N_2637,N_1269,N_1702);
nor U2638 (N_2638,N_1415,N_1700);
xor U2639 (N_2639,N_1210,N_1091);
nand U2640 (N_2640,N_1648,N_1011);
and U2641 (N_2641,N_1886,N_1002);
nand U2642 (N_2642,N_1962,N_1016);
and U2643 (N_2643,N_1851,N_1953);
xor U2644 (N_2644,N_1038,N_1512);
nor U2645 (N_2645,N_1541,N_1652);
nand U2646 (N_2646,N_1648,N_1088);
nand U2647 (N_2647,N_1478,N_1882);
xnor U2648 (N_2648,N_1157,N_1604);
and U2649 (N_2649,N_1260,N_1057);
or U2650 (N_2650,N_1863,N_1852);
xor U2651 (N_2651,N_1072,N_1909);
nor U2652 (N_2652,N_1890,N_1651);
xor U2653 (N_2653,N_1680,N_1967);
xor U2654 (N_2654,N_1081,N_1069);
nand U2655 (N_2655,N_1698,N_1539);
nand U2656 (N_2656,N_1622,N_1997);
and U2657 (N_2657,N_1255,N_1057);
nor U2658 (N_2658,N_1105,N_1425);
nand U2659 (N_2659,N_1938,N_1793);
and U2660 (N_2660,N_1023,N_1764);
and U2661 (N_2661,N_1318,N_1743);
xnor U2662 (N_2662,N_1247,N_1281);
or U2663 (N_2663,N_1473,N_1459);
nor U2664 (N_2664,N_1381,N_1442);
nor U2665 (N_2665,N_1709,N_1941);
nand U2666 (N_2666,N_1149,N_1875);
nand U2667 (N_2667,N_1060,N_1013);
xnor U2668 (N_2668,N_1725,N_1313);
and U2669 (N_2669,N_1960,N_1367);
nand U2670 (N_2670,N_1678,N_1103);
nor U2671 (N_2671,N_1483,N_1521);
nand U2672 (N_2672,N_1607,N_1645);
or U2673 (N_2673,N_1143,N_1948);
nand U2674 (N_2674,N_1486,N_1162);
nand U2675 (N_2675,N_1771,N_1365);
nand U2676 (N_2676,N_1624,N_1099);
xnor U2677 (N_2677,N_1779,N_1920);
and U2678 (N_2678,N_1978,N_1935);
or U2679 (N_2679,N_1052,N_1802);
and U2680 (N_2680,N_1574,N_1476);
nand U2681 (N_2681,N_1770,N_1366);
nor U2682 (N_2682,N_1100,N_1820);
nand U2683 (N_2683,N_1122,N_1524);
and U2684 (N_2684,N_1032,N_1284);
or U2685 (N_2685,N_1211,N_1420);
or U2686 (N_2686,N_1991,N_1235);
and U2687 (N_2687,N_1672,N_1502);
xnor U2688 (N_2688,N_1363,N_1110);
nor U2689 (N_2689,N_1128,N_1974);
or U2690 (N_2690,N_1870,N_1931);
or U2691 (N_2691,N_1702,N_1283);
and U2692 (N_2692,N_1399,N_1209);
nand U2693 (N_2693,N_1405,N_1129);
nand U2694 (N_2694,N_1194,N_1403);
xor U2695 (N_2695,N_1661,N_1316);
nor U2696 (N_2696,N_1841,N_1513);
nand U2697 (N_2697,N_1054,N_1004);
xnor U2698 (N_2698,N_1142,N_1523);
and U2699 (N_2699,N_1526,N_1238);
and U2700 (N_2700,N_1249,N_1428);
nor U2701 (N_2701,N_1232,N_1672);
and U2702 (N_2702,N_1155,N_1412);
and U2703 (N_2703,N_1914,N_1149);
nand U2704 (N_2704,N_1958,N_1174);
nand U2705 (N_2705,N_1794,N_1295);
and U2706 (N_2706,N_1487,N_1423);
or U2707 (N_2707,N_1894,N_1113);
xnor U2708 (N_2708,N_1133,N_1004);
and U2709 (N_2709,N_1596,N_1114);
or U2710 (N_2710,N_1180,N_1369);
and U2711 (N_2711,N_1996,N_1295);
xor U2712 (N_2712,N_1749,N_1895);
and U2713 (N_2713,N_1215,N_1302);
or U2714 (N_2714,N_1716,N_1603);
or U2715 (N_2715,N_1076,N_1531);
and U2716 (N_2716,N_1417,N_1985);
nand U2717 (N_2717,N_1510,N_1514);
xor U2718 (N_2718,N_1107,N_1398);
nor U2719 (N_2719,N_1715,N_1237);
xnor U2720 (N_2720,N_1260,N_1247);
and U2721 (N_2721,N_1689,N_1536);
nor U2722 (N_2722,N_1261,N_1877);
or U2723 (N_2723,N_1679,N_1282);
nor U2724 (N_2724,N_1996,N_1647);
nand U2725 (N_2725,N_1625,N_1501);
or U2726 (N_2726,N_1381,N_1186);
nand U2727 (N_2727,N_1201,N_1622);
and U2728 (N_2728,N_1753,N_1488);
and U2729 (N_2729,N_1913,N_1089);
or U2730 (N_2730,N_1210,N_1297);
or U2731 (N_2731,N_1123,N_1630);
nand U2732 (N_2732,N_1737,N_1026);
nor U2733 (N_2733,N_1048,N_1095);
and U2734 (N_2734,N_1412,N_1705);
nand U2735 (N_2735,N_1633,N_1077);
nor U2736 (N_2736,N_1556,N_1375);
nor U2737 (N_2737,N_1420,N_1336);
and U2738 (N_2738,N_1085,N_1057);
nor U2739 (N_2739,N_1982,N_1704);
nor U2740 (N_2740,N_1004,N_1776);
nor U2741 (N_2741,N_1230,N_1313);
and U2742 (N_2742,N_1758,N_1783);
nor U2743 (N_2743,N_1158,N_1091);
or U2744 (N_2744,N_1059,N_1032);
nand U2745 (N_2745,N_1235,N_1740);
nor U2746 (N_2746,N_1961,N_1478);
nand U2747 (N_2747,N_1955,N_1302);
nor U2748 (N_2748,N_1599,N_1331);
nand U2749 (N_2749,N_1675,N_1269);
nor U2750 (N_2750,N_1504,N_1422);
xor U2751 (N_2751,N_1137,N_1046);
nand U2752 (N_2752,N_1594,N_1988);
nand U2753 (N_2753,N_1841,N_1401);
nand U2754 (N_2754,N_1893,N_1996);
and U2755 (N_2755,N_1317,N_1295);
or U2756 (N_2756,N_1471,N_1126);
or U2757 (N_2757,N_1490,N_1048);
nor U2758 (N_2758,N_1633,N_1978);
nand U2759 (N_2759,N_1836,N_1359);
or U2760 (N_2760,N_1504,N_1727);
xor U2761 (N_2761,N_1759,N_1719);
nor U2762 (N_2762,N_1043,N_1345);
nand U2763 (N_2763,N_1448,N_1782);
nand U2764 (N_2764,N_1684,N_1394);
nor U2765 (N_2765,N_1198,N_1463);
and U2766 (N_2766,N_1158,N_1728);
and U2767 (N_2767,N_1366,N_1369);
nand U2768 (N_2768,N_1954,N_1316);
and U2769 (N_2769,N_1959,N_1126);
or U2770 (N_2770,N_1681,N_1330);
nor U2771 (N_2771,N_1943,N_1402);
or U2772 (N_2772,N_1519,N_1160);
nor U2773 (N_2773,N_1730,N_1673);
and U2774 (N_2774,N_1510,N_1914);
and U2775 (N_2775,N_1100,N_1765);
xnor U2776 (N_2776,N_1662,N_1850);
or U2777 (N_2777,N_1063,N_1904);
or U2778 (N_2778,N_1568,N_1654);
or U2779 (N_2779,N_1750,N_1525);
or U2780 (N_2780,N_1433,N_1864);
or U2781 (N_2781,N_1500,N_1309);
or U2782 (N_2782,N_1851,N_1164);
and U2783 (N_2783,N_1758,N_1927);
xor U2784 (N_2784,N_1680,N_1735);
nand U2785 (N_2785,N_1520,N_1492);
and U2786 (N_2786,N_1980,N_1471);
or U2787 (N_2787,N_1962,N_1613);
nand U2788 (N_2788,N_1353,N_1974);
and U2789 (N_2789,N_1839,N_1681);
nor U2790 (N_2790,N_1682,N_1611);
nand U2791 (N_2791,N_1723,N_1811);
nand U2792 (N_2792,N_1352,N_1501);
nand U2793 (N_2793,N_1837,N_1413);
and U2794 (N_2794,N_1943,N_1339);
nor U2795 (N_2795,N_1108,N_1897);
or U2796 (N_2796,N_1284,N_1553);
nand U2797 (N_2797,N_1717,N_1601);
nand U2798 (N_2798,N_1148,N_1606);
and U2799 (N_2799,N_1208,N_1894);
nor U2800 (N_2800,N_1423,N_1377);
nor U2801 (N_2801,N_1152,N_1868);
xor U2802 (N_2802,N_1477,N_1877);
or U2803 (N_2803,N_1989,N_1282);
xnor U2804 (N_2804,N_1395,N_1494);
xor U2805 (N_2805,N_1702,N_1542);
or U2806 (N_2806,N_1945,N_1866);
nor U2807 (N_2807,N_1591,N_1286);
and U2808 (N_2808,N_1461,N_1441);
and U2809 (N_2809,N_1565,N_1234);
or U2810 (N_2810,N_1579,N_1694);
and U2811 (N_2811,N_1839,N_1547);
and U2812 (N_2812,N_1084,N_1751);
and U2813 (N_2813,N_1577,N_1861);
or U2814 (N_2814,N_1973,N_1800);
nor U2815 (N_2815,N_1222,N_1365);
nor U2816 (N_2816,N_1925,N_1795);
xor U2817 (N_2817,N_1324,N_1297);
or U2818 (N_2818,N_1761,N_1035);
xor U2819 (N_2819,N_1736,N_1783);
or U2820 (N_2820,N_1647,N_1809);
nor U2821 (N_2821,N_1817,N_1678);
nand U2822 (N_2822,N_1242,N_1868);
nor U2823 (N_2823,N_1666,N_1194);
and U2824 (N_2824,N_1327,N_1439);
nor U2825 (N_2825,N_1894,N_1027);
or U2826 (N_2826,N_1024,N_1632);
nor U2827 (N_2827,N_1752,N_1265);
nor U2828 (N_2828,N_1479,N_1718);
nor U2829 (N_2829,N_1759,N_1065);
and U2830 (N_2830,N_1442,N_1540);
or U2831 (N_2831,N_1646,N_1168);
xor U2832 (N_2832,N_1883,N_1781);
nand U2833 (N_2833,N_1312,N_1550);
nand U2834 (N_2834,N_1516,N_1073);
nor U2835 (N_2835,N_1084,N_1674);
and U2836 (N_2836,N_1853,N_1022);
or U2837 (N_2837,N_1273,N_1425);
or U2838 (N_2838,N_1297,N_1199);
or U2839 (N_2839,N_1600,N_1644);
nor U2840 (N_2840,N_1277,N_1704);
or U2841 (N_2841,N_1112,N_1877);
or U2842 (N_2842,N_1277,N_1877);
or U2843 (N_2843,N_1558,N_1867);
or U2844 (N_2844,N_1730,N_1837);
nand U2845 (N_2845,N_1528,N_1261);
nor U2846 (N_2846,N_1412,N_1465);
and U2847 (N_2847,N_1155,N_1211);
nor U2848 (N_2848,N_1733,N_1163);
nand U2849 (N_2849,N_1257,N_1659);
nor U2850 (N_2850,N_1762,N_1639);
and U2851 (N_2851,N_1147,N_1298);
nor U2852 (N_2852,N_1018,N_1127);
nor U2853 (N_2853,N_1183,N_1476);
xor U2854 (N_2854,N_1290,N_1213);
nand U2855 (N_2855,N_1919,N_1305);
and U2856 (N_2856,N_1040,N_1918);
nand U2857 (N_2857,N_1641,N_1654);
nor U2858 (N_2858,N_1838,N_1589);
xnor U2859 (N_2859,N_1824,N_1466);
or U2860 (N_2860,N_1500,N_1771);
nand U2861 (N_2861,N_1046,N_1703);
and U2862 (N_2862,N_1864,N_1443);
and U2863 (N_2863,N_1885,N_1033);
or U2864 (N_2864,N_1133,N_1337);
and U2865 (N_2865,N_1206,N_1388);
or U2866 (N_2866,N_1360,N_1826);
and U2867 (N_2867,N_1421,N_1249);
and U2868 (N_2868,N_1001,N_1350);
or U2869 (N_2869,N_1573,N_1113);
or U2870 (N_2870,N_1725,N_1708);
nand U2871 (N_2871,N_1191,N_1848);
or U2872 (N_2872,N_1227,N_1005);
and U2873 (N_2873,N_1703,N_1516);
or U2874 (N_2874,N_1780,N_1033);
nand U2875 (N_2875,N_1763,N_1181);
or U2876 (N_2876,N_1776,N_1748);
or U2877 (N_2877,N_1465,N_1138);
or U2878 (N_2878,N_1661,N_1771);
and U2879 (N_2879,N_1429,N_1607);
nor U2880 (N_2880,N_1649,N_1371);
nand U2881 (N_2881,N_1264,N_1577);
or U2882 (N_2882,N_1781,N_1380);
nand U2883 (N_2883,N_1098,N_1741);
and U2884 (N_2884,N_1754,N_1395);
nor U2885 (N_2885,N_1080,N_1343);
or U2886 (N_2886,N_1339,N_1810);
nand U2887 (N_2887,N_1653,N_1634);
nand U2888 (N_2888,N_1094,N_1270);
nor U2889 (N_2889,N_1343,N_1319);
or U2890 (N_2890,N_1234,N_1463);
nand U2891 (N_2891,N_1537,N_1822);
and U2892 (N_2892,N_1596,N_1001);
nand U2893 (N_2893,N_1031,N_1199);
nor U2894 (N_2894,N_1661,N_1574);
nor U2895 (N_2895,N_1231,N_1981);
xor U2896 (N_2896,N_1746,N_1552);
nand U2897 (N_2897,N_1334,N_1123);
and U2898 (N_2898,N_1790,N_1709);
or U2899 (N_2899,N_1274,N_1939);
or U2900 (N_2900,N_1469,N_1452);
nor U2901 (N_2901,N_1889,N_1246);
nand U2902 (N_2902,N_1854,N_1771);
nor U2903 (N_2903,N_1006,N_1455);
or U2904 (N_2904,N_1192,N_1749);
nand U2905 (N_2905,N_1755,N_1575);
nand U2906 (N_2906,N_1740,N_1481);
nand U2907 (N_2907,N_1400,N_1562);
nor U2908 (N_2908,N_1992,N_1921);
xnor U2909 (N_2909,N_1149,N_1535);
or U2910 (N_2910,N_1672,N_1390);
nor U2911 (N_2911,N_1150,N_1583);
xor U2912 (N_2912,N_1503,N_1268);
nor U2913 (N_2913,N_1433,N_1586);
and U2914 (N_2914,N_1730,N_1995);
and U2915 (N_2915,N_1772,N_1241);
nand U2916 (N_2916,N_1923,N_1324);
nand U2917 (N_2917,N_1295,N_1631);
nor U2918 (N_2918,N_1620,N_1014);
and U2919 (N_2919,N_1902,N_1075);
nand U2920 (N_2920,N_1177,N_1203);
nand U2921 (N_2921,N_1926,N_1950);
or U2922 (N_2922,N_1244,N_1090);
and U2923 (N_2923,N_1449,N_1837);
nor U2924 (N_2924,N_1572,N_1934);
nor U2925 (N_2925,N_1745,N_1551);
or U2926 (N_2926,N_1871,N_1845);
nor U2927 (N_2927,N_1508,N_1958);
nor U2928 (N_2928,N_1532,N_1974);
nor U2929 (N_2929,N_1793,N_1988);
and U2930 (N_2930,N_1889,N_1677);
nor U2931 (N_2931,N_1504,N_1645);
xnor U2932 (N_2932,N_1310,N_1085);
nor U2933 (N_2933,N_1681,N_1925);
xnor U2934 (N_2934,N_1006,N_1079);
or U2935 (N_2935,N_1359,N_1857);
nor U2936 (N_2936,N_1212,N_1047);
nor U2937 (N_2937,N_1997,N_1815);
xnor U2938 (N_2938,N_1447,N_1671);
nand U2939 (N_2939,N_1825,N_1624);
nand U2940 (N_2940,N_1563,N_1526);
nor U2941 (N_2941,N_1883,N_1831);
and U2942 (N_2942,N_1828,N_1289);
xnor U2943 (N_2943,N_1827,N_1394);
nand U2944 (N_2944,N_1524,N_1794);
nor U2945 (N_2945,N_1751,N_1777);
or U2946 (N_2946,N_1073,N_1654);
xor U2947 (N_2947,N_1171,N_1150);
and U2948 (N_2948,N_1412,N_1131);
nor U2949 (N_2949,N_1219,N_1888);
or U2950 (N_2950,N_1810,N_1421);
nor U2951 (N_2951,N_1132,N_1021);
nand U2952 (N_2952,N_1196,N_1600);
nand U2953 (N_2953,N_1492,N_1552);
and U2954 (N_2954,N_1886,N_1923);
and U2955 (N_2955,N_1662,N_1328);
nor U2956 (N_2956,N_1588,N_1357);
nor U2957 (N_2957,N_1829,N_1946);
nand U2958 (N_2958,N_1932,N_1905);
nor U2959 (N_2959,N_1403,N_1522);
nand U2960 (N_2960,N_1652,N_1051);
nand U2961 (N_2961,N_1351,N_1564);
nand U2962 (N_2962,N_1974,N_1765);
nand U2963 (N_2963,N_1357,N_1557);
or U2964 (N_2964,N_1311,N_1596);
nor U2965 (N_2965,N_1877,N_1669);
nand U2966 (N_2966,N_1302,N_1227);
or U2967 (N_2967,N_1982,N_1536);
nor U2968 (N_2968,N_1014,N_1636);
nand U2969 (N_2969,N_1227,N_1341);
nand U2970 (N_2970,N_1343,N_1895);
and U2971 (N_2971,N_1276,N_1036);
or U2972 (N_2972,N_1096,N_1416);
nand U2973 (N_2973,N_1217,N_1057);
or U2974 (N_2974,N_1160,N_1143);
nand U2975 (N_2975,N_1099,N_1298);
or U2976 (N_2976,N_1078,N_1614);
nand U2977 (N_2977,N_1571,N_1696);
xor U2978 (N_2978,N_1768,N_1523);
nand U2979 (N_2979,N_1302,N_1171);
or U2980 (N_2980,N_1555,N_1867);
or U2981 (N_2981,N_1918,N_1013);
nand U2982 (N_2982,N_1944,N_1276);
or U2983 (N_2983,N_1908,N_1938);
or U2984 (N_2984,N_1682,N_1410);
nor U2985 (N_2985,N_1566,N_1428);
and U2986 (N_2986,N_1022,N_1046);
nand U2987 (N_2987,N_1539,N_1509);
nor U2988 (N_2988,N_1061,N_1861);
nor U2989 (N_2989,N_1076,N_1211);
nor U2990 (N_2990,N_1144,N_1426);
nand U2991 (N_2991,N_1150,N_1716);
or U2992 (N_2992,N_1101,N_1511);
xnor U2993 (N_2993,N_1836,N_1541);
or U2994 (N_2994,N_1054,N_1789);
nor U2995 (N_2995,N_1858,N_1450);
or U2996 (N_2996,N_1927,N_1754);
nand U2997 (N_2997,N_1375,N_1317);
or U2998 (N_2998,N_1048,N_1793);
and U2999 (N_2999,N_1493,N_1245);
nand U3000 (N_3000,N_2006,N_2372);
nor U3001 (N_3001,N_2499,N_2961);
nor U3002 (N_3002,N_2406,N_2503);
xor U3003 (N_3003,N_2253,N_2160);
or U3004 (N_3004,N_2690,N_2319);
nor U3005 (N_3005,N_2075,N_2935);
xor U3006 (N_3006,N_2665,N_2479);
or U3007 (N_3007,N_2857,N_2305);
nor U3008 (N_3008,N_2177,N_2807);
nand U3009 (N_3009,N_2995,N_2063);
or U3010 (N_3010,N_2072,N_2200);
and U3011 (N_3011,N_2929,N_2512);
and U3012 (N_3012,N_2909,N_2489);
nand U3013 (N_3013,N_2614,N_2097);
nand U3014 (N_3014,N_2147,N_2481);
nor U3015 (N_3015,N_2783,N_2007);
and U3016 (N_3016,N_2603,N_2394);
or U3017 (N_3017,N_2440,N_2657);
nand U3018 (N_3018,N_2326,N_2618);
and U3019 (N_3019,N_2140,N_2718);
and U3020 (N_3020,N_2050,N_2798);
or U3021 (N_3021,N_2809,N_2528);
or U3022 (N_3022,N_2327,N_2679);
xor U3023 (N_3023,N_2056,N_2547);
nand U3024 (N_3024,N_2136,N_2170);
or U3025 (N_3025,N_2633,N_2012);
nand U3026 (N_3026,N_2716,N_2014);
xnor U3027 (N_3027,N_2506,N_2087);
and U3028 (N_3028,N_2281,N_2786);
nand U3029 (N_3029,N_2088,N_2445);
nor U3030 (N_3030,N_2367,N_2708);
nand U3031 (N_3031,N_2846,N_2686);
nor U3032 (N_3032,N_2987,N_2685);
and U3033 (N_3033,N_2859,N_2167);
nor U3034 (N_3034,N_2599,N_2661);
and U3035 (N_3035,N_2758,N_2399);
nand U3036 (N_3036,N_2335,N_2328);
and U3037 (N_3037,N_2789,N_2055);
xor U3038 (N_3038,N_2849,N_2856);
nor U3039 (N_3039,N_2704,N_2689);
nor U3040 (N_3040,N_2184,N_2794);
nor U3041 (N_3041,N_2196,N_2141);
nor U3042 (N_3042,N_2076,N_2299);
nor U3043 (N_3043,N_2166,N_2617);
and U3044 (N_3044,N_2418,N_2414);
nor U3045 (N_3045,N_2611,N_2060);
and U3046 (N_3046,N_2377,N_2483);
nor U3047 (N_3047,N_2575,N_2344);
nand U3048 (N_3048,N_2877,N_2897);
nor U3049 (N_3049,N_2062,N_2355);
or U3050 (N_3050,N_2962,N_2641);
xor U3051 (N_3051,N_2952,N_2924);
and U3052 (N_3052,N_2415,N_2890);
or U3053 (N_3053,N_2564,N_2040);
and U3054 (N_3054,N_2997,N_2828);
or U3055 (N_3055,N_2571,N_2941);
nand U3056 (N_3056,N_2537,N_2265);
and U3057 (N_3057,N_2153,N_2780);
or U3058 (N_3058,N_2687,N_2683);
or U3059 (N_3059,N_2968,N_2039);
nor U3060 (N_3060,N_2357,N_2519);
and U3061 (N_3061,N_2886,N_2317);
nor U3062 (N_3062,N_2126,N_2517);
or U3063 (N_3063,N_2465,N_2002);
nand U3064 (N_3064,N_2252,N_2260);
nor U3065 (N_3065,N_2323,N_2871);
nor U3066 (N_3066,N_2225,N_2868);
xnor U3067 (N_3067,N_2521,N_2923);
and U3068 (N_3068,N_2610,N_2982);
or U3069 (N_3069,N_2092,N_2037);
and U3070 (N_3070,N_2156,N_2241);
or U3071 (N_3071,N_2436,N_2590);
xnor U3072 (N_3072,N_2284,N_2349);
nand U3073 (N_3073,N_2159,N_2747);
nand U3074 (N_3074,N_2172,N_2237);
or U3075 (N_3075,N_2484,N_2870);
nand U3076 (N_3076,N_2762,N_2467);
xor U3077 (N_3077,N_2879,N_2812);
nand U3078 (N_3078,N_2231,N_2423);
nand U3079 (N_3079,N_2824,N_2373);
or U3080 (N_3080,N_2573,N_2726);
or U3081 (N_3081,N_2815,N_2619);
nand U3082 (N_3082,N_2792,N_2214);
nor U3083 (N_3083,N_2767,N_2644);
or U3084 (N_3084,N_2822,N_2179);
and U3085 (N_3085,N_2965,N_2194);
nor U3086 (N_3086,N_2622,N_2643);
xnor U3087 (N_3087,N_2400,N_2369);
xor U3088 (N_3088,N_2460,N_2648);
or U3089 (N_3089,N_2883,N_2667);
nor U3090 (N_3090,N_2473,N_2916);
nand U3091 (N_3091,N_2266,N_2866);
xnor U3092 (N_3092,N_2201,N_2301);
nor U3093 (N_3093,N_2496,N_2675);
nor U3094 (N_3094,N_2936,N_2303);
nor U3095 (N_3095,N_2784,N_2024);
nand U3096 (N_3096,N_2522,N_2663);
or U3097 (N_3097,N_2535,N_2278);
nand U3098 (N_3098,N_2884,N_2861);
and U3099 (N_3099,N_2294,N_2624);
xor U3100 (N_3100,N_2351,N_2984);
nor U3101 (N_3101,N_2920,N_2138);
nand U3102 (N_3102,N_2598,N_2613);
and U3103 (N_3103,N_2739,N_2931);
nor U3104 (N_3104,N_2977,N_2645);
and U3105 (N_3105,N_2205,N_2137);
or U3106 (N_3106,N_2454,N_2158);
xor U3107 (N_3107,N_2606,N_2958);
nor U3108 (N_3108,N_2382,N_2600);
nor U3109 (N_3109,N_2232,N_2998);
or U3110 (N_3110,N_2673,N_2559);
or U3111 (N_3111,N_2550,N_2081);
or U3112 (N_3112,N_2152,N_2124);
or U3113 (N_3113,N_2276,N_2251);
and U3114 (N_3114,N_2270,N_2042);
and U3115 (N_3115,N_2878,N_2086);
nand U3116 (N_3116,N_2412,N_2873);
nand U3117 (N_3117,N_2154,N_2735);
nand U3118 (N_3118,N_2381,N_2209);
nor U3119 (N_3119,N_2130,N_2476);
nor U3120 (N_3120,N_2485,N_2765);
or U3121 (N_3121,N_2132,N_2829);
and U3122 (N_3122,N_2963,N_2826);
or U3123 (N_3123,N_2967,N_2477);
and U3124 (N_3124,N_2761,N_2810);
nand U3125 (N_3125,N_2020,N_2469);
or U3126 (N_3126,N_2329,N_2478);
nor U3127 (N_3127,N_2486,N_2234);
and U3128 (N_3128,N_2175,N_2430);
or U3129 (N_3129,N_2751,N_2664);
nand U3130 (N_3130,N_2227,N_2696);
nor U3131 (N_3131,N_2555,N_2511);
and U3132 (N_3132,N_2533,N_2855);
nand U3133 (N_3133,N_2892,N_2101);
nor U3134 (N_3134,N_2360,N_2283);
or U3135 (N_3135,N_2971,N_2576);
or U3136 (N_3136,N_2438,N_2578);
nand U3137 (N_3137,N_2717,N_2678);
nand U3138 (N_3138,N_2255,N_2321);
and U3139 (N_3139,N_2821,N_2356);
nor U3140 (N_3140,N_2364,N_2119);
and U3141 (N_3141,N_2374,N_2461);
or U3142 (N_3142,N_2368,N_2658);
or U3143 (N_3143,N_2019,N_2706);
and U3144 (N_3144,N_2799,N_2051);
and U3145 (N_3145,N_2894,N_2552);
xnor U3146 (N_3146,N_2411,N_2992);
nand U3147 (N_3147,N_2831,N_2102);
and U3148 (N_3148,N_2947,N_2629);
or U3149 (N_3149,N_2836,N_2443);
nand U3150 (N_3150,N_2366,N_2388);
nor U3151 (N_3151,N_2435,N_2981);
nand U3152 (N_3152,N_2651,N_2401);
and U3153 (N_3153,N_2514,N_2094);
nor U3154 (N_3154,N_2649,N_2804);
nor U3155 (N_3155,N_2026,N_2509);
nand U3156 (N_3156,N_2990,N_2106);
nand U3157 (N_3157,N_2422,N_2249);
nand U3158 (N_3158,N_2405,N_2580);
nor U3159 (N_3159,N_2398,N_2502);
nor U3160 (N_3160,N_2588,N_2009);
nand U3161 (N_3161,N_2937,N_2380);
or U3162 (N_3162,N_2906,N_2727);
nand U3163 (N_3163,N_2769,N_2748);
nand U3164 (N_3164,N_2688,N_2236);
nor U3165 (N_3165,N_2383,N_2500);
nand U3166 (N_3166,N_2410,N_2532);
xor U3167 (N_3167,N_2448,N_2248);
xor U3168 (N_3168,N_2803,N_2976);
or U3169 (N_3169,N_2218,N_2637);
nor U3170 (N_3170,N_2286,N_2551);
and U3171 (N_3171,N_2585,N_2053);
and U3172 (N_3172,N_2887,N_2833);
nor U3173 (N_3173,N_2691,N_2721);
or U3174 (N_3174,N_2090,N_2934);
nor U3175 (N_3175,N_2654,N_2202);
and U3176 (N_3176,N_2989,N_2332);
and U3177 (N_3177,N_2457,N_2539);
nand U3178 (N_3178,N_2882,N_2290);
and U3179 (N_3179,N_2946,N_2577);
nor U3180 (N_3180,N_2067,N_2697);
or U3181 (N_3181,N_2216,N_2318);
and U3182 (N_3182,N_2757,N_2015);
nor U3183 (N_3183,N_2304,N_2437);
xor U3184 (N_3184,N_2386,N_2843);
nand U3185 (N_3185,N_2907,N_2560);
or U3186 (N_3186,N_2455,N_2729);
nor U3187 (N_3187,N_2495,N_2818);
and U3188 (N_3188,N_2518,N_2562);
or U3189 (N_3189,N_2546,N_2116);
and U3190 (N_3190,N_2434,N_2280);
nor U3191 (N_3191,N_2921,N_2226);
nand U3192 (N_3192,N_2764,N_2681);
and U3193 (N_3193,N_2943,N_2523);
and U3194 (N_3194,N_2439,N_2703);
nand U3195 (N_3195,N_2942,N_2979);
or U3196 (N_3196,N_2129,N_2404);
nor U3197 (N_3197,N_2066,N_2324);
and U3198 (N_3198,N_2653,N_2805);
nand U3199 (N_3199,N_2919,N_2197);
and U3200 (N_3200,N_2722,N_2001);
or U3201 (N_3201,N_2309,N_2994);
and U3202 (N_3202,N_2526,N_2928);
and U3203 (N_3203,N_2608,N_2507);
xnor U3204 (N_3204,N_2151,N_2903);
nand U3205 (N_3205,N_2628,N_2224);
nor U3206 (N_3206,N_2701,N_2025);
nand U3207 (N_3207,N_2736,N_2582);
or U3208 (N_3208,N_2070,N_2734);
or U3209 (N_3209,N_2482,N_2397);
and U3210 (N_3210,N_2827,N_2966);
nand U3211 (N_3211,N_2379,N_2820);
nand U3212 (N_3212,N_2516,N_2269);
or U3213 (N_3213,N_2340,N_2145);
and U3214 (N_3214,N_2973,N_2350);
nor U3215 (N_3215,N_2035,N_2389);
nand U3216 (N_3216,N_2361,N_2331);
nor U3217 (N_3217,N_2755,N_2999);
nand U3218 (N_3218,N_2858,N_2221);
nand U3219 (N_3219,N_2813,N_2785);
or U3220 (N_3220,N_2096,N_2911);
or U3221 (N_3221,N_2162,N_2313);
nand U3222 (N_3222,N_2168,N_2135);
nor U3223 (N_3223,N_2148,N_2844);
and U3224 (N_3224,N_2932,N_2626);
and U3225 (N_3225,N_2195,N_2680);
or U3226 (N_3226,N_2874,N_2534);
and U3227 (N_3227,N_2071,N_2058);
nor U3228 (N_3228,N_2817,N_2563);
and U3229 (N_3229,N_2190,N_2545);
or U3230 (N_3230,N_2558,N_2872);
and U3231 (N_3231,N_2267,N_2548);
or U3232 (N_3232,N_2845,N_2904);
xnor U3233 (N_3233,N_2307,N_2938);
xor U3234 (N_3234,N_2308,N_2186);
nand U3235 (N_3235,N_2951,N_2095);
nand U3236 (N_3236,N_2760,N_2046);
and U3237 (N_3237,N_2052,N_2763);
nor U3238 (N_3238,N_2416,N_2542);
and U3239 (N_3239,N_2948,N_2017);
and U3240 (N_3240,N_2230,N_2268);
or U3241 (N_3241,N_2692,N_2334);
nand U3242 (N_3242,N_2811,N_2432);
or U3243 (N_3243,N_2442,N_2876);
xor U3244 (N_3244,N_2352,N_2605);
nand U3245 (N_3245,N_2640,N_2032);
or U3246 (N_3246,N_2745,N_2896);
nand U3247 (N_3247,N_2851,N_2082);
nand U3248 (N_3248,N_2737,N_2834);
nor U3249 (N_3249,N_2615,N_2295);
and U3250 (N_3250,N_2793,N_2744);
nor U3251 (N_3251,N_2217,N_2581);
and U3252 (N_3252,N_2421,N_2320);
and U3253 (N_3253,N_2459,N_2010);
or U3254 (N_3254,N_2425,N_2464);
nor U3255 (N_3255,N_2099,N_2568);
nor U3256 (N_3256,N_2074,N_2292);
or U3257 (N_3257,N_2417,N_2393);
and U3258 (N_3258,N_2927,N_2263);
or U3259 (N_3259,N_2530,N_2801);
nor U3260 (N_3260,N_2376,N_2497);
and U3261 (N_3261,N_2011,N_2456);
nor U3262 (N_3262,N_2322,N_2752);
nor U3263 (N_3263,N_2165,N_2501);
nor U3264 (N_3264,N_2191,N_2342);
and U3265 (N_3265,N_2244,N_2144);
or U3266 (N_3266,N_2969,N_2392);
and U3267 (N_3267,N_2554,N_2312);
or U3268 (N_3268,N_2616,N_2655);
nor U3269 (N_3269,N_2193,N_2491);
xnor U3270 (N_3270,N_2347,N_2970);
and U3271 (N_3271,N_2529,N_2450);
nand U3272 (N_3272,N_2709,N_2210);
nand U3273 (N_3273,N_2541,N_2122);
or U3274 (N_3274,N_2353,N_2754);
nand U3275 (N_3275,N_2213,N_2770);
nand U3276 (N_3276,N_2084,N_2128);
nor U3277 (N_3277,N_2285,N_2583);
nor U3278 (N_3278,N_2893,N_2228);
xnor U3279 (N_3279,N_2261,N_2864);
nor U3280 (N_3280,N_2370,N_2220);
and U3281 (N_3281,N_2515,N_2384);
nor U3282 (N_3282,N_2738,N_2944);
or U3283 (N_3283,N_2490,N_2107);
nor U3284 (N_3284,N_2189,N_2198);
nor U3285 (N_3285,N_2746,N_2279);
nand U3286 (N_3286,N_2723,N_2354);
and U3287 (N_3287,N_2662,N_2902);
and U3288 (N_3288,N_2781,N_2345);
nor U3289 (N_3289,N_2905,N_2695);
nand U3290 (N_3290,N_2593,N_2111);
nand U3291 (N_3291,N_2957,N_2142);
or U3292 (N_3292,N_2378,N_2540);
or U3293 (N_3293,N_2720,N_2488);
and U3294 (N_3294,N_2787,N_2642);
and U3295 (N_3295,N_2901,N_2779);
and U3296 (N_3296,N_2004,N_2108);
nand U3297 (N_3297,N_2297,N_2566);
or U3298 (N_3298,N_2885,N_2574);
nor U3299 (N_3299,N_2636,N_2579);
nor U3300 (N_3300,N_2634,N_2143);
and U3301 (N_3301,N_2359,N_2259);
nor U3302 (N_3302,N_2264,N_2631);
nand U3303 (N_3303,N_2114,N_2671);
nor U3304 (N_3304,N_2365,N_2204);
nand U3305 (N_3305,N_2113,N_2996);
and U3306 (N_3306,N_2869,N_2756);
nand U3307 (N_3307,N_2693,N_2390);
nand U3308 (N_3308,N_2713,N_2607);
nor U3309 (N_3309,N_2556,N_2257);
or U3310 (N_3310,N_2570,N_2073);
nand U3311 (N_3311,N_2079,N_2271);
nor U3312 (N_3312,N_2823,N_2110);
or U3313 (N_3313,N_2044,N_2527);
xor U3314 (N_3314,N_2049,N_2800);
xnor U3315 (N_3315,N_2569,N_2043);
nand U3316 (N_3316,N_2089,N_2387);
xnor U3317 (N_3317,N_2632,N_2930);
nand U3318 (N_3318,N_2041,N_2852);
and U3319 (N_3319,N_2841,N_2620);
nor U3320 (N_3320,N_2925,N_2510);
nand U3321 (N_3321,N_2033,N_2498);
nand U3322 (N_3322,N_2022,N_2098);
or U3323 (N_3323,N_2048,N_2949);
nor U3324 (N_3324,N_2715,N_2336);
nand U3325 (N_3325,N_2561,N_2699);
and U3326 (N_3326,N_2358,N_2091);
and U3327 (N_3327,N_2741,N_2293);
or U3328 (N_3328,N_2468,N_2176);
nor U3329 (N_3329,N_2339,N_2668);
nor U3330 (N_3330,N_2847,N_2211);
nand U3331 (N_3331,N_2660,N_2531);
or U3332 (N_3332,N_2121,N_2112);
or U3333 (N_3333,N_2480,N_2830);
or U3334 (N_3334,N_2553,N_2447);
or U3335 (N_3335,N_2922,N_2000);
nand U3336 (N_3336,N_2174,N_2420);
or U3337 (N_3337,N_2391,N_2325);
and U3338 (N_3338,N_2750,N_2077);
or U3339 (N_3339,N_2212,N_2466);
nand U3340 (N_3340,N_2171,N_2505);
or U3341 (N_3341,N_2407,N_2867);
or U3342 (N_3342,N_2700,N_2972);
nand U3343 (N_3343,N_2115,N_2163);
or U3344 (N_3344,N_2061,N_2743);
and U3345 (N_3345,N_2282,N_2808);
nand U3346 (N_3346,N_2275,N_2832);
nand U3347 (N_3347,N_2330,N_2702);
nor U3348 (N_3348,N_2774,N_2912);
or U3349 (N_3349,N_2986,N_2900);
nor U3350 (N_3350,N_2650,N_2003);
and U3351 (N_3351,N_2712,N_2272);
nand U3352 (N_3352,N_2954,N_2589);
and U3353 (N_3353,N_2258,N_2601);
nand U3354 (N_3354,N_2229,N_2005);
nand U3355 (N_3355,N_2725,N_2740);
nor U3356 (N_3356,N_2247,N_2188);
xor U3357 (N_3357,N_2402,N_2104);
nor U3358 (N_3358,N_2880,N_2433);
or U3359 (N_3359,N_2806,N_2848);
xnor U3360 (N_3360,N_2837,N_2300);
nand U3361 (N_3361,N_2038,N_2240);
nor U3362 (N_3362,N_2639,N_2233);
and U3363 (N_3363,N_2453,N_2068);
and U3364 (N_3364,N_2638,N_2474);
and U3365 (N_3365,N_2594,N_2109);
or U3366 (N_3366,N_2223,N_2842);
nand U3367 (N_3367,N_2016,N_2471);
nand U3368 (N_3368,N_2031,N_2064);
or U3369 (N_3369,N_2045,N_2596);
nand U3370 (N_3370,N_2980,N_2630);
or U3371 (N_3371,N_2666,N_2707);
or U3372 (N_3372,N_2778,N_2396);
nor U3373 (N_3373,N_2612,N_2462);
xor U3374 (N_3374,N_2623,N_2239);
nand U3375 (N_3375,N_2338,N_2782);
and U3376 (N_3376,N_2157,N_2215);
nand U3377 (N_3377,N_2134,N_2120);
nand U3378 (N_3378,N_2875,N_2592);
nand U3379 (N_3379,N_2908,N_2103);
and U3380 (N_3380,N_2889,N_2475);
or U3381 (N_3381,N_2888,N_2918);
nor U3382 (N_3382,N_2235,N_2635);
nor U3383 (N_3383,N_2431,N_2449);
and U3384 (N_3384,N_2910,N_2424);
and U3385 (N_3385,N_2926,N_2538);
nor U3386 (N_3386,N_2536,N_2173);
and U3387 (N_3387,N_2337,N_2773);
or U3388 (N_3388,N_2825,N_2508);
and U3389 (N_3389,N_2960,N_2802);
nor U3390 (N_3390,N_2775,N_2395);
nand U3391 (N_3391,N_2771,N_2891);
xor U3392 (N_3392,N_2023,N_2034);
xnor U3393 (N_3393,N_2835,N_2021);
or U3394 (N_3394,N_2371,N_2672);
nand U3395 (N_3395,N_2595,N_2669);
nand U3396 (N_3396,N_2985,N_2940);
nand U3397 (N_3397,N_2428,N_2427);
xnor U3398 (N_3398,N_2100,N_2557);
and U3399 (N_3399,N_2161,N_2730);
or U3400 (N_3400,N_2953,N_2083);
nor U3401 (N_3401,N_2059,N_2203);
and U3402 (N_3402,N_2544,N_2853);
nand U3403 (N_3403,N_2768,N_2187);
and U3404 (N_3404,N_2238,N_2549);
and U3405 (N_3405,N_2452,N_2346);
and U3406 (N_3406,N_2451,N_2816);
or U3407 (N_3407,N_2242,N_2008);
and U3408 (N_3408,N_2621,N_2978);
or U3409 (N_3409,N_2311,N_2597);
and U3410 (N_3410,N_2105,N_2047);
nor U3411 (N_3411,N_2458,N_2155);
xor U3412 (N_3412,N_2945,N_2408);
or U3413 (N_3413,N_2494,N_2567);
nand U3414 (N_3414,N_2192,N_2054);
nand U3415 (N_3415,N_2791,N_2819);
nor U3416 (N_3416,N_2470,N_2080);
nor U3417 (N_3417,N_2013,N_2917);
or U3418 (N_3418,N_2343,N_2419);
nand U3419 (N_3419,N_2287,N_2964);
or U3420 (N_3420,N_2207,N_2674);
and U3421 (N_3421,N_2341,N_2839);
nand U3422 (N_3422,N_2254,N_2444);
or U3423 (N_3423,N_2296,N_2310);
or U3424 (N_3424,N_2123,N_2604);
nand U3425 (N_3425,N_2777,N_2670);
or U3426 (N_3426,N_2065,N_2790);
and U3427 (N_3427,N_2914,N_2895);
or U3428 (N_3428,N_2487,N_2733);
or U3429 (N_3429,N_2409,N_2446);
nor U3430 (N_3430,N_2742,N_2705);
nand U3431 (N_3431,N_2766,N_2602);
nor U3432 (N_3432,N_2975,N_2245);
xor U3433 (N_3433,N_2647,N_2850);
nand U3434 (N_3434,N_2125,N_2246);
or U3435 (N_3435,N_2753,N_2854);
nand U3436 (N_3436,N_2749,N_2028);
nor U3437 (N_3437,N_2572,N_2274);
or U3438 (N_3438,N_2262,N_2587);
nand U3439 (N_3439,N_2315,N_2298);
nor U3440 (N_3440,N_2732,N_2860);
or U3441 (N_3441,N_2796,N_2788);
nand U3442 (N_3442,N_2676,N_2127);
xor U3443 (N_3443,N_2714,N_2881);
nand U3444 (N_3444,N_2719,N_2513);
and U3445 (N_3445,N_2069,N_2362);
nand U3446 (N_3446,N_2899,N_2933);
or U3447 (N_3447,N_2256,N_2429);
nor U3448 (N_3448,N_2913,N_2139);
nor U3449 (N_3449,N_2492,N_2180);
nand U3450 (N_3450,N_2289,N_2316);
or U3451 (N_3451,N_2243,N_2306);
and U3452 (N_3452,N_2333,N_2375);
nor U3453 (N_3453,N_2565,N_2840);
xor U3454 (N_3454,N_2504,N_2724);
and U3455 (N_3455,N_2472,N_2199);
or U3456 (N_3456,N_2524,N_2525);
nor U3457 (N_3457,N_2915,N_2993);
nand U3458 (N_3458,N_2795,N_2169);
and U3459 (N_3459,N_2609,N_2797);
and U3460 (N_3460,N_2441,N_2164);
nor U3461 (N_3461,N_2772,N_2117);
nand U3462 (N_3462,N_2898,N_2950);
nand U3463 (N_3463,N_2277,N_2991);
nor U3464 (N_3464,N_2463,N_2627);
and U3465 (N_3465,N_2036,N_2677);
and U3466 (N_3466,N_2426,N_2178);
nor U3467 (N_3467,N_2956,N_2288);
nor U3468 (N_3468,N_2591,N_2027);
nor U3469 (N_3469,N_2694,N_2493);
or U3470 (N_3470,N_2029,N_2181);
nand U3471 (N_3471,N_2146,N_2862);
nand U3472 (N_3472,N_2988,N_2291);
nand U3473 (N_3473,N_2939,N_2625);
nand U3474 (N_3474,N_2185,N_2085);
nor U3475 (N_3475,N_2865,N_2646);
and U3476 (N_3476,N_2057,N_2814);
nor U3477 (N_3477,N_2149,N_2131);
nor U3478 (N_3478,N_2150,N_2974);
or U3479 (N_3479,N_2273,N_2183);
and U3480 (N_3480,N_2543,N_2219);
nand U3481 (N_3481,N_2078,N_2863);
or U3482 (N_3482,N_2118,N_2698);
nor U3483 (N_3483,N_2838,N_2728);
nor U3484 (N_3484,N_2093,N_2302);
and U3485 (N_3485,N_2711,N_2684);
nand U3486 (N_3486,N_2955,N_2363);
and U3487 (N_3487,N_2133,N_2314);
nor U3488 (N_3488,N_2208,N_2659);
and U3489 (N_3489,N_2776,N_2385);
and U3490 (N_3490,N_2030,N_2759);
nor U3491 (N_3491,N_2403,N_2731);
nand U3492 (N_3492,N_2206,N_2586);
nor U3493 (N_3493,N_2182,N_2250);
and U3494 (N_3494,N_2656,N_2682);
or U3495 (N_3495,N_2348,N_2018);
nor U3496 (N_3496,N_2584,N_2222);
xnor U3497 (N_3497,N_2710,N_2520);
or U3498 (N_3498,N_2983,N_2959);
nand U3499 (N_3499,N_2413,N_2652);
xor U3500 (N_3500,N_2259,N_2665);
nand U3501 (N_3501,N_2894,N_2867);
or U3502 (N_3502,N_2454,N_2046);
or U3503 (N_3503,N_2727,N_2355);
nand U3504 (N_3504,N_2002,N_2731);
nand U3505 (N_3505,N_2177,N_2308);
and U3506 (N_3506,N_2970,N_2896);
or U3507 (N_3507,N_2624,N_2541);
or U3508 (N_3508,N_2075,N_2631);
nor U3509 (N_3509,N_2710,N_2473);
nand U3510 (N_3510,N_2907,N_2943);
nor U3511 (N_3511,N_2872,N_2867);
nand U3512 (N_3512,N_2516,N_2643);
nor U3513 (N_3513,N_2855,N_2983);
or U3514 (N_3514,N_2446,N_2140);
nor U3515 (N_3515,N_2984,N_2252);
nor U3516 (N_3516,N_2743,N_2613);
nand U3517 (N_3517,N_2648,N_2061);
nor U3518 (N_3518,N_2745,N_2079);
nor U3519 (N_3519,N_2202,N_2972);
nor U3520 (N_3520,N_2841,N_2746);
nand U3521 (N_3521,N_2578,N_2163);
or U3522 (N_3522,N_2672,N_2978);
or U3523 (N_3523,N_2363,N_2433);
nor U3524 (N_3524,N_2568,N_2032);
and U3525 (N_3525,N_2892,N_2914);
nor U3526 (N_3526,N_2775,N_2260);
nor U3527 (N_3527,N_2893,N_2352);
or U3528 (N_3528,N_2216,N_2716);
and U3529 (N_3529,N_2872,N_2208);
and U3530 (N_3530,N_2204,N_2455);
or U3531 (N_3531,N_2996,N_2224);
nand U3532 (N_3532,N_2913,N_2108);
nor U3533 (N_3533,N_2175,N_2964);
nand U3534 (N_3534,N_2115,N_2807);
xnor U3535 (N_3535,N_2471,N_2487);
and U3536 (N_3536,N_2117,N_2423);
nand U3537 (N_3537,N_2204,N_2051);
nor U3538 (N_3538,N_2305,N_2703);
nor U3539 (N_3539,N_2257,N_2682);
or U3540 (N_3540,N_2094,N_2323);
or U3541 (N_3541,N_2895,N_2434);
or U3542 (N_3542,N_2224,N_2612);
nor U3543 (N_3543,N_2845,N_2956);
or U3544 (N_3544,N_2648,N_2546);
nor U3545 (N_3545,N_2395,N_2043);
nand U3546 (N_3546,N_2543,N_2675);
nand U3547 (N_3547,N_2532,N_2302);
and U3548 (N_3548,N_2150,N_2518);
nor U3549 (N_3549,N_2703,N_2101);
xnor U3550 (N_3550,N_2813,N_2965);
nand U3551 (N_3551,N_2949,N_2739);
nand U3552 (N_3552,N_2437,N_2977);
nor U3553 (N_3553,N_2340,N_2422);
nor U3554 (N_3554,N_2250,N_2917);
and U3555 (N_3555,N_2909,N_2275);
xor U3556 (N_3556,N_2851,N_2666);
nand U3557 (N_3557,N_2228,N_2381);
and U3558 (N_3558,N_2658,N_2915);
and U3559 (N_3559,N_2208,N_2743);
nor U3560 (N_3560,N_2570,N_2472);
nor U3561 (N_3561,N_2006,N_2060);
or U3562 (N_3562,N_2234,N_2875);
nand U3563 (N_3563,N_2011,N_2990);
nor U3564 (N_3564,N_2401,N_2933);
or U3565 (N_3565,N_2414,N_2157);
nand U3566 (N_3566,N_2195,N_2053);
xor U3567 (N_3567,N_2247,N_2535);
nor U3568 (N_3568,N_2461,N_2999);
xor U3569 (N_3569,N_2602,N_2622);
and U3570 (N_3570,N_2375,N_2573);
nand U3571 (N_3571,N_2788,N_2554);
and U3572 (N_3572,N_2067,N_2348);
nand U3573 (N_3573,N_2304,N_2517);
or U3574 (N_3574,N_2203,N_2727);
xor U3575 (N_3575,N_2412,N_2975);
nand U3576 (N_3576,N_2151,N_2385);
or U3577 (N_3577,N_2871,N_2595);
xnor U3578 (N_3578,N_2454,N_2088);
nand U3579 (N_3579,N_2833,N_2751);
or U3580 (N_3580,N_2215,N_2302);
nand U3581 (N_3581,N_2124,N_2321);
or U3582 (N_3582,N_2101,N_2707);
nand U3583 (N_3583,N_2223,N_2296);
xor U3584 (N_3584,N_2485,N_2905);
and U3585 (N_3585,N_2027,N_2041);
nand U3586 (N_3586,N_2473,N_2153);
nor U3587 (N_3587,N_2976,N_2797);
xor U3588 (N_3588,N_2786,N_2022);
nand U3589 (N_3589,N_2028,N_2321);
nor U3590 (N_3590,N_2274,N_2290);
or U3591 (N_3591,N_2463,N_2797);
nor U3592 (N_3592,N_2256,N_2693);
nand U3593 (N_3593,N_2807,N_2852);
nor U3594 (N_3594,N_2601,N_2109);
xor U3595 (N_3595,N_2593,N_2259);
xnor U3596 (N_3596,N_2400,N_2656);
and U3597 (N_3597,N_2226,N_2038);
xnor U3598 (N_3598,N_2663,N_2080);
nand U3599 (N_3599,N_2117,N_2249);
and U3600 (N_3600,N_2320,N_2831);
nor U3601 (N_3601,N_2308,N_2721);
nor U3602 (N_3602,N_2223,N_2478);
and U3603 (N_3603,N_2763,N_2857);
or U3604 (N_3604,N_2951,N_2210);
nand U3605 (N_3605,N_2746,N_2213);
nor U3606 (N_3606,N_2514,N_2223);
nand U3607 (N_3607,N_2926,N_2420);
nor U3608 (N_3608,N_2171,N_2203);
nand U3609 (N_3609,N_2386,N_2068);
or U3610 (N_3610,N_2241,N_2556);
or U3611 (N_3611,N_2459,N_2915);
or U3612 (N_3612,N_2659,N_2773);
nor U3613 (N_3613,N_2616,N_2748);
or U3614 (N_3614,N_2765,N_2940);
nand U3615 (N_3615,N_2035,N_2173);
nor U3616 (N_3616,N_2657,N_2000);
nand U3617 (N_3617,N_2059,N_2715);
and U3618 (N_3618,N_2464,N_2018);
or U3619 (N_3619,N_2812,N_2215);
nand U3620 (N_3620,N_2033,N_2095);
nand U3621 (N_3621,N_2028,N_2301);
nor U3622 (N_3622,N_2099,N_2806);
xnor U3623 (N_3623,N_2515,N_2731);
nand U3624 (N_3624,N_2209,N_2180);
nand U3625 (N_3625,N_2522,N_2437);
or U3626 (N_3626,N_2789,N_2073);
xnor U3627 (N_3627,N_2141,N_2798);
nand U3628 (N_3628,N_2289,N_2934);
nand U3629 (N_3629,N_2260,N_2800);
nor U3630 (N_3630,N_2111,N_2628);
or U3631 (N_3631,N_2295,N_2992);
nand U3632 (N_3632,N_2762,N_2148);
or U3633 (N_3633,N_2629,N_2111);
xnor U3634 (N_3634,N_2630,N_2735);
and U3635 (N_3635,N_2494,N_2165);
or U3636 (N_3636,N_2791,N_2633);
nand U3637 (N_3637,N_2096,N_2473);
and U3638 (N_3638,N_2465,N_2087);
nor U3639 (N_3639,N_2953,N_2586);
or U3640 (N_3640,N_2658,N_2474);
or U3641 (N_3641,N_2399,N_2148);
nand U3642 (N_3642,N_2571,N_2001);
and U3643 (N_3643,N_2693,N_2289);
and U3644 (N_3644,N_2599,N_2165);
or U3645 (N_3645,N_2001,N_2660);
and U3646 (N_3646,N_2352,N_2752);
nand U3647 (N_3647,N_2578,N_2486);
nand U3648 (N_3648,N_2973,N_2395);
or U3649 (N_3649,N_2905,N_2497);
or U3650 (N_3650,N_2306,N_2152);
or U3651 (N_3651,N_2281,N_2910);
nor U3652 (N_3652,N_2791,N_2103);
or U3653 (N_3653,N_2081,N_2610);
nand U3654 (N_3654,N_2087,N_2108);
and U3655 (N_3655,N_2230,N_2333);
nand U3656 (N_3656,N_2387,N_2444);
nand U3657 (N_3657,N_2842,N_2347);
nor U3658 (N_3658,N_2455,N_2660);
nand U3659 (N_3659,N_2889,N_2505);
nand U3660 (N_3660,N_2266,N_2567);
or U3661 (N_3661,N_2479,N_2104);
or U3662 (N_3662,N_2827,N_2267);
and U3663 (N_3663,N_2580,N_2848);
nor U3664 (N_3664,N_2128,N_2386);
xnor U3665 (N_3665,N_2808,N_2309);
nand U3666 (N_3666,N_2288,N_2944);
and U3667 (N_3667,N_2223,N_2141);
nand U3668 (N_3668,N_2415,N_2578);
nor U3669 (N_3669,N_2458,N_2006);
and U3670 (N_3670,N_2585,N_2235);
or U3671 (N_3671,N_2599,N_2637);
nand U3672 (N_3672,N_2905,N_2920);
and U3673 (N_3673,N_2786,N_2398);
xor U3674 (N_3674,N_2907,N_2993);
nor U3675 (N_3675,N_2474,N_2501);
nand U3676 (N_3676,N_2040,N_2496);
or U3677 (N_3677,N_2683,N_2707);
and U3678 (N_3678,N_2475,N_2051);
nor U3679 (N_3679,N_2148,N_2840);
nand U3680 (N_3680,N_2304,N_2651);
nand U3681 (N_3681,N_2110,N_2347);
nor U3682 (N_3682,N_2062,N_2843);
nand U3683 (N_3683,N_2140,N_2962);
nand U3684 (N_3684,N_2738,N_2332);
or U3685 (N_3685,N_2448,N_2377);
nand U3686 (N_3686,N_2185,N_2648);
and U3687 (N_3687,N_2186,N_2402);
or U3688 (N_3688,N_2706,N_2737);
and U3689 (N_3689,N_2781,N_2401);
xnor U3690 (N_3690,N_2238,N_2648);
nand U3691 (N_3691,N_2781,N_2994);
and U3692 (N_3692,N_2240,N_2287);
nor U3693 (N_3693,N_2903,N_2509);
or U3694 (N_3694,N_2314,N_2820);
or U3695 (N_3695,N_2581,N_2484);
nand U3696 (N_3696,N_2564,N_2395);
nor U3697 (N_3697,N_2364,N_2547);
and U3698 (N_3698,N_2736,N_2487);
nand U3699 (N_3699,N_2976,N_2030);
or U3700 (N_3700,N_2440,N_2180);
nand U3701 (N_3701,N_2088,N_2922);
xor U3702 (N_3702,N_2713,N_2784);
nand U3703 (N_3703,N_2079,N_2615);
or U3704 (N_3704,N_2019,N_2683);
or U3705 (N_3705,N_2077,N_2274);
or U3706 (N_3706,N_2418,N_2130);
or U3707 (N_3707,N_2734,N_2193);
nand U3708 (N_3708,N_2575,N_2350);
nor U3709 (N_3709,N_2436,N_2779);
xor U3710 (N_3710,N_2653,N_2837);
nand U3711 (N_3711,N_2025,N_2403);
or U3712 (N_3712,N_2250,N_2903);
nand U3713 (N_3713,N_2168,N_2790);
nor U3714 (N_3714,N_2087,N_2454);
nand U3715 (N_3715,N_2746,N_2996);
nand U3716 (N_3716,N_2921,N_2420);
nor U3717 (N_3717,N_2851,N_2447);
xnor U3718 (N_3718,N_2046,N_2724);
and U3719 (N_3719,N_2464,N_2653);
nor U3720 (N_3720,N_2974,N_2462);
nor U3721 (N_3721,N_2595,N_2830);
nand U3722 (N_3722,N_2010,N_2843);
nand U3723 (N_3723,N_2795,N_2701);
and U3724 (N_3724,N_2094,N_2048);
nor U3725 (N_3725,N_2963,N_2891);
nand U3726 (N_3726,N_2524,N_2019);
or U3727 (N_3727,N_2723,N_2443);
nor U3728 (N_3728,N_2420,N_2382);
or U3729 (N_3729,N_2566,N_2492);
nor U3730 (N_3730,N_2348,N_2204);
nor U3731 (N_3731,N_2031,N_2654);
nand U3732 (N_3732,N_2696,N_2087);
nor U3733 (N_3733,N_2846,N_2856);
xnor U3734 (N_3734,N_2869,N_2617);
nor U3735 (N_3735,N_2054,N_2393);
nor U3736 (N_3736,N_2412,N_2022);
or U3737 (N_3737,N_2631,N_2326);
nand U3738 (N_3738,N_2139,N_2302);
nor U3739 (N_3739,N_2016,N_2303);
or U3740 (N_3740,N_2787,N_2260);
nand U3741 (N_3741,N_2661,N_2691);
nor U3742 (N_3742,N_2527,N_2121);
nand U3743 (N_3743,N_2173,N_2915);
xnor U3744 (N_3744,N_2329,N_2287);
nor U3745 (N_3745,N_2749,N_2175);
and U3746 (N_3746,N_2101,N_2979);
xor U3747 (N_3747,N_2514,N_2074);
nand U3748 (N_3748,N_2564,N_2285);
nor U3749 (N_3749,N_2093,N_2643);
or U3750 (N_3750,N_2418,N_2861);
and U3751 (N_3751,N_2157,N_2470);
xnor U3752 (N_3752,N_2819,N_2573);
and U3753 (N_3753,N_2184,N_2921);
nor U3754 (N_3754,N_2748,N_2680);
nor U3755 (N_3755,N_2667,N_2725);
nor U3756 (N_3756,N_2659,N_2634);
xor U3757 (N_3757,N_2665,N_2217);
nor U3758 (N_3758,N_2350,N_2018);
or U3759 (N_3759,N_2850,N_2865);
xor U3760 (N_3760,N_2269,N_2977);
or U3761 (N_3761,N_2128,N_2808);
or U3762 (N_3762,N_2795,N_2880);
and U3763 (N_3763,N_2813,N_2029);
nand U3764 (N_3764,N_2130,N_2046);
nor U3765 (N_3765,N_2727,N_2639);
and U3766 (N_3766,N_2925,N_2888);
nand U3767 (N_3767,N_2362,N_2827);
nor U3768 (N_3768,N_2819,N_2671);
nand U3769 (N_3769,N_2901,N_2333);
nor U3770 (N_3770,N_2613,N_2476);
nor U3771 (N_3771,N_2604,N_2736);
and U3772 (N_3772,N_2088,N_2892);
nand U3773 (N_3773,N_2631,N_2341);
or U3774 (N_3774,N_2141,N_2052);
nand U3775 (N_3775,N_2277,N_2945);
or U3776 (N_3776,N_2344,N_2333);
nor U3777 (N_3777,N_2506,N_2163);
nand U3778 (N_3778,N_2293,N_2039);
nand U3779 (N_3779,N_2270,N_2400);
or U3780 (N_3780,N_2881,N_2381);
nand U3781 (N_3781,N_2668,N_2191);
or U3782 (N_3782,N_2636,N_2858);
xor U3783 (N_3783,N_2963,N_2912);
nor U3784 (N_3784,N_2717,N_2418);
xor U3785 (N_3785,N_2641,N_2447);
nand U3786 (N_3786,N_2017,N_2445);
nand U3787 (N_3787,N_2901,N_2584);
nand U3788 (N_3788,N_2494,N_2199);
xor U3789 (N_3789,N_2518,N_2289);
nand U3790 (N_3790,N_2902,N_2422);
nor U3791 (N_3791,N_2953,N_2761);
or U3792 (N_3792,N_2570,N_2249);
nor U3793 (N_3793,N_2505,N_2546);
or U3794 (N_3794,N_2465,N_2893);
nand U3795 (N_3795,N_2578,N_2810);
and U3796 (N_3796,N_2806,N_2021);
and U3797 (N_3797,N_2766,N_2562);
nand U3798 (N_3798,N_2088,N_2982);
nand U3799 (N_3799,N_2455,N_2409);
nor U3800 (N_3800,N_2197,N_2761);
xnor U3801 (N_3801,N_2053,N_2078);
xnor U3802 (N_3802,N_2002,N_2493);
nand U3803 (N_3803,N_2580,N_2852);
nor U3804 (N_3804,N_2465,N_2634);
nor U3805 (N_3805,N_2623,N_2310);
and U3806 (N_3806,N_2815,N_2719);
nor U3807 (N_3807,N_2379,N_2721);
and U3808 (N_3808,N_2959,N_2963);
xnor U3809 (N_3809,N_2152,N_2186);
and U3810 (N_3810,N_2639,N_2451);
and U3811 (N_3811,N_2769,N_2787);
nor U3812 (N_3812,N_2734,N_2455);
or U3813 (N_3813,N_2968,N_2653);
or U3814 (N_3814,N_2813,N_2905);
or U3815 (N_3815,N_2212,N_2169);
or U3816 (N_3816,N_2854,N_2987);
and U3817 (N_3817,N_2299,N_2580);
and U3818 (N_3818,N_2436,N_2997);
or U3819 (N_3819,N_2352,N_2948);
nand U3820 (N_3820,N_2645,N_2958);
xor U3821 (N_3821,N_2263,N_2071);
or U3822 (N_3822,N_2604,N_2294);
and U3823 (N_3823,N_2562,N_2592);
or U3824 (N_3824,N_2773,N_2543);
nand U3825 (N_3825,N_2843,N_2944);
xor U3826 (N_3826,N_2562,N_2658);
nor U3827 (N_3827,N_2090,N_2533);
and U3828 (N_3828,N_2477,N_2675);
nor U3829 (N_3829,N_2026,N_2018);
or U3830 (N_3830,N_2963,N_2806);
xor U3831 (N_3831,N_2905,N_2078);
and U3832 (N_3832,N_2134,N_2904);
nor U3833 (N_3833,N_2245,N_2500);
nand U3834 (N_3834,N_2780,N_2569);
nor U3835 (N_3835,N_2868,N_2749);
xor U3836 (N_3836,N_2634,N_2556);
nand U3837 (N_3837,N_2122,N_2059);
and U3838 (N_3838,N_2243,N_2553);
and U3839 (N_3839,N_2437,N_2887);
and U3840 (N_3840,N_2046,N_2176);
and U3841 (N_3841,N_2606,N_2128);
nand U3842 (N_3842,N_2949,N_2414);
xnor U3843 (N_3843,N_2783,N_2192);
nor U3844 (N_3844,N_2537,N_2506);
nand U3845 (N_3845,N_2294,N_2210);
nand U3846 (N_3846,N_2522,N_2796);
nand U3847 (N_3847,N_2203,N_2535);
and U3848 (N_3848,N_2445,N_2102);
nor U3849 (N_3849,N_2435,N_2024);
xor U3850 (N_3850,N_2700,N_2609);
and U3851 (N_3851,N_2416,N_2898);
nand U3852 (N_3852,N_2529,N_2742);
nor U3853 (N_3853,N_2737,N_2358);
xnor U3854 (N_3854,N_2053,N_2320);
nand U3855 (N_3855,N_2983,N_2354);
or U3856 (N_3856,N_2789,N_2456);
nand U3857 (N_3857,N_2865,N_2493);
nand U3858 (N_3858,N_2084,N_2702);
nand U3859 (N_3859,N_2502,N_2785);
nor U3860 (N_3860,N_2106,N_2531);
or U3861 (N_3861,N_2918,N_2081);
and U3862 (N_3862,N_2441,N_2439);
nor U3863 (N_3863,N_2127,N_2185);
nand U3864 (N_3864,N_2020,N_2582);
and U3865 (N_3865,N_2709,N_2030);
nand U3866 (N_3866,N_2671,N_2834);
nor U3867 (N_3867,N_2269,N_2232);
xnor U3868 (N_3868,N_2363,N_2869);
and U3869 (N_3869,N_2043,N_2235);
nand U3870 (N_3870,N_2450,N_2699);
nor U3871 (N_3871,N_2789,N_2123);
nor U3872 (N_3872,N_2907,N_2106);
or U3873 (N_3873,N_2676,N_2341);
and U3874 (N_3874,N_2775,N_2991);
or U3875 (N_3875,N_2697,N_2155);
xnor U3876 (N_3876,N_2499,N_2503);
and U3877 (N_3877,N_2824,N_2060);
or U3878 (N_3878,N_2162,N_2657);
or U3879 (N_3879,N_2570,N_2946);
nand U3880 (N_3880,N_2371,N_2366);
and U3881 (N_3881,N_2549,N_2208);
nand U3882 (N_3882,N_2745,N_2987);
nor U3883 (N_3883,N_2858,N_2301);
and U3884 (N_3884,N_2509,N_2033);
or U3885 (N_3885,N_2846,N_2465);
and U3886 (N_3886,N_2416,N_2607);
nand U3887 (N_3887,N_2992,N_2578);
nor U3888 (N_3888,N_2744,N_2467);
nand U3889 (N_3889,N_2616,N_2165);
nand U3890 (N_3890,N_2808,N_2015);
or U3891 (N_3891,N_2847,N_2358);
nor U3892 (N_3892,N_2704,N_2711);
and U3893 (N_3893,N_2328,N_2106);
nand U3894 (N_3894,N_2544,N_2573);
and U3895 (N_3895,N_2575,N_2638);
and U3896 (N_3896,N_2413,N_2462);
nor U3897 (N_3897,N_2655,N_2743);
nor U3898 (N_3898,N_2214,N_2921);
nand U3899 (N_3899,N_2064,N_2763);
or U3900 (N_3900,N_2083,N_2299);
nor U3901 (N_3901,N_2456,N_2633);
nand U3902 (N_3902,N_2674,N_2071);
or U3903 (N_3903,N_2973,N_2991);
and U3904 (N_3904,N_2782,N_2387);
nand U3905 (N_3905,N_2057,N_2644);
nand U3906 (N_3906,N_2495,N_2432);
and U3907 (N_3907,N_2675,N_2448);
and U3908 (N_3908,N_2519,N_2558);
and U3909 (N_3909,N_2150,N_2216);
xnor U3910 (N_3910,N_2395,N_2965);
and U3911 (N_3911,N_2960,N_2943);
nand U3912 (N_3912,N_2340,N_2658);
nand U3913 (N_3913,N_2403,N_2575);
nand U3914 (N_3914,N_2042,N_2857);
or U3915 (N_3915,N_2459,N_2990);
and U3916 (N_3916,N_2629,N_2116);
nand U3917 (N_3917,N_2067,N_2536);
nand U3918 (N_3918,N_2891,N_2924);
nand U3919 (N_3919,N_2480,N_2834);
nor U3920 (N_3920,N_2351,N_2817);
nand U3921 (N_3921,N_2742,N_2002);
or U3922 (N_3922,N_2413,N_2578);
or U3923 (N_3923,N_2611,N_2323);
nor U3924 (N_3924,N_2495,N_2107);
nand U3925 (N_3925,N_2201,N_2383);
or U3926 (N_3926,N_2805,N_2973);
nand U3927 (N_3927,N_2497,N_2365);
or U3928 (N_3928,N_2448,N_2231);
xor U3929 (N_3929,N_2989,N_2288);
nand U3930 (N_3930,N_2326,N_2653);
nor U3931 (N_3931,N_2642,N_2970);
and U3932 (N_3932,N_2029,N_2739);
or U3933 (N_3933,N_2849,N_2810);
nand U3934 (N_3934,N_2951,N_2944);
nand U3935 (N_3935,N_2796,N_2977);
or U3936 (N_3936,N_2057,N_2692);
and U3937 (N_3937,N_2632,N_2348);
nand U3938 (N_3938,N_2620,N_2582);
nand U3939 (N_3939,N_2531,N_2098);
nor U3940 (N_3940,N_2669,N_2967);
nand U3941 (N_3941,N_2374,N_2888);
and U3942 (N_3942,N_2909,N_2463);
nor U3943 (N_3943,N_2323,N_2791);
nand U3944 (N_3944,N_2106,N_2740);
nor U3945 (N_3945,N_2233,N_2160);
nand U3946 (N_3946,N_2460,N_2204);
nor U3947 (N_3947,N_2269,N_2592);
and U3948 (N_3948,N_2798,N_2102);
or U3949 (N_3949,N_2481,N_2968);
xor U3950 (N_3950,N_2370,N_2290);
or U3951 (N_3951,N_2802,N_2315);
and U3952 (N_3952,N_2723,N_2136);
nand U3953 (N_3953,N_2222,N_2544);
nand U3954 (N_3954,N_2624,N_2469);
and U3955 (N_3955,N_2403,N_2091);
or U3956 (N_3956,N_2166,N_2104);
or U3957 (N_3957,N_2400,N_2700);
or U3958 (N_3958,N_2152,N_2840);
or U3959 (N_3959,N_2114,N_2947);
or U3960 (N_3960,N_2944,N_2040);
or U3961 (N_3961,N_2000,N_2092);
or U3962 (N_3962,N_2678,N_2978);
and U3963 (N_3963,N_2631,N_2940);
and U3964 (N_3964,N_2255,N_2200);
nand U3965 (N_3965,N_2629,N_2934);
and U3966 (N_3966,N_2377,N_2948);
xor U3967 (N_3967,N_2080,N_2212);
nor U3968 (N_3968,N_2735,N_2468);
or U3969 (N_3969,N_2133,N_2735);
and U3970 (N_3970,N_2937,N_2991);
and U3971 (N_3971,N_2017,N_2064);
nand U3972 (N_3972,N_2138,N_2843);
or U3973 (N_3973,N_2702,N_2390);
nand U3974 (N_3974,N_2398,N_2539);
and U3975 (N_3975,N_2164,N_2719);
and U3976 (N_3976,N_2764,N_2344);
or U3977 (N_3977,N_2455,N_2047);
or U3978 (N_3978,N_2857,N_2585);
xor U3979 (N_3979,N_2821,N_2024);
and U3980 (N_3980,N_2718,N_2028);
nand U3981 (N_3981,N_2735,N_2975);
and U3982 (N_3982,N_2281,N_2658);
or U3983 (N_3983,N_2989,N_2884);
nor U3984 (N_3984,N_2694,N_2960);
nand U3985 (N_3985,N_2641,N_2029);
or U3986 (N_3986,N_2931,N_2413);
nor U3987 (N_3987,N_2471,N_2637);
nand U3988 (N_3988,N_2867,N_2537);
or U3989 (N_3989,N_2619,N_2497);
or U3990 (N_3990,N_2406,N_2194);
or U3991 (N_3991,N_2427,N_2293);
or U3992 (N_3992,N_2261,N_2482);
and U3993 (N_3993,N_2607,N_2991);
and U3994 (N_3994,N_2400,N_2029);
nor U3995 (N_3995,N_2653,N_2027);
xnor U3996 (N_3996,N_2452,N_2820);
xor U3997 (N_3997,N_2453,N_2814);
nand U3998 (N_3998,N_2964,N_2331);
and U3999 (N_3999,N_2116,N_2715);
nor U4000 (N_4000,N_3195,N_3463);
nor U4001 (N_4001,N_3217,N_3082);
nor U4002 (N_4002,N_3087,N_3444);
xor U4003 (N_4003,N_3155,N_3038);
nand U4004 (N_4004,N_3852,N_3273);
and U4005 (N_4005,N_3141,N_3828);
or U4006 (N_4006,N_3146,N_3788);
and U4007 (N_4007,N_3533,N_3691);
and U4008 (N_4008,N_3968,N_3016);
nor U4009 (N_4009,N_3306,N_3292);
xor U4010 (N_4010,N_3561,N_3367);
nand U4011 (N_4011,N_3938,N_3687);
or U4012 (N_4012,N_3308,N_3879);
or U4013 (N_4013,N_3934,N_3536);
and U4014 (N_4014,N_3936,N_3895);
nor U4015 (N_4015,N_3291,N_3330);
or U4016 (N_4016,N_3889,N_3102);
and U4017 (N_4017,N_3211,N_3052);
xor U4018 (N_4018,N_3126,N_3707);
and U4019 (N_4019,N_3992,N_3605);
xnor U4020 (N_4020,N_3021,N_3452);
and U4021 (N_4021,N_3910,N_3476);
and U4022 (N_4022,N_3702,N_3805);
or U4023 (N_4023,N_3088,N_3675);
nand U4024 (N_4024,N_3401,N_3109);
or U4025 (N_4025,N_3315,N_3656);
or U4026 (N_4026,N_3012,N_3623);
nand U4027 (N_4027,N_3190,N_3985);
or U4028 (N_4028,N_3064,N_3447);
nor U4029 (N_4029,N_3795,N_3699);
nor U4030 (N_4030,N_3518,N_3836);
nor U4031 (N_4031,N_3056,N_3194);
xnor U4032 (N_4032,N_3201,N_3983);
and U4033 (N_4033,N_3744,N_3074);
or U4034 (N_4034,N_3681,N_3753);
nor U4035 (N_4035,N_3193,N_3551);
and U4036 (N_4036,N_3739,N_3418);
nor U4037 (N_4037,N_3133,N_3579);
and U4038 (N_4038,N_3804,N_3724);
or U4039 (N_4039,N_3178,N_3270);
nor U4040 (N_4040,N_3426,N_3034);
nor U4041 (N_4041,N_3116,N_3013);
or U4042 (N_4042,N_3337,N_3247);
xnor U4043 (N_4043,N_3888,N_3669);
or U4044 (N_4044,N_3776,N_3598);
and U4045 (N_4045,N_3479,N_3660);
and U4046 (N_4046,N_3617,N_3398);
nand U4047 (N_4047,N_3477,N_3670);
or U4048 (N_4048,N_3854,N_3348);
or U4049 (N_4049,N_3122,N_3483);
or U4050 (N_4050,N_3467,N_3297);
nand U4051 (N_4051,N_3131,N_3290);
and U4052 (N_4052,N_3906,N_3184);
and U4053 (N_4053,N_3372,N_3902);
nand U4054 (N_4054,N_3263,N_3345);
or U4055 (N_4055,N_3809,N_3180);
and U4056 (N_4056,N_3473,N_3898);
or U4057 (N_4057,N_3262,N_3731);
nand U4058 (N_4058,N_3487,N_3633);
and U4059 (N_4059,N_3559,N_3510);
nor U4060 (N_4060,N_3972,N_3912);
or U4061 (N_4061,N_3168,N_3358);
and U4062 (N_4062,N_3550,N_3838);
nor U4063 (N_4063,N_3755,N_3264);
and U4064 (N_4064,N_3875,N_3606);
nor U4065 (N_4065,N_3079,N_3908);
or U4066 (N_4066,N_3923,N_3918);
nand U4067 (N_4067,N_3090,N_3949);
and U4068 (N_4068,N_3349,N_3392);
nand U4069 (N_4069,N_3100,N_3406);
xnor U4070 (N_4070,N_3404,N_3111);
and U4071 (N_4071,N_3229,N_3973);
and U4072 (N_4072,N_3148,N_3864);
nand U4073 (N_4073,N_3176,N_3803);
nand U4074 (N_4074,N_3227,N_3932);
or U4075 (N_4075,N_3523,N_3431);
nand U4076 (N_4076,N_3611,N_3218);
and U4077 (N_4077,N_3407,N_3640);
and U4078 (N_4078,N_3981,N_3061);
and U4079 (N_4079,N_3583,N_3192);
nor U4080 (N_4080,N_3365,N_3482);
xnor U4081 (N_4081,N_3671,N_3204);
or U4082 (N_4082,N_3442,N_3999);
nand U4083 (N_4083,N_3465,N_3573);
and U4084 (N_4084,N_3959,N_3435);
nor U4085 (N_4085,N_3587,N_3894);
and U4086 (N_4086,N_3667,N_3811);
and U4087 (N_4087,N_3892,N_3443);
or U4088 (N_4088,N_3051,N_3784);
nor U4089 (N_4089,N_3872,N_3503);
xnor U4090 (N_4090,N_3553,N_3230);
nand U4091 (N_4091,N_3036,N_3083);
nor U4092 (N_4092,N_3493,N_3976);
nor U4093 (N_4093,N_3858,N_3314);
and U4094 (N_4094,N_3953,N_3585);
nor U4095 (N_4095,N_3271,N_3066);
and U4096 (N_4096,N_3831,N_3882);
or U4097 (N_4097,N_3272,N_3620);
or U4098 (N_4098,N_3848,N_3441);
xor U4099 (N_4099,N_3539,N_3351);
or U4100 (N_4100,N_3065,N_3245);
nor U4101 (N_4101,N_3387,N_3806);
nor U4102 (N_4102,N_3224,N_3929);
and U4103 (N_4103,N_3220,N_3377);
or U4104 (N_4104,N_3185,N_3323);
and U4105 (N_4105,N_3097,N_3887);
or U4106 (N_4106,N_3615,N_3039);
nand U4107 (N_4107,N_3866,N_3957);
nand U4108 (N_4108,N_3798,N_3198);
and U4109 (N_4109,N_3975,N_3708);
and U4110 (N_4110,N_3527,N_3495);
or U4111 (N_4111,N_3604,N_3233);
nor U4112 (N_4112,N_3873,N_3395);
and U4113 (N_4113,N_3943,N_3215);
or U4114 (N_4114,N_3931,N_3106);
nor U4115 (N_4115,N_3117,N_3746);
and U4116 (N_4116,N_3951,N_3678);
and U4117 (N_4117,N_3399,N_3686);
or U4118 (N_4118,N_3555,N_3375);
nand U4119 (N_4119,N_3967,N_3704);
nand U4120 (N_4120,N_3020,N_3715);
nand U4121 (N_4121,N_3995,N_3538);
nand U4122 (N_4122,N_3793,N_3797);
nor U4123 (N_4123,N_3517,N_3814);
and U4124 (N_4124,N_3305,N_3319);
nor U4125 (N_4125,N_3763,N_3733);
nor U4126 (N_4126,N_3842,N_3504);
xnor U4127 (N_4127,N_3352,N_3453);
nor U4128 (N_4128,N_3316,N_3214);
and U4129 (N_4129,N_3093,N_3607);
nand U4130 (N_4130,N_3693,N_3762);
and U4131 (N_4131,N_3400,N_3557);
xnor U4132 (N_4132,N_3528,N_3584);
nand U4133 (N_4133,N_3312,N_3274);
nor U4134 (N_4134,N_3252,N_3979);
or U4135 (N_4135,N_3490,N_3823);
and U4136 (N_4136,N_3022,N_3175);
and U4137 (N_4137,N_3451,N_3756);
or U4138 (N_4138,N_3129,N_3149);
and U4139 (N_4139,N_3718,N_3159);
and U4140 (N_4140,N_3904,N_3698);
or U4141 (N_4141,N_3840,N_3602);
nor U4142 (N_4142,N_3960,N_3549);
and U4143 (N_4143,N_3472,N_3621);
xnor U4144 (N_4144,N_3712,N_3903);
or U4145 (N_4145,N_3145,N_3388);
and U4146 (N_4146,N_3935,N_3046);
nor U4147 (N_4147,N_3260,N_3385);
xnor U4148 (N_4148,N_3091,N_3857);
and U4149 (N_4149,N_3354,N_3248);
and U4150 (N_4150,N_3727,N_3276);
and U4151 (N_4151,N_3015,N_3940);
nand U4152 (N_4152,N_3522,N_3474);
and U4153 (N_4153,N_3566,N_3662);
and U4154 (N_4154,N_3028,N_3160);
and U4155 (N_4155,N_3958,N_3657);
xor U4156 (N_4156,N_3807,N_3771);
and U4157 (N_4157,N_3464,N_3984);
and U4158 (N_4158,N_3648,N_3344);
nand U4159 (N_4159,N_3721,N_3361);
nand U4160 (N_4160,N_3757,N_3379);
nand U4161 (N_4161,N_3049,N_3471);
or U4162 (N_4162,N_3187,N_3360);
and U4163 (N_4163,N_3547,N_3208);
and U4164 (N_4164,N_3458,N_3210);
nor U4165 (N_4165,N_3537,N_3861);
nor U4166 (N_4166,N_3941,N_3868);
nor U4167 (N_4167,N_3334,N_3595);
or U4168 (N_4168,N_3989,N_3519);
nor U4169 (N_4169,N_3371,N_3173);
nand U4170 (N_4170,N_3780,N_3120);
or U4171 (N_4171,N_3832,N_3901);
or U4172 (N_4172,N_3688,N_3318);
and U4173 (N_4173,N_3608,N_3130);
nand U4174 (N_4174,N_3412,N_3513);
or U4175 (N_4175,N_3964,N_3563);
nor U4176 (N_4176,N_3156,N_3496);
or U4177 (N_4177,N_3042,N_3711);
and U4178 (N_4178,N_3679,N_3055);
nor U4179 (N_4179,N_3800,N_3884);
nor U4180 (N_4180,N_3096,N_3044);
or U4181 (N_4181,N_3256,N_3397);
xnor U4182 (N_4182,N_3860,N_3317);
nand U4183 (N_4183,N_3589,N_3965);
and U4184 (N_4184,N_3963,N_3103);
and U4185 (N_4185,N_3336,N_3642);
nand U4186 (N_4186,N_3877,N_3764);
or U4187 (N_4187,N_3845,N_3653);
nand U4188 (N_4188,N_3294,N_3209);
nor U4189 (N_4189,N_3134,N_3244);
and U4190 (N_4190,N_3729,N_3646);
xnor U4191 (N_4191,N_3356,N_3520);
or U4192 (N_4192,N_3535,N_3766);
nor U4193 (N_4193,N_3614,N_3694);
or U4194 (N_4194,N_3922,N_3783);
xnor U4195 (N_4195,N_3592,N_3683);
or U4196 (N_4196,N_3630,N_3541);
and U4197 (N_4197,N_3138,N_3622);
nand U4198 (N_4198,N_3081,N_3005);
or U4199 (N_4199,N_3424,N_3137);
and U4200 (N_4200,N_3110,N_3680);
or U4201 (N_4201,N_3768,N_3433);
and U4202 (N_4202,N_3706,N_3759);
and U4203 (N_4203,N_3213,N_3505);
nor U4204 (N_4204,N_3280,N_3971);
and U4205 (N_4205,N_3355,N_3597);
nand U4206 (N_4206,N_3534,N_3303);
or U4207 (N_4207,N_3859,N_3177);
and U4208 (N_4208,N_3728,N_3978);
xor U4209 (N_4209,N_3414,N_3121);
nor U4210 (N_4210,N_3825,N_3569);
and U4211 (N_4211,N_3144,N_3363);
and U4212 (N_4212,N_3499,N_3112);
and U4213 (N_4213,N_3885,N_3909);
or U4214 (N_4214,N_3413,N_3668);
nor U4215 (N_4215,N_3002,N_3147);
or U4216 (N_4216,N_3249,N_3659);
nand U4217 (N_4217,N_3251,N_3277);
nor U4218 (N_4218,N_3543,N_3509);
nor U4219 (N_4219,N_3455,N_3301);
nor U4220 (N_4220,N_3043,N_3332);
and U4221 (N_4221,N_3827,N_3059);
or U4222 (N_4222,N_3734,N_3037);
and U4223 (N_4223,N_3114,N_3461);
and U4224 (N_4224,N_3293,N_3078);
nor U4225 (N_4225,N_3339,N_3010);
and U4226 (N_4226,N_3639,N_3415);
xnor U4227 (N_4227,N_3874,N_3286);
and U4228 (N_4228,N_3063,N_3747);
or U4229 (N_4229,N_3370,N_3911);
and U4230 (N_4230,N_3516,N_3690);
nor U4231 (N_4231,N_3713,N_3599);
and U4232 (N_4232,N_3007,N_3239);
xnor U4233 (N_4233,N_3478,N_3710);
nor U4234 (N_4234,N_3024,N_3644);
nor U4235 (N_4235,N_3603,N_3641);
and U4236 (N_4236,N_3950,N_3207);
nor U4237 (N_4237,N_3779,N_3267);
or U4238 (N_4238,N_3636,N_3423);
nand U4239 (N_4239,N_3627,N_3626);
and U4240 (N_4240,N_3011,N_3778);
nand U4241 (N_4241,N_3824,N_3900);
and U4242 (N_4242,N_3933,N_3484);
xor U4243 (N_4243,N_3457,N_3115);
nor U4244 (N_4244,N_3761,N_3409);
or U4245 (N_4245,N_3427,N_3741);
or U4246 (N_4246,N_3946,N_3231);
nor U4247 (N_4247,N_3525,N_3158);
nand U4248 (N_4248,N_3925,N_3829);
or U4249 (N_4249,N_3228,N_3616);
xnor U4250 (N_4250,N_3266,N_3250);
nor U4251 (N_4251,N_3035,N_3440);
nand U4252 (N_4252,N_3930,N_3000);
nand U4253 (N_4253,N_3692,N_3919);
nand U4254 (N_4254,N_3677,N_3076);
and U4255 (N_4255,N_3311,N_3546);
nand U4256 (N_4256,N_3926,N_3309);
nor U4257 (N_4257,N_3770,N_3696);
nor U4258 (N_4258,N_3382,N_3890);
and U4259 (N_4259,N_3645,N_3003);
or U4260 (N_4260,N_3990,N_3335);
and U4261 (N_4261,N_3221,N_3058);
nor U4262 (N_4262,N_3855,N_3577);
nor U4263 (N_4263,N_3053,N_3099);
nor U4264 (N_4264,N_3456,N_3165);
nor U4265 (N_4265,N_3026,N_3593);
nand U4266 (N_4266,N_3665,N_3815);
xor U4267 (N_4267,N_3944,N_3637);
nand U4268 (N_4268,N_3402,N_3374);
nor U4269 (N_4269,N_3281,N_3284);
xnor U4270 (N_4270,N_3390,N_3353);
or U4271 (N_4271,N_3299,N_3086);
nand U4272 (N_4272,N_3647,N_3410);
xor U4273 (N_4273,N_3916,N_3222);
or U4274 (N_4274,N_3501,N_3568);
and U4275 (N_4275,N_3571,N_3773);
and U4276 (N_4276,N_3329,N_3181);
nor U4277 (N_4277,N_3977,N_3961);
and U4278 (N_4278,N_3253,N_3748);
nor U4279 (N_4279,N_3403,N_3853);
nand U4280 (N_4280,N_3655,N_3416);
nor U4281 (N_4281,N_3171,N_3167);
nor U4282 (N_4282,N_3774,N_3001);
nand U4283 (N_4283,N_3802,N_3462);
nor U4284 (N_4284,N_3142,N_3432);
or U4285 (N_4285,N_3196,N_3663);
nand U4286 (N_4286,N_3434,N_3069);
nor U4287 (N_4287,N_3969,N_3869);
or U4288 (N_4288,N_3749,N_3591);
and U4289 (N_4289,N_3428,N_3162);
and U4290 (N_4290,N_3880,N_3150);
or U4291 (N_4291,N_3542,N_3014);
or U4292 (N_4292,N_3140,N_3179);
and U4293 (N_4293,N_3450,N_3048);
nand U4294 (N_4294,N_3040,N_3532);
and U4295 (N_4295,N_3350,N_3275);
and U4296 (N_4296,N_3781,N_3841);
and U4297 (N_4297,N_3917,N_3008);
and U4298 (N_4298,N_3072,N_3170);
nor U4299 (N_4299,N_3369,N_3151);
and U4300 (N_4300,N_3760,N_3004);
nor U4301 (N_4301,N_3554,N_3937);
and U4302 (N_4302,N_3974,N_3886);
or U4303 (N_4303,N_3393,N_3676);
xnor U4304 (N_4304,N_3018,N_3526);
or U4305 (N_4305,N_3241,N_3684);
nor U4306 (N_4306,N_3135,N_3907);
and U4307 (N_4307,N_3666,N_3742);
and U4308 (N_4308,N_3552,N_3067);
nand U4309 (N_4309,N_3321,N_3674);
nor U4310 (N_4310,N_3300,N_3856);
or U4311 (N_4311,N_3320,N_3095);
xnor U4312 (N_4312,N_3512,N_3982);
nand U4313 (N_4313,N_3871,N_3792);
nand U4314 (N_4314,N_3590,N_3257);
and U4315 (N_4315,N_3327,N_3326);
and U4316 (N_4316,N_3826,N_3719);
nand U4317 (N_4317,N_3124,N_3835);
nor U4318 (N_4318,N_3153,N_3169);
nand U4319 (N_4319,N_3649,N_3313);
xor U4320 (N_4320,N_3796,N_3027);
nor U4321 (N_4321,N_3436,N_3524);
nand U4322 (N_4322,N_3485,N_3246);
and U4323 (N_4323,N_3980,N_3019);
nor U4324 (N_4324,N_3896,N_3629);
and U4325 (N_4325,N_3123,N_3928);
nand U4326 (N_4326,N_3071,N_3883);
or U4327 (N_4327,N_3325,N_3157);
and U4328 (N_4328,N_3785,N_3765);
nor U4329 (N_4329,N_3288,N_3628);
or U4330 (N_4330,N_3240,N_3575);
or U4331 (N_4331,N_3988,N_3689);
nand U4332 (N_4332,N_3047,N_3163);
and U4333 (N_4333,N_3651,N_3006);
nor U4334 (N_4334,N_3127,N_3394);
or U4335 (N_4335,N_3799,N_3791);
or U4336 (N_4336,N_3366,N_3128);
nor U4337 (N_4337,N_3787,N_3564);
and U4338 (N_4338,N_3673,N_3279);
nor U4339 (N_4339,N_3511,N_3962);
xnor U4340 (N_4340,N_3897,N_3740);
nor U4341 (N_4341,N_3234,N_3914);
nand U4342 (N_4342,N_3556,N_3986);
and U4343 (N_4343,N_3188,N_3255);
nor U4344 (N_4344,N_3948,N_3421);
nand U4345 (N_4345,N_3632,N_3998);
or U4346 (N_4346,N_3736,N_3488);
and U4347 (N_4347,N_3716,N_3023);
nor U4348 (N_4348,N_3031,N_3816);
nor U4349 (N_4349,N_3261,N_3212);
and U4350 (N_4350,N_3700,N_3068);
or U4351 (N_4351,N_3927,N_3030);
nor U4352 (N_4352,N_3152,N_3839);
nor U4353 (N_4353,N_3437,N_3189);
nor U4354 (N_4354,N_3343,N_3565);
nor U4355 (N_4355,N_3834,N_3610);
xnor U4356 (N_4356,N_3405,N_3243);
xnor U4357 (N_4357,N_3619,N_3658);
nor U4358 (N_4358,N_3775,N_3322);
and U4359 (N_4359,N_3506,N_3723);
and U4360 (N_4360,N_3391,N_3362);
nand U4361 (N_4361,N_3101,N_3143);
nand U4362 (N_4362,N_3430,N_3077);
and U4363 (N_4363,N_3705,N_3161);
nand U4364 (N_4364,N_3492,N_3481);
nand U4365 (N_4365,N_3235,N_3468);
and U4366 (N_4366,N_3205,N_3782);
nand U4367 (N_4367,N_3216,N_3567);
or U4368 (N_4368,N_3899,N_3576);
or U4369 (N_4369,N_3786,N_3062);
nor U4370 (N_4370,N_3638,N_3843);
xnor U4371 (N_4371,N_3480,N_3380);
nand U4372 (N_4372,N_3594,N_3324);
nor U4373 (N_4373,N_3737,N_3174);
nor U4374 (N_4374,N_3098,N_3844);
nor U4375 (N_4375,N_3454,N_3381);
nor U4376 (N_4376,N_3601,N_3050);
nand U4377 (N_4377,N_3199,N_3970);
xnor U4378 (N_4378,N_3794,N_3132);
nand U4379 (N_4379,N_3772,N_3119);
and U4380 (N_4380,N_3588,N_3994);
and U4381 (N_4381,N_3108,N_3225);
or U4382 (N_4382,N_3259,N_3738);
and U4383 (N_4383,N_3060,N_3905);
nand U4384 (N_4384,N_3341,N_3609);
and U4385 (N_4385,N_3219,N_3089);
or U4386 (N_4386,N_3265,N_3743);
nand U4387 (N_4387,N_3384,N_3878);
nor U4388 (N_4388,N_3701,N_3714);
or U4389 (N_4389,N_3833,N_3913);
nor U4390 (N_4390,N_3408,N_3769);
nor U4391 (N_4391,N_3863,N_3813);
nor U4392 (N_4392,N_3634,N_3333);
nand U4393 (N_4393,N_3808,N_3475);
nand U4394 (N_4394,N_3304,N_3232);
and U4395 (N_4395,N_3236,N_3891);
nand U4396 (N_4396,N_3893,N_3347);
nand U4397 (N_4397,N_3494,N_3945);
or U4398 (N_4398,N_3183,N_3438);
nor U4399 (N_4399,N_3997,N_3789);
and U4400 (N_4400,N_3545,N_3777);
xor U4401 (N_4401,N_3439,N_3497);
xor U4402 (N_4402,N_3164,N_3238);
nor U4403 (N_4403,N_3295,N_3466);
nor U4404 (N_4404,N_3531,N_3041);
nor U4405 (N_4405,N_3498,N_3750);
and U4406 (N_4406,N_3821,N_3955);
nor U4407 (N_4407,N_3203,N_3338);
or U4408 (N_4408,N_3489,N_3624);
and U4409 (N_4409,N_3486,N_3104);
or U4410 (N_4410,N_3191,N_3287);
and U4411 (N_4411,N_3947,N_3491);
xor U4412 (N_4412,N_3752,N_3996);
nor U4413 (N_4413,N_3118,N_3847);
xor U4414 (N_4414,N_3200,N_3172);
and U4415 (N_4415,N_3635,N_3810);
nor U4416 (N_4416,N_3672,N_3993);
nor U4417 (N_4417,N_3530,N_3730);
and U4418 (N_4418,N_3340,N_3182);
xor U4419 (N_4419,N_3448,N_3223);
or U4420 (N_4420,N_3376,N_3202);
nand U4421 (N_4421,N_3682,N_3717);
nand U4422 (N_4422,N_3029,N_3278);
or U4423 (N_4423,N_3073,N_3726);
nand U4424 (N_4424,N_3876,N_3386);
xnor U4425 (N_4425,N_3529,N_3618);
or U4426 (N_4426,N_3725,N_3302);
nor U4427 (N_4427,N_3417,N_3449);
and U4428 (N_4428,N_3446,N_3732);
and U4429 (N_4429,N_3954,N_3865);
xor U4430 (N_4430,N_3703,N_3581);
nand U4431 (N_4431,N_3094,N_3500);
nand U4432 (N_4432,N_3425,N_3722);
nor U4433 (N_4433,N_3357,N_3801);
nor U4434 (N_4434,N_3560,N_3952);
and U4435 (N_4435,N_3767,N_3364);
and U4436 (N_4436,N_3862,N_3818);
or U4437 (N_4437,N_3820,N_3307);
nand U4438 (N_4438,N_3664,N_3057);
xnor U4439 (N_4439,N_3507,N_3924);
or U4440 (N_4440,N_3054,N_3654);
or U4441 (N_4441,N_3389,N_3631);
xnor U4442 (N_4442,N_3881,N_3469);
nor U4443 (N_4443,N_3092,N_3470);
or U4444 (N_4444,N_3758,N_3643);
nor U4445 (N_4445,N_3697,N_3359);
nor U4446 (N_4446,N_3735,N_3396);
or U4447 (N_4447,N_3817,N_3502);
or U4448 (N_4448,N_3017,N_3226);
nor U4449 (N_4449,N_3080,N_3136);
and U4450 (N_4450,N_3650,N_3572);
and U4451 (N_4451,N_3025,N_3846);
nor U4452 (N_4452,N_3009,N_3661);
nand U4453 (N_4453,N_3920,N_3613);
nand U4454 (N_4454,N_3419,N_3258);
nand U4455 (N_4455,N_3107,N_3745);
and U4456 (N_4456,N_3851,N_3346);
xor U4457 (N_4457,N_3459,N_3580);
nor U4458 (N_4458,N_3139,N_3237);
nor U4459 (N_4459,N_3956,N_3373);
and U4460 (N_4460,N_3328,N_3586);
or U4461 (N_4461,N_3268,N_3915);
nor U4462 (N_4462,N_3070,N_3045);
nor U4463 (N_4463,N_3849,N_3269);
and U4464 (N_4464,N_3166,N_3429);
and U4465 (N_4465,N_3342,N_3105);
and U4466 (N_4466,N_3197,N_3751);
and U4467 (N_4467,N_3075,N_3445);
and U4468 (N_4468,N_3685,N_3383);
and U4469 (N_4469,N_3837,N_3521);
and U4470 (N_4470,N_3460,N_3422);
xnor U4471 (N_4471,N_3420,N_3289);
and U4472 (N_4472,N_3186,N_3032);
nor U4473 (N_4473,N_3695,N_3508);
and U4474 (N_4474,N_3867,N_3154);
or U4475 (N_4475,N_3652,N_3514);
nor U4476 (N_4476,N_3830,N_3378);
or U4477 (N_4477,N_3870,N_3206);
or U4478 (N_4478,N_3242,N_3966);
and U4479 (N_4479,N_3033,N_3720);
nand U4480 (N_4480,N_3544,N_3331);
nand U4481 (N_4481,N_3850,N_3125);
nand U4482 (N_4482,N_3596,N_3113);
and U4483 (N_4483,N_3822,N_3939);
or U4484 (N_4484,N_3515,N_3625);
nand U4485 (N_4485,N_3570,N_3562);
nand U4486 (N_4486,N_3819,N_3582);
and U4487 (N_4487,N_3754,N_3254);
xnor U4488 (N_4488,N_3283,N_3987);
and U4489 (N_4489,N_3921,N_3084);
xnor U4490 (N_4490,N_3540,N_3942);
nand U4491 (N_4491,N_3600,N_3085);
nand U4492 (N_4492,N_3790,N_3411);
or U4493 (N_4493,N_3368,N_3578);
xor U4494 (N_4494,N_3991,N_3612);
nor U4495 (N_4495,N_3548,N_3296);
nor U4496 (N_4496,N_3812,N_3310);
xor U4497 (N_4497,N_3282,N_3298);
and U4498 (N_4498,N_3285,N_3558);
nor U4499 (N_4499,N_3709,N_3574);
and U4500 (N_4500,N_3250,N_3443);
nor U4501 (N_4501,N_3182,N_3796);
xor U4502 (N_4502,N_3684,N_3167);
and U4503 (N_4503,N_3280,N_3577);
nor U4504 (N_4504,N_3401,N_3445);
and U4505 (N_4505,N_3201,N_3453);
or U4506 (N_4506,N_3892,N_3543);
nand U4507 (N_4507,N_3116,N_3586);
nor U4508 (N_4508,N_3862,N_3078);
or U4509 (N_4509,N_3773,N_3937);
nor U4510 (N_4510,N_3754,N_3565);
or U4511 (N_4511,N_3689,N_3655);
nand U4512 (N_4512,N_3396,N_3495);
xor U4513 (N_4513,N_3586,N_3365);
nor U4514 (N_4514,N_3724,N_3723);
and U4515 (N_4515,N_3958,N_3863);
nor U4516 (N_4516,N_3102,N_3006);
nand U4517 (N_4517,N_3532,N_3045);
and U4518 (N_4518,N_3215,N_3752);
nor U4519 (N_4519,N_3105,N_3834);
and U4520 (N_4520,N_3845,N_3617);
nand U4521 (N_4521,N_3122,N_3564);
nor U4522 (N_4522,N_3992,N_3668);
xnor U4523 (N_4523,N_3807,N_3762);
xnor U4524 (N_4524,N_3979,N_3418);
and U4525 (N_4525,N_3135,N_3889);
nor U4526 (N_4526,N_3863,N_3920);
nand U4527 (N_4527,N_3015,N_3552);
nor U4528 (N_4528,N_3999,N_3507);
nor U4529 (N_4529,N_3928,N_3033);
and U4530 (N_4530,N_3777,N_3005);
nor U4531 (N_4531,N_3354,N_3726);
xor U4532 (N_4532,N_3566,N_3712);
nor U4533 (N_4533,N_3350,N_3904);
nand U4534 (N_4534,N_3097,N_3620);
nand U4535 (N_4535,N_3671,N_3338);
nor U4536 (N_4536,N_3202,N_3785);
and U4537 (N_4537,N_3300,N_3398);
nand U4538 (N_4538,N_3480,N_3537);
or U4539 (N_4539,N_3744,N_3378);
nor U4540 (N_4540,N_3451,N_3625);
and U4541 (N_4541,N_3266,N_3437);
nor U4542 (N_4542,N_3059,N_3034);
nor U4543 (N_4543,N_3458,N_3464);
or U4544 (N_4544,N_3689,N_3014);
and U4545 (N_4545,N_3101,N_3014);
or U4546 (N_4546,N_3932,N_3354);
xor U4547 (N_4547,N_3729,N_3523);
nand U4548 (N_4548,N_3499,N_3705);
nand U4549 (N_4549,N_3900,N_3453);
nor U4550 (N_4550,N_3829,N_3012);
and U4551 (N_4551,N_3215,N_3040);
xnor U4552 (N_4552,N_3128,N_3546);
or U4553 (N_4553,N_3746,N_3660);
or U4554 (N_4554,N_3196,N_3652);
xor U4555 (N_4555,N_3078,N_3587);
nand U4556 (N_4556,N_3246,N_3123);
nand U4557 (N_4557,N_3123,N_3684);
or U4558 (N_4558,N_3620,N_3984);
and U4559 (N_4559,N_3096,N_3855);
or U4560 (N_4560,N_3555,N_3575);
xor U4561 (N_4561,N_3475,N_3238);
nor U4562 (N_4562,N_3330,N_3647);
nand U4563 (N_4563,N_3035,N_3356);
nand U4564 (N_4564,N_3791,N_3329);
nand U4565 (N_4565,N_3802,N_3625);
or U4566 (N_4566,N_3662,N_3666);
and U4567 (N_4567,N_3115,N_3529);
or U4568 (N_4568,N_3499,N_3254);
and U4569 (N_4569,N_3089,N_3945);
nor U4570 (N_4570,N_3379,N_3822);
nand U4571 (N_4571,N_3302,N_3543);
or U4572 (N_4572,N_3042,N_3238);
nor U4573 (N_4573,N_3978,N_3673);
and U4574 (N_4574,N_3832,N_3147);
nor U4575 (N_4575,N_3649,N_3481);
nor U4576 (N_4576,N_3227,N_3572);
nor U4577 (N_4577,N_3051,N_3578);
or U4578 (N_4578,N_3964,N_3359);
nor U4579 (N_4579,N_3660,N_3404);
nor U4580 (N_4580,N_3348,N_3110);
xnor U4581 (N_4581,N_3299,N_3736);
nand U4582 (N_4582,N_3119,N_3219);
nor U4583 (N_4583,N_3652,N_3148);
nor U4584 (N_4584,N_3286,N_3457);
or U4585 (N_4585,N_3265,N_3324);
or U4586 (N_4586,N_3492,N_3927);
nand U4587 (N_4587,N_3984,N_3219);
or U4588 (N_4588,N_3521,N_3166);
or U4589 (N_4589,N_3926,N_3455);
nand U4590 (N_4590,N_3801,N_3113);
and U4591 (N_4591,N_3107,N_3683);
nor U4592 (N_4592,N_3947,N_3473);
nand U4593 (N_4593,N_3194,N_3634);
and U4594 (N_4594,N_3878,N_3092);
nor U4595 (N_4595,N_3960,N_3060);
and U4596 (N_4596,N_3902,N_3809);
or U4597 (N_4597,N_3847,N_3006);
nand U4598 (N_4598,N_3010,N_3056);
xor U4599 (N_4599,N_3263,N_3330);
and U4600 (N_4600,N_3788,N_3747);
xnor U4601 (N_4601,N_3114,N_3489);
nor U4602 (N_4602,N_3395,N_3142);
and U4603 (N_4603,N_3759,N_3776);
or U4604 (N_4604,N_3890,N_3981);
and U4605 (N_4605,N_3010,N_3090);
and U4606 (N_4606,N_3098,N_3185);
and U4607 (N_4607,N_3337,N_3369);
and U4608 (N_4608,N_3394,N_3204);
or U4609 (N_4609,N_3143,N_3842);
xnor U4610 (N_4610,N_3847,N_3453);
nor U4611 (N_4611,N_3220,N_3518);
or U4612 (N_4612,N_3285,N_3390);
nor U4613 (N_4613,N_3380,N_3942);
nand U4614 (N_4614,N_3360,N_3763);
nand U4615 (N_4615,N_3019,N_3916);
nor U4616 (N_4616,N_3983,N_3447);
and U4617 (N_4617,N_3638,N_3559);
xor U4618 (N_4618,N_3532,N_3962);
nor U4619 (N_4619,N_3040,N_3893);
nand U4620 (N_4620,N_3604,N_3732);
and U4621 (N_4621,N_3446,N_3815);
and U4622 (N_4622,N_3914,N_3394);
nor U4623 (N_4623,N_3513,N_3961);
and U4624 (N_4624,N_3195,N_3816);
nand U4625 (N_4625,N_3334,N_3130);
nor U4626 (N_4626,N_3752,N_3056);
nand U4627 (N_4627,N_3006,N_3234);
or U4628 (N_4628,N_3546,N_3437);
nand U4629 (N_4629,N_3000,N_3727);
nor U4630 (N_4630,N_3478,N_3594);
and U4631 (N_4631,N_3317,N_3778);
nor U4632 (N_4632,N_3380,N_3811);
nor U4633 (N_4633,N_3252,N_3211);
nor U4634 (N_4634,N_3213,N_3791);
nand U4635 (N_4635,N_3656,N_3464);
nand U4636 (N_4636,N_3984,N_3122);
or U4637 (N_4637,N_3887,N_3413);
xnor U4638 (N_4638,N_3956,N_3154);
and U4639 (N_4639,N_3421,N_3176);
or U4640 (N_4640,N_3661,N_3712);
nand U4641 (N_4641,N_3471,N_3246);
xnor U4642 (N_4642,N_3582,N_3866);
and U4643 (N_4643,N_3883,N_3537);
and U4644 (N_4644,N_3133,N_3213);
xnor U4645 (N_4645,N_3299,N_3494);
or U4646 (N_4646,N_3582,N_3825);
nor U4647 (N_4647,N_3698,N_3175);
or U4648 (N_4648,N_3697,N_3194);
or U4649 (N_4649,N_3213,N_3307);
nand U4650 (N_4650,N_3373,N_3393);
or U4651 (N_4651,N_3285,N_3875);
nor U4652 (N_4652,N_3339,N_3978);
and U4653 (N_4653,N_3136,N_3460);
nand U4654 (N_4654,N_3948,N_3710);
xnor U4655 (N_4655,N_3780,N_3828);
nand U4656 (N_4656,N_3739,N_3927);
and U4657 (N_4657,N_3380,N_3794);
and U4658 (N_4658,N_3029,N_3059);
and U4659 (N_4659,N_3955,N_3994);
nor U4660 (N_4660,N_3192,N_3807);
nor U4661 (N_4661,N_3045,N_3168);
and U4662 (N_4662,N_3421,N_3606);
nor U4663 (N_4663,N_3910,N_3893);
xnor U4664 (N_4664,N_3823,N_3232);
xnor U4665 (N_4665,N_3925,N_3124);
or U4666 (N_4666,N_3214,N_3172);
nand U4667 (N_4667,N_3936,N_3592);
or U4668 (N_4668,N_3546,N_3117);
or U4669 (N_4669,N_3204,N_3854);
or U4670 (N_4670,N_3619,N_3114);
xnor U4671 (N_4671,N_3679,N_3906);
or U4672 (N_4672,N_3330,N_3309);
nand U4673 (N_4673,N_3902,N_3318);
nand U4674 (N_4674,N_3642,N_3545);
nor U4675 (N_4675,N_3285,N_3045);
xnor U4676 (N_4676,N_3275,N_3664);
or U4677 (N_4677,N_3586,N_3396);
nand U4678 (N_4678,N_3214,N_3726);
or U4679 (N_4679,N_3132,N_3337);
and U4680 (N_4680,N_3917,N_3408);
and U4681 (N_4681,N_3310,N_3999);
nand U4682 (N_4682,N_3429,N_3712);
and U4683 (N_4683,N_3732,N_3619);
and U4684 (N_4684,N_3290,N_3853);
xnor U4685 (N_4685,N_3660,N_3834);
and U4686 (N_4686,N_3826,N_3635);
and U4687 (N_4687,N_3233,N_3283);
or U4688 (N_4688,N_3688,N_3678);
or U4689 (N_4689,N_3637,N_3965);
nor U4690 (N_4690,N_3591,N_3053);
nor U4691 (N_4691,N_3142,N_3803);
nand U4692 (N_4692,N_3389,N_3509);
and U4693 (N_4693,N_3095,N_3098);
nand U4694 (N_4694,N_3888,N_3385);
nand U4695 (N_4695,N_3035,N_3794);
nand U4696 (N_4696,N_3006,N_3422);
and U4697 (N_4697,N_3715,N_3686);
nor U4698 (N_4698,N_3227,N_3272);
or U4699 (N_4699,N_3814,N_3171);
or U4700 (N_4700,N_3384,N_3083);
nand U4701 (N_4701,N_3496,N_3389);
nand U4702 (N_4702,N_3822,N_3812);
nand U4703 (N_4703,N_3085,N_3920);
nand U4704 (N_4704,N_3099,N_3123);
nor U4705 (N_4705,N_3016,N_3536);
nor U4706 (N_4706,N_3328,N_3345);
nor U4707 (N_4707,N_3361,N_3288);
xnor U4708 (N_4708,N_3821,N_3271);
or U4709 (N_4709,N_3638,N_3146);
or U4710 (N_4710,N_3423,N_3409);
nand U4711 (N_4711,N_3577,N_3734);
nor U4712 (N_4712,N_3094,N_3012);
nor U4713 (N_4713,N_3454,N_3511);
nor U4714 (N_4714,N_3315,N_3370);
nand U4715 (N_4715,N_3566,N_3149);
nand U4716 (N_4716,N_3043,N_3111);
nor U4717 (N_4717,N_3249,N_3204);
nor U4718 (N_4718,N_3553,N_3214);
nor U4719 (N_4719,N_3357,N_3656);
nand U4720 (N_4720,N_3661,N_3517);
and U4721 (N_4721,N_3842,N_3712);
and U4722 (N_4722,N_3534,N_3502);
and U4723 (N_4723,N_3297,N_3173);
and U4724 (N_4724,N_3516,N_3752);
or U4725 (N_4725,N_3019,N_3889);
xor U4726 (N_4726,N_3113,N_3703);
nand U4727 (N_4727,N_3082,N_3505);
nand U4728 (N_4728,N_3203,N_3729);
nor U4729 (N_4729,N_3673,N_3498);
and U4730 (N_4730,N_3073,N_3233);
and U4731 (N_4731,N_3550,N_3151);
or U4732 (N_4732,N_3088,N_3400);
and U4733 (N_4733,N_3676,N_3423);
and U4734 (N_4734,N_3318,N_3035);
and U4735 (N_4735,N_3497,N_3737);
and U4736 (N_4736,N_3452,N_3331);
and U4737 (N_4737,N_3004,N_3994);
or U4738 (N_4738,N_3014,N_3124);
xnor U4739 (N_4739,N_3481,N_3098);
xor U4740 (N_4740,N_3463,N_3192);
nor U4741 (N_4741,N_3952,N_3138);
or U4742 (N_4742,N_3717,N_3246);
and U4743 (N_4743,N_3593,N_3559);
nor U4744 (N_4744,N_3413,N_3801);
nand U4745 (N_4745,N_3942,N_3162);
and U4746 (N_4746,N_3851,N_3341);
or U4747 (N_4747,N_3820,N_3537);
nand U4748 (N_4748,N_3733,N_3091);
nand U4749 (N_4749,N_3263,N_3690);
nand U4750 (N_4750,N_3314,N_3378);
nand U4751 (N_4751,N_3479,N_3870);
nand U4752 (N_4752,N_3467,N_3899);
nor U4753 (N_4753,N_3790,N_3289);
nand U4754 (N_4754,N_3235,N_3872);
nand U4755 (N_4755,N_3953,N_3943);
nor U4756 (N_4756,N_3228,N_3841);
xor U4757 (N_4757,N_3029,N_3277);
nor U4758 (N_4758,N_3237,N_3792);
xnor U4759 (N_4759,N_3893,N_3532);
nor U4760 (N_4760,N_3732,N_3182);
and U4761 (N_4761,N_3199,N_3234);
nand U4762 (N_4762,N_3766,N_3624);
and U4763 (N_4763,N_3341,N_3641);
or U4764 (N_4764,N_3587,N_3098);
nor U4765 (N_4765,N_3988,N_3828);
and U4766 (N_4766,N_3278,N_3170);
xnor U4767 (N_4767,N_3338,N_3091);
and U4768 (N_4768,N_3529,N_3023);
nor U4769 (N_4769,N_3334,N_3330);
or U4770 (N_4770,N_3849,N_3759);
nand U4771 (N_4771,N_3105,N_3115);
or U4772 (N_4772,N_3428,N_3549);
and U4773 (N_4773,N_3361,N_3591);
nand U4774 (N_4774,N_3547,N_3906);
and U4775 (N_4775,N_3854,N_3572);
nand U4776 (N_4776,N_3489,N_3835);
or U4777 (N_4777,N_3191,N_3446);
nor U4778 (N_4778,N_3977,N_3703);
nor U4779 (N_4779,N_3494,N_3548);
nand U4780 (N_4780,N_3815,N_3417);
nand U4781 (N_4781,N_3201,N_3826);
nor U4782 (N_4782,N_3583,N_3404);
xnor U4783 (N_4783,N_3950,N_3492);
and U4784 (N_4784,N_3827,N_3808);
or U4785 (N_4785,N_3618,N_3003);
and U4786 (N_4786,N_3019,N_3458);
and U4787 (N_4787,N_3838,N_3435);
nor U4788 (N_4788,N_3998,N_3586);
and U4789 (N_4789,N_3812,N_3738);
nand U4790 (N_4790,N_3634,N_3760);
or U4791 (N_4791,N_3785,N_3982);
nand U4792 (N_4792,N_3989,N_3038);
nor U4793 (N_4793,N_3097,N_3564);
or U4794 (N_4794,N_3273,N_3813);
or U4795 (N_4795,N_3729,N_3600);
or U4796 (N_4796,N_3387,N_3973);
and U4797 (N_4797,N_3106,N_3766);
nand U4798 (N_4798,N_3506,N_3135);
nor U4799 (N_4799,N_3852,N_3615);
and U4800 (N_4800,N_3268,N_3787);
nor U4801 (N_4801,N_3074,N_3547);
and U4802 (N_4802,N_3430,N_3200);
nor U4803 (N_4803,N_3743,N_3658);
and U4804 (N_4804,N_3400,N_3580);
nand U4805 (N_4805,N_3151,N_3559);
or U4806 (N_4806,N_3312,N_3917);
or U4807 (N_4807,N_3792,N_3881);
nand U4808 (N_4808,N_3627,N_3817);
and U4809 (N_4809,N_3985,N_3009);
and U4810 (N_4810,N_3499,N_3729);
nor U4811 (N_4811,N_3912,N_3007);
nor U4812 (N_4812,N_3987,N_3319);
and U4813 (N_4813,N_3301,N_3045);
nor U4814 (N_4814,N_3485,N_3849);
nor U4815 (N_4815,N_3443,N_3357);
nor U4816 (N_4816,N_3964,N_3227);
or U4817 (N_4817,N_3150,N_3000);
nand U4818 (N_4818,N_3441,N_3808);
and U4819 (N_4819,N_3751,N_3256);
nand U4820 (N_4820,N_3369,N_3335);
and U4821 (N_4821,N_3749,N_3945);
xor U4822 (N_4822,N_3581,N_3724);
or U4823 (N_4823,N_3818,N_3949);
and U4824 (N_4824,N_3116,N_3133);
nor U4825 (N_4825,N_3961,N_3045);
nand U4826 (N_4826,N_3347,N_3503);
nor U4827 (N_4827,N_3276,N_3010);
nor U4828 (N_4828,N_3384,N_3397);
and U4829 (N_4829,N_3187,N_3496);
nor U4830 (N_4830,N_3104,N_3174);
xnor U4831 (N_4831,N_3491,N_3347);
and U4832 (N_4832,N_3568,N_3173);
nand U4833 (N_4833,N_3416,N_3037);
xor U4834 (N_4834,N_3448,N_3227);
or U4835 (N_4835,N_3837,N_3465);
nor U4836 (N_4836,N_3994,N_3708);
nor U4837 (N_4837,N_3108,N_3183);
and U4838 (N_4838,N_3146,N_3204);
or U4839 (N_4839,N_3228,N_3550);
or U4840 (N_4840,N_3308,N_3475);
and U4841 (N_4841,N_3559,N_3152);
and U4842 (N_4842,N_3083,N_3612);
and U4843 (N_4843,N_3710,N_3064);
nand U4844 (N_4844,N_3371,N_3209);
and U4845 (N_4845,N_3211,N_3530);
xnor U4846 (N_4846,N_3986,N_3945);
or U4847 (N_4847,N_3163,N_3808);
nor U4848 (N_4848,N_3395,N_3232);
nor U4849 (N_4849,N_3264,N_3643);
and U4850 (N_4850,N_3478,N_3296);
xor U4851 (N_4851,N_3460,N_3990);
or U4852 (N_4852,N_3285,N_3406);
nor U4853 (N_4853,N_3795,N_3203);
nor U4854 (N_4854,N_3280,N_3664);
or U4855 (N_4855,N_3759,N_3930);
and U4856 (N_4856,N_3617,N_3172);
nand U4857 (N_4857,N_3385,N_3144);
xnor U4858 (N_4858,N_3696,N_3074);
xnor U4859 (N_4859,N_3633,N_3021);
or U4860 (N_4860,N_3565,N_3344);
or U4861 (N_4861,N_3812,N_3506);
nand U4862 (N_4862,N_3277,N_3229);
and U4863 (N_4863,N_3463,N_3356);
and U4864 (N_4864,N_3710,N_3034);
nand U4865 (N_4865,N_3262,N_3215);
and U4866 (N_4866,N_3584,N_3229);
nor U4867 (N_4867,N_3888,N_3136);
nor U4868 (N_4868,N_3198,N_3239);
or U4869 (N_4869,N_3753,N_3747);
or U4870 (N_4870,N_3616,N_3103);
and U4871 (N_4871,N_3503,N_3751);
nor U4872 (N_4872,N_3251,N_3497);
nor U4873 (N_4873,N_3307,N_3344);
nor U4874 (N_4874,N_3074,N_3478);
and U4875 (N_4875,N_3403,N_3949);
or U4876 (N_4876,N_3341,N_3252);
nand U4877 (N_4877,N_3058,N_3183);
or U4878 (N_4878,N_3182,N_3192);
or U4879 (N_4879,N_3116,N_3872);
or U4880 (N_4880,N_3168,N_3200);
or U4881 (N_4881,N_3550,N_3359);
and U4882 (N_4882,N_3925,N_3177);
xnor U4883 (N_4883,N_3562,N_3805);
nand U4884 (N_4884,N_3110,N_3852);
nand U4885 (N_4885,N_3537,N_3629);
or U4886 (N_4886,N_3353,N_3995);
xnor U4887 (N_4887,N_3038,N_3325);
and U4888 (N_4888,N_3771,N_3769);
nor U4889 (N_4889,N_3493,N_3686);
or U4890 (N_4890,N_3424,N_3207);
nand U4891 (N_4891,N_3470,N_3199);
and U4892 (N_4892,N_3054,N_3906);
nand U4893 (N_4893,N_3057,N_3767);
nand U4894 (N_4894,N_3855,N_3074);
nor U4895 (N_4895,N_3814,N_3573);
nor U4896 (N_4896,N_3399,N_3573);
or U4897 (N_4897,N_3698,N_3743);
and U4898 (N_4898,N_3375,N_3223);
or U4899 (N_4899,N_3751,N_3157);
xor U4900 (N_4900,N_3006,N_3204);
nand U4901 (N_4901,N_3415,N_3143);
xor U4902 (N_4902,N_3011,N_3760);
nand U4903 (N_4903,N_3807,N_3439);
and U4904 (N_4904,N_3524,N_3998);
nor U4905 (N_4905,N_3902,N_3805);
nand U4906 (N_4906,N_3905,N_3423);
nand U4907 (N_4907,N_3686,N_3805);
xnor U4908 (N_4908,N_3901,N_3326);
nor U4909 (N_4909,N_3555,N_3901);
and U4910 (N_4910,N_3497,N_3030);
nor U4911 (N_4911,N_3542,N_3065);
nor U4912 (N_4912,N_3706,N_3741);
nor U4913 (N_4913,N_3370,N_3731);
xor U4914 (N_4914,N_3690,N_3062);
nor U4915 (N_4915,N_3400,N_3154);
xnor U4916 (N_4916,N_3322,N_3837);
or U4917 (N_4917,N_3112,N_3386);
nand U4918 (N_4918,N_3038,N_3950);
nand U4919 (N_4919,N_3960,N_3578);
and U4920 (N_4920,N_3225,N_3289);
and U4921 (N_4921,N_3724,N_3008);
xor U4922 (N_4922,N_3072,N_3146);
xor U4923 (N_4923,N_3764,N_3480);
nor U4924 (N_4924,N_3847,N_3234);
and U4925 (N_4925,N_3117,N_3187);
nand U4926 (N_4926,N_3255,N_3286);
nor U4927 (N_4927,N_3964,N_3090);
xor U4928 (N_4928,N_3030,N_3366);
xnor U4929 (N_4929,N_3087,N_3986);
or U4930 (N_4930,N_3989,N_3741);
nor U4931 (N_4931,N_3656,N_3109);
or U4932 (N_4932,N_3932,N_3298);
xnor U4933 (N_4933,N_3265,N_3883);
nand U4934 (N_4934,N_3472,N_3898);
nor U4935 (N_4935,N_3580,N_3242);
or U4936 (N_4936,N_3862,N_3071);
nand U4937 (N_4937,N_3962,N_3952);
nand U4938 (N_4938,N_3371,N_3983);
or U4939 (N_4939,N_3459,N_3738);
nor U4940 (N_4940,N_3849,N_3974);
or U4941 (N_4941,N_3823,N_3277);
or U4942 (N_4942,N_3041,N_3868);
nor U4943 (N_4943,N_3042,N_3998);
nor U4944 (N_4944,N_3741,N_3251);
and U4945 (N_4945,N_3412,N_3644);
and U4946 (N_4946,N_3726,N_3690);
nand U4947 (N_4947,N_3208,N_3036);
xor U4948 (N_4948,N_3155,N_3523);
nand U4949 (N_4949,N_3573,N_3023);
xnor U4950 (N_4950,N_3022,N_3308);
xor U4951 (N_4951,N_3047,N_3395);
nor U4952 (N_4952,N_3152,N_3037);
or U4953 (N_4953,N_3149,N_3593);
or U4954 (N_4954,N_3872,N_3688);
and U4955 (N_4955,N_3801,N_3457);
or U4956 (N_4956,N_3881,N_3744);
nor U4957 (N_4957,N_3113,N_3708);
xor U4958 (N_4958,N_3517,N_3665);
nand U4959 (N_4959,N_3686,N_3757);
xor U4960 (N_4960,N_3459,N_3632);
nor U4961 (N_4961,N_3503,N_3715);
or U4962 (N_4962,N_3830,N_3360);
or U4963 (N_4963,N_3919,N_3670);
or U4964 (N_4964,N_3450,N_3078);
nand U4965 (N_4965,N_3296,N_3416);
or U4966 (N_4966,N_3001,N_3213);
nor U4967 (N_4967,N_3128,N_3438);
and U4968 (N_4968,N_3347,N_3650);
nor U4969 (N_4969,N_3701,N_3236);
and U4970 (N_4970,N_3462,N_3658);
nand U4971 (N_4971,N_3015,N_3144);
or U4972 (N_4972,N_3242,N_3147);
nand U4973 (N_4973,N_3292,N_3244);
or U4974 (N_4974,N_3047,N_3934);
or U4975 (N_4975,N_3407,N_3526);
nor U4976 (N_4976,N_3144,N_3487);
and U4977 (N_4977,N_3849,N_3040);
or U4978 (N_4978,N_3861,N_3427);
nor U4979 (N_4979,N_3721,N_3733);
nor U4980 (N_4980,N_3808,N_3343);
or U4981 (N_4981,N_3353,N_3997);
nor U4982 (N_4982,N_3397,N_3599);
and U4983 (N_4983,N_3012,N_3648);
and U4984 (N_4984,N_3269,N_3069);
and U4985 (N_4985,N_3463,N_3518);
and U4986 (N_4986,N_3736,N_3417);
and U4987 (N_4987,N_3108,N_3444);
and U4988 (N_4988,N_3673,N_3052);
or U4989 (N_4989,N_3074,N_3027);
and U4990 (N_4990,N_3499,N_3534);
xor U4991 (N_4991,N_3581,N_3134);
nand U4992 (N_4992,N_3210,N_3755);
xor U4993 (N_4993,N_3896,N_3492);
or U4994 (N_4994,N_3012,N_3436);
nand U4995 (N_4995,N_3119,N_3089);
nand U4996 (N_4996,N_3503,N_3611);
and U4997 (N_4997,N_3990,N_3229);
nand U4998 (N_4998,N_3094,N_3616);
or U4999 (N_4999,N_3653,N_3401);
or U5000 (N_5000,N_4195,N_4181);
and U5001 (N_5001,N_4267,N_4005);
nor U5002 (N_5002,N_4228,N_4535);
nand U5003 (N_5003,N_4752,N_4276);
nor U5004 (N_5004,N_4473,N_4901);
nand U5005 (N_5005,N_4614,N_4140);
or U5006 (N_5006,N_4282,N_4873);
nand U5007 (N_5007,N_4877,N_4676);
nand U5008 (N_5008,N_4116,N_4413);
or U5009 (N_5009,N_4899,N_4943);
nor U5010 (N_5010,N_4438,N_4170);
and U5011 (N_5011,N_4346,N_4744);
nand U5012 (N_5012,N_4792,N_4514);
xor U5013 (N_5013,N_4059,N_4644);
and U5014 (N_5014,N_4259,N_4906);
nor U5015 (N_5015,N_4671,N_4100);
or U5016 (N_5016,N_4757,N_4232);
nor U5017 (N_5017,N_4057,N_4331);
nor U5018 (N_5018,N_4117,N_4250);
nand U5019 (N_5019,N_4333,N_4600);
or U5020 (N_5020,N_4749,N_4482);
nand U5021 (N_5021,N_4640,N_4764);
and U5022 (N_5022,N_4270,N_4283);
and U5023 (N_5023,N_4420,N_4012);
nor U5024 (N_5024,N_4824,N_4762);
and U5025 (N_5025,N_4302,N_4495);
nand U5026 (N_5026,N_4870,N_4596);
nor U5027 (N_5027,N_4936,N_4225);
nand U5028 (N_5028,N_4506,N_4039);
nor U5029 (N_5029,N_4650,N_4108);
nor U5030 (N_5030,N_4446,N_4975);
or U5031 (N_5031,N_4791,N_4165);
and U5032 (N_5032,N_4982,N_4867);
nor U5033 (N_5033,N_4444,N_4390);
nor U5034 (N_5034,N_4103,N_4325);
nand U5035 (N_5035,N_4903,N_4106);
nand U5036 (N_5036,N_4552,N_4178);
nor U5037 (N_5037,N_4935,N_4942);
nor U5038 (N_5038,N_4743,N_4229);
nand U5039 (N_5039,N_4980,N_4998);
xor U5040 (N_5040,N_4448,N_4349);
nand U5041 (N_5041,N_4487,N_4431);
or U5042 (N_5042,N_4869,N_4911);
nand U5043 (N_5043,N_4782,N_4344);
nand U5044 (N_5044,N_4890,N_4766);
nand U5045 (N_5045,N_4385,N_4434);
nor U5046 (N_5046,N_4518,N_4281);
or U5047 (N_5047,N_4001,N_4714);
and U5048 (N_5048,N_4391,N_4995);
or U5049 (N_5049,N_4511,N_4131);
and U5050 (N_5050,N_4287,N_4688);
and U5051 (N_5051,N_4698,N_4311);
nand U5052 (N_5052,N_4529,N_4266);
or U5053 (N_5053,N_4043,N_4696);
xor U5054 (N_5054,N_4635,N_4082);
or U5055 (N_5055,N_4423,N_4254);
nand U5056 (N_5056,N_4990,N_4395);
and U5057 (N_5057,N_4636,N_4891);
nand U5058 (N_5058,N_4104,N_4148);
and U5059 (N_5059,N_4667,N_4685);
nor U5060 (N_5060,N_4860,N_4780);
nor U5061 (N_5061,N_4755,N_4433);
nand U5062 (N_5062,N_4244,N_4306);
nand U5063 (N_5063,N_4855,N_4846);
and U5064 (N_5064,N_4414,N_4121);
nor U5065 (N_5065,N_4162,N_4214);
or U5066 (N_5066,N_4775,N_4411);
and U5067 (N_5067,N_4294,N_4656);
xnor U5068 (N_5068,N_4280,N_4701);
nor U5069 (N_5069,N_4258,N_4295);
and U5070 (N_5070,N_4209,N_4004);
and U5071 (N_5071,N_4392,N_4985);
and U5072 (N_5072,N_4566,N_4272);
or U5073 (N_5073,N_4692,N_4951);
nor U5074 (N_5074,N_4927,N_4018);
or U5075 (N_5075,N_4763,N_4958);
and U5076 (N_5076,N_4526,N_4620);
nand U5077 (N_5077,N_4547,N_4924);
or U5078 (N_5078,N_4954,N_4442);
and U5079 (N_5079,N_4727,N_4885);
nand U5080 (N_5080,N_4095,N_4425);
and U5081 (N_5081,N_4492,N_4088);
and U5082 (N_5082,N_4008,N_4955);
xnor U5083 (N_5083,N_4109,N_4594);
nor U5084 (N_5084,N_4872,N_4080);
and U5085 (N_5085,N_4686,N_4101);
or U5086 (N_5086,N_4388,N_4613);
nand U5087 (N_5087,N_4092,N_4716);
nand U5088 (N_5088,N_4062,N_4205);
nand U5089 (N_5089,N_4753,N_4125);
xnor U5090 (N_5090,N_4319,N_4499);
nor U5091 (N_5091,N_4628,N_4601);
or U5092 (N_5092,N_4257,N_4748);
nand U5093 (N_5093,N_4187,N_4112);
xnor U5094 (N_5094,N_4723,N_4718);
nor U5095 (N_5095,N_4141,N_4300);
nor U5096 (N_5096,N_4687,N_4216);
nor U5097 (N_5097,N_4668,N_4907);
and U5098 (N_5098,N_4163,N_4624);
or U5099 (N_5099,N_4631,N_4772);
or U5100 (N_5100,N_4738,N_4470);
nor U5101 (N_5101,N_4750,N_4188);
nand U5102 (N_5102,N_4622,N_4050);
nand U5103 (N_5103,N_4273,N_4003);
and U5104 (N_5104,N_4618,N_4263);
or U5105 (N_5105,N_4831,N_4251);
or U5106 (N_5106,N_4290,N_4794);
nor U5107 (N_5107,N_4567,N_4900);
or U5108 (N_5108,N_4673,N_4669);
xor U5109 (N_5109,N_4948,N_4969);
nand U5110 (N_5110,N_4445,N_4450);
xnor U5111 (N_5111,N_4505,N_4934);
nor U5112 (N_5112,N_4172,N_4652);
and U5113 (N_5113,N_4069,N_4467);
and U5114 (N_5114,N_4953,N_4834);
nor U5115 (N_5115,N_4706,N_4666);
xor U5116 (N_5116,N_4968,N_4611);
and U5117 (N_5117,N_4974,N_4055);
nor U5118 (N_5118,N_4902,N_4369);
nor U5119 (N_5119,N_4862,N_4503);
and U5120 (N_5120,N_4602,N_4771);
or U5121 (N_5121,N_4457,N_4852);
nand U5122 (N_5122,N_4805,N_4580);
and U5123 (N_5123,N_4387,N_4724);
nor U5124 (N_5124,N_4704,N_4127);
nand U5125 (N_5125,N_4115,N_4058);
and U5126 (N_5126,N_4049,N_4068);
nand U5127 (N_5127,N_4756,N_4139);
xnor U5128 (N_5128,N_4695,N_4374);
nand U5129 (N_5129,N_4219,N_4021);
and U5130 (N_5130,N_4277,N_4405);
nand U5131 (N_5131,N_4575,N_4983);
or U5132 (N_5132,N_4383,N_4019);
or U5133 (N_5133,N_4715,N_4284);
and U5134 (N_5134,N_4449,N_4785);
xor U5135 (N_5135,N_4167,N_4452);
nand U5136 (N_5136,N_4774,N_4017);
and U5137 (N_5137,N_4957,N_4584);
and U5138 (N_5138,N_4813,N_4340);
nor U5139 (N_5139,N_4986,N_4469);
and U5140 (N_5140,N_4120,N_4963);
nand U5141 (N_5141,N_4978,N_4320);
and U5142 (N_5142,N_4142,N_4326);
nand U5143 (N_5143,N_4626,N_4767);
and U5144 (N_5144,N_4956,N_4658);
nor U5145 (N_5145,N_4558,N_4910);
nor U5146 (N_5146,N_4398,N_4278);
xnor U5147 (N_5147,N_4321,N_4905);
nand U5148 (N_5148,N_4833,N_4897);
nor U5149 (N_5149,N_4048,N_4539);
xor U5150 (N_5150,N_4838,N_4328);
nand U5151 (N_5151,N_4670,N_4230);
or U5152 (N_5152,N_4150,N_4989);
nor U5153 (N_5153,N_4816,N_4481);
and U5154 (N_5154,N_4574,N_4587);
nand U5155 (N_5155,N_4593,N_4410);
or U5156 (N_5156,N_4304,N_4962);
and U5157 (N_5157,N_4072,N_4751);
nor U5158 (N_5158,N_4546,N_4617);
and U5159 (N_5159,N_4061,N_4923);
nor U5160 (N_5160,N_4474,N_4381);
xnor U5161 (N_5161,N_4002,N_4754);
nor U5162 (N_5162,N_4498,N_4261);
and U5163 (N_5163,N_4418,N_4376);
and U5164 (N_5164,N_4168,N_4478);
nor U5165 (N_5165,N_4486,N_4305);
nand U5166 (N_5166,N_4342,N_4238);
and U5167 (N_5167,N_4107,N_4880);
xor U5168 (N_5168,N_4534,N_4472);
nand U5169 (N_5169,N_4235,N_4682);
nand U5170 (N_5170,N_4513,N_4582);
nand U5171 (N_5171,N_4299,N_4159);
xnor U5172 (N_5172,N_4661,N_4459);
xnor U5173 (N_5173,N_4157,N_4347);
or U5174 (N_5174,N_4933,N_4076);
nand U5175 (N_5175,N_4521,N_4352);
or U5176 (N_5176,N_4770,N_4013);
nand U5177 (N_5177,N_4407,N_4997);
xor U5178 (N_5178,N_4553,N_4011);
nand U5179 (N_5179,N_4154,N_4536);
xnor U5180 (N_5180,N_4458,N_4932);
nand U5181 (N_5181,N_4071,N_4056);
or U5182 (N_5182,N_4060,N_4843);
and U5183 (N_5183,N_4703,N_4312);
or U5184 (N_5184,N_4204,N_4460);
nor U5185 (N_5185,N_4079,N_4882);
nand U5186 (N_5186,N_4881,N_4585);
and U5187 (N_5187,N_4190,N_4525);
nand U5188 (N_5188,N_4045,N_4175);
nand U5189 (N_5189,N_4412,N_4330);
nand U5190 (N_5190,N_4179,N_4726);
or U5191 (N_5191,N_4865,N_4086);
nor U5192 (N_5192,N_4914,N_4679);
nand U5193 (N_5193,N_4237,N_4675);
nand U5194 (N_5194,N_4711,N_4965);
and U5195 (N_5195,N_4221,N_4629);
or U5196 (N_5196,N_4074,N_4158);
nor U5197 (N_5197,N_4067,N_4586);
nor U5198 (N_5198,N_4416,N_4657);
xor U5199 (N_5199,N_4836,N_4211);
and U5200 (N_5200,N_4156,N_4694);
nand U5201 (N_5201,N_4776,N_4191);
or U5202 (N_5202,N_4806,N_4099);
nand U5203 (N_5203,N_4977,N_4083);
or U5204 (N_5204,N_4393,N_4879);
nor U5205 (N_5205,N_4515,N_4046);
nand U5206 (N_5206,N_4761,N_4377);
and U5207 (N_5207,N_4429,N_4875);
and U5208 (N_5208,N_4246,N_4610);
nand U5209 (N_5209,N_4397,N_4378);
nand U5210 (N_5210,N_4528,N_4297);
and U5211 (N_5211,N_4143,N_4360);
nand U5212 (N_5212,N_4262,N_4712);
nand U5213 (N_5213,N_4615,N_4196);
nand U5214 (N_5214,N_4928,N_4527);
or U5215 (N_5215,N_4683,N_4819);
and U5216 (N_5216,N_4700,N_4365);
nand U5217 (N_5217,N_4721,N_4144);
and U5218 (N_5218,N_4677,N_4085);
and U5219 (N_5219,N_4363,N_4884);
nor U5220 (N_5220,N_4020,N_4950);
or U5221 (N_5221,N_4130,N_4415);
nand U5222 (N_5222,N_4522,N_4781);
nor U5223 (N_5223,N_4691,N_4542);
nand U5224 (N_5224,N_4268,N_4041);
nand U5225 (N_5225,N_4409,N_4801);
and U5226 (N_5226,N_4063,N_4355);
xor U5227 (N_5227,N_4009,N_4680);
or U5228 (N_5228,N_4913,N_4912);
nand U5229 (N_5229,N_4798,N_4549);
and U5230 (N_5230,N_4742,N_4389);
and U5231 (N_5231,N_4840,N_4541);
nor U5232 (N_5232,N_4672,N_4337);
nand U5233 (N_5233,N_4252,N_4984);
and U5234 (N_5234,N_4078,N_4576);
xnor U5235 (N_5235,N_4314,N_4236);
nor U5236 (N_5236,N_4630,N_4098);
or U5237 (N_5237,N_4560,N_4126);
or U5238 (N_5238,N_4197,N_4634);
and U5239 (N_5239,N_4096,N_4128);
or U5240 (N_5240,N_4462,N_4973);
xor U5241 (N_5241,N_4255,N_4269);
or U5242 (N_5242,N_4184,N_4937);
nor U5243 (N_5243,N_4023,N_4684);
xor U5244 (N_5244,N_4571,N_4638);
nor U5245 (N_5245,N_4186,N_4802);
and U5246 (N_5246,N_4896,N_4339);
xor U5247 (N_5247,N_4815,N_4137);
nor U5248 (N_5248,N_4026,N_4359);
and U5249 (N_5249,N_4783,N_4737);
or U5250 (N_5250,N_4941,N_4508);
nand U5251 (N_5251,N_4435,N_4940);
nor U5252 (N_5252,N_4199,N_4662);
nand U5253 (N_5253,N_4437,N_4678);
nor U5254 (N_5254,N_4105,N_4345);
nor U5255 (N_5255,N_4952,N_4090);
and U5256 (N_5256,N_4837,N_4177);
or U5257 (N_5257,N_4133,N_4849);
xnor U5258 (N_5258,N_4510,N_4155);
and U5259 (N_5259,N_4579,N_4741);
xnor U5260 (N_5260,N_4648,N_4303);
xor U5261 (N_5261,N_4544,N_4562);
and U5262 (N_5262,N_4129,N_4296);
nor U5263 (N_5263,N_4256,N_4189);
nor U5264 (N_5264,N_4279,N_4520);
or U5265 (N_5265,N_4859,N_4489);
xor U5266 (N_5266,N_4599,N_4947);
and U5267 (N_5267,N_4336,N_4605);
or U5268 (N_5268,N_4681,N_4275);
nand U5269 (N_5269,N_4348,N_4226);
nor U5270 (N_5270,N_4193,N_4334);
or U5271 (N_5271,N_4739,N_4722);
nand U5272 (N_5272,N_4024,N_4145);
and U5273 (N_5273,N_4639,N_4967);
and U5274 (N_5274,N_4176,N_4709);
nor U5275 (N_5275,N_4335,N_4151);
and U5276 (N_5276,N_4945,N_4091);
and U5277 (N_5277,N_4301,N_4271);
xor U5278 (N_5278,N_4590,N_4164);
xnor U5279 (N_5279,N_4111,N_4641);
nand U5280 (N_5280,N_4298,N_4243);
xnor U5281 (N_5281,N_4814,N_4245);
nor U5282 (N_5282,N_4035,N_4915);
and U5283 (N_5283,N_4317,N_4033);
nor U5284 (N_5284,N_4689,N_4044);
nand U5285 (N_5285,N_4572,N_4364);
nand U5286 (N_5286,N_4358,N_4182);
xnor U5287 (N_5287,N_4608,N_4971);
nand U5288 (N_5288,N_4642,N_4516);
and U5289 (N_5289,N_4356,N_4779);
or U5290 (N_5290,N_4789,N_4198);
nand U5291 (N_5291,N_4519,N_4871);
and U5292 (N_5292,N_4408,N_4203);
xnor U5293 (N_5293,N_4493,N_4494);
or U5294 (N_5294,N_4240,N_4597);
nor U5295 (N_5295,N_4394,N_4166);
nor U5296 (N_5296,N_4491,N_4454);
nor U5297 (N_5297,N_4451,N_4939);
and U5298 (N_5298,N_4598,N_4417);
and U5299 (N_5299,N_4220,N_4561);
and U5300 (N_5300,N_4064,N_4274);
nand U5301 (N_5301,N_4066,N_4595);
nand U5302 (N_5302,N_4479,N_4160);
nand U5303 (N_5303,N_4892,N_4353);
or U5304 (N_5304,N_4288,N_4291);
or U5305 (N_5305,N_4808,N_4070);
nand U5306 (N_5306,N_4464,N_4351);
nand U5307 (N_5307,N_4665,N_4894);
or U5308 (N_5308,N_4745,N_4324);
nand U5309 (N_5309,N_4740,N_4909);
or U5310 (N_5310,N_4822,N_4570);
nor U5311 (N_5311,N_4223,N_4996);
xor U5312 (N_5312,N_4361,N_4428);
or U5313 (N_5313,N_4366,N_4404);
and U5314 (N_5314,N_4769,N_4465);
xor U5315 (N_5315,N_4800,N_4565);
and U5316 (N_5316,N_4874,N_4135);
xnor U5317 (N_5317,N_4842,N_4732);
nor U5318 (N_5318,N_4208,N_4619);
nand U5319 (N_5319,N_4367,N_4322);
nor U5320 (N_5320,N_4372,N_4403);
nor U5321 (N_5321,N_4264,N_4400);
nand U5322 (N_5322,N_4147,N_4114);
xnor U5323 (N_5323,N_4916,N_4646);
nor U5324 (N_5324,N_4093,N_4202);
and U5325 (N_5325,N_4592,N_4654);
or U5326 (N_5326,N_4134,N_4215);
nor U5327 (N_5327,N_4921,N_4530);
and U5328 (N_5328,N_4222,N_4876);
and U5329 (N_5329,N_4286,N_4746);
nand U5330 (N_5330,N_4375,N_4292);
or U5331 (N_5331,N_4893,N_4858);
nor U5332 (N_5332,N_4559,N_4632);
nor U5333 (N_5333,N_4674,N_4655);
or U5334 (N_5334,N_4702,N_4509);
or U5335 (N_5335,N_4864,N_4988);
nand U5336 (N_5336,N_4224,N_4563);
nand U5337 (N_5337,N_4710,N_4730);
nor U5338 (N_5338,N_4427,N_4382);
nand U5339 (N_5339,N_4790,N_4419);
xnor U5340 (N_5340,N_4550,N_4007);
nor U5341 (N_5341,N_4854,N_4153);
xor U5342 (N_5342,N_4373,N_4664);
and U5343 (N_5343,N_4315,N_4979);
nor U5344 (N_5344,N_4606,N_4239);
nor U5345 (N_5345,N_4758,N_4247);
and U5346 (N_5346,N_4917,N_4323);
and U5347 (N_5347,N_4327,N_4637);
and U5348 (N_5348,N_4828,N_4016);
or U5349 (N_5349,N_4734,N_4850);
nor U5350 (N_5350,N_4699,N_4354);
or U5351 (N_5351,N_4210,N_4659);
nor U5352 (N_5352,N_4384,N_4185);
nand U5353 (N_5353,N_4054,N_4468);
nand U5354 (N_5354,N_4543,N_4386);
or U5355 (N_5355,N_4826,N_4436);
or U5356 (N_5356,N_4000,N_4797);
nand U5357 (N_5357,N_4094,N_4138);
or U5358 (N_5358,N_4338,N_4643);
nand U5359 (N_5359,N_4500,N_4441);
nand U5360 (N_5360,N_4488,N_4625);
and U5361 (N_5361,N_4904,N_4633);
nand U5362 (N_5362,N_4787,N_4960);
or U5363 (N_5363,N_4777,N_4042);
nand U5364 (N_5364,N_4047,N_4231);
nand U5365 (N_5365,N_4930,N_4075);
nor U5366 (N_5366,N_4693,N_4192);
or U5367 (N_5367,N_4040,N_4490);
nand U5368 (N_5368,N_4118,N_4554);
or U5369 (N_5369,N_4249,N_4293);
or U5370 (N_5370,N_4310,N_4289);
or U5371 (N_5371,N_4329,N_4647);
nor U5372 (N_5372,N_4201,N_4728);
or U5373 (N_5373,N_4523,N_4030);
or U5374 (N_5374,N_4476,N_4213);
nand U5375 (N_5375,N_4820,N_4545);
nor U5376 (N_5376,N_4084,N_4512);
nand U5377 (N_5377,N_4132,N_4014);
or U5378 (N_5378,N_4052,N_4113);
nand U5379 (N_5379,N_4218,N_4747);
nor U5380 (N_5380,N_4583,N_4847);
and U5381 (N_5381,N_4406,N_4788);
nor U5382 (N_5382,N_4949,N_4961);
xnor U5383 (N_5383,N_4999,N_4217);
nand U5384 (N_5384,N_4690,N_4817);
nand U5385 (N_5385,N_4697,N_4540);
nand U5386 (N_5386,N_4430,N_4485);
nand U5387 (N_5387,N_4759,N_4357);
nor U5388 (N_5388,N_4573,N_4920);
nand U5389 (N_5389,N_4557,N_4038);
nor U5390 (N_5390,N_4316,N_4623);
or U5391 (N_5391,N_4649,N_4895);
nand U5392 (N_5392,N_4350,N_4604);
or U5393 (N_5393,N_4396,N_4736);
nor U5394 (N_5394,N_4480,N_4929);
and U5395 (N_5395,N_4857,N_4786);
nand U5396 (N_5396,N_4851,N_4966);
and U5397 (N_5397,N_4053,N_4853);
nand U5398 (N_5398,N_4110,N_4309);
or U5399 (N_5399,N_4760,N_4421);
nand U5400 (N_5400,N_4171,N_4032);
nor U5401 (N_5401,N_4705,N_4926);
and U5402 (N_5402,N_4371,N_4102);
nand U5403 (N_5403,N_4380,N_4821);
and U5404 (N_5404,N_4022,N_4343);
or U5405 (N_5405,N_4399,N_4856);
or U5406 (N_5406,N_4073,N_4987);
and U5407 (N_5407,N_4568,N_4253);
or U5408 (N_5408,N_4898,N_4015);
and U5409 (N_5409,N_4795,N_4830);
or U5410 (N_5410,N_4878,N_4006);
xnor U5411 (N_5411,N_4889,N_4194);
nor U5412 (N_5412,N_4768,N_4578);
and U5413 (N_5413,N_4773,N_4887);
nor U5414 (N_5414,N_4461,N_4811);
xnor U5415 (N_5415,N_4517,N_4832);
nor U5416 (N_5416,N_4796,N_4081);
or U5417 (N_5417,N_4200,N_4136);
and U5418 (N_5418,N_4551,N_4234);
nor U5419 (N_5419,N_4401,N_4180);
nand U5420 (N_5420,N_4065,N_4097);
nand U5421 (N_5421,N_4025,N_4720);
nor U5422 (N_5422,N_4207,N_4051);
and U5423 (N_5423,N_4981,N_4959);
and U5424 (N_5424,N_4970,N_4663);
nor U5425 (N_5425,N_4807,N_4588);
nand U5426 (N_5426,N_4537,N_4556);
and U5427 (N_5427,N_4612,N_4242);
nand U5428 (N_5428,N_4812,N_4616);
xor U5429 (N_5429,N_4161,N_4443);
nor U5430 (N_5430,N_4803,N_4835);
and U5431 (N_5431,N_4603,N_4206);
nor U5432 (N_5432,N_4471,N_4034);
and U5433 (N_5433,N_4332,N_4784);
and U5434 (N_5434,N_4868,N_4863);
nand U5435 (N_5435,N_4653,N_4029);
nor U5436 (N_5436,N_4976,N_4028);
nand U5437 (N_5437,N_4627,N_4861);
nor U5438 (N_5438,N_4524,N_4841);
nand U5439 (N_5439,N_4439,N_4123);
nor U5440 (N_5440,N_4719,N_4260);
nand U5441 (N_5441,N_4607,N_4233);
and U5442 (N_5442,N_4532,N_4037);
nor U5443 (N_5443,N_4504,N_4149);
nand U5444 (N_5444,N_4426,N_4483);
nor U5445 (N_5445,N_4848,N_4124);
or U5446 (N_5446,N_4845,N_4591);
or U5447 (N_5447,N_4285,N_4502);
and U5448 (N_5448,N_4501,N_4432);
nor U5449 (N_5449,N_4827,N_4466);
or U5450 (N_5450,N_4918,N_4645);
nand U5451 (N_5451,N_4725,N_4829);
nor U5452 (N_5452,N_4765,N_4538);
xnor U5453 (N_5453,N_4818,N_4531);
or U5454 (N_5454,N_4651,N_4077);
nand U5455 (N_5455,N_4031,N_4341);
and U5456 (N_5456,N_4866,N_4122);
or U5457 (N_5457,N_4908,N_4455);
nand U5458 (N_5458,N_4799,N_4318);
nor U5459 (N_5459,N_4825,N_4475);
or U5460 (N_5460,N_4569,N_4424);
nand U5461 (N_5461,N_4609,N_4484);
and U5462 (N_5462,N_4152,N_4946);
nor U5463 (N_5463,N_4422,N_4507);
and U5464 (N_5464,N_4735,N_4992);
nor U5465 (N_5465,N_4146,N_4844);
or U5466 (N_5466,N_4731,N_4440);
nand U5467 (N_5467,N_4173,N_4362);
or U5468 (N_5468,N_4227,N_4778);
nor U5469 (N_5469,N_4307,N_4174);
nand U5470 (N_5470,N_4886,N_4087);
nor U5471 (N_5471,N_4804,N_4379);
xnor U5472 (N_5472,N_4212,N_4477);
or U5473 (N_5473,N_4497,N_4447);
nor U5474 (N_5474,N_4402,N_4938);
xor U5475 (N_5475,N_4729,N_4993);
xor U5476 (N_5476,N_4089,N_4707);
or U5477 (N_5477,N_4621,N_4308);
and U5478 (N_5478,N_4036,N_4555);
or U5479 (N_5479,N_4717,N_4991);
or U5480 (N_5480,N_4823,N_4883);
nor U5481 (N_5481,N_4888,N_4533);
or U5482 (N_5482,N_4010,N_4922);
or U5483 (N_5483,N_4810,N_4944);
and U5484 (N_5484,N_4119,N_4456);
nand U5485 (N_5485,N_4581,N_4931);
nand U5486 (N_5486,N_4241,N_4964);
nand U5487 (N_5487,N_4994,N_4370);
nor U5488 (N_5488,N_4733,N_4548);
nand U5489 (N_5489,N_4577,N_4793);
nand U5490 (N_5490,N_4496,N_4708);
or U5491 (N_5491,N_4589,N_4027);
nand U5492 (N_5492,N_4839,N_4169);
nor U5493 (N_5493,N_4564,N_4463);
or U5494 (N_5494,N_4368,N_4972);
and U5495 (N_5495,N_4919,N_4248);
nor U5496 (N_5496,N_4925,N_4453);
nor U5497 (N_5497,N_4660,N_4809);
and U5498 (N_5498,N_4183,N_4713);
and U5499 (N_5499,N_4313,N_4265);
nand U5500 (N_5500,N_4915,N_4904);
and U5501 (N_5501,N_4979,N_4305);
nor U5502 (N_5502,N_4309,N_4851);
nand U5503 (N_5503,N_4312,N_4569);
nand U5504 (N_5504,N_4364,N_4006);
or U5505 (N_5505,N_4459,N_4838);
xor U5506 (N_5506,N_4739,N_4316);
or U5507 (N_5507,N_4926,N_4307);
xnor U5508 (N_5508,N_4418,N_4360);
nor U5509 (N_5509,N_4712,N_4422);
and U5510 (N_5510,N_4960,N_4361);
and U5511 (N_5511,N_4256,N_4155);
and U5512 (N_5512,N_4307,N_4002);
and U5513 (N_5513,N_4760,N_4516);
and U5514 (N_5514,N_4505,N_4105);
or U5515 (N_5515,N_4892,N_4181);
nor U5516 (N_5516,N_4655,N_4243);
and U5517 (N_5517,N_4146,N_4867);
nand U5518 (N_5518,N_4659,N_4938);
nand U5519 (N_5519,N_4049,N_4052);
nand U5520 (N_5520,N_4618,N_4344);
or U5521 (N_5521,N_4153,N_4650);
nand U5522 (N_5522,N_4626,N_4413);
and U5523 (N_5523,N_4482,N_4497);
or U5524 (N_5524,N_4034,N_4993);
or U5525 (N_5525,N_4858,N_4888);
nor U5526 (N_5526,N_4536,N_4311);
or U5527 (N_5527,N_4191,N_4476);
and U5528 (N_5528,N_4347,N_4345);
or U5529 (N_5529,N_4930,N_4935);
or U5530 (N_5530,N_4570,N_4417);
nand U5531 (N_5531,N_4946,N_4353);
nand U5532 (N_5532,N_4725,N_4405);
nand U5533 (N_5533,N_4122,N_4144);
and U5534 (N_5534,N_4400,N_4604);
nand U5535 (N_5535,N_4758,N_4334);
nand U5536 (N_5536,N_4377,N_4161);
and U5537 (N_5537,N_4393,N_4791);
or U5538 (N_5538,N_4661,N_4133);
and U5539 (N_5539,N_4005,N_4760);
and U5540 (N_5540,N_4567,N_4187);
nand U5541 (N_5541,N_4902,N_4439);
or U5542 (N_5542,N_4658,N_4572);
or U5543 (N_5543,N_4845,N_4101);
nand U5544 (N_5544,N_4856,N_4662);
or U5545 (N_5545,N_4118,N_4972);
nor U5546 (N_5546,N_4486,N_4448);
or U5547 (N_5547,N_4370,N_4922);
or U5548 (N_5548,N_4638,N_4117);
and U5549 (N_5549,N_4770,N_4119);
and U5550 (N_5550,N_4541,N_4564);
and U5551 (N_5551,N_4306,N_4245);
and U5552 (N_5552,N_4102,N_4839);
nand U5553 (N_5553,N_4169,N_4442);
nor U5554 (N_5554,N_4610,N_4770);
nand U5555 (N_5555,N_4963,N_4790);
nand U5556 (N_5556,N_4682,N_4623);
nor U5557 (N_5557,N_4620,N_4317);
or U5558 (N_5558,N_4191,N_4053);
nand U5559 (N_5559,N_4278,N_4353);
or U5560 (N_5560,N_4596,N_4721);
nor U5561 (N_5561,N_4505,N_4184);
and U5562 (N_5562,N_4080,N_4791);
and U5563 (N_5563,N_4029,N_4536);
or U5564 (N_5564,N_4415,N_4661);
or U5565 (N_5565,N_4377,N_4442);
nor U5566 (N_5566,N_4970,N_4380);
nand U5567 (N_5567,N_4167,N_4590);
nor U5568 (N_5568,N_4511,N_4328);
nand U5569 (N_5569,N_4791,N_4577);
nand U5570 (N_5570,N_4760,N_4918);
and U5571 (N_5571,N_4053,N_4583);
nand U5572 (N_5572,N_4203,N_4734);
nand U5573 (N_5573,N_4480,N_4324);
and U5574 (N_5574,N_4788,N_4766);
nand U5575 (N_5575,N_4600,N_4328);
or U5576 (N_5576,N_4079,N_4066);
nor U5577 (N_5577,N_4843,N_4494);
and U5578 (N_5578,N_4577,N_4764);
nand U5579 (N_5579,N_4358,N_4614);
nand U5580 (N_5580,N_4985,N_4394);
or U5581 (N_5581,N_4972,N_4374);
and U5582 (N_5582,N_4480,N_4182);
or U5583 (N_5583,N_4488,N_4486);
xnor U5584 (N_5584,N_4649,N_4887);
or U5585 (N_5585,N_4360,N_4818);
or U5586 (N_5586,N_4489,N_4298);
nor U5587 (N_5587,N_4710,N_4513);
or U5588 (N_5588,N_4826,N_4806);
nand U5589 (N_5589,N_4925,N_4295);
xnor U5590 (N_5590,N_4861,N_4925);
nor U5591 (N_5591,N_4887,N_4670);
nor U5592 (N_5592,N_4325,N_4809);
and U5593 (N_5593,N_4600,N_4026);
nand U5594 (N_5594,N_4333,N_4585);
or U5595 (N_5595,N_4340,N_4596);
xnor U5596 (N_5596,N_4525,N_4763);
or U5597 (N_5597,N_4606,N_4413);
nor U5598 (N_5598,N_4499,N_4313);
nand U5599 (N_5599,N_4192,N_4956);
nor U5600 (N_5600,N_4518,N_4916);
nor U5601 (N_5601,N_4832,N_4693);
or U5602 (N_5602,N_4354,N_4678);
nor U5603 (N_5603,N_4814,N_4440);
and U5604 (N_5604,N_4545,N_4610);
or U5605 (N_5605,N_4891,N_4680);
and U5606 (N_5606,N_4749,N_4886);
nor U5607 (N_5607,N_4416,N_4128);
and U5608 (N_5608,N_4645,N_4507);
nor U5609 (N_5609,N_4615,N_4851);
nor U5610 (N_5610,N_4568,N_4935);
nor U5611 (N_5611,N_4084,N_4605);
nor U5612 (N_5612,N_4753,N_4303);
nand U5613 (N_5613,N_4561,N_4421);
and U5614 (N_5614,N_4480,N_4439);
xor U5615 (N_5615,N_4219,N_4838);
or U5616 (N_5616,N_4047,N_4402);
nor U5617 (N_5617,N_4306,N_4036);
nand U5618 (N_5618,N_4347,N_4128);
and U5619 (N_5619,N_4192,N_4591);
and U5620 (N_5620,N_4069,N_4886);
and U5621 (N_5621,N_4977,N_4384);
and U5622 (N_5622,N_4713,N_4190);
nor U5623 (N_5623,N_4385,N_4653);
nand U5624 (N_5624,N_4486,N_4047);
xor U5625 (N_5625,N_4194,N_4668);
or U5626 (N_5626,N_4797,N_4734);
nor U5627 (N_5627,N_4496,N_4906);
nand U5628 (N_5628,N_4246,N_4009);
and U5629 (N_5629,N_4922,N_4558);
xor U5630 (N_5630,N_4603,N_4402);
or U5631 (N_5631,N_4416,N_4503);
or U5632 (N_5632,N_4493,N_4799);
nand U5633 (N_5633,N_4305,N_4181);
or U5634 (N_5634,N_4366,N_4972);
or U5635 (N_5635,N_4983,N_4570);
nor U5636 (N_5636,N_4216,N_4185);
or U5637 (N_5637,N_4984,N_4509);
xnor U5638 (N_5638,N_4764,N_4502);
nand U5639 (N_5639,N_4724,N_4274);
and U5640 (N_5640,N_4604,N_4884);
or U5641 (N_5641,N_4421,N_4067);
nand U5642 (N_5642,N_4643,N_4583);
and U5643 (N_5643,N_4187,N_4972);
nor U5644 (N_5644,N_4325,N_4551);
nor U5645 (N_5645,N_4449,N_4368);
xor U5646 (N_5646,N_4692,N_4638);
nor U5647 (N_5647,N_4888,N_4429);
and U5648 (N_5648,N_4896,N_4271);
and U5649 (N_5649,N_4201,N_4237);
and U5650 (N_5650,N_4684,N_4676);
nand U5651 (N_5651,N_4870,N_4444);
and U5652 (N_5652,N_4940,N_4934);
and U5653 (N_5653,N_4397,N_4486);
or U5654 (N_5654,N_4241,N_4540);
xor U5655 (N_5655,N_4375,N_4025);
nand U5656 (N_5656,N_4673,N_4749);
and U5657 (N_5657,N_4148,N_4780);
or U5658 (N_5658,N_4546,N_4189);
or U5659 (N_5659,N_4774,N_4544);
and U5660 (N_5660,N_4788,N_4634);
and U5661 (N_5661,N_4531,N_4226);
nand U5662 (N_5662,N_4148,N_4865);
or U5663 (N_5663,N_4310,N_4369);
or U5664 (N_5664,N_4428,N_4925);
nor U5665 (N_5665,N_4587,N_4565);
and U5666 (N_5666,N_4204,N_4955);
nor U5667 (N_5667,N_4594,N_4258);
nand U5668 (N_5668,N_4120,N_4380);
or U5669 (N_5669,N_4683,N_4947);
nor U5670 (N_5670,N_4380,N_4780);
xnor U5671 (N_5671,N_4368,N_4308);
xnor U5672 (N_5672,N_4057,N_4763);
xnor U5673 (N_5673,N_4215,N_4471);
or U5674 (N_5674,N_4982,N_4663);
nor U5675 (N_5675,N_4713,N_4739);
and U5676 (N_5676,N_4259,N_4898);
nand U5677 (N_5677,N_4819,N_4500);
or U5678 (N_5678,N_4495,N_4769);
and U5679 (N_5679,N_4046,N_4432);
nor U5680 (N_5680,N_4881,N_4857);
nor U5681 (N_5681,N_4715,N_4156);
nor U5682 (N_5682,N_4649,N_4118);
and U5683 (N_5683,N_4134,N_4900);
and U5684 (N_5684,N_4048,N_4731);
nand U5685 (N_5685,N_4131,N_4973);
nand U5686 (N_5686,N_4691,N_4702);
nor U5687 (N_5687,N_4284,N_4030);
nor U5688 (N_5688,N_4700,N_4814);
nor U5689 (N_5689,N_4348,N_4510);
xor U5690 (N_5690,N_4430,N_4026);
or U5691 (N_5691,N_4034,N_4384);
nand U5692 (N_5692,N_4177,N_4751);
and U5693 (N_5693,N_4665,N_4682);
and U5694 (N_5694,N_4202,N_4068);
and U5695 (N_5695,N_4578,N_4319);
nand U5696 (N_5696,N_4951,N_4249);
nand U5697 (N_5697,N_4847,N_4841);
nand U5698 (N_5698,N_4976,N_4463);
or U5699 (N_5699,N_4334,N_4694);
and U5700 (N_5700,N_4581,N_4970);
xnor U5701 (N_5701,N_4373,N_4085);
nor U5702 (N_5702,N_4130,N_4576);
and U5703 (N_5703,N_4091,N_4267);
or U5704 (N_5704,N_4968,N_4794);
xor U5705 (N_5705,N_4257,N_4853);
or U5706 (N_5706,N_4278,N_4991);
and U5707 (N_5707,N_4333,N_4749);
nor U5708 (N_5708,N_4985,N_4729);
nor U5709 (N_5709,N_4010,N_4916);
and U5710 (N_5710,N_4476,N_4252);
nor U5711 (N_5711,N_4039,N_4562);
and U5712 (N_5712,N_4759,N_4243);
or U5713 (N_5713,N_4477,N_4373);
xor U5714 (N_5714,N_4078,N_4416);
nand U5715 (N_5715,N_4675,N_4509);
nor U5716 (N_5716,N_4439,N_4198);
and U5717 (N_5717,N_4157,N_4203);
nand U5718 (N_5718,N_4184,N_4501);
and U5719 (N_5719,N_4577,N_4677);
or U5720 (N_5720,N_4829,N_4098);
or U5721 (N_5721,N_4253,N_4626);
and U5722 (N_5722,N_4929,N_4241);
nand U5723 (N_5723,N_4815,N_4299);
xnor U5724 (N_5724,N_4947,N_4952);
and U5725 (N_5725,N_4707,N_4357);
nand U5726 (N_5726,N_4178,N_4757);
or U5727 (N_5727,N_4110,N_4075);
or U5728 (N_5728,N_4096,N_4884);
and U5729 (N_5729,N_4696,N_4197);
xor U5730 (N_5730,N_4791,N_4799);
or U5731 (N_5731,N_4645,N_4252);
and U5732 (N_5732,N_4454,N_4719);
and U5733 (N_5733,N_4141,N_4630);
nand U5734 (N_5734,N_4698,N_4144);
nor U5735 (N_5735,N_4292,N_4491);
nand U5736 (N_5736,N_4698,N_4366);
or U5737 (N_5737,N_4904,N_4712);
nor U5738 (N_5738,N_4535,N_4919);
or U5739 (N_5739,N_4950,N_4273);
or U5740 (N_5740,N_4296,N_4970);
nor U5741 (N_5741,N_4325,N_4957);
nor U5742 (N_5742,N_4867,N_4434);
or U5743 (N_5743,N_4172,N_4593);
or U5744 (N_5744,N_4453,N_4980);
and U5745 (N_5745,N_4382,N_4999);
nor U5746 (N_5746,N_4196,N_4958);
nand U5747 (N_5747,N_4946,N_4180);
or U5748 (N_5748,N_4610,N_4231);
or U5749 (N_5749,N_4046,N_4379);
nand U5750 (N_5750,N_4618,N_4276);
nand U5751 (N_5751,N_4986,N_4812);
and U5752 (N_5752,N_4513,N_4758);
or U5753 (N_5753,N_4629,N_4663);
and U5754 (N_5754,N_4507,N_4803);
nand U5755 (N_5755,N_4295,N_4547);
and U5756 (N_5756,N_4962,N_4996);
nand U5757 (N_5757,N_4089,N_4950);
nand U5758 (N_5758,N_4968,N_4888);
or U5759 (N_5759,N_4196,N_4373);
or U5760 (N_5760,N_4870,N_4951);
nor U5761 (N_5761,N_4369,N_4302);
or U5762 (N_5762,N_4254,N_4884);
nor U5763 (N_5763,N_4225,N_4418);
nand U5764 (N_5764,N_4384,N_4677);
xnor U5765 (N_5765,N_4162,N_4586);
or U5766 (N_5766,N_4378,N_4411);
xnor U5767 (N_5767,N_4615,N_4564);
xnor U5768 (N_5768,N_4842,N_4963);
and U5769 (N_5769,N_4831,N_4435);
and U5770 (N_5770,N_4952,N_4783);
nand U5771 (N_5771,N_4470,N_4271);
nor U5772 (N_5772,N_4408,N_4133);
nor U5773 (N_5773,N_4940,N_4812);
nand U5774 (N_5774,N_4170,N_4654);
nand U5775 (N_5775,N_4983,N_4777);
xor U5776 (N_5776,N_4962,N_4764);
or U5777 (N_5777,N_4702,N_4687);
nor U5778 (N_5778,N_4138,N_4420);
xor U5779 (N_5779,N_4444,N_4707);
nor U5780 (N_5780,N_4852,N_4175);
and U5781 (N_5781,N_4715,N_4143);
nor U5782 (N_5782,N_4362,N_4782);
nor U5783 (N_5783,N_4561,N_4070);
nor U5784 (N_5784,N_4754,N_4054);
nor U5785 (N_5785,N_4620,N_4587);
and U5786 (N_5786,N_4579,N_4470);
nand U5787 (N_5787,N_4711,N_4790);
or U5788 (N_5788,N_4822,N_4416);
and U5789 (N_5789,N_4856,N_4021);
and U5790 (N_5790,N_4907,N_4316);
nor U5791 (N_5791,N_4242,N_4419);
xnor U5792 (N_5792,N_4154,N_4720);
nor U5793 (N_5793,N_4050,N_4547);
xor U5794 (N_5794,N_4660,N_4737);
nor U5795 (N_5795,N_4037,N_4402);
or U5796 (N_5796,N_4947,N_4176);
nand U5797 (N_5797,N_4966,N_4737);
and U5798 (N_5798,N_4787,N_4390);
xor U5799 (N_5799,N_4365,N_4616);
and U5800 (N_5800,N_4155,N_4083);
and U5801 (N_5801,N_4614,N_4177);
nand U5802 (N_5802,N_4953,N_4767);
nor U5803 (N_5803,N_4117,N_4752);
and U5804 (N_5804,N_4988,N_4860);
nor U5805 (N_5805,N_4717,N_4589);
and U5806 (N_5806,N_4050,N_4413);
nand U5807 (N_5807,N_4235,N_4990);
nor U5808 (N_5808,N_4760,N_4090);
nor U5809 (N_5809,N_4819,N_4333);
nor U5810 (N_5810,N_4886,N_4439);
and U5811 (N_5811,N_4783,N_4924);
and U5812 (N_5812,N_4990,N_4683);
and U5813 (N_5813,N_4740,N_4250);
and U5814 (N_5814,N_4689,N_4850);
nand U5815 (N_5815,N_4743,N_4570);
nand U5816 (N_5816,N_4344,N_4085);
nor U5817 (N_5817,N_4097,N_4076);
nor U5818 (N_5818,N_4205,N_4065);
nand U5819 (N_5819,N_4616,N_4078);
nand U5820 (N_5820,N_4910,N_4991);
or U5821 (N_5821,N_4318,N_4438);
nor U5822 (N_5822,N_4929,N_4582);
nand U5823 (N_5823,N_4086,N_4802);
nand U5824 (N_5824,N_4260,N_4692);
and U5825 (N_5825,N_4725,N_4332);
or U5826 (N_5826,N_4914,N_4217);
nor U5827 (N_5827,N_4086,N_4059);
nor U5828 (N_5828,N_4970,N_4561);
and U5829 (N_5829,N_4212,N_4713);
or U5830 (N_5830,N_4497,N_4651);
nand U5831 (N_5831,N_4476,N_4162);
nand U5832 (N_5832,N_4419,N_4420);
nand U5833 (N_5833,N_4137,N_4046);
nand U5834 (N_5834,N_4685,N_4281);
xnor U5835 (N_5835,N_4078,N_4193);
and U5836 (N_5836,N_4280,N_4164);
or U5837 (N_5837,N_4055,N_4342);
and U5838 (N_5838,N_4272,N_4670);
or U5839 (N_5839,N_4965,N_4702);
xor U5840 (N_5840,N_4755,N_4866);
and U5841 (N_5841,N_4529,N_4103);
and U5842 (N_5842,N_4758,N_4545);
nor U5843 (N_5843,N_4108,N_4860);
nor U5844 (N_5844,N_4652,N_4386);
and U5845 (N_5845,N_4045,N_4273);
xor U5846 (N_5846,N_4865,N_4336);
nor U5847 (N_5847,N_4643,N_4485);
and U5848 (N_5848,N_4988,N_4371);
nor U5849 (N_5849,N_4845,N_4761);
nor U5850 (N_5850,N_4321,N_4274);
or U5851 (N_5851,N_4859,N_4500);
or U5852 (N_5852,N_4039,N_4551);
nor U5853 (N_5853,N_4946,N_4497);
and U5854 (N_5854,N_4384,N_4581);
nor U5855 (N_5855,N_4930,N_4579);
nor U5856 (N_5856,N_4210,N_4955);
and U5857 (N_5857,N_4700,N_4164);
nor U5858 (N_5858,N_4632,N_4335);
and U5859 (N_5859,N_4778,N_4192);
nor U5860 (N_5860,N_4393,N_4475);
and U5861 (N_5861,N_4092,N_4329);
or U5862 (N_5862,N_4883,N_4505);
and U5863 (N_5863,N_4767,N_4867);
nor U5864 (N_5864,N_4291,N_4865);
nor U5865 (N_5865,N_4088,N_4070);
or U5866 (N_5866,N_4430,N_4806);
and U5867 (N_5867,N_4997,N_4806);
and U5868 (N_5868,N_4069,N_4726);
or U5869 (N_5869,N_4782,N_4049);
or U5870 (N_5870,N_4274,N_4570);
nor U5871 (N_5871,N_4486,N_4285);
nor U5872 (N_5872,N_4235,N_4654);
nand U5873 (N_5873,N_4765,N_4232);
nand U5874 (N_5874,N_4490,N_4689);
nand U5875 (N_5875,N_4798,N_4378);
and U5876 (N_5876,N_4239,N_4045);
nor U5877 (N_5877,N_4851,N_4138);
nor U5878 (N_5878,N_4857,N_4408);
or U5879 (N_5879,N_4390,N_4369);
and U5880 (N_5880,N_4792,N_4016);
nor U5881 (N_5881,N_4204,N_4499);
nand U5882 (N_5882,N_4115,N_4027);
nand U5883 (N_5883,N_4162,N_4581);
nand U5884 (N_5884,N_4603,N_4510);
nor U5885 (N_5885,N_4523,N_4277);
nor U5886 (N_5886,N_4222,N_4402);
xnor U5887 (N_5887,N_4523,N_4967);
and U5888 (N_5888,N_4867,N_4277);
nand U5889 (N_5889,N_4133,N_4753);
nor U5890 (N_5890,N_4091,N_4766);
and U5891 (N_5891,N_4858,N_4086);
and U5892 (N_5892,N_4763,N_4283);
xor U5893 (N_5893,N_4517,N_4794);
and U5894 (N_5894,N_4072,N_4809);
xnor U5895 (N_5895,N_4274,N_4884);
xnor U5896 (N_5896,N_4884,N_4440);
nor U5897 (N_5897,N_4683,N_4700);
or U5898 (N_5898,N_4605,N_4216);
and U5899 (N_5899,N_4062,N_4442);
nand U5900 (N_5900,N_4749,N_4288);
nor U5901 (N_5901,N_4054,N_4651);
and U5902 (N_5902,N_4477,N_4906);
nor U5903 (N_5903,N_4299,N_4706);
nand U5904 (N_5904,N_4088,N_4403);
or U5905 (N_5905,N_4703,N_4334);
or U5906 (N_5906,N_4320,N_4103);
and U5907 (N_5907,N_4909,N_4816);
or U5908 (N_5908,N_4097,N_4441);
nand U5909 (N_5909,N_4520,N_4940);
nor U5910 (N_5910,N_4113,N_4046);
nand U5911 (N_5911,N_4922,N_4011);
xnor U5912 (N_5912,N_4927,N_4986);
nand U5913 (N_5913,N_4744,N_4092);
nor U5914 (N_5914,N_4728,N_4415);
and U5915 (N_5915,N_4688,N_4259);
xor U5916 (N_5916,N_4645,N_4150);
xor U5917 (N_5917,N_4913,N_4420);
nand U5918 (N_5918,N_4265,N_4492);
nor U5919 (N_5919,N_4791,N_4115);
and U5920 (N_5920,N_4171,N_4111);
and U5921 (N_5921,N_4004,N_4603);
nor U5922 (N_5922,N_4187,N_4568);
and U5923 (N_5923,N_4567,N_4917);
xnor U5924 (N_5924,N_4323,N_4779);
nand U5925 (N_5925,N_4391,N_4944);
nor U5926 (N_5926,N_4788,N_4118);
nand U5927 (N_5927,N_4968,N_4463);
xor U5928 (N_5928,N_4763,N_4221);
or U5929 (N_5929,N_4284,N_4913);
nand U5930 (N_5930,N_4898,N_4521);
nor U5931 (N_5931,N_4587,N_4051);
nand U5932 (N_5932,N_4254,N_4206);
and U5933 (N_5933,N_4751,N_4863);
nor U5934 (N_5934,N_4184,N_4800);
and U5935 (N_5935,N_4719,N_4278);
or U5936 (N_5936,N_4284,N_4151);
nor U5937 (N_5937,N_4593,N_4572);
and U5938 (N_5938,N_4869,N_4813);
xnor U5939 (N_5939,N_4890,N_4325);
nor U5940 (N_5940,N_4414,N_4967);
nor U5941 (N_5941,N_4983,N_4613);
nand U5942 (N_5942,N_4084,N_4402);
xor U5943 (N_5943,N_4273,N_4961);
nor U5944 (N_5944,N_4021,N_4641);
and U5945 (N_5945,N_4966,N_4621);
nand U5946 (N_5946,N_4663,N_4365);
or U5947 (N_5947,N_4595,N_4199);
nand U5948 (N_5948,N_4677,N_4076);
nor U5949 (N_5949,N_4742,N_4549);
or U5950 (N_5950,N_4922,N_4039);
or U5951 (N_5951,N_4943,N_4414);
and U5952 (N_5952,N_4130,N_4166);
nand U5953 (N_5953,N_4985,N_4473);
or U5954 (N_5954,N_4492,N_4635);
nand U5955 (N_5955,N_4217,N_4483);
and U5956 (N_5956,N_4770,N_4530);
or U5957 (N_5957,N_4013,N_4559);
nand U5958 (N_5958,N_4191,N_4220);
nand U5959 (N_5959,N_4874,N_4424);
nand U5960 (N_5960,N_4618,N_4897);
and U5961 (N_5961,N_4291,N_4775);
nand U5962 (N_5962,N_4419,N_4974);
or U5963 (N_5963,N_4960,N_4744);
and U5964 (N_5964,N_4683,N_4384);
xor U5965 (N_5965,N_4130,N_4017);
nand U5966 (N_5966,N_4885,N_4044);
or U5967 (N_5967,N_4252,N_4191);
nor U5968 (N_5968,N_4741,N_4168);
or U5969 (N_5969,N_4152,N_4474);
nand U5970 (N_5970,N_4152,N_4142);
and U5971 (N_5971,N_4492,N_4329);
nand U5972 (N_5972,N_4025,N_4806);
nor U5973 (N_5973,N_4323,N_4098);
nor U5974 (N_5974,N_4386,N_4950);
and U5975 (N_5975,N_4269,N_4365);
and U5976 (N_5976,N_4768,N_4620);
and U5977 (N_5977,N_4654,N_4210);
nand U5978 (N_5978,N_4240,N_4968);
and U5979 (N_5979,N_4828,N_4101);
or U5980 (N_5980,N_4602,N_4957);
or U5981 (N_5981,N_4931,N_4937);
nand U5982 (N_5982,N_4805,N_4697);
and U5983 (N_5983,N_4379,N_4036);
and U5984 (N_5984,N_4943,N_4250);
and U5985 (N_5985,N_4965,N_4097);
or U5986 (N_5986,N_4871,N_4675);
and U5987 (N_5987,N_4996,N_4719);
and U5988 (N_5988,N_4482,N_4719);
nor U5989 (N_5989,N_4372,N_4205);
nor U5990 (N_5990,N_4366,N_4056);
nand U5991 (N_5991,N_4168,N_4201);
or U5992 (N_5992,N_4173,N_4177);
or U5993 (N_5993,N_4696,N_4382);
xor U5994 (N_5994,N_4130,N_4789);
nand U5995 (N_5995,N_4609,N_4051);
nor U5996 (N_5996,N_4081,N_4924);
nand U5997 (N_5997,N_4791,N_4380);
nand U5998 (N_5998,N_4042,N_4806);
nand U5999 (N_5999,N_4810,N_4617);
nand U6000 (N_6000,N_5031,N_5674);
nand U6001 (N_6001,N_5096,N_5286);
and U6002 (N_6002,N_5394,N_5464);
and U6003 (N_6003,N_5379,N_5959);
nor U6004 (N_6004,N_5566,N_5429);
or U6005 (N_6005,N_5458,N_5479);
nand U6006 (N_6006,N_5795,N_5625);
nand U6007 (N_6007,N_5956,N_5687);
nor U6008 (N_6008,N_5125,N_5537);
nand U6009 (N_6009,N_5898,N_5772);
nor U6010 (N_6010,N_5565,N_5536);
xor U6011 (N_6011,N_5268,N_5299);
nand U6012 (N_6012,N_5645,N_5166);
or U6013 (N_6013,N_5076,N_5719);
and U6014 (N_6014,N_5315,N_5177);
or U6015 (N_6015,N_5685,N_5235);
nor U6016 (N_6016,N_5401,N_5095);
nand U6017 (N_6017,N_5936,N_5468);
or U6018 (N_6018,N_5373,N_5875);
and U6019 (N_6019,N_5688,N_5664);
nor U6020 (N_6020,N_5984,N_5253);
nand U6021 (N_6021,N_5261,N_5508);
nand U6022 (N_6022,N_5994,N_5644);
and U6023 (N_6023,N_5215,N_5162);
nand U6024 (N_6024,N_5525,N_5749);
xnor U6025 (N_6025,N_5143,N_5917);
and U6026 (N_6026,N_5836,N_5060);
and U6027 (N_6027,N_5927,N_5758);
nand U6028 (N_6028,N_5196,N_5888);
nor U6029 (N_6029,N_5928,N_5078);
nand U6030 (N_6030,N_5856,N_5652);
and U6031 (N_6031,N_5270,N_5399);
nand U6032 (N_6032,N_5336,N_5209);
nor U6033 (N_6033,N_5707,N_5668);
xor U6034 (N_6034,N_5939,N_5821);
or U6035 (N_6035,N_5460,N_5382);
nand U6036 (N_6036,N_5179,N_5037);
xnor U6037 (N_6037,N_5459,N_5388);
nor U6038 (N_6038,N_5280,N_5436);
or U6039 (N_6039,N_5481,N_5937);
or U6040 (N_6040,N_5365,N_5509);
nor U6041 (N_6041,N_5904,N_5183);
nor U6042 (N_6042,N_5922,N_5540);
nand U6043 (N_6043,N_5755,N_5395);
or U6044 (N_6044,N_5328,N_5899);
and U6045 (N_6045,N_5249,N_5977);
xnor U6046 (N_6046,N_5543,N_5329);
and U6047 (N_6047,N_5036,N_5351);
nand U6048 (N_6048,N_5194,N_5971);
or U6049 (N_6049,N_5420,N_5594);
or U6050 (N_6050,N_5488,N_5042);
or U6051 (N_6051,N_5045,N_5083);
xnor U6052 (N_6052,N_5406,N_5014);
nand U6053 (N_6053,N_5756,N_5841);
nor U6054 (N_6054,N_5448,N_5062);
nor U6055 (N_6055,N_5752,N_5891);
nand U6056 (N_6056,N_5578,N_5846);
xnor U6057 (N_6057,N_5414,N_5759);
or U6058 (N_6058,N_5628,N_5112);
and U6059 (N_6059,N_5829,N_5575);
nor U6060 (N_6060,N_5943,N_5346);
or U6061 (N_6061,N_5156,N_5483);
or U6062 (N_6062,N_5213,N_5326);
xor U6063 (N_6063,N_5485,N_5848);
nor U6064 (N_6064,N_5728,N_5616);
nor U6065 (N_6065,N_5981,N_5426);
nand U6066 (N_6066,N_5779,N_5562);
nor U6067 (N_6067,N_5858,N_5808);
and U6068 (N_6068,N_5761,N_5195);
nor U6069 (N_6069,N_5202,N_5842);
and U6070 (N_6070,N_5504,N_5149);
nor U6071 (N_6071,N_5544,N_5725);
nand U6072 (N_6072,N_5600,N_5975);
and U6073 (N_6073,N_5925,N_5090);
nand U6074 (N_6074,N_5558,N_5840);
or U6075 (N_6075,N_5234,N_5965);
nor U6076 (N_6076,N_5265,N_5358);
and U6077 (N_6077,N_5513,N_5774);
or U6078 (N_6078,N_5952,N_5340);
nand U6079 (N_6079,N_5785,N_5053);
xor U6080 (N_6080,N_5342,N_5816);
nor U6081 (N_6081,N_5665,N_5659);
and U6082 (N_6082,N_5757,N_5839);
and U6083 (N_6083,N_5080,N_5916);
nor U6084 (N_6084,N_5963,N_5622);
or U6085 (N_6085,N_5325,N_5990);
nand U6086 (N_6086,N_5244,N_5519);
nor U6087 (N_6087,N_5911,N_5822);
nor U6088 (N_6088,N_5626,N_5692);
and U6089 (N_6089,N_5029,N_5642);
and U6090 (N_6090,N_5871,N_5114);
nand U6091 (N_6091,N_5735,N_5109);
nor U6092 (N_6092,N_5180,N_5199);
and U6093 (N_6093,N_5577,N_5022);
and U6094 (N_6094,N_5750,N_5237);
or U6095 (N_6095,N_5775,N_5371);
or U6096 (N_6096,N_5520,N_5119);
nand U6097 (N_6097,N_5410,N_5876);
or U6098 (N_6098,N_5833,N_5717);
nor U6099 (N_6099,N_5059,N_5834);
xor U6100 (N_6100,N_5219,N_5563);
nor U6101 (N_6101,N_5417,N_5592);
nor U6102 (N_6102,N_5776,N_5976);
nand U6103 (N_6103,N_5847,N_5352);
nand U6104 (N_6104,N_5857,N_5948);
and U6105 (N_6105,N_5350,N_5819);
nor U6106 (N_6106,N_5689,N_5812);
or U6107 (N_6107,N_5356,N_5013);
or U6108 (N_6108,N_5434,N_5670);
nand U6109 (N_6109,N_5500,N_5309);
nor U6110 (N_6110,N_5285,N_5661);
and U6111 (N_6111,N_5969,N_5451);
or U6112 (N_6112,N_5453,N_5103);
or U6113 (N_6113,N_5556,N_5535);
nor U6114 (N_6114,N_5027,N_5683);
nor U6115 (N_6115,N_5100,N_5548);
xor U6116 (N_6116,N_5933,N_5903);
or U6117 (N_6117,N_5621,N_5318);
nand U6118 (N_6118,N_5967,N_5257);
or U6119 (N_6119,N_5361,N_5985);
nor U6120 (N_6120,N_5929,N_5258);
nand U6121 (N_6121,N_5667,N_5026);
or U6122 (N_6122,N_5307,N_5678);
nand U6123 (N_6123,N_5501,N_5471);
or U6124 (N_6124,N_5455,N_5657);
or U6125 (N_6125,N_5810,N_5961);
nand U6126 (N_6126,N_5355,N_5383);
and U6127 (N_6127,N_5363,N_5568);
nor U6128 (N_6128,N_5739,N_5989);
xnor U6129 (N_6129,N_5153,N_5113);
nor U6130 (N_6130,N_5514,N_5945);
or U6131 (N_6131,N_5206,N_5806);
xnor U6132 (N_6132,N_5901,N_5999);
nor U6133 (N_6133,N_5389,N_5932);
nand U6134 (N_6134,N_5102,N_5276);
or U6135 (N_6135,N_5730,N_5020);
nor U6136 (N_6136,N_5854,N_5518);
nor U6137 (N_6137,N_5175,N_5762);
or U6138 (N_6138,N_5482,N_5324);
or U6139 (N_6139,N_5962,N_5597);
and U6140 (N_6140,N_5546,N_5450);
or U6141 (N_6141,N_5827,N_5461);
and U6142 (N_6142,N_5416,N_5765);
nor U6143 (N_6143,N_5569,N_5243);
nor U6144 (N_6144,N_5647,N_5691);
xor U6145 (N_6145,N_5151,N_5968);
or U6146 (N_6146,N_5317,N_5279);
or U6147 (N_6147,N_5579,N_5002);
and U6148 (N_6148,N_5905,N_5353);
and U6149 (N_6149,N_5127,N_5487);
or U6150 (N_6150,N_5145,N_5710);
nor U6151 (N_6151,N_5019,N_5826);
or U6152 (N_6152,N_5718,N_5696);
xnor U6153 (N_6153,N_5559,N_5646);
and U6154 (N_6154,N_5748,N_5233);
nor U6155 (N_6155,N_5190,N_5720);
nand U6156 (N_6156,N_5295,N_5079);
and U6157 (N_6157,N_5220,N_5596);
and U6158 (N_6158,N_5672,N_5723);
or U6159 (N_6159,N_5385,N_5239);
and U6160 (N_6160,N_5919,N_5470);
nor U6161 (N_6161,N_5906,N_5517);
nand U6162 (N_6162,N_5868,N_5413);
and U6163 (N_6163,N_5030,N_5666);
and U6164 (N_6164,N_5960,N_5835);
or U6165 (N_6165,N_5791,N_5660);
or U6166 (N_6166,N_5466,N_5275);
xor U6167 (N_6167,N_5743,N_5915);
and U6168 (N_6168,N_5955,N_5217);
and U6169 (N_6169,N_5516,N_5110);
and U6170 (N_6170,N_5882,N_5530);
nor U6171 (N_6171,N_5944,N_5983);
or U6172 (N_6172,N_5675,N_5040);
xor U6173 (N_6173,N_5116,N_5377);
nand U6174 (N_6174,N_5094,N_5506);
or U6175 (N_6175,N_5585,N_5527);
xor U6176 (N_6176,N_5640,N_5910);
nor U6177 (N_6177,N_5368,N_5804);
nor U6178 (N_6178,N_5015,N_5740);
xnor U6179 (N_6179,N_5892,N_5281);
nand U6180 (N_6180,N_5551,N_5139);
and U6181 (N_6181,N_5278,N_5005);
or U6182 (N_6182,N_5751,N_5337);
nor U6183 (N_6183,N_5150,N_5447);
or U6184 (N_6184,N_5711,N_5864);
nor U6185 (N_6185,N_5953,N_5421);
nand U6186 (N_6186,N_5082,N_5669);
and U6187 (N_6187,N_5160,N_5742);
xnor U6188 (N_6188,N_5721,N_5753);
nand U6189 (N_6189,N_5218,N_5115);
nor U6190 (N_6190,N_5547,N_5741);
nand U6191 (N_6191,N_5402,N_5860);
nor U6192 (N_6192,N_5247,N_5021);
nand U6193 (N_6193,N_5084,N_5849);
nand U6194 (N_6194,N_5574,N_5273);
and U6195 (N_6195,N_5690,N_5771);
or U6196 (N_6196,N_5529,N_5148);
or U6197 (N_6197,N_5679,N_5250);
nand U6198 (N_6198,N_5226,N_5722);
nor U6199 (N_6199,N_5267,N_5809);
or U6200 (N_6200,N_5706,N_5161);
nor U6201 (N_6201,N_5651,N_5634);
nand U6202 (N_6202,N_5372,N_5503);
and U6203 (N_6203,N_5798,N_5302);
and U6204 (N_6204,N_5982,N_5935);
or U6205 (N_6205,N_5497,N_5957);
and U6206 (N_6206,N_5445,N_5890);
or U6207 (N_6207,N_5044,N_5418);
nand U6208 (N_6208,N_5778,N_5400);
and U6209 (N_6209,N_5843,N_5381);
and U6210 (N_6210,N_5908,N_5222);
nor U6211 (N_6211,N_5629,N_5820);
or U6212 (N_6212,N_5870,N_5088);
or U6213 (N_6213,N_5242,N_5620);
nor U6214 (N_6214,N_5940,N_5705);
nor U6215 (N_6215,N_5462,N_5437);
nand U6216 (N_6216,N_5442,N_5091);
nand U6217 (N_6217,N_5913,N_5004);
or U6218 (N_6218,N_5224,N_5476);
nand U6219 (N_6219,N_5188,N_5931);
xor U6220 (N_6220,N_5205,N_5650);
and U6221 (N_6221,N_5522,N_5154);
nand U6222 (N_6222,N_5131,N_5073);
nand U6223 (N_6223,N_5996,N_5000);
or U6224 (N_6224,N_5554,N_5713);
and U6225 (N_6225,N_5168,N_5902);
or U6226 (N_6226,N_5287,N_5251);
or U6227 (N_6227,N_5736,N_5425);
nor U6228 (N_6228,N_5700,N_5282);
nor U6229 (N_6229,N_5502,N_5314);
and U6230 (N_6230,N_5704,N_5814);
nand U6231 (N_6231,N_5452,N_5256);
nor U6232 (N_6232,N_5946,N_5375);
nand U6233 (N_6233,N_5232,N_5298);
nand U6234 (N_6234,N_5553,N_5972);
and U6235 (N_6235,N_5889,N_5731);
nor U6236 (N_6236,N_5283,N_5354);
and U6237 (N_6237,N_5055,N_5874);
and U6238 (N_6238,N_5435,N_5788);
and U6239 (N_6239,N_5011,N_5494);
nor U6240 (N_6240,N_5297,N_5631);
and U6241 (N_6241,N_5069,N_5693);
xor U6242 (N_6242,N_5316,N_5245);
nand U6243 (N_6243,N_5167,N_5321);
nand U6244 (N_6244,N_5236,N_5894);
and U6245 (N_6245,N_5310,N_5066);
or U6246 (N_6246,N_5998,N_5225);
nor U6247 (N_6247,N_5305,N_5699);
and U6248 (N_6248,N_5893,N_5773);
nand U6249 (N_6249,N_5920,N_5058);
or U6250 (N_6250,N_5763,N_5942);
nor U6251 (N_6251,N_5813,N_5465);
nor U6252 (N_6252,N_5591,N_5724);
or U6253 (N_6253,N_5863,N_5671);
nor U6254 (N_6254,N_5319,N_5648);
nor U6255 (N_6255,N_5051,N_5701);
nand U6256 (N_6256,N_5738,N_5880);
or U6257 (N_6257,N_5580,N_5786);
nor U6258 (N_6258,N_5266,N_5797);
and U6259 (N_6259,N_5469,N_5018);
or U6260 (N_6260,N_5056,N_5966);
and U6261 (N_6261,N_5680,N_5432);
nor U6262 (N_6262,N_5627,N_5170);
xor U6263 (N_6263,N_5312,N_5122);
or U6264 (N_6264,N_5292,N_5539);
nand U6265 (N_6265,N_5612,N_5284);
nand U6266 (N_6266,N_5768,N_5092);
and U6267 (N_6267,N_5837,N_5567);
nor U6268 (N_6268,N_5866,N_5089);
or U6269 (N_6269,N_5885,N_5008);
nor U6270 (N_6270,N_5802,N_5473);
and U6271 (N_6271,N_5490,N_5698);
nand U6272 (N_6272,N_5048,N_5493);
or U6273 (N_6273,N_5884,N_5941);
or U6274 (N_6274,N_5238,N_5992);
nor U6275 (N_6275,N_5979,N_5193);
nor U6276 (N_6276,N_5611,N_5964);
nand U6277 (N_6277,N_5378,N_5737);
nand U6278 (N_6278,N_5534,N_5189);
or U6279 (N_6279,N_5792,N_5587);
and U6280 (N_6280,N_5552,N_5571);
or U6281 (N_6281,N_5409,N_5017);
and U6282 (N_6282,N_5440,N_5364);
nand U6283 (N_6283,N_5330,N_5398);
and U6284 (N_6284,N_5872,N_5344);
or U6285 (N_6285,N_5277,N_5221);
nand U6286 (N_6286,N_5576,N_5049);
and U6287 (N_6287,N_5780,N_5853);
nor U6288 (N_6288,N_5496,N_5191);
and U6289 (N_6289,N_5097,N_5178);
or U6290 (N_6290,N_5947,N_5491);
nand U6291 (N_6291,N_5844,N_5702);
xnor U6292 (N_6292,N_5246,N_5396);
and U6293 (N_6293,N_5431,N_5216);
nor U6294 (N_6294,N_5142,N_5995);
xor U6295 (N_6295,N_5101,N_5783);
or U6296 (N_6296,N_5181,N_5619);
nor U6297 (N_6297,N_5028,N_5137);
or U6298 (N_6298,N_5682,N_5229);
nor U6299 (N_6299,N_5201,N_5449);
nand U6300 (N_6300,N_5341,N_5584);
or U6301 (N_6301,N_5393,N_5130);
xor U6302 (N_6302,N_5173,N_5367);
nor U6303 (N_6303,N_5993,N_5643);
nor U6304 (N_6304,N_5370,N_5545);
xnor U6305 (N_6305,N_5478,N_5803);
or U6306 (N_6306,N_5815,N_5290);
xnor U6307 (N_6307,N_5974,N_5147);
and U6308 (N_6308,N_5007,N_5129);
nand U6309 (N_6309,N_5210,N_5230);
xnor U6310 (N_6310,N_5662,N_5046);
xnor U6311 (N_6311,N_5851,N_5446);
and U6312 (N_6312,N_5726,N_5988);
nand U6313 (N_6313,N_5697,N_5411);
nor U6314 (N_6314,N_5391,N_5121);
or U6315 (N_6315,N_5673,N_5086);
nand U6316 (N_6316,N_5009,N_5272);
nor U6317 (N_6317,N_5495,N_5676);
and U6318 (N_6318,N_5601,N_5288);
nor U6319 (N_6319,N_5729,N_5144);
xor U6320 (N_6320,N_5422,N_5289);
nand U6321 (N_6321,N_5050,N_5986);
or U6322 (N_6322,N_5163,N_5824);
or U6323 (N_6323,N_5572,N_5590);
xnor U6324 (N_6324,N_5524,N_5376);
xnor U6325 (N_6325,N_5560,N_5474);
nor U6326 (N_6326,N_5348,N_5010);
or U6327 (N_6327,N_5306,N_5200);
and U6328 (N_6328,N_5323,N_5632);
xor U6329 (N_6329,N_5227,N_5146);
or U6330 (N_6330,N_5746,N_5061);
or U6331 (N_6331,N_5862,N_5869);
or U6332 (N_6332,N_5604,N_5589);
xor U6333 (N_6333,N_5549,N_5374);
nand U6334 (N_6334,N_5633,N_5107);
xnor U6335 (N_6335,N_5311,N_5024);
and U6336 (N_6336,N_5228,N_5745);
nor U6337 (N_6337,N_5801,N_5542);
and U6338 (N_6338,N_5171,N_5515);
nand U6339 (N_6339,N_5507,N_5970);
and U6340 (N_6340,N_5118,N_5438);
nand U6341 (N_6341,N_5521,N_5387);
and U6342 (N_6342,N_5255,N_5214);
and U6343 (N_6343,N_5164,N_5203);
nand U6344 (N_6344,N_5924,N_5293);
xnor U6345 (N_6345,N_5793,N_5583);
xnor U6346 (N_6346,N_5038,N_5909);
nand U6347 (N_6347,N_5703,N_5182);
and U6348 (N_6348,N_5254,N_5807);
and U6349 (N_6349,N_5208,N_5322);
nor U6350 (N_6350,N_5655,N_5897);
nor U6351 (N_6351,N_5057,N_5561);
nor U6352 (N_6352,N_5071,N_5430);
and U6353 (N_6353,N_5630,N_5532);
and U6354 (N_6354,N_5052,N_5850);
xor U6355 (N_6355,N_5263,N_5065);
nor U6356 (N_6356,N_5064,N_5954);
or U6357 (N_6357,N_5618,N_5879);
and U6358 (N_6358,N_5878,N_5035);
xor U6359 (N_6359,N_5949,N_5923);
or U6360 (N_6360,N_5605,N_5296);
or U6361 (N_6361,N_5380,N_5248);
xnor U6362 (N_6362,N_5198,N_5390);
and U6363 (N_6363,N_5912,N_5138);
or U6364 (N_6364,N_5359,N_5638);
nor U6365 (N_6365,N_5754,N_5881);
and U6366 (N_6366,N_5769,N_5694);
nor U6367 (N_6367,N_5712,N_5855);
and U6368 (N_6368,N_5800,N_5427);
and U6369 (N_6369,N_5658,N_5204);
nor U6370 (N_6370,N_5108,N_5075);
and U6371 (N_6371,N_5054,N_5172);
nand U6372 (N_6372,N_5796,N_5407);
nand U6373 (N_6373,N_5001,N_5764);
and U6374 (N_6374,N_5747,N_5093);
or U6375 (N_6375,N_5304,N_5997);
nor U6376 (N_6376,N_5439,N_5259);
xnor U6377 (N_6377,N_5260,N_5338);
nand U6378 (N_6378,N_5041,N_5294);
xnor U6379 (N_6379,N_5777,N_5252);
and U6380 (N_6380,N_5357,N_5320);
and U6381 (N_6381,N_5106,N_5811);
nor U6382 (N_6382,N_5165,N_5973);
nand U6383 (N_6383,N_5538,N_5262);
or U6384 (N_6384,N_5852,N_5155);
nand U6385 (N_6385,N_5012,N_5291);
and U6386 (N_6386,N_5444,N_5303);
nand U6387 (N_6387,N_5602,N_5463);
and U6388 (N_6388,N_5555,N_5211);
nand U6389 (N_6389,N_5158,N_5523);
or U6390 (N_6390,N_5475,N_5157);
or U6391 (N_6391,N_5641,N_5550);
nor U6392 (N_6392,N_5126,N_5950);
nand U6393 (N_6393,N_5918,N_5386);
and U6394 (N_6394,N_5805,N_5117);
or U6395 (N_6395,N_5404,N_5921);
xnor U6396 (N_6396,N_5825,N_5865);
and U6397 (N_6397,N_5343,N_5264);
and U6398 (N_6398,N_5653,N_5588);
nor U6399 (N_6399,N_5831,N_5987);
and U6400 (N_6400,N_5714,N_5767);
or U6401 (N_6401,N_5895,N_5197);
nor U6402 (N_6402,N_5345,N_5557);
nand U6403 (N_6403,N_5790,N_5067);
and U6404 (N_6404,N_5308,N_5369);
and U6405 (N_6405,N_5489,N_5511);
or U6406 (N_6406,N_5859,N_5081);
and U6407 (N_6407,N_5043,N_5938);
and U6408 (N_6408,N_5105,N_5300);
nor U6409 (N_6409,N_5456,N_5174);
nor U6410 (N_6410,N_5528,N_5654);
and U6411 (N_6411,N_5039,N_5362);
nor U6412 (N_6412,N_5609,N_5686);
and U6413 (N_6413,N_5134,N_5104);
nand U6414 (N_6414,N_5457,N_5124);
or U6415 (N_6415,N_5033,N_5656);
and U6416 (N_6416,N_5510,N_5708);
and U6417 (N_6417,N_5614,N_5240);
nor U6418 (N_6418,N_5499,N_5684);
or U6419 (N_6419,N_5727,N_5184);
nand U6420 (N_6420,N_5087,N_5883);
nand U6421 (N_6421,N_5681,N_5598);
nand U6422 (N_6422,N_5599,N_5454);
nor U6423 (N_6423,N_5828,N_5782);
nor U6424 (N_6424,N_5486,N_5072);
xor U6425 (N_6425,N_5787,N_5709);
nand U6426 (N_6426,N_5241,N_5784);
or U6427 (N_6427,N_5606,N_5123);
and U6428 (N_6428,N_5185,N_5135);
or U6429 (N_6429,N_5732,N_5152);
and U6430 (N_6430,N_5789,N_5934);
nor U6431 (N_6431,N_5593,N_5140);
nor U6432 (N_6432,N_5582,N_5132);
nand U6433 (N_6433,N_5492,N_5615);
nor U6434 (N_6434,N_5926,N_5360);
or U6435 (N_6435,N_5951,N_5472);
or U6436 (N_6436,N_5744,N_5034);
and U6437 (N_6437,N_5958,N_5331);
or U6438 (N_6438,N_5991,N_5845);
and U6439 (N_6439,N_5613,N_5120);
or U6440 (N_6440,N_5068,N_5327);
nand U6441 (N_6441,N_5570,N_5159);
nand U6442 (N_6442,N_5006,N_5635);
nor U6443 (N_6443,N_5887,N_5900);
and U6444 (N_6444,N_5760,N_5443);
nand U6445 (N_6445,N_5867,N_5624);
nor U6446 (N_6446,N_5467,N_5334);
or U6447 (N_6447,N_5136,N_5832);
nand U6448 (N_6448,N_5715,N_5269);
and U6449 (N_6449,N_5271,N_5223);
xnor U6450 (N_6450,N_5823,N_5818);
xor U6451 (N_6451,N_5610,N_5301);
or U6452 (N_6452,N_5586,N_5141);
nor U6453 (N_6453,N_5663,N_5025);
nor U6454 (N_6454,N_5274,N_5581);
xnor U6455 (N_6455,N_5128,N_5541);
nor U6456 (N_6456,N_5099,N_5781);
or U6457 (N_6457,N_5063,N_5980);
and U6458 (N_6458,N_5403,N_5077);
nor U6459 (N_6459,N_5133,N_5192);
or U6460 (N_6460,N_5649,N_5480);
and U6461 (N_6461,N_5433,N_5512);
or U6462 (N_6462,N_5169,N_5313);
nor U6463 (N_6463,N_5734,N_5412);
nand U6464 (N_6464,N_5392,N_5070);
nor U6465 (N_6465,N_5886,N_5873);
and U6466 (N_6466,N_5607,N_5817);
xor U6467 (N_6467,N_5799,N_5637);
nor U6468 (N_6468,N_5914,N_5861);
nor U6469 (N_6469,N_5186,N_5023);
or U6470 (N_6470,N_5907,N_5636);
nand U6471 (N_6471,N_5347,N_5733);
or U6472 (N_6472,N_5896,N_5032);
or U6473 (N_6473,N_5212,N_5016);
and U6474 (N_6474,N_5349,N_5617);
or U6475 (N_6475,N_5423,N_5505);
nand U6476 (N_6476,N_5838,N_5533);
nand U6477 (N_6477,N_5639,N_5770);
or U6478 (N_6478,N_5978,N_5573);
or U6479 (N_6479,N_5335,N_5766);
xnor U6480 (N_6480,N_5498,N_5441);
or U6481 (N_6481,N_5526,N_5424);
and U6482 (N_6482,N_5187,N_5716);
and U6483 (N_6483,N_5231,N_5677);
or U6484 (N_6484,N_5877,N_5930);
and U6485 (N_6485,N_5408,N_5176);
nand U6486 (N_6486,N_5477,N_5047);
nor U6487 (N_6487,N_5085,N_5415);
nand U6488 (N_6488,N_5332,N_5098);
nor U6489 (N_6489,N_5531,N_5830);
nand U6490 (N_6490,N_5595,N_5339);
or U6491 (N_6491,N_5384,N_5623);
nand U6492 (N_6492,N_5397,N_5695);
nor U6493 (N_6493,N_5564,N_5603);
xor U6494 (N_6494,N_5608,N_5405);
or U6495 (N_6495,N_5333,N_5419);
and U6496 (N_6496,N_5074,N_5484);
and U6497 (N_6497,N_5794,N_5003);
nor U6498 (N_6498,N_5428,N_5207);
and U6499 (N_6499,N_5366,N_5111);
nand U6500 (N_6500,N_5549,N_5294);
or U6501 (N_6501,N_5415,N_5899);
xnor U6502 (N_6502,N_5012,N_5142);
or U6503 (N_6503,N_5732,N_5903);
or U6504 (N_6504,N_5760,N_5111);
nand U6505 (N_6505,N_5703,N_5434);
or U6506 (N_6506,N_5453,N_5792);
xnor U6507 (N_6507,N_5481,N_5689);
nand U6508 (N_6508,N_5692,N_5561);
or U6509 (N_6509,N_5279,N_5344);
xor U6510 (N_6510,N_5652,N_5425);
xor U6511 (N_6511,N_5432,N_5571);
nor U6512 (N_6512,N_5133,N_5046);
nand U6513 (N_6513,N_5845,N_5897);
and U6514 (N_6514,N_5121,N_5607);
or U6515 (N_6515,N_5613,N_5234);
and U6516 (N_6516,N_5964,N_5602);
and U6517 (N_6517,N_5660,N_5074);
nand U6518 (N_6518,N_5805,N_5390);
nor U6519 (N_6519,N_5636,N_5022);
or U6520 (N_6520,N_5219,N_5424);
nor U6521 (N_6521,N_5470,N_5992);
or U6522 (N_6522,N_5213,N_5468);
and U6523 (N_6523,N_5053,N_5281);
and U6524 (N_6524,N_5355,N_5198);
nor U6525 (N_6525,N_5532,N_5360);
nand U6526 (N_6526,N_5276,N_5285);
and U6527 (N_6527,N_5166,N_5413);
or U6528 (N_6528,N_5878,N_5014);
xor U6529 (N_6529,N_5440,N_5481);
and U6530 (N_6530,N_5943,N_5281);
xnor U6531 (N_6531,N_5665,N_5055);
nor U6532 (N_6532,N_5586,N_5754);
and U6533 (N_6533,N_5527,N_5039);
nand U6534 (N_6534,N_5315,N_5191);
nor U6535 (N_6535,N_5174,N_5326);
and U6536 (N_6536,N_5836,N_5736);
and U6537 (N_6537,N_5239,N_5118);
and U6538 (N_6538,N_5837,N_5463);
or U6539 (N_6539,N_5610,N_5189);
or U6540 (N_6540,N_5118,N_5181);
or U6541 (N_6541,N_5723,N_5507);
and U6542 (N_6542,N_5324,N_5399);
nor U6543 (N_6543,N_5327,N_5270);
or U6544 (N_6544,N_5456,N_5688);
or U6545 (N_6545,N_5000,N_5343);
nand U6546 (N_6546,N_5308,N_5534);
nor U6547 (N_6547,N_5185,N_5959);
and U6548 (N_6548,N_5829,N_5866);
or U6549 (N_6549,N_5111,N_5850);
and U6550 (N_6550,N_5067,N_5355);
and U6551 (N_6551,N_5324,N_5920);
nor U6552 (N_6552,N_5122,N_5444);
or U6553 (N_6553,N_5399,N_5796);
or U6554 (N_6554,N_5811,N_5696);
nor U6555 (N_6555,N_5881,N_5067);
nor U6556 (N_6556,N_5972,N_5851);
and U6557 (N_6557,N_5969,N_5977);
nor U6558 (N_6558,N_5362,N_5764);
or U6559 (N_6559,N_5270,N_5710);
xor U6560 (N_6560,N_5031,N_5995);
and U6561 (N_6561,N_5414,N_5987);
xor U6562 (N_6562,N_5229,N_5350);
or U6563 (N_6563,N_5475,N_5084);
or U6564 (N_6564,N_5556,N_5511);
and U6565 (N_6565,N_5867,N_5652);
nand U6566 (N_6566,N_5200,N_5503);
xnor U6567 (N_6567,N_5343,N_5441);
and U6568 (N_6568,N_5796,N_5946);
or U6569 (N_6569,N_5043,N_5584);
nand U6570 (N_6570,N_5980,N_5416);
or U6571 (N_6571,N_5718,N_5785);
nand U6572 (N_6572,N_5515,N_5717);
nand U6573 (N_6573,N_5170,N_5918);
nand U6574 (N_6574,N_5244,N_5830);
and U6575 (N_6575,N_5321,N_5968);
nor U6576 (N_6576,N_5982,N_5675);
nand U6577 (N_6577,N_5596,N_5195);
nor U6578 (N_6578,N_5162,N_5684);
or U6579 (N_6579,N_5570,N_5139);
xor U6580 (N_6580,N_5175,N_5122);
nor U6581 (N_6581,N_5540,N_5148);
or U6582 (N_6582,N_5837,N_5499);
and U6583 (N_6583,N_5396,N_5466);
and U6584 (N_6584,N_5976,N_5182);
nor U6585 (N_6585,N_5837,N_5453);
nor U6586 (N_6586,N_5743,N_5954);
or U6587 (N_6587,N_5285,N_5506);
nor U6588 (N_6588,N_5819,N_5630);
nand U6589 (N_6589,N_5458,N_5722);
and U6590 (N_6590,N_5121,N_5124);
or U6591 (N_6591,N_5845,N_5071);
xor U6592 (N_6592,N_5055,N_5938);
nand U6593 (N_6593,N_5291,N_5055);
nand U6594 (N_6594,N_5515,N_5896);
and U6595 (N_6595,N_5901,N_5917);
xor U6596 (N_6596,N_5073,N_5046);
nor U6597 (N_6597,N_5969,N_5507);
and U6598 (N_6598,N_5770,N_5073);
and U6599 (N_6599,N_5213,N_5080);
nand U6600 (N_6600,N_5192,N_5197);
and U6601 (N_6601,N_5732,N_5199);
nor U6602 (N_6602,N_5511,N_5453);
nor U6603 (N_6603,N_5599,N_5419);
nand U6604 (N_6604,N_5154,N_5442);
or U6605 (N_6605,N_5015,N_5102);
and U6606 (N_6606,N_5646,N_5319);
nand U6607 (N_6607,N_5255,N_5232);
xor U6608 (N_6608,N_5451,N_5157);
nor U6609 (N_6609,N_5643,N_5685);
or U6610 (N_6610,N_5463,N_5938);
and U6611 (N_6611,N_5894,N_5917);
and U6612 (N_6612,N_5722,N_5019);
nand U6613 (N_6613,N_5153,N_5859);
nor U6614 (N_6614,N_5074,N_5779);
nor U6615 (N_6615,N_5990,N_5348);
nor U6616 (N_6616,N_5256,N_5880);
and U6617 (N_6617,N_5149,N_5560);
nor U6618 (N_6618,N_5744,N_5452);
nand U6619 (N_6619,N_5812,N_5256);
and U6620 (N_6620,N_5266,N_5241);
or U6621 (N_6621,N_5296,N_5386);
and U6622 (N_6622,N_5299,N_5514);
and U6623 (N_6623,N_5215,N_5513);
nand U6624 (N_6624,N_5935,N_5168);
nor U6625 (N_6625,N_5263,N_5632);
nand U6626 (N_6626,N_5817,N_5798);
nand U6627 (N_6627,N_5100,N_5212);
and U6628 (N_6628,N_5705,N_5787);
and U6629 (N_6629,N_5580,N_5889);
and U6630 (N_6630,N_5929,N_5332);
nand U6631 (N_6631,N_5283,N_5072);
nor U6632 (N_6632,N_5670,N_5284);
nor U6633 (N_6633,N_5789,N_5078);
nor U6634 (N_6634,N_5787,N_5117);
and U6635 (N_6635,N_5500,N_5268);
xor U6636 (N_6636,N_5220,N_5078);
or U6637 (N_6637,N_5267,N_5121);
xor U6638 (N_6638,N_5616,N_5770);
or U6639 (N_6639,N_5113,N_5332);
or U6640 (N_6640,N_5278,N_5190);
nor U6641 (N_6641,N_5673,N_5285);
and U6642 (N_6642,N_5346,N_5206);
and U6643 (N_6643,N_5320,N_5818);
and U6644 (N_6644,N_5107,N_5818);
xnor U6645 (N_6645,N_5256,N_5839);
or U6646 (N_6646,N_5431,N_5389);
nand U6647 (N_6647,N_5585,N_5213);
nand U6648 (N_6648,N_5862,N_5671);
nor U6649 (N_6649,N_5486,N_5580);
and U6650 (N_6650,N_5158,N_5520);
nand U6651 (N_6651,N_5402,N_5510);
nand U6652 (N_6652,N_5105,N_5065);
or U6653 (N_6653,N_5997,N_5848);
nand U6654 (N_6654,N_5787,N_5041);
or U6655 (N_6655,N_5956,N_5614);
nand U6656 (N_6656,N_5417,N_5692);
nor U6657 (N_6657,N_5827,N_5138);
nand U6658 (N_6658,N_5600,N_5997);
nand U6659 (N_6659,N_5180,N_5185);
or U6660 (N_6660,N_5771,N_5265);
and U6661 (N_6661,N_5635,N_5199);
nor U6662 (N_6662,N_5674,N_5323);
or U6663 (N_6663,N_5455,N_5966);
nand U6664 (N_6664,N_5697,N_5298);
nand U6665 (N_6665,N_5312,N_5268);
nand U6666 (N_6666,N_5697,N_5402);
nor U6667 (N_6667,N_5330,N_5251);
xor U6668 (N_6668,N_5469,N_5931);
or U6669 (N_6669,N_5884,N_5152);
and U6670 (N_6670,N_5510,N_5569);
nand U6671 (N_6671,N_5094,N_5718);
and U6672 (N_6672,N_5400,N_5231);
and U6673 (N_6673,N_5898,N_5301);
xor U6674 (N_6674,N_5916,N_5027);
or U6675 (N_6675,N_5243,N_5466);
or U6676 (N_6676,N_5301,N_5683);
and U6677 (N_6677,N_5913,N_5750);
nand U6678 (N_6678,N_5231,N_5166);
nand U6679 (N_6679,N_5561,N_5969);
nor U6680 (N_6680,N_5423,N_5981);
nor U6681 (N_6681,N_5237,N_5784);
or U6682 (N_6682,N_5166,N_5872);
nand U6683 (N_6683,N_5171,N_5152);
or U6684 (N_6684,N_5526,N_5264);
nor U6685 (N_6685,N_5394,N_5475);
nor U6686 (N_6686,N_5970,N_5245);
and U6687 (N_6687,N_5312,N_5254);
and U6688 (N_6688,N_5747,N_5244);
or U6689 (N_6689,N_5064,N_5151);
nor U6690 (N_6690,N_5330,N_5432);
nor U6691 (N_6691,N_5072,N_5583);
or U6692 (N_6692,N_5754,N_5424);
and U6693 (N_6693,N_5232,N_5776);
nor U6694 (N_6694,N_5901,N_5404);
nand U6695 (N_6695,N_5083,N_5516);
or U6696 (N_6696,N_5992,N_5320);
or U6697 (N_6697,N_5919,N_5039);
nand U6698 (N_6698,N_5806,N_5158);
or U6699 (N_6699,N_5961,N_5199);
xor U6700 (N_6700,N_5424,N_5863);
xnor U6701 (N_6701,N_5757,N_5299);
nand U6702 (N_6702,N_5334,N_5211);
or U6703 (N_6703,N_5959,N_5015);
and U6704 (N_6704,N_5249,N_5845);
and U6705 (N_6705,N_5762,N_5966);
nand U6706 (N_6706,N_5829,N_5147);
nand U6707 (N_6707,N_5166,N_5864);
and U6708 (N_6708,N_5153,N_5018);
or U6709 (N_6709,N_5430,N_5855);
nor U6710 (N_6710,N_5090,N_5621);
nor U6711 (N_6711,N_5726,N_5144);
nor U6712 (N_6712,N_5251,N_5213);
nand U6713 (N_6713,N_5891,N_5280);
or U6714 (N_6714,N_5627,N_5027);
nand U6715 (N_6715,N_5829,N_5891);
xor U6716 (N_6716,N_5142,N_5078);
and U6717 (N_6717,N_5151,N_5622);
xor U6718 (N_6718,N_5280,N_5841);
or U6719 (N_6719,N_5921,N_5768);
xnor U6720 (N_6720,N_5676,N_5936);
nor U6721 (N_6721,N_5841,N_5473);
or U6722 (N_6722,N_5273,N_5465);
or U6723 (N_6723,N_5163,N_5182);
xnor U6724 (N_6724,N_5570,N_5683);
nand U6725 (N_6725,N_5503,N_5405);
xor U6726 (N_6726,N_5275,N_5028);
or U6727 (N_6727,N_5085,N_5552);
nor U6728 (N_6728,N_5835,N_5936);
nor U6729 (N_6729,N_5974,N_5702);
or U6730 (N_6730,N_5417,N_5044);
nor U6731 (N_6731,N_5333,N_5283);
and U6732 (N_6732,N_5317,N_5328);
xor U6733 (N_6733,N_5142,N_5784);
and U6734 (N_6734,N_5985,N_5186);
and U6735 (N_6735,N_5782,N_5379);
nor U6736 (N_6736,N_5065,N_5546);
and U6737 (N_6737,N_5793,N_5417);
and U6738 (N_6738,N_5265,N_5520);
or U6739 (N_6739,N_5729,N_5685);
nor U6740 (N_6740,N_5124,N_5551);
and U6741 (N_6741,N_5800,N_5460);
or U6742 (N_6742,N_5794,N_5031);
xor U6743 (N_6743,N_5283,N_5530);
nor U6744 (N_6744,N_5645,N_5959);
or U6745 (N_6745,N_5916,N_5053);
nand U6746 (N_6746,N_5527,N_5648);
or U6747 (N_6747,N_5010,N_5847);
nand U6748 (N_6748,N_5946,N_5513);
nor U6749 (N_6749,N_5478,N_5071);
and U6750 (N_6750,N_5632,N_5383);
or U6751 (N_6751,N_5013,N_5528);
nor U6752 (N_6752,N_5082,N_5022);
nand U6753 (N_6753,N_5220,N_5821);
nor U6754 (N_6754,N_5383,N_5058);
and U6755 (N_6755,N_5426,N_5715);
nor U6756 (N_6756,N_5570,N_5393);
and U6757 (N_6757,N_5067,N_5066);
nand U6758 (N_6758,N_5185,N_5155);
xor U6759 (N_6759,N_5362,N_5256);
or U6760 (N_6760,N_5655,N_5771);
nand U6761 (N_6761,N_5783,N_5343);
and U6762 (N_6762,N_5248,N_5865);
or U6763 (N_6763,N_5381,N_5293);
or U6764 (N_6764,N_5854,N_5210);
or U6765 (N_6765,N_5667,N_5063);
nand U6766 (N_6766,N_5156,N_5108);
nor U6767 (N_6767,N_5792,N_5986);
nand U6768 (N_6768,N_5051,N_5204);
nand U6769 (N_6769,N_5210,N_5004);
and U6770 (N_6770,N_5013,N_5974);
nor U6771 (N_6771,N_5692,N_5544);
nand U6772 (N_6772,N_5764,N_5394);
or U6773 (N_6773,N_5526,N_5693);
nor U6774 (N_6774,N_5689,N_5059);
nand U6775 (N_6775,N_5756,N_5378);
nor U6776 (N_6776,N_5482,N_5595);
or U6777 (N_6777,N_5475,N_5150);
nand U6778 (N_6778,N_5341,N_5774);
and U6779 (N_6779,N_5873,N_5398);
or U6780 (N_6780,N_5605,N_5436);
or U6781 (N_6781,N_5460,N_5577);
and U6782 (N_6782,N_5552,N_5222);
xnor U6783 (N_6783,N_5587,N_5622);
and U6784 (N_6784,N_5651,N_5716);
nor U6785 (N_6785,N_5858,N_5514);
nor U6786 (N_6786,N_5423,N_5732);
xnor U6787 (N_6787,N_5497,N_5483);
or U6788 (N_6788,N_5328,N_5680);
nor U6789 (N_6789,N_5400,N_5584);
or U6790 (N_6790,N_5313,N_5711);
or U6791 (N_6791,N_5312,N_5026);
nor U6792 (N_6792,N_5570,N_5826);
and U6793 (N_6793,N_5639,N_5874);
nor U6794 (N_6794,N_5146,N_5997);
nor U6795 (N_6795,N_5845,N_5680);
xor U6796 (N_6796,N_5075,N_5404);
nor U6797 (N_6797,N_5812,N_5429);
nand U6798 (N_6798,N_5113,N_5659);
and U6799 (N_6799,N_5349,N_5364);
xor U6800 (N_6800,N_5571,N_5345);
or U6801 (N_6801,N_5218,N_5423);
or U6802 (N_6802,N_5758,N_5423);
nand U6803 (N_6803,N_5583,N_5470);
and U6804 (N_6804,N_5031,N_5617);
or U6805 (N_6805,N_5888,N_5035);
or U6806 (N_6806,N_5718,N_5786);
or U6807 (N_6807,N_5995,N_5344);
or U6808 (N_6808,N_5972,N_5347);
and U6809 (N_6809,N_5890,N_5309);
nor U6810 (N_6810,N_5082,N_5969);
xnor U6811 (N_6811,N_5551,N_5807);
and U6812 (N_6812,N_5861,N_5296);
and U6813 (N_6813,N_5597,N_5767);
or U6814 (N_6814,N_5173,N_5954);
and U6815 (N_6815,N_5501,N_5189);
nor U6816 (N_6816,N_5427,N_5994);
and U6817 (N_6817,N_5215,N_5414);
nand U6818 (N_6818,N_5721,N_5307);
xor U6819 (N_6819,N_5093,N_5278);
nand U6820 (N_6820,N_5288,N_5274);
nor U6821 (N_6821,N_5842,N_5005);
nor U6822 (N_6822,N_5271,N_5378);
or U6823 (N_6823,N_5532,N_5391);
and U6824 (N_6824,N_5890,N_5623);
nor U6825 (N_6825,N_5854,N_5472);
xnor U6826 (N_6826,N_5440,N_5963);
or U6827 (N_6827,N_5254,N_5001);
nand U6828 (N_6828,N_5869,N_5271);
nand U6829 (N_6829,N_5598,N_5959);
nand U6830 (N_6830,N_5058,N_5143);
xnor U6831 (N_6831,N_5309,N_5595);
or U6832 (N_6832,N_5024,N_5190);
xor U6833 (N_6833,N_5780,N_5745);
nor U6834 (N_6834,N_5042,N_5543);
or U6835 (N_6835,N_5612,N_5020);
or U6836 (N_6836,N_5419,N_5617);
nor U6837 (N_6837,N_5933,N_5962);
xor U6838 (N_6838,N_5060,N_5375);
nand U6839 (N_6839,N_5032,N_5858);
nand U6840 (N_6840,N_5101,N_5828);
and U6841 (N_6841,N_5641,N_5003);
and U6842 (N_6842,N_5182,N_5075);
nor U6843 (N_6843,N_5565,N_5755);
or U6844 (N_6844,N_5401,N_5996);
nor U6845 (N_6845,N_5103,N_5716);
nand U6846 (N_6846,N_5928,N_5258);
or U6847 (N_6847,N_5186,N_5506);
nor U6848 (N_6848,N_5159,N_5225);
nand U6849 (N_6849,N_5252,N_5503);
or U6850 (N_6850,N_5152,N_5454);
and U6851 (N_6851,N_5915,N_5250);
nand U6852 (N_6852,N_5714,N_5189);
nor U6853 (N_6853,N_5272,N_5443);
nor U6854 (N_6854,N_5401,N_5502);
and U6855 (N_6855,N_5813,N_5413);
nor U6856 (N_6856,N_5487,N_5964);
and U6857 (N_6857,N_5085,N_5208);
and U6858 (N_6858,N_5231,N_5317);
or U6859 (N_6859,N_5118,N_5123);
and U6860 (N_6860,N_5498,N_5830);
and U6861 (N_6861,N_5396,N_5509);
or U6862 (N_6862,N_5212,N_5666);
nand U6863 (N_6863,N_5618,N_5829);
and U6864 (N_6864,N_5765,N_5895);
nor U6865 (N_6865,N_5520,N_5305);
xnor U6866 (N_6866,N_5041,N_5815);
nor U6867 (N_6867,N_5127,N_5148);
and U6868 (N_6868,N_5320,N_5964);
nor U6869 (N_6869,N_5836,N_5866);
and U6870 (N_6870,N_5989,N_5906);
nor U6871 (N_6871,N_5472,N_5243);
xor U6872 (N_6872,N_5236,N_5856);
nor U6873 (N_6873,N_5377,N_5123);
and U6874 (N_6874,N_5379,N_5164);
nor U6875 (N_6875,N_5596,N_5000);
or U6876 (N_6876,N_5721,N_5793);
nand U6877 (N_6877,N_5760,N_5385);
nor U6878 (N_6878,N_5217,N_5265);
and U6879 (N_6879,N_5968,N_5697);
nand U6880 (N_6880,N_5831,N_5733);
nand U6881 (N_6881,N_5270,N_5299);
and U6882 (N_6882,N_5520,N_5287);
nor U6883 (N_6883,N_5343,N_5567);
and U6884 (N_6884,N_5257,N_5350);
nor U6885 (N_6885,N_5068,N_5677);
and U6886 (N_6886,N_5163,N_5097);
or U6887 (N_6887,N_5249,N_5239);
nand U6888 (N_6888,N_5140,N_5056);
nor U6889 (N_6889,N_5699,N_5497);
nor U6890 (N_6890,N_5687,N_5039);
or U6891 (N_6891,N_5285,N_5147);
xnor U6892 (N_6892,N_5926,N_5325);
nor U6893 (N_6893,N_5976,N_5536);
and U6894 (N_6894,N_5724,N_5412);
nand U6895 (N_6895,N_5813,N_5181);
nand U6896 (N_6896,N_5138,N_5610);
or U6897 (N_6897,N_5849,N_5331);
nor U6898 (N_6898,N_5819,N_5254);
nor U6899 (N_6899,N_5136,N_5469);
and U6900 (N_6900,N_5306,N_5148);
nor U6901 (N_6901,N_5561,N_5160);
xor U6902 (N_6902,N_5655,N_5105);
and U6903 (N_6903,N_5584,N_5663);
and U6904 (N_6904,N_5136,N_5165);
nor U6905 (N_6905,N_5011,N_5191);
and U6906 (N_6906,N_5065,N_5948);
nor U6907 (N_6907,N_5235,N_5446);
and U6908 (N_6908,N_5438,N_5705);
nor U6909 (N_6909,N_5341,N_5191);
or U6910 (N_6910,N_5576,N_5660);
xnor U6911 (N_6911,N_5020,N_5251);
or U6912 (N_6912,N_5525,N_5384);
and U6913 (N_6913,N_5072,N_5239);
nand U6914 (N_6914,N_5357,N_5438);
and U6915 (N_6915,N_5566,N_5858);
nor U6916 (N_6916,N_5548,N_5462);
nor U6917 (N_6917,N_5575,N_5826);
or U6918 (N_6918,N_5445,N_5713);
nand U6919 (N_6919,N_5720,N_5230);
xor U6920 (N_6920,N_5897,N_5721);
nor U6921 (N_6921,N_5987,N_5470);
nor U6922 (N_6922,N_5380,N_5268);
nand U6923 (N_6923,N_5446,N_5530);
nand U6924 (N_6924,N_5748,N_5775);
nand U6925 (N_6925,N_5338,N_5169);
or U6926 (N_6926,N_5249,N_5252);
nand U6927 (N_6927,N_5101,N_5258);
nor U6928 (N_6928,N_5849,N_5169);
and U6929 (N_6929,N_5800,N_5522);
nand U6930 (N_6930,N_5798,N_5010);
nor U6931 (N_6931,N_5830,N_5312);
nor U6932 (N_6932,N_5445,N_5086);
and U6933 (N_6933,N_5819,N_5565);
nor U6934 (N_6934,N_5169,N_5828);
and U6935 (N_6935,N_5188,N_5833);
and U6936 (N_6936,N_5361,N_5423);
or U6937 (N_6937,N_5605,N_5760);
and U6938 (N_6938,N_5005,N_5246);
and U6939 (N_6939,N_5670,N_5923);
nor U6940 (N_6940,N_5258,N_5384);
nor U6941 (N_6941,N_5192,N_5935);
nand U6942 (N_6942,N_5462,N_5134);
or U6943 (N_6943,N_5473,N_5905);
nor U6944 (N_6944,N_5116,N_5995);
and U6945 (N_6945,N_5224,N_5289);
or U6946 (N_6946,N_5380,N_5454);
nand U6947 (N_6947,N_5742,N_5385);
nor U6948 (N_6948,N_5279,N_5990);
nand U6949 (N_6949,N_5648,N_5209);
and U6950 (N_6950,N_5264,N_5629);
xnor U6951 (N_6951,N_5849,N_5673);
and U6952 (N_6952,N_5209,N_5730);
or U6953 (N_6953,N_5264,N_5506);
xor U6954 (N_6954,N_5160,N_5757);
and U6955 (N_6955,N_5072,N_5393);
nand U6956 (N_6956,N_5173,N_5175);
nand U6957 (N_6957,N_5293,N_5979);
nor U6958 (N_6958,N_5908,N_5389);
nor U6959 (N_6959,N_5693,N_5212);
nand U6960 (N_6960,N_5711,N_5720);
and U6961 (N_6961,N_5502,N_5799);
nand U6962 (N_6962,N_5819,N_5308);
nor U6963 (N_6963,N_5831,N_5250);
or U6964 (N_6964,N_5298,N_5229);
or U6965 (N_6965,N_5542,N_5669);
nand U6966 (N_6966,N_5126,N_5807);
nand U6967 (N_6967,N_5284,N_5337);
nor U6968 (N_6968,N_5948,N_5748);
nor U6969 (N_6969,N_5241,N_5907);
nand U6970 (N_6970,N_5640,N_5952);
xor U6971 (N_6971,N_5760,N_5705);
nand U6972 (N_6972,N_5628,N_5532);
and U6973 (N_6973,N_5514,N_5700);
nand U6974 (N_6974,N_5049,N_5994);
nor U6975 (N_6975,N_5800,N_5030);
or U6976 (N_6976,N_5372,N_5230);
and U6977 (N_6977,N_5825,N_5623);
nand U6978 (N_6978,N_5254,N_5082);
nand U6979 (N_6979,N_5358,N_5413);
nor U6980 (N_6980,N_5817,N_5633);
nor U6981 (N_6981,N_5341,N_5194);
or U6982 (N_6982,N_5254,N_5747);
nor U6983 (N_6983,N_5920,N_5530);
nand U6984 (N_6984,N_5252,N_5977);
or U6985 (N_6985,N_5637,N_5706);
or U6986 (N_6986,N_5944,N_5515);
nand U6987 (N_6987,N_5484,N_5036);
and U6988 (N_6988,N_5693,N_5427);
or U6989 (N_6989,N_5113,N_5469);
or U6990 (N_6990,N_5889,N_5372);
nand U6991 (N_6991,N_5177,N_5380);
or U6992 (N_6992,N_5648,N_5759);
xnor U6993 (N_6993,N_5149,N_5077);
or U6994 (N_6994,N_5394,N_5206);
nor U6995 (N_6995,N_5093,N_5959);
nand U6996 (N_6996,N_5394,N_5068);
nand U6997 (N_6997,N_5005,N_5685);
and U6998 (N_6998,N_5816,N_5129);
and U6999 (N_6999,N_5759,N_5559);
and U7000 (N_7000,N_6597,N_6606);
and U7001 (N_7001,N_6442,N_6813);
or U7002 (N_7002,N_6109,N_6629);
and U7003 (N_7003,N_6080,N_6217);
nor U7004 (N_7004,N_6904,N_6415);
or U7005 (N_7005,N_6522,N_6538);
nand U7006 (N_7006,N_6725,N_6095);
nand U7007 (N_7007,N_6701,N_6125);
nor U7008 (N_7008,N_6089,N_6698);
nand U7009 (N_7009,N_6667,N_6285);
xor U7010 (N_7010,N_6842,N_6039);
and U7011 (N_7011,N_6818,N_6118);
nand U7012 (N_7012,N_6933,N_6705);
or U7013 (N_7013,N_6047,N_6750);
and U7014 (N_7014,N_6954,N_6059);
and U7015 (N_7015,N_6846,N_6441);
nand U7016 (N_7016,N_6308,N_6588);
and U7017 (N_7017,N_6645,N_6835);
nor U7018 (N_7018,N_6638,N_6689);
and U7019 (N_7019,N_6578,N_6609);
or U7020 (N_7020,N_6897,N_6599);
nor U7021 (N_7021,N_6706,N_6622);
xnor U7022 (N_7022,N_6240,N_6476);
nor U7023 (N_7023,N_6860,N_6583);
nor U7024 (N_7024,N_6016,N_6045);
or U7025 (N_7025,N_6070,N_6389);
nand U7026 (N_7026,N_6970,N_6124);
and U7027 (N_7027,N_6021,N_6873);
nand U7028 (N_7028,N_6322,N_6466);
and U7029 (N_7029,N_6816,N_6778);
xor U7030 (N_7030,N_6349,N_6533);
nor U7031 (N_7031,N_6026,N_6603);
or U7032 (N_7032,N_6277,N_6675);
nand U7033 (N_7033,N_6791,N_6140);
nand U7034 (N_7034,N_6458,N_6516);
nand U7035 (N_7035,N_6265,N_6719);
and U7036 (N_7036,N_6865,N_6207);
nor U7037 (N_7037,N_6450,N_6529);
and U7038 (N_7038,N_6895,N_6808);
or U7039 (N_7039,N_6112,N_6024);
nor U7040 (N_7040,N_6684,N_6562);
or U7041 (N_7041,N_6327,N_6312);
and U7042 (N_7042,N_6162,N_6823);
and U7043 (N_7043,N_6081,N_6608);
and U7044 (N_7044,N_6158,N_6448);
xnor U7045 (N_7045,N_6592,N_6113);
and U7046 (N_7046,N_6116,N_6214);
nand U7047 (N_7047,N_6446,N_6774);
and U7048 (N_7048,N_6014,N_6971);
nand U7049 (N_7049,N_6484,N_6145);
and U7050 (N_7050,N_6500,N_6812);
nor U7051 (N_7051,N_6878,N_6176);
or U7052 (N_7052,N_6917,N_6224);
nor U7053 (N_7053,N_6934,N_6932);
nor U7054 (N_7054,N_6163,N_6786);
and U7055 (N_7055,N_6135,N_6286);
nor U7056 (N_7056,N_6883,N_6067);
and U7057 (N_7057,N_6715,N_6863);
or U7058 (N_7058,N_6087,N_6427);
or U7059 (N_7059,N_6682,N_6000);
xor U7060 (N_7060,N_6197,N_6749);
nand U7061 (N_7061,N_6663,N_6837);
nand U7062 (N_7062,N_6394,N_6198);
xor U7063 (N_7063,N_6807,N_6976);
nor U7064 (N_7064,N_6685,N_6790);
and U7065 (N_7065,N_6637,N_6077);
xor U7066 (N_7066,N_6230,N_6041);
or U7067 (N_7067,N_6734,N_6150);
and U7068 (N_7068,N_6797,N_6004);
and U7069 (N_7069,N_6102,N_6413);
xor U7070 (N_7070,N_6074,N_6297);
nand U7071 (N_7071,N_6462,N_6439);
nor U7072 (N_7072,N_6517,N_6788);
nor U7073 (N_7073,N_6683,N_6962);
or U7074 (N_7074,N_6806,N_6338);
nor U7075 (N_7075,N_6209,N_6890);
or U7076 (N_7076,N_6872,N_6433);
and U7077 (N_7077,N_6619,N_6810);
or U7078 (N_7078,N_6346,N_6747);
or U7079 (N_7079,N_6287,N_6704);
nor U7080 (N_7080,N_6770,N_6351);
or U7081 (N_7081,N_6121,N_6900);
or U7082 (N_7082,N_6753,N_6334);
or U7083 (N_7083,N_6025,N_6249);
nor U7084 (N_7084,N_6258,N_6677);
nand U7085 (N_7085,N_6553,N_6919);
nand U7086 (N_7086,N_6844,N_6984);
and U7087 (N_7087,N_6115,N_6979);
nand U7088 (N_7088,N_6022,N_6306);
and U7089 (N_7089,N_6365,N_6231);
xor U7090 (N_7090,N_6160,N_6511);
nand U7091 (N_7091,N_6172,N_6615);
and U7092 (N_7092,N_6856,N_6502);
nor U7093 (N_7093,N_6709,N_6229);
nand U7094 (N_7094,N_6730,N_6443);
or U7095 (N_7095,N_6552,N_6395);
nor U7096 (N_7096,N_6050,N_6953);
nand U7097 (N_7097,N_6591,N_6726);
nor U7098 (N_7098,N_6916,N_6589);
and U7099 (N_7099,N_6999,N_6069);
nand U7100 (N_7100,N_6417,N_6513);
and U7101 (N_7101,N_6772,N_6487);
and U7102 (N_7102,N_6027,N_6071);
xnor U7103 (N_7103,N_6370,N_6617);
and U7104 (N_7104,N_6988,N_6002);
nor U7105 (N_7105,N_6980,N_6590);
nand U7106 (N_7106,N_6064,N_6721);
nor U7107 (N_7107,N_6802,N_6536);
nand U7108 (N_7108,N_6870,N_6180);
nor U7109 (N_7109,N_6983,N_6927);
or U7110 (N_7110,N_6570,N_6489);
xnor U7111 (N_7111,N_6822,N_6323);
nor U7112 (N_7112,N_6783,N_6042);
nor U7113 (N_7113,N_6898,N_6833);
xor U7114 (N_7114,N_6903,N_6992);
xnor U7115 (N_7115,N_6029,N_6139);
and U7116 (N_7116,N_6151,N_6354);
nand U7117 (N_7117,N_6142,N_6482);
or U7118 (N_7118,N_6357,N_6880);
and U7119 (N_7119,N_6935,N_6119);
xnor U7120 (N_7120,N_6132,N_6248);
or U7121 (N_7121,N_6094,N_6657);
nand U7122 (N_7122,N_6781,N_6820);
nand U7123 (N_7123,N_6393,N_6170);
nor U7124 (N_7124,N_6751,N_6134);
nand U7125 (N_7125,N_6961,N_6038);
nand U7126 (N_7126,N_6337,N_6366);
and U7127 (N_7127,N_6696,N_6741);
or U7128 (N_7128,N_6396,N_6771);
and U7129 (N_7129,N_6573,N_6264);
xnor U7130 (N_7130,N_6969,N_6879);
or U7131 (N_7131,N_6843,N_6141);
or U7132 (N_7132,N_6815,N_6035);
nor U7133 (N_7133,N_6133,N_6550);
xor U7134 (N_7134,N_6196,N_6792);
or U7135 (N_7135,N_6864,N_6990);
nor U7136 (N_7136,N_6716,N_6665);
nor U7137 (N_7137,N_6329,N_6031);
nand U7138 (N_7138,N_6210,N_6686);
or U7139 (N_7139,N_6510,N_6801);
nand U7140 (N_7140,N_6278,N_6326);
xor U7141 (N_7141,N_6593,N_6471);
xor U7142 (N_7142,N_6130,N_6015);
nand U7143 (N_7143,N_6244,N_6567);
nor U7144 (N_7144,N_6032,N_6204);
nor U7145 (N_7145,N_6496,N_6332);
nand U7146 (N_7146,N_6459,N_6956);
or U7147 (N_7147,N_6656,N_6646);
nand U7148 (N_7148,N_6347,N_6085);
and U7149 (N_7149,N_6915,N_6161);
xor U7150 (N_7150,N_6653,N_6554);
xor U7151 (N_7151,N_6019,N_6273);
and U7152 (N_7152,N_6493,N_6710);
and U7153 (N_7153,N_6524,N_6044);
xor U7154 (N_7154,N_6681,N_6950);
and U7155 (N_7155,N_6449,N_6551);
xor U7156 (N_7156,N_6690,N_6416);
nand U7157 (N_7157,N_6598,N_6614);
nand U7158 (N_7158,N_6455,N_6159);
nand U7159 (N_7159,N_6626,N_6829);
or U7160 (N_7160,N_6260,N_6404);
nor U7161 (N_7161,N_6795,N_6520);
nor U7162 (N_7162,N_6558,N_6110);
and U7163 (N_7163,N_6886,N_6485);
nor U7164 (N_7164,N_6147,N_6291);
nor U7165 (N_7165,N_6222,N_6964);
xnor U7166 (N_7166,N_6530,N_6671);
and U7167 (N_7167,N_6007,N_6930);
or U7168 (N_7168,N_6876,N_6758);
xor U7169 (N_7169,N_6831,N_6321);
or U7170 (N_7170,N_6505,N_6361);
and U7171 (N_7171,N_6635,N_6952);
and U7172 (N_7172,N_6202,N_6669);
and U7173 (N_7173,N_6840,N_6921);
xor U7174 (N_7174,N_6695,N_6862);
nor U7175 (N_7175,N_6699,N_6083);
xor U7176 (N_7176,N_6242,N_6371);
nand U7177 (N_7177,N_6168,N_6114);
or U7178 (N_7178,N_6392,N_6281);
nand U7179 (N_7179,N_6090,N_6785);
nand U7180 (N_7180,N_6798,N_6046);
or U7181 (N_7181,N_6528,N_6020);
nand U7182 (N_7182,N_6908,N_6169);
nand U7183 (N_7183,N_6092,N_6010);
and U7184 (N_7184,N_6804,N_6624);
or U7185 (N_7185,N_6850,N_6457);
nor U7186 (N_7186,N_6634,N_6834);
and U7187 (N_7187,N_6303,N_6532);
nor U7188 (N_7188,N_6430,N_6909);
nor U7189 (N_7189,N_6282,N_6664);
and U7190 (N_7190,N_6407,N_6099);
or U7191 (N_7191,N_6912,N_6193);
nor U7192 (N_7192,N_6208,N_6581);
nor U7193 (N_7193,N_6494,N_6256);
nor U7194 (N_7194,N_6474,N_6707);
and U7195 (N_7195,N_6399,N_6991);
and U7196 (N_7196,N_6154,N_6410);
xor U7197 (N_7197,N_6541,N_6146);
or U7198 (N_7198,N_6166,N_6429);
nor U7199 (N_7199,N_6727,N_6018);
and U7200 (N_7200,N_6661,N_6993);
xor U7201 (N_7201,N_6218,N_6955);
nor U7202 (N_7202,N_6216,N_6377);
or U7203 (N_7203,N_6509,N_6672);
nor U7204 (N_7204,N_6495,N_6143);
nor U7205 (N_7205,N_6678,N_6717);
or U7206 (N_7206,N_6001,N_6654);
and U7207 (N_7207,N_6560,N_6960);
and U7208 (N_7208,N_6649,N_6518);
nor U7209 (N_7209,N_6616,N_6913);
and U7210 (N_7210,N_6737,N_6828);
nand U7211 (N_7211,N_6742,N_6212);
or U7212 (N_7212,N_6565,N_6131);
nand U7213 (N_7213,N_6011,N_6333);
or U7214 (N_7214,N_6033,N_6793);
nand U7215 (N_7215,N_6756,N_6313);
and U7216 (N_7216,N_6219,N_6129);
xnor U7217 (N_7217,N_6561,N_6623);
nor U7218 (N_7218,N_6799,N_6227);
or U7219 (N_7219,N_6939,N_6058);
and U7220 (N_7220,N_6680,N_6650);
or U7221 (N_7221,N_6779,N_6259);
nand U7222 (N_7222,N_6963,N_6182);
and U7223 (N_7223,N_6787,N_6486);
nand U7224 (N_7224,N_6926,N_6745);
nor U7225 (N_7225,N_6296,N_6073);
nor U7226 (N_7226,N_6643,N_6720);
or U7227 (N_7227,N_6279,N_6838);
or U7228 (N_7228,N_6435,N_6702);
or U7229 (N_7229,N_6907,N_6580);
nand U7230 (N_7230,N_6272,N_6107);
and U7231 (N_7231,N_6929,N_6868);
or U7232 (N_7232,N_6901,N_6363);
or U7233 (N_7233,N_6780,N_6187);
and U7234 (N_7234,N_6171,N_6456);
nor U7235 (N_7235,N_6402,N_6884);
nand U7236 (N_7236,N_6968,N_6275);
and U7237 (N_7237,N_6009,N_6658);
nor U7238 (N_7238,N_6061,N_6488);
and U7239 (N_7239,N_6854,N_6848);
and U7240 (N_7240,N_6521,N_6630);
xor U7241 (N_7241,N_6388,N_6445);
and U7242 (N_7242,N_6703,N_6483);
nand U7243 (N_7243,N_6362,N_6691);
and U7244 (N_7244,N_6899,N_6226);
and U7245 (N_7245,N_6996,N_6319);
and U7246 (N_7246,N_6276,N_6299);
xnor U7247 (N_7247,N_6465,N_6847);
and U7248 (N_7248,N_6266,N_6568);
nor U7249 (N_7249,N_6738,N_6403);
and U7250 (N_7250,N_6576,N_6364);
nor U7251 (N_7251,N_6386,N_6490);
nand U7252 (N_7252,N_6540,N_6111);
nand U7253 (N_7253,N_6397,N_6128);
nor U7254 (N_7254,N_6673,N_6440);
nor U7255 (N_7255,N_6767,N_6243);
nor U7256 (N_7256,N_6674,N_6173);
or U7257 (N_7257,N_6352,N_6460);
nor U7258 (N_7258,N_6559,N_6777);
and U7259 (N_7259,N_6755,N_6937);
and U7260 (N_7260,N_6692,N_6421);
xor U7261 (N_7261,N_6238,N_6017);
or U7262 (N_7262,N_6262,N_6414);
nor U7263 (N_7263,N_6424,N_6350);
nand U7264 (N_7264,N_6066,N_6481);
and U7265 (N_7265,N_6028,N_6431);
xnor U7266 (N_7266,N_6632,N_6263);
nor U7267 (N_7267,N_6467,N_6304);
and U7268 (N_7268,N_6894,N_6451);
or U7269 (N_7269,N_6255,N_6651);
nor U7270 (N_7270,N_6866,N_6062);
or U7271 (N_7271,N_6875,N_6406);
and U7272 (N_7272,N_6881,N_6931);
nand U7273 (N_7273,N_6784,N_6295);
and U7274 (N_7274,N_6858,N_6251);
nand U7275 (N_7275,N_6924,N_6454);
xor U7276 (N_7276,N_6311,N_6628);
nand U7277 (N_7277,N_6340,N_6049);
and U7278 (N_7278,N_6300,N_6839);
or U7279 (N_7279,N_6030,N_6174);
nor U7280 (N_7280,N_6736,N_6076);
xor U7281 (N_7281,N_6579,N_6379);
nor U7282 (N_7282,N_6827,N_6461);
nor U7283 (N_7283,N_6891,N_6239);
or U7284 (N_7284,N_6607,N_6499);
and U7285 (N_7285,N_6809,N_6535);
xor U7286 (N_7286,N_6766,N_6475);
nand U7287 (N_7287,N_6966,N_6679);
nand U7288 (N_7288,N_6012,N_6195);
nor U7289 (N_7289,N_6213,N_6283);
or U7290 (N_7290,N_6054,N_6288);
xnor U7291 (N_7291,N_6572,N_6662);
and U7292 (N_7292,N_6434,N_6225);
xnor U7293 (N_7293,N_6501,N_6743);
or U7294 (N_7294,N_6527,N_6359);
and U7295 (N_7295,N_6605,N_6398);
nand U7296 (N_7296,N_6641,N_6382);
xor U7297 (N_7297,N_6192,N_6302);
xor U7298 (N_7298,N_6353,N_6892);
and U7299 (N_7299,N_6339,N_6164);
xnor U7300 (N_7300,N_6307,N_6611);
or U7301 (N_7301,N_6688,N_6660);
and U7302 (N_7302,N_6639,N_6335);
nand U7303 (N_7303,N_6108,N_6188);
or U7304 (N_7304,N_6068,N_6504);
and U7305 (N_7305,N_6343,N_6411);
nor U7306 (N_7306,N_6888,N_6497);
xor U7307 (N_7307,N_6355,N_6419);
nand U7308 (N_7308,N_6436,N_6995);
nor U7309 (N_7309,N_6051,N_6604);
or U7310 (N_7310,N_6267,N_6974);
nand U7311 (N_7311,N_6760,N_6585);
or U7312 (N_7312,N_6345,N_6789);
xor U7313 (N_7313,N_6472,N_6563);
nor U7314 (N_7314,N_6280,N_6373);
or U7315 (N_7315,N_6923,N_6542);
or U7316 (N_7316,N_6910,N_6728);
nor U7317 (N_7317,N_6391,N_6384);
and U7318 (N_7318,N_6712,N_6882);
and U7319 (N_7319,N_6423,N_6261);
nand U7320 (N_7320,N_6194,N_6814);
or U7321 (N_7321,N_6694,N_6556);
or U7322 (N_7322,N_6473,N_6056);
xor U7323 (N_7323,N_6776,N_6006);
or U7324 (N_7324,N_6444,N_6564);
nand U7325 (N_7325,N_6714,N_6422);
xor U7326 (N_7326,N_6317,N_6203);
nand U7327 (N_7327,N_6228,N_6998);
xnor U7328 (N_7328,N_6945,N_6079);
nor U7329 (N_7329,N_6724,N_6739);
or U7330 (N_7330,N_6763,N_6469);
xor U7331 (N_7331,N_6997,N_6084);
and U7332 (N_7332,N_6948,N_6127);
nor U7333 (N_7333,N_6468,N_6137);
and U7334 (N_7334,N_6796,N_6148);
and U7335 (N_7335,N_6418,N_6246);
nand U7336 (N_7336,N_6136,N_6036);
nand U7337 (N_7337,N_6331,N_6156);
nand U7338 (N_7338,N_6902,N_6986);
and U7339 (N_7339,N_6744,N_6367);
and U7340 (N_7340,N_6254,N_6477);
nor U7341 (N_7341,N_6060,N_6922);
or U7342 (N_7342,N_6794,N_6234);
nand U7343 (N_7343,N_6905,N_6775);
nor U7344 (N_7344,N_6896,N_6186);
nor U7345 (N_7345,N_6072,N_6093);
xnor U7346 (N_7346,N_6723,N_6268);
nor U7347 (N_7347,N_6342,N_6078);
nor U7348 (N_7348,N_6601,N_6048);
nand U7349 (N_7349,N_6514,N_6479);
or U7350 (N_7350,N_6096,N_6324);
nand U7351 (N_7351,N_6874,N_6817);
nor U7352 (N_7352,N_6571,N_6023);
or U7353 (N_7353,N_6943,N_6985);
and U7354 (N_7354,N_6401,N_6356);
nand U7355 (N_7355,N_6757,N_6523);
and U7356 (N_7356,N_6091,N_6700);
and U7357 (N_7357,N_6369,N_6941);
xnor U7358 (N_7358,N_6232,N_6236);
nor U7359 (N_7359,N_6857,N_6117);
nor U7360 (N_7360,N_6100,N_6223);
and U7361 (N_7361,N_6566,N_6625);
nor U7362 (N_7362,N_6869,N_6426);
nor U7363 (N_7363,N_6765,N_6718);
xor U7364 (N_7364,N_6183,N_6453);
nand U7365 (N_7365,N_6034,N_6512);
nor U7366 (N_7366,N_6711,N_6729);
nor U7367 (N_7367,N_6408,N_6185);
xor U7368 (N_7368,N_6503,N_6138);
or U7369 (N_7369,N_6480,N_6447);
nand U7370 (N_7370,N_6959,N_6088);
xor U7371 (N_7371,N_6586,N_6320);
and U7372 (N_7372,N_6199,N_6867);
nor U7373 (N_7373,N_6206,N_6432);
nand U7374 (N_7374,N_6086,N_6305);
nor U7375 (N_7375,N_6005,N_6537);
nand U7376 (N_7376,N_6746,N_6252);
nand U7377 (N_7377,N_6636,N_6201);
and U7378 (N_7378,N_6438,N_6506);
and U7379 (N_7379,N_6211,N_6697);
nand U7380 (N_7380,N_6105,N_6544);
xnor U7381 (N_7381,N_6235,N_6972);
nand U7382 (N_7382,N_6942,N_6250);
or U7383 (N_7383,N_6861,N_6768);
nor U7384 (N_7384,N_6314,N_6097);
and U7385 (N_7385,N_6824,N_6341);
nand U7386 (N_7386,N_6761,N_6740);
xor U7387 (N_7387,N_6152,N_6547);
nor U7388 (N_7388,N_6053,N_6515);
nand U7389 (N_7389,N_6855,N_6676);
xor U7390 (N_7390,N_6375,N_6368);
or U7391 (N_7391,N_6437,N_6759);
nor U7392 (N_7392,N_6981,N_6325);
and U7393 (N_7393,N_6944,N_6595);
xnor U7394 (N_7394,N_6507,N_6310);
and U7395 (N_7395,N_6819,N_6233);
and U7396 (N_7396,N_6400,N_6877);
nor U7397 (N_7397,N_6428,N_6247);
and U7398 (N_7398,N_6845,N_6574);
nor U7399 (N_7399,N_6220,N_6811);
nand U7400 (N_7400,N_6374,N_6836);
or U7401 (N_7401,N_6647,N_6178);
nand U7402 (N_7402,N_6965,N_6270);
nand U7403 (N_7403,N_6189,N_6271);
nor U7404 (N_7404,N_6491,N_6106);
and U7405 (N_7405,N_6889,N_6463);
nor U7406 (N_7406,N_6621,N_6525);
nand U7407 (N_7407,N_6748,N_6498);
nor U7408 (N_7408,N_6290,N_6713);
nand U7409 (N_7409,N_6887,N_6762);
or U7410 (N_7410,N_6175,N_6949);
or U7411 (N_7411,N_6994,N_6938);
nand U7412 (N_7412,N_6973,N_6659);
nand U7413 (N_7413,N_6425,N_6644);
and U7414 (N_7414,N_6733,N_6191);
or U7415 (N_7415,N_6947,N_6805);
nand U7416 (N_7416,N_6803,N_6732);
xnor U7417 (N_7417,N_6545,N_6063);
nand U7418 (N_7418,N_6769,N_6853);
and U7419 (N_7419,N_6849,N_6298);
nand U7420 (N_7420,N_6800,N_6555);
and U7421 (N_7421,N_6378,N_6906);
nor U7422 (N_7422,N_6951,N_6620);
nor U7423 (N_7423,N_6582,N_6731);
xor U7424 (N_7424,N_6631,N_6316);
nand U7425 (N_7425,N_6925,N_6409);
or U7426 (N_7426,N_6052,N_6978);
or U7427 (N_7427,N_6412,N_6420);
and U7428 (N_7428,N_6975,N_6652);
or U7429 (N_7429,N_6390,N_6508);
and U7430 (N_7430,N_6253,N_6782);
nor U7431 (N_7431,N_6557,N_6008);
and U7432 (N_7432,N_6754,N_6526);
nor U7433 (N_7433,N_6989,N_6764);
and U7434 (N_7434,N_6315,N_6982);
nor U7435 (N_7435,N_6967,N_6977);
xor U7436 (N_7436,N_6722,N_6830);
xor U7437 (N_7437,N_6852,N_6832);
nand U7438 (N_7438,N_6257,N_6376);
nand U7439 (N_7439,N_6383,N_6752);
or U7440 (N_7440,N_6309,N_6452);
nor U7441 (N_7441,N_6821,N_6387);
nand U7442 (N_7442,N_6548,N_6104);
and U7443 (N_7443,N_6911,N_6274);
nand U7444 (N_7444,N_6773,N_6549);
nand U7445 (N_7445,N_6825,N_6184);
and U7446 (N_7446,N_6284,N_6618);
nor U7447 (N_7447,N_6534,N_6057);
and U7448 (N_7448,N_6575,N_6602);
nor U7449 (N_7449,N_6826,N_6958);
nor U7450 (N_7450,N_6241,N_6179);
nand U7451 (N_7451,N_6655,N_6666);
or U7452 (N_7452,N_6144,N_6360);
and U7453 (N_7453,N_6693,N_6120);
nand U7454 (N_7454,N_6330,N_6841);
or U7455 (N_7455,N_6200,N_6940);
nand U7456 (N_7456,N_6914,N_6040);
nand U7457 (N_7457,N_6013,N_6946);
nor U7458 (N_7458,N_6292,N_6587);
nand U7459 (N_7459,N_6600,N_6584);
and U7460 (N_7460,N_6957,N_6043);
or U7461 (N_7461,N_6082,N_6155);
nor U7462 (N_7462,N_6936,N_6577);
or U7463 (N_7463,N_6928,N_6075);
nor U7464 (N_7464,N_6687,N_6987);
or U7465 (N_7465,N_6478,N_6670);
xor U7466 (N_7466,N_6642,N_6464);
and U7467 (N_7467,N_6708,N_6613);
and U7468 (N_7468,N_6851,N_6037);
nor U7469 (N_7469,N_6205,N_6149);
nand U7470 (N_7470,N_6385,N_6596);
nand U7471 (N_7471,N_6519,N_6294);
and U7472 (N_7472,N_6301,N_6237);
nor U7473 (N_7473,N_6181,N_6470);
nand U7474 (N_7474,N_6165,N_6531);
nor U7475 (N_7475,N_6381,N_6167);
nand U7476 (N_7476,N_6640,N_6177);
or U7477 (N_7477,N_6492,N_6289);
or U7478 (N_7478,N_6633,N_6328);
nand U7479 (N_7479,N_6735,N_6215);
and U7480 (N_7480,N_6405,N_6348);
and U7481 (N_7481,N_6648,N_6539);
nand U7482 (N_7482,N_6221,N_6885);
nand U7483 (N_7483,N_6101,N_6269);
nor U7484 (N_7484,N_6871,N_6893);
nor U7485 (N_7485,N_6610,N_6126);
xnor U7486 (N_7486,N_6668,N_6612);
nand U7487 (N_7487,N_6003,N_6245);
and U7488 (N_7488,N_6380,N_6594);
and U7489 (N_7489,N_6569,N_6103);
and U7490 (N_7490,N_6372,N_6123);
nand U7491 (N_7491,N_6153,N_6157);
nand U7492 (N_7492,N_6190,N_6920);
nor U7493 (N_7493,N_6543,N_6318);
or U7494 (N_7494,N_6098,N_6055);
nor U7495 (N_7495,N_6358,N_6336);
and U7496 (N_7496,N_6293,N_6122);
and U7497 (N_7497,N_6627,N_6546);
nor U7498 (N_7498,N_6859,N_6918);
nand U7499 (N_7499,N_6065,N_6344);
or U7500 (N_7500,N_6134,N_6742);
nor U7501 (N_7501,N_6266,N_6017);
nor U7502 (N_7502,N_6894,N_6159);
and U7503 (N_7503,N_6386,N_6694);
nand U7504 (N_7504,N_6099,N_6558);
and U7505 (N_7505,N_6218,N_6849);
nor U7506 (N_7506,N_6425,N_6974);
and U7507 (N_7507,N_6201,N_6232);
nor U7508 (N_7508,N_6742,N_6844);
xnor U7509 (N_7509,N_6574,N_6122);
nand U7510 (N_7510,N_6964,N_6744);
nor U7511 (N_7511,N_6547,N_6774);
xor U7512 (N_7512,N_6836,N_6812);
nand U7513 (N_7513,N_6885,N_6801);
or U7514 (N_7514,N_6510,N_6414);
nand U7515 (N_7515,N_6438,N_6294);
or U7516 (N_7516,N_6916,N_6582);
or U7517 (N_7517,N_6231,N_6136);
nor U7518 (N_7518,N_6179,N_6651);
and U7519 (N_7519,N_6260,N_6705);
nor U7520 (N_7520,N_6777,N_6432);
and U7521 (N_7521,N_6127,N_6950);
nor U7522 (N_7522,N_6039,N_6304);
and U7523 (N_7523,N_6817,N_6643);
and U7524 (N_7524,N_6988,N_6336);
nand U7525 (N_7525,N_6456,N_6308);
and U7526 (N_7526,N_6721,N_6636);
nand U7527 (N_7527,N_6566,N_6435);
nor U7528 (N_7528,N_6741,N_6095);
and U7529 (N_7529,N_6692,N_6717);
nor U7530 (N_7530,N_6483,N_6677);
nor U7531 (N_7531,N_6530,N_6401);
nor U7532 (N_7532,N_6056,N_6511);
or U7533 (N_7533,N_6420,N_6333);
and U7534 (N_7534,N_6771,N_6962);
nand U7535 (N_7535,N_6542,N_6099);
nor U7536 (N_7536,N_6223,N_6603);
nor U7537 (N_7537,N_6122,N_6536);
nor U7538 (N_7538,N_6265,N_6361);
nand U7539 (N_7539,N_6456,N_6862);
and U7540 (N_7540,N_6695,N_6952);
or U7541 (N_7541,N_6009,N_6357);
and U7542 (N_7542,N_6099,N_6618);
nand U7543 (N_7543,N_6973,N_6049);
and U7544 (N_7544,N_6531,N_6957);
or U7545 (N_7545,N_6001,N_6940);
nor U7546 (N_7546,N_6424,N_6274);
xor U7547 (N_7547,N_6306,N_6718);
nand U7548 (N_7548,N_6362,N_6303);
and U7549 (N_7549,N_6223,N_6974);
and U7550 (N_7550,N_6398,N_6395);
nor U7551 (N_7551,N_6998,N_6504);
and U7552 (N_7552,N_6384,N_6219);
nand U7553 (N_7553,N_6048,N_6969);
xnor U7554 (N_7554,N_6281,N_6293);
nor U7555 (N_7555,N_6741,N_6945);
nor U7556 (N_7556,N_6886,N_6594);
nor U7557 (N_7557,N_6265,N_6509);
and U7558 (N_7558,N_6065,N_6911);
and U7559 (N_7559,N_6081,N_6688);
xor U7560 (N_7560,N_6544,N_6451);
or U7561 (N_7561,N_6639,N_6399);
nand U7562 (N_7562,N_6974,N_6377);
nor U7563 (N_7563,N_6906,N_6917);
nor U7564 (N_7564,N_6318,N_6920);
nand U7565 (N_7565,N_6969,N_6608);
nor U7566 (N_7566,N_6624,N_6872);
or U7567 (N_7567,N_6320,N_6108);
nand U7568 (N_7568,N_6747,N_6487);
xor U7569 (N_7569,N_6362,N_6247);
and U7570 (N_7570,N_6617,N_6738);
nand U7571 (N_7571,N_6066,N_6640);
or U7572 (N_7572,N_6028,N_6023);
and U7573 (N_7573,N_6383,N_6514);
nor U7574 (N_7574,N_6781,N_6702);
nand U7575 (N_7575,N_6422,N_6104);
nor U7576 (N_7576,N_6847,N_6828);
xor U7577 (N_7577,N_6134,N_6417);
nor U7578 (N_7578,N_6671,N_6845);
and U7579 (N_7579,N_6713,N_6031);
or U7580 (N_7580,N_6812,N_6670);
nand U7581 (N_7581,N_6495,N_6058);
and U7582 (N_7582,N_6532,N_6761);
nand U7583 (N_7583,N_6238,N_6441);
nand U7584 (N_7584,N_6778,N_6680);
and U7585 (N_7585,N_6762,N_6893);
nand U7586 (N_7586,N_6387,N_6139);
nand U7587 (N_7587,N_6304,N_6952);
nand U7588 (N_7588,N_6618,N_6202);
nor U7589 (N_7589,N_6803,N_6529);
or U7590 (N_7590,N_6405,N_6607);
nand U7591 (N_7591,N_6546,N_6628);
nand U7592 (N_7592,N_6887,N_6384);
and U7593 (N_7593,N_6382,N_6090);
nand U7594 (N_7594,N_6704,N_6282);
or U7595 (N_7595,N_6196,N_6089);
xor U7596 (N_7596,N_6897,N_6248);
nand U7597 (N_7597,N_6166,N_6337);
or U7598 (N_7598,N_6467,N_6444);
or U7599 (N_7599,N_6645,N_6795);
and U7600 (N_7600,N_6885,N_6746);
nand U7601 (N_7601,N_6895,N_6009);
xnor U7602 (N_7602,N_6977,N_6959);
nor U7603 (N_7603,N_6646,N_6649);
and U7604 (N_7604,N_6359,N_6838);
nor U7605 (N_7605,N_6313,N_6281);
nand U7606 (N_7606,N_6257,N_6000);
nor U7607 (N_7607,N_6090,N_6916);
and U7608 (N_7608,N_6275,N_6689);
nor U7609 (N_7609,N_6031,N_6146);
and U7610 (N_7610,N_6885,N_6056);
or U7611 (N_7611,N_6462,N_6026);
nand U7612 (N_7612,N_6725,N_6073);
xor U7613 (N_7613,N_6704,N_6569);
xnor U7614 (N_7614,N_6741,N_6796);
nor U7615 (N_7615,N_6838,N_6617);
and U7616 (N_7616,N_6996,N_6086);
nor U7617 (N_7617,N_6414,N_6031);
or U7618 (N_7618,N_6309,N_6158);
nand U7619 (N_7619,N_6860,N_6807);
nand U7620 (N_7620,N_6709,N_6287);
and U7621 (N_7621,N_6714,N_6708);
nor U7622 (N_7622,N_6314,N_6416);
and U7623 (N_7623,N_6551,N_6597);
and U7624 (N_7624,N_6445,N_6964);
nor U7625 (N_7625,N_6805,N_6592);
nor U7626 (N_7626,N_6315,N_6233);
nand U7627 (N_7627,N_6684,N_6598);
xor U7628 (N_7628,N_6874,N_6893);
nor U7629 (N_7629,N_6743,N_6671);
or U7630 (N_7630,N_6781,N_6791);
and U7631 (N_7631,N_6444,N_6576);
nor U7632 (N_7632,N_6415,N_6638);
nor U7633 (N_7633,N_6891,N_6729);
xor U7634 (N_7634,N_6298,N_6624);
nand U7635 (N_7635,N_6445,N_6873);
or U7636 (N_7636,N_6858,N_6492);
and U7637 (N_7637,N_6341,N_6610);
nor U7638 (N_7638,N_6908,N_6512);
nor U7639 (N_7639,N_6457,N_6009);
or U7640 (N_7640,N_6835,N_6444);
and U7641 (N_7641,N_6944,N_6624);
or U7642 (N_7642,N_6783,N_6008);
nor U7643 (N_7643,N_6915,N_6773);
nor U7644 (N_7644,N_6708,N_6528);
or U7645 (N_7645,N_6032,N_6517);
or U7646 (N_7646,N_6557,N_6495);
nand U7647 (N_7647,N_6947,N_6543);
and U7648 (N_7648,N_6024,N_6625);
and U7649 (N_7649,N_6842,N_6328);
nor U7650 (N_7650,N_6209,N_6207);
nand U7651 (N_7651,N_6186,N_6615);
xor U7652 (N_7652,N_6888,N_6168);
or U7653 (N_7653,N_6829,N_6739);
nand U7654 (N_7654,N_6319,N_6716);
nand U7655 (N_7655,N_6891,N_6920);
or U7656 (N_7656,N_6741,N_6449);
nand U7657 (N_7657,N_6247,N_6994);
or U7658 (N_7658,N_6134,N_6340);
and U7659 (N_7659,N_6523,N_6351);
and U7660 (N_7660,N_6353,N_6398);
and U7661 (N_7661,N_6779,N_6484);
or U7662 (N_7662,N_6193,N_6239);
and U7663 (N_7663,N_6473,N_6233);
nor U7664 (N_7664,N_6476,N_6873);
nand U7665 (N_7665,N_6589,N_6581);
and U7666 (N_7666,N_6040,N_6757);
and U7667 (N_7667,N_6282,N_6202);
or U7668 (N_7668,N_6652,N_6957);
nand U7669 (N_7669,N_6316,N_6825);
nor U7670 (N_7670,N_6536,N_6091);
and U7671 (N_7671,N_6787,N_6300);
and U7672 (N_7672,N_6361,N_6282);
nand U7673 (N_7673,N_6911,N_6484);
nor U7674 (N_7674,N_6611,N_6591);
and U7675 (N_7675,N_6554,N_6581);
nor U7676 (N_7676,N_6512,N_6375);
and U7677 (N_7677,N_6302,N_6578);
xor U7678 (N_7678,N_6738,N_6990);
nor U7679 (N_7679,N_6381,N_6712);
nand U7680 (N_7680,N_6581,N_6269);
and U7681 (N_7681,N_6969,N_6258);
nor U7682 (N_7682,N_6445,N_6919);
xnor U7683 (N_7683,N_6433,N_6110);
nor U7684 (N_7684,N_6341,N_6530);
or U7685 (N_7685,N_6426,N_6886);
and U7686 (N_7686,N_6566,N_6582);
nand U7687 (N_7687,N_6439,N_6932);
and U7688 (N_7688,N_6733,N_6381);
nor U7689 (N_7689,N_6714,N_6945);
nor U7690 (N_7690,N_6016,N_6012);
nand U7691 (N_7691,N_6493,N_6010);
or U7692 (N_7692,N_6329,N_6487);
or U7693 (N_7693,N_6285,N_6051);
nand U7694 (N_7694,N_6411,N_6160);
nand U7695 (N_7695,N_6920,N_6100);
nand U7696 (N_7696,N_6349,N_6453);
nor U7697 (N_7697,N_6911,N_6777);
nor U7698 (N_7698,N_6793,N_6815);
or U7699 (N_7699,N_6308,N_6440);
xor U7700 (N_7700,N_6985,N_6489);
xnor U7701 (N_7701,N_6516,N_6251);
xnor U7702 (N_7702,N_6489,N_6801);
nand U7703 (N_7703,N_6561,N_6411);
or U7704 (N_7704,N_6831,N_6101);
nor U7705 (N_7705,N_6386,N_6222);
nor U7706 (N_7706,N_6636,N_6663);
nand U7707 (N_7707,N_6032,N_6128);
and U7708 (N_7708,N_6207,N_6699);
nor U7709 (N_7709,N_6242,N_6251);
nand U7710 (N_7710,N_6873,N_6024);
nand U7711 (N_7711,N_6516,N_6080);
and U7712 (N_7712,N_6809,N_6165);
and U7713 (N_7713,N_6941,N_6088);
nand U7714 (N_7714,N_6275,N_6688);
and U7715 (N_7715,N_6472,N_6253);
nand U7716 (N_7716,N_6292,N_6863);
nor U7717 (N_7717,N_6732,N_6674);
or U7718 (N_7718,N_6587,N_6709);
or U7719 (N_7719,N_6294,N_6949);
nand U7720 (N_7720,N_6009,N_6302);
and U7721 (N_7721,N_6988,N_6634);
nor U7722 (N_7722,N_6773,N_6599);
nor U7723 (N_7723,N_6488,N_6300);
nor U7724 (N_7724,N_6676,N_6233);
or U7725 (N_7725,N_6999,N_6848);
or U7726 (N_7726,N_6131,N_6322);
nor U7727 (N_7727,N_6077,N_6455);
or U7728 (N_7728,N_6525,N_6756);
and U7729 (N_7729,N_6205,N_6555);
nand U7730 (N_7730,N_6567,N_6416);
and U7731 (N_7731,N_6365,N_6915);
nor U7732 (N_7732,N_6854,N_6739);
nor U7733 (N_7733,N_6919,N_6614);
and U7734 (N_7734,N_6925,N_6281);
nor U7735 (N_7735,N_6506,N_6368);
nand U7736 (N_7736,N_6801,N_6498);
or U7737 (N_7737,N_6677,N_6631);
xor U7738 (N_7738,N_6394,N_6404);
nor U7739 (N_7739,N_6643,N_6046);
and U7740 (N_7740,N_6114,N_6093);
nor U7741 (N_7741,N_6842,N_6095);
or U7742 (N_7742,N_6211,N_6246);
and U7743 (N_7743,N_6127,N_6456);
or U7744 (N_7744,N_6804,N_6393);
and U7745 (N_7745,N_6706,N_6473);
or U7746 (N_7746,N_6838,N_6381);
xor U7747 (N_7747,N_6587,N_6787);
and U7748 (N_7748,N_6863,N_6184);
nor U7749 (N_7749,N_6819,N_6312);
or U7750 (N_7750,N_6754,N_6377);
nor U7751 (N_7751,N_6760,N_6429);
nand U7752 (N_7752,N_6185,N_6485);
nor U7753 (N_7753,N_6153,N_6477);
nand U7754 (N_7754,N_6201,N_6959);
nor U7755 (N_7755,N_6133,N_6056);
or U7756 (N_7756,N_6919,N_6370);
nand U7757 (N_7757,N_6107,N_6162);
nand U7758 (N_7758,N_6440,N_6428);
or U7759 (N_7759,N_6287,N_6767);
and U7760 (N_7760,N_6145,N_6343);
nor U7761 (N_7761,N_6398,N_6085);
nand U7762 (N_7762,N_6438,N_6142);
and U7763 (N_7763,N_6306,N_6218);
nor U7764 (N_7764,N_6271,N_6604);
nand U7765 (N_7765,N_6306,N_6213);
nand U7766 (N_7766,N_6832,N_6474);
and U7767 (N_7767,N_6867,N_6414);
or U7768 (N_7768,N_6200,N_6068);
or U7769 (N_7769,N_6263,N_6866);
nand U7770 (N_7770,N_6235,N_6762);
nand U7771 (N_7771,N_6462,N_6625);
nand U7772 (N_7772,N_6232,N_6287);
nor U7773 (N_7773,N_6656,N_6072);
nor U7774 (N_7774,N_6134,N_6414);
and U7775 (N_7775,N_6953,N_6855);
nor U7776 (N_7776,N_6038,N_6183);
nand U7777 (N_7777,N_6299,N_6999);
nand U7778 (N_7778,N_6398,N_6998);
and U7779 (N_7779,N_6353,N_6123);
nor U7780 (N_7780,N_6645,N_6140);
nand U7781 (N_7781,N_6296,N_6542);
or U7782 (N_7782,N_6743,N_6474);
nand U7783 (N_7783,N_6123,N_6323);
nand U7784 (N_7784,N_6423,N_6757);
nand U7785 (N_7785,N_6343,N_6965);
or U7786 (N_7786,N_6263,N_6003);
nor U7787 (N_7787,N_6826,N_6088);
nor U7788 (N_7788,N_6399,N_6747);
nand U7789 (N_7789,N_6334,N_6170);
and U7790 (N_7790,N_6885,N_6180);
nand U7791 (N_7791,N_6464,N_6038);
nand U7792 (N_7792,N_6625,N_6404);
nor U7793 (N_7793,N_6041,N_6665);
or U7794 (N_7794,N_6981,N_6500);
xnor U7795 (N_7795,N_6986,N_6278);
and U7796 (N_7796,N_6543,N_6525);
nand U7797 (N_7797,N_6200,N_6443);
and U7798 (N_7798,N_6291,N_6717);
nor U7799 (N_7799,N_6220,N_6849);
nand U7800 (N_7800,N_6993,N_6028);
xnor U7801 (N_7801,N_6051,N_6599);
nand U7802 (N_7802,N_6901,N_6833);
and U7803 (N_7803,N_6932,N_6693);
nand U7804 (N_7804,N_6178,N_6068);
nor U7805 (N_7805,N_6981,N_6124);
nor U7806 (N_7806,N_6758,N_6083);
or U7807 (N_7807,N_6839,N_6899);
nor U7808 (N_7808,N_6753,N_6397);
nand U7809 (N_7809,N_6340,N_6483);
and U7810 (N_7810,N_6827,N_6847);
and U7811 (N_7811,N_6753,N_6198);
xor U7812 (N_7812,N_6769,N_6678);
nor U7813 (N_7813,N_6289,N_6852);
or U7814 (N_7814,N_6174,N_6660);
nor U7815 (N_7815,N_6370,N_6442);
or U7816 (N_7816,N_6664,N_6790);
or U7817 (N_7817,N_6378,N_6221);
and U7818 (N_7818,N_6387,N_6571);
nor U7819 (N_7819,N_6523,N_6330);
nand U7820 (N_7820,N_6901,N_6395);
nand U7821 (N_7821,N_6581,N_6123);
nand U7822 (N_7822,N_6944,N_6529);
nand U7823 (N_7823,N_6830,N_6074);
or U7824 (N_7824,N_6942,N_6107);
or U7825 (N_7825,N_6242,N_6971);
and U7826 (N_7826,N_6431,N_6631);
and U7827 (N_7827,N_6259,N_6711);
nand U7828 (N_7828,N_6007,N_6202);
nor U7829 (N_7829,N_6147,N_6331);
nand U7830 (N_7830,N_6177,N_6446);
or U7831 (N_7831,N_6022,N_6944);
nor U7832 (N_7832,N_6600,N_6745);
or U7833 (N_7833,N_6870,N_6189);
or U7834 (N_7834,N_6854,N_6289);
nor U7835 (N_7835,N_6886,N_6766);
and U7836 (N_7836,N_6127,N_6450);
and U7837 (N_7837,N_6095,N_6473);
nand U7838 (N_7838,N_6790,N_6987);
and U7839 (N_7839,N_6667,N_6892);
nor U7840 (N_7840,N_6056,N_6639);
and U7841 (N_7841,N_6209,N_6962);
xor U7842 (N_7842,N_6017,N_6262);
nand U7843 (N_7843,N_6230,N_6890);
or U7844 (N_7844,N_6473,N_6146);
nor U7845 (N_7845,N_6849,N_6422);
nor U7846 (N_7846,N_6725,N_6182);
nand U7847 (N_7847,N_6028,N_6416);
nor U7848 (N_7848,N_6897,N_6594);
nand U7849 (N_7849,N_6784,N_6109);
or U7850 (N_7850,N_6520,N_6709);
xnor U7851 (N_7851,N_6647,N_6309);
nor U7852 (N_7852,N_6158,N_6678);
nor U7853 (N_7853,N_6178,N_6285);
nor U7854 (N_7854,N_6572,N_6053);
nor U7855 (N_7855,N_6629,N_6292);
nand U7856 (N_7856,N_6970,N_6187);
nor U7857 (N_7857,N_6592,N_6744);
or U7858 (N_7858,N_6855,N_6497);
nor U7859 (N_7859,N_6314,N_6636);
and U7860 (N_7860,N_6870,N_6064);
and U7861 (N_7861,N_6080,N_6496);
and U7862 (N_7862,N_6443,N_6967);
xnor U7863 (N_7863,N_6959,N_6321);
nand U7864 (N_7864,N_6877,N_6907);
nor U7865 (N_7865,N_6329,N_6730);
xnor U7866 (N_7866,N_6395,N_6601);
nor U7867 (N_7867,N_6117,N_6987);
nand U7868 (N_7868,N_6930,N_6635);
nand U7869 (N_7869,N_6696,N_6962);
or U7870 (N_7870,N_6955,N_6635);
xor U7871 (N_7871,N_6836,N_6682);
nor U7872 (N_7872,N_6094,N_6140);
xnor U7873 (N_7873,N_6568,N_6996);
and U7874 (N_7874,N_6473,N_6137);
nor U7875 (N_7875,N_6184,N_6071);
or U7876 (N_7876,N_6585,N_6112);
nor U7877 (N_7877,N_6883,N_6376);
or U7878 (N_7878,N_6920,N_6654);
nand U7879 (N_7879,N_6373,N_6069);
nand U7880 (N_7880,N_6243,N_6315);
nand U7881 (N_7881,N_6133,N_6359);
and U7882 (N_7882,N_6200,N_6523);
nor U7883 (N_7883,N_6704,N_6372);
nand U7884 (N_7884,N_6680,N_6757);
and U7885 (N_7885,N_6636,N_6261);
nor U7886 (N_7886,N_6398,N_6007);
nor U7887 (N_7887,N_6717,N_6031);
nand U7888 (N_7888,N_6358,N_6447);
nor U7889 (N_7889,N_6032,N_6614);
or U7890 (N_7890,N_6367,N_6751);
nand U7891 (N_7891,N_6082,N_6028);
and U7892 (N_7892,N_6940,N_6672);
nor U7893 (N_7893,N_6783,N_6591);
and U7894 (N_7894,N_6267,N_6327);
nor U7895 (N_7895,N_6087,N_6915);
or U7896 (N_7896,N_6234,N_6722);
and U7897 (N_7897,N_6256,N_6459);
or U7898 (N_7898,N_6705,N_6041);
nor U7899 (N_7899,N_6871,N_6270);
and U7900 (N_7900,N_6490,N_6787);
nor U7901 (N_7901,N_6820,N_6911);
and U7902 (N_7902,N_6534,N_6441);
nand U7903 (N_7903,N_6035,N_6698);
nand U7904 (N_7904,N_6972,N_6148);
nor U7905 (N_7905,N_6053,N_6741);
nor U7906 (N_7906,N_6293,N_6300);
nand U7907 (N_7907,N_6341,N_6722);
nor U7908 (N_7908,N_6926,N_6499);
and U7909 (N_7909,N_6296,N_6189);
nor U7910 (N_7910,N_6124,N_6419);
and U7911 (N_7911,N_6577,N_6597);
nand U7912 (N_7912,N_6535,N_6114);
nand U7913 (N_7913,N_6243,N_6816);
or U7914 (N_7914,N_6523,N_6015);
or U7915 (N_7915,N_6100,N_6951);
and U7916 (N_7916,N_6958,N_6913);
and U7917 (N_7917,N_6715,N_6839);
or U7918 (N_7918,N_6664,N_6264);
and U7919 (N_7919,N_6938,N_6084);
nand U7920 (N_7920,N_6664,N_6904);
nand U7921 (N_7921,N_6285,N_6938);
and U7922 (N_7922,N_6496,N_6010);
nor U7923 (N_7923,N_6407,N_6428);
nor U7924 (N_7924,N_6925,N_6425);
nand U7925 (N_7925,N_6122,N_6513);
nor U7926 (N_7926,N_6484,N_6162);
or U7927 (N_7927,N_6441,N_6336);
nor U7928 (N_7928,N_6642,N_6907);
nand U7929 (N_7929,N_6112,N_6236);
or U7930 (N_7930,N_6574,N_6165);
nor U7931 (N_7931,N_6707,N_6997);
and U7932 (N_7932,N_6065,N_6281);
nor U7933 (N_7933,N_6396,N_6261);
or U7934 (N_7934,N_6802,N_6553);
or U7935 (N_7935,N_6635,N_6295);
nand U7936 (N_7936,N_6419,N_6482);
nor U7937 (N_7937,N_6650,N_6710);
and U7938 (N_7938,N_6779,N_6414);
xnor U7939 (N_7939,N_6793,N_6389);
nor U7940 (N_7940,N_6639,N_6062);
nand U7941 (N_7941,N_6452,N_6125);
and U7942 (N_7942,N_6488,N_6707);
and U7943 (N_7943,N_6600,N_6929);
and U7944 (N_7944,N_6388,N_6248);
or U7945 (N_7945,N_6971,N_6543);
and U7946 (N_7946,N_6508,N_6256);
or U7947 (N_7947,N_6787,N_6371);
nand U7948 (N_7948,N_6120,N_6605);
nand U7949 (N_7949,N_6002,N_6127);
and U7950 (N_7950,N_6448,N_6676);
and U7951 (N_7951,N_6100,N_6591);
xnor U7952 (N_7952,N_6921,N_6190);
or U7953 (N_7953,N_6377,N_6876);
and U7954 (N_7954,N_6979,N_6717);
xor U7955 (N_7955,N_6310,N_6264);
or U7956 (N_7956,N_6359,N_6818);
and U7957 (N_7957,N_6498,N_6729);
nor U7958 (N_7958,N_6000,N_6464);
or U7959 (N_7959,N_6629,N_6044);
nand U7960 (N_7960,N_6136,N_6409);
nand U7961 (N_7961,N_6632,N_6303);
xnor U7962 (N_7962,N_6201,N_6574);
nor U7963 (N_7963,N_6862,N_6510);
and U7964 (N_7964,N_6047,N_6202);
and U7965 (N_7965,N_6017,N_6765);
nand U7966 (N_7966,N_6424,N_6178);
nand U7967 (N_7967,N_6499,N_6527);
or U7968 (N_7968,N_6162,N_6755);
and U7969 (N_7969,N_6785,N_6252);
nand U7970 (N_7970,N_6415,N_6135);
nor U7971 (N_7971,N_6829,N_6048);
or U7972 (N_7972,N_6279,N_6294);
or U7973 (N_7973,N_6449,N_6662);
and U7974 (N_7974,N_6492,N_6669);
or U7975 (N_7975,N_6521,N_6308);
nor U7976 (N_7976,N_6330,N_6509);
or U7977 (N_7977,N_6504,N_6861);
nand U7978 (N_7978,N_6682,N_6760);
and U7979 (N_7979,N_6688,N_6744);
nand U7980 (N_7980,N_6646,N_6050);
and U7981 (N_7981,N_6075,N_6829);
or U7982 (N_7982,N_6009,N_6523);
nand U7983 (N_7983,N_6047,N_6595);
and U7984 (N_7984,N_6735,N_6641);
nand U7985 (N_7985,N_6184,N_6475);
nand U7986 (N_7986,N_6951,N_6085);
xnor U7987 (N_7987,N_6185,N_6369);
and U7988 (N_7988,N_6685,N_6864);
nor U7989 (N_7989,N_6230,N_6046);
nand U7990 (N_7990,N_6570,N_6515);
and U7991 (N_7991,N_6742,N_6287);
or U7992 (N_7992,N_6573,N_6600);
and U7993 (N_7993,N_6710,N_6520);
or U7994 (N_7994,N_6975,N_6532);
and U7995 (N_7995,N_6542,N_6462);
and U7996 (N_7996,N_6204,N_6890);
or U7997 (N_7997,N_6668,N_6946);
and U7998 (N_7998,N_6942,N_6486);
or U7999 (N_7999,N_6083,N_6439);
or U8000 (N_8000,N_7061,N_7534);
and U8001 (N_8001,N_7063,N_7227);
nor U8002 (N_8002,N_7810,N_7753);
nand U8003 (N_8003,N_7032,N_7192);
xnor U8004 (N_8004,N_7423,N_7215);
nor U8005 (N_8005,N_7079,N_7676);
and U8006 (N_8006,N_7732,N_7953);
nor U8007 (N_8007,N_7211,N_7783);
xor U8008 (N_8008,N_7619,N_7538);
nand U8009 (N_8009,N_7963,N_7266);
or U8010 (N_8010,N_7555,N_7915);
or U8011 (N_8011,N_7411,N_7491);
and U8012 (N_8012,N_7735,N_7277);
nand U8013 (N_8013,N_7900,N_7134);
or U8014 (N_8014,N_7582,N_7125);
nand U8015 (N_8015,N_7451,N_7090);
nor U8016 (N_8016,N_7165,N_7999);
or U8017 (N_8017,N_7151,N_7637);
nor U8018 (N_8018,N_7180,N_7386);
or U8019 (N_8019,N_7575,N_7808);
and U8020 (N_8020,N_7271,N_7099);
nor U8021 (N_8021,N_7991,N_7472);
and U8022 (N_8022,N_7527,N_7996);
or U8023 (N_8023,N_7250,N_7967);
or U8024 (N_8024,N_7843,N_7228);
or U8025 (N_8025,N_7235,N_7458);
xor U8026 (N_8026,N_7248,N_7425);
nand U8027 (N_8027,N_7142,N_7096);
and U8028 (N_8028,N_7364,N_7412);
nor U8029 (N_8029,N_7340,N_7093);
and U8030 (N_8030,N_7357,N_7368);
and U8031 (N_8031,N_7195,N_7471);
nand U8032 (N_8032,N_7204,N_7485);
nor U8033 (N_8033,N_7954,N_7322);
nand U8034 (N_8034,N_7818,N_7421);
nand U8035 (N_8035,N_7070,N_7443);
nor U8036 (N_8036,N_7223,N_7780);
or U8037 (N_8037,N_7932,N_7758);
xor U8038 (N_8038,N_7716,N_7001);
nand U8039 (N_8039,N_7764,N_7292);
or U8040 (N_8040,N_7429,N_7087);
xnor U8041 (N_8041,N_7601,N_7157);
xor U8042 (N_8042,N_7489,N_7349);
nor U8043 (N_8043,N_7715,N_7072);
and U8044 (N_8044,N_7759,N_7171);
and U8045 (N_8045,N_7650,N_7994);
nand U8046 (N_8046,N_7182,N_7435);
or U8047 (N_8047,N_7671,N_7642);
and U8048 (N_8048,N_7988,N_7413);
nand U8049 (N_8049,N_7950,N_7144);
and U8050 (N_8050,N_7960,N_7338);
or U8051 (N_8051,N_7749,N_7444);
and U8052 (N_8052,N_7921,N_7640);
and U8053 (N_8053,N_7437,N_7146);
xor U8054 (N_8054,N_7710,N_7867);
nor U8055 (N_8055,N_7889,N_7612);
nand U8056 (N_8056,N_7969,N_7310);
xor U8057 (N_8057,N_7073,N_7104);
nor U8058 (N_8058,N_7822,N_7975);
and U8059 (N_8059,N_7559,N_7707);
or U8060 (N_8060,N_7321,N_7914);
xor U8061 (N_8061,N_7567,N_7805);
xor U8062 (N_8062,N_7268,N_7863);
nor U8063 (N_8063,N_7939,N_7795);
and U8064 (N_8064,N_7592,N_7419);
or U8065 (N_8065,N_7557,N_7771);
nand U8066 (N_8066,N_7272,N_7560);
or U8067 (N_8067,N_7137,N_7378);
nand U8068 (N_8068,N_7325,N_7839);
nor U8069 (N_8069,N_7660,N_7428);
and U8070 (N_8070,N_7877,N_7332);
nand U8071 (N_8071,N_7649,N_7750);
and U8072 (N_8072,N_7673,N_7447);
and U8073 (N_8073,N_7633,N_7085);
nand U8074 (N_8074,N_7162,N_7442);
and U8075 (N_8075,N_7845,N_7012);
nand U8076 (N_8076,N_7956,N_7462);
nor U8077 (N_8077,N_7488,N_7351);
nand U8078 (N_8078,N_7704,N_7329);
nor U8079 (N_8079,N_7029,N_7422);
xnor U8080 (N_8080,N_7686,N_7053);
or U8081 (N_8081,N_7264,N_7047);
nor U8082 (N_8082,N_7404,N_7634);
nor U8083 (N_8083,N_7212,N_7852);
nand U8084 (N_8084,N_7806,N_7885);
nor U8085 (N_8085,N_7232,N_7761);
nor U8086 (N_8086,N_7393,N_7200);
nand U8087 (N_8087,N_7928,N_7618);
nand U8088 (N_8088,N_7553,N_7479);
and U8089 (N_8089,N_7807,N_7525);
and U8090 (N_8090,N_7821,N_7345);
xor U8091 (N_8091,N_7974,N_7729);
or U8092 (N_8092,N_7734,N_7544);
nand U8093 (N_8093,N_7628,N_7667);
nor U8094 (N_8094,N_7895,N_7418);
nand U8095 (N_8095,N_7275,N_7907);
nor U8096 (N_8096,N_7240,N_7997);
xor U8097 (N_8097,N_7978,N_7888);
nor U8098 (N_8098,N_7905,N_7456);
and U8099 (N_8099,N_7789,N_7820);
and U8100 (N_8100,N_7782,N_7655);
nand U8101 (N_8101,N_7880,N_7778);
or U8102 (N_8102,N_7962,N_7762);
or U8103 (N_8103,N_7840,N_7376);
or U8104 (N_8104,N_7247,N_7936);
or U8105 (N_8105,N_7593,N_7835);
nor U8106 (N_8106,N_7656,N_7587);
nor U8107 (N_8107,N_7518,N_7058);
and U8108 (N_8108,N_7140,N_7241);
and U8109 (N_8109,N_7218,N_7927);
xnor U8110 (N_8110,N_7955,N_7632);
or U8111 (N_8111,N_7003,N_7493);
and U8112 (N_8112,N_7385,N_7558);
nor U8113 (N_8113,N_7849,N_7167);
or U8114 (N_8114,N_7006,N_7893);
and U8115 (N_8115,N_7505,N_7647);
nor U8116 (N_8116,N_7887,N_7375);
and U8117 (N_8117,N_7258,N_7536);
nand U8118 (N_8118,N_7233,N_7478);
xor U8119 (N_8119,N_7293,N_7653);
and U8120 (N_8120,N_7082,N_7530);
or U8121 (N_8121,N_7949,N_7688);
or U8122 (N_8122,N_7133,N_7797);
or U8123 (N_8123,N_7754,N_7743);
nand U8124 (N_8124,N_7202,N_7139);
nand U8125 (N_8125,N_7516,N_7860);
nand U8126 (N_8126,N_7498,N_7513);
or U8127 (N_8127,N_7665,N_7940);
nand U8128 (N_8128,N_7737,N_7288);
nand U8129 (N_8129,N_7508,N_7579);
nand U8130 (N_8130,N_7366,N_7751);
and U8131 (N_8131,N_7919,N_7842);
nor U8132 (N_8132,N_7021,N_7685);
or U8133 (N_8133,N_7023,N_7580);
nor U8134 (N_8134,N_7123,N_7262);
xor U8135 (N_8135,N_7205,N_7234);
nor U8136 (N_8136,N_7229,N_7563);
or U8137 (N_8137,N_7920,N_7050);
nand U8138 (N_8138,N_7521,N_7600);
xnor U8139 (N_8139,N_7630,N_7452);
nand U8140 (N_8140,N_7038,N_7353);
or U8141 (N_8141,N_7341,N_7448);
nand U8142 (N_8142,N_7858,N_7196);
nand U8143 (N_8143,N_7018,N_7209);
xnor U8144 (N_8144,N_7347,N_7473);
or U8145 (N_8145,N_7106,N_7668);
and U8146 (N_8146,N_7257,N_7725);
xor U8147 (N_8147,N_7186,N_7365);
nand U8148 (N_8148,N_7147,N_7613);
or U8149 (N_8149,N_7982,N_7851);
nor U8150 (N_8150,N_7691,N_7168);
nand U8151 (N_8151,N_7705,N_7625);
and U8152 (N_8152,N_7026,N_7416);
xnor U8153 (N_8153,N_7817,N_7014);
or U8154 (N_8154,N_7239,N_7581);
xnor U8155 (N_8155,N_7740,N_7254);
and U8156 (N_8156,N_7057,N_7361);
or U8157 (N_8157,N_7721,N_7203);
or U8158 (N_8158,N_7551,N_7689);
and U8159 (N_8159,N_7602,N_7641);
and U8160 (N_8160,N_7577,N_7924);
nand U8161 (N_8161,N_7410,N_7497);
and U8162 (N_8162,N_7078,N_7221);
or U8163 (N_8163,N_7285,N_7523);
nor U8164 (N_8164,N_7185,N_7874);
and U8165 (N_8165,N_7714,N_7399);
nand U8166 (N_8166,N_7446,N_7155);
or U8167 (N_8167,N_7496,N_7048);
nand U8168 (N_8168,N_7501,N_7396);
xor U8169 (N_8169,N_7315,N_7515);
and U8170 (N_8170,N_7738,N_7263);
or U8171 (N_8171,N_7397,N_7319);
xor U8172 (N_8172,N_7701,N_7979);
or U8173 (N_8173,N_7039,N_7220);
nor U8174 (N_8174,N_7894,N_7379);
and U8175 (N_8175,N_7346,N_7219);
nor U8176 (N_8176,N_7164,N_7583);
or U8177 (N_8177,N_7105,N_7430);
nor U8178 (N_8178,N_7426,N_7286);
nand U8179 (N_8179,N_7143,N_7794);
nor U8180 (N_8180,N_7111,N_7985);
nor U8181 (N_8181,N_7645,N_7486);
nand U8182 (N_8182,N_7015,N_7398);
nor U8183 (N_8183,N_7333,N_7069);
nor U8184 (N_8184,N_7432,N_7279);
or U8185 (N_8185,N_7269,N_7377);
nand U8186 (N_8186,N_7942,N_7776);
or U8187 (N_8187,N_7722,N_7261);
nor U8188 (N_8188,N_7083,N_7627);
nand U8189 (N_8189,N_7094,N_7173);
nor U8190 (N_8190,N_7296,N_7054);
nand U8191 (N_8191,N_7311,N_7862);
nand U8192 (N_8192,N_7302,N_7502);
and U8193 (N_8193,N_7194,N_7826);
and U8194 (N_8194,N_7779,N_7475);
nand U8195 (N_8195,N_7372,N_7120);
or U8196 (N_8196,N_7700,N_7813);
and U8197 (N_8197,N_7896,N_7482);
and U8198 (N_8198,N_7713,N_7910);
and U8199 (N_8199,N_7103,N_7121);
xnor U8200 (N_8200,N_7415,N_7884);
and U8201 (N_8201,N_7855,N_7336);
nand U8202 (N_8202,N_7499,N_7916);
and U8203 (N_8203,N_7098,N_7533);
and U8204 (N_8204,N_7854,N_7868);
nand U8205 (N_8205,N_7477,N_7403);
nand U8206 (N_8206,N_7687,N_7830);
nor U8207 (N_8207,N_7067,N_7998);
nor U8208 (N_8208,N_7864,N_7253);
or U8209 (N_8209,N_7675,N_7586);
xnor U8210 (N_8210,N_7214,N_7131);
nor U8211 (N_8211,N_7929,N_7781);
nor U8212 (N_8212,N_7334,N_7730);
nand U8213 (N_8213,N_7175,N_7948);
nor U8214 (N_8214,N_7681,N_7574);
and U8215 (N_8215,N_7951,N_7007);
or U8216 (N_8216,N_7172,N_7037);
nor U8217 (N_8217,N_7484,N_7829);
nor U8218 (N_8218,N_7387,N_7958);
and U8219 (N_8219,N_7439,N_7692);
or U8220 (N_8220,N_7408,N_7362);
and U8221 (N_8221,N_7210,N_7395);
and U8222 (N_8222,N_7152,N_7252);
and U8223 (N_8223,N_7961,N_7135);
nor U8224 (N_8224,N_7976,N_7166);
nand U8225 (N_8225,N_7947,N_7548);
and U8226 (N_8226,N_7391,N_7331);
or U8227 (N_8227,N_7453,N_7766);
or U8228 (N_8228,N_7564,N_7184);
and U8229 (N_8229,N_7774,N_7149);
nand U8230 (N_8230,N_7610,N_7249);
and U8231 (N_8231,N_7595,N_7657);
nor U8232 (N_8232,N_7305,N_7791);
or U8233 (N_8233,N_7284,N_7912);
xnor U8234 (N_8234,N_7622,N_7646);
nand U8235 (N_8235,N_7492,N_7370);
nand U8236 (N_8236,N_7526,N_7925);
and U8237 (N_8237,N_7599,N_7011);
xor U8238 (N_8238,N_7320,N_7158);
or U8239 (N_8239,N_7741,N_7876);
and U8240 (N_8240,N_7040,N_7460);
nor U8241 (N_8241,N_7666,N_7303);
nor U8242 (N_8242,N_7578,N_7883);
and U8243 (N_8243,N_7267,N_7828);
nor U8244 (N_8244,N_7242,N_7405);
nand U8245 (N_8245,N_7697,N_7207);
nor U8246 (N_8246,N_7841,N_7314);
and U8247 (N_8247,N_7494,N_7181);
nand U8248 (N_8248,N_7763,N_7980);
nor U8249 (N_8249,N_7307,N_7931);
or U8250 (N_8250,N_7658,N_7068);
and U8251 (N_8251,N_7222,N_7720);
xor U8252 (N_8252,N_7785,N_7313);
nor U8253 (N_8253,N_7208,N_7875);
nor U8254 (N_8254,N_7765,N_7108);
nand U8255 (N_8255,N_7092,N_7684);
and U8256 (N_8256,N_7065,N_7406);
xor U8257 (N_8257,N_7431,N_7596);
nand U8258 (N_8258,N_7572,N_7190);
nor U8259 (N_8259,N_7116,N_7076);
nand U8260 (N_8260,N_7114,N_7971);
or U8261 (N_8261,N_7747,N_7295);
nor U8262 (N_8262,N_7230,N_7170);
xnor U8263 (N_8263,N_7348,N_7873);
nor U8264 (N_8264,N_7352,N_7441);
or U8265 (N_8265,N_7424,N_7831);
nor U8266 (N_8266,N_7274,N_7723);
nand U8267 (N_8267,N_7464,N_7191);
and U8268 (N_8268,N_7597,N_7787);
nand U8269 (N_8269,N_7651,N_7708);
or U8270 (N_8270,N_7016,N_7746);
or U8271 (N_8271,N_7588,N_7838);
nor U8272 (N_8272,N_7992,N_7861);
or U8273 (N_8273,N_7752,N_7614);
xnor U8274 (N_8274,N_7519,N_7363);
and U8275 (N_8275,N_7051,N_7183);
nand U8276 (N_8276,N_7324,N_7000);
nand U8277 (N_8277,N_7524,N_7512);
or U8278 (N_8278,N_7100,N_7540);
nor U8279 (N_8279,N_7127,N_7719);
nand U8280 (N_8280,N_7299,N_7727);
or U8281 (N_8281,N_7077,N_7966);
nor U8282 (N_8282,N_7318,N_7846);
nor U8283 (N_8283,N_7584,N_7476);
xnor U8284 (N_8284,N_7224,N_7853);
or U8285 (N_8285,N_7811,N_7480);
nor U8286 (N_8286,N_7280,N_7554);
xor U8287 (N_8287,N_7672,N_7522);
and U8288 (N_8288,N_7045,N_7129);
nand U8289 (N_8289,N_7031,N_7033);
or U8290 (N_8290,N_7606,N_7993);
or U8291 (N_8291,N_7008,N_7436);
nand U8292 (N_8292,N_7273,N_7744);
nand U8293 (N_8293,N_7815,N_7798);
nor U8294 (N_8294,N_7312,N_7836);
and U8295 (N_8295,N_7690,N_7825);
xnor U8296 (N_8296,N_7381,N_7661);
nor U8297 (N_8297,N_7400,N_7968);
xor U8298 (N_8298,N_7897,N_7847);
nor U8299 (N_8299,N_7682,N_7944);
and U8300 (N_8300,N_7648,N_7055);
xor U8301 (N_8301,N_7027,N_7814);
and U8302 (N_8302,N_7308,N_7504);
nand U8303 (N_8303,N_7298,N_7760);
nor U8304 (N_8304,N_7878,N_7454);
xor U8305 (N_8305,N_7392,N_7706);
nor U8306 (N_8306,N_7095,N_7696);
xor U8307 (N_8307,N_7793,N_7904);
and U8308 (N_8308,N_7118,N_7569);
and U8309 (N_8309,N_7693,N_7571);
or U8310 (N_8310,N_7898,N_7112);
and U8311 (N_8311,N_7260,N_7490);
nand U8312 (N_8312,N_7128,N_7695);
nor U8313 (N_8313,N_7407,N_7136);
nor U8314 (N_8314,N_7470,N_7297);
or U8315 (N_8315,N_7122,N_7259);
and U8316 (N_8316,N_7117,N_7736);
and U8317 (N_8317,N_7394,N_7709);
nand U8318 (N_8318,N_7281,N_7495);
nand U8319 (N_8319,N_7193,N_7344);
or U8320 (N_8320,N_7834,N_7265);
nor U8321 (N_8321,N_7644,N_7570);
nor U8322 (N_8322,N_7019,N_7433);
and U8323 (N_8323,N_7388,N_7141);
xnor U8324 (N_8324,N_7276,N_7371);
nor U8325 (N_8325,N_7631,N_7350);
nor U8326 (N_8326,N_7323,N_7603);
xor U8327 (N_8327,N_7742,N_7621);
or U8328 (N_8328,N_7585,N_7624);
nor U8329 (N_8329,N_7532,N_7608);
or U8330 (N_8330,N_7995,N_7035);
nand U8331 (N_8331,N_7169,N_7154);
or U8332 (N_8332,N_7594,N_7237);
nor U8333 (N_8333,N_7984,N_7198);
nand U8334 (N_8334,N_7153,N_7132);
xor U8335 (N_8335,N_7110,N_7881);
xnor U8336 (N_8336,N_7679,N_7773);
or U8337 (N_8337,N_7552,N_7712);
nand U8338 (N_8338,N_7503,N_7531);
nand U8339 (N_8339,N_7483,N_7420);
and U8340 (N_8340,N_7699,N_7517);
nor U8341 (N_8341,N_7549,N_7440);
nand U8342 (N_8342,N_7529,N_7043);
nand U8343 (N_8343,N_7089,N_7163);
xnor U8344 (N_8344,N_7964,N_7358);
nor U8345 (N_8345,N_7010,N_7300);
nor U8346 (N_8346,N_7803,N_7837);
and U8347 (N_8347,N_7243,N_7663);
or U8348 (N_8348,N_7983,N_7882);
nand U8349 (N_8349,N_7355,N_7786);
and U8350 (N_8350,N_7115,N_7102);
and U8351 (N_8351,N_7041,N_7449);
and U8352 (N_8352,N_7629,N_7981);
and U8353 (N_8353,N_7251,N_7330);
nor U8354 (N_8354,N_7062,N_7680);
xnor U8355 (N_8355,N_7414,N_7568);
nor U8356 (N_8356,N_7772,N_7565);
xnor U8357 (N_8357,N_7977,N_7930);
xor U8358 (N_8358,N_7866,N_7130);
or U8359 (N_8359,N_7450,N_7457);
nand U8360 (N_8360,N_7463,N_7282);
and U8361 (N_8361,N_7402,N_7389);
nor U8362 (N_8362,N_7197,N_7711);
xor U8363 (N_8363,N_7635,N_7075);
nor U8364 (N_8364,N_7790,N_7879);
or U8365 (N_8365,N_7002,N_7788);
xnor U8366 (N_8366,N_7150,N_7466);
nor U8367 (N_8367,N_7659,N_7683);
xor U8368 (N_8368,N_7620,N_7187);
nor U8369 (N_8369,N_7703,N_7617);
or U8370 (N_8370,N_7986,N_7113);
and U8371 (N_8371,N_7445,N_7824);
nor U8372 (N_8372,N_7856,N_7309);
or U8373 (N_8373,N_7890,N_7176);
or U8374 (N_8374,N_7091,N_7832);
nor U8375 (N_8375,N_7046,N_7913);
and U8376 (N_8376,N_7674,N_7935);
nand U8377 (N_8377,N_7028,N_7812);
or U8378 (N_8378,N_7796,N_7561);
nor U8379 (N_8379,N_7800,N_7294);
xor U8380 (N_8380,N_7576,N_7246);
nand U8381 (N_8381,N_7064,N_7605);
nand U8382 (N_8382,N_7946,N_7654);
xor U8383 (N_8383,N_7459,N_7731);
nand U8384 (N_8384,N_7317,N_7071);
or U8385 (N_8385,N_7970,N_7899);
or U8386 (N_8386,N_7636,N_7052);
xnor U8387 (N_8387,N_7022,N_7188);
or U8388 (N_8388,N_7909,N_7342);
and U8389 (N_8389,N_7335,N_7256);
nand U8390 (N_8390,N_7179,N_7590);
or U8391 (N_8391,N_7550,N_7678);
nor U8392 (N_8392,N_7804,N_7107);
xnor U8393 (N_8393,N_7020,N_7066);
nand U8394 (N_8394,N_7161,N_7865);
and U8395 (N_8395,N_7859,N_7231);
or U8396 (N_8396,N_7409,N_7145);
and U8397 (N_8397,N_7468,N_7922);
and U8398 (N_8398,N_7417,N_7049);
nor U8399 (N_8399,N_7373,N_7367);
and U8400 (N_8400,N_7156,N_7500);
nand U8401 (N_8401,N_7160,N_7304);
or U8402 (N_8402,N_7514,N_7662);
nor U8403 (N_8403,N_7081,N_7034);
nor U8404 (N_8404,N_7802,N_7987);
nand U8405 (N_8405,N_7702,N_7535);
and U8406 (N_8406,N_7573,N_7957);
and U8407 (N_8407,N_7965,N_7902);
nand U8408 (N_8408,N_7086,N_7611);
and U8409 (N_8409,N_7384,N_7427);
nand U8410 (N_8410,N_7626,N_7748);
nor U8411 (N_8411,N_7101,N_7886);
nor U8412 (N_8412,N_7326,N_7537);
nor U8413 (N_8413,N_7546,N_7343);
nor U8414 (N_8414,N_7777,N_7848);
and U8415 (N_8415,N_7255,N_7545);
nand U8416 (N_8416,N_7177,N_7467);
nand U8417 (N_8417,N_7465,N_7871);
or U8418 (N_8418,N_7278,N_7327);
and U8419 (N_8419,N_7652,N_7088);
or U8420 (N_8420,N_7383,N_7434);
or U8421 (N_8421,N_7784,N_7543);
nor U8422 (N_8422,N_7566,N_7301);
xnor U8423 (N_8423,N_7174,N_7005);
and U8424 (N_8424,N_7918,N_7287);
xnor U8425 (N_8425,N_7827,N_7556);
nand U8426 (N_8426,N_7507,N_7756);
or U8427 (N_8427,N_7542,N_7178);
and U8428 (N_8428,N_7474,N_7892);
nand U8429 (N_8429,N_7717,N_7669);
nor U8430 (N_8430,N_7639,N_7004);
and U8431 (N_8431,N_7289,N_7044);
and U8432 (N_8432,N_7726,N_7908);
nand U8433 (N_8433,N_7799,N_7316);
nand U8434 (N_8434,N_7511,N_7213);
nand U8435 (N_8435,N_7792,N_7591);
and U8436 (N_8436,N_7872,N_7850);
nand U8437 (N_8437,N_7733,N_7901);
nand U8438 (N_8438,N_7917,N_7767);
or U8439 (N_8439,N_7891,N_7934);
and U8440 (N_8440,N_7816,N_7923);
or U8441 (N_8441,N_7159,N_7670);
or U8442 (N_8442,N_7306,N_7952);
or U8443 (N_8443,N_7017,N_7819);
or U8444 (N_8444,N_7903,N_7718);
xnor U8445 (N_8445,N_7060,N_7124);
nand U8446 (N_8446,N_7926,N_7487);
nor U8447 (N_8447,N_7959,N_7539);
or U8448 (N_8448,N_7481,N_7643);
nand U8449 (N_8449,N_7933,N_7937);
or U8450 (N_8450,N_7080,N_7339);
and U8451 (N_8451,N_7359,N_7598);
xnor U8452 (N_8452,N_7990,N_7290);
and U8453 (N_8453,N_7199,N_7972);
nand U8454 (N_8454,N_7401,N_7024);
nor U8455 (N_8455,N_7109,N_7455);
nand U8456 (N_8456,N_7911,N_7461);
or U8457 (N_8457,N_7030,N_7469);
xnor U8458 (N_8458,N_7724,N_7236);
xnor U8459 (N_8459,N_7547,N_7506);
nor U8460 (N_8460,N_7056,N_7074);
xnor U8461 (N_8461,N_7616,N_7438);
nor U8462 (N_8462,N_7941,N_7084);
or U8463 (N_8463,N_7216,N_7768);
xor U8464 (N_8464,N_7036,N_7745);
or U8465 (N_8465,N_7906,N_7238);
xnor U8466 (N_8466,N_7380,N_7677);
xor U8467 (N_8467,N_7694,N_7541);
and U8468 (N_8468,N_7801,N_7328);
nand U8469 (N_8469,N_7360,N_7189);
nand U8470 (N_8470,N_7528,N_7698);
nand U8471 (N_8471,N_7138,N_7206);
or U8472 (N_8472,N_7770,N_7869);
nor U8473 (N_8473,N_7217,N_7382);
nor U8474 (N_8474,N_7755,N_7943);
nand U8475 (N_8475,N_7739,N_7025);
and U8476 (N_8476,N_7291,N_7226);
nor U8477 (N_8477,N_7520,N_7009);
or U8478 (N_8478,N_7757,N_7148);
nand U8479 (N_8479,N_7973,N_7270);
or U8480 (N_8480,N_7604,N_7201);
or U8481 (N_8481,N_7938,N_7609);
xnor U8482 (N_8482,N_7775,N_7059);
nand U8483 (N_8483,N_7097,N_7615);
and U8484 (N_8484,N_7509,N_7283);
and U8485 (N_8485,N_7245,N_7042);
nand U8486 (N_8486,N_7607,N_7809);
nor U8487 (N_8487,N_7623,N_7989);
nor U8488 (N_8488,N_7374,N_7225);
nand U8489 (N_8489,N_7638,N_7510);
and U8490 (N_8490,N_7013,N_7870);
or U8491 (N_8491,N_7390,N_7562);
or U8492 (N_8492,N_7356,N_7119);
and U8493 (N_8493,N_7833,N_7354);
and U8494 (N_8494,N_7769,N_7664);
and U8495 (N_8495,N_7857,N_7589);
nand U8496 (N_8496,N_7728,N_7823);
nand U8497 (N_8497,N_7844,N_7244);
and U8498 (N_8498,N_7369,N_7945);
nor U8499 (N_8499,N_7337,N_7126);
or U8500 (N_8500,N_7546,N_7393);
nand U8501 (N_8501,N_7016,N_7542);
and U8502 (N_8502,N_7765,N_7014);
nand U8503 (N_8503,N_7074,N_7874);
xnor U8504 (N_8504,N_7317,N_7247);
and U8505 (N_8505,N_7018,N_7316);
or U8506 (N_8506,N_7549,N_7747);
or U8507 (N_8507,N_7429,N_7306);
and U8508 (N_8508,N_7904,N_7940);
xor U8509 (N_8509,N_7096,N_7998);
or U8510 (N_8510,N_7379,N_7467);
nor U8511 (N_8511,N_7450,N_7139);
or U8512 (N_8512,N_7242,N_7871);
xor U8513 (N_8513,N_7121,N_7045);
nor U8514 (N_8514,N_7652,N_7191);
nand U8515 (N_8515,N_7861,N_7847);
xnor U8516 (N_8516,N_7618,N_7041);
nor U8517 (N_8517,N_7712,N_7440);
nand U8518 (N_8518,N_7492,N_7495);
and U8519 (N_8519,N_7973,N_7211);
or U8520 (N_8520,N_7707,N_7333);
or U8521 (N_8521,N_7600,N_7622);
or U8522 (N_8522,N_7737,N_7010);
and U8523 (N_8523,N_7992,N_7111);
or U8524 (N_8524,N_7493,N_7519);
nor U8525 (N_8525,N_7141,N_7246);
or U8526 (N_8526,N_7635,N_7091);
and U8527 (N_8527,N_7197,N_7635);
xnor U8528 (N_8528,N_7501,N_7128);
nor U8529 (N_8529,N_7847,N_7608);
nor U8530 (N_8530,N_7604,N_7029);
or U8531 (N_8531,N_7103,N_7251);
nor U8532 (N_8532,N_7197,N_7092);
and U8533 (N_8533,N_7373,N_7780);
and U8534 (N_8534,N_7817,N_7943);
nand U8535 (N_8535,N_7609,N_7210);
xnor U8536 (N_8536,N_7033,N_7886);
nor U8537 (N_8537,N_7050,N_7477);
or U8538 (N_8538,N_7906,N_7209);
nor U8539 (N_8539,N_7211,N_7739);
and U8540 (N_8540,N_7469,N_7027);
nor U8541 (N_8541,N_7269,N_7571);
nor U8542 (N_8542,N_7719,N_7694);
xnor U8543 (N_8543,N_7671,N_7675);
nor U8544 (N_8544,N_7601,N_7114);
or U8545 (N_8545,N_7553,N_7042);
nor U8546 (N_8546,N_7943,N_7701);
xnor U8547 (N_8547,N_7229,N_7585);
and U8548 (N_8548,N_7285,N_7095);
and U8549 (N_8549,N_7177,N_7724);
xor U8550 (N_8550,N_7121,N_7521);
nand U8551 (N_8551,N_7094,N_7068);
nand U8552 (N_8552,N_7471,N_7645);
and U8553 (N_8553,N_7075,N_7630);
and U8554 (N_8554,N_7481,N_7992);
or U8555 (N_8555,N_7046,N_7534);
or U8556 (N_8556,N_7742,N_7134);
and U8557 (N_8557,N_7002,N_7711);
xor U8558 (N_8558,N_7463,N_7496);
nand U8559 (N_8559,N_7216,N_7839);
nand U8560 (N_8560,N_7079,N_7274);
and U8561 (N_8561,N_7149,N_7412);
or U8562 (N_8562,N_7717,N_7264);
nand U8563 (N_8563,N_7673,N_7608);
or U8564 (N_8564,N_7531,N_7112);
nand U8565 (N_8565,N_7968,N_7579);
or U8566 (N_8566,N_7979,N_7607);
nor U8567 (N_8567,N_7381,N_7590);
and U8568 (N_8568,N_7698,N_7437);
nand U8569 (N_8569,N_7575,N_7881);
and U8570 (N_8570,N_7939,N_7872);
nor U8571 (N_8571,N_7465,N_7111);
and U8572 (N_8572,N_7534,N_7716);
nand U8573 (N_8573,N_7644,N_7287);
nor U8574 (N_8574,N_7288,N_7776);
and U8575 (N_8575,N_7263,N_7854);
nor U8576 (N_8576,N_7109,N_7144);
nand U8577 (N_8577,N_7268,N_7614);
nor U8578 (N_8578,N_7342,N_7422);
and U8579 (N_8579,N_7350,N_7173);
and U8580 (N_8580,N_7623,N_7948);
and U8581 (N_8581,N_7242,N_7270);
xnor U8582 (N_8582,N_7904,N_7630);
and U8583 (N_8583,N_7963,N_7855);
nand U8584 (N_8584,N_7236,N_7159);
or U8585 (N_8585,N_7112,N_7528);
nand U8586 (N_8586,N_7023,N_7425);
nor U8587 (N_8587,N_7840,N_7859);
nor U8588 (N_8588,N_7322,N_7002);
or U8589 (N_8589,N_7357,N_7329);
and U8590 (N_8590,N_7326,N_7536);
nand U8591 (N_8591,N_7450,N_7371);
nand U8592 (N_8592,N_7479,N_7982);
and U8593 (N_8593,N_7016,N_7322);
nor U8594 (N_8594,N_7664,N_7343);
and U8595 (N_8595,N_7402,N_7007);
or U8596 (N_8596,N_7756,N_7850);
or U8597 (N_8597,N_7691,N_7343);
nor U8598 (N_8598,N_7819,N_7890);
xor U8599 (N_8599,N_7015,N_7552);
and U8600 (N_8600,N_7116,N_7592);
or U8601 (N_8601,N_7421,N_7823);
or U8602 (N_8602,N_7931,N_7743);
nand U8603 (N_8603,N_7183,N_7096);
nand U8604 (N_8604,N_7252,N_7416);
nor U8605 (N_8605,N_7184,N_7475);
nor U8606 (N_8606,N_7923,N_7486);
or U8607 (N_8607,N_7310,N_7870);
and U8608 (N_8608,N_7870,N_7319);
and U8609 (N_8609,N_7345,N_7707);
and U8610 (N_8610,N_7859,N_7594);
nand U8611 (N_8611,N_7343,N_7875);
xnor U8612 (N_8612,N_7545,N_7413);
and U8613 (N_8613,N_7856,N_7634);
nand U8614 (N_8614,N_7428,N_7566);
and U8615 (N_8615,N_7075,N_7123);
xnor U8616 (N_8616,N_7490,N_7847);
nand U8617 (N_8617,N_7038,N_7986);
xor U8618 (N_8618,N_7823,N_7673);
xor U8619 (N_8619,N_7578,N_7778);
nand U8620 (N_8620,N_7612,N_7766);
nor U8621 (N_8621,N_7417,N_7817);
nor U8622 (N_8622,N_7615,N_7928);
xor U8623 (N_8623,N_7434,N_7129);
nand U8624 (N_8624,N_7563,N_7016);
and U8625 (N_8625,N_7268,N_7167);
and U8626 (N_8626,N_7494,N_7618);
nand U8627 (N_8627,N_7588,N_7856);
or U8628 (N_8628,N_7761,N_7454);
nand U8629 (N_8629,N_7690,N_7753);
nand U8630 (N_8630,N_7338,N_7696);
and U8631 (N_8631,N_7085,N_7386);
and U8632 (N_8632,N_7410,N_7050);
or U8633 (N_8633,N_7204,N_7214);
or U8634 (N_8634,N_7480,N_7292);
or U8635 (N_8635,N_7125,N_7295);
xnor U8636 (N_8636,N_7187,N_7952);
nor U8637 (N_8637,N_7362,N_7119);
and U8638 (N_8638,N_7291,N_7782);
nand U8639 (N_8639,N_7073,N_7149);
nor U8640 (N_8640,N_7540,N_7120);
nor U8641 (N_8641,N_7699,N_7025);
and U8642 (N_8642,N_7156,N_7643);
nor U8643 (N_8643,N_7105,N_7763);
nand U8644 (N_8644,N_7647,N_7161);
nand U8645 (N_8645,N_7997,N_7324);
or U8646 (N_8646,N_7149,N_7583);
or U8647 (N_8647,N_7396,N_7013);
and U8648 (N_8648,N_7124,N_7360);
nor U8649 (N_8649,N_7029,N_7302);
or U8650 (N_8650,N_7775,N_7937);
or U8651 (N_8651,N_7125,N_7782);
and U8652 (N_8652,N_7764,N_7981);
or U8653 (N_8653,N_7007,N_7144);
nand U8654 (N_8654,N_7650,N_7501);
nor U8655 (N_8655,N_7124,N_7659);
and U8656 (N_8656,N_7588,N_7401);
and U8657 (N_8657,N_7094,N_7116);
nor U8658 (N_8658,N_7117,N_7835);
nor U8659 (N_8659,N_7478,N_7660);
or U8660 (N_8660,N_7651,N_7254);
nor U8661 (N_8661,N_7032,N_7899);
xnor U8662 (N_8662,N_7958,N_7255);
xnor U8663 (N_8663,N_7634,N_7942);
nor U8664 (N_8664,N_7225,N_7584);
or U8665 (N_8665,N_7096,N_7251);
and U8666 (N_8666,N_7345,N_7450);
nand U8667 (N_8667,N_7840,N_7725);
nand U8668 (N_8668,N_7834,N_7185);
or U8669 (N_8669,N_7794,N_7912);
and U8670 (N_8670,N_7446,N_7616);
and U8671 (N_8671,N_7560,N_7924);
or U8672 (N_8672,N_7925,N_7513);
and U8673 (N_8673,N_7310,N_7880);
nand U8674 (N_8674,N_7826,N_7255);
nor U8675 (N_8675,N_7800,N_7967);
and U8676 (N_8676,N_7330,N_7625);
and U8677 (N_8677,N_7394,N_7074);
xnor U8678 (N_8678,N_7723,N_7726);
nand U8679 (N_8679,N_7809,N_7663);
nand U8680 (N_8680,N_7671,N_7244);
or U8681 (N_8681,N_7590,N_7834);
nor U8682 (N_8682,N_7221,N_7817);
and U8683 (N_8683,N_7978,N_7525);
or U8684 (N_8684,N_7896,N_7898);
nor U8685 (N_8685,N_7511,N_7550);
or U8686 (N_8686,N_7799,N_7425);
nand U8687 (N_8687,N_7223,N_7829);
and U8688 (N_8688,N_7130,N_7050);
nor U8689 (N_8689,N_7538,N_7822);
nor U8690 (N_8690,N_7907,N_7736);
and U8691 (N_8691,N_7960,N_7274);
or U8692 (N_8692,N_7199,N_7245);
and U8693 (N_8693,N_7194,N_7695);
and U8694 (N_8694,N_7528,N_7244);
nand U8695 (N_8695,N_7831,N_7027);
xor U8696 (N_8696,N_7147,N_7296);
or U8697 (N_8697,N_7015,N_7294);
and U8698 (N_8698,N_7336,N_7880);
or U8699 (N_8699,N_7844,N_7833);
nand U8700 (N_8700,N_7536,N_7567);
xnor U8701 (N_8701,N_7730,N_7925);
xnor U8702 (N_8702,N_7344,N_7371);
nand U8703 (N_8703,N_7537,N_7154);
or U8704 (N_8704,N_7519,N_7037);
nand U8705 (N_8705,N_7394,N_7496);
and U8706 (N_8706,N_7282,N_7651);
and U8707 (N_8707,N_7850,N_7362);
nor U8708 (N_8708,N_7194,N_7046);
or U8709 (N_8709,N_7557,N_7937);
nand U8710 (N_8710,N_7880,N_7244);
or U8711 (N_8711,N_7563,N_7874);
or U8712 (N_8712,N_7570,N_7115);
and U8713 (N_8713,N_7114,N_7705);
nor U8714 (N_8714,N_7558,N_7428);
or U8715 (N_8715,N_7891,N_7230);
nand U8716 (N_8716,N_7431,N_7122);
nor U8717 (N_8717,N_7132,N_7567);
nor U8718 (N_8718,N_7116,N_7863);
nand U8719 (N_8719,N_7583,N_7454);
and U8720 (N_8720,N_7105,N_7221);
or U8721 (N_8721,N_7972,N_7773);
nor U8722 (N_8722,N_7362,N_7159);
and U8723 (N_8723,N_7788,N_7444);
and U8724 (N_8724,N_7917,N_7022);
nand U8725 (N_8725,N_7788,N_7819);
nand U8726 (N_8726,N_7052,N_7761);
nand U8727 (N_8727,N_7025,N_7632);
or U8728 (N_8728,N_7508,N_7526);
or U8729 (N_8729,N_7463,N_7891);
and U8730 (N_8730,N_7586,N_7372);
nor U8731 (N_8731,N_7623,N_7895);
or U8732 (N_8732,N_7596,N_7368);
or U8733 (N_8733,N_7956,N_7241);
and U8734 (N_8734,N_7268,N_7615);
nand U8735 (N_8735,N_7543,N_7801);
or U8736 (N_8736,N_7928,N_7997);
or U8737 (N_8737,N_7905,N_7348);
nand U8738 (N_8738,N_7605,N_7752);
nand U8739 (N_8739,N_7594,N_7461);
xnor U8740 (N_8740,N_7604,N_7341);
or U8741 (N_8741,N_7090,N_7371);
and U8742 (N_8742,N_7368,N_7490);
and U8743 (N_8743,N_7424,N_7004);
xor U8744 (N_8744,N_7324,N_7458);
or U8745 (N_8745,N_7304,N_7517);
nand U8746 (N_8746,N_7804,N_7186);
nor U8747 (N_8747,N_7632,N_7021);
and U8748 (N_8748,N_7597,N_7608);
or U8749 (N_8749,N_7854,N_7296);
or U8750 (N_8750,N_7249,N_7883);
and U8751 (N_8751,N_7021,N_7852);
xnor U8752 (N_8752,N_7495,N_7177);
nand U8753 (N_8753,N_7088,N_7234);
and U8754 (N_8754,N_7217,N_7954);
or U8755 (N_8755,N_7775,N_7852);
nor U8756 (N_8756,N_7657,N_7739);
or U8757 (N_8757,N_7461,N_7663);
nand U8758 (N_8758,N_7295,N_7296);
and U8759 (N_8759,N_7549,N_7778);
nor U8760 (N_8760,N_7734,N_7299);
nand U8761 (N_8761,N_7180,N_7024);
xnor U8762 (N_8762,N_7269,N_7982);
nor U8763 (N_8763,N_7826,N_7984);
nand U8764 (N_8764,N_7807,N_7733);
nand U8765 (N_8765,N_7041,N_7258);
nor U8766 (N_8766,N_7479,N_7292);
nor U8767 (N_8767,N_7025,N_7191);
nand U8768 (N_8768,N_7146,N_7674);
or U8769 (N_8769,N_7814,N_7053);
nand U8770 (N_8770,N_7278,N_7536);
and U8771 (N_8771,N_7915,N_7849);
xor U8772 (N_8772,N_7771,N_7894);
nand U8773 (N_8773,N_7385,N_7303);
nor U8774 (N_8774,N_7780,N_7430);
xor U8775 (N_8775,N_7844,N_7548);
or U8776 (N_8776,N_7369,N_7246);
xor U8777 (N_8777,N_7940,N_7659);
or U8778 (N_8778,N_7378,N_7046);
nand U8779 (N_8779,N_7267,N_7062);
or U8780 (N_8780,N_7996,N_7282);
nand U8781 (N_8781,N_7396,N_7196);
or U8782 (N_8782,N_7220,N_7763);
or U8783 (N_8783,N_7855,N_7041);
or U8784 (N_8784,N_7214,N_7461);
nand U8785 (N_8785,N_7279,N_7666);
and U8786 (N_8786,N_7512,N_7193);
nor U8787 (N_8787,N_7136,N_7388);
and U8788 (N_8788,N_7819,N_7396);
nand U8789 (N_8789,N_7860,N_7711);
or U8790 (N_8790,N_7674,N_7661);
or U8791 (N_8791,N_7659,N_7317);
nand U8792 (N_8792,N_7768,N_7439);
nand U8793 (N_8793,N_7530,N_7826);
nand U8794 (N_8794,N_7083,N_7915);
or U8795 (N_8795,N_7750,N_7386);
nor U8796 (N_8796,N_7454,N_7604);
xnor U8797 (N_8797,N_7268,N_7108);
or U8798 (N_8798,N_7040,N_7048);
or U8799 (N_8799,N_7697,N_7056);
and U8800 (N_8800,N_7187,N_7869);
nand U8801 (N_8801,N_7117,N_7899);
nor U8802 (N_8802,N_7461,N_7393);
or U8803 (N_8803,N_7974,N_7523);
xnor U8804 (N_8804,N_7845,N_7361);
nand U8805 (N_8805,N_7297,N_7055);
or U8806 (N_8806,N_7427,N_7167);
and U8807 (N_8807,N_7166,N_7104);
nor U8808 (N_8808,N_7031,N_7378);
or U8809 (N_8809,N_7955,N_7453);
or U8810 (N_8810,N_7649,N_7600);
or U8811 (N_8811,N_7143,N_7665);
or U8812 (N_8812,N_7846,N_7443);
and U8813 (N_8813,N_7487,N_7863);
or U8814 (N_8814,N_7812,N_7140);
nand U8815 (N_8815,N_7404,N_7422);
and U8816 (N_8816,N_7594,N_7944);
or U8817 (N_8817,N_7746,N_7064);
and U8818 (N_8818,N_7999,N_7445);
or U8819 (N_8819,N_7502,N_7862);
nand U8820 (N_8820,N_7790,N_7093);
nand U8821 (N_8821,N_7524,N_7867);
nor U8822 (N_8822,N_7765,N_7744);
or U8823 (N_8823,N_7879,N_7401);
xnor U8824 (N_8824,N_7801,N_7034);
or U8825 (N_8825,N_7406,N_7448);
or U8826 (N_8826,N_7397,N_7354);
or U8827 (N_8827,N_7191,N_7941);
xnor U8828 (N_8828,N_7048,N_7279);
and U8829 (N_8829,N_7112,N_7271);
nand U8830 (N_8830,N_7925,N_7026);
nor U8831 (N_8831,N_7714,N_7741);
or U8832 (N_8832,N_7875,N_7045);
nor U8833 (N_8833,N_7856,N_7784);
nor U8834 (N_8834,N_7515,N_7782);
nand U8835 (N_8835,N_7010,N_7352);
and U8836 (N_8836,N_7288,N_7635);
nor U8837 (N_8837,N_7473,N_7156);
nor U8838 (N_8838,N_7923,N_7518);
nand U8839 (N_8839,N_7070,N_7927);
and U8840 (N_8840,N_7590,N_7264);
or U8841 (N_8841,N_7189,N_7785);
and U8842 (N_8842,N_7881,N_7025);
and U8843 (N_8843,N_7476,N_7123);
or U8844 (N_8844,N_7479,N_7236);
xnor U8845 (N_8845,N_7751,N_7029);
or U8846 (N_8846,N_7460,N_7872);
nor U8847 (N_8847,N_7823,N_7190);
or U8848 (N_8848,N_7234,N_7582);
and U8849 (N_8849,N_7021,N_7836);
nand U8850 (N_8850,N_7185,N_7361);
nand U8851 (N_8851,N_7327,N_7990);
and U8852 (N_8852,N_7111,N_7810);
and U8853 (N_8853,N_7167,N_7151);
or U8854 (N_8854,N_7189,N_7657);
or U8855 (N_8855,N_7500,N_7793);
xnor U8856 (N_8856,N_7571,N_7010);
nor U8857 (N_8857,N_7559,N_7931);
and U8858 (N_8858,N_7924,N_7890);
or U8859 (N_8859,N_7405,N_7625);
nand U8860 (N_8860,N_7724,N_7358);
nand U8861 (N_8861,N_7924,N_7043);
xor U8862 (N_8862,N_7020,N_7489);
and U8863 (N_8863,N_7495,N_7002);
nand U8864 (N_8864,N_7996,N_7584);
nor U8865 (N_8865,N_7689,N_7413);
nand U8866 (N_8866,N_7090,N_7655);
nand U8867 (N_8867,N_7563,N_7679);
nor U8868 (N_8868,N_7870,N_7171);
nor U8869 (N_8869,N_7672,N_7285);
or U8870 (N_8870,N_7894,N_7066);
nand U8871 (N_8871,N_7033,N_7699);
nand U8872 (N_8872,N_7638,N_7927);
nor U8873 (N_8873,N_7038,N_7112);
and U8874 (N_8874,N_7314,N_7696);
nor U8875 (N_8875,N_7887,N_7400);
or U8876 (N_8876,N_7138,N_7691);
and U8877 (N_8877,N_7820,N_7946);
or U8878 (N_8878,N_7913,N_7877);
and U8879 (N_8879,N_7547,N_7797);
nand U8880 (N_8880,N_7662,N_7842);
and U8881 (N_8881,N_7018,N_7089);
nor U8882 (N_8882,N_7655,N_7990);
nand U8883 (N_8883,N_7152,N_7871);
or U8884 (N_8884,N_7211,N_7771);
nand U8885 (N_8885,N_7473,N_7236);
nand U8886 (N_8886,N_7647,N_7121);
or U8887 (N_8887,N_7244,N_7608);
or U8888 (N_8888,N_7854,N_7478);
or U8889 (N_8889,N_7624,N_7159);
and U8890 (N_8890,N_7370,N_7569);
xnor U8891 (N_8891,N_7369,N_7814);
nor U8892 (N_8892,N_7385,N_7731);
and U8893 (N_8893,N_7849,N_7431);
or U8894 (N_8894,N_7612,N_7626);
xnor U8895 (N_8895,N_7337,N_7247);
and U8896 (N_8896,N_7143,N_7467);
nand U8897 (N_8897,N_7255,N_7905);
nor U8898 (N_8898,N_7455,N_7732);
and U8899 (N_8899,N_7918,N_7748);
nand U8900 (N_8900,N_7052,N_7886);
and U8901 (N_8901,N_7941,N_7816);
and U8902 (N_8902,N_7388,N_7497);
or U8903 (N_8903,N_7755,N_7929);
and U8904 (N_8904,N_7080,N_7167);
and U8905 (N_8905,N_7217,N_7014);
or U8906 (N_8906,N_7534,N_7793);
or U8907 (N_8907,N_7768,N_7228);
xnor U8908 (N_8908,N_7554,N_7694);
or U8909 (N_8909,N_7196,N_7167);
nor U8910 (N_8910,N_7319,N_7108);
nor U8911 (N_8911,N_7970,N_7626);
and U8912 (N_8912,N_7048,N_7510);
xor U8913 (N_8913,N_7728,N_7735);
xor U8914 (N_8914,N_7817,N_7304);
or U8915 (N_8915,N_7150,N_7872);
nor U8916 (N_8916,N_7508,N_7386);
xnor U8917 (N_8917,N_7405,N_7834);
nor U8918 (N_8918,N_7614,N_7673);
xor U8919 (N_8919,N_7350,N_7754);
nor U8920 (N_8920,N_7625,N_7346);
nor U8921 (N_8921,N_7400,N_7310);
nand U8922 (N_8922,N_7547,N_7055);
nand U8923 (N_8923,N_7299,N_7174);
nand U8924 (N_8924,N_7283,N_7424);
nor U8925 (N_8925,N_7596,N_7053);
nand U8926 (N_8926,N_7742,N_7369);
and U8927 (N_8927,N_7062,N_7282);
nand U8928 (N_8928,N_7240,N_7620);
and U8929 (N_8929,N_7198,N_7970);
xnor U8930 (N_8930,N_7067,N_7443);
or U8931 (N_8931,N_7976,N_7781);
nand U8932 (N_8932,N_7313,N_7869);
nand U8933 (N_8933,N_7176,N_7879);
or U8934 (N_8934,N_7073,N_7580);
nor U8935 (N_8935,N_7325,N_7044);
and U8936 (N_8936,N_7582,N_7538);
nand U8937 (N_8937,N_7577,N_7797);
nor U8938 (N_8938,N_7919,N_7187);
nor U8939 (N_8939,N_7518,N_7244);
nor U8940 (N_8940,N_7097,N_7088);
nor U8941 (N_8941,N_7584,N_7975);
nor U8942 (N_8942,N_7180,N_7020);
xnor U8943 (N_8943,N_7592,N_7511);
or U8944 (N_8944,N_7729,N_7413);
or U8945 (N_8945,N_7246,N_7041);
nand U8946 (N_8946,N_7203,N_7928);
nor U8947 (N_8947,N_7366,N_7405);
nor U8948 (N_8948,N_7222,N_7980);
and U8949 (N_8949,N_7560,N_7201);
nor U8950 (N_8950,N_7896,N_7221);
nand U8951 (N_8951,N_7706,N_7871);
nor U8952 (N_8952,N_7177,N_7973);
nor U8953 (N_8953,N_7211,N_7574);
xor U8954 (N_8954,N_7098,N_7185);
and U8955 (N_8955,N_7976,N_7162);
or U8956 (N_8956,N_7592,N_7633);
nand U8957 (N_8957,N_7084,N_7847);
nor U8958 (N_8958,N_7083,N_7137);
or U8959 (N_8959,N_7951,N_7841);
and U8960 (N_8960,N_7795,N_7362);
nor U8961 (N_8961,N_7401,N_7793);
and U8962 (N_8962,N_7148,N_7427);
and U8963 (N_8963,N_7154,N_7502);
nor U8964 (N_8964,N_7596,N_7636);
xor U8965 (N_8965,N_7330,N_7708);
nand U8966 (N_8966,N_7069,N_7348);
and U8967 (N_8967,N_7951,N_7701);
nor U8968 (N_8968,N_7093,N_7020);
and U8969 (N_8969,N_7683,N_7900);
and U8970 (N_8970,N_7819,N_7871);
nand U8971 (N_8971,N_7221,N_7475);
nand U8972 (N_8972,N_7460,N_7790);
nor U8973 (N_8973,N_7304,N_7887);
nor U8974 (N_8974,N_7347,N_7838);
and U8975 (N_8975,N_7272,N_7488);
nor U8976 (N_8976,N_7762,N_7166);
and U8977 (N_8977,N_7295,N_7319);
xnor U8978 (N_8978,N_7187,N_7349);
or U8979 (N_8979,N_7002,N_7971);
nor U8980 (N_8980,N_7066,N_7573);
or U8981 (N_8981,N_7186,N_7488);
nand U8982 (N_8982,N_7362,N_7648);
or U8983 (N_8983,N_7135,N_7864);
nor U8984 (N_8984,N_7084,N_7268);
nand U8985 (N_8985,N_7257,N_7017);
or U8986 (N_8986,N_7357,N_7695);
and U8987 (N_8987,N_7838,N_7457);
nand U8988 (N_8988,N_7441,N_7319);
nand U8989 (N_8989,N_7063,N_7057);
nor U8990 (N_8990,N_7751,N_7606);
and U8991 (N_8991,N_7550,N_7525);
nand U8992 (N_8992,N_7473,N_7183);
nand U8993 (N_8993,N_7919,N_7066);
or U8994 (N_8994,N_7017,N_7735);
or U8995 (N_8995,N_7677,N_7726);
and U8996 (N_8996,N_7294,N_7942);
or U8997 (N_8997,N_7791,N_7148);
and U8998 (N_8998,N_7483,N_7827);
nor U8999 (N_8999,N_7281,N_7185);
nand U9000 (N_9000,N_8509,N_8498);
or U9001 (N_9001,N_8315,N_8520);
and U9002 (N_9002,N_8206,N_8596);
nor U9003 (N_9003,N_8467,N_8199);
xor U9004 (N_9004,N_8667,N_8378);
and U9005 (N_9005,N_8502,N_8601);
and U9006 (N_9006,N_8176,N_8203);
and U9007 (N_9007,N_8582,N_8974);
nand U9008 (N_9008,N_8134,N_8123);
nand U9009 (N_9009,N_8441,N_8468);
or U9010 (N_9010,N_8487,N_8102);
nor U9011 (N_9011,N_8618,N_8141);
and U9012 (N_9012,N_8617,N_8299);
xnor U9013 (N_9013,N_8595,N_8615);
or U9014 (N_9014,N_8774,N_8685);
or U9015 (N_9015,N_8218,N_8909);
nand U9016 (N_9016,N_8439,N_8513);
xor U9017 (N_9017,N_8651,N_8319);
and U9018 (N_9018,N_8503,N_8827);
and U9019 (N_9019,N_8526,N_8122);
xnor U9020 (N_9020,N_8566,N_8172);
nand U9021 (N_9021,N_8057,N_8668);
nor U9022 (N_9022,N_8627,N_8769);
or U9023 (N_9023,N_8935,N_8921);
xor U9024 (N_9024,N_8383,N_8939);
or U9025 (N_9025,N_8585,N_8320);
or U9026 (N_9026,N_8519,N_8648);
xnor U9027 (N_9027,N_8281,N_8660);
and U9028 (N_9028,N_8340,N_8157);
xnor U9029 (N_9029,N_8870,N_8525);
and U9030 (N_9030,N_8204,N_8738);
and U9031 (N_9031,N_8599,N_8308);
nor U9032 (N_9032,N_8830,N_8094);
nor U9033 (N_9033,N_8722,N_8676);
or U9034 (N_9034,N_8592,N_8112);
nor U9035 (N_9035,N_8014,N_8765);
or U9036 (N_9036,N_8611,N_8273);
nor U9037 (N_9037,N_8540,N_8843);
xnor U9038 (N_9038,N_8543,N_8715);
nand U9039 (N_9039,N_8853,N_8705);
xnor U9040 (N_9040,N_8028,N_8198);
or U9041 (N_9041,N_8449,N_8817);
or U9042 (N_9042,N_8524,N_8781);
nor U9043 (N_9043,N_8447,N_8174);
and U9044 (N_9044,N_8753,N_8576);
or U9045 (N_9045,N_8614,N_8744);
and U9046 (N_9046,N_8026,N_8532);
nand U9047 (N_9047,N_8562,N_8456);
and U9048 (N_9048,N_8200,N_8868);
nand U9049 (N_9049,N_8162,N_8160);
nor U9050 (N_9050,N_8878,N_8838);
nor U9051 (N_9051,N_8401,N_8732);
or U9052 (N_9052,N_8042,N_8326);
nand U9053 (N_9053,N_8314,N_8077);
and U9054 (N_9054,N_8953,N_8686);
or U9055 (N_9055,N_8457,N_8871);
nand U9056 (N_9056,N_8922,N_8081);
or U9057 (N_9057,N_8171,N_8639);
xnor U9058 (N_9058,N_8849,N_8716);
and U9059 (N_9059,N_8496,N_8404);
nor U9060 (N_9060,N_8644,N_8995);
and U9061 (N_9061,N_8891,N_8548);
or U9062 (N_9062,N_8845,N_8850);
nand U9063 (N_9063,N_8772,N_8387);
nand U9064 (N_9064,N_8947,N_8733);
nand U9065 (N_9065,N_8445,N_8504);
or U9066 (N_9066,N_8636,N_8580);
or U9067 (N_9067,N_8183,N_8139);
nor U9068 (N_9068,N_8969,N_8224);
or U9069 (N_9069,N_8279,N_8377);
and U9070 (N_9070,N_8034,N_8285);
nor U9071 (N_9071,N_8129,N_8235);
and U9072 (N_9072,N_8393,N_8675);
or U9073 (N_9073,N_8429,N_8723);
or U9074 (N_9074,N_8238,N_8666);
or U9075 (N_9075,N_8215,N_8254);
and U9076 (N_9076,N_8142,N_8926);
and U9077 (N_9077,N_8563,N_8937);
and U9078 (N_9078,N_8180,N_8929);
and U9079 (N_9079,N_8262,N_8444);
or U9080 (N_9080,N_8284,N_8465);
or U9081 (N_9081,N_8464,N_8770);
and U9082 (N_9082,N_8343,N_8653);
nor U9083 (N_9083,N_8328,N_8622);
nand U9084 (N_9084,N_8571,N_8763);
nor U9085 (N_9085,N_8434,N_8084);
nor U9086 (N_9086,N_8471,N_8346);
xnor U9087 (N_9087,N_8096,N_8036);
xor U9088 (N_9088,N_8414,N_8810);
nor U9089 (N_9089,N_8996,N_8743);
nor U9090 (N_9090,N_8016,N_8248);
nand U9091 (N_9091,N_8261,N_8448);
or U9092 (N_9092,N_8641,N_8071);
nand U9093 (N_9093,N_8957,N_8597);
nor U9094 (N_9094,N_8435,N_8181);
nand U9095 (N_9095,N_8135,N_8959);
nor U9096 (N_9096,N_8395,N_8373);
or U9097 (N_9097,N_8984,N_8438);
nand U9098 (N_9098,N_8230,N_8428);
and U9099 (N_9099,N_8606,N_8100);
or U9100 (N_9100,N_8133,N_8777);
or U9101 (N_9101,N_8758,N_8820);
and U9102 (N_9102,N_8334,N_8593);
nand U9103 (N_9103,N_8126,N_8903);
nand U9104 (N_9104,N_8874,N_8952);
nand U9105 (N_9105,N_8547,N_8250);
nand U9106 (N_9106,N_8745,N_8397);
nor U9107 (N_9107,N_8313,N_8083);
nor U9108 (N_9108,N_8523,N_8251);
xor U9109 (N_9109,N_8815,N_8053);
and U9110 (N_9110,N_8054,N_8494);
or U9111 (N_9111,N_8389,N_8229);
xnor U9112 (N_9112,N_8915,N_8099);
nor U9113 (N_9113,N_8460,N_8741);
or U9114 (N_9114,N_8259,N_8792);
nand U9115 (N_9115,N_8073,N_8689);
or U9116 (N_9116,N_8029,N_8746);
nand U9117 (N_9117,N_8747,N_8185);
nand U9118 (N_9118,N_8706,N_8872);
nand U9119 (N_9119,N_8294,N_8293);
and U9120 (N_9120,N_8092,N_8799);
or U9121 (N_9121,N_8696,N_8749);
nor U9122 (N_9122,N_8633,N_8040);
xnor U9123 (N_9123,N_8304,N_8784);
nor U9124 (N_9124,N_8078,N_8537);
xnor U9125 (N_9125,N_8316,N_8234);
nand U9126 (N_9126,N_8156,N_8275);
or U9127 (N_9127,N_8702,N_8737);
and U9128 (N_9128,N_8348,N_8193);
or U9129 (N_9129,N_8158,N_8413);
xor U9130 (N_9130,N_8466,N_8037);
or U9131 (N_9131,N_8086,N_8165);
nor U9132 (N_9132,N_8347,N_8219);
and U9133 (N_9133,N_8545,N_8754);
nor U9134 (N_9134,N_8202,N_8717);
or U9135 (N_9135,N_8662,N_8088);
nand U9136 (N_9136,N_8698,N_8842);
nor U9137 (N_9137,N_8361,N_8453);
nor U9138 (N_9138,N_8881,N_8865);
or U9139 (N_9139,N_8568,N_8610);
nand U9140 (N_9140,N_8479,N_8298);
nor U9141 (N_9141,N_8296,N_8282);
nor U9142 (N_9142,N_8712,N_8327);
and U9143 (N_9143,N_8768,N_8803);
nand U9144 (N_9144,N_8427,N_8860);
or U9145 (N_9145,N_8007,N_8694);
nor U9146 (N_9146,N_8458,N_8687);
and U9147 (N_9147,N_8551,N_8679);
or U9148 (N_9148,N_8927,N_8398);
or U9149 (N_9149,N_8791,N_8958);
nand U9150 (N_9150,N_8127,N_8128);
nor U9151 (N_9151,N_8267,N_8629);
and U9152 (N_9152,N_8677,N_8965);
and U9153 (N_9153,N_8039,N_8533);
and U9154 (N_9154,N_8191,N_8242);
or U9155 (N_9155,N_8473,N_8538);
or U9156 (N_9156,N_8474,N_8748);
nand U9157 (N_9157,N_8020,N_8031);
xor U9158 (N_9158,N_8276,N_8925);
or U9159 (N_9159,N_8938,N_8011);
nand U9160 (N_9160,N_8883,N_8443);
and U9161 (N_9161,N_8528,N_8064);
nand U9162 (N_9162,N_8659,N_8167);
nor U9163 (N_9163,N_8661,N_8233);
nor U9164 (N_9164,N_8977,N_8987);
nand U9165 (N_9165,N_8402,N_8944);
and U9166 (N_9166,N_8833,N_8518);
or U9167 (N_9167,N_8998,N_8151);
nor U9168 (N_9168,N_8982,N_8895);
or U9169 (N_9169,N_8650,N_8249);
xnor U9170 (N_9170,N_8381,N_8756);
xnor U9171 (N_9171,N_8501,N_8634);
and U9172 (N_9172,N_8119,N_8352);
nor U9173 (N_9173,N_8796,N_8022);
nand U9174 (N_9174,N_8695,N_8762);
and U9175 (N_9175,N_8517,N_8683);
and U9176 (N_9176,N_8153,N_8412);
nand U9177 (N_9177,N_8417,N_8840);
or U9178 (N_9178,N_8055,N_8385);
nor U9179 (N_9179,N_8409,N_8400);
nor U9180 (N_9180,N_8967,N_8931);
xnor U9181 (N_9181,N_8056,N_8673);
nor U9182 (N_9182,N_8554,N_8709);
nor U9183 (N_9183,N_8452,N_8900);
or U9184 (N_9184,N_8638,N_8589);
and U9185 (N_9185,N_8300,N_8557);
nand U9186 (N_9186,N_8310,N_8463);
nand U9187 (N_9187,N_8530,N_8970);
and U9188 (N_9188,N_8258,N_8396);
nor U9189 (N_9189,N_8047,N_8424);
and U9190 (N_9190,N_8188,N_8560);
and U9191 (N_9191,N_8800,N_8701);
or U9192 (N_9192,N_8069,N_8368);
or U9193 (N_9193,N_8577,N_8643);
and U9194 (N_9194,N_8236,N_8207);
nand U9195 (N_9195,N_8573,N_8270);
nand U9196 (N_9196,N_8008,N_8063);
and U9197 (N_9197,N_8949,N_8898);
or U9198 (N_9198,N_8472,N_8693);
nor U9199 (N_9199,N_8149,N_8090);
nand U9200 (N_9200,N_8807,N_8834);
nand U9201 (N_9201,N_8164,N_8710);
nor U9202 (N_9202,N_8121,N_8943);
nor U9203 (N_9203,N_8681,N_8887);
or U9204 (N_9204,N_8354,N_8866);
and U9205 (N_9205,N_8355,N_8642);
nand U9206 (N_9206,N_8357,N_8613);
nand U9207 (N_9207,N_8060,N_8936);
or U9208 (N_9208,N_8671,N_8425);
and U9209 (N_9209,N_8836,N_8535);
and U9210 (N_9210,N_8682,N_8721);
nand U9211 (N_9211,N_8621,N_8835);
nand U9212 (N_9212,N_8363,N_8110);
and U9213 (N_9213,N_8497,N_8893);
and U9214 (N_9214,N_8814,N_8885);
nand U9215 (N_9215,N_8286,N_8801);
nor U9216 (N_9216,N_8844,N_8522);
xnor U9217 (N_9217,N_8358,N_8990);
or U9218 (N_9218,N_8773,N_8038);
and U9219 (N_9219,N_8244,N_8052);
xor U9220 (N_9220,N_8306,N_8812);
nand U9221 (N_9221,N_8684,N_8002);
xnor U9222 (N_9222,N_8272,N_8217);
and U9223 (N_9223,N_8163,N_8075);
or U9224 (N_9224,N_8558,N_8231);
or U9225 (N_9225,N_8266,N_8044);
and U9226 (N_9226,N_8534,N_8764);
and U9227 (N_9227,N_8109,N_8976);
nor U9228 (N_9228,N_8362,N_8000);
xnor U9229 (N_9229,N_8919,N_8003);
nand U9230 (N_9230,N_8718,N_8894);
xnor U9231 (N_9231,N_8051,N_8486);
nor U9232 (N_9232,N_8742,N_8116);
and U9233 (N_9233,N_8968,N_8041);
nand U9234 (N_9234,N_8847,N_8674);
or U9235 (N_9235,N_8901,N_8461);
nor U9236 (N_9236,N_8019,N_8050);
or U9237 (N_9237,N_8418,N_8113);
or U9238 (N_9238,N_8818,N_8107);
nor U9239 (N_9239,N_8988,N_8212);
or U9240 (N_9240,N_8783,N_8731);
nand U9241 (N_9241,N_8735,N_8946);
nand U9242 (N_9242,N_8336,N_8980);
or U9243 (N_9243,N_8391,N_8205);
and U9244 (N_9244,N_8291,N_8423);
nor U9245 (N_9245,N_8646,N_8290);
or U9246 (N_9246,N_8906,N_8469);
or U9247 (N_9247,N_8154,N_8345);
and U9248 (N_9248,N_8657,N_8567);
nor U9249 (N_9249,N_8059,N_8822);
nor U9250 (N_9250,N_8572,N_8225);
or U9251 (N_9251,N_8410,N_8076);
nand U9252 (N_9252,N_8546,N_8432);
nand U9253 (N_9253,N_8370,N_8095);
nand U9254 (N_9254,N_8208,N_8426);
nand U9255 (N_9255,N_8280,N_8147);
and U9256 (N_9256,N_8979,N_8321);
and U9257 (N_9257,N_8416,N_8030);
nor U9258 (N_9258,N_8899,N_8260);
nand U9259 (N_9259,N_8570,N_8852);
nor U9260 (N_9260,N_8691,N_8975);
nand U9261 (N_9261,N_8337,N_8697);
or U9262 (N_9262,N_8612,N_8405);
nand U9263 (N_9263,N_8776,N_8986);
nand U9264 (N_9264,N_8117,N_8655);
and U9265 (N_9265,N_8159,N_8954);
or U9266 (N_9266,N_8161,N_8289);
nor U9267 (N_9267,N_8263,N_8480);
and U9268 (N_9268,N_8455,N_8879);
or U9269 (N_9269,N_8569,N_8483);
and U9270 (N_9270,N_8910,N_8484);
xnor U9271 (N_9271,N_8598,N_8018);
nand U9272 (N_9272,N_8148,N_8928);
nor U9273 (N_9273,N_8588,N_8714);
and U9274 (N_9274,N_8492,N_8010);
xor U9275 (N_9275,N_8993,N_8009);
and U9276 (N_9276,N_8024,N_8491);
nand U9277 (N_9277,N_8415,N_8325);
nand U9278 (N_9278,N_8097,N_8854);
nor U9279 (N_9279,N_8145,N_8583);
nor U9280 (N_9280,N_8933,N_8561);
and U9281 (N_9281,N_8072,N_8004);
xnor U9282 (N_9282,N_8876,N_8670);
nor U9283 (N_9283,N_8364,N_8708);
nand U9284 (N_9284,N_8246,N_8816);
or U9285 (N_9285,N_8353,N_8278);
nand U9286 (N_9286,N_8788,N_8992);
or U9287 (N_9287,N_8237,N_8292);
nor U9288 (N_9288,N_8515,N_8759);
nor U9289 (N_9289,N_8586,N_8727);
xor U9290 (N_9290,N_8924,N_8283);
and U9291 (N_9291,N_8640,N_8440);
nor U9292 (N_9292,N_8376,N_8195);
nor U9293 (N_9293,N_8608,N_8374);
nor U9294 (N_9294,N_8948,N_8837);
and U9295 (N_9295,N_8902,N_8062);
nor U9296 (N_9296,N_8889,N_8529);
or U9297 (N_9297,N_8779,N_8859);
xor U9298 (N_9298,N_8755,N_8940);
nand U9299 (N_9299,N_8624,N_8918);
nor U9300 (N_9300,N_8690,N_8856);
nor U9301 (N_9301,N_8809,N_8602);
nor U9302 (N_9302,N_8239,N_8493);
nand U9303 (N_9303,N_8170,N_8350);
nand U9304 (N_9304,N_8625,N_8322);
and U9305 (N_9305,N_8584,N_8462);
or U9306 (N_9306,N_8407,N_8521);
xor U9307 (N_9307,N_8600,N_8136);
nor U9308 (N_9308,N_8390,N_8678);
or U9309 (N_9309,N_8297,N_8553);
nand U9310 (N_9310,N_8507,N_8228);
or U9311 (N_9311,N_8963,N_8317);
or U9312 (N_9312,N_8399,N_8032);
or U9313 (N_9313,N_8620,N_8371);
nand U9314 (N_9314,N_8761,N_8305);
and U9315 (N_9315,N_8021,N_8005);
nor U9316 (N_9316,N_8500,N_8880);
nor U9317 (N_9317,N_8475,N_8630);
xor U9318 (N_9318,N_8531,N_8911);
or U9319 (N_9319,N_8711,N_8851);
or U9320 (N_9320,N_8861,N_8826);
nand U9321 (N_9321,N_8961,N_8813);
or U9322 (N_9322,N_8966,N_8632);
nand U9323 (N_9323,N_8130,N_8672);
or U9324 (N_9324,N_8780,N_8999);
xnor U9325 (N_9325,N_8489,N_8908);
and U9326 (N_9326,N_8105,N_8559);
or U9327 (N_9327,N_8027,N_8386);
nand U9328 (N_9328,N_8067,N_8221);
nand U9329 (N_9329,N_8912,N_8828);
or U9330 (N_9330,N_8775,N_8477);
nor U9331 (N_9331,N_8594,N_8506);
nor U9332 (N_9332,N_8823,N_8066);
nand U9333 (N_9333,N_8581,N_8408);
nor U9334 (N_9334,N_8886,N_8647);
xor U9335 (N_9335,N_8790,N_8144);
nor U9336 (N_9336,N_8339,N_8983);
or U9337 (N_9337,N_8247,N_8210);
nand U9338 (N_9338,N_8527,N_8307);
and U9339 (N_9339,N_8025,N_8956);
nor U9340 (N_9340,N_8649,N_8544);
nand U9341 (N_9341,N_8349,N_8365);
nand U9342 (N_9342,N_8132,N_8725);
nand U9343 (N_9343,N_8274,N_8446);
or U9344 (N_9344,N_8825,N_8541);
or U9345 (N_9345,N_8867,N_8587);
nand U9346 (N_9346,N_8771,N_8512);
nand U9347 (N_9347,N_8227,N_8795);
and U9348 (N_9348,N_8369,N_8819);
nand U9349 (N_9349,N_8539,N_8451);
xor U9350 (N_9350,N_8245,N_8726);
or U9351 (N_9351,N_8431,N_8955);
nand U9352 (N_9352,N_8991,N_8888);
or U9353 (N_9353,N_8388,N_8190);
nand U9354 (N_9354,N_8394,N_8663);
and U9355 (N_9355,N_8150,N_8216);
and U9356 (N_9356,N_8068,N_8751);
or U9357 (N_9357,N_8222,N_8536);
nor U9358 (N_9358,N_8579,N_8516);
and U9359 (N_9359,N_8877,N_8108);
xor U9360 (N_9360,N_8923,N_8740);
and U9361 (N_9361,N_8436,N_8897);
or U9362 (N_9362,N_8971,N_8973);
and U9363 (N_9363,N_8688,N_8137);
or U9364 (N_9364,N_8704,N_8192);
xnor U9365 (N_9365,N_8699,N_8269);
nand U9366 (N_9366,N_8680,N_8470);
and U9367 (N_9367,N_8232,N_8264);
nor U9368 (N_9368,N_8045,N_8713);
nor U9369 (N_9369,N_8012,N_8187);
nand U9370 (N_9370,N_8268,N_8125);
and U9371 (N_9371,N_8006,N_8197);
and U9372 (N_9372,N_8213,N_8542);
nor U9373 (N_9373,N_8226,N_8301);
xor U9374 (N_9374,N_8832,N_8786);
nor U9375 (N_9375,N_8080,N_8626);
or U9376 (N_9376,N_8514,N_8730);
and U9377 (N_9377,N_8766,N_8411);
and U9378 (N_9378,N_8510,N_8013);
nor U9379 (N_9379,N_8619,N_8857);
nand U9380 (N_9380,N_8907,N_8890);
nor U9381 (N_9381,N_8904,N_8808);
or U9382 (N_9382,N_8295,N_8214);
nand U9383 (N_9383,N_8302,N_8333);
or U9384 (N_9384,N_8994,N_8802);
nand U9385 (N_9385,N_8035,N_8309);
nor U9386 (N_9386,N_8173,N_8511);
nand U9387 (N_9387,N_8945,N_8609);
or U9388 (N_9388,N_8177,N_8366);
nand U9389 (N_9389,N_8916,N_8637);
and U9390 (N_9390,N_8841,N_8419);
nand U9391 (N_9391,N_8015,N_8288);
or U9392 (N_9392,N_8603,N_8082);
nand U9393 (N_9393,N_8757,N_8243);
nand U9394 (N_9394,N_8089,N_8104);
or U9395 (N_9395,N_8482,N_8329);
and U9396 (N_9396,N_8578,N_8997);
nor U9397 (N_9397,N_8169,N_8960);
xor U9398 (N_9398,N_8848,N_8488);
nand U9399 (N_9399,N_8778,N_8422);
and U9400 (N_9400,N_8070,N_8972);
nor U9401 (N_9401,N_8782,N_8178);
or U9402 (N_9402,N_8989,N_8332);
and U9403 (N_9403,N_8656,N_8182);
xor U9404 (N_9404,N_8669,N_8131);
and U9405 (N_9405,N_8351,N_8074);
or U9406 (N_9406,N_8420,N_8869);
nand U9407 (N_9407,N_8917,N_8481);
or U9408 (N_9408,N_8379,N_8892);
nand U9409 (N_9409,N_8556,N_8138);
nor U9410 (N_9410,N_8384,N_8767);
xor U9411 (N_9411,N_8049,N_8964);
or U9412 (N_9412,N_8257,N_8478);
and U9413 (N_9413,N_8442,N_8862);
xnor U9414 (N_9414,N_8896,N_8985);
nor U9415 (N_9415,N_8829,N_8454);
nand U9416 (N_9416,N_8382,N_8591);
nand U9417 (N_9417,N_8962,N_8652);
or U9418 (N_9418,N_8882,N_8324);
nor U9419 (N_9419,N_8085,N_8367);
and U9420 (N_9420,N_8140,N_8664);
or U9421 (N_9421,N_8403,N_8564);
xnor U9422 (N_9422,N_8111,N_8739);
nand U9423 (N_9423,N_8476,N_8805);
nand U9424 (N_9424,N_8485,N_8490);
nor U9425 (N_9425,N_8433,N_8079);
or U9426 (N_9426,N_8342,N_8914);
and U9427 (N_9427,N_8654,N_8091);
nor U9428 (N_9428,N_8430,N_8794);
and U9429 (N_9429,N_8590,N_8913);
nand U9430 (N_9430,N_8700,N_8372);
and U9431 (N_9431,N_8421,N_8785);
or U9432 (N_9432,N_8846,N_8168);
or U9433 (N_9433,N_8811,N_8981);
nor U9434 (N_9434,N_8920,N_8750);
or U9435 (N_9435,N_8941,N_8392);
and U9436 (N_9436,N_8752,N_8665);
nand U9437 (N_9437,N_8437,N_8189);
nand U9438 (N_9438,N_8821,N_8101);
and U9439 (N_9439,N_8905,N_8356);
xnor U9440 (N_9440,N_8495,N_8604);
and U9441 (N_9441,N_8864,N_8277);
nand U9442 (N_9442,N_8152,N_8023);
nor U9443 (N_9443,N_8331,N_8175);
nor U9444 (N_9444,N_8798,N_8508);
and U9445 (N_9445,N_8806,N_8875);
and U9446 (N_9446,N_8549,N_8196);
nor U9447 (N_9447,N_8505,N_8114);
xor U9448 (N_9448,N_8184,N_8058);
nor U9449 (N_9449,N_8303,N_8499);
nand U9450 (N_9450,N_8255,N_8033);
and U9451 (N_9451,N_8793,N_8932);
nor U9452 (N_9452,N_8001,N_8450);
or U9453 (N_9453,N_8863,N_8724);
nor U9454 (N_9454,N_8065,N_8804);
or U9455 (N_9455,N_8311,N_8605);
xor U9456 (N_9456,N_8375,N_8555);
and U9457 (N_9457,N_8093,N_8789);
xor U9458 (N_9458,N_8115,N_8720);
nor U9459 (N_9459,N_8344,N_8120);
xnor U9460 (N_9460,N_8143,N_8194);
and U9461 (N_9461,N_8360,N_8824);
xnor U9462 (N_9462,N_8760,N_8118);
nand U9463 (N_9463,N_8106,N_8574);
nand U9464 (N_9464,N_8645,N_8628);
nand U9465 (N_9465,N_8265,N_8978);
nand U9466 (N_9466,N_8406,N_8635);
nand U9467 (N_9467,N_8951,N_8380);
nor U9468 (N_9468,N_8155,N_8312);
or U9469 (N_9469,N_8241,N_8046);
nor U9470 (N_9470,N_8103,N_8692);
nand U9471 (N_9471,N_8873,N_8884);
and U9472 (N_9472,N_8146,N_8223);
and U9473 (N_9473,N_8338,N_8240);
and U9474 (N_9474,N_8459,N_8930);
and U9475 (N_9475,N_8719,N_8565);
nor U9476 (N_9476,N_8550,N_8209);
or U9477 (N_9477,N_8256,N_8552);
nor U9478 (N_9478,N_8318,N_8098);
or U9479 (N_9479,N_8061,N_8607);
xnor U9480 (N_9480,N_8048,N_8707);
or U9481 (N_9481,N_8623,N_8703);
nor U9482 (N_9482,N_8831,N_8201);
and U9483 (N_9483,N_8220,N_8043);
and U9484 (N_9484,N_8855,N_8341);
xnor U9485 (N_9485,N_8616,N_8335);
and U9486 (N_9486,N_8211,N_8734);
xor U9487 (N_9487,N_8253,N_8252);
or U9488 (N_9488,N_8166,N_8858);
nand U9489 (N_9489,N_8934,N_8271);
nor U9490 (N_9490,N_8797,N_8287);
xor U9491 (N_9491,N_8575,N_8736);
nand U9492 (N_9492,N_8186,N_8179);
nand U9493 (N_9493,N_8787,N_8729);
nor U9494 (N_9494,N_8017,N_8359);
nand U9495 (N_9495,N_8950,N_8942);
nor U9496 (N_9496,N_8839,N_8124);
nand U9497 (N_9497,N_8631,N_8087);
and U9498 (N_9498,N_8323,N_8330);
nor U9499 (N_9499,N_8728,N_8658);
or U9500 (N_9500,N_8159,N_8433);
nor U9501 (N_9501,N_8530,N_8478);
nor U9502 (N_9502,N_8850,N_8787);
nand U9503 (N_9503,N_8571,N_8316);
or U9504 (N_9504,N_8740,N_8449);
nand U9505 (N_9505,N_8030,N_8456);
or U9506 (N_9506,N_8118,N_8180);
nand U9507 (N_9507,N_8587,N_8392);
and U9508 (N_9508,N_8174,N_8491);
nor U9509 (N_9509,N_8931,N_8858);
and U9510 (N_9510,N_8359,N_8230);
and U9511 (N_9511,N_8761,N_8301);
nor U9512 (N_9512,N_8764,N_8566);
and U9513 (N_9513,N_8243,N_8993);
xor U9514 (N_9514,N_8073,N_8431);
nand U9515 (N_9515,N_8744,N_8156);
or U9516 (N_9516,N_8086,N_8664);
and U9517 (N_9517,N_8809,N_8387);
xnor U9518 (N_9518,N_8386,N_8159);
or U9519 (N_9519,N_8813,N_8271);
and U9520 (N_9520,N_8617,N_8302);
and U9521 (N_9521,N_8260,N_8591);
or U9522 (N_9522,N_8484,N_8313);
or U9523 (N_9523,N_8485,N_8925);
or U9524 (N_9524,N_8731,N_8698);
nand U9525 (N_9525,N_8050,N_8156);
nand U9526 (N_9526,N_8158,N_8009);
nor U9527 (N_9527,N_8899,N_8976);
and U9528 (N_9528,N_8329,N_8773);
and U9529 (N_9529,N_8047,N_8158);
and U9530 (N_9530,N_8635,N_8399);
and U9531 (N_9531,N_8341,N_8353);
or U9532 (N_9532,N_8936,N_8703);
and U9533 (N_9533,N_8412,N_8133);
nor U9534 (N_9534,N_8504,N_8306);
nor U9535 (N_9535,N_8370,N_8434);
or U9536 (N_9536,N_8628,N_8243);
or U9537 (N_9537,N_8322,N_8737);
nand U9538 (N_9538,N_8448,N_8791);
and U9539 (N_9539,N_8214,N_8134);
and U9540 (N_9540,N_8491,N_8504);
nand U9541 (N_9541,N_8637,N_8776);
and U9542 (N_9542,N_8940,N_8238);
nand U9543 (N_9543,N_8671,N_8424);
nand U9544 (N_9544,N_8837,N_8936);
and U9545 (N_9545,N_8288,N_8202);
nor U9546 (N_9546,N_8826,N_8788);
and U9547 (N_9547,N_8684,N_8057);
nor U9548 (N_9548,N_8424,N_8277);
nor U9549 (N_9549,N_8093,N_8303);
or U9550 (N_9550,N_8319,N_8968);
nor U9551 (N_9551,N_8452,N_8439);
or U9552 (N_9552,N_8861,N_8621);
or U9553 (N_9553,N_8523,N_8805);
or U9554 (N_9554,N_8546,N_8068);
or U9555 (N_9555,N_8640,N_8080);
nand U9556 (N_9556,N_8077,N_8484);
nand U9557 (N_9557,N_8014,N_8352);
or U9558 (N_9558,N_8116,N_8587);
and U9559 (N_9559,N_8076,N_8679);
and U9560 (N_9560,N_8384,N_8437);
nor U9561 (N_9561,N_8358,N_8497);
nor U9562 (N_9562,N_8900,N_8454);
or U9563 (N_9563,N_8017,N_8656);
and U9564 (N_9564,N_8353,N_8885);
nor U9565 (N_9565,N_8181,N_8862);
and U9566 (N_9566,N_8796,N_8856);
or U9567 (N_9567,N_8134,N_8170);
nor U9568 (N_9568,N_8284,N_8564);
or U9569 (N_9569,N_8461,N_8108);
nand U9570 (N_9570,N_8501,N_8242);
or U9571 (N_9571,N_8761,N_8196);
nand U9572 (N_9572,N_8048,N_8445);
nor U9573 (N_9573,N_8920,N_8566);
nor U9574 (N_9574,N_8015,N_8353);
and U9575 (N_9575,N_8704,N_8738);
nor U9576 (N_9576,N_8016,N_8474);
nand U9577 (N_9577,N_8614,N_8655);
nor U9578 (N_9578,N_8242,N_8605);
or U9579 (N_9579,N_8788,N_8967);
and U9580 (N_9580,N_8095,N_8457);
xor U9581 (N_9581,N_8447,N_8421);
nor U9582 (N_9582,N_8447,N_8038);
nand U9583 (N_9583,N_8851,N_8971);
and U9584 (N_9584,N_8079,N_8454);
or U9585 (N_9585,N_8936,N_8119);
or U9586 (N_9586,N_8124,N_8596);
xnor U9587 (N_9587,N_8590,N_8807);
nand U9588 (N_9588,N_8588,N_8124);
nor U9589 (N_9589,N_8811,N_8236);
nor U9590 (N_9590,N_8731,N_8657);
nand U9591 (N_9591,N_8005,N_8083);
and U9592 (N_9592,N_8081,N_8594);
or U9593 (N_9593,N_8439,N_8210);
and U9594 (N_9594,N_8045,N_8274);
or U9595 (N_9595,N_8739,N_8492);
nor U9596 (N_9596,N_8033,N_8664);
nand U9597 (N_9597,N_8216,N_8879);
or U9598 (N_9598,N_8524,N_8859);
nand U9599 (N_9599,N_8793,N_8517);
or U9600 (N_9600,N_8683,N_8610);
and U9601 (N_9601,N_8663,N_8165);
nand U9602 (N_9602,N_8609,N_8630);
nor U9603 (N_9603,N_8121,N_8485);
or U9604 (N_9604,N_8272,N_8916);
and U9605 (N_9605,N_8263,N_8485);
xor U9606 (N_9606,N_8654,N_8105);
or U9607 (N_9607,N_8658,N_8072);
nor U9608 (N_9608,N_8466,N_8992);
or U9609 (N_9609,N_8531,N_8515);
nand U9610 (N_9610,N_8603,N_8051);
and U9611 (N_9611,N_8638,N_8751);
xor U9612 (N_9612,N_8261,N_8876);
nor U9613 (N_9613,N_8989,N_8286);
nor U9614 (N_9614,N_8570,N_8688);
nor U9615 (N_9615,N_8436,N_8195);
or U9616 (N_9616,N_8826,N_8755);
nand U9617 (N_9617,N_8709,N_8517);
xnor U9618 (N_9618,N_8344,N_8138);
nor U9619 (N_9619,N_8345,N_8570);
and U9620 (N_9620,N_8070,N_8708);
and U9621 (N_9621,N_8477,N_8061);
nor U9622 (N_9622,N_8930,N_8623);
and U9623 (N_9623,N_8798,N_8453);
or U9624 (N_9624,N_8079,N_8644);
and U9625 (N_9625,N_8218,N_8167);
nand U9626 (N_9626,N_8275,N_8607);
and U9627 (N_9627,N_8638,N_8167);
and U9628 (N_9628,N_8572,N_8220);
xor U9629 (N_9629,N_8822,N_8521);
or U9630 (N_9630,N_8802,N_8202);
or U9631 (N_9631,N_8019,N_8518);
nor U9632 (N_9632,N_8986,N_8261);
nor U9633 (N_9633,N_8281,N_8435);
and U9634 (N_9634,N_8151,N_8292);
nor U9635 (N_9635,N_8708,N_8693);
or U9636 (N_9636,N_8133,N_8427);
nand U9637 (N_9637,N_8572,N_8651);
and U9638 (N_9638,N_8937,N_8203);
or U9639 (N_9639,N_8686,N_8020);
nand U9640 (N_9640,N_8843,N_8461);
and U9641 (N_9641,N_8651,N_8038);
or U9642 (N_9642,N_8629,N_8811);
xnor U9643 (N_9643,N_8737,N_8969);
nand U9644 (N_9644,N_8308,N_8530);
or U9645 (N_9645,N_8276,N_8545);
or U9646 (N_9646,N_8983,N_8702);
nand U9647 (N_9647,N_8190,N_8844);
and U9648 (N_9648,N_8558,N_8491);
nor U9649 (N_9649,N_8675,N_8097);
xnor U9650 (N_9650,N_8254,N_8376);
nand U9651 (N_9651,N_8031,N_8743);
nor U9652 (N_9652,N_8940,N_8809);
and U9653 (N_9653,N_8806,N_8165);
xnor U9654 (N_9654,N_8489,N_8152);
or U9655 (N_9655,N_8317,N_8928);
and U9656 (N_9656,N_8023,N_8622);
and U9657 (N_9657,N_8388,N_8914);
nand U9658 (N_9658,N_8854,N_8834);
and U9659 (N_9659,N_8912,N_8135);
and U9660 (N_9660,N_8723,N_8323);
or U9661 (N_9661,N_8799,N_8075);
or U9662 (N_9662,N_8588,N_8637);
nor U9663 (N_9663,N_8382,N_8776);
and U9664 (N_9664,N_8534,N_8220);
nand U9665 (N_9665,N_8804,N_8616);
and U9666 (N_9666,N_8994,N_8827);
and U9667 (N_9667,N_8384,N_8873);
nor U9668 (N_9668,N_8008,N_8616);
or U9669 (N_9669,N_8676,N_8518);
nand U9670 (N_9670,N_8084,N_8738);
or U9671 (N_9671,N_8079,N_8389);
nor U9672 (N_9672,N_8984,N_8497);
or U9673 (N_9673,N_8509,N_8395);
nand U9674 (N_9674,N_8192,N_8631);
or U9675 (N_9675,N_8424,N_8399);
nand U9676 (N_9676,N_8978,N_8642);
xor U9677 (N_9677,N_8909,N_8678);
or U9678 (N_9678,N_8708,N_8373);
nand U9679 (N_9679,N_8566,N_8719);
nand U9680 (N_9680,N_8819,N_8303);
or U9681 (N_9681,N_8265,N_8846);
nand U9682 (N_9682,N_8657,N_8184);
nor U9683 (N_9683,N_8429,N_8191);
nand U9684 (N_9684,N_8082,N_8925);
xnor U9685 (N_9685,N_8249,N_8795);
and U9686 (N_9686,N_8701,N_8568);
or U9687 (N_9687,N_8406,N_8908);
nand U9688 (N_9688,N_8729,N_8420);
nand U9689 (N_9689,N_8452,N_8069);
or U9690 (N_9690,N_8961,N_8920);
or U9691 (N_9691,N_8235,N_8618);
nor U9692 (N_9692,N_8195,N_8120);
xnor U9693 (N_9693,N_8675,N_8878);
and U9694 (N_9694,N_8338,N_8975);
and U9695 (N_9695,N_8764,N_8186);
nor U9696 (N_9696,N_8896,N_8965);
or U9697 (N_9697,N_8030,N_8061);
or U9698 (N_9698,N_8936,N_8437);
nor U9699 (N_9699,N_8800,N_8806);
and U9700 (N_9700,N_8575,N_8498);
nand U9701 (N_9701,N_8101,N_8071);
or U9702 (N_9702,N_8690,N_8550);
and U9703 (N_9703,N_8530,N_8586);
or U9704 (N_9704,N_8052,N_8799);
or U9705 (N_9705,N_8970,N_8448);
xor U9706 (N_9706,N_8883,N_8235);
and U9707 (N_9707,N_8654,N_8502);
nor U9708 (N_9708,N_8735,N_8787);
or U9709 (N_9709,N_8423,N_8930);
nand U9710 (N_9710,N_8932,N_8652);
or U9711 (N_9711,N_8652,N_8692);
nor U9712 (N_9712,N_8799,N_8045);
xnor U9713 (N_9713,N_8121,N_8027);
and U9714 (N_9714,N_8417,N_8977);
nand U9715 (N_9715,N_8562,N_8436);
xor U9716 (N_9716,N_8035,N_8385);
and U9717 (N_9717,N_8991,N_8077);
xor U9718 (N_9718,N_8726,N_8826);
nor U9719 (N_9719,N_8460,N_8237);
nand U9720 (N_9720,N_8698,N_8646);
nor U9721 (N_9721,N_8511,N_8836);
nor U9722 (N_9722,N_8408,N_8855);
xor U9723 (N_9723,N_8377,N_8626);
and U9724 (N_9724,N_8130,N_8238);
and U9725 (N_9725,N_8204,N_8769);
and U9726 (N_9726,N_8774,N_8023);
or U9727 (N_9727,N_8969,N_8090);
nand U9728 (N_9728,N_8652,N_8981);
xor U9729 (N_9729,N_8313,N_8585);
and U9730 (N_9730,N_8060,N_8103);
and U9731 (N_9731,N_8188,N_8060);
or U9732 (N_9732,N_8938,N_8023);
xor U9733 (N_9733,N_8560,N_8553);
nand U9734 (N_9734,N_8379,N_8624);
and U9735 (N_9735,N_8177,N_8388);
and U9736 (N_9736,N_8019,N_8293);
xor U9737 (N_9737,N_8877,N_8865);
nor U9738 (N_9738,N_8198,N_8193);
or U9739 (N_9739,N_8428,N_8693);
and U9740 (N_9740,N_8090,N_8156);
and U9741 (N_9741,N_8678,N_8146);
or U9742 (N_9742,N_8915,N_8664);
nand U9743 (N_9743,N_8462,N_8631);
nor U9744 (N_9744,N_8666,N_8971);
nor U9745 (N_9745,N_8325,N_8896);
nand U9746 (N_9746,N_8991,N_8612);
nand U9747 (N_9747,N_8727,N_8896);
nor U9748 (N_9748,N_8221,N_8852);
and U9749 (N_9749,N_8009,N_8871);
nor U9750 (N_9750,N_8557,N_8670);
nand U9751 (N_9751,N_8404,N_8807);
nand U9752 (N_9752,N_8306,N_8773);
nand U9753 (N_9753,N_8124,N_8994);
xor U9754 (N_9754,N_8142,N_8204);
nor U9755 (N_9755,N_8132,N_8555);
nor U9756 (N_9756,N_8897,N_8957);
nor U9757 (N_9757,N_8322,N_8685);
nor U9758 (N_9758,N_8915,N_8197);
or U9759 (N_9759,N_8082,N_8493);
nor U9760 (N_9760,N_8179,N_8577);
nand U9761 (N_9761,N_8095,N_8552);
nor U9762 (N_9762,N_8320,N_8827);
nor U9763 (N_9763,N_8825,N_8146);
xor U9764 (N_9764,N_8886,N_8954);
or U9765 (N_9765,N_8715,N_8309);
nand U9766 (N_9766,N_8941,N_8909);
or U9767 (N_9767,N_8724,N_8780);
nand U9768 (N_9768,N_8098,N_8677);
and U9769 (N_9769,N_8397,N_8047);
nand U9770 (N_9770,N_8337,N_8969);
nor U9771 (N_9771,N_8161,N_8621);
xnor U9772 (N_9772,N_8818,N_8085);
or U9773 (N_9773,N_8668,N_8214);
nand U9774 (N_9774,N_8898,N_8611);
and U9775 (N_9775,N_8316,N_8315);
nand U9776 (N_9776,N_8286,N_8493);
nand U9777 (N_9777,N_8373,N_8821);
nand U9778 (N_9778,N_8339,N_8807);
nand U9779 (N_9779,N_8922,N_8058);
or U9780 (N_9780,N_8426,N_8528);
nor U9781 (N_9781,N_8762,N_8792);
and U9782 (N_9782,N_8766,N_8043);
xor U9783 (N_9783,N_8931,N_8837);
nand U9784 (N_9784,N_8250,N_8432);
nand U9785 (N_9785,N_8388,N_8083);
and U9786 (N_9786,N_8648,N_8577);
or U9787 (N_9787,N_8360,N_8715);
nand U9788 (N_9788,N_8128,N_8177);
and U9789 (N_9789,N_8176,N_8094);
nor U9790 (N_9790,N_8982,N_8163);
xor U9791 (N_9791,N_8572,N_8563);
or U9792 (N_9792,N_8760,N_8267);
and U9793 (N_9793,N_8693,N_8231);
and U9794 (N_9794,N_8816,N_8801);
nor U9795 (N_9795,N_8230,N_8109);
nor U9796 (N_9796,N_8828,N_8846);
nand U9797 (N_9797,N_8316,N_8092);
or U9798 (N_9798,N_8767,N_8110);
or U9799 (N_9799,N_8857,N_8470);
or U9800 (N_9800,N_8950,N_8907);
nand U9801 (N_9801,N_8732,N_8720);
nor U9802 (N_9802,N_8729,N_8580);
nand U9803 (N_9803,N_8453,N_8263);
and U9804 (N_9804,N_8229,N_8825);
or U9805 (N_9805,N_8715,N_8742);
or U9806 (N_9806,N_8679,N_8533);
nand U9807 (N_9807,N_8910,N_8653);
and U9808 (N_9808,N_8757,N_8683);
and U9809 (N_9809,N_8925,N_8159);
or U9810 (N_9810,N_8111,N_8495);
or U9811 (N_9811,N_8549,N_8521);
or U9812 (N_9812,N_8387,N_8562);
and U9813 (N_9813,N_8000,N_8994);
nor U9814 (N_9814,N_8071,N_8504);
nand U9815 (N_9815,N_8346,N_8260);
or U9816 (N_9816,N_8916,N_8315);
xor U9817 (N_9817,N_8876,N_8062);
and U9818 (N_9818,N_8481,N_8914);
nand U9819 (N_9819,N_8325,N_8405);
or U9820 (N_9820,N_8025,N_8523);
nand U9821 (N_9821,N_8126,N_8654);
or U9822 (N_9822,N_8383,N_8301);
xnor U9823 (N_9823,N_8639,N_8354);
and U9824 (N_9824,N_8567,N_8924);
or U9825 (N_9825,N_8844,N_8121);
nand U9826 (N_9826,N_8476,N_8007);
xnor U9827 (N_9827,N_8099,N_8651);
nand U9828 (N_9828,N_8276,N_8491);
xor U9829 (N_9829,N_8950,N_8793);
or U9830 (N_9830,N_8668,N_8782);
nand U9831 (N_9831,N_8617,N_8717);
nor U9832 (N_9832,N_8250,N_8224);
nand U9833 (N_9833,N_8907,N_8857);
nor U9834 (N_9834,N_8878,N_8107);
nor U9835 (N_9835,N_8063,N_8458);
and U9836 (N_9836,N_8192,N_8196);
and U9837 (N_9837,N_8203,N_8901);
and U9838 (N_9838,N_8760,N_8344);
and U9839 (N_9839,N_8864,N_8037);
and U9840 (N_9840,N_8292,N_8995);
or U9841 (N_9841,N_8051,N_8699);
and U9842 (N_9842,N_8677,N_8790);
xor U9843 (N_9843,N_8545,N_8087);
and U9844 (N_9844,N_8856,N_8052);
xor U9845 (N_9845,N_8898,N_8806);
nor U9846 (N_9846,N_8231,N_8737);
or U9847 (N_9847,N_8981,N_8821);
and U9848 (N_9848,N_8564,N_8207);
or U9849 (N_9849,N_8742,N_8284);
nor U9850 (N_9850,N_8659,N_8715);
nand U9851 (N_9851,N_8996,N_8993);
and U9852 (N_9852,N_8542,N_8174);
nand U9853 (N_9853,N_8827,N_8166);
nand U9854 (N_9854,N_8372,N_8748);
nand U9855 (N_9855,N_8339,N_8789);
and U9856 (N_9856,N_8199,N_8691);
and U9857 (N_9857,N_8341,N_8817);
nand U9858 (N_9858,N_8023,N_8002);
or U9859 (N_9859,N_8883,N_8706);
and U9860 (N_9860,N_8562,N_8511);
nor U9861 (N_9861,N_8012,N_8164);
nor U9862 (N_9862,N_8332,N_8329);
and U9863 (N_9863,N_8256,N_8866);
xnor U9864 (N_9864,N_8065,N_8474);
nand U9865 (N_9865,N_8186,N_8606);
xor U9866 (N_9866,N_8034,N_8879);
nor U9867 (N_9867,N_8426,N_8736);
xnor U9868 (N_9868,N_8457,N_8907);
xor U9869 (N_9869,N_8838,N_8611);
nand U9870 (N_9870,N_8057,N_8992);
or U9871 (N_9871,N_8421,N_8143);
or U9872 (N_9872,N_8911,N_8135);
or U9873 (N_9873,N_8625,N_8924);
or U9874 (N_9874,N_8425,N_8214);
nand U9875 (N_9875,N_8853,N_8504);
nor U9876 (N_9876,N_8970,N_8164);
or U9877 (N_9877,N_8153,N_8692);
or U9878 (N_9878,N_8969,N_8999);
or U9879 (N_9879,N_8597,N_8106);
nor U9880 (N_9880,N_8895,N_8843);
xor U9881 (N_9881,N_8372,N_8648);
nor U9882 (N_9882,N_8073,N_8120);
and U9883 (N_9883,N_8264,N_8434);
and U9884 (N_9884,N_8428,N_8023);
xor U9885 (N_9885,N_8209,N_8780);
nor U9886 (N_9886,N_8759,N_8134);
and U9887 (N_9887,N_8630,N_8126);
xnor U9888 (N_9888,N_8890,N_8851);
nor U9889 (N_9889,N_8488,N_8526);
or U9890 (N_9890,N_8815,N_8855);
or U9891 (N_9891,N_8502,N_8645);
and U9892 (N_9892,N_8037,N_8190);
xor U9893 (N_9893,N_8334,N_8738);
nor U9894 (N_9894,N_8600,N_8916);
nor U9895 (N_9895,N_8968,N_8226);
and U9896 (N_9896,N_8599,N_8347);
xnor U9897 (N_9897,N_8903,N_8082);
nand U9898 (N_9898,N_8735,N_8324);
or U9899 (N_9899,N_8441,N_8762);
or U9900 (N_9900,N_8809,N_8081);
xnor U9901 (N_9901,N_8768,N_8955);
nor U9902 (N_9902,N_8812,N_8445);
nand U9903 (N_9903,N_8880,N_8343);
nor U9904 (N_9904,N_8457,N_8939);
xor U9905 (N_9905,N_8715,N_8665);
or U9906 (N_9906,N_8030,N_8727);
xnor U9907 (N_9907,N_8058,N_8376);
nor U9908 (N_9908,N_8991,N_8590);
nor U9909 (N_9909,N_8381,N_8595);
nor U9910 (N_9910,N_8174,N_8180);
nor U9911 (N_9911,N_8257,N_8009);
nand U9912 (N_9912,N_8879,N_8412);
and U9913 (N_9913,N_8432,N_8209);
xor U9914 (N_9914,N_8361,N_8750);
xnor U9915 (N_9915,N_8932,N_8632);
or U9916 (N_9916,N_8634,N_8931);
nand U9917 (N_9917,N_8496,N_8645);
and U9918 (N_9918,N_8356,N_8390);
xor U9919 (N_9919,N_8019,N_8580);
xnor U9920 (N_9920,N_8521,N_8814);
nand U9921 (N_9921,N_8956,N_8497);
or U9922 (N_9922,N_8092,N_8691);
and U9923 (N_9923,N_8471,N_8588);
xor U9924 (N_9924,N_8357,N_8723);
xor U9925 (N_9925,N_8676,N_8868);
and U9926 (N_9926,N_8873,N_8953);
or U9927 (N_9927,N_8382,N_8559);
nand U9928 (N_9928,N_8789,N_8979);
xor U9929 (N_9929,N_8787,N_8717);
nor U9930 (N_9930,N_8294,N_8598);
nor U9931 (N_9931,N_8754,N_8857);
or U9932 (N_9932,N_8854,N_8428);
or U9933 (N_9933,N_8419,N_8629);
nor U9934 (N_9934,N_8887,N_8278);
nor U9935 (N_9935,N_8448,N_8871);
nor U9936 (N_9936,N_8865,N_8697);
or U9937 (N_9937,N_8220,N_8689);
xor U9938 (N_9938,N_8264,N_8095);
and U9939 (N_9939,N_8086,N_8357);
nand U9940 (N_9940,N_8422,N_8309);
nand U9941 (N_9941,N_8268,N_8409);
nand U9942 (N_9942,N_8765,N_8615);
nor U9943 (N_9943,N_8590,N_8870);
nor U9944 (N_9944,N_8027,N_8389);
or U9945 (N_9945,N_8317,N_8613);
and U9946 (N_9946,N_8219,N_8380);
or U9947 (N_9947,N_8849,N_8154);
nor U9948 (N_9948,N_8839,N_8184);
xor U9949 (N_9949,N_8812,N_8593);
nand U9950 (N_9950,N_8823,N_8835);
nor U9951 (N_9951,N_8419,N_8680);
and U9952 (N_9952,N_8633,N_8840);
nand U9953 (N_9953,N_8196,N_8259);
nor U9954 (N_9954,N_8136,N_8226);
nand U9955 (N_9955,N_8345,N_8792);
nand U9956 (N_9956,N_8456,N_8659);
or U9957 (N_9957,N_8105,N_8271);
or U9958 (N_9958,N_8840,N_8062);
or U9959 (N_9959,N_8900,N_8119);
or U9960 (N_9960,N_8922,N_8174);
nor U9961 (N_9961,N_8218,N_8888);
nor U9962 (N_9962,N_8752,N_8740);
nor U9963 (N_9963,N_8780,N_8575);
or U9964 (N_9964,N_8862,N_8587);
nor U9965 (N_9965,N_8868,N_8703);
nor U9966 (N_9966,N_8018,N_8198);
nor U9967 (N_9967,N_8225,N_8725);
nor U9968 (N_9968,N_8895,N_8606);
xnor U9969 (N_9969,N_8088,N_8003);
nor U9970 (N_9970,N_8378,N_8327);
and U9971 (N_9971,N_8475,N_8669);
and U9972 (N_9972,N_8128,N_8891);
nand U9973 (N_9973,N_8372,N_8671);
and U9974 (N_9974,N_8643,N_8552);
nor U9975 (N_9975,N_8603,N_8468);
nor U9976 (N_9976,N_8242,N_8374);
and U9977 (N_9977,N_8963,N_8934);
nand U9978 (N_9978,N_8739,N_8225);
and U9979 (N_9979,N_8006,N_8789);
nand U9980 (N_9980,N_8672,N_8185);
and U9981 (N_9981,N_8819,N_8931);
nor U9982 (N_9982,N_8855,N_8197);
nand U9983 (N_9983,N_8342,N_8383);
nand U9984 (N_9984,N_8399,N_8230);
and U9985 (N_9985,N_8261,N_8507);
and U9986 (N_9986,N_8278,N_8316);
or U9987 (N_9987,N_8397,N_8237);
nor U9988 (N_9988,N_8901,N_8401);
or U9989 (N_9989,N_8058,N_8850);
and U9990 (N_9990,N_8508,N_8725);
nor U9991 (N_9991,N_8519,N_8121);
xnor U9992 (N_9992,N_8386,N_8325);
nor U9993 (N_9993,N_8212,N_8494);
and U9994 (N_9994,N_8043,N_8192);
and U9995 (N_9995,N_8036,N_8414);
nand U9996 (N_9996,N_8643,N_8754);
nor U9997 (N_9997,N_8216,N_8472);
or U9998 (N_9998,N_8331,N_8596);
nand U9999 (N_9999,N_8838,N_8199);
nor UO_0 (O_0,N_9825,N_9438);
nand UO_1 (O_1,N_9840,N_9395);
nand UO_2 (O_2,N_9106,N_9744);
nand UO_3 (O_3,N_9482,N_9291);
nor UO_4 (O_4,N_9435,N_9972);
or UO_5 (O_5,N_9186,N_9533);
nor UO_6 (O_6,N_9779,N_9928);
or UO_7 (O_7,N_9300,N_9866);
nand UO_8 (O_8,N_9181,N_9777);
xor UO_9 (O_9,N_9970,N_9556);
or UO_10 (O_10,N_9770,N_9303);
xnor UO_11 (O_11,N_9297,N_9999);
nand UO_12 (O_12,N_9974,N_9256);
xor UO_13 (O_13,N_9439,N_9322);
nand UO_14 (O_14,N_9233,N_9028);
xnor UO_15 (O_15,N_9656,N_9286);
or UO_16 (O_16,N_9477,N_9512);
or UO_17 (O_17,N_9728,N_9400);
and UO_18 (O_18,N_9516,N_9369);
nand UO_19 (O_19,N_9195,N_9150);
nor UO_20 (O_20,N_9610,N_9007);
nor UO_21 (O_21,N_9714,N_9382);
nand UO_22 (O_22,N_9469,N_9496);
nand UO_23 (O_23,N_9151,N_9807);
and UO_24 (O_24,N_9733,N_9391);
or UO_25 (O_25,N_9888,N_9585);
or UO_26 (O_26,N_9555,N_9843);
and UO_27 (O_27,N_9984,N_9913);
nand UO_28 (O_28,N_9763,N_9097);
and UO_29 (O_29,N_9667,N_9146);
or UO_30 (O_30,N_9328,N_9713);
and UO_31 (O_31,N_9758,N_9942);
nor UO_32 (O_32,N_9488,N_9899);
nand UO_33 (O_33,N_9910,N_9637);
and UO_34 (O_34,N_9990,N_9611);
xor UO_35 (O_35,N_9451,N_9618);
nor UO_36 (O_36,N_9077,N_9874);
or UO_37 (O_37,N_9992,N_9677);
and UO_38 (O_38,N_9155,N_9827);
nand UO_39 (O_39,N_9732,N_9617);
xor UO_40 (O_40,N_9952,N_9364);
nor UO_41 (O_41,N_9137,N_9887);
nand UO_42 (O_42,N_9634,N_9564);
or UO_43 (O_43,N_9312,N_9117);
nand UO_44 (O_44,N_9706,N_9852);
nor UO_45 (O_45,N_9093,N_9276);
and UO_46 (O_46,N_9778,N_9110);
or UO_47 (O_47,N_9380,N_9842);
nor UO_48 (O_48,N_9072,N_9554);
and UO_49 (O_49,N_9659,N_9804);
xnor UO_50 (O_50,N_9370,N_9232);
nand UO_51 (O_51,N_9480,N_9129);
or UO_52 (O_52,N_9615,N_9107);
nand UO_53 (O_53,N_9069,N_9803);
or UO_54 (O_54,N_9115,N_9021);
nor UO_55 (O_55,N_9812,N_9414);
or UO_56 (O_56,N_9649,N_9524);
or UO_57 (O_57,N_9546,N_9586);
or UO_58 (O_58,N_9343,N_9755);
and UO_59 (O_59,N_9540,N_9294);
or UO_60 (O_60,N_9773,N_9444);
or UO_61 (O_61,N_9063,N_9962);
xor UO_62 (O_62,N_9141,N_9495);
and UO_63 (O_63,N_9219,N_9349);
nand UO_64 (O_64,N_9004,N_9589);
nor UO_65 (O_65,N_9044,N_9998);
xor UO_66 (O_66,N_9494,N_9473);
nand UO_67 (O_67,N_9961,N_9111);
nor UO_68 (O_68,N_9227,N_9719);
nand UO_69 (O_69,N_9994,N_9797);
nand UO_70 (O_70,N_9440,N_9737);
or UO_71 (O_71,N_9434,N_9768);
and UO_72 (O_72,N_9317,N_9164);
and UO_73 (O_73,N_9404,N_9491);
or UO_74 (O_74,N_9387,N_9614);
nor UO_75 (O_75,N_9454,N_9739);
and UO_76 (O_76,N_9230,N_9749);
nand UO_77 (O_77,N_9809,N_9158);
nor UO_78 (O_78,N_9314,N_9581);
nand UO_79 (O_79,N_9679,N_9075);
or UO_80 (O_80,N_9192,N_9392);
nor UO_81 (O_81,N_9800,N_9460);
nor UO_82 (O_82,N_9967,N_9693);
or UO_83 (O_83,N_9764,N_9787);
nand UO_84 (O_84,N_9453,N_9025);
xnor UO_85 (O_85,N_9327,N_9968);
nand UO_86 (O_86,N_9424,N_9616);
or UO_87 (O_87,N_9786,N_9258);
nand UO_88 (O_88,N_9736,N_9022);
nand UO_89 (O_89,N_9302,N_9034);
xnor UO_90 (O_90,N_9223,N_9049);
or UO_91 (O_91,N_9929,N_9675);
or UO_92 (O_92,N_9879,N_9838);
nor UO_93 (O_93,N_9318,N_9660);
nand UO_94 (O_94,N_9165,N_9521);
xor UO_95 (O_95,N_9224,N_9776);
nand UO_96 (O_96,N_9828,N_9249);
nor UO_97 (O_97,N_9864,N_9356);
and UO_98 (O_98,N_9092,N_9731);
xor UO_99 (O_99,N_9470,N_9848);
and UO_100 (O_100,N_9363,N_9507);
xor UO_101 (O_101,N_9368,N_9694);
nand UO_102 (O_102,N_9397,N_9096);
or UO_103 (O_103,N_9619,N_9854);
nand UO_104 (O_104,N_9071,N_9089);
and UO_105 (O_105,N_9431,N_9310);
nor UO_106 (O_106,N_9598,N_9877);
and UO_107 (O_107,N_9121,N_9673);
nor UO_108 (O_108,N_9166,N_9362);
nand UO_109 (O_109,N_9134,N_9518);
xor UO_110 (O_110,N_9243,N_9196);
nor UO_111 (O_111,N_9251,N_9650);
nor UO_112 (O_112,N_9215,N_9187);
nor UO_113 (O_113,N_9350,N_9133);
nor UO_114 (O_114,N_9130,N_9508);
and UO_115 (O_115,N_9837,N_9411);
or UO_116 (O_116,N_9427,N_9690);
xnor UO_117 (O_117,N_9290,N_9892);
nor UO_118 (O_118,N_9449,N_9452);
or UO_119 (O_119,N_9640,N_9287);
or UO_120 (O_120,N_9037,N_9475);
nor UO_121 (O_121,N_9216,N_9261);
or UO_122 (O_122,N_9558,N_9509);
or UO_123 (O_123,N_9798,N_9979);
nand UO_124 (O_124,N_9419,N_9398);
and UO_125 (O_125,N_9883,N_9279);
and UO_126 (O_126,N_9943,N_9484);
and UO_127 (O_127,N_9934,N_9868);
nor UO_128 (O_128,N_9461,N_9780);
and UO_129 (O_129,N_9231,N_9337);
and UO_130 (O_130,N_9070,N_9964);
or UO_131 (O_131,N_9059,N_9666);
xor UO_132 (O_132,N_9720,N_9283);
or UO_133 (O_133,N_9281,N_9594);
nor UO_134 (O_134,N_9055,N_9793);
xnor UO_135 (O_135,N_9207,N_9824);
nand UO_136 (O_136,N_9857,N_9735);
and UO_137 (O_137,N_9523,N_9561);
xnor UO_138 (O_138,N_9923,N_9293);
and UO_139 (O_139,N_9008,N_9336);
or UO_140 (O_140,N_9271,N_9474);
nor UO_141 (O_141,N_9050,N_9466);
and UO_142 (O_142,N_9018,N_9331);
nand UO_143 (O_143,N_9194,N_9926);
nor UO_144 (O_144,N_9909,N_9250);
or UO_145 (O_145,N_9774,N_9959);
or UO_146 (O_146,N_9851,N_9607);
or UO_147 (O_147,N_9725,N_9278);
and UO_148 (O_148,N_9685,N_9260);
nand UO_149 (O_149,N_9818,N_9376);
nor UO_150 (O_150,N_9576,N_9174);
and UO_151 (O_151,N_9753,N_9307);
nor UO_152 (O_152,N_9632,N_9032);
or UO_153 (O_153,N_9612,N_9428);
and UO_154 (O_154,N_9856,N_9064);
nor UO_155 (O_155,N_9654,N_9661);
nand UO_156 (O_156,N_9423,N_9889);
and UO_157 (O_157,N_9026,N_9145);
and UO_158 (O_158,N_9846,N_9361);
nand UO_159 (O_159,N_9479,N_9273);
nand UO_160 (O_160,N_9575,N_9394);
and UO_161 (O_161,N_9039,N_9354);
nor UO_162 (O_162,N_9078,N_9308);
or UO_163 (O_163,N_9099,N_9299);
nor UO_164 (O_164,N_9052,N_9939);
and UO_165 (O_165,N_9360,N_9978);
or UO_166 (O_166,N_9221,N_9834);
xnor UO_167 (O_167,N_9220,N_9405);
nand UO_168 (O_168,N_9020,N_9662);
or UO_169 (O_169,N_9432,N_9647);
and UO_170 (O_170,N_9919,N_9547);
nor UO_171 (O_171,N_9638,N_9526);
or UO_172 (O_172,N_9655,N_9298);
or UO_173 (O_173,N_9264,N_9762);
nor UO_174 (O_174,N_9599,N_9886);
and UO_175 (O_175,N_9855,N_9272);
and UO_176 (O_176,N_9241,N_9152);
or UO_177 (O_177,N_9003,N_9206);
and UO_178 (O_178,N_9065,N_9329);
nand UO_179 (O_179,N_9501,N_9965);
or UO_180 (O_180,N_9949,N_9748);
and UO_181 (O_181,N_9458,N_9105);
nand UO_182 (O_182,N_9709,N_9016);
nor UO_183 (O_183,N_9161,N_9184);
nor UO_184 (O_184,N_9193,N_9365);
xnor UO_185 (O_185,N_9352,N_9613);
nand UO_186 (O_186,N_9930,N_9759);
or UO_187 (O_187,N_9073,N_9023);
nand UO_188 (O_188,N_9315,N_9882);
or UO_189 (O_189,N_9875,N_9399);
nor UO_190 (O_190,N_9173,N_9410);
nor UO_191 (O_191,N_9426,N_9788);
and UO_192 (O_192,N_9031,N_9863);
or UO_193 (O_193,N_9334,N_9171);
nand UO_194 (O_194,N_9548,N_9204);
nand UO_195 (O_195,N_9682,N_9982);
nand UO_196 (O_196,N_9963,N_9157);
and UO_197 (O_197,N_9269,N_9375);
and UO_198 (O_198,N_9333,N_9727);
and UO_199 (O_199,N_9353,N_9374);
and UO_200 (O_200,N_9019,N_9305);
or UO_201 (O_201,N_9179,N_9715);
nand UO_202 (O_202,N_9823,N_9583);
nand UO_203 (O_203,N_9498,N_9188);
and UO_204 (O_204,N_9056,N_9805);
nand UO_205 (O_205,N_9723,N_9741);
nor UO_206 (O_206,N_9902,N_9606);
xnor UO_207 (O_207,N_9492,N_9525);
and UO_208 (O_208,N_9528,N_9344);
nor UO_209 (O_209,N_9531,N_9274);
nand UO_210 (O_210,N_9483,N_9320);
or UO_211 (O_211,N_9865,N_9148);
and UO_212 (O_212,N_9562,N_9620);
nor UO_213 (O_213,N_9593,N_9701);
and UO_214 (O_214,N_9955,N_9489);
or UO_215 (O_215,N_9808,N_9149);
or UO_216 (O_216,N_9257,N_9631);
nand UO_217 (O_217,N_9960,N_9202);
nand UO_218 (O_218,N_9420,N_9436);
or UO_219 (O_219,N_9784,N_9678);
or UO_220 (O_220,N_9912,N_9047);
nand UO_221 (O_221,N_9014,N_9917);
nand UO_222 (O_222,N_9935,N_9476);
nand UO_223 (O_223,N_9750,N_9568);
nor UO_224 (O_224,N_9009,N_9806);
or UO_225 (O_225,N_9580,N_9502);
or UO_226 (O_226,N_9871,N_9658);
or UO_227 (O_227,N_9467,N_9132);
and UO_228 (O_228,N_9408,N_9513);
nand UO_229 (O_229,N_9313,N_9275);
nor UO_230 (O_230,N_9574,N_9625);
nand UO_231 (O_231,N_9170,N_9058);
or UO_232 (O_232,N_9756,N_9462);
or UO_233 (O_233,N_9550,N_9190);
or UO_234 (O_234,N_9729,N_9730);
or UO_235 (O_235,N_9602,N_9153);
or UO_236 (O_236,N_9332,N_9384);
nand UO_237 (O_237,N_9218,N_9745);
or UO_238 (O_238,N_9835,N_9120);
nand UO_239 (O_239,N_9648,N_9029);
xor UO_240 (O_240,N_9708,N_9103);
nor UO_241 (O_241,N_9543,N_9005);
and UO_242 (O_242,N_9908,N_9506);
and UO_243 (O_243,N_9213,N_9168);
or UO_244 (O_244,N_9989,N_9163);
nand UO_245 (O_245,N_9139,N_9988);
xnor UO_246 (O_246,N_9185,N_9895);
and UO_247 (O_247,N_9535,N_9747);
nand UO_248 (O_248,N_9873,N_9811);
and UO_249 (O_249,N_9916,N_9493);
or UO_250 (O_250,N_9742,N_9140);
nand UO_251 (O_251,N_9043,N_9381);
nand UO_252 (O_252,N_9683,N_9932);
nor UO_253 (O_253,N_9890,N_9478);
nand UO_254 (O_254,N_9945,N_9629);
nor UO_255 (O_255,N_9347,N_9503);
xnor UO_256 (O_256,N_9570,N_9002);
nand UO_257 (O_257,N_9053,N_9761);
nand UO_258 (O_258,N_9627,N_9674);
and UO_259 (O_259,N_9027,N_9514);
xnor UO_260 (O_260,N_9635,N_9704);
and UO_261 (O_261,N_9721,N_9520);
or UO_262 (O_262,N_9696,N_9255);
nor UO_263 (O_263,N_9515,N_9421);
or UO_264 (O_264,N_9288,N_9101);
xor UO_265 (O_265,N_9699,N_9335);
nand UO_266 (O_266,N_9552,N_9931);
nor UO_267 (O_267,N_9358,N_9127);
nor UO_268 (O_268,N_9124,N_9373);
and UO_269 (O_269,N_9641,N_9829);
nand UO_270 (O_270,N_9534,N_9270);
or UO_271 (O_271,N_9794,N_9630);
nand UO_272 (O_272,N_9084,N_9191);
xnor UO_273 (O_273,N_9712,N_9359);
nor UO_274 (O_274,N_9481,N_9536);
and UO_275 (O_275,N_9497,N_9248);
or UO_276 (O_276,N_9118,N_9850);
nand UO_277 (O_277,N_9790,N_9549);
nand UO_278 (O_278,N_9878,N_9413);
nor UO_279 (O_279,N_9406,N_9109);
or UO_280 (O_280,N_9819,N_9956);
and UO_281 (O_281,N_9572,N_9057);
nand UO_282 (O_282,N_9321,N_9772);
nor UO_283 (O_283,N_9012,N_9156);
and UO_284 (O_284,N_9209,N_9876);
or UO_285 (O_285,N_9858,N_9891);
and UO_286 (O_286,N_9323,N_9950);
or UO_287 (O_287,N_9813,N_9817);
or UO_288 (O_288,N_9011,N_9401);
nor UO_289 (O_289,N_9205,N_9030);
or UO_290 (O_290,N_9517,N_9292);
or UO_291 (O_291,N_9901,N_9821);
xor UO_292 (O_292,N_9541,N_9212);
or UO_293 (O_293,N_9425,N_9180);
or UO_294 (O_294,N_9355,N_9076);
nand UO_295 (O_295,N_9162,N_9144);
nor UO_296 (O_296,N_9437,N_9665);
nor UO_297 (O_297,N_9237,N_9210);
nor UO_298 (O_298,N_9054,N_9228);
or UO_299 (O_299,N_9529,N_9407);
or UO_300 (O_300,N_9765,N_9836);
nand UO_301 (O_301,N_9885,N_9379);
nand UO_302 (O_302,N_9252,N_9176);
xnor UO_303 (O_303,N_9083,N_9486);
nand UO_304 (O_304,N_9282,N_9867);
and UO_305 (O_305,N_9903,N_9849);
and UO_306 (O_306,N_9367,N_9826);
or UO_307 (O_307,N_9688,N_9505);
xnor UO_308 (O_308,N_9692,N_9060);
xor UO_309 (O_309,N_9563,N_9954);
nor UO_310 (O_310,N_9081,N_9760);
nand UO_311 (O_311,N_9040,N_9062);
nand UO_312 (O_312,N_9681,N_9986);
and UO_313 (O_313,N_9082,N_9448);
and UO_314 (O_314,N_9389,N_9993);
nor UO_315 (O_315,N_9079,N_9893);
and UO_316 (O_316,N_9944,N_9415);
and UO_317 (O_317,N_9707,N_9691);
or UO_318 (O_318,N_9485,N_9734);
and UO_319 (O_319,N_9208,N_9642);
nand UO_320 (O_320,N_9985,N_9403);
or UO_321 (O_321,N_9510,N_9015);
nand UO_322 (O_322,N_9265,N_9262);
nand UO_323 (O_323,N_9981,N_9663);
xnor UO_324 (O_324,N_9628,N_9457);
xnor UO_325 (O_325,N_9569,N_9222);
nor UO_326 (O_326,N_9348,N_9519);
or UO_327 (O_327,N_9061,N_9046);
and UO_328 (O_328,N_9927,N_9687);
or UO_329 (O_329,N_9412,N_9722);
or UO_330 (O_330,N_9087,N_9242);
nand UO_331 (O_331,N_9296,N_9409);
and UO_332 (O_332,N_9511,N_9142);
nand UO_333 (O_333,N_9238,N_9560);
or UO_334 (O_334,N_9587,N_9048);
nor UO_335 (O_335,N_9090,N_9138);
and UO_336 (O_336,N_9443,N_9244);
or UO_337 (O_337,N_9422,N_9740);
nor UO_338 (O_338,N_9689,N_9402);
and UO_339 (O_339,N_9487,N_9983);
or UO_340 (O_340,N_9504,N_9557);
or UO_341 (O_341,N_9114,N_9905);
xnor UO_342 (O_342,N_9446,N_9383);
xor UO_343 (O_343,N_9203,N_9769);
or UO_344 (O_344,N_9143,N_9676);
nor UO_345 (O_345,N_9941,N_9066);
and UO_346 (O_346,N_9253,N_9102);
and UO_347 (O_347,N_9936,N_9668);
xor UO_348 (O_348,N_9924,N_9464);
nand UO_349 (O_349,N_9544,N_9418);
or UO_350 (O_350,N_9860,N_9259);
nand UO_351 (O_351,N_9500,N_9175);
and UO_352 (O_352,N_9135,N_9766);
nand UO_353 (O_353,N_9633,N_9605);
nand UO_354 (O_354,N_9268,N_9442);
nor UO_355 (O_355,N_9757,N_9160);
nand UO_356 (O_356,N_9859,N_9995);
nor UO_357 (O_357,N_9921,N_9746);
nor UO_358 (O_358,N_9814,N_9167);
and UO_359 (O_359,N_9670,N_9664);
nor UO_360 (O_360,N_9338,N_9671);
nor UO_361 (O_361,N_9789,N_9122);
or UO_362 (O_362,N_9128,N_9033);
nand UO_363 (O_363,N_9450,N_9068);
and UO_364 (O_364,N_9263,N_9906);
nand UO_365 (O_365,N_9957,N_9100);
and UO_366 (O_366,N_9372,N_9559);
nor UO_367 (O_367,N_9830,N_9869);
nand UO_368 (O_368,N_9782,N_9571);
and UO_369 (O_369,N_9001,N_9754);
and UO_370 (O_370,N_9006,N_9038);
or UO_371 (O_371,N_9499,N_9710);
nor UO_372 (O_372,N_9247,N_9000);
nor UO_373 (O_373,N_9997,N_9975);
and UO_374 (O_374,N_9816,N_9904);
and UO_375 (O_375,N_9199,N_9226);
nand UO_376 (O_376,N_9578,N_9266);
and UO_377 (O_377,N_9582,N_9847);
nand UO_378 (O_378,N_9197,N_9169);
nor UO_379 (O_379,N_9447,N_9468);
and UO_380 (O_380,N_9697,N_9366);
or UO_381 (O_381,N_9703,N_9136);
nor UO_382 (O_382,N_9345,N_9393);
nor UO_383 (O_383,N_9545,N_9178);
nand UO_384 (O_384,N_9898,N_9098);
nand UO_385 (O_385,N_9796,N_9767);
and UO_386 (O_386,N_9839,N_9940);
nor UO_387 (O_387,N_9159,N_9459);
and UO_388 (O_388,N_9853,N_9783);
and UO_389 (O_389,N_9894,N_9831);
nor UO_390 (O_390,N_9621,N_9880);
nand UO_391 (O_391,N_9214,N_9907);
nor UO_392 (O_392,N_9626,N_9378);
nand UO_393 (O_393,N_9680,N_9522);
nor UO_394 (O_394,N_9112,N_9539);
or UO_395 (O_395,N_9591,N_9669);
and UO_396 (O_396,N_9472,N_9126);
and UO_397 (O_397,N_9608,N_9751);
and UO_398 (O_398,N_9726,N_9225);
or UO_399 (O_399,N_9551,N_9958);
or UO_400 (O_400,N_9235,N_9042);
and UO_401 (O_401,N_9700,N_9815);
nor UO_402 (O_402,N_9911,N_9088);
nor UO_403 (O_403,N_9284,N_9781);
or UO_404 (O_404,N_9651,N_9810);
nand UO_405 (O_405,N_9588,N_9537);
nand UO_406 (O_406,N_9396,N_9987);
or UO_407 (O_407,N_9324,N_9319);
or UO_408 (O_408,N_9953,N_9316);
nor UO_409 (O_409,N_9377,N_9596);
or UO_410 (O_410,N_9991,N_9937);
and UO_411 (O_411,N_9445,N_9925);
and UO_412 (O_412,N_9340,N_9116);
nand UO_413 (O_413,N_9716,N_9922);
or UO_414 (O_414,N_9711,N_9200);
xor UO_415 (O_415,N_9280,N_9182);
nand UO_416 (O_416,N_9657,N_9080);
xnor UO_417 (O_417,N_9743,N_9604);
or UO_418 (O_418,N_9024,N_9386);
and UO_419 (O_419,N_9429,N_9017);
nand UO_420 (O_420,N_9698,N_9330);
or UO_421 (O_421,N_9326,N_9051);
nand UO_422 (O_422,N_9718,N_9490);
nor UO_423 (O_423,N_9609,N_9624);
nor UO_424 (O_424,N_9802,N_9938);
xnor UO_425 (O_425,N_9357,N_9236);
or UO_426 (O_426,N_9915,N_9897);
nor UO_427 (O_427,N_9653,N_9652);
and UO_428 (O_428,N_9091,N_9872);
nand UO_429 (O_429,N_9900,N_9577);
xor UO_430 (O_430,N_9104,N_9579);
nor UO_431 (O_431,N_9346,N_9013);
nor UO_432 (O_432,N_9565,N_9918);
xnor UO_433 (O_433,N_9566,N_9074);
nand UO_434 (O_434,N_9844,N_9695);
and UO_435 (O_435,N_9785,N_9198);
nor UO_436 (O_436,N_9306,N_9775);
or UO_437 (O_437,N_9590,N_9969);
nor UO_438 (O_438,N_9822,N_9455);
nor UO_439 (O_439,N_9234,N_9177);
nor UO_440 (O_440,N_9430,N_9841);
or UO_441 (O_441,N_9933,N_9646);
nand UO_442 (O_442,N_9795,N_9045);
nor UO_443 (O_443,N_9036,N_9245);
xor UO_444 (O_444,N_9035,N_9342);
nor UO_445 (O_445,N_9645,N_9201);
and UO_446 (O_446,N_9131,N_9010);
nand UO_447 (O_447,N_9724,N_9799);
xor UO_448 (O_448,N_9977,N_9976);
and UO_449 (O_449,N_9623,N_9189);
xnor UO_450 (O_450,N_9239,N_9341);
or UO_451 (O_451,N_9833,N_9217);
or UO_452 (O_452,N_9301,N_9771);
and UO_453 (O_453,N_9870,N_9801);
or UO_454 (O_454,N_9832,N_9947);
nand UO_455 (O_455,N_9304,N_9289);
nor UO_456 (O_456,N_9684,N_9456);
nor UO_457 (O_457,N_9295,N_9966);
xnor UO_458 (O_458,N_9532,N_9636);
or UO_459 (O_459,N_9417,N_9530);
and UO_460 (O_460,N_9738,N_9996);
nand UO_461 (O_461,N_9119,N_9527);
or UO_462 (O_462,N_9125,N_9946);
nor UO_463 (O_463,N_9971,N_9573);
and UO_464 (O_464,N_9211,N_9433);
nand UO_465 (O_465,N_9311,N_9644);
nor UO_466 (O_466,N_9085,N_9686);
nor UO_467 (O_467,N_9086,N_9861);
nand UO_468 (O_468,N_9948,N_9538);
or UO_469 (O_469,N_9385,N_9862);
or UO_470 (O_470,N_9094,N_9095);
nor UO_471 (O_471,N_9567,N_9603);
or UO_472 (O_472,N_9584,N_9240);
nor UO_473 (O_473,N_9172,N_9553);
nor UO_474 (O_474,N_9914,N_9416);
and UO_475 (O_475,N_9717,N_9267);
and UO_476 (O_476,N_9388,N_9277);
and UO_477 (O_477,N_9702,N_9309);
nand UO_478 (O_478,N_9672,N_9592);
nor UO_479 (O_479,N_9113,N_9597);
or UO_480 (O_480,N_9639,N_9067);
and UO_481 (O_481,N_9465,N_9154);
nor UO_482 (O_482,N_9123,N_9600);
nor UO_483 (O_483,N_9351,N_9339);
or UO_484 (O_484,N_9471,N_9845);
nor UO_485 (O_485,N_9791,N_9108);
and UO_486 (O_486,N_9881,N_9601);
and UO_487 (O_487,N_9980,N_9183);
xnor UO_488 (O_488,N_9792,N_9441);
nand UO_489 (O_489,N_9041,N_9390);
xnor UO_490 (O_490,N_9285,N_9371);
and UO_491 (O_491,N_9229,N_9973);
nand UO_492 (O_492,N_9622,N_9246);
or UO_493 (O_493,N_9325,N_9920);
nor UO_494 (O_494,N_9884,N_9705);
and UO_495 (O_495,N_9542,N_9147);
nor UO_496 (O_496,N_9752,N_9896);
nand UO_497 (O_497,N_9254,N_9820);
and UO_498 (O_498,N_9951,N_9595);
or UO_499 (O_499,N_9643,N_9463);
and UO_500 (O_500,N_9180,N_9102);
nand UO_501 (O_501,N_9158,N_9369);
nor UO_502 (O_502,N_9844,N_9525);
nand UO_503 (O_503,N_9718,N_9239);
or UO_504 (O_504,N_9059,N_9470);
and UO_505 (O_505,N_9524,N_9821);
and UO_506 (O_506,N_9683,N_9876);
and UO_507 (O_507,N_9681,N_9300);
and UO_508 (O_508,N_9710,N_9790);
and UO_509 (O_509,N_9723,N_9081);
and UO_510 (O_510,N_9764,N_9542);
and UO_511 (O_511,N_9957,N_9618);
xnor UO_512 (O_512,N_9006,N_9870);
and UO_513 (O_513,N_9146,N_9644);
nor UO_514 (O_514,N_9620,N_9143);
or UO_515 (O_515,N_9978,N_9755);
or UO_516 (O_516,N_9702,N_9679);
and UO_517 (O_517,N_9691,N_9851);
and UO_518 (O_518,N_9982,N_9892);
nand UO_519 (O_519,N_9796,N_9854);
or UO_520 (O_520,N_9038,N_9690);
nand UO_521 (O_521,N_9877,N_9302);
nand UO_522 (O_522,N_9992,N_9818);
and UO_523 (O_523,N_9461,N_9012);
nand UO_524 (O_524,N_9959,N_9831);
and UO_525 (O_525,N_9494,N_9977);
nand UO_526 (O_526,N_9980,N_9751);
or UO_527 (O_527,N_9279,N_9571);
nand UO_528 (O_528,N_9102,N_9309);
and UO_529 (O_529,N_9752,N_9002);
nand UO_530 (O_530,N_9613,N_9148);
nor UO_531 (O_531,N_9540,N_9100);
and UO_532 (O_532,N_9341,N_9048);
or UO_533 (O_533,N_9086,N_9636);
nand UO_534 (O_534,N_9651,N_9266);
nor UO_535 (O_535,N_9049,N_9199);
or UO_536 (O_536,N_9900,N_9277);
xor UO_537 (O_537,N_9517,N_9793);
and UO_538 (O_538,N_9467,N_9244);
nor UO_539 (O_539,N_9690,N_9744);
or UO_540 (O_540,N_9298,N_9023);
or UO_541 (O_541,N_9242,N_9967);
and UO_542 (O_542,N_9248,N_9178);
nand UO_543 (O_543,N_9835,N_9303);
nor UO_544 (O_544,N_9061,N_9995);
and UO_545 (O_545,N_9300,N_9742);
and UO_546 (O_546,N_9693,N_9126);
or UO_547 (O_547,N_9014,N_9978);
nand UO_548 (O_548,N_9644,N_9780);
nand UO_549 (O_549,N_9566,N_9159);
or UO_550 (O_550,N_9042,N_9243);
and UO_551 (O_551,N_9547,N_9771);
xnor UO_552 (O_552,N_9082,N_9953);
or UO_553 (O_553,N_9865,N_9809);
and UO_554 (O_554,N_9964,N_9165);
or UO_555 (O_555,N_9900,N_9541);
or UO_556 (O_556,N_9202,N_9560);
nand UO_557 (O_557,N_9467,N_9022);
and UO_558 (O_558,N_9382,N_9486);
and UO_559 (O_559,N_9090,N_9555);
and UO_560 (O_560,N_9046,N_9414);
nand UO_561 (O_561,N_9512,N_9735);
nand UO_562 (O_562,N_9261,N_9649);
and UO_563 (O_563,N_9951,N_9793);
nand UO_564 (O_564,N_9529,N_9847);
and UO_565 (O_565,N_9348,N_9999);
nand UO_566 (O_566,N_9268,N_9149);
nor UO_567 (O_567,N_9269,N_9245);
xor UO_568 (O_568,N_9381,N_9976);
nand UO_569 (O_569,N_9678,N_9979);
xnor UO_570 (O_570,N_9514,N_9044);
or UO_571 (O_571,N_9074,N_9199);
or UO_572 (O_572,N_9222,N_9322);
nor UO_573 (O_573,N_9229,N_9709);
and UO_574 (O_574,N_9267,N_9410);
and UO_575 (O_575,N_9671,N_9658);
xor UO_576 (O_576,N_9427,N_9439);
xnor UO_577 (O_577,N_9550,N_9037);
or UO_578 (O_578,N_9719,N_9590);
and UO_579 (O_579,N_9249,N_9403);
nand UO_580 (O_580,N_9517,N_9766);
nand UO_581 (O_581,N_9728,N_9922);
or UO_582 (O_582,N_9418,N_9976);
and UO_583 (O_583,N_9556,N_9717);
and UO_584 (O_584,N_9545,N_9630);
and UO_585 (O_585,N_9106,N_9467);
nand UO_586 (O_586,N_9411,N_9896);
nor UO_587 (O_587,N_9417,N_9683);
and UO_588 (O_588,N_9854,N_9275);
xnor UO_589 (O_589,N_9894,N_9670);
nor UO_590 (O_590,N_9730,N_9685);
nand UO_591 (O_591,N_9947,N_9559);
xor UO_592 (O_592,N_9770,N_9080);
or UO_593 (O_593,N_9513,N_9783);
or UO_594 (O_594,N_9730,N_9904);
nand UO_595 (O_595,N_9349,N_9836);
nor UO_596 (O_596,N_9113,N_9799);
nand UO_597 (O_597,N_9688,N_9407);
and UO_598 (O_598,N_9148,N_9968);
nand UO_599 (O_599,N_9334,N_9025);
and UO_600 (O_600,N_9277,N_9481);
or UO_601 (O_601,N_9012,N_9425);
and UO_602 (O_602,N_9860,N_9452);
or UO_603 (O_603,N_9173,N_9614);
nand UO_604 (O_604,N_9986,N_9789);
or UO_605 (O_605,N_9299,N_9005);
and UO_606 (O_606,N_9634,N_9978);
and UO_607 (O_607,N_9191,N_9647);
and UO_608 (O_608,N_9071,N_9737);
or UO_609 (O_609,N_9606,N_9849);
or UO_610 (O_610,N_9450,N_9709);
nor UO_611 (O_611,N_9534,N_9706);
nand UO_612 (O_612,N_9149,N_9161);
and UO_613 (O_613,N_9810,N_9506);
nand UO_614 (O_614,N_9232,N_9342);
and UO_615 (O_615,N_9837,N_9149);
and UO_616 (O_616,N_9814,N_9732);
nor UO_617 (O_617,N_9996,N_9588);
and UO_618 (O_618,N_9975,N_9288);
nor UO_619 (O_619,N_9155,N_9872);
nor UO_620 (O_620,N_9121,N_9163);
or UO_621 (O_621,N_9614,N_9526);
xnor UO_622 (O_622,N_9990,N_9097);
or UO_623 (O_623,N_9609,N_9399);
nand UO_624 (O_624,N_9088,N_9258);
nor UO_625 (O_625,N_9968,N_9686);
xnor UO_626 (O_626,N_9656,N_9398);
and UO_627 (O_627,N_9979,N_9884);
or UO_628 (O_628,N_9059,N_9826);
xnor UO_629 (O_629,N_9687,N_9956);
or UO_630 (O_630,N_9337,N_9862);
nor UO_631 (O_631,N_9253,N_9220);
nor UO_632 (O_632,N_9558,N_9648);
and UO_633 (O_633,N_9981,N_9339);
nand UO_634 (O_634,N_9653,N_9451);
and UO_635 (O_635,N_9251,N_9411);
or UO_636 (O_636,N_9283,N_9418);
or UO_637 (O_637,N_9011,N_9307);
and UO_638 (O_638,N_9568,N_9698);
or UO_639 (O_639,N_9221,N_9956);
and UO_640 (O_640,N_9581,N_9385);
or UO_641 (O_641,N_9265,N_9758);
or UO_642 (O_642,N_9121,N_9495);
and UO_643 (O_643,N_9317,N_9763);
nor UO_644 (O_644,N_9673,N_9182);
and UO_645 (O_645,N_9485,N_9131);
or UO_646 (O_646,N_9993,N_9346);
or UO_647 (O_647,N_9564,N_9673);
or UO_648 (O_648,N_9912,N_9520);
and UO_649 (O_649,N_9855,N_9302);
or UO_650 (O_650,N_9247,N_9225);
or UO_651 (O_651,N_9678,N_9032);
nand UO_652 (O_652,N_9628,N_9303);
nand UO_653 (O_653,N_9129,N_9608);
and UO_654 (O_654,N_9067,N_9277);
nand UO_655 (O_655,N_9050,N_9083);
or UO_656 (O_656,N_9936,N_9869);
nor UO_657 (O_657,N_9304,N_9518);
nand UO_658 (O_658,N_9859,N_9819);
or UO_659 (O_659,N_9283,N_9416);
nand UO_660 (O_660,N_9115,N_9049);
nand UO_661 (O_661,N_9197,N_9906);
and UO_662 (O_662,N_9665,N_9378);
xnor UO_663 (O_663,N_9468,N_9493);
nand UO_664 (O_664,N_9929,N_9140);
xor UO_665 (O_665,N_9309,N_9388);
nor UO_666 (O_666,N_9381,N_9462);
or UO_667 (O_667,N_9113,N_9138);
nor UO_668 (O_668,N_9689,N_9378);
nor UO_669 (O_669,N_9561,N_9717);
or UO_670 (O_670,N_9894,N_9414);
xnor UO_671 (O_671,N_9774,N_9546);
or UO_672 (O_672,N_9206,N_9960);
nor UO_673 (O_673,N_9002,N_9970);
nor UO_674 (O_674,N_9416,N_9545);
nand UO_675 (O_675,N_9723,N_9138);
xor UO_676 (O_676,N_9751,N_9784);
or UO_677 (O_677,N_9008,N_9252);
nor UO_678 (O_678,N_9880,N_9345);
nand UO_679 (O_679,N_9636,N_9540);
nor UO_680 (O_680,N_9749,N_9928);
nor UO_681 (O_681,N_9251,N_9599);
nor UO_682 (O_682,N_9246,N_9198);
nand UO_683 (O_683,N_9212,N_9258);
and UO_684 (O_684,N_9577,N_9115);
or UO_685 (O_685,N_9937,N_9373);
nor UO_686 (O_686,N_9104,N_9834);
nand UO_687 (O_687,N_9436,N_9503);
nand UO_688 (O_688,N_9376,N_9921);
and UO_689 (O_689,N_9652,N_9207);
or UO_690 (O_690,N_9198,N_9206);
and UO_691 (O_691,N_9358,N_9190);
and UO_692 (O_692,N_9329,N_9930);
nand UO_693 (O_693,N_9282,N_9587);
nand UO_694 (O_694,N_9369,N_9065);
nor UO_695 (O_695,N_9790,N_9111);
or UO_696 (O_696,N_9373,N_9181);
nand UO_697 (O_697,N_9872,N_9865);
and UO_698 (O_698,N_9213,N_9126);
nand UO_699 (O_699,N_9758,N_9899);
or UO_700 (O_700,N_9757,N_9897);
and UO_701 (O_701,N_9282,N_9486);
xor UO_702 (O_702,N_9007,N_9103);
and UO_703 (O_703,N_9229,N_9401);
nand UO_704 (O_704,N_9396,N_9174);
xor UO_705 (O_705,N_9236,N_9135);
and UO_706 (O_706,N_9128,N_9655);
nand UO_707 (O_707,N_9146,N_9981);
nand UO_708 (O_708,N_9283,N_9329);
nand UO_709 (O_709,N_9997,N_9959);
xnor UO_710 (O_710,N_9719,N_9310);
nor UO_711 (O_711,N_9545,N_9851);
and UO_712 (O_712,N_9864,N_9464);
or UO_713 (O_713,N_9785,N_9316);
nor UO_714 (O_714,N_9789,N_9592);
nor UO_715 (O_715,N_9766,N_9455);
nor UO_716 (O_716,N_9596,N_9807);
nor UO_717 (O_717,N_9521,N_9082);
xor UO_718 (O_718,N_9987,N_9577);
and UO_719 (O_719,N_9194,N_9465);
nand UO_720 (O_720,N_9997,N_9397);
nand UO_721 (O_721,N_9417,N_9222);
nand UO_722 (O_722,N_9781,N_9525);
or UO_723 (O_723,N_9516,N_9253);
or UO_724 (O_724,N_9546,N_9115);
and UO_725 (O_725,N_9956,N_9138);
xnor UO_726 (O_726,N_9777,N_9877);
or UO_727 (O_727,N_9402,N_9862);
and UO_728 (O_728,N_9153,N_9387);
nand UO_729 (O_729,N_9689,N_9736);
nor UO_730 (O_730,N_9645,N_9926);
nand UO_731 (O_731,N_9847,N_9405);
nor UO_732 (O_732,N_9963,N_9290);
and UO_733 (O_733,N_9503,N_9467);
nand UO_734 (O_734,N_9944,N_9066);
and UO_735 (O_735,N_9245,N_9891);
nand UO_736 (O_736,N_9325,N_9966);
and UO_737 (O_737,N_9645,N_9613);
and UO_738 (O_738,N_9581,N_9351);
nor UO_739 (O_739,N_9519,N_9478);
nand UO_740 (O_740,N_9566,N_9711);
nand UO_741 (O_741,N_9716,N_9519);
or UO_742 (O_742,N_9306,N_9209);
xor UO_743 (O_743,N_9052,N_9846);
and UO_744 (O_744,N_9086,N_9376);
nand UO_745 (O_745,N_9870,N_9606);
nor UO_746 (O_746,N_9170,N_9214);
and UO_747 (O_747,N_9972,N_9328);
and UO_748 (O_748,N_9667,N_9730);
nor UO_749 (O_749,N_9909,N_9324);
nor UO_750 (O_750,N_9214,N_9319);
or UO_751 (O_751,N_9508,N_9166);
nor UO_752 (O_752,N_9987,N_9771);
or UO_753 (O_753,N_9924,N_9946);
or UO_754 (O_754,N_9336,N_9474);
or UO_755 (O_755,N_9116,N_9743);
and UO_756 (O_756,N_9839,N_9229);
nor UO_757 (O_757,N_9174,N_9883);
nand UO_758 (O_758,N_9743,N_9068);
xor UO_759 (O_759,N_9508,N_9955);
nor UO_760 (O_760,N_9275,N_9109);
nor UO_761 (O_761,N_9068,N_9997);
or UO_762 (O_762,N_9620,N_9122);
nand UO_763 (O_763,N_9343,N_9906);
nor UO_764 (O_764,N_9934,N_9017);
nor UO_765 (O_765,N_9661,N_9579);
and UO_766 (O_766,N_9414,N_9193);
and UO_767 (O_767,N_9825,N_9629);
nor UO_768 (O_768,N_9310,N_9073);
or UO_769 (O_769,N_9638,N_9017);
and UO_770 (O_770,N_9988,N_9498);
and UO_771 (O_771,N_9268,N_9816);
xnor UO_772 (O_772,N_9822,N_9354);
nand UO_773 (O_773,N_9499,N_9980);
nor UO_774 (O_774,N_9398,N_9597);
nor UO_775 (O_775,N_9669,N_9596);
nor UO_776 (O_776,N_9541,N_9143);
nor UO_777 (O_777,N_9908,N_9520);
or UO_778 (O_778,N_9677,N_9068);
nand UO_779 (O_779,N_9232,N_9579);
and UO_780 (O_780,N_9756,N_9046);
xnor UO_781 (O_781,N_9085,N_9851);
nand UO_782 (O_782,N_9487,N_9364);
nand UO_783 (O_783,N_9045,N_9581);
nand UO_784 (O_784,N_9163,N_9316);
nor UO_785 (O_785,N_9084,N_9628);
nor UO_786 (O_786,N_9219,N_9901);
nand UO_787 (O_787,N_9325,N_9004);
nor UO_788 (O_788,N_9436,N_9822);
xor UO_789 (O_789,N_9544,N_9837);
or UO_790 (O_790,N_9138,N_9740);
or UO_791 (O_791,N_9111,N_9254);
nand UO_792 (O_792,N_9374,N_9253);
nor UO_793 (O_793,N_9147,N_9403);
nor UO_794 (O_794,N_9732,N_9944);
nand UO_795 (O_795,N_9104,N_9199);
nand UO_796 (O_796,N_9810,N_9162);
nand UO_797 (O_797,N_9349,N_9037);
nand UO_798 (O_798,N_9352,N_9881);
and UO_799 (O_799,N_9265,N_9727);
xor UO_800 (O_800,N_9575,N_9468);
xnor UO_801 (O_801,N_9869,N_9201);
or UO_802 (O_802,N_9844,N_9636);
and UO_803 (O_803,N_9324,N_9344);
nand UO_804 (O_804,N_9703,N_9462);
nand UO_805 (O_805,N_9969,N_9589);
or UO_806 (O_806,N_9347,N_9483);
xor UO_807 (O_807,N_9538,N_9434);
nand UO_808 (O_808,N_9425,N_9262);
and UO_809 (O_809,N_9471,N_9535);
xor UO_810 (O_810,N_9407,N_9427);
or UO_811 (O_811,N_9773,N_9223);
and UO_812 (O_812,N_9709,N_9996);
nand UO_813 (O_813,N_9974,N_9969);
nor UO_814 (O_814,N_9248,N_9010);
xor UO_815 (O_815,N_9551,N_9132);
nor UO_816 (O_816,N_9773,N_9006);
nand UO_817 (O_817,N_9948,N_9935);
nand UO_818 (O_818,N_9327,N_9712);
or UO_819 (O_819,N_9445,N_9652);
nand UO_820 (O_820,N_9774,N_9380);
nand UO_821 (O_821,N_9010,N_9841);
and UO_822 (O_822,N_9158,N_9839);
nor UO_823 (O_823,N_9183,N_9726);
and UO_824 (O_824,N_9665,N_9897);
or UO_825 (O_825,N_9185,N_9519);
nor UO_826 (O_826,N_9976,N_9117);
and UO_827 (O_827,N_9066,N_9627);
nand UO_828 (O_828,N_9265,N_9210);
and UO_829 (O_829,N_9458,N_9087);
nor UO_830 (O_830,N_9084,N_9667);
nor UO_831 (O_831,N_9312,N_9128);
nor UO_832 (O_832,N_9537,N_9246);
or UO_833 (O_833,N_9747,N_9003);
or UO_834 (O_834,N_9528,N_9744);
nor UO_835 (O_835,N_9779,N_9737);
nor UO_836 (O_836,N_9760,N_9841);
nand UO_837 (O_837,N_9109,N_9833);
or UO_838 (O_838,N_9840,N_9333);
xor UO_839 (O_839,N_9850,N_9066);
nor UO_840 (O_840,N_9668,N_9868);
and UO_841 (O_841,N_9537,N_9511);
xnor UO_842 (O_842,N_9109,N_9607);
nand UO_843 (O_843,N_9057,N_9387);
and UO_844 (O_844,N_9501,N_9735);
nor UO_845 (O_845,N_9547,N_9573);
or UO_846 (O_846,N_9603,N_9992);
and UO_847 (O_847,N_9894,N_9594);
and UO_848 (O_848,N_9022,N_9087);
or UO_849 (O_849,N_9802,N_9509);
xor UO_850 (O_850,N_9344,N_9071);
nor UO_851 (O_851,N_9896,N_9026);
or UO_852 (O_852,N_9785,N_9416);
nand UO_853 (O_853,N_9339,N_9669);
nand UO_854 (O_854,N_9264,N_9292);
or UO_855 (O_855,N_9064,N_9868);
xnor UO_856 (O_856,N_9289,N_9305);
nand UO_857 (O_857,N_9770,N_9977);
or UO_858 (O_858,N_9237,N_9923);
or UO_859 (O_859,N_9824,N_9973);
nand UO_860 (O_860,N_9482,N_9422);
and UO_861 (O_861,N_9278,N_9429);
nor UO_862 (O_862,N_9696,N_9455);
or UO_863 (O_863,N_9344,N_9374);
nor UO_864 (O_864,N_9251,N_9930);
nand UO_865 (O_865,N_9613,N_9455);
nor UO_866 (O_866,N_9945,N_9952);
or UO_867 (O_867,N_9233,N_9582);
or UO_868 (O_868,N_9601,N_9981);
nand UO_869 (O_869,N_9897,N_9331);
and UO_870 (O_870,N_9402,N_9544);
and UO_871 (O_871,N_9966,N_9724);
nor UO_872 (O_872,N_9157,N_9124);
xnor UO_873 (O_873,N_9257,N_9568);
nor UO_874 (O_874,N_9497,N_9209);
and UO_875 (O_875,N_9333,N_9684);
and UO_876 (O_876,N_9434,N_9870);
and UO_877 (O_877,N_9710,N_9795);
nor UO_878 (O_878,N_9332,N_9497);
and UO_879 (O_879,N_9344,N_9391);
nand UO_880 (O_880,N_9523,N_9421);
or UO_881 (O_881,N_9356,N_9273);
and UO_882 (O_882,N_9274,N_9432);
nand UO_883 (O_883,N_9244,N_9130);
and UO_884 (O_884,N_9645,N_9265);
or UO_885 (O_885,N_9641,N_9609);
or UO_886 (O_886,N_9053,N_9278);
nor UO_887 (O_887,N_9540,N_9400);
and UO_888 (O_888,N_9703,N_9606);
nand UO_889 (O_889,N_9740,N_9752);
or UO_890 (O_890,N_9054,N_9129);
and UO_891 (O_891,N_9844,N_9617);
nand UO_892 (O_892,N_9142,N_9281);
nand UO_893 (O_893,N_9583,N_9620);
nor UO_894 (O_894,N_9001,N_9375);
nand UO_895 (O_895,N_9167,N_9417);
or UO_896 (O_896,N_9844,N_9985);
or UO_897 (O_897,N_9787,N_9247);
nor UO_898 (O_898,N_9524,N_9411);
or UO_899 (O_899,N_9881,N_9149);
nand UO_900 (O_900,N_9363,N_9627);
nand UO_901 (O_901,N_9159,N_9430);
xnor UO_902 (O_902,N_9285,N_9884);
xor UO_903 (O_903,N_9545,N_9021);
and UO_904 (O_904,N_9858,N_9214);
or UO_905 (O_905,N_9462,N_9794);
nor UO_906 (O_906,N_9978,N_9283);
and UO_907 (O_907,N_9586,N_9961);
and UO_908 (O_908,N_9576,N_9755);
nor UO_909 (O_909,N_9734,N_9230);
nor UO_910 (O_910,N_9030,N_9320);
nand UO_911 (O_911,N_9898,N_9874);
nor UO_912 (O_912,N_9791,N_9700);
and UO_913 (O_913,N_9153,N_9768);
nor UO_914 (O_914,N_9121,N_9207);
or UO_915 (O_915,N_9053,N_9248);
and UO_916 (O_916,N_9363,N_9160);
or UO_917 (O_917,N_9781,N_9346);
nand UO_918 (O_918,N_9047,N_9504);
and UO_919 (O_919,N_9493,N_9044);
nor UO_920 (O_920,N_9451,N_9017);
nand UO_921 (O_921,N_9147,N_9341);
nor UO_922 (O_922,N_9234,N_9865);
nor UO_923 (O_923,N_9629,N_9250);
or UO_924 (O_924,N_9502,N_9163);
and UO_925 (O_925,N_9562,N_9727);
or UO_926 (O_926,N_9754,N_9417);
and UO_927 (O_927,N_9241,N_9529);
nand UO_928 (O_928,N_9130,N_9766);
nor UO_929 (O_929,N_9847,N_9726);
nor UO_930 (O_930,N_9404,N_9476);
nor UO_931 (O_931,N_9965,N_9599);
and UO_932 (O_932,N_9471,N_9624);
nor UO_933 (O_933,N_9982,N_9921);
and UO_934 (O_934,N_9634,N_9723);
or UO_935 (O_935,N_9351,N_9867);
nor UO_936 (O_936,N_9490,N_9805);
nand UO_937 (O_937,N_9500,N_9802);
nand UO_938 (O_938,N_9084,N_9889);
nor UO_939 (O_939,N_9639,N_9072);
nand UO_940 (O_940,N_9237,N_9313);
and UO_941 (O_941,N_9025,N_9784);
nand UO_942 (O_942,N_9992,N_9880);
nor UO_943 (O_943,N_9794,N_9756);
or UO_944 (O_944,N_9874,N_9220);
and UO_945 (O_945,N_9718,N_9700);
and UO_946 (O_946,N_9330,N_9437);
or UO_947 (O_947,N_9130,N_9090);
xnor UO_948 (O_948,N_9540,N_9130);
and UO_949 (O_949,N_9768,N_9511);
and UO_950 (O_950,N_9688,N_9767);
nand UO_951 (O_951,N_9834,N_9965);
and UO_952 (O_952,N_9469,N_9869);
nand UO_953 (O_953,N_9299,N_9535);
or UO_954 (O_954,N_9150,N_9699);
or UO_955 (O_955,N_9897,N_9415);
and UO_956 (O_956,N_9286,N_9758);
nor UO_957 (O_957,N_9876,N_9947);
or UO_958 (O_958,N_9071,N_9235);
or UO_959 (O_959,N_9495,N_9395);
or UO_960 (O_960,N_9093,N_9810);
and UO_961 (O_961,N_9711,N_9119);
nand UO_962 (O_962,N_9071,N_9489);
xor UO_963 (O_963,N_9191,N_9311);
nor UO_964 (O_964,N_9991,N_9360);
nand UO_965 (O_965,N_9576,N_9319);
nand UO_966 (O_966,N_9312,N_9756);
or UO_967 (O_967,N_9435,N_9087);
nor UO_968 (O_968,N_9485,N_9187);
nor UO_969 (O_969,N_9763,N_9417);
and UO_970 (O_970,N_9102,N_9390);
and UO_971 (O_971,N_9122,N_9989);
nor UO_972 (O_972,N_9929,N_9384);
nand UO_973 (O_973,N_9671,N_9278);
and UO_974 (O_974,N_9531,N_9883);
or UO_975 (O_975,N_9583,N_9901);
xnor UO_976 (O_976,N_9926,N_9566);
nand UO_977 (O_977,N_9958,N_9837);
nand UO_978 (O_978,N_9570,N_9135);
nor UO_979 (O_979,N_9447,N_9052);
nor UO_980 (O_980,N_9530,N_9380);
or UO_981 (O_981,N_9605,N_9890);
xor UO_982 (O_982,N_9265,N_9705);
nand UO_983 (O_983,N_9536,N_9752);
xnor UO_984 (O_984,N_9277,N_9831);
and UO_985 (O_985,N_9633,N_9767);
or UO_986 (O_986,N_9977,N_9883);
nand UO_987 (O_987,N_9041,N_9122);
nand UO_988 (O_988,N_9486,N_9362);
nor UO_989 (O_989,N_9395,N_9625);
nand UO_990 (O_990,N_9149,N_9128);
nor UO_991 (O_991,N_9920,N_9018);
nor UO_992 (O_992,N_9113,N_9918);
nor UO_993 (O_993,N_9988,N_9572);
nor UO_994 (O_994,N_9631,N_9389);
or UO_995 (O_995,N_9692,N_9460);
and UO_996 (O_996,N_9284,N_9024);
nand UO_997 (O_997,N_9176,N_9086);
nand UO_998 (O_998,N_9242,N_9561);
or UO_999 (O_999,N_9712,N_9651);
nand UO_1000 (O_1000,N_9072,N_9187);
xnor UO_1001 (O_1001,N_9491,N_9948);
nor UO_1002 (O_1002,N_9544,N_9591);
nand UO_1003 (O_1003,N_9181,N_9028);
nand UO_1004 (O_1004,N_9760,N_9504);
or UO_1005 (O_1005,N_9526,N_9743);
and UO_1006 (O_1006,N_9608,N_9506);
nand UO_1007 (O_1007,N_9702,N_9685);
nand UO_1008 (O_1008,N_9951,N_9083);
or UO_1009 (O_1009,N_9929,N_9499);
nand UO_1010 (O_1010,N_9978,N_9259);
nand UO_1011 (O_1011,N_9294,N_9230);
or UO_1012 (O_1012,N_9038,N_9164);
xor UO_1013 (O_1013,N_9585,N_9418);
xnor UO_1014 (O_1014,N_9428,N_9323);
nor UO_1015 (O_1015,N_9997,N_9802);
or UO_1016 (O_1016,N_9146,N_9101);
nor UO_1017 (O_1017,N_9334,N_9423);
or UO_1018 (O_1018,N_9053,N_9166);
and UO_1019 (O_1019,N_9102,N_9511);
and UO_1020 (O_1020,N_9018,N_9583);
xor UO_1021 (O_1021,N_9066,N_9866);
nor UO_1022 (O_1022,N_9333,N_9008);
or UO_1023 (O_1023,N_9940,N_9920);
and UO_1024 (O_1024,N_9879,N_9414);
xnor UO_1025 (O_1025,N_9423,N_9248);
or UO_1026 (O_1026,N_9868,N_9287);
nor UO_1027 (O_1027,N_9481,N_9202);
and UO_1028 (O_1028,N_9632,N_9685);
nor UO_1029 (O_1029,N_9298,N_9811);
nor UO_1030 (O_1030,N_9634,N_9592);
or UO_1031 (O_1031,N_9485,N_9443);
and UO_1032 (O_1032,N_9628,N_9891);
nor UO_1033 (O_1033,N_9515,N_9015);
or UO_1034 (O_1034,N_9557,N_9742);
or UO_1035 (O_1035,N_9331,N_9711);
and UO_1036 (O_1036,N_9526,N_9261);
and UO_1037 (O_1037,N_9125,N_9620);
or UO_1038 (O_1038,N_9075,N_9316);
or UO_1039 (O_1039,N_9881,N_9469);
nand UO_1040 (O_1040,N_9269,N_9201);
nand UO_1041 (O_1041,N_9113,N_9726);
nand UO_1042 (O_1042,N_9141,N_9780);
or UO_1043 (O_1043,N_9158,N_9643);
nor UO_1044 (O_1044,N_9686,N_9708);
nand UO_1045 (O_1045,N_9357,N_9174);
nor UO_1046 (O_1046,N_9170,N_9694);
and UO_1047 (O_1047,N_9478,N_9278);
nand UO_1048 (O_1048,N_9650,N_9860);
nand UO_1049 (O_1049,N_9651,N_9032);
and UO_1050 (O_1050,N_9842,N_9941);
or UO_1051 (O_1051,N_9771,N_9940);
nor UO_1052 (O_1052,N_9303,N_9159);
or UO_1053 (O_1053,N_9367,N_9757);
xnor UO_1054 (O_1054,N_9965,N_9020);
and UO_1055 (O_1055,N_9475,N_9539);
and UO_1056 (O_1056,N_9480,N_9467);
xnor UO_1057 (O_1057,N_9550,N_9344);
and UO_1058 (O_1058,N_9026,N_9020);
and UO_1059 (O_1059,N_9608,N_9885);
xnor UO_1060 (O_1060,N_9432,N_9161);
xor UO_1061 (O_1061,N_9088,N_9544);
nor UO_1062 (O_1062,N_9307,N_9144);
xnor UO_1063 (O_1063,N_9029,N_9703);
and UO_1064 (O_1064,N_9606,N_9576);
and UO_1065 (O_1065,N_9856,N_9912);
nor UO_1066 (O_1066,N_9444,N_9949);
or UO_1067 (O_1067,N_9108,N_9086);
and UO_1068 (O_1068,N_9958,N_9981);
xnor UO_1069 (O_1069,N_9989,N_9507);
nor UO_1070 (O_1070,N_9834,N_9235);
nor UO_1071 (O_1071,N_9996,N_9626);
or UO_1072 (O_1072,N_9645,N_9933);
or UO_1073 (O_1073,N_9403,N_9808);
xor UO_1074 (O_1074,N_9003,N_9655);
or UO_1075 (O_1075,N_9674,N_9315);
and UO_1076 (O_1076,N_9466,N_9253);
nor UO_1077 (O_1077,N_9815,N_9826);
and UO_1078 (O_1078,N_9108,N_9080);
or UO_1079 (O_1079,N_9136,N_9151);
xnor UO_1080 (O_1080,N_9094,N_9809);
and UO_1081 (O_1081,N_9908,N_9454);
nand UO_1082 (O_1082,N_9332,N_9020);
nand UO_1083 (O_1083,N_9684,N_9511);
and UO_1084 (O_1084,N_9352,N_9032);
or UO_1085 (O_1085,N_9694,N_9387);
and UO_1086 (O_1086,N_9498,N_9938);
and UO_1087 (O_1087,N_9275,N_9571);
and UO_1088 (O_1088,N_9195,N_9728);
and UO_1089 (O_1089,N_9358,N_9079);
and UO_1090 (O_1090,N_9941,N_9245);
nor UO_1091 (O_1091,N_9831,N_9747);
or UO_1092 (O_1092,N_9726,N_9577);
nor UO_1093 (O_1093,N_9782,N_9495);
or UO_1094 (O_1094,N_9806,N_9682);
nand UO_1095 (O_1095,N_9027,N_9802);
and UO_1096 (O_1096,N_9904,N_9010);
xor UO_1097 (O_1097,N_9514,N_9141);
nand UO_1098 (O_1098,N_9478,N_9942);
or UO_1099 (O_1099,N_9561,N_9784);
nor UO_1100 (O_1100,N_9204,N_9742);
and UO_1101 (O_1101,N_9412,N_9422);
nand UO_1102 (O_1102,N_9034,N_9714);
nor UO_1103 (O_1103,N_9502,N_9510);
or UO_1104 (O_1104,N_9190,N_9321);
nand UO_1105 (O_1105,N_9161,N_9197);
and UO_1106 (O_1106,N_9308,N_9938);
and UO_1107 (O_1107,N_9270,N_9048);
xnor UO_1108 (O_1108,N_9697,N_9862);
or UO_1109 (O_1109,N_9584,N_9020);
nor UO_1110 (O_1110,N_9270,N_9262);
and UO_1111 (O_1111,N_9527,N_9921);
or UO_1112 (O_1112,N_9092,N_9687);
nor UO_1113 (O_1113,N_9228,N_9657);
nand UO_1114 (O_1114,N_9416,N_9987);
or UO_1115 (O_1115,N_9128,N_9903);
xnor UO_1116 (O_1116,N_9971,N_9972);
and UO_1117 (O_1117,N_9703,N_9245);
nor UO_1118 (O_1118,N_9093,N_9587);
nor UO_1119 (O_1119,N_9337,N_9889);
nor UO_1120 (O_1120,N_9928,N_9173);
nand UO_1121 (O_1121,N_9849,N_9851);
nor UO_1122 (O_1122,N_9236,N_9044);
nand UO_1123 (O_1123,N_9249,N_9855);
nand UO_1124 (O_1124,N_9540,N_9844);
nand UO_1125 (O_1125,N_9018,N_9880);
and UO_1126 (O_1126,N_9147,N_9935);
or UO_1127 (O_1127,N_9538,N_9853);
nor UO_1128 (O_1128,N_9034,N_9042);
and UO_1129 (O_1129,N_9562,N_9054);
nand UO_1130 (O_1130,N_9635,N_9508);
nand UO_1131 (O_1131,N_9755,N_9990);
nand UO_1132 (O_1132,N_9019,N_9950);
or UO_1133 (O_1133,N_9664,N_9996);
or UO_1134 (O_1134,N_9254,N_9497);
and UO_1135 (O_1135,N_9622,N_9617);
and UO_1136 (O_1136,N_9594,N_9975);
or UO_1137 (O_1137,N_9944,N_9793);
nand UO_1138 (O_1138,N_9055,N_9329);
and UO_1139 (O_1139,N_9460,N_9909);
nor UO_1140 (O_1140,N_9894,N_9918);
nand UO_1141 (O_1141,N_9787,N_9582);
or UO_1142 (O_1142,N_9840,N_9316);
nor UO_1143 (O_1143,N_9545,N_9892);
and UO_1144 (O_1144,N_9050,N_9183);
or UO_1145 (O_1145,N_9476,N_9200);
and UO_1146 (O_1146,N_9219,N_9211);
nor UO_1147 (O_1147,N_9184,N_9140);
nor UO_1148 (O_1148,N_9796,N_9280);
or UO_1149 (O_1149,N_9266,N_9073);
nor UO_1150 (O_1150,N_9234,N_9829);
or UO_1151 (O_1151,N_9064,N_9834);
and UO_1152 (O_1152,N_9682,N_9053);
and UO_1153 (O_1153,N_9038,N_9074);
nand UO_1154 (O_1154,N_9145,N_9666);
and UO_1155 (O_1155,N_9492,N_9644);
xnor UO_1156 (O_1156,N_9120,N_9027);
nor UO_1157 (O_1157,N_9575,N_9355);
nor UO_1158 (O_1158,N_9253,N_9884);
or UO_1159 (O_1159,N_9629,N_9918);
nor UO_1160 (O_1160,N_9753,N_9737);
nor UO_1161 (O_1161,N_9918,N_9739);
nand UO_1162 (O_1162,N_9159,N_9178);
nor UO_1163 (O_1163,N_9299,N_9478);
and UO_1164 (O_1164,N_9730,N_9746);
or UO_1165 (O_1165,N_9214,N_9910);
and UO_1166 (O_1166,N_9368,N_9457);
nor UO_1167 (O_1167,N_9985,N_9826);
or UO_1168 (O_1168,N_9644,N_9245);
and UO_1169 (O_1169,N_9557,N_9649);
or UO_1170 (O_1170,N_9231,N_9050);
or UO_1171 (O_1171,N_9546,N_9238);
and UO_1172 (O_1172,N_9045,N_9405);
nand UO_1173 (O_1173,N_9586,N_9985);
nand UO_1174 (O_1174,N_9529,N_9563);
nand UO_1175 (O_1175,N_9490,N_9858);
nor UO_1176 (O_1176,N_9094,N_9199);
nor UO_1177 (O_1177,N_9184,N_9574);
or UO_1178 (O_1178,N_9624,N_9570);
and UO_1179 (O_1179,N_9881,N_9542);
nand UO_1180 (O_1180,N_9624,N_9851);
nand UO_1181 (O_1181,N_9291,N_9762);
and UO_1182 (O_1182,N_9691,N_9949);
or UO_1183 (O_1183,N_9093,N_9843);
or UO_1184 (O_1184,N_9518,N_9948);
nand UO_1185 (O_1185,N_9855,N_9017);
xnor UO_1186 (O_1186,N_9136,N_9443);
or UO_1187 (O_1187,N_9990,N_9123);
or UO_1188 (O_1188,N_9863,N_9077);
and UO_1189 (O_1189,N_9808,N_9968);
nand UO_1190 (O_1190,N_9336,N_9007);
xor UO_1191 (O_1191,N_9185,N_9842);
xnor UO_1192 (O_1192,N_9768,N_9234);
and UO_1193 (O_1193,N_9370,N_9429);
nand UO_1194 (O_1194,N_9402,N_9239);
nand UO_1195 (O_1195,N_9681,N_9720);
nand UO_1196 (O_1196,N_9092,N_9775);
or UO_1197 (O_1197,N_9896,N_9244);
and UO_1198 (O_1198,N_9723,N_9254);
and UO_1199 (O_1199,N_9987,N_9999);
and UO_1200 (O_1200,N_9178,N_9490);
and UO_1201 (O_1201,N_9053,N_9876);
nand UO_1202 (O_1202,N_9998,N_9279);
and UO_1203 (O_1203,N_9377,N_9927);
nor UO_1204 (O_1204,N_9004,N_9145);
and UO_1205 (O_1205,N_9888,N_9746);
nor UO_1206 (O_1206,N_9743,N_9936);
nand UO_1207 (O_1207,N_9687,N_9439);
nand UO_1208 (O_1208,N_9043,N_9698);
nand UO_1209 (O_1209,N_9785,N_9415);
and UO_1210 (O_1210,N_9078,N_9582);
nand UO_1211 (O_1211,N_9433,N_9863);
xnor UO_1212 (O_1212,N_9885,N_9227);
or UO_1213 (O_1213,N_9150,N_9886);
nor UO_1214 (O_1214,N_9094,N_9273);
and UO_1215 (O_1215,N_9088,N_9409);
or UO_1216 (O_1216,N_9976,N_9610);
nor UO_1217 (O_1217,N_9916,N_9301);
nand UO_1218 (O_1218,N_9583,N_9104);
nand UO_1219 (O_1219,N_9856,N_9415);
nor UO_1220 (O_1220,N_9653,N_9260);
or UO_1221 (O_1221,N_9878,N_9950);
nor UO_1222 (O_1222,N_9541,N_9637);
xnor UO_1223 (O_1223,N_9717,N_9990);
and UO_1224 (O_1224,N_9164,N_9388);
nand UO_1225 (O_1225,N_9293,N_9052);
nor UO_1226 (O_1226,N_9541,N_9996);
nor UO_1227 (O_1227,N_9563,N_9538);
nand UO_1228 (O_1228,N_9936,N_9234);
or UO_1229 (O_1229,N_9076,N_9616);
nand UO_1230 (O_1230,N_9271,N_9006);
and UO_1231 (O_1231,N_9036,N_9244);
nand UO_1232 (O_1232,N_9010,N_9170);
nand UO_1233 (O_1233,N_9870,N_9873);
nand UO_1234 (O_1234,N_9329,N_9979);
and UO_1235 (O_1235,N_9648,N_9863);
and UO_1236 (O_1236,N_9569,N_9681);
and UO_1237 (O_1237,N_9081,N_9407);
and UO_1238 (O_1238,N_9399,N_9490);
nand UO_1239 (O_1239,N_9602,N_9540);
and UO_1240 (O_1240,N_9634,N_9211);
or UO_1241 (O_1241,N_9267,N_9275);
xor UO_1242 (O_1242,N_9529,N_9072);
xor UO_1243 (O_1243,N_9020,N_9075);
or UO_1244 (O_1244,N_9132,N_9765);
nand UO_1245 (O_1245,N_9351,N_9911);
nor UO_1246 (O_1246,N_9524,N_9461);
nand UO_1247 (O_1247,N_9310,N_9262);
nor UO_1248 (O_1248,N_9178,N_9282);
xnor UO_1249 (O_1249,N_9596,N_9440);
and UO_1250 (O_1250,N_9661,N_9498);
and UO_1251 (O_1251,N_9196,N_9828);
nor UO_1252 (O_1252,N_9436,N_9808);
nand UO_1253 (O_1253,N_9881,N_9923);
and UO_1254 (O_1254,N_9531,N_9859);
nand UO_1255 (O_1255,N_9927,N_9133);
nor UO_1256 (O_1256,N_9093,N_9550);
nand UO_1257 (O_1257,N_9899,N_9969);
or UO_1258 (O_1258,N_9888,N_9323);
or UO_1259 (O_1259,N_9650,N_9129);
and UO_1260 (O_1260,N_9875,N_9889);
and UO_1261 (O_1261,N_9599,N_9533);
nand UO_1262 (O_1262,N_9923,N_9308);
xnor UO_1263 (O_1263,N_9674,N_9150);
or UO_1264 (O_1264,N_9331,N_9771);
xor UO_1265 (O_1265,N_9536,N_9092);
and UO_1266 (O_1266,N_9987,N_9509);
xnor UO_1267 (O_1267,N_9843,N_9834);
and UO_1268 (O_1268,N_9589,N_9011);
or UO_1269 (O_1269,N_9485,N_9830);
and UO_1270 (O_1270,N_9152,N_9606);
or UO_1271 (O_1271,N_9960,N_9272);
or UO_1272 (O_1272,N_9692,N_9099);
and UO_1273 (O_1273,N_9030,N_9468);
nand UO_1274 (O_1274,N_9500,N_9626);
nand UO_1275 (O_1275,N_9508,N_9237);
nor UO_1276 (O_1276,N_9850,N_9553);
nand UO_1277 (O_1277,N_9937,N_9105);
nor UO_1278 (O_1278,N_9590,N_9295);
nand UO_1279 (O_1279,N_9017,N_9076);
nand UO_1280 (O_1280,N_9136,N_9727);
or UO_1281 (O_1281,N_9219,N_9911);
nand UO_1282 (O_1282,N_9601,N_9617);
nor UO_1283 (O_1283,N_9666,N_9465);
nor UO_1284 (O_1284,N_9748,N_9909);
or UO_1285 (O_1285,N_9665,N_9598);
nor UO_1286 (O_1286,N_9994,N_9033);
and UO_1287 (O_1287,N_9803,N_9422);
nor UO_1288 (O_1288,N_9142,N_9403);
xnor UO_1289 (O_1289,N_9839,N_9409);
or UO_1290 (O_1290,N_9049,N_9537);
nor UO_1291 (O_1291,N_9255,N_9312);
nor UO_1292 (O_1292,N_9902,N_9248);
nor UO_1293 (O_1293,N_9815,N_9863);
nand UO_1294 (O_1294,N_9408,N_9411);
nand UO_1295 (O_1295,N_9205,N_9533);
or UO_1296 (O_1296,N_9396,N_9989);
xnor UO_1297 (O_1297,N_9561,N_9387);
nand UO_1298 (O_1298,N_9277,N_9582);
nand UO_1299 (O_1299,N_9576,N_9286);
nand UO_1300 (O_1300,N_9645,N_9603);
nor UO_1301 (O_1301,N_9717,N_9858);
xnor UO_1302 (O_1302,N_9589,N_9021);
or UO_1303 (O_1303,N_9740,N_9075);
xor UO_1304 (O_1304,N_9042,N_9321);
nand UO_1305 (O_1305,N_9758,N_9113);
or UO_1306 (O_1306,N_9805,N_9542);
and UO_1307 (O_1307,N_9934,N_9986);
and UO_1308 (O_1308,N_9502,N_9478);
nand UO_1309 (O_1309,N_9031,N_9557);
nand UO_1310 (O_1310,N_9240,N_9916);
and UO_1311 (O_1311,N_9430,N_9383);
or UO_1312 (O_1312,N_9711,N_9913);
or UO_1313 (O_1313,N_9232,N_9956);
nor UO_1314 (O_1314,N_9592,N_9402);
xor UO_1315 (O_1315,N_9085,N_9682);
or UO_1316 (O_1316,N_9144,N_9100);
xnor UO_1317 (O_1317,N_9347,N_9540);
xor UO_1318 (O_1318,N_9472,N_9080);
nor UO_1319 (O_1319,N_9029,N_9180);
nor UO_1320 (O_1320,N_9650,N_9657);
or UO_1321 (O_1321,N_9427,N_9831);
and UO_1322 (O_1322,N_9641,N_9601);
and UO_1323 (O_1323,N_9905,N_9713);
or UO_1324 (O_1324,N_9512,N_9858);
or UO_1325 (O_1325,N_9617,N_9840);
or UO_1326 (O_1326,N_9300,N_9503);
or UO_1327 (O_1327,N_9638,N_9674);
nand UO_1328 (O_1328,N_9148,N_9798);
nor UO_1329 (O_1329,N_9758,N_9739);
nor UO_1330 (O_1330,N_9105,N_9742);
nor UO_1331 (O_1331,N_9222,N_9946);
nor UO_1332 (O_1332,N_9086,N_9014);
and UO_1333 (O_1333,N_9462,N_9214);
or UO_1334 (O_1334,N_9726,N_9904);
nand UO_1335 (O_1335,N_9614,N_9294);
or UO_1336 (O_1336,N_9575,N_9417);
nor UO_1337 (O_1337,N_9612,N_9824);
nor UO_1338 (O_1338,N_9889,N_9998);
and UO_1339 (O_1339,N_9680,N_9394);
or UO_1340 (O_1340,N_9042,N_9576);
xor UO_1341 (O_1341,N_9259,N_9348);
nor UO_1342 (O_1342,N_9391,N_9591);
nor UO_1343 (O_1343,N_9192,N_9558);
and UO_1344 (O_1344,N_9362,N_9829);
or UO_1345 (O_1345,N_9216,N_9326);
or UO_1346 (O_1346,N_9326,N_9981);
nand UO_1347 (O_1347,N_9621,N_9599);
nor UO_1348 (O_1348,N_9491,N_9993);
nor UO_1349 (O_1349,N_9767,N_9250);
nand UO_1350 (O_1350,N_9463,N_9354);
nand UO_1351 (O_1351,N_9453,N_9485);
nand UO_1352 (O_1352,N_9951,N_9261);
nand UO_1353 (O_1353,N_9156,N_9405);
nand UO_1354 (O_1354,N_9128,N_9827);
nor UO_1355 (O_1355,N_9941,N_9256);
or UO_1356 (O_1356,N_9079,N_9689);
nor UO_1357 (O_1357,N_9412,N_9086);
or UO_1358 (O_1358,N_9878,N_9111);
and UO_1359 (O_1359,N_9915,N_9574);
xor UO_1360 (O_1360,N_9363,N_9025);
and UO_1361 (O_1361,N_9027,N_9928);
nor UO_1362 (O_1362,N_9835,N_9923);
or UO_1363 (O_1363,N_9696,N_9470);
nor UO_1364 (O_1364,N_9460,N_9148);
xor UO_1365 (O_1365,N_9006,N_9382);
and UO_1366 (O_1366,N_9894,N_9608);
and UO_1367 (O_1367,N_9611,N_9331);
xnor UO_1368 (O_1368,N_9581,N_9978);
nor UO_1369 (O_1369,N_9763,N_9298);
and UO_1370 (O_1370,N_9714,N_9724);
xnor UO_1371 (O_1371,N_9385,N_9671);
and UO_1372 (O_1372,N_9076,N_9888);
and UO_1373 (O_1373,N_9880,N_9006);
nand UO_1374 (O_1374,N_9865,N_9221);
nor UO_1375 (O_1375,N_9708,N_9073);
and UO_1376 (O_1376,N_9227,N_9934);
or UO_1377 (O_1377,N_9995,N_9808);
or UO_1378 (O_1378,N_9323,N_9761);
or UO_1379 (O_1379,N_9207,N_9722);
xnor UO_1380 (O_1380,N_9095,N_9905);
and UO_1381 (O_1381,N_9792,N_9227);
or UO_1382 (O_1382,N_9546,N_9142);
nand UO_1383 (O_1383,N_9391,N_9499);
or UO_1384 (O_1384,N_9940,N_9259);
and UO_1385 (O_1385,N_9339,N_9952);
nor UO_1386 (O_1386,N_9609,N_9318);
nand UO_1387 (O_1387,N_9045,N_9529);
nor UO_1388 (O_1388,N_9965,N_9440);
and UO_1389 (O_1389,N_9654,N_9755);
nor UO_1390 (O_1390,N_9093,N_9478);
nand UO_1391 (O_1391,N_9795,N_9879);
nand UO_1392 (O_1392,N_9337,N_9404);
nor UO_1393 (O_1393,N_9681,N_9555);
and UO_1394 (O_1394,N_9401,N_9255);
nand UO_1395 (O_1395,N_9827,N_9387);
nand UO_1396 (O_1396,N_9149,N_9980);
or UO_1397 (O_1397,N_9078,N_9549);
and UO_1398 (O_1398,N_9320,N_9552);
and UO_1399 (O_1399,N_9527,N_9058);
nor UO_1400 (O_1400,N_9654,N_9240);
nor UO_1401 (O_1401,N_9045,N_9616);
xnor UO_1402 (O_1402,N_9399,N_9575);
or UO_1403 (O_1403,N_9334,N_9492);
or UO_1404 (O_1404,N_9682,N_9853);
or UO_1405 (O_1405,N_9501,N_9999);
and UO_1406 (O_1406,N_9224,N_9447);
or UO_1407 (O_1407,N_9822,N_9830);
and UO_1408 (O_1408,N_9011,N_9324);
nand UO_1409 (O_1409,N_9740,N_9757);
xnor UO_1410 (O_1410,N_9256,N_9171);
or UO_1411 (O_1411,N_9071,N_9003);
or UO_1412 (O_1412,N_9520,N_9953);
nand UO_1413 (O_1413,N_9756,N_9857);
xor UO_1414 (O_1414,N_9758,N_9090);
and UO_1415 (O_1415,N_9016,N_9248);
nor UO_1416 (O_1416,N_9913,N_9254);
nor UO_1417 (O_1417,N_9279,N_9059);
or UO_1418 (O_1418,N_9648,N_9915);
nand UO_1419 (O_1419,N_9973,N_9799);
and UO_1420 (O_1420,N_9441,N_9748);
nand UO_1421 (O_1421,N_9231,N_9380);
nor UO_1422 (O_1422,N_9238,N_9435);
and UO_1423 (O_1423,N_9890,N_9396);
or UO_1424 (O_1424,N_9551,N_9634);
nand UO_1425 (O_1425,N_9700,N_9030);
nand UO_1426 (O_1426,N_9701,N_9534);
nor UO_1427 (O_1427,N_9017,N_9350);
and UO_1428 (O_1428,N_9863,N_9851);
xor UO_1429 (O_1429,N_9529,N_9838);
nor UO_1430 (O_1430,N_9410,N_9964);
and UO_1431 (O_1431,N_9548,N_9922);
nor UO_1432 (O_1432,N_9685,N_9938);
or UO_1433 (O_1433,N_9558,N_9520);
or UO_1434 (O_1434,N_9636,N_9148);
and UO_1435 (O_1435,N_9888,N_9675);
nand UO_1436 (O_1436,N_9058,N_9137);
or UO_1437 (O_1437,N_9194,N_9847);
and UO_1438 (O_1438,N_9226,N_9762);
nor UO_1439 (O_1439,N_9988,N_9365);
nand UO_1440 (O_1440,N_9837,N_9762);
nor UO_1441 (O_1441,N_9911,N_9623);
nor UO_1442 (O_1442,N_9592,N_9351);
nor UO_1443 (O_1443,N_9968,N_9893);
nor UO_1444 (O_1444,N_9175,N_9828);
nand UO_1445 (O_1445,N_9390,N_9538);
nand UO_1446 (O_1446,N_9727,N_9086);
and UO_1447 (O_1447,N_9523,N_9267);
or UO_1448 (O_1448,N_9576,N_9990);
or UO_1449 (O_1449,N_9747,N_9975);
or UO_1450 (O_1450,N_9320,N_9322);
xnor UO_1451 (O_1451,N_9574,N_9650);
nand UO_1452 (O_1452,N_9033,N_9514);
xor UO_1453 (O_1453,N_9504,N_9245);
nand UO_1454 (O_1454,N_9596,N_9066);
nor UO_1455 (O_1455,N_9633,N_9320);
nand UO_1456 (O_1456,N_9926,N_9876);
xnor UO_1457 (O_1457,N_9204,N_9233);
or UO_1458 (O_1458,N_9449,N_9058);
nand UO_1459 (O_1459,N_9148,N_9540);
and UO_1460 (O_1460,N_9108,N_9912);
nand UO_1461 (O_1461,N_9293,N_9710);
nor UO_1462 (O_1462,N_9535,N_9870);
nor UO_1463 (O_1463,N_9266,N_9118);
xnor UO_1464 (O_1464,N_9835,N_9033);
and UO_1465 (O_1465,N_9390,N_9939);
xnor UO_1466 (O_1466,N_9041,N_9233);
and UO_1467 (O_1467,N_9351,N_9997);
or UO_1468 (O_1468,N_9699,N_9116);
or UO_1469 (O_1469,N_9756,N_9865);
or UO_1470 (O_1470,N_9143,N_9970);
xor UO_1471 (O_1471,N_9145,N_9544);
or UO_1472 (O_1472,N_9584,N_9318);
and UO_1473 (O_1473,N_9542,N_9535);
nor UO_1474 (O_1474,N_9373,N_9591);
or UO_1475 (O_1475,N_9980,N_9577);
or UO_1476 (O_1476,N_9020,N_9036);
or UO_1477 (O_1477,N_9101,N_9089);
or UO_1478 (O_1478,N_9293,N_9384);
nor UO_1479 (O_1479,N_9786,N_9599);
or UO_1480 (O_1480,N_9619,N_9695);
or UO_1481 (O_1481,N_9417,N_9676);
or UO_1482 (O_1482,N_9436,N_9012);
nand UO_1483 (O_1483,N_9202,N_9612);
nand UO_1484 (O_1484,N_9405,N_9861);
nand UO_1485 (O_1485,N_9403,N_9934);
and UO_1486 (O_1486,N_9107,N_9225);
and UO_1487 (O_1487,N_9937,N_9716);
and UO_1488 (O_1488,N_9783,N_9294);
xnor UO_1489 (O_1489,N_9203,N_9156);
or UO_1490 (O_1490,N_9380,N_9261);
nor UO_1491 (O_1491,N_9274,N_9416);
or UO_1492 (O_1492,N_9364,N_9486);
or UO_1493 (O_1493,N_9193,N_9310);
or UO_1494 (O_1494,N_9069,N_9937);
nor UO_1495 (O_1495,N_9830,N_9848);
and UO_1496 (O_1496,N_9602,N_9906);
nor UO_1497 (O_1497,N_9524,N_9968);
and UO_1498 (O_1498,N_9450,N_9476);
nor UO_1499 (O_1499,N_9268,N_9100);
endmodule